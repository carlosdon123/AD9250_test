// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:20 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mQHrSsKXcAaikwLmzAxI/44s+bgsjcUOoQtRu1Ddz/bPHuSwTbCH6GrPqEgvy5Tb
CICnvfwoLsYkkYgQjsWWLSmJEP5qmUiL2d87Pbqs40fwh80JhvPgT5wcCbNa5jBE
hwXw8aCY6GbY6K3NCpUW6b5RN3VsAtUjockA9D8PR94=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36832)
ABrhg+Crjw+namycmn5Z/pweBAam50F2ghLxV7spSMtiSDCqV+EwZJ/MFGRbvvYI
uWAK6W5N2r0y6Zts+CSPdLJiOlK7o+b0bEPjShBnwkUlvdHa/AJ+rJEGCdsxYS61
kc0U17KEJ/OxljE+O3xYsyNsZ76+id8mxV49RxTIjY0gmvBy1BKFxDaxkwvijYDP
k9VjqzmxvJ4VIgh5EMlfSWms3dVE0J5nlL0tuAOFFaAVNRzk/wTHSylBBfCOQizl
P3ZUcCN67N7oC/Uwn8OtpFEay/266V/Zay3lgRJzT72pB1qCzQrvRtVmQ/NPW23d
gKUx95W7QarwrS3acjpvCM8MBiJM2lfNX0jG3V8uC4QBo8tJ22C5F9MW5iM3HY36
U3xVz5/HdNtYkY1bCCEu584Hqmf384KUlmjprkR86fTQSR+EK3LCOvbc+23qV1Z3
sVjv/aoGbr+ZTriRld7CSUHvnaHfyIMofpP/NeChjOnmx/HgrBdvCmEDTNxIjuae
sSNjCh1ukrMk8zfjFaPjfnocanpmsSN0Yp4SUiP/SkpZxh0VvrcDyg17DDBMKJWN
oNve/abyGxETMC+fgTojq1cZacY8oXJPFh5NkxeL4iHFs6lieucbgQw5kUdbtlq2
0+vrwbxJFkl929kDxS18/oCbQFElm/BWcLt2bHA9WpEJZg/wl7pBLs8Rmt2eCa2v
lbi2Ij2eKlU/7IXGu/iaWKgYI962xTNAGFpT3rBGVU3E3rh8DYF1G1as6wX//iYn
+Y0z5LmNzJpCKA9Tk6SGhX8eSouyyUw8+IKkq2aGWod979fE1b4OdRzDD1BdNOfM
/C65qvk+I5kgllZjq51XQIt3I10FfLVZeCXLfWdXcK/vNg89EUm1M3ASB1Il4+/a
Y0mXw4q4hJozgLoCl0Fy5SBSk0IVPh17JUW91OEcapgBKdyhKCQdMtl2GpaXZOiG
8T+87ujaPND/D+OCFfcoFIFC29ljIeg1Y0scRDfnmWtRwAmosaYyKqHiaoCpR2F7
oN1HJMcGuVty7A4Y7cYwnWZCuwI+UVW6yvlCFRa4MuS6OKxRIC0jSU1XkjC6ekN6
YgdvsmCS0BJFPAOyAk1P0NcvKM/Rio9eZSpolT++cqEDFGw3AgkFa75kW0QqEhcQ
LCccr2IjxQ1q7yx05ArhbDH3EcJDd7qf4cEtXz0nfdz68+ikJ0m0cqgynVxvHJIL
K1nBsjhRgqp5N7hxa1UHzkHezDZvbWTU0a0Y7lwKxjucaXkMoEQ8Eu/b3gx8z4aP
5IPHj2ryDEnyzPShxnh1LMfMU+LBGgOPRlEh42hL8GGr6FuvgO7V0XSk60dV2pPX
pCxH5rD/+G0Po14KImX+7pPaXKZ/hGC7rygh1f974BUstyXeLJ/dc6HG/Qhq+0lO
VIjX4+A7ftEM4DFvvgor89S3B4aVJfk3VYN0qPEUD3nggZqKNTy5vUyqvCXXu2iK
BMeKjK51yZQ1Q2GhfcHL+kbHwE+Qqzh6h6VeBE7DKt5MatKJLT7YFoKi9PtFJolk
7lnw6R68PB381/qv5gaPo+EcvOezAdPxI+JALP27whDsuuU7zE0QYXU931Ws/PNY
0ZDCPeWPcy2g5og4RHTp9aqJID6LXHXJahFjJ47/qV3ATBY8k0FKQm9c0CRd9u1z
ui502ZUeuLnatO99HZWIdjZos2m/QTSGPiQX6i2MqP6N8/xQrqTvR8wOI3QqFFd4
sdbwUdAs74mXPWCCGH6oiRnTaCE4kK45GMSMOyUvaVO7b9wMf4ab7cfGoqaQ2jBo
8/cFDJuecgQndj7iLXttFB1pTu8v4tHbS4DVQP80ULA29vVBUwFBiMcYaj+SYvGJ
ZmDXHJK4CqMulhZ8W+UjHdaMsZhxJkElRNxwDkhAAoONcvC48NnOwfErcgr0GDKl
gND/imIvBJL2fj9PfywgU9GsB2zXKptCza6r1DUCD7SSSBfvv/b3Sn6J2EGf75V6
KfzCi9P4QQ0WXnThAYpWKqGP/iYwTTEHAsmCRKvK9unYQMWtZ2lOG+WYZ68S8U90
jQIS9XloVT8i2UZS/3/fJ9YWOjNPA9nhj+6edrRGlg9df8P7JIUThQTBCjsG48Dv
YboDRghKGohZcHT1Cl1gAM3Wqfk7+eu2BMSlH4LM1NBj9RjZpo242V+BxK39y+f+
5bszYlI9yC+cSPKmbXGEukMm3MF/f0cEcJRqm5CFJPtGg6bVSJOcnXNneT/1h1rz
if15B8lJjAZYii4CpSefReuWSQk0TelcJe6vZHAcqJjhjd5ax1UkixZaoHjpkh3D
117nzAEze1Jg1wXskEHOiGhRV9WYPjsCmIMwDRul/WJWytTpJYnnP9g5X+7rJNz7
ojzzEdCqTPfNIMKDNZGxFEdMdzpmBreLObCxu3zO2fsiPMyUvfgivbyaqJmnmd6V
MgvfrBV96q1npfHs1LZFFKfVPIKP4xC6w9wKa3qJe0mjxXOwVEV51BumuBAHckkI
iO+XlK5XQQpk4CcFnpewOkxWA80aOqSphrtw9pFqvyz116M37+qT5jZJu4eHTWac
iajXXssS1usnK8+Q6neqKTMD9fvXGhY71fSm6/jjtcqq9P9FbRhgbOVzkBX8+5zp
BCcVxh4W4Kq3JK+2QQq4YEK2s+UKgFR4NveNHeoVLsrTlGGebk6k/hbSTdxTtYBm
2SmNZ2WWtH0DGN774QV/d9aL0D6tKxxafI0LvIZzCx5TEif2AJykOSaGFpVozUbc
C7sO0M3Uo5NdMp0vFV8Y91TVIkgAm33+9J8N1dPd1rwdlZDQXS/Utt1xhG88T/WI
e60eYCp5vWbc7rqjRLQ+tSx2tJymJzixVaQH4zefjwPdDhTRaRJGkHK/99e896X7
EfqZFMiybjZ0f98c+yQHLB4l5WwRsmJtU8hNyHhIlJuypxPXDvGNW4Xo0zNET+/j
2fJQFmlTXfxe/z+waKNaS16RhqUya26SecNr8KdE2K5h1p1R+FktCsltP7h6wPSo
pEymefcGzEJkhvoBt7h2i52a2wrPI4kL5iHW2PJ4oNULZv25Ec7tyy9piG+uMYGI
ijdQBZYEK9OrWexyEXMpqC3xpPb6Nu4dr1h2flpzRMbWu2u2f7ZTZHOSBjMHxNeJ
MrOWMt9Ug6FMErZlKlETEQ7kZ5EeKqrNVfg+hCexDcwNnF9+JAOC6SkayTdDFIh2
+TpDHW8vzDoMQZyFGw2p8NoxgOjr/5ZfvFryp7WaQT1DgIRhKsVQtEbja7ryx84H
9WFicyAca3H1/HTc/IKjQ68BNbSKdKVC7o62RQpX/TkbAogCG0Sykcwusk1PUXiE
G2X3rAxif4IZgLxv+xsunL32fC5/zfPJDuI9U0DHxnNK0spF7iCK25KnLuJQbafJ
HETXVlZEym90b413vztPAgrkdXVmyLvQH/4H58v0uxYIoCLwFV/E90RBfg3pvWn6
bdoyrR/LqXegRdK4OpTgXOr0cp/6zikMEuIgO/2Ef64ZbfvXt2vnXPcUrGuT94z/
sRgfFpqFXxzapdLNucO6AFOZn80kw2dAxw1Deqohw8hA6QdzePBztbFDA1//8IGd
wTFabiFLQKiVkW0f6EFa6P3gl2Jc3Nl+QOoeJU6an8rMh+AFHXeJtIoHSAs2h//C
sOgJvxCiknsTh7iBZSt3b4i4gfG1SY7PO1zqSavUosEDNhVbLnH7jYjdLROcxgcA
bNfGiU4as1bUxAhbC2ooik9nFnC5Q5mdQDHGLDLZRXIrLpTVY2OqEwc0aBvsBHOs
2SVNwt5QAuG7wEB1B8Pe+QkzSVfa7J5vpG/HkQ4NmVmbVTY4gDWYYfBgKZ3PrqYU
knd0+Oa3B9LJjCIMaxFIDaoZqwvwdhDxxgtAsgg79iCD/9kqf/DGkXu6S3ZWndja
Saf8cudD6FlyvpufXqAlIFYrep0JmCaZj+e+WYtoYt0tGIHmi+mrthK0DLzy2d7a
Ld5AdbtfOy+axgbb4+ItrQN/iT+uuwwY5Q9itpKn2lgCJljBLcM6QcunAOqWegu9
fE3Ijm19njtP8gRJMomSESLhhPUqn1ISftV2uiBS9KI9rDGL2JA72OjgMunW1EWb
peDcitz/DqNOiMre76Wvkcdo75KlFP67savg0HF2MDQMWD67gxHAcjCNVkmlKq+3
reqiMEQRjpV2cf6KcikWid4VAyrdLkt3fBuc4CcpAzbZCDa45RKz2pheFnoz+Awd
O3DPP0teHQlFG/h5MD/q3VZqpKd2KO4HDhEi8RFriDgeHHqN8pvWvTZuzIfQ7eZk
VTMM4GxQ7RnSwuZV6iHguq6uXlxdsLAxdp1Ayjm4a4e2ybxFMt69+IYn4O31aVAf
m6koiuRWsDK1myP5QdLToNUH70moU0I3NXH9kljA/z7Vru9eei/YxPao/F3c+RK4
zBhmu6I893TguSWlueUAupFtTJEn/Jr17sdotcI4rBRc7PHTaadbYxP0bjNX4H7C
mDpb8ZoThfAIrwlpCyXOAyu4VptPyE5BWcLjYnNDvAE9035sIQTwBZ2v2N34ZAQB
WGLgtw8i7HQVaoJFIqWn2RUsa0I31NTzY173HHaYX53zPm8jSNPlk5j2nJjZ01dq
M3qa3KqXL2rYvlsuvz0gykwPlKQfm6hif5oTPUK3iJmrUk5xMhWowoeAAWfbzxk0
bCIPy1Q9T56MeKY6DENUkN1P/LhlCk+/RqUY/wsD+i7rBLVZae1pAx5BYD9Yceir
xVgJz0ij+jrJHkHEm5QfBbP5bMekDENGQ/qsR6wC4YlslW1vYmUg5YoHU8QZm653
clEgbqOaXee0/7paleQtWh3XJU1AD9ZT9NMRkWzRToy2GGdaDFviqKfcb+8bLnvX
vd/na+3o3crxf6RQM/27p/8RgwvbeE6UfFM+sAwp/vERQxYO5Ma5CqmgEE2BYMaa
8nK/e8Idj+aXX+SQXfsBupmlCyT68O77mHrTg2qMPJySZZBgaYTqph1B7/q5Uj6G
Ffw2f695OZDT1Fx/tiZtQxfgwWJ/rHZ3OkNlNXbKYhvmsULJQn+hGKJEBQ03nRni
LQrjhpZEFV/uHzjMsHRLeQGBc7dPh6Ob2mW4i0CwYbhln7Iex7K82JFqnPZUMdKP
70j7ytI7g9ZXio7uQwRIsPR8zOQ564ju6y6fDWJeWTxEVtA1x2w5cjlru2RiewLw
0jEv/GF/qpl+3MwwCpetWW2Hvaxvti4krS7U1TDrM62uZ5AnKp6VB306voN14cay
XYIjkNKhYVU+omSWRVe9JmMIKnxJqYMrTEgcuizswCWLQ0fGCF58kbL+C6hQPok2
vhWCzpiXtnnSNdRFzMNlxsekjWHA0f6eURObvdgKJ0INlfHDkPE6xlipBW4tUMt8
veCKNQtVqJyTLJOe5/LTTbuWRk/vLcr+AbmINO7lK/doAQtms3IPWSgNHrLZY6KI
pZ47LCp+oMV3WPkuAfh4BPRxiCTXkHpa8uRBXkd2Cgq2/NSVGxi941pcsgQW038Z
IF/s/gy4oX0KeoQLdfHl4IG0clbcgi8yU4bSEZ/cOeCoNmcCAncEre9bd6IPkJML
nu6R5NeFCXCDIGkVQmP4uUIuaGzSRBm1N4CASGy7nMKKBJemOAWPMrFd/cxkyK0N
xKX3hqUlHeXVEczTlu/nzrn1Xhh1EWOrCeNWIE81jJQzdzBfqlsm7ArbJaMVwCBO
3YYTiQiCuCcgEzN7hHWjCWRbDiJPX45JUomSP2FXrE3YXS0wpXAUq91uV7B6z0+V
E2Dsc+JWSHsikdhnAktuYXAO7UXlXbe+vmRjn/Zt0Dx3pYlBjRxssELknXXDh5Ot
fYQ3K4aLxP0l6QP4m/IiCfeQ9I3UrKLNX0+d2gCYH9oDAo0ammOry5oNVnCQxx4A
9kXA9ZTyclr7ynFufealNvDmAK5PEqkLEuTzR5g6Dg9SzQmcfrG/6lg8p/bA1cMf
SbOP3noA0VHbImF8nRPsU4fxxCOX75nB0DuTbPX5f4J+av0EJfnuAqEHN2W8lhSV
hSkbuyAUlsV2EQb/rwDgak5xcA0tGFgSUDnUC6MZtpYVg/eUqnG10sEnHXtsWF9H
s4fDtMbh4FPw4QuwEz3Vcp+/00/nBmV2xONG3GTwknQYUEtwJqzm0yium6s4ZgS7
N8Ou7XPD9ORrSlK4w2zptZGjF3efUb/XuI3wuJqYZCEK1sTTip6sCq6BylYx+zXx
lTycMsw9UnEfdEc8gXNQ3p3LrEYEq6yvmy4vLuVzVjjaPoKn5qm/p0KB6ODSD44G
phv04MOEp7scKt29WG0eSFNpbxyJ2iQARhxQFm+kiXr18kguACa0kZRHRC/mIQSi
19EYWTRZWL53bJenIuhml+BszbR+QdxrF2MgJy5huf45gsSfb+zNNaYL4dzyz7f+
ay1FNKpxcAhO4N5X2vQTSZ6xJV5t6GojktZ1t/FZc0CYkMAlZ3FLZKKsbvswd4Yk
kTEz53V8PwVhJSGiVB/SQM3lWylIZf2FBrvj9htFzWEhyO96YQW+o4H9oQQjd1zA
zmeWGVly9QOAveAD83Vw1q/ZC0RV4l6eIoFSikSe9SX3O4A36V/0W5sfmTz4oeF9
JEW+M5cLtJ+7vpLHLQE29tDmqD9VXRaBOfIIK7lhAxF43BZV6+xrvTAiId+kbbzV
g0X5dVwB0SynVodWnM6cDAWoSQocBv/QnGascBgsiv58B4y2/yb1AsrequYdNf1T
lP3CcbnBzhYpD0Qo52A7Xxa5WlUH7Yh5QlrboWjnCCVxRjRvZIGMjKBLGVKppwN4
OQEiSKIw5yJbbgMg/1VH3pCLXnb/9IlFQ7BBgCD+UyBWFkTWTeu3uRbIYHrHdP0x
2awDuyoF5sWzkySntAbrejVL8wy9GgHQ8Tt8lBVh44jVEKcPoavGlFXJceNmKoQD
ismSytVctyGAuDolaT88O24143JyXE/UyG4QDK6j7jL+LBpZNO7XukdcwY9q1s3y
6H25Hmco9Q9d/bJMWrLN+Bc5O2MgakXX3DAyHsnyzC7JuU9iG0uJwzJarbGibE5n
wS4Hr34dOlxFfsZjSZn0sdoHG7iezwFZ1GdiPnoLXnx4ycAgwbicgfamCWdMYL2N
C8WA5o0UyOMNVsFHo2V+SN6J/6ZiqzOh8oSzb/FKP33i5sZ6cmPb0V2KVE6ZgKfX
Ol0MAKXNy+A0BhtKE3RcmXAjJ9S0UovG9HbNKMStU2Q/cHPvvMqGaTT2MGCDxC9i
/YQbW93wv0fpRst9B7JMvmRysHJhdBcYVCGQKJD+LWRMQ7F9im7nWuD1ojpZo/nw
XwpN7f4RtQQYANLTSWjy33R6CK1aVltkmUVVDVrRRR/q7MYddd8a4i9TWkhYMxFn
ka4qBXd6LlPkBPz7F7AWtjtHd+tIKgI21ehR+XjAtXBLhbW8Rrzx8fVcJFKplPfk
ySzNaY66IQgkUCPTRVzaIuqg2aWPs5BIeDIKuxIJM6W+3l1dwL2X/GcUfcWUYtOi
uNR6FUFV/F7g6MfJtYYnC+v+Iros8IjHqDKxBVbc1I9/j7jho0INTQFKt3DouBGm
lFOpvZ7sRkYzew2Gx00Lk/INT3pl9YbVFUu/uqXs79YK8vfRcVdq/lgLMNCzHfgl
STyxm2x2VP9ISMyQlGGJitS0IwmT54hUQYDOT/q4DFXmMSkRUOcxz7axPnmOAORP
YMUVNZGxlwyzNDZaTFWn9R3fBgXfmdjYz36prwSFFVs8FMAQH1IOdqkN9QTlqoW5
Vpi1mXGwZHBCfSznZAY/tTBSI0nyw3gvm6MlqBngZwUedMhSaSXrsgsMtw4DVk2+
vpV5Opyb1DBlsssEHpLujDr9ZELP5im6K9l7tBocU0GbxGnOLGXyyrvHeRpI4ShB
G8sqWm0i2vW23XgEPIWRi2ULg3QutvViXnv6SZkrs/TzPFOoMuU/aztdk6PQx3zU
oJ5AVh1x1Hn3WsQ1fgCyMhugMe8NxeZgCsRnRYuvArhWlMgCKal8szG3GrxNNihS
tjPBvlS23bdecmgUdJxlea/D90q1bLMR84g1E2+l1bNReNCvsubjEqtcjSDPnOI0
fttumNm7X9usCbNYUs91HiNMFL+L1D043rft3VJ9K/lkJvLqOh+l8LYf1q3HUwqM
ZMrlOlLswUirTuzrld9mHNsqTzXTtWi7CFxO6fCTIuNx4r4BYvzpc4qOyZZuJwgn
popH+sLMs5p5eDfF/1EgKbjx0+0MHa1hJrDYD+pGSWqbOlAII5dNP201HnwuYSx6
9EZARHNfYwAKYAfKgBE4N3jyj7uEgFXdeKRHyZPoGL4eM8gg1ZUlCouBZBjJhuCu
U5y9H84H5K6BgzMoArTu0faBL8jsrNhwJenw/yGjQjgVVO3B7dEj72JcXT9zSLLy
+sNQpZcpGRZ1GRdW+zkh+a8a+/50me6slU/oaCiydWyLiEvSXn+PPYbC/U7Cy0uX
OxqThyh511QBwTpetHNCH/4fxyGjXHXATlRg46/seXwv0a+umNHY963ctTCwSkkV
uk4blxhBr46TYKljGu0vMlGjHvIX+bCG7kM7RG81nGsO6ftVdkRqrWf1HtyxD2Pe
aHWXbsL82WSP/Rp+QQgtKPB/zZ/t6GlLhR1CL4wh5olPHaaV5/90omAhixBX4ixC
vTHVTECCYQkRMKRJYJD3f6fr+He++ipybI4EMt83mM264+I3sx/r71QPazErXu0t
YJ9d66UzSfM6sWs3fwG6vSCghEEH0VK6tWidZOvMAlQG8cv8GdFKkPOIh/gGwRhW
GwbwODbIfIuPD/jvcOr0hWZjm58OZVkJAk6gOZY8iXalgMZgxEKPCO3Dk57QRGfr
dsSU8D/Y5P0s6GEXI7OCJIsMVSt4wfqpaWQrwsyqYEsMzwPh8wo0C34OCzFkrk3C
B/zVMZCAVA0tQaM8zoUnUeKh3+7Bcu8LA4ge+m+WbATF0JVKYnV+t2/jpje/kuVO
QUDwq5hcPeS0ZeQx99cHOSDBpiroau/ZZ4HqG4b+b9ndvKUCv/d5MbT5PChsVo9b
W6dckE30V/hGyCndqTaC2t9bQKs0SS9q4q11n8aiKR2Us17Z7KgOT1MKtkt9K/Vy
1bQytIDDFgXrqHNcYdELsys5VsR0GFqS3rY0NAftgGY9H0VdhNy7b86OKT/DdIoC
1/PZml4NiwgvtHKVTYs/TLL6LwjXEi6fPZ9fXq0AR5soUZcntlLhEan/mbqmObiQ
Ts4bsybMK1BCxrqI5Dwm/4MFd+fl+Lqn5L8KGYCN1yLiBQdZwTmA2jCDEVjTp8cY
lC91t12PGRu5zXNLnAT0LkDwe84+abBeOuKqEVYQcxNDsPxb1TmU16KxI38V3YXO
XCBb3VZddm6Kruuh+oY9Qkn+a1gZzhmUkHYTOCcVuM/GVyy98rDOGlqmb+1VVIww
yZSqK7lMupdSf8qN5Pi7KV6nYACfMnMXUZYtD3ehy+PvCxttyyx4FnNPU9ADG/EC
Z+VhpsBkESAddW5WBjcmCZv2eRyRHBazS2+SMK6xSlicdz5aJWsm+rgHQUjqeqh/
i51DMk/emHVhIKOTioGyr0akPS2/IipMFCeniaKmXcc1eFD3L20jtaoUvSA5nIBE
5T1Yt3u9PuR7o70BLOPmVDPeqOdb73KkCoCVv+9QCLqCtrKJTwUIDct0/BEdpNnY
+Tt2TOT1XJ9dEDG6XQ7uHZjkGB1qfGL6MyPWFXMXTbpJSPbR03aKQUvlfctL0X9G
o2UKQ2uiRzAKZET9h5ElXXJFOoDLY0dt42kSJnrsm39ddh8bWOKYzKCx6WXeeEJ5
LSJy4oT0tI8FxNp7jMP4VC70ocQaaOiwRaWeC7znkd5gjayCpkLicoiLWr+dliP8
FwkSqK1BPGGrcN2KCzFNu3iVeS64dYGtmg0TfcXLjQ5MDtNMJMhMVM+9NiqLjYkw
nYAwopSETJrWHhze7aDVtHoSQ4wLWKQqui+QkIvigYq8OOMsjVpqUa3UkuD9+NB9
RMX4MTieA2rqqiVO7W+W/NHQEsabONCnUWuXwpX0biQzYDKg15U/IsOMPs772Tuh
8bIgoZ9kIHdHcDDDtMD9XzZbd9zVGOrmK6wvlc4f0P2dJvW+7HVWdX4dbSWGHzFj
JRF1OWHhHvZ5Wm2kWBj/fjf5iYp/hZrvHVYvoQyn+utB1FOoscuaDh7cnHu5TYkz
n/alv0ybB2wu+EUZUWTXE8rbMUryqpxyh6c3MHGhE8BoYoWfXvRpW8TiZs0ZtlU8
IdVddffmT6HSCfINIHjCIAhC7HGFwxornNdEQH1q6WIIQ+seFd3JpclwUk3xUH7C
BSQFFpKLaro6Nht5xNGZ/bEaSR1liiAznjsynGul7+EI3PkxRCZsKWrLYIrRKjh/
+4mNWbWPECCahHzwoZCE/NS4iDMAMTIfPYmlPZocXqwrI45RJsCDQgFS6dbUXEIR
c1Wztr9F1buQZZwvs2K9XA5vbd95Fi3AWjBE0do/ZVDjZTxbxjVoX9WcTuJ6ySW5
LAnbVWzJ3Lys22YCAug6K9U6HULf5+JcpMtXPFRcOm7VcgyAWURxs+xKAMtbGsTC
IjRlnNSAPN6GmmkMXvuboHZ36J6RUT5twibtMFetZZlhtR4IFN35ypYy059gBSD0
jhP4IubAhOb6CRR7elHFhNQ5O0RD8GaqqHixakn9IbsUfvA08iFXHD0IbykJTLB4
HINiJ5y9e+9pasrT7KBg54yDl4G+NT39aokt6tTyyMVx5Y48t319SsNqtlf45A58
SA2rgn3FCZIJfYieKfyGrLia4oaacdZrcSNYt2hMVltfixIndyv/i+p7gk2SE7Uo
6jssyl44etlE5Hl4TsMtEX1yEQmCcyElWGvBOKL5K4B1AlBoTKm3wBPqct+nqdZo
z/GrHjy+/9WsqWYONUak97JRi6zPsWl9Z36HQyTcDiuJNaBep1e0dy/rUVSwB3Ys
lsGqX9XuHFpRd7tdeYMY4wmZ+Bifp7UJ9wdqyOA/NgVz+WJcRVu/GsT+BUkrZ4Qp
MqXuk59CcsBAjV4LGF+xZ0cZU2C6bMAF/92UK/B3/UwVPWI5d4mHzk/nFFOtwBTP
vsXdxlTjWHUtjgl6VEBJOoicZ8hRWgt2+F89etF0B6LyIRqVJo+u2wg5AAFJAPhc
Xyx1GaIv4ihm9Hsyb/9l33bxf7qpfkSoOrRwzZxos7V9Qf7Qe96LdEvX02AAn5/f
zpyK35MxO5XVa5Jy+8eCLOA92WB+8K4YoJV/w/Q8xZrAne5gpLpo5g6H86ak/jeT
LtVEOuQo7pHX9UJrhPxq8u0yFQVHdwHfUvdbWh+9oSQacBHS0mSKfOxmAT+bXd4T
trrqv3vvZoKuQTI7tBURTgXdFDjmYNMtsVnW+3TEMganzhaKt6dprrPyVKLGpkM6
qAujUp5vP5nSVNBKFM03i+fiWTobRCHBxodDkEQ7GlRbtil11VhmecDe60MUjwLs
3H26+ET//hQsuMDOYNcEoE7GqGoeT+NUhAJhO1zyn79qd6FuHz/aIwAalL36vpxh
Jj0pIVubaKWoixntD6udeoKDlf33D3+rwCxpBLlQuc58TjCOaiBHyfj9vPltO00t
2P9recOyPZ5c38Lya4COkpvm15cZ7sd3Kh4EvSGlR+gQAabs05164IzBXBODz30O
4rVhzcIMgXvLWmQ6xrddBagg9P4qn/eAdbwUMvf1uV+GGMry0fBF1eXllXkslooH
sgGpIB6Xrq5ONX2jcNDRa431La3CD/6PfjkTYt3qOWSMeJCI895AxLtVuyjq20D/
1hAw3maPTiKXrxV23F1KahxLbgQP/rwtsHBrXPf7ZpRDoh+PbB3NIVv+yijfWkjP
2mEGWWvy0DTcNG8W7XRF1+p4vBlgdfpIup/MO+1JdoR+MMCYsudqrPTg/ZejLW7q
63s4GpGlcynvEntetBr7CaGBIxA20acgU21MmZ5uD1MG8kYzk6s5xa75hyV96XEP
3/DAU/Ad6iSwqJ1okazssJFr4ozumO9wGF9IHHuzrYCHFoV/KiVOj0O6IhcbvbHu
k2QYDjFH2Hqf2uMc5tAmLqoN6m5jIH0Sg3nMuMBGY/WfTIW8/MOjhdWCNNBk+JWU
suJgN0iT6LOQwlem4Ifn0m5w2Ikfya6kZEEYUGgCYi1lPS2saU/nvQCGkDtO49QW
bZF5+5mYNNHeuqbOlQ//T9tS+q09sDgIDtFu7BXkRUWdDGLJ0z+WTZDztDJFpoji
qRylrBrezpIXZL8M+iICnCgIPLDbEKm2Cju+HKA8imWSHNIYoaOIQOKYsrsge6b8
JhJOjVNVhebS67G2c/FomGM5MVIjlFpR9mtloJapiOc4qp4sHxGL+BcRZA7FaJln
QpAh/OerQDjNOiUOuiu2r+1j6fULIJsqHz13nDVrXUe9n9pCQUnsskFFbcia3cc7
NHRMIJT8Ybuvmo/ZiFC9vGCtjMq4UI0Fjgnu4FUuOMQqUdCaK7GJnJ3yka+D54Ty
e6IIjDiJyB9knIBsR/TmXr9qFWWS6IZWeYGwgTTiMn9N40FQzULyRVHm1J3QJl7x
oyCqRvn8nZuczW7Zk+7/tdfDk1+9YgkKG2NyReXn3h57tZMP2zmD6Lvn28H1yXmI
CKlDBjSDa1Ondm4sSiqU7KNMgyWHDoXWcPDebIWJOG9VhVd/gMagQLRBc2eJuXJ6
dMi2jfHk1Dx2aDOFt4whYl4EMduWA6MAUEbnOopGIVyxzJSK/ENpe5D/eiUaSt4N
apAGoIw77Bj08trVUhdAiHfEAw9mgkdYMg4p3KbyOD6vxM5LdY1YEpaCjmP+stNE
4UbZP2Tfoqh3qDNGPHIqpQvLSCfnLczREYe4CaIq17wk8LJqJYXxazYp0uG4qUyl
a3FQjZUXVK0cv4adVNWLoguf6LZGMpI4my39Qxf/nKgUCO6javfBPti8ICnjD3mU
Tj/UobOYo27lOrKTGYouZKa2XS4clIVjAVEgrbaqHmb8sicolNKV/kQmOeHg63dk
V/pYJ75aiHj1XUf63R770VVNtvWp+eYQhPaJrv1upRh1MXVv41I+xy0jbgiE6HXr
z6El8SbrckCiCZviFeH5lLMxy/hZRWdrnB9FUZjQYxncj/aqMj4FODsPZanzzqaa
mCvGckCiiT5pfxppMUJdJ33PNEnXDzy6INZpVWYJwkj55jjKONkUrgU6vc0tWldu
K5lF3AielNWcdUuzzysLSiNbrbdN+uIog0A0hoc3us95Po1EeMMHzhCaJsoWsl4V
ZenUIba+fynHS4uGcqOtW1wsCyBfVpQJLBarYp9FiMzGz4sfBR4XsQIB2nKIeTAA
K7ioppoxulawymnkkx/w847V20pHFLHCiIWHmVOQD79KHhvKPDrUapuASL1BpExE
le0eSd9jA++uItZcm3e5wqnSIDhSrC0mzQX/oBl5g6ecWs9y6VgeE62+Pwoupx1u
lQCwKO1WAR+HKkrfJu+499QsgSariQSl+bmpQHDVBmSD3qSNQ0KT9SY4S5marnox
K88hX56SGH09NBR7actKW2u5GFenGKtiDP9Z/S6CUI2HnytTQrMSChaqdPX+Fyxw
mIAn6aP6bKUC7c/5KiXqW3UBrgMpEU7e8P2Gd0xn9Fll6RJwOJyQbSIHC4VL64wT
qmQchQKp/B9OBJumYpRr3Po3rCXnYZBSh3meKVU5THDJ/52/Pn1yuWCejpwGAg7A
mMwQkW01C0vYMfSygQfUMpvosIN80FJDvYp5086TM/qcgaHneor1WzLfVj5eMkzO
wuQcl5uiQTcFnRyGIlzFFAz50h0QzgBXGRc+037AWPlL0+xOoq9l9T3dOCOKQUBs
SgaaDBY3h5ISdviapATLonA1cZZUKUY68Z3SOhpGRa/ytGJZcTx6SSHdg6MJbzyl
DWnwNzxdrz1RUcg3O5LQTlZKPqe7NxlLu99NgMWeNrvN1RIsZ8JQvIQLJMUWMnYF
4296yrgLRmp/G2Twz8+NWKvf18sz5k5P9Qc5iSuWBKGYyz7lH/uiN0aperO7GqhE
7ntRz4GhCisWTjakbUa0PTqnhZSR75dzlNNF/kd3BLiv96VRrUY8yvFsVM1o9/fA
c/o1KifXas2hSnok4rCDFHRxPwne60/TjzD18n44ET0PLa4Kd1xZzjOz2ZIXh6lU
v+TI6ipT4cYJy1avBAEaIJpjkwgsp2tf6zcC2tZuVpNbcvFzSygPRNkMygQYR0zf
QsvYR+ukUesXu/anOxqop3I1ta1V+EmEmm3tj3tTPNbD5GwhrBS5Ko7DJg5pnLbL
kP7uniRtgetcoQW94MCVvKDnT9UCewEJ753Pp6gp7mrtR/ZFKmps3NxNof9ktVW6
LtHCZdOD6rgTuSfSc9qaEcrwZ/jBiu91aoCzVvdxF3WYoKZ2i0pO6P6i0+O/hBB/
HTNciUZP9eLMjGAYoEYuXE6cRlGwq3GRviOKJLCrojItPjpghCFtEKm0hfE95yKQ
AEKCytaFT4wCwUju/SyqJwrBUvoFZm6wx43SwSku8b/eedQRf2g4kg7KnzepDl7I
dwA7zKsSulZtO/OaLStmWoLfJHeqIYmAcDa8MV9ijlPlVwra3cLoaKXu7yXBsF++
M4OaPQoatPYXpHUmZKJx/qVjR5pSYvKv9clysxZxyQX9giWDt9CIzRLCxsr29u7d
urFS0k/LBt0ynkdPzOvAD42bSKBO832SKHNcBmqERmrWx3E0oQp77rp2WS1unOhE
mkMW+jcb8vpbce/sjKU1lsI0a21qrXUu6kAwNcHAz5BJWhc19ALh4kPSxRD0uQ0e
kP784C+F1+O1nDQcdaG81W/yDp3jXAu4bi9q/7DUs8TNu9a+cPhMQgViU4xpjPyr
5ycoUY8bLfbhPM73NZCjnSLpvsejH51mhwJOxA2YR/j24Jhdw6OYriffvDYsVGGQ
ftDxsc33DgzVHIZIkkbnRn3w5b3SV5ulDjf+htb0PKesWTAPdywxtLc8fIc0tEje
kmADcfaNSPhLgQk3jiVHvpl5GAaTg7XU+9qsKL+VVEFMu7zEIFguX/HwQkk8cw+G
cmLsB6ZgrA0fG0IIXrEoqY7c2GLwOzB3YrnoOnE86Qr5OQaVxWhpjrrFw170StHw
B+HwoEwBHX7Tfupw6VJCY1I2keMbJiAyGPc3XiaVlaWEwz4CY1JrJbjDOB/F8DeS
kEhIoesFVbDrr6UBIP2iSHzScv7Fz0BcM9O9flL33NVvQL0llMTNYUTfjH7eexTA
kqoRvsF/aKX31VO+LUJWYYTKq2VZFOdCSM86zroLWNHLboWB3jY+ch0HIeQ3DSDD
sTqowu3bW3AI9de29ByJ7KVapTzea6AGrZmAuvTBhxgnAVRkDnttjqsKb6kumz/7
eAGC3HrsCG3gmdPmOwziTAjMEzb16zNS9PaBv0pEBRp9fLpWY7BsSpLg8egzY5w3
OAI4UrE7UTPaAfJyy4VJc0sgsBf97teWksNfm8ii4a6U+kkzPzLL3AuASg2beByB
78VLLqdqyVdLX3zU5/xJw3K3kONpHryUO16FPVw+YjtV1P3ti50FNaRtbD3HAUVx
8ubC8yOVdx2PtlXQG3BDptOiVtrOxeOsXbpFQIhMVFUVr0rhMsSA/vsr2cjiPivh
ZiWV56z+EEajWofFxAmDjCgbANUJXsmwWz4+MHtZI/Zisx1O1IMqey9+0WNPRv2S
Z5qeYU44bxnn6ff4n+KLO90uMDK9MBBum8+HC8uPWFKyR8hCI8R5KlB+Nbgffgme
PtR7kkThEGj/LGKJ2QmaemnOy6Mtz00OZQIrpxbVmPwql/l6mMkwN75QF0xqA1BA
xCephdo6w94cgCEn22VckIrPVNsFxNQI2RRJUXag5NBA3Kq5wvc5O/YwbN5hLY9X
ySavAB4/tW62PsxFStiXz4ahAhJGssv+VvMYc7hnHyLFheqDhPwt6ljKXPgI2Kgm
wub+QGgMqmdN0quaAv6VRy6xu4s3mZDkm/p01WFckO2WjmK1PWK5E8hxLr8QBkdP
u8FRPCnCugfDhxpLc+T8GSidwtB/AT0RtVhGPQU+1T1IZRZF4d5OetPbFH8NqGip
c9nQQ5T46eYVv9iOWLPjVCP/Z9qPMBIgJogPrgkDbFrhTDuJkgyWfOHfDiG+SA3k
Ld9IYgeoWl3bkF0v+U6ViW02Np9LBNc8lOVWFyELCrYwLS5yurbCtXS6ujxgRTJB
sg480iqXDelJSzIkKh1mChqeoxVR8NnFOeimFnUQoJx2JdGVgqQ6fY03nSBvhq84
+BQ3OKwk3jgRDjKtNzXl5ktsK3djq4og/1DB8LDHz2CBM33xffBQNfbhAhjpREZZ
EGeMV6sm80aY7SamMAQ5csq1PByJLTZRh4NKHwsos1ZKSuAym7rk+FHMo9DkhAPD
f+KvJ/4MdidVdwsMlrYSb4eV6AETxgzjam7ok/FHWeiE9QWzPaV+ORlLUYb675/O
EWo4sr8z7dQvGjuxk4irtQAxN9CY7kI73J3YLP9smQZTJfW8y8FJcXGp1o+hZHsQ
kX5s/Y0V0/Ht/E67TjBDMmdxjMYGRCsS/7ei6gDU1CM7bgfQi+p9ZZiW0NPlyVPa
nkOInHJJ0hRIjQ9wTKJeVxcdL77TZtGZaW60CbEg3PS5HYmFarDEMWsce+V6gbcd
EvJ4L2ewLkqVePGPu+I7vsxWbCVNSJySOIXkHFFv9XFq656y8vaZuaaJCPzmSG1f
luO/1jhPyEVDaiO+r3O+NsQQsgLsgfQlkdYVyHbAtfAbPHaPyWiq67cYN5J65qEM
IjESRyvd7rIfjKvwoBmmWykKmc9FD5TZGX79WfQLJ7NZjsLIHsuiExyrcQBbP8F1
OZhsEgrgZnlE9GcmMk/vjTgfyFlBLYO3612W/J5QncEVJi9SWWnKJ089h5XTueV3
oPUwipey7SBdEcm+cR77GSTSb4qjoPSSmXUZ43epw4qrJxdUvdvSzspMPGnOhde8
WinTXqE3Tok+/ia1QLUu2SPCRV8dA7hqhUm4/loHguj03vLRqYAv+hWHbrIOpnYv
LSFKNQhBsUJL9P3t5IpvaTkKrYz3AAycx5t2Yi2YgXVzH2eQAADWkLyFSu1Ldujw
lxQ5uO9PPW+tTypmldofR/znvWZ8bmTe6YxdIK7tAz3N2+12da2M0TPXxsB8W63g
ZkXsYmJYXFPWVY+YgTkGaZ1Be3a42j2Wps2gtlQCKbunNt2hYFCXgKPR8Z/3gN0r
UCnC/6SxZ0KsYRk31irocej6kCK8a4B5MeePUJLnOCr5aVSzErKLQp9Uea7av9bn
6VN+yEmIPWSiBF1EsGhdyUvGoPOIw+nZvhY0/3xLTBsloEJ7YJKKAWoftnHiXjAK
oeaifrxVOSWD6acQM551hKUcSrmHfb1zeJalvSlj3tswsGs4u5/pvV1F9S8eOEfz
oMXS2yFqq2A+3S9D7qiOtphzt0rXYEsTrljyXOF4MWrfjvXY9SFbxNwjrhxUt9mw
rea7ug6fq2myMpKoVk1SDz5SHxBPxhKS1QuvSfElVVECVeQTjyh4kIJ7pcYL5+g2
J6KN4hQUM5xHdGV4+k7koqLMoOteKaEQVB7A+O67IGcD83X+1Uz0l9rZB8Lr/yzZ
peoSD2H+fdriKFdoJf3raN6YFGGWcBoaeaBK8lftnZI8mkoECjZYDyasJatWLTIe
Okue7uESmSZBZgGzxlICvXCIalmeMI4MxAXnQqIFvYWAFtBxvi45zoAqv+tmKaS3
vHnfOcIAp8tls3xvPYc98Z3tFXSvfjeAXB7h0ruTXFuGAUfma+vGYuFonlRxzLoZ
vjNxCT2au3u4vsZ/OYRMs9CXNzqdigUm/hrMVsHBHKgdkuQbGNPAoA88uvsU0DZu
6EilW1Gs6OcHFg7NNbQ8fMZvHwW3Y2z2uwJMRq9rWVQHXOqf47OqqIeR5epQhGUr
jNDt6ah0wMcoT6zf6u/TbOD++nBx8TNc+cevw9jIaMN//yZEX/V7zm34X9YBKgz+
hmAwEi9QE6TnE6WKRAptKRK9tCUjjPrlTHfo/Km6Up1v3If4QD5fPxbARfB/YSK9
xX5f5q/SdfmyU58koKv4zXmMv2NNnLFXL+XErjuq9qovFP0t/APKRqFXJUhMoc5h
yeCQ/ZO0vKAyDWeJSK6mzo97Riwv9T4V8jKn6boZ6CrTRQgZFsRCY2LFHtE1W0Cj
eHYStu+IE6OFVq8bSS5zDcmWTR043lqdX2MkxH1U30OutdghvwHOVcWfDgnGmPci
xPB3IvQBob1ytjvv6yRkuezPFQCtLvzjtI9qu1L1ixgiTGtn4D9QPlXNCzvMTSsW
/CDcmNz9UMTsz5hqxblPN2v4n/9R708nVfjDdteGJFlzLUpbuqNqFVUHhMFMKzgv
J25FW5Ufk8cGODDRysRPzhIrLMek+MQhLsKD7OlhalhkzWm9xmQMr+nEkkr68l4v
sb7xJ6CnyNdptxrtc6c+F3mo/gZADGAIDqwMo/WtEoa553lYRSevC5/KJajD2MnZ
1Ziytb4Fq4/W0NXOBmFBG5RJEA64rAecBil371wQT1vwqo721Bs5AJOWnm2TPQVy
OO7PSq0A/L6ZvtLG14ZRd+s2SO21KzGZVpu0a3URjYOYP9l6f2G/Fu/CsJFYvGqG
rWTiDW+4crz3qfmZwSNBJj76j6GEDsbpb1s4w7NHy+brVrXaMliA0v836r+OX5Hk
na7pCzw9kbGYyFRGSRDf2XCrIIy/atM89su5A/7WHUa4QP2yQZULi6Dw6UuVBE3K
W3t8tOpf3Nguf+4NO+H+ARCQdUGC5NaVdCG1KZCQpp/OceRzUrfLTB7nqFptvZSU
1Lctc0K5Z61gzaRvOvjIvwudur5DYkYLuJUEsjoeZ9WCNck0fhgIB0sz7InyIFt4
J+LQ0V+pq+aoUPNqYtjQ9LbldkW/pN2MXPQlUmXs11LpBE9S2JA0hU+bQ6eYukPd
/5FUYeIVqh8PN4jGCVcjHz+93z/DcYw1b/b8+PzcMvjvICV+AkVEd6STLkTxXzRS
x2RkMgES97ZayNzc6VysB7HNqKAXBd8g0FTbebiY8cKjl2xlCNzI3rpjXS84yoow
Te15YZAAWQBTSv2Dn30Ss0aSaCfL5M64DwcT0pBZt25syJ8Y4EfNEdS4l5bIi7dI
qPSl1Y0lAOZRlu5mauKcitU714/d58+5VIiIxF/5ClxE461l1Y0jpgzlVNBohMYb
/z3+wZHro1lVWf8z5SwOU4Ffd7I+q54Drtd6kzEO0aA2AA3fEdQ6kEuqUdsvPEua
RmugeCxVXfvlEkSxYT2FTjKEvHhSgbMiGYG5+h9T/u7CK443LaEtNzOHnOTiKDms
IGaKVmacGa/O67VU+H1ziV8y31KAsIrCXgwpEBzwzDkWGZoRlD/VoHoGafbVvpbu
T85KaplXZOrOdmx/xbsadbAu0S2Q3UTWffafqHNl9MN2oIWuHpHmd0O7APdEdBvK
3y60kmRTMR3tn7RM8XxMGCHhpPrhZX3+kMhNiGpZ4yBS1OARfCEIYEeVKXle8tmL
58y9BqIbqcO4hBcboU7YbK67mCHVzYrt+hjQfEeuoP/yyxroZzYQ1DbhHkVALDKU
TmN1wNpqWjBaL13YASnXkaXdS+5OXP7qG84G9fZh+QCLonaNJnOc/999eSCk1liU
dtq05E4zQzkLt+mpCi0Npw0PIqDFGo9uxJQrUbh2jzBeOF1AYkAFHbdalP+IajW0
NO+uvaEtrP414V9XeUa3YjYr9hZJFwVO+VvJ0a9sFP3aG2Rzd5NiuCu9nIkbTdpt
gzaonnWvvavMYeDcTHiM+o1+Vi2Jeq7dhJfWJi5Uv/QyVucZzSlIK3vVb4CeePSB
3Vkta8+3yaYaDctkKQignrka6EzbrBk/mxOAtnojaRTbMLY1vpAImsCBODZIRiCg
TaZ2YjQvWSxUhQ6/Ke6+UNqhuQ6cHGC+B3iAaKlhU+LFzGU+htfYSQjqUKP1trKN
l5W9Dj8YKPgbI81OzszFpY74zy4EPG3UhALq3s9TS9ZyNkx386+TtDgRYMa0Ua5q
oiIpOucX7Oem0pMJrhVwCe6QiYDeGlbRpezGwSMvJy8BbVutxzYb/1cqoREWrtwn
MvfPG72NAptAkIvABDEjoxSpD2dwRe7NR6uQhf5fLTz2z0YinChXUKcI+zF2+hnl
VyYYUj0t9a2faqXJtldd8C3Hbc0cArz4qiXRGrfcBCkgz6cIsMlLyxQiHr/x/RmJ
pBjq3e05BZ+O5gsDF71VAKXPmxPPDReUNZZnMuOQk0TRXrg5LYI3+yrOyACRk9DX
eBLnWrRUUvRZK9qzF/m+xtjHDiBUeOnl44WZH2d8IFzODsyQJZH2RpJk8RGxFyPi
zeEKx4s5e6WjKcgunX/It1xeLka5ZwQ4Uhnhzekwj+TskEgJddp615/MYxRdKd+2
ufGYTQJ4CEDPHvLQOO6M1qsWnZ8PSi4Rq5b/MOr/pnWAvhYppp/vL99gPjyUw3R0
seimEYCsafuSS3PIGmOKWLjUT+g/baoprKLXe8RvL/lBS9WjAXRyAHPd88qyCfrm
ib15ig6ahTZJlXCAD51J3Z9nGi3i/Zlc6+bpYe25V/t+p7RMePb38W0OJTV7Wfrg
pXWSoV2LFy6optndzAbZbsajg1JU+xkw+robzmyqcPc7a4qfGEGzhfK5oidxJ1Du
gSBJ07i+MjJ/+r1dIC1pKciqT1GTMn9a1XG9aMrXng5/8QUSvzBovWzfnoyhNru3
Xt5hAMZZUSdtgPSpJ1gS0Ld6uzK/Y69gvVMYsse03i/qJWNDbeyFOTdVQhd6NFOF
0xCgOARFffT65Si/TcEzlZEh0sKRCOqvUxkzllkuJIXook2hXqlrBSRuMvHJUlka
kE/7hQyzdZIo2moFIoCHwbR3cEbz1Kns4dS0UXGNYqlwa/yngKpfwQwblgBWuJHs
F6hA+ugaPUMypqICDk1a7wiSRSUClwJiiZChcXrIKWurgjyMQPdS1x9/ixCrRabZ
jAiwhTB2zIMXQ1cn9KeuB96qhJgyjHqHEWraMTFSLGH8dBJJGVE/5IoXFDap21jg
dYRPc124eCzxNoVhTlDButVYQDYivqA4rcIiTiEMtQ2Ms854ndCVjyUmuU8aqkvg
KcuYJtuMZ6Jt00puxTPaUdz4FX5qwDTXqfFZDUIhCwHRbZF5or6RifcPZREo2JHs
FbI+h1EIcNdLN8pLzebDQRQHQ3QbO4vNkeirDW+TlI2aW4IM2+pCQDWc6d3dLD6z
245MHIRySROaDsBMxxNdI06B16/YVV6bcic6RiE0ciw3GmAI0tbgFV2CtGAxkLCI
H3adBILBbgVO89qOS4Bvjgz+EwNtQ0m0YXXwXPPiqRBwTzKF+L74cNFzrCU7WCrD
6P1KIMJP8ACVFbp9BGEqnhM7kT+OZZ21E0yw8RxmeHjPl8D1+ypyEYVK1dmsqyi2
mL+020K6PQmTb0aTHXXVTYsnnRopJwu2AInJV9NsWOhQ/wJzwHd/qPwSx8V4cJmF
deJFIgBgJDnK66IO7Yg6HwPDtC6qJUrOTSzcmMXuCPVG/b94cQFJiT9w1HgdOCoc
uUdGEtaVpdNOxGXtWSkqjLritRz5uwnUe49S9tqjaNYihr2+xMAwqBgFXpieVs5c
BA/bBOrik5xRcuxwmpcuY0f1zvzP32/aVB+VfYjy4emOtSHaRoObThuWIeix7h45
jt+dUuDJ0YiLnsm/edD6LINYemRtdczc1mcTceIdnZSKV6g0/+FY2RPTL+wsjP4q
eC4ku49jNuWPdWa2Org3eCsT6Dfhx4HC2QurUm5SrSyxpm52qIqdiHVUjKZvtaom
PFMug+ZIaIbLv4MpnvPvBPVZ/JPWSL5lRuzOwtPZzUryHaKUEbmqjvwm9dRrTli4
+qhfNV8qafAobbBXgo+kKwz2xpyYE3vH6V0fUzfHW7MAs42CI/7+gd0ok95E7Fn3
DQ+Cd0pzv7bm0BTon4YNy6VHY+pz0Sm+d1he9JIBvo4gbvzuh8YC6YhBSrSebtOx
FH7O6ERyL/2MI1n0XzUwTwNBeBzpwKKflzQaZda0+R6skcT7Tg8PFqZ4SwGUucw0
YFGgvxKuUAbgjgKVTOIrkfeF8oPs1XCnFaaLPYoqVaVoTnFtcC1HWpPGa0NMJ2Yw
uwzi8rIDWP7m2QVNKR/azehhabezbfyVr6QTp+gkoBX6QpkNGKeqm/naeGM8F99x
0NxysXb3RmCK+LYH6Qt+/kSRFfa70AbKSqe+kwITb2SJwDKita6X+rtV9Lneq7dY
tJHe3mOhJgCr22nvVeSbhR0XnpO3UbzbJFnwD8j3DxnhEJhhqREw5OLgZ3hJg3Uh
d9KHRH/p3fLcE6qyOsCDonRXxdyAlK5nO6RzZfzhCzLMe1ycclPjtnOK/rVtaute
vnDekh6r3zjMFgqEEFntPeskLKA3wPoXua6/1KI79GZ2r2DSZF4koJWF1ux2jAH4
7Nx4tSDsg1sFBMSAlM+lAEQHo2waY6W8hjGjWlZmVHm3uehniylQQBAAOsFEXW4+
7Htxd9Wes5T51Vdqk3MVDM4/Lhqg01WfeZMy/+JbfEt8obYMiFJXefPYGaZOeSPs
g/dRExBbpbQ89X4uLXpWBkzsgfqxG66NqbuyXihXUIhudT4PkmSQfACb7ExlhKu+
3YKqu4Qn2z6pjZr+dcQoK340NcJd3nXE8s+4jxTVMQLwqllS22qo1IW50mNvdu61
59ATDslEkUjkR8kffjmtBUuYqjLM2dGJEB/OmpdjYeG6+IxX6LIm7+frQBfTaQbT
wb6yNWQ/qJnwEpss3jjM+gfQ/8WJXROvpi9rYFDtau9etCBEFOLgoSFnPhfzbzn3
hhz6ecz9dMcSrP3s9M6mlUss8zzWPjGMZRZfVbUYydwsAXKP9Pj20t2zRQ6U1VmJ
DLfSwf6XduSqnGpOf1ospJ79NqVzgsgg2InZuL6mhkfP9sz2RxbLkaKdqQrl1qIA
YLiqKqhjt060FfwqGF2if79H33tMAyrQQT/y6t6NFGxunkVR9Xjw1rXM4QrDxmKq
8QghJWb4/62doNkXtZiAVpzpzonQtna7iwWOoRP0NDEKBGQu7vKN73xnqzGzxaqc
sFeM9s4A/GUtFh1KIWuRDytv0IyeOsoJIwyD4pc189x2MAOx740gkTqSscbilt0d
JP94X4xMvBhYOFxkNF9Y8ObXyTeZPiP88/Z9tSyVOzq5LGQCVnryQTr8lLQA6tRD
olttLJfQu7Cj07Vc7lfhNmhOK48P3SzOj9KIVu7EksP91hbbnECxhIKiXppgeUfA
8PR1+9v8xn7I2pGLAFA+WCcsN1nx4YTpgL5DEU3qPG/sF2xU7r5qyMNSXthRsfLr
zy7Kk6MQPrk4Il9VSAfAaGRKOCjSuyKZFJlubEWmKblTEAo28wO/CuFPC/YmhGVN
bE+awwa0w9Ssmipo5sldQQUPiIdVMZWHwcrVlq3cVbqYsSjC2Q7yYx/i23aZRPne
/yW8Ena8iCPsOCnKahD4DcHkUQ+JQFaGovGKKCTcVL02ovg2oUo5c5CAbskMp6V7
qmi7b1HYaKuHEfYi+GcyZf+DIdhYhpuX2TiV3sBHy5k55R37AX6MK2T7wWiIyMpK
9RjCdoE2hHsNYamIbeKr4ICgJIMInANF8OX8bYlVDEG0/ZeUZummMbqVPCNMOjIh
WkU1QltFBR4Jrla6rBwCuKBwkQ5hpxRNpOGhneQB6MEfoKGa5YoRD0okqK3hYINg
SVzuwJZxoBh6MsBCVi86DJbRqbaZ+wmFTAO5tcmbSEoRrtlSgJZd2wMSVsOUKzWl
2QygQB1WD4Dx9JV4OzTbBVpJVpT0SqjTZMyM5MWFKSFa9uuxYjuryE2OqEeRKjP5
hMjPOd8NrWPganH+Lq7TDM3nF6Hupi6CmWHdRaHOpbAaSRbSq3l3qU/1E24JZoOk
gfVVEp7IGLE5POHp2BYqwq7MAsiarqaZoubQHxmw6hkKtk7mcg0s8yaOETosG+/4
xxfhMBnYudsjl5rt7iTWOIeRL6FKIYyhWhwy4VCb4t0BGUIxNEAQA+EKcVTzBXiX
i1aX+Jp0YMnfnsWnPY37gXOare0jN4lodaqmvT+reF5H5VFfJtAMU0u5R/RS/LNg
rZJMhRL02ZTbeN5y7/Dn4gqyiZugHoldoPG/D/K2fRm2pc/ltt3UsRvLm08/zn4j
TlhFZBdZOSVpPr7OAw7xFksvinLZc7w2BAOXcYbpBenUiQxTPwWb7Gigy+omnmIR
7gkRimERrkGac5MOG7hPkur62ERuFtulfqK1V0N9SOi2JiD5i+UbXyfpMdgTmScY
2wxC92C+GqlVsi9q2KixEYv5emkLbTkBmylCV04Uq2JWjDVrxZamBDYQY4YNLUaN
OlZd5XGSxJyd8ajJuIhk+HsadCFbJjqm2M+Qq4fJm+IHKWZTtXQr5cq0hR9dyJhP
EMUxggd3uTy7FwMgzDtkJwlzJd5ggWi74r5YUhtuVNlvM1HNClWhiBKWpVubC2Hj
cFHM+MK77QKNY0nrnrIRZVCVYhcMmD3AiarS2XHoH3VtNEa/KfaPgJ8hzVcGzT8p
jcREVhRnyCoDUZcfGZbJ/3nDETNT2m4EBSMIK9fzV7+KKOriY1hHOluXERa+Fj0+
TKx9Zap+oGVq0f6dM99pN39gbIBmggO7PDWixWlsZ+pT1F3IfEhWAjp4nMic2eRn
ejZwWnBPJiIALOKOp7Op1Dnwy2BujOHaxOvv/otNYGJmd3h6tq/AcWeTU/mOIeeo
Da7tqk0jYRK9Ngg+PDHvGkZbZso8F+uLNwRNL0qEMkt0VNpwAtYqcZdTH0GbiJUm
gBIlsTj+7b6HijrxBU7b2X0SFAdlLTtTbC/fmoVEwp76c6z/xDGrdepigWG3L+sl
zG9PG3n8Y+NUj0jTUNY2mCY2AH10yN/Gj+s3xHZT1tMCWfBmnUrcDeFzyGh7NN91
CG6LPtaEQsycEKSEQs7s20cBxWsh0IcEGgQKiD52g+8JbNUL3HL7BeygtWlyu8Jh
Ul4+13Et+1iNXGPjCnBbwtRitAr77UhEULISCjgFtIaHrnqfoPH23Xlo4yd1/ej3
Cp5juuC1mpLYZelT07ZGhxa0MQSTXj9HPEBncFnXl7FavANH3KceXRQag3uAeVPh
K0cvRGbozM9CKwGdYLjNyDT2kVDF1YhwLB7OnWevwGxMPJMLtYqyw2QxjNzu//fD
o8LP94daj38TL/pFA7gIf2nezuErv+fdT/H5vWeYuXli9Fb+duJ6dyOS+0OHv+sI
TPSGArIWNF4BLGITExYtqnEeKNpcUTZ24CO+GoK7dOMIqLgUrjCr0m+8396Rv3rj
t+W9pNKyVs3mA5k+XGx0ib10zwPBEl3DRZV8FZoQiEGkS0xvoYAkG9hL2Pg+elz4
R6LK2KDN4fZaWFLnI7Bmyj0GKrojzFhJaQ0aBEw/A+LQBK68IR+vMYZlnF22vL1d
sXSy2H2sYpMPx64VBrCUjFRtrrGmbUSvXCOQiSj1AkuhOXbUZ9N7fCLE0qBq9bJC
GwQgE6BqLzHSPr2m3qOlvlXgMrRhHamQBHv5eEruaOWrMMMe9CgARDYkXmwe32Zx
EAw/d8t6VQxK3w6z3bfW7VvcTbE7L3FHtqYv/VUAIcZeNS13JRFMt6Ro8zNsj+Tc
XdLKsL5KSawVxz40xE/iGOflr2lNQ3iPc7faHS5VDgT8Gr1LzwaFnCxc2eMFsE94
0l8aGeB0lLxkFEX8Y5qZyxmjAQpYy2Ivpfzfdep9dooR0KD9xD56hepT2M/DNgSh
JY6S0e4TAsTebpudW0QZJxnHOjbNe+DnPIyZ1KD04myXT+/I6XO7ZV8KRi+9zeGH
Apdxqofl4KfEtsRDL6F79IWfa5XaCafLqwov5tanbdRPhII4F5R04eoyZ4Rqh1Mk
CKV7u2TziMWC0TIeJHdr0QIkaN7YDHuq0+iQc/6yMY50Oq37jqeLWibW0Wf8pDjX
3UfRHU7ZwRmnn2lDRrMty1N0tYTFwMCUQPc3cpaXvnb5gahufEQow0jQ38NTK/7c
bP8Za/XaQu1T6ubo6KNmu4IVBcNbd9QDK4YCfqpoeysDVyKhZxv3E8AXDw3MsrE0
wTabM20/QgYziDO63EUxijEEOtaqkVe5jUkaS9yTJhvcsNAzAss5HIDzsqr6+TK6
WTm7lzbh1GVEkjE2TJ3xgfj9JQ2oG+iuHadVnvHeW0QjK7v2EXkfpbQeZl22wlLB
tfeJl1obLnHrYEK7kJns0nLD6dBEVhMVKahZRbJLLiKu8Un/wdOEd5rgOhd3dxzs
dsNnpN+p/3tuvifn9BpcMA5RTZn3KC19736W8RV4vWoiVJDrcHX/ZWni5bk9f2jp
mT56cq4WNCWpGXMbbQZHrldfwcLTDHiTY+gwNR97JmjN1N+ScXoFSX/Z7eYy8+5N
sgolzZJ70YE9wSDrOycZzxDernyKX75JFDlfQh2SMLXhyMm4kEEp9Hy65FWJZE2f
OtKyPWoeeV7bRCTfWjRs+mTEK8ARemXDwx7TD+S9VSF0/Ec6HIFJrOWgIZ7LjaAD
lVL19EmY7ETfJeRdgRfOZsSoc2dZj3/7E4YBvjTdlmegkum72qfjficxgBLJbBys
Ibi7J/LJi06nUcVcLyNz5WfHbQZjwmVp3QqtIAAg0j6ezrFdu3ThqSe0YH00Trmm
+R6XpFgnBX4AxdSDzAvzo8Nw7A4wBCoHnJWdC0dJ9eZvFkiLqhZsXQ76lvt5hvAm
3nJUMQ+GIBGGvlmEd6wv0G0TWtfrCNXatRCqgeQX0Ily7dvn7fpMpaBV5mbqNf6h
za7vsDKtF2mzvdpJFQs+CBiE1oQOJ1YnFHE9jtHYgkier//w255x3vG2zWA0P+RK
h9g8Hi8RFehKQOpiG1GJQuwG3/ySeK0ZmUDkB7Pb6ZQlwbIFtbf+8wGnIBSa/ND8
SDV5abHWyrzIbvntke484Q3kX0/vmNKmdHltBzJqFtiFd+FkbQcfDgMQ0VGIWS/+
VF+8bO4NQ+i6emwiNaGiLDOFIr1c3O3vlTiJVoRAiDMEXxTHO+l7GwUy412dyt0S
8ErQ4fwvvxoWOLUKDIs17mX5KrHM0+wUqnKx/HHnxS/tQ3x1L7OJNwhl92NvR1VR
VJFArmTLhQ036NT7u8bpA47HtUwh254KUjvWrMnDy+M959bmcLPlbPAbdc+jJfAS
fIb8EM9ZEPLPQDnd4H3q7/cmEot5xS/+RbPkyTRDsXKGGKoJjNwVyt1G5/Cp89Bp
EKfUmsDDubxaW3mo/mJQZf0IPXjUGP+uuftY7ERoAasFvkYisiMx8G1qSfp2CYPM
5C8+oiYdwx9Aj7TWChy86jTTX4kXFizMkNYUIHbkqPEtQYKP/6q9UO4rz2H+bRIJ
pqfoc6Xi2OW3R9DKJmyUQDC0ZS96a88QhDt0ztoBNtWAJzW9beSxALuijDmXUAXy
o40vo+wq+9h6O/lBhpp2n3ikWWrW7gxQDvGvk62Ue9wzpLk7fohJ1kyhMameaG5f
1JamyAKnmUsx9iuKdcsaEpt6kAo4N1dWQeie1z/WxME4iDCjd5nlB5HjPSlZOJxD
5SyOP417NTh96lF6gJq4dPZJ4aRkuFunCntNuc4k/lVqDyEHBWn2c7P0E20bUw+/
Ut/VcWOShhTvC959Z7OoC6aQuxsKyZedqkMxYqGF6ZVlqOBl9XJ5Xgpb6i9T+v79
8lgT3bbr6jmdRHdcJysIRg4da/AaqwEh0uJn0wa+5taEk+zDkljXGRI0ipfXFoFv
H2tWNo8nLqROgj/zsM6nThBq6RlWSReMF5b+itZhT4++6McQ/hhLPZWx8phUO3ne
zB+vT1YzCQF828V+39GmNwf1kjS4Q1GJ6g031pNJywc594mStOAI+it2h8IcVXjr
E4UOhOOW+1R+dkT4Q6K+COPIZ1ioe4r+bOPPrbevw2qPtEW7mNpxdO/itFS2XxRP
G/HSpW113oF0XMVEcY7z31u3Pe0wQMzYgiks64gFl3UJ6nVL9lbPt2uOwgxfF8QE
dvb4ehaVPH7/9i2OL5nINcikyMgYBBf5+VGchxCvKaFDtxc7CcY3MiU7gt+pDGqX
i/wRU9Ofsr57umiGatS/1mIBkgNkj589uxG8oXB0s17usn1KBBrYPkt6JrxJN118
VtyJKwgow/y7jb8Fzx/ewWDiP3ajyBEJhUQEETYW98j4io2KuWEkGfGRAGh94MoD
g2/57WTtZ3qGPAnocl+NZQdVIvITLofgmXauWN02HeiDc6S1cdQIyuoufaXnWRBD
fNfCNvWzRHfchBfYlFHbyhUoC2NxOIahRbToRQOdGArXwXP/Dot9+oFpOrrm8Q1H
01FDqrkfgkpV28+zv4WwaWyWUDXfgjkkNjGjWNnH7WlfeBJ9VOIqPAkWVTBcT5PV
BGGyaI/leMbvxHB3v/zmo9B9yN4IlkjhDF3u9tgVfsFVfBTZpFSW8/e+Z7f2mMvx
DPGlclzTRydfn6jyREHAE+K+S/RDH3RvicrAfgTQx+ngaK+XP/xSHtTIqERMz6bU
I+6m4sxG2wKanY3fGcJEdeDqSrA0qKL8p2o+8APgzCyk59d4ebPbGyp1IMcryXXV
RE2s5IfRfP01I/iHt3mDLj/CEDQWJdiCA+x/TS/SPfD4Tqn0y9X2nANoP346qHxF
8FnXLf8qsX6FF2De4chL2UsLMHfRhAXI5d2QOqz4acbjL1AhreLy1qzrh9wE7ijL
10tKMEhnG7zSLf0oMykt4RzktFjcM1ZfvRNg2rZKOsD3pJNM9y3IK917B1/zMGij
SLokxkHAwddHMymcaFeg+AqR9DYEYr6+m7QTndvRLvcZIwzrWc0z5MI5b854RPtt
tUx7f8f+mFi0wPXOKm013YsPu2ZjGi6ucWI5k8j60VMM218xoBbzSGMxAo+L1KY/
FriF4x0hTdnKoTzJvvYWWmUwQ23sGzSqZllKSeQG3AYHWFB234Sx5UPWNHs/kk+6
J0zo0uvLT3oCJTCKlN7MYM5fwujzc9FAT/Vu0BZIvoWCU4bPETMKQgYwJpddkdO2
4Oa4/ZoIhpOi71zyucA4lxKjjKwU0CX6n8t5cYhWMVt0ub3kby4CDYG82mnx4vfs
y3P9KRVtKHhl6XlLsmR0aG+jyLRIwSLaVzsUggPKduLdtOn+Xc5CD61HAyTrnS3Y
E8n45ha0gj8qAE+gBL2RtsLBXdZXAcCFaLlk0pfnPTor+k5mVEB7DCHE44LqgvzR
SUYehzMGFMM+GrBCw0Qu+toKEQk7UBVxVfA1H6ZbjTCU3YAMTKOC/+R2tewfmZBL
AJA6ORgLgJ0Z68VT/T4elNwNQOoMmFawfHVvjW9IOr35rIS5DLbgFkaEx6YQ4Uzl
p2yqJ1eRpVqTQkNW1auARgjWdk6J+yIwRKVJM0gZ1UMxFLfauQfajxfglKYGRsZM
4ywS0Tq9nHFZK/jmR9k24eXcqscSV+K2qzV/DQVoLi5BqecfqGosoI6YcB1aK7uS
GPA1qKMvDdUUOfhwuJF09viZf04CxoCMR+5wch9IVC29ZZFDX9Z9qjeQzdUDhic3
CbYnCz7l76jOVEtz59nn4Z6IWuJBvYP3kg60SGuNf/nobJdOznlI5sFuhIiD+q26
YRa1GSLCK5DAr+9VwmVFPS3kXNkKy8O55W82ihdQ5YIYzQuMt9onbYrgH091X6y0
cLlC8qmY3Dqwf58qt8EK8FDFLBu9MC0VeQoHGDMS0WLYAobaS6QCh2wZ1KW8/UJD
aLNQLZZJA2izACM+qYUaYCPWM1iMstAePxn4dsIRIZ8Lcr4IAuT0hrd+mH2r3nwF
qJCK/HoeRzFcBGokxChXwLHDmFSOzFhMrZk93xq2X/qxQXiGARXjXYnl31P2DuZY
YJmOHZraXgjB2Lvx4GdTOySr2dnpG+5pTNAxUMTB8606qgy+7/chTZFfEUkII4pg
TmimVae4s7TALz7Qyj8WDO8nmDgRjiSejvrqEUq+W0z8TBrHiqNDk/U/LD12Le4I
6F3vPWuRPJMGJ4X3zO93NfY08WuW6usrpGOQB13R21sjC2n1kZnK7vOoxXVOTqZa
GheyawbI9V+av2j3KpiKWRJbWdUK2XY0YH2vn87RXYBdHLz20MfnQv56DMFQ3oZp
zdehdyey9JXuqIxH7OeqYGPpoqhhzHJpP9cYiQWfESASOQwyvUbqxfhV48k4hiU1
4gczp2WU2EiCgQoB6+gMWx+WepoDJFFZi5QtCJ37GPYMgG8J6wAjrhxWE/U3uOn4
XZ/sahWbKjXI3ieg8cGvQ3Y0Qjn5+RxI1TtDmfwQQ81yg+PvAsbzkbmeSLS1iUWR
h2sEKQ4DbuwQsxMIUqDRknH+mC8VO33y/pDTHYshhKIC3zg525FJokt8iMDuoioY
4BhatRcXJUf2iES7lLmFzYFkTmN8B7dLromAiYEg5ZP4TfehUqCo8sHZzv1jdPZJ
Q9Jrn2D0K7EVK2YkxhMTYMzs0pBGb35sKnm2g1qQfKnfOx6FaqO/9a9cCxdjWgit
r3YmqmG3AcIfMoCY1t8I3zfNpbJQGwRBxwhb+ln0gsCYjMGXVVwTnnJ91Hyo7pcl
DKVqNpSOw8t27L2YXP3+uKyDBkXXIEkGtxE3BURvS7NeRLpzIJaXCtzb5F4HD7LY
kRYVr3a+FoP1+ffn26kZnSt5jor3aKSQSQnHqutXKNUU93DqKVvwYlGZsWHoO86+
ESgbgJr0lEtw49Ky7x5J67Rbg/w75FrGeVIEavdB20kUlQF+QQD7esJubM+WNuTl
0dXGOiqIwWPYTeyCx/lIlFWb+mhxYYFU2lO00uZ1XD6qezhvarbT90vI/WipQ1dJ
jEpL/Cuklt71S/OBEaOu/8KIsSOS9TFcrQ4GS5ZBaQQMDGQ8kEIkw31J2o0rEnnT
LfDU4pOBOiYTgfpW5cUStJQVEUEh200KQD9x+7CmxqtzRHbibKEDTy3gZvPnrl6B
VG3q2ZYRZGrdPdtw01dp/Qad4wkkW0XRQyD9ZIGX8A3FRwb5H4bjq+Eiqikw4aVo
rWJ2cFqlBosWXi36rcbAf2mnBl5Jqfch5mVHscdCRBwhMrLPtjJ3XJGfCGaq4ayS
wfyYP1P+eN82L4snDlou3DtPEt3sEJ+WEs0lATc9h6EF7D2Syzrf4CeA5IhV+nbJ
8dQcuwtM8iI3VYE/gautDlZtI9V/uCURZ+zCHRIGQnv9t5oGPCyhUPirAohwxLwP
99Qi/L4ybO38vcW1BNys6i8EBE/GxiHmqDFlrn9mMfji9qjGTxaiciqmwhS4xR8t
kN3JmaOLobX5P/SgQmiwo90MO2e4eUjnWJ1F5SVq/gtUPmf3FZzViMJnonQ88EKp
ZN2dCTTTFNEMGaeyy+DGSFlI5aLaHoSBFiUSiVtTGMhn9/YWHOUyuJR96tPzf03O
9ORKWjOx8kjNX6hZ52/nQvaBxu5xpW2L0noxSPY5DLH9oXd800bZ9Ko7T5SnNn4M
HKkT3WRh1E9vehg4A4rNOM8FE5hNL1z7M5QoYwLt3ncLEAPW+B4WBV6LPB/9AdVO
a7LqrH3AxyzlXSKD7Jpcxt2XEFmepnUqerTvsKbcPitMY3WqKsTYvn1YRSXMAQjM
diUsf91St1roJ180mWnLBVXMpf2M9RfXljNERx6YR3XOMBQnAcl04CgkhFVi+HA4
CECpRUJmHV7qH7L0E+W2Be8pfmLU5KhrU9x05BOjHppMKIdod9ffcLy+XARys4dv
T5YLFVUoIDqaiAwnEAWJu1fxBKGe9cfBALeAUihu6Pqft0KobYMP6ymGdzBj8xdq
7wk7ZwTHx8J2FFbbh28OafiJ7XiJ7pn8K8INlxmU0PPCY0fFinxBZLBujPSO9pSZ
GXMAQ2XjujdoF6jnpG0H+xqxVDS6BKiZvBJARrAABle4P6GBNdr2orGcC89+dTcL
T5LoIJKnaTESUiqXezEafODffFs62QVSm3MiudFhDY+FifOrx36fPWOyO249SM9K
isxvndYjCI+EspSjW5IZGlmizsr2uNAtQvEDg9/GYZDGorLRElWCGIYnAMKyug40
zuQ7twZL8sc+zovuOHH2KU1dQRnEbipXOeHIwLLrPBFPwZgO8uvHQX5qdjbHMlcF
Nujy042RN0hz1i6+mp4ZwgDbIkLzrGtBMSM4s+ekoPbpYg91csUrhsVkbY7Jgn7B
tVEd56UzyJpd8X7JXpf/q6pZvk9/xUVdP+aTssrD6X3A4LM4RdoCXbtWJ4KhGwe9
yCJwzLdA1w5ZDPkHDavgJsKe91IgFSPQ2ah6SNyv72TFP35F8f4ie4Esa7s53v9d
3epcTbAcJcvSn1BWRkhCkn3mkR10eS0FJiYTOUF1hkn1m+7ckETsEbsBVRLVEtfj
/HLJJ2Go7GVk7shHr8sC7U5pDK6GOhchoxSeaVInOnEs0hj9cSWoXgVgPLKjyPNb
8JBdkb5Ozxu2MhuVyPxeavGEux+8FjNC1FiAUWHpBrocMaVsnn1UEnYgqa0tkCLI
n9k1fArei2ffczT6FqLxzLyxp2VB+6b2ge32gdh69+cP04S+iyVUpl1qjEGuyL/s
ZiOJG3Xw0/lO1b33ZGEDcJw49PSqSL+AQ0P1Lc4m10qkUFYBCSajhWthe3jnwjs2
U3W1chJxgFdGgjp8qF2w2xJ1zqWyGWMeHJ0LqLucuEz+evB3/mY7xORaK2wVepno
Ed9ds56UBz1Ku6FOVlhv71CDUc3bolAlINsT4wbxfGWajI6vBcwb4cLOFleOA2y5
mGL5pkTUrMxJUdnVnLYVHxSBnF6T8+eMBERYlrNj3BJAbpcWXOijXHn2ojjGIMWY
TTYNVG6k/rxVQqAIgauIdRZpW48y3PltHM2kKOcxE0oBg5vtdOCQfGDwSVTqMY7e
+NViwWnfzw3ogsDkYO7U3F+uFVU6KYM9bQOW39BL3Q6GeVyQvt9T7s4sqe1aYCT9
+yzRWltus0KWBWh0NdEqzCE3b7+WlwB4m5TbQtLvJHMw7kCQDhN4XjmZyFmm4dXL
WZ23Jdwz8PpzRow2sXSMt7FrSWUmd5WUfelyF3cbHMtG8gYRC685HowSgEmgXHuF
9uvIb/weADTQHkhRR6D57iSN9yupEOfHvvKGj599gkP3x2xtfhL9bRttwR3CqHvT
W2y3aev7VoJIy0MuprqvlAX6WGHwA4UNRcmDlouZ1s2KV7nSC6cfSkfDOl5Lis2a
uv148hKcYH6du0JFV8s6bGsCJqp/2iVvAZ+7PnyftmumbVr/qFKBe3Om3Qc4jAGD
gKOE9MSky5lUr1+dlz+9gKMkCwKEC8hAUJRGhI5U9ISp0NkWEqKWS3pJzGg0IRDf
wX/2pj/Zw2dMb7jyjH5FKwmeY9A9SJuWROiARLGK+gY0Z1oem4plQQ72wpW3fPPd
aiViq7d2APfdH2yZleBNzymHUPHav0+hM2SsOfRDG83pFX9eSL6wStw6/OUJN4FG
M22MoARW8ej3giYbG6oGIXBGWQo1Tmu80MZE1U7/k1EKXqvVzAMlXhvJYj63DFqV
DXzxBP3GqygiPq4VLHasAAHoGeoBaZkLF3vZfLLUPnGUmUPXp4QOgbe7eJDchm4E
XNvQyXtHgkYauh7gG6LIFzlJkVVR2GBhn9NEfJBbT5qCrBl83oXLIjByg2KtQLKe
WY03OUXQ2GxOXlZDXC3nr8YoJGO12YhxWcS/0yKkPd2C74OZTKSNg382sZpiiW0e
bwndl1DednTmVZh1d1wj31yDsg70NsGzkTkIf5zsxMmVL3mAt+fHUq8U6kD5j1XA
Ww7T7H9LRPVJy7cCg6Bd2aRFuMjXwkDDO40/g+0kRY4RRfQuWSbLF2QZmuTFSy2W
ivgaA98iwV5y9V4P34pdNODfRmatFeIHMurDZkYYM7hYHFC2RfC31/J7fXPjb/S2
7ATHueN4fpyTrcSSftg87X0frmB7+CfcOPO1ra6b0r41j86nA8k7ubXcPkFO/RQl
64X0dzdw0x5gqJyiWkLSXLtkAzkEuopdEz7s/ZlooSh7sUlGcb9LQLkfoI/azwX3
Plqhm5z6ye20wHyE1+fLqv6mIFgJUKerSC00l0uFphcg8EAwSZDi/34YPecmV1Ac
+nZSocoCFBmL9tWlCoD2SlV4NaUAAu/KkTgFUPZnQ/REryeHTYV4gthKlSPjxDri
snT2QmjbNusYvjRUx6rP60Y2Dy8hvy8ZbJrrkRQrglMNikyyoN4E1S8UopZ+QwyQ
IOSULFfBLEPSyfRyyXqhtuLF1/sLtXL+Mr2dBi8AhAedpP/J9MjztUH37TLkpJpm
gIUbfdQw9E+5lQNiUdFyULlZmDiICyQoR5p+dX3S5LQc2QKIwNAShm5AnHyTh4au
dKqiPl0upzelDxxa0IpUJUNwNdEgQNLsJN+7achFcnecmF2iDx2aAf9AegHGzxdR
Q83+sCl9lQDX+xMmrKPZ2TBYqjU7/UwoPDosyZm4UHyNSVNSGPR0tDXBomiddChh
4SFJ3B+Md4HK/jxqj9nJO6OR/MOT1Oypts8Tulvo00n0b1FR7mCLvTSHf+BVfl47
lvVqsdxRv7ZtvLgHI4AcXNM28P23teIqTtp/sbqaadx9NyLD61gTzTDUX5o2cvan
u534qySuqqsunLAACvr2AYxooVHG/TD8Ye3CFuAXJbuhIDj0iqvH5yRQvWeBlvwe
5nCIxaP3Yul1uVCT6ygJoLe0tTW7Wt1y3Odh0oRTXIxTcqxMXa45xtYGIV4d6OF5
flvvTm/PrlRSfMpO5shVM7E5Ac3gq2A7EjxKnMEEnOV2jQov+bmH7aQP9YrSNvGF
he0BJrkfG6NFlslhXn7P9TtlP5Ze44MGZpWXBOIfBgvl7TGMXFP2k79Te9X4MmxO
cWXj2m5YaGsycBsjS99p3VBR/f3/gh0q1OdHKJkDj6xpv5JX+IKtsMUsNTRsmwUh
QZzm3da8JgA7jw0RXSwCnmYMagH6DKuXiLec+L+5bhQJRWzPwJgQKOz7QCl0DHd8
j9KrkPJhUKPjdCLdlVVXGpJYBO/reBgUg2JxllY1NgQSxnK9p6OkJbT8xOquHbct
bR04Es+U/P+AzzcbAGudCkzYt/DtqRwJZVrTc+T/XT8LvwbPJmpbAWjpZY25odOj
eDdxAA2G8cVJnxz2XNuBaQy7IfqHyzGvkMEUWx1Q7Ru58wxqkYZpAozmhbyI17Gr
lPc6yxLq5ruksKSgj1JZZAgQa28AWxCyK+HDZLDHhDL+mBbw2gycZMSnOdCDOxJ+
au2XNtg9hwnmtJ+EkWXFFQyI6UcBU2SM7napChPlVmlz7FIBNxJNRrrF78Cllifg
ZuStkGDLzE9TlSXVA/Vq+/D8u5AAWGGKpY1/g96WdU02zJswt57Q1VWm4WNh3YDS
UmwCjRIDUtbysLe/QQiSszBK/WCokvh27eVmVr0isOcnTenPi8eh1Kbk6VzMMCY4
gxvJST9ouduWRAYstTIFHxTJYsCWMMRCavtugGrCc9w+SbT7j7p25KKTtXTc4ypA
sV3zkJBB3Ul+2Ex214QrBkf8azAnh0jXCiK8Q6/Cz91lwYzjtEmRMiY3M+EkzTBE
XgHAyegmBppZsikVrghfv4Di2kLD1XWCV3p2iwpdvQyV5bFk37q1luXDnUPE843N
28N1EX04KCg3tD9NKCkaOERfYrXawJ1MWbnLZROOdUD0Uw7FGY9wV6oPDAnbiDS8
HpV9CxYctUcb7FekzuRB+JDRfINAtwuyNLBOYzk5QXgAWYtuAnb+ckdcKPVn9KRX
9tJVBOJE1pwrUMDjTG8o0WtwChnCrqlo7whc1yf5n/l5JV25U32sWd/Jq64MuuR3
TgOtP507niNdurtq45v5XujtWKPkgetiFEtlWb9Kykzc6jPdxFftk6WTq+u80Xu4
9vR8Xww8CwBlUG/9JIwOBcus8ZrzdvoD9Ehwe+m1lRBN4RFeRSZcpeJTyzStfxCC
EbjqlGYh4IChmTbBap7XDpaGiwt7huKKVHn50PnTpMsYYXxWfL2XflmsgfwgFbdQ
zHbsdsK16iCCeYN5kYyYU8OmOYomv1eVTFg2fNC86761T0evtHtGhnI27r5mDTH7
V+rWtKNii0xIa96iIHzTaIja5MJkAFGziot5PG7QqiYEBl78Cn1vR0VyAM2nXfuX
JFG1lxSm9jTbeqIh8WgaT/CbpuRuw8eUxBwzU01N6BLYMiTlA6SCydlFVvGJpxjw
T3ETFUpqhP41R1Hf5XazjuUebzekcHvmFMk2xNO+1I8mjjNUlER13zbcAGc3nMi5
nbcPAKmfbMFUahiWUVqcPdMTAD1Nje4DShk7O7vj20uBZFlM3XQbB7bOvcAI7eJy
uPRBQbpbP9P3LyAYIM19UjVd2h75tJm3nQkmIfjcUopV9eS++2HVK5NXe6LEh09I
ZASIwDcA2Io67bVGAV3nE91qcuNiYIAp416MWU8vUxP/oYQ0Nnpq3PPWdKD1JCBl
uoJS/b2tlubaJX6D0tujXqupefN0zxQop36U1TLyOXKgmT+yIsn4Y9H9yB1tIgUf
UJP63JiQXTHaxmydsjDHKiE7PD9tHSdXu8BocFm0zEnJb0LRrioxr5i+eTVWxpGA
8OeaJU/6MSglcH0CfVxBW4bO936KDPBeSzC9hk6UvXfrl6kSrwLvde3/IjCv0UGJ
SN662bCfo1Aga+zSJFrvY32rNUfX24xQCSV9THi5sA968OZ1LlqW6LtVCiDMQJDW
vVYYgz0LbYTkuy3JUcnyCw3mbNR1j/YT4uazXSMHFq5QE/VtOQ2g87UtVt/cfhe0
wdsdfYrPU+L9WbdXTO+ME17ftMWkCeDodPuCWn6FN/F8Lra8b2mrKTbqTMNB1uXV
p42uyxhUfaIAWM7DiEMF0t8EWOkLfJ226QLs/rXgqGG9nvLeYqTlNFu79kQA6t/B
mU/dLbF7NZsxtts/MCalQsn+oKINhjpZU2Nqi9medbnmCzO5SuRvSJ0K6hIu2Mcs
t09i4pVan5zAlp8NIbHeEgI+z7+cVr76Kykg5y4yxR1GsGWqzPAaBZvP5+GiZcUs
K5KcGx1VaMIOzvF9yeUadjBiwB8GoMjX1j8Me8/uvzLxsuO26GEywaCrnu7KceTV
1mO0SDxL4ZzZX2DpOT2zQd0W2lYm8+i7UvKiIfTdfAZNia9dqGpzbjJSnRJZVNZe
WnFzDrIwG8JvDuDHgMDruSJTQQyQsRBVOiV8UkN/rMwyfdzqbdeLZHussAR0dtTK
iN/2TYL9Cd0RMFVPibIkj+EAYHi8Q+xRT/sT5wnIYL4+t3NgPJtdWkzbJDyD7mi+
HVi12lcBDVHnZ/lZZ19bIutoRibapLb05/NIVFhCXKadL+wqgGERkaW43pJgQkwh
RKL+b0SAUmeH4j+Xr1SlPhtYN3nElR6Oj35TOp05jeQlHO0bbZ13qHxYuXuNh8KM
sFus3/IGCBXEIuhpO4mbD/BhCsAHFyiH9XTTqogWp2nLymYlujuO2t/p1njZHAlq
RMXFW9rT7Qg5Rt4EQuN1eoC3WcPmfGKhPhAiWwRdxVs3GVK+Vxz8aEIVtb+oylBF
UYC1MoSxDCmlqmDO3hiPKuI1O5yKZZPqGNF/s9eTSgChrmNsoF/GDW+6KohDMsBR
2CDOt8TwuZ3uxNFVlK+10eA/knPPNQBFu3ft+xg1bDyT0qhqHJ7SuyFAoDIUTTI5
51q72K08FHYKyfXK/zVKh9y8yJYvGhon8CJNGlflt93OpAE/vPBHXIU12+O1RP6/
gmOHaEYgIeIPakIy/yOflnmVut39p3bL0uA4XbHCdTvf1JG9vDGzQLu7xy+3HBQi
qyXDmINRk4BRuir+08yJpbMOaICAXdjTV5qIopYBODt2UMZC5Pns5COZYlTTc75e
xUkza8HqlacGdjBl7kNeEWuDLR1DRBpCFWMAijt80HCS3IRZBjygJmu9kv47ZTqG
MyDz54XCac0RhIamZIYYtOSrZ8s/bPDBcmeRah3Gqi5HYGmug4bHyER+21QeOz33
niXbvJv4Hmz2jdi/Q1pI2RH02dgYjDFuaM8E+NzWEH26VuRFqRYgZcM92GZmF3PV
mM2TWp2LakkSVF07x8fJVQBcUQizx1KL+Bm+bFQQES7Ih1BH/mTbIYkcXm0JLWYk
vjtFZE2WOtf7HcssumKr8A9g9eQ1F6Xw4vDIBT1xetgwU3gMDcW33qQzP5f5Pca4
all6ZlKD8g33EAH3KGwhKoV7b4JrJDWvzajiWGl/llShnuUekxb2q1sYZm9I+2b/
3LrZSKt5+QUFGsmztHnmxvpXLvqk+Mu8L07YvqEKn1L9JnOjZTWnv0qDEOCTTpI1
YWpmLWYXUNWI1mHf+xbjvbJo2FKCyl/Blaq18HHSkvKbHMZgJZYwRJaqZHSAhh5t
hSxVmUXzqbD95fBbCtXwgpa4jOPA3/ogK54zXq1p8Gx0kgyN7evbsfye9+ig6LKD
umpCuennBO9Py0NIQEmDzzUX0W4HJZpaSfcA5G5Ria5Up4MHmXzM/7bbl6csJ01k
oDsltk0qWg84mKQFq35hoN6jNpxbOCaBmdl4R2BlEPL73pPacehv9TC4R9qM3BN6
K5clCOA9marOdOv0KzUNd1pSjmzspQv/AMIvNlt4aagPs491KYyMtfKHcQ+AV6SY
OdYDThR+sQnfVzD3J5E3qVbcx12pH8BTzkMy3dbFFIdyN3UjHicn8RYcX7DZymWD
J0Dvv0c72TW1n9r2ZImJzGXxVh6/kbNoHkiQC+uBDEpoi19dMRpbBJXmSCy7Xj2f
x7XLWtAKZSSaSyEek9XjThCWzMaye4ewMRyzB0zsJlTivuw3N4TilwTHnd/ChiVB
CHcq0Jx7Wr24ASGgE8tvX6/vYAWB3SdFsFn6tnX/b1sgfpYdzMj7YbY85oeuUl0M
l1O8jVVXw4VPy3zeHD29QnjIDnrHB3TsRkKeFsr1uYflI/GZIEiiBB3lJAonOqNY
TTPyB++7ZrfMJQf1ke8tJXibQ5YsyGLSaFz5Zbf6QzySDnCGt54rNQJ1YoPiEvT0
oRn/tyQGBhvX3V6y0v9tXdWWUjcdt4cyyCu5lhklSgPZRLyp9tJIpZSDw/3fJACa
tBLgoiOm8m8yMgeQpiwe7WrrU2/Ikv8mi7g1XS3SteaJgDFWYqxtcnbH65Ut9hZo
pH+KEv8p0Zj/47OC9/jOWv91cwoQyUNMlyBE83sXwvdArD+dEnTy01si+LrC6Isg
E6HvfVSEhr/QQxnvOG6X+JLuKZs2cK+JNWhn1BdHmOg/jQ0OTQN29L0obCexzdOt
3qHLTymd+SB8w5PEtwEWeGxe4H9tH1YshNg+DuR7Cx+6v+hTa/eJycDC7zc5BqRa
RfJogg8UQjs6VeA1Wi2jmyZM+csgmVCzxqfuZFwy4lb4AkCFeErMbw/fBIDzGv2s
z1VForBJQU+VGiNJEohOdR1a40kEeVAXF3Tu6E25io5YRZVT2EvZLMPBZ88dhVyu
VEL88q4apaVGMymET+0O0D7y1RceFdrpyAfAA/f0pwu8bKTiGxRxbQkjQxJVfQos
KvmSMHVNLdtKtNZSYgRmXdeDuQwD5hsNVHWMuT2Zz7IuSKK42lFerLDkf0ZtXul1
bsOCC96Si+1x0GHRazhAlnSWR2ik7S57ld/vj+M4FlJO+VKFQKJpa9Htow9jnF/h
EqeKGwqR3BzmJT+v47Y9CwHSTgQe4F03iB8gu6w65Eut46d73fpVApIaRx4qa/Rf
UOVoGoPjHC2DkqQc0Q6Uf80yTusqVZ/GUVkoPb+ZRKVJ+XsLc1KtyOPJR8G4/JD1
PS09tuPj9exWYs0NoAtgA2crlRkuze3hxThOw3rWeEfL67q5uHrbvvaWv6DzK3gw
dKm4cqLTECyIsJmZ0QUC6FxjRJWRUUayXgeowGY8yGrQrL2WjoDdskQdhI2hxxeJ
iHchNEIaRXPsBJTuxDhnSB6HT9wDw1wAOASjVL3m+EuA+AfaE/2ZzTWDjryNppgj
5l3W4yfQik7UXLds7FlHtdPEajwO0Uyb1lYI2bMxjcelqIJJA0st+tFAPmhafuym
5JeuhOMcmapw/hcNguKUkZLRmJwKqQzkvu4r3gWUAygHy7QUyufPUDoWEhjSrdgj
8hx+xflXf5eK6SGBBVg7r02T8ytvbRiq1fFXzKB95MxhxkemC5zhBFqWTDl25eqm
ir5rGjLVlk6fXuCehVqVSM8TAWoNB3CIVg0pMu1YVYqw2EdGgE5H1SUOKpAODJBW
krIVdRsh/qVKmLdklMIdqamTS42mjy6FNkoI4kL05ljl31HDrVxI+H3wnpD9hG6N
VSsdrbK75NNGE1AJu5SnJR8efcQSuo8TWGZHQYWzvINP/YYMdjrNbyQIU5dyYXpb
au350TNGPx1L0GRyILvoDT+G2Fc3QwXQUabdwDc/AHvOTfdLa8SuFgXqID82nStc
fsT5Gb//YigO7s8Xjq2JSdRT78746/zeEAMgjB0zIOsE6ymOlIR4ot8vMA7K+Xgy
S5v4k7A70N7/Mnb9Iw0+a5ro9E1GXPQv3IeNuNeOMhXwgTtJ8W/xYHT7+8a1p2ha
L4FHssqQTyJENeTDpXo4Ci6Yergr2rdJlFDYpJtiUWciPydYlQDsYNfbFMGGt3xT
aCNR5bwLR471Icv4sLPC/I8mgdAHMfkohRqdseA1X6cb2JKrPTYaVm+FmGS5y9gx
6OFM4optXEQKdnPZqXV28fVDcfqZphUGM1HgnBH/i3xzgntWdxfILZjM/th6PIM2
UHsfDsebh7/AoE/aDV4wYz6gM9oLjynQyg8CeMIJ5Lw+8McvyZ5rQCSzSnL8EtnN
sLEsODqFwCNQvJQ6oGe8N/Uv0Yu+iyu4G6+4lL2qqmFTK5Z2X1Z6X985sR2R8ojx
egjXVIU9fb/HkJNGVeQVGgqtVzTsYRMSJv6zLFH7cg3L9eU+8bD/RITyIAka11gI
8PUSpUNA88IiJfDSMvMyggoShOe9+z7dXBNErCDan+S3S+IRf8dwWLCi2ylUYNpw
775ucj5YIB1Tok5Ow23NtRzuzJeyBnLyd6jo5dynh2AUIhOZ2X1qCOyXEgx853Wk
r4xpoW/1DT6ZBzOnb1FmjcAjWguRPlEw/sVLBDYIpHoQRoNF48zAaQMvBaVE2RVz
fUZ12wy0RldcwuQvldlPPGEXJxGVGND/6t3etFn+rRSkoUYcgUrNNKPXpYo8wWu2
WvJcE6Nr1TmXn73LJCfM9l5am5G/jnfe+dorqqjVF2Bve7ieLx2G0+i1OKmKRLya
EeZSZZXIANEIxu3dNMYe96Mns49y6GTU2AsEMWqQ5ePFD7o7pMzeknct79jWJqhM
5mu5CZZCQeM0CsEYqbHsR8Y4f78iZobMA6lORkFzQ5B+Hh7QJCmVbFDAN7EondR0
ARltvsUs7Is84H+Yhv/AA22i0kpDl9zQyAOw9Dh9TjxQTkpsCt+a0q3aMFx9zANp
n8j+M0H4ABKLcHwQ5K0PUCPgbAgNDrOgG7u8kFCFRGCVuisuXjl0n0B+MYRLrOfB
X8EzM3wsIH02mwmgnt3dex7BOGfAhh/AQHAK/O/YcZyj/4VjDjiiCh6BFWyJIpDz
MCcIVZ/23ap68CaSI3LgzAfDUCVXAQI90MU9DFooQXr/mZtf3PkuNf9a8SsVZZrp
DZ11AUQWMHmpisi7jEofAL8P3skwyvWgNggAIDNvMqI06JJGvIXPF4WVSfW9fAtU
M8C7Oc90qcHbsq2nVR1K4NGNcToTTkKpJTU+NF0Y1AzJOembP8f/qqS4agshFttY
wtjwFwCEm6HKMYlSKT0ohRyXZuU+KPNyIVLjfxFDp2Op4J8Z9j5v5XJVLlxKBvWV
5uDzyBbbtL3kj+TCrnl9Ev/3t+428gl/UNiNEVBZeD+ljTqqgjc2nzjk/86SwGVD
prTcI8ikvPBqyzoQK5sQg8vgsJIjU/kQ6hJXE7Txs/3Yrb1wuIGmw4BEy+TeBbqb
39Equ3TSGuryqPsAqdEjlq3GS6IAtbYY4AJeCtB12PhEWOr7A0C9pld2dSxoTBhc
Zknmw7jZW3HKe4Bqip5xl2mumEHlIzAVXOE2MLesL5naYYDjOXc+j+1v9HZuPUxg
0w0kf0AU+IwE9ulU/DOlB6kqIu8SkOqc0CUzVBIZiombnRKXyn/IC4rliNvANsJC
rmuzcsnB4N7GACzLH0toqEmV6Mw7YOTjQscCR3ujOW71ZJ79WV5KX9ahgwtdZkZ/
QY1JHQxjleGHU01hYeaEa0FzaZ6GI617+opNhQezI6gCjxdaiiNy8n2GZ9b4PecU
+5opgxBC2PdC7NygfR5razSqvOUmEGKkgialjv6SmSQPl5lZNZE137jWVA+XpT+7
6RHBSZTuXRe8wVELXOABYAdrg11hfi+joe5OgeZ8WYCvw3/HmOg/yT2+kmikbsBE
7EdlZ5Xyp3PrMHn+mA9e1BnLqriYEJeahMEQRmK3lKCZENBJBR2GQojEodZjq6vq
pu8+6DEZ1y+a9uQS8nW8tEdRTmJ3oB5c+/uuvudyqgBM+cq3OiLveqHM50Hy5V6f
8qmv86qzkwD+zOCdEr2QyP66bmJJrNsBuKle5lOCIjwYRDYZhjEa/x+Zgae+mzO8
5xsxFfb6WvBr/qBL5q7fusOeY+ORqJfFG5uJosjBwSJyHq/xJ3xhJ2/SDMahkY60
+fOoEEQ9ulLTP9zfMYMIcQHGt99mpdoacKftAYa0ocf3cPvOlGjzbZvH6wLCnj/7
XS8NlX3w75l9+Hf71vCgGCX4rdURA2ch8ejoUaXgKBtHn5Rims6aLr5e9cvXYZkx
vxlgDeB0Z/9K+/iamkHapEvo02FNEiguqKYBEua1nMbSGa0Ftpnks4rBWwlTH9We
CgwN7TPcrpGIbwo97ivH24AD0By/HKsQCSNdVG5F1f6w81D9wFp6cCk/fNR6ZJub
DF2m+5A1OeshpFAd382RJKx4BGQ04kr7SnYosdXIKxn4umHlpSreCvUMzMh7z4DL
+zwx3HWL0LCgz10a30G2oukpzArCSBs4l7T9Ot5oLTqWvlM4kCH1nmyZGnC5uX9V
nxSZguriqSKr+tokslwLIAHoxpes4V1qa9/vAFb0u2paC0O4x0Ow239VlRo06I+1
6+BJhOvcJd9jkP07/QopixdpTgStVUltslwV6gumJvTNKMhO8Ik2FTckSHC6jFpd
jJJdHSZqY1m0XsQIr7Y07DKdcVHqFzgZtCBkMSa8Mm/b6tCwjUEMAla35nNNbvUQ
q9cViH1WYSsyB9cxGIPBWEQHwpOYIFVl7MysWv3oYt8/yYhTahZu9E2gpe7MK3Op
WKQDG24fPmsqC88NeCqlzf83dJSLNh6qokxfopVFhZtv0NEyTt0/5xcxYIFZgEiA
TIg+VpgEGZ8lVd1pGSYoM5IuwuCZ3DPzUPG09vvEkDis4+BXQAAZn2poUAuJ1X06
RDTXglB6jIYH082MTZljk4reha0uycv9PqcR0ACCX89wU+SONqfzIqI9vYf8VwN6
SSGAWLE6KtJQ7OpQs6avKPv7u0GCH6QMbCfdzvp9+QsEjaUBUaV1V3Fh1mmTiM8w
A2A3MQzvagGWHo+w/h5in3EIQnAFyXvQNMrR2WsKg6MgobndQk7OZemtXdFe9XSO
ipZ+tJfOHP/QDwbGcH4t2Ux+QfelPJA8Mhc5PYJANbIbWzJN0IIqI/lAWZFaBSAN
d5MugQKXpPTQ+qrdttzesx8mcop78g/xnYZNxPGPTors5D/Yl8gosWvbu+8sNbFq
3V2DjV5+fjcXcHKRKqS7saIVQBmfQPCPXNNsNdmAY00Or9RmSFmuSzi4rLkRJWaJ
/a6/Fou++dlWkN7K1WdS+ZHSzv1XLhOxXehSjsVW+zlU4hLujJJg5hbH+M0AwucJ
l6cGya/tBJWYxoOGFPjzERcoCPReXK4s0O4iYmcUk8SO5QcYQCLKCX+pjekTL1hE
UbV0kH6CRnQWPLOtoQRt0vHGEm2EmFKNAv+xozvzIUF1ZXayxJMYTfUhbl93OQMR
OiLleOm4cywC+FQD0hq2tLVndIMu2FaLpZ+t3wftvPVZBAOpXPSs8kQUaK5kFvih
O3O8qkh97Ic9g+1WbySZkweGP38eVfKtVC36t1zG7ieaIimleWiUNhmX8RU5RDZx
crSUGrCGo86BgNkqIxDNqwlt8k+YG3skS4mXhkE6CWP6+KZ6csT86Zt/H8imWSOc
wGH9UgSKHGM2cCG3IVqhStQO2KWGwQI82maYxKuZh79167y8lJ6hinLuujIa0KmD
21cjRhP5RWlcdifO8oqRkA7+AA6vhEBdyM3ruM1XNL7/eAe+bk53zjTJDQeMPnKJ
iQWMeXmyoXez4F7DqpUkXhsyTZl6HDq5uI8qLvgXy1LD0vWytp/NdWWcKcLk+hf9
kvFq66JQ2AwVTTDMnxrSq0k7SHRbO69UOXJJhgOosnCPxKNIc231YDbt0GjZXW5y
m7VuOtmeH9jaTgYdaghtjrnKa38LyUPwfH1HFrzmivScUgQ7m4MFoonUApG0yxWB
zgAMYKhWbPF78dFdmPwjcVmp74sMZ7AuuYJjLhCiq7GzhbAzjLruRzxPZJ/yE5G9
BShypB4mSAHyIz7w8AiVneUSOuo2hiYPQ1NbhBHJ2r3i6qRwysuMEoXTEQw7V3y8
vxuVTnjW/CBbg9nJ6KJ9Azw6e76fAxQfzOGzWXaOtpIDruC2hEh+9w3Lv4ybWkrM
V0vIJxUtXUMDCOw60GzXnDm9UWmyl7pjTOwyIuBH/bKvqtk+KuOADukcN4QX8w4A
TUHgqp8VI8osX3i3HB4Scq5tPF/gdDxVuNAQcWEmHNmSSSuGm6ulWlyAux3/5WRo
Ltz93i6PnYF+67El/pizYB4AXPWs/CNl2B0BhW4A7FvOX/1NbDMdHWZZUfzWJEUm
wk763U/uUxprcXTB5z6tn7p1LBbhl+se/DI/cADnsg7gt+BYwCZABxyxtNfdtGzM
4mNow3PTfq2iJEFnK3eliK5usreQ+9hLoSyKo43IM8cdV2+feX7Rry4gjjIMLYPQ
9LbJlLA6+7q4hhAC736DttDpGYGfznTyVYai5FmpqdoBJvSKtiDgA4VdXTm2v2M7
oMuM3pe46dkzhfGho9THTQEqhoYxqk8JwZLHZ9jLM6GiQOTSdV5sBVf+FwQP+9JH
JMBDFtv9SHWSYJ0feP8KNk7dJicDJzkoPR51nyk+wYJSHR1O398TuTfIMUk19b3X
eWZrogevjb79eK6+wE7CQ/LlcdvyTq0MmwID5OVvTTq4RT4mwhXaPh5mWr17V7+l
AkbKziqgIPttulVHp9UFoZ3kT/qCTdmhlQ0w26cA1x7NCJWsbiMwEOU4v5r6dXdi
bxZIh2Q13rrWNyfR380P9+ikS7EEQAVIjdbiEjnYG7rANzdCs/1zcIoz4Fc9J2fk
GtV4zOvM0ygJtRmTYbjSGfWAPA2hBWe9z1Wgx/E9v/5Jhwxfo+f90KQgwUvltzDZ
EPo/U99M0XqrBI2XrIn3nid8p+63gHCLZqIQzlAq88a71Pg8zVG+WCJYMAAsR836
UOUYPtdELD/Ah8tEVX8CO7hK76WTLv67dstEwAx5nlRydOPQA5CM4luQsmz8CJCd
fVXD0w5KJpX49UOanQcMLROpsuDs07klQ+t3M9iOXkRS6J8WoQXLDKqf2uOtKLvC
zv8CKn5YByvgbgVtPUaxXW6fjr3kFuvSCSHmeGQy6dSlt0wjUHpefN6KVMtGUhCk
e7fhGXi6eEe6DDVQG01RivfWHGxqvZDFtXk92IS/HoB8tVJif7LV/URn08WFGCpo
uKAPI2xlESWTn/vvA9pS2Mi9sJpNcRZb3pYuL4ARJHvW3aaP525RFEQRsjMDq8nT
lRlQwxeUBJPt/U0iH9GOppK8+N660w9m+ZCUgbI9CRLIa4ajSzYXWHliRPXON48y
Qfv5mva7P+QIi2RVuXAO53RCIZ8TfX+nWAKG2XCkMbC2SJjcT9fTe/rnLoOg/QMz
Eqr/3xgARS88ylI7CAgrPdbUao7fqHpNuEmw/ESWwn4ptI37sj69/5ZWdBMukxQB
fFobCXwXnTNbhQ4943wf06M+T9dPV67/vWitrNwKvXQ09fyLSg18N7AgQQZZzFlp
pxSp4l5n4Tyk6QBtg7StlwrD1lpq0neadMGnAy3Haps4Xw6zPjWwAPzLzpAhpgve
UyxCLD2qsYjGoo6uoBkkY7RobufflBFT7YSptT0M2M3fFKu6zb8x3a8RTQu6L/jc
1DrhKx3UDa7Hvcrpc7Y7pdkXKajBJ6cgxVJo9Mu7HRatuPrKcr8NCYrTaa/vA4h8
ICkVCCaERhXA7DeuXNCH7gI7FNpDbYM0d3A9vLzuyUXFTK38OGHAkv/yUB3hKtQJ
6NbBmdMoCRXGel5XnM6nfjEaMais0X8f4RYZ4AJTrIV1siI/2qQmPmFttq5ORd54
PhyP4fZdWDu1mxOMmKC2ZUU2gq06ZndikwKlny0fBIbhhvNhH7dDk2lyIsAaYYIk
qUEj204wbmRtUdeHXmOSCA41BPu/dqUKLvFdWgQyTHxpTnFLLS0qk9HQirTNHwYN
HDsV436J5BHcp2eo6oS9jntndXpEzJ6ijpqbRUwGriZDraG3GWrhb+UJkW3LVNM7
B6YCtfEhgsb3EjfbwpaP9SnK4SQG7x1O4Fp09/tub+Tn9Q2cee6de6g+jcgazJoG
XwJGKVY3osLLtBZW6ExoGD9J6PdgKA6acjjp6316lFBX9XD137/KNoc754iYHOb7
JyPtXQR3CQOTJqksE7Aq/kh82MENUgADownSClkjLN3JBLGXIVEliGgMPpO1brkc
Z+djtPMfgUqbw61zPBEdwkHdx3Mx18JRcYnk62oRLE5ZUYlANbVv4KbLTDAI/3vq
Iyik/AG/31EVDcI4Z4xiVKqjcriCvYZydszUFWcgPkhQrmYN21By2RLQxLxW0s9u
K0Fze7BZexntJQS3Lhcw58LHmKVOfn2NqfQOIHviBRkymLKuaibO+t57eyCf7/MF
8xbGW3MZTzvHGe96298djxAUdao/c4iG4V5uyMO+TIN6dkB9uAFWYp/r4p3Q3peb
4opFINmHLYPpsMJMYGIkm7SrKBKgplIhn+ZNIi/w2VNVmwyL88OIlXDU3Tb3Qtrw
9KeXOPVYxfJ98eZY88SracDHTGgSKY+FNpxvdaMPfjkMscUTb5V+wKTivWSbwv7+
4/VtijBW0cZimBAQQbx49YeDLybJaNb6HeoCVY7LDurN7aa9lNzrLFo6nyq3iLBT
rPoNfcu0JHB1Dt9UWGd6iMdKhmzkqIOZobLgWOuSCGbE6qYFPnombMjsYrJ8cbrk
KSKHkVXQPN2HSat8v/+uu5YGIuG75zJpthOu+DUOnBYxTb3PCr6ks+M/7zZa7Ekf
EXpRJsKyPUo5pu45ZrsQJEQQ49o0pQNO6/qcojTgMt9HIE5G083XA4EQAuxY8Vj3
cr9Vm5z3i8YF7vU+BA9zu3vl2+QpcFgegIar4wOsBvcOOiZ4kbq5bG+jh0mm1rnP
FkT9X7nxHB4fyq7MP3KcTCu0Kl8CkmbYE0Ze4Ryy8OKM0ZXV8TSdpFnNhgMhbUnq
XVy45yplBI+2cow11z58LDxWiDQ/PTvwuvAQ3GP9PX8XdLPpVnxXkgL5f3FNymJB
QcNOcKXXyHJBg3VnmJW4rhah0AHVHx/bEfBuPSGRZfkMoM96k7Y9Cu4AlMpqbznC
DsSWVSOcwxLDMv0J+tOF0RiU+66FpHSj8/PBYtZLEq+sHe0DOoUPHmcZhpiJlYfC
vtrqTiq6MlLe5V06DLXORCeA8AOl2Qa1s+bgcJ7focA2gJcReS51fuaBcH2zjXY5
XywIbAKFXyaxZm+ZYwHFu4FlpXfQieINHYVeoO8hO3pNAvjfpji/CwNmOPn00Yjr
PzVqlXznp9XfbvYmNwYjaOisuxqBhEGwcN1DXT4Z56iOpMI3moJROWSr1V7IaV0f
vvubxox/CuieG8VTjxBSR59yrdJaS3zD3O/INwvaaE9gkuFAC25r44gzXcIHuDPR
HGI8aK5l7ER4V6ytloghHUidk8g/thnxgjFbI8kB1XMgqs5IVJiNpaOOv0Ns6DBr
5hxgPUz/leukOBkCD5zJA/UGIlJmqiwrCLqO2auiWv7qudhTXAoUUW1HmAlY4BpR
n9F01hoNoSiTzhhkALcdF1N6r6xlmcwW9nguhNGvs4h1IdRCobAyhml7bpq4SIxM
SdZYiROPYcM1BEX3BlvXsZiJ+iU/6VCtg70vptUUQBrCpk2+z12VE0zXRkHYjHEA
l8P71NN/NzzWqKIxD6MgAmtwUw+72yEJVwL4TGB2mzHRt8lPuKle4SDGw/XbzJKM
zjpBBVp1Xq3WAsCAVkitbcdIKWoCjCjKtbhP7wfq1Q/eA9BF3F2xhh/3NzT46euu
jGCE7IjP4lxsYdL02wwpfZAHeTes2xCAfhKe/awyc0e1IrNvUwySkjx1nXfqaZ5D
6yiHavFejx8BLZbhHIIo8KC04ucW48ZGJlImDFgIWnnKK72VVCMnLNnbm/tPHvOe
0AjLvdOBmEnzH4vrwAYr17Zoj19MPW9NRVQPK+PtmzDCKeSXl8fXBVq10LmEDB7I
4YJae4Vkoh5/QBY0D3tpyfgODOieCT5bzm9GEqgsMxZfZQllGcu1ReREiREVKfxZ
MI9xpmdKXb2Mlc7vjop+Ej04dkdMBQlZvJnaxFH0fdhfABDkBBl4eFJRLLsQL3/D
zepE0jgC5sIZQcdqpBjjqCFRSTEgQGUkLnp/48NmEcmzDBdXARPmnviiHBM9SytF
6KPupSucTsJdUNdYG//ntyui7geAlVlVSXEyb/eaBitwu3B4IFKfGWh6qUFPB8yq
D0rKCN3devN+npkit07oQBb+1iv2WfSA24zW755GG48VaLavmb91ydYlJ4EnjxK6
DygeckbI3iNAuEADC9cteBafz50FyG2R9WNgkmy3RDazW+HIIE0xAfy4+QevlOLD
03YArJxLJEUihLt4yI/TxRaKUOMkeczv/oKYE36EEfz+IeI8qshc1j7oEl6ppHUv
V1m3I83wZh+x/B3L9jhB6w==
`pragma protect end_protected
