// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:20 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mAVgSeDWZMY2r4+HuPL9s190F4FwX/dOGiQVkJdSYnx1Y9C/wZzbf+glNenIil8w
udafCK4Cnl5c2vxJuQxaTGKtahUYB6m7HkV24xPp4qZiZmFatAsVmTXfUu+ahYQD
7RWnKIKOlSIF2c86WEfDbPETKYdecIb0nnpftWIBMAw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
ClMi16JgcTEc6f8mMi0LJG+4j49voqTTFG0MaqBvb3MTN46rAzbRYL+m/3L7JF3J
URQFJd3gYBLGxqlvythmr3onkIpHughGvguC9GIq+Z5LCWoxUhS3QhYHwSvAeDe9
z5l02Ov8UUDxEbVqPK5wDnn9lt/l6OubSS8g4bkwIKdCwzokaeLFbo0cm3khnd0O
YUppXOMes+A17XPXgmgVosxWVLGjfAnEcB+qVTK+cvuhYG7q9NWda0a5q5/i1A3J
nYIqBvIERKRzl51zjqxlhA/jEz8acQhnIlyHKg7vyyt81maYr1omrEhYcqMXEERy
HX+Z7jcVkjMk9DfQld59H0rDqDdtGQC32yVI2GAL2o3uyeYfXb6FODHyRVCv7Kq3
h4xFbv4Wy1tA1kOZ+C/q0nX64pP7I2trCUL0sc3iakD7tU0xIpsLLycFALS8WCHR
DI1XEGnSUt74mjxg6cZz7t+gkLd1ZHvFlNd+a1hjcYQQ3v5xW/RqT05W1/oZTQND
OcHnfgmIDNxq/VUYSUy839XLCoi1WQTAh2bt/C24MHsJRwuKxZ52hi/+e7gq6mEb
dhTZfvvic17Vj+dmEbvMRgguojy7S9lFAgedcw2x4FWOH2YMlDGEfNYcrhscPzJQ
jtJnYiX2It1Be27usvrU2lnDeyBqW+8w+MS83ZUeRLYWqqMQvn7tME/3cuQL2BeP
dGNexkrh6n2lqxvsuOkLXcaHCtNgq9Q3t90pZXSwaJTm6wSR2lBh/KMm6couA0dA
DwhXvxw6/kosljAC57XRLfcVtqhJ9eGqdiEdCcf5WnOk5OvwK6DtqAs8DqsDxlR/
YfCVHcBn1PQAxME2cpkCVKXZPLdV5L0RDwR6D/aMMNHktYyn+7PfFULsnRxNg7Ix
0JhtKDu1UZyGbwqRkrzy9di+bqk+x/pfMOgLSBa82c//rw/DZIb5u52ssS54OyZu
YBhjV0zIN904jS+eKJzCWpZxl2P47WOnpNXOV358MUYGvATw+EKW4EVv379mhqr2
kCpRRAg3FaXFUy887z9y5r8tEokfJWZYuidOtbqb7upETEe9lp2HxAyE4tY7Aq5d
oDbFdJYlj13td8ufywmfBOrh1huRZgOXi65LE340+PTEltoCLgvaE66iNw5vIcgy
uiVMGWSYDPbx3OSpSYjYnUlf5gIjQs6H3bqi7uCSju1jEGvRvs9JbCkKW8KwVpV+
1VW+V8HS1s3sRN3gxk7XmW/gCZd7BMHO+FurgD40w4CRHHwrRHoeAxhcnuVl8omc
EtXcLXBz2Wk7QQ3xcrNURrjO3+YyiunWE+RKvYISS9so9/ZVy4XnjXpFM0Mzc4Fk
AkDDXBdhqKbQvMxypQUxVI+lnYUVWug8B2+G8ZSYvQcet7JUwuXKmZ48vFSNYcaL
LDaw2J8NA0UkB1XjgU89fxMvKEUtCnC4xbZocyz5tX1lnax0hMqW+uL6iQiPRgqC
h/WFM6QQfsrrsLKWGaJfVzPoW7h/HT0ZOPzyStBIhAV+nH/hsFUUYhPEH84/oUHZ
Ku3tZ0Q7eTjObmZnMk6eTR9/wgEdqm2Bjjru0e37rgGZOOeYV3ntJ6I69lBCCDeF
JvfRcyfGz1W/JYxvgDdExJFYpyjvTbJbhHDH20Gr0WwDeTH0kBiQvwfs8oEx8q15
+m75EcbBDUqHa/C88SgtAcq+p0ZlOagqX7Bfg5I93gRMKCGKTId+bJcXlainJDuF
O5cJzmmHxfGatq92zi0A2fZ6GSezg+Y+Bv4Yiinrmedqmq43CSCbs+65cag5ZJ5t
E4qEeGImPDU3VpdTNCL8q77G/ST/ipk4iP8T6Zhc9O8hzglF4a5BsjaWGjvWOiww
hRcY6K2/h5AWeDAQ2G6WzTzL30xpvCuNa7dYV43mks/bytnSpRb+IcAAXW3Zo+Qs
cGqTGTeXqkM1BHwFbg/dWiBxqsNsY4PiTUa12ZA6MpDBj/PQwIDElmfjmWCysqE6
ch3c/O0Yd+ZFDf/uLhpeWBVbt1jNcL1ew9/9SS7QKhOPkDK5WUOZhhNR9HgR+V4G
CiWIKNmd5QOpeyg6Oy3E2m0lI0Yb2w3i6KBT5KFZYTlxWUz3XvpfFDhzySUn5JgU
rmr1Q0pK98Gjg9mu2dGQTcbInu5y5gLAIpM4W+fjXt4gi2SCIdH7wgoJ4jv2BlLy
na2Cfad6g+z25lP7+8Oo9Tgc/2qo3ojvzrD8id9kVRCw5E5ur6bT/isrR9XIwJVl
I14kQd0Wg6wsxuda4tcdipuvx4S39hDt+/xR62G98dCAzmxnzVbYzg3TBXuACuXf
cmoTuNHGMNrGkthZ/kNK1Q/Vi9HADFE4Kx1XtwvvzlG80+AFGV9cL3M/u0WvaKtJ
ZAd2U1psdG1X7CCtrhct5OSmddtR7ibEzxP5KixrYKzqx7zIxvrBTshaQhPqbISh
ONo+ZZGJrKDOm+3lwuxDxq7SGAAKkTUBVWEo4sfHFfLMu8lr9zzEKn+Q2DBEwP+8
oeFs/3I1pN3DKc8R/MxDy1bbjVVyaI3sdfuvYqvnsMRzcqqpdG0LO628BIa4lz/n
gzKGJ1oxw50rZVz9Bj8HIqPP4Rj9DmPG3RKQAuO4CLJmetzmoJ0oFBkODblOmyPp
n51zcui90LfUZfLLd2jo/0Caak7JcpEF66ULLJBgP6KUK/Eyaz28sDGRuzx6F+/H
07hJ54cbIJHZio0II0lscFZo8wSsiWHGAkcKx4dvli29vNSan8IuDokZZShas5vH
7Y5HVSsPt/rVnu14/PZcWoQ4xnKwwjyxPDaaqd9J/p+wsSHees0hKwaf2PQVfgC2
7am096tasMj/aNT6dZkmPjADUkFdWvKTX1ME1r0AXU+sv/xy5n0VZDevOK2U8ZZB
FkCmaZDdsM+UTI4mdmtTuGbAr0GVfcqinbsP3qaqxxAB4hvtaGJMya8yxaLjf64L
wlv0ViOyWOi5YRZcNkdqCHce/t3kog0puUTOSr9G/Kd1IXxCBMw3MARNG7W/azoq
1ayyuS3hK0JWk8UI0FMN+F4Do8X8goup8U+44l5Zc+47+jhqv285KVsxqG//gCVv
6OwVztVPoT9hYg0iYrN9y92gwvaTWmfX5H3HxCdbr/gM/a1hvS5pVtP+s9RpJIGb
4WFUBk4BYeUxG5axn52bNQ2p/OgR0L0JvbeCFY7fJzlan/YYY3+mqKJpmQvZJE0h
hodAYR4B/4pyH9EDWyq828KZid2yFNBpNkGPq1kXDynUSBHGYBE+eIlVn30HxJuC
/WhXJA3jY9fMqLZsTPKeOfYdgqnnb2CoqiCmjYsFCa0q/Ql15GzcauHPuR9A22Jf
Pr7pHqiWIc+pMvF/Xr2Xc5IfDJp/7bSut4xyKJOn+8htm95X5U24cYRke32oBxjI
/lRBNQDT647BzQuL+0akYsDmnLDPAsEvf5oudL4Tbu3Acem44nIJxv6M5vFuakDc
H5NjApwZw5GFDBgMZtKoXvnUogZ4of34860awiFmBEdvQTqGiY5eFgk9QSUEjgB4
Bx92fdNKxWHLgDKVTjUWabyj84eOhyJPkipNvafEbz3L9X6kIL3L7PnzRKMx1jXY
AcSfbzKtcYl8TNyX9iE4nhDC8gdM/LYST4dRmRM0CDSFHu/It/08AOshvqqkk25g
5ww+kuosiQYC1VoFWJsAHe5ssFVVTHF2vyQdp4GJ93/QwYb5ogGlLkFdWW1BDhnx
372xjMaq28ZpeD8XvxmijhA83oTlc6GjzlHBH8kE+UrxTcMdNBOLXv3250K9QXYI
BNLOuLB4fCMzLd4dxAEQxctSf0B+ZoilNZRRe7Z3TSxmNH6YgX7YQDMzeeik9E4E
3IikNjJ6lVpCdiCHFKGU8bTsAgnLLseA2iAFmzLu807+JoU0/mdOOmZTPv0z5AqV
apJcZeJOPqs+XujYsdc1ByYyLMGU2nzenOpwjhzct+mNPNAITvpiq2gqPV2pyC5/
UGL+S3ouUVJzeu3TurJkdfrmRH83kg/Mzmgy3OXgDgOMpf/n6P1F+uwYgQRoFOhJ
ssJefTP6h0gKoxdYPSXvgliR9IeUk4kGdCJikHpj3mQZcV6Gmnnr1rqBUlJejM43
Vi5LxHiOkUMM6UyO0LY4VPlbOoLUD6mxbH9/f7P3DVOiPn54Si+PB1suqT5wGHVB
ySLhsB/mtbidK3pqKPHO6Se28mh0DsdGbm0jDH53FS+PGyv6TQd4Daut47H2n3GJ
BT9eoaIKreo5TRnQ7g13xpyimyKKk28bnCzlLkpR6XxFm54jk2SYD/BS7NMEFmVy
wtbnhcktBAv5zAAfY2MEkzOgssuoDwsEth7goRtGImDUcyvdGxLTqnuAfP/uRa8T
mHSoTc4Ekkf6slQJTJyUyYuqVMa0r7T03U4df7DKvIRwxfws4D9+pcYKqOxOEeDa
P3ZbaY8UgRxjDK4fmOs9uAJ1G02fTWUCR+h5BHzxc0JbT8Ju3TNhXl9sgVPSalOg
GCDeey4lTiS3/KQw8iH3EYCSvE2lS+Epr+XyEi5ebZZDBu70O0fwsHYigFrkg2Jw
cJV1yIeibv06t8BzUacZI9ClxoXe7GHXpVjIAGiNZgZayu+CNb+TS3cMKEMpehcj
Arnexvwq7mwUxVTaaTVuG/ANNQioWSma1A2Jqn6PKVznsDRbwnVqXl1yqE7VpQH7
h0+/yddBo76sokphvqZ26oXHS/Yei7OaFAAOOvV5dZZjgNxE+gZElkkkPhkGNdB8
x7+9aOeVFdcIyhP9Wnnp011FAzkY+IaaLU+LI4ShNbYYD/CgU9Ek4EWxN1cf+ki6
6NyU+6Ku+koKF8ow9yt1roJ8r9G/38rBYyzwaeg0mybjYlxnOa91fmWzCiJW3bWK
yBH4NKRYsEm+k/hbgvRHtbeSAvj/hzKS0PU0498vYVKj3gbdDNAIycZcFNvjVtcO
Ck2Fvk8f1XjIzGOerNnlKXo9xtIVo+f2DFZoDTH4E9PSEKBhVWvvoOJg8hfiYSK2
duEvxGZcsAoX26s2dHcMr79pYU931JAaA9VjAhzZvGZkuad2Q5Oe9NPOKTsvUDDV
IyzbvBJaadFues7BjdYZoHJwiBAXnDxTpAJiElGy0QwDFlvjBPg6VGopG5JXnDHg
4kWPbZDH21vL6kiEXSTuWzaodPEnyrOEC7ekEtbyIHbvW1gX8FS0/y0LNNs2Kafl
0gNiUea3baVv1gE+bj7TNi2IS5Ji1kweItMoyMV5XBsGf0jkZO+Oc+oNBN4hfBQj
RAdKYEsbYNYlhHsxTdNygHHVTp57Hm0HBfTcyt01qWVBPe6NXUGvUH04xF+Ln+zB
Fk92CttQS/NqQ694mdFRPL29yUkTY/4Z4jUtRfTdyZlnieXbuG+Y9OjGVvW8qgJ5
bQgQXKaR1BBNdg+7GLCNlDIi3oMAOIitvABjol/zMzW5TUj4fM3K2SJEZTA3bIOu
3ISv+w4U7l0rMxzWc3dsUyc1+QuWjbut8d5uUUq9PuagGCL3b1eJGXs2LOD4NCCp
tkkga2zsazpgKwFbVr+fDXt4f1f2EhspCZeGPKimJTGWfE1hLi/lOyjJbOlYYNdR
hkBt+6yJNSN00xbFCYmmOrOK9HSJ2TVYkL+ZCOsQPQ7Z2BLkloB099MudprijiOt
8PSoeEbAnDsUnBRbtEFW0cfqvGcoX/sSK0WMezAwQ4mC0ZQ/3XDEmRFncjU6HuNh
j+rfa8nMF4YhOLR1Y7rMCZNxTjioQriaXZjyoFWH8XKwgt2BWyFIw0/RR+4Wp+3S
HSECrgAEcBJQdbCI5uM416vxCzXzorfuc6OzHqauuHzyloFcw1QcfsFUMKDW//V1
Tquu6adPCAbBYXcR7yewdkQYIEGCiwjPiaT9kSi96Ysh1H4zoWlqACA98jdpaRuw
AQPJ22feCsSmMjx7jVasGyJReupln9GRpYBP/tXQi6Lm25xR9sP06kX6hY4YG1F9
q4tXYyyEpH3bA+pYJQCry/Jbpx2a1bL36ZhsqH8W52NsZZtECT3yGCN0AbdzCqoY
sVQvQoBy4YuisLJIRHy4IGe89oe1SsZerUa+6nN7Djkd0KsEEn/ob1+bHfajfrEK
eG33/uu+kCayNmlTLOqSv6ju12O0diN1jCWcTAA+WFy9Qc9qRk2ySEH05UHTtusY
Fp8BePgVJXuObUGkGZOzjlE1yDa9nqRERJYMXWTMiYmO5zB5guHGLeW+7ItVtBrz
wrxol4RbHwjiYUasC8w5XB8bcqn5ifSfwOEp9sYbx0DG4H/UJ0zLNIa3Uo9c7iOQ
99pUBeKZy+aKhDvGnim6UVKxD5vB77VlDkkFwTUK9eygIeMDNwtneAEaRxVJ9ehx
pumfj1BDnOC+H1xcU07+/aMJq7aSo+UQw3FwVksaGtVBqIhkh788/oZLR8MMZl+K
DhyCTWmQndYwbJxizOMRE4Q3jMC5mhkNjYBwtFpascQy3jE34x+teUcxaI7/5vcG
mcP2e4sj0WyQ1vTwq4/cHsGrYxW+s/l6mkuICrbZvSNYoyQAw4Lnv7KLh35WSUBR
jfdCvy3UiQ5DWWqYTU/ckhDJfAIo0pjJfP0HH09plAxnc/XSWCx7/D7jt7YXUnLE
G9vO6s1DcsAZhxo/raJvGQjWG/6Z864Onx46HP1QNH9RWC1w8FZk3Zx5jRrPrJu5
yTFda/FWXkP3xrL3M25jIQTDF247crZJvCaC7fWU1Se44s6roFOB71OoedJREczT
2ZzjCqvPQeV2mVibgEfREk/gMrU3enQDNgr1rGL1YAzcpmdeA28f6hJmj24tkDtH
uiv0vvhANAYO2TVYbOPrftXUut5Wp5zJ/Lku7H9l1B9KJ8wSqPOLqYto3snQq4/h
pwHMZitGfywWMmlKRAlHeqZfylM2Wbr8VClQiJEakBWv3+NVgs7HfyjSahmqOd7T
2+p5+CbI7Kh8uFKSqqAAuCgsOtUqS/wQvwz50t3zu2Mm+5UgW3t6ai+Xy9l5sWlw
hMCoPWNpSNDrpvXvHUj+vdFA5NLRTX+x5B2DY3QcGW0YXAjgcgfYKenFn2ijx+7V
YhJbXV3RAlSSZM+48mYZM8pqTE9uYosg/7BPvIKsLw+5PDAOyxedYnB6NouscgNK
yag78Qw6LNFQXl+0ZBE6LyG+/bcBcx1So8+rJ7kgvPTCo3O5S5T46psYUl5VfZFB
xoWMw+2UA+J3QRm7EHOLCEGamB9L30XX91pZ+ciiCK9ARbv283E0s9G68NtoYt6c
W3G0z1HAI6sRJPQdvb2kvZ8BjqxLpsGnnD3g8+ZPLUZ1k+9fKjJT6bQ5krvtvFJD
31kR/YRzRbMJTRXTQkXy1v2mdzG+gsR1EUvQsDIxdfHwCqMQXJ6nocbHC3rn+vaX
JMaIr7We0kySbawcsBP2zUOJmyjTB4enUxxJpT6n/1zyaLvFt4zCFgk7YUFzDm9F
hQ4xfDDrIvb5I42SifLgAVyxBvGYPUECy9J0fbA00T9lclXqo57ZLurJ+z7jCuDY
uVMbnWe4leuZUNsVxR83yn7HYlan+A+WD6ebn8rFAqyeDShOUJt8Bmvn9yWTgUlC
jb8Kr9svLAX24Lku91xfNwwlYPvKKAJbkQhTMx3PX+Bl9nNYNvOu90zsOKUoCd3v
FgFejMF1Q/25t2GRCbrhtLo7wayydgezmNmSEqQCoZVShb6zgsgzTm0ATXKimG0O
iyWOoeioZiTNRP78QQ+j2e1nGalHJAL/lkIJPpIuorXgP0VtpR5HbLRIY1vm6wH1
u0j96K3/dg6kcaVx7+ThTUHMGKC76MA7xWhCGXeGhC5DDkeDMi78HCTIclZzKE0r
5F/ImZCN/vHJCR1sPVFWEbgb9eERGtWixrg6VQrmfKFjVRrFZFpL/AiAmWIxhXZi
pF+EuOVEMONOyYBv99yibcA2Xv2xJ7qFcnLb/IVAiN4Wy1eIxEZ22w7F/QYSVIvC
L58Xdx75HBmu4Z5DldaRp/Ks8DT/Pe99kLPpVsyD7d3Mh/HtfLsC+oGarpogDHyC
Jiv5V2zDaGwCPTv/5yw64xVu/rZDzPj26M7f0bHI3KE0QSZOcoONghIctxZBbxn+
8JQnHX/GCPBSUFpiG4bWTOFxaoXxe4OUIqyLAscsPPTwr+2t8FyGjkDt+CbtG0kO
WQmaTDdG8g75DKRUbtvVLMBSFulEyMobAGRgX4wY/euDuyCpGG0Q5mfLswQIlUDa
mnsBlQXKSrvrFk0L+9fSC4iHLoB8U7nzOHMn4CrtTsNzjYSmKP339U8yAjw5aWpu
Tg4i5PPJmBBLRZH9NmYh6cGesxQgFpuisxUDnsg7Cm0SYskUtGr5jA0NBmtV54lk
TQmaYiYE6QENX6PWKdYKrUN/WXt544jcgIyGgLRmTAPXnOdKx2MzHqsTtwVobRto
pay8ufK42zQsd1shGSkO7q8XzjPIzcEnYsVHV4ZAoooW6Ywgrvu9ABHlTGX/u7O0
`pragma protect end_protected
