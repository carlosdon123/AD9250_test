// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:20 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l19LVkaNXet4wY2nV6Ar6thiNiD2FO2CCrj5l2Q2jzSj3nXLA6ywQy4wUexfOre6
unmAbZKwjDk570YoXjNh6MBJOqFN3BloOeQy5pVcVywXnW32qDlpAIuP5RW+w4fT
sjLLsJSgqMpt5bDMiBextrV9LV8NVdYk8g4cC3bKpiM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3072)
Se4R+d1G0N1qJffsny8W43xXihwJ4KM6kTfktm1DyRz8UEqzcBSBfkvLgK6JWhNI
9yFfb+BZlwr6D5R/398pFMRNzrNrJqrllxhFMb1PlKY7I1TEP6hpdpYgHVK90pQv
CU1+3afx5lDRB6Rao1tbQ2FJpoU85r1MAA1o8Bk/dR5sJkkgzk/qBcnavSXTFlni
hKcxdYJ8s9ZYzZLZnpVEw2rXUYDoau1eQQPAGi3/rCAipWZ9Rza5bmXQKXKRvOjo
Gjh56/hxVFfHIJbaOSLnHkX3EPthJHLWL4npoKIioim6aaPkQO4wIYU6RHHFV700
+XSJa1g6ysfOZPdMjWSb+VhyU+EIhA19P+4na5E8KWHGk0lBsBGNRU5Mtp59F9hb
LsLp2gfJtbiCAjtQV7H94sC66I09X5Vq4XnhIsdDLG98Og7cSSnL+n83+/fYTNEQ
nAaYgalGQYdHhJPEtljwKvxcKHU0C4IF/qtFxKgXtNQ8IzBxWv7/JOqeYgVOMdUS
qWnwWaL4PLavXkdsc78Ngw5o6PG37i6d/w0ovl5SYAai2TnD/H9uYzCUwauCIscd
9c2SJCZG6VVYiKkVbWWdTec+th10a2+NVLT5xlYH7KvGdxwKH+bU//+iEh3XVIGW
J2jlP/mTyZl9cvwndP0YXQUgcW79ej/OkJtkNe4Yibtn19mI57kDm7QevDPub8f3
DvM7WHJhOMr1AG4XvBLhFLT0GYXHZ3jvn6c/BRp4OtMsCSFm0mdg5t/YVHzU16uF
p+2KeX2Mhu9mZ7Uy0LlsgoaN6BSsFchxmBr7YzmadMp6QryQwrWaDTO1BzY8MaBk
9qWNLttcT5gpFdaullPAb1GT4riZzFvrwcaZdGnITO6EKvH+czgaclI32NniOxW2
Ob+0ufRUD2xzc/s9HWEB8IxjPSHj06RCyXlP3XplAIggJPu0j+hiuIEDC5tDffiQ
pQB9Jmo4NXRQpVGW3e2A5PoKyWkqgzJMJ/Pbv1WJLn0ViXwnXvVQOY3QAYTpHuS5
mlc85MmODohO1PMwtRmk+00I7TbTCwSPCiZf9NoCtVbmnZ81IczrHbwZZBVPR2JF
Kib43jeuWgcy+Wakq6uvdSDrJG446vw0ruP7ZdvNuq6m075zmeI9kJdQU6M08a0M
mDewgTvsogXcdo0H898YMAV1wme8ojrD2gpi6MOMTeK1oavUHS4fZFjFBTY0TpEX
dBQdVJFEKkjnO+sSGk9KTm0m98G3teFK4fWZArlE6L9lIKvmdYDIKNyDuLUREaaA
fn0ZVIogqSSdKzcg72soX+v3rv+aLNdXr29uj44Pi83IHI944/HYK6wNIQpTRbvZ
64mf7UZ6eS6FbxK/JYVzhmkdC62d4WJBunb7URGaGe3rdKG+s4upUm8Vk9YCTroj
6psCTeMAUa0euT/vq17nCLFVzNegqxHNf2LY52A22a8Jt0IjvBpRWyw5QpY1LCcn
AVGoUFgyU2x9Ln/ezKt3+IVcXULjcyZS39AhEFFwEzbVaiDjnYhHuFzKWtFNx6wK
yGgliZ042CohmbF8/by856hEvg0fBLMoBdVvLjWEW6b95sy57p1YONIJmv0+Omak
umo0sVO7FVB2bZUD8GcneC/GFgwfpzovv0vqzuZxnte2HyLVAyhsvo9kY61MvdtM
R7spV+KL+3CldO2XMsv3HgTBeNBfQyhwe0iIma5XuPARUl8BPAfyCChi4NNHy/td
UgU5TcdX93ZjiIldGQzte+ZVBF28II4mkX3sVF5TxqqJDKBSCE0qYLgJate2z9Wr
N7DSZtOy1Uii1z/T7OwnF02La4vmHXzq+EbNk0I4UUGFOHK7uVIcRC7ZM/gwWxL+
IFXMTaT3jOsCc2PwoweYpqn+QuGEBHgAamhm3QSXkcVBmaxtcUZO/kjxHAvVrvGH
ISQXRcCHHl0PKTy2ZRh0A8rJlU6+50MwuJ2qrGaRN/PnT6SpBQmDwxnGND7EoTle
jczmeDgTQucntkgIHXUBIi97l1JAoY34spVdIHQj8/m7dvHZWuXB3sEWvcpbRL8L
ADPQ9LGoIBxBn//qD2ABFFIqle++EHzDVuS9yk6DZuqkewWgA+Jn8L9QxFwG3uht
2PAsqf6G0IVifx8vCJ5tcKLBeohICCZ9mVkvZvX89bt3/Ig+OyKgNnGKq3RCPhl2
oDZHKIMYW7fm5zn6cOqll3kAOgkKWhrBVjddTb92eYP8ylkSgmj7WqMTHxb0paNC
MzWgb3C1Q649iv/e1esEn0D+OcjFNXasoKMi3RlrhwKXxgCV0Vh20IzQTWEcUySf
aou2i8+fsE2jRCfMYSQRU+PtXmGC2M0jk54T4UstN1W+5uEOyYVRfvuWRCZI8kZd
4GwlzDfEnYFOM3NO2x6XZXcAUZDxfhgg1Jju/l34kqYP3M/Nr/jb1iqmhYtnE7xT
ZtsvjVfgN/LYFvooUufreFGhF1+69qdKzz3sk0/Ld5GJbsQ/Cq4qPPYHYCmhJeVg
2wnM47nzFS8UfFZZZ+nnOmFuxq9MNSP0p6uQmoHlgWI2nVszER6ugE0tHzHL7LM8
WXR3rgj67zG00OflWGA8Xp5jnLkKW/z8lxoZfbuHn1jd5raJLaGB7tMgodklT/US
lXq4i5mH0zJSCsQVpKspozw6ngsNhkVLVT7TV9GghchIfbHsCmryV2UvqWWU+nlj
ND0X+cTe+kMnEZufBxr7Eh5uYrYeCIOfNaKkHsuWT0PtLxQoqqsnoLayggRdDFeJ
tk2/JHq0gZB3dfkLMy7mAQKmeueqGuYdPJmdBdldh2BMEy4iMGX1I5glSOJOXNCx
reTl4DEo7AKZK4ASQZTl3YXgyw5aLbTu4LBTWJTdehi+XNIRYzlJ58L2QIbj6EKR
AuLqiE6vRNScanEPB3DAdluMRVvow5gq+ppoe+nf5Lcq4iYCBcdlKpvJucacRY3y
uN6h8TnBURUWvnFVWeapF0aMhkQf80nSm8hw3PWbOwwCOXyFe9ufX3kBlPhkeMRy
YKJ93UsngMPvtPk4HZcx6cmoqUBtb+iG06yw08D11s270mviAVI8bMMTp9MLmhgO
AiwMZt50UvxTAODfRzCjpEdAa+OOHo5+7TcTTJLvHTjRwfO6q3xhxq2tG+xIa0uE
UKjtgFWCvH6nKS50z8eCVlpXSyQLYviAavqbjE74x4b2W4xRI//itTuukY2SH6T6
UR8r6u5hZRPV0PwQftG/lJfa70zO6bbM+9xpKCA3nahbid19Pq27KkclLBpstJlH
jIo4MgPuTpb22/ugq2rkMcN9vgIcEUqpl9WsflR3xzjpO3gfNLAYquTmBusC2NoY
okxr/F/bZkhtVDXtUlr8YTvE5cYCY0yTasUvfBLecp9NMVzPqFjWnzRAD7BtS9kh
eWlMWLi8OgE0vN30U7Hje1VJRJBl7Q/5JennPWlRUyN3Cr5iC17eICi4FVuYdoXy
QFU7ZHHHQHED+kMjNpx7aoAwvz3U0PLVdA3PEExpnb6ixdUXuLA5567x2FvOE7MP
aR3SiTwjPkri1h8L0S8Zx+dqmVCP4FA62864a896dDPxq5VCnzTvQe1tXAUTlhOH
kJHZxpIFa6I09RzkE/JmdoI8xaKEUWlKK+3Dy3Av+QEso+QA2nQUBjXVMd4oasqF
d80bOQ6T+0ZXAchN3GMAEC03hN6UAG8j38YSVQzO4Lh0owEAb9lJYYY8B6FVcuvD
Mm/IrJO1SguJ4WNWinEJgEtXnoPVS4IYTOa3HLj56xp+89VBv+TIi3t+UFILlUe0
SVclM30YJYG636ibqbKcDyrsHEukp0OrDe2Bxx7+fM7FmacILz2p/7GjLCouoIXr
66j6/+gmY1uAKFyzLNJQaA7Sc7ubTteAdueSfqzbgJpMwJSd1HsquHo7AryM2+5n
sEbb58Tcud+ETC7PuojQYOA3HVv0iUe4RPdS7WS6Khk3+0NWlIkgKULoX+BKWXS0
wAtNk/jpJziv+hT4mLp0316ZwTEdHDOITzTai41h7E0ZOzsLATGRq+xY+SFUITqE
GyCWTSmszpuNPir8db86RaDIm+FvRTKWCNQMPQ0qwMz8vgf4mNH8KMXLUvRDI+58
`pragma protect end_protected
