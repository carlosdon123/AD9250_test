// phyrst_controller.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module phyrst_controller (
		input  wire       clock,              //              clock.clk
		input  wire       reset,              //              reset.reset
		output wire [1:0] rx_analogreset,     //     rx_analogreset.rx_analogreset
		input  wire [1:0] rx_cal_busy,        //        rx_cal_busy.rx_cal_busy
		output wire [1:0] rx_digitalreset,    //    rx_digitalreset.rx_digitalreset
		input  wire [1:0] rx_is_lockedtodata, // rx_is_lockedtodata.rx_is_lockedtodata
		output wire [1:0] rx_ready            //           rx_ready.rx_ready
	);

	altera_xcvr_reset_control #(
		.CHANNELS              (2),
		.PLLS                  (1),
		.SYS_CLK_IN_MHZ        (100),
		.SYNCHRONIZE_RESET     (1),
		.REDUCED_SIM_TIME      (1),
		.TX_PLL_ENABLE         (0),
		.T_PLL_POWERDOWN       (1000),
		.SYNCHRONIZE_PLL_RESET (0),
		.TX_ENABLE             (0),
		.TX_PER_CHANNEL        (0),
		.T_TX_ANALOGRESET      (70000),
		.T_TX_DIGITALRESET     (70000),
		.T_PLL_LOCK_HYST       (0),
		.EN_PLL_CAL_BUSY       (0),
		.RX_ENABLE             (1),
		.RX_PER_CHANNEL        (0),
		.T_RX_ANALOGRESET      (70000),
		.T_RX_DIGITALRESET     (4000)
	) xcvr_reset_control_0 (
		.clock              (clock),              //              clock.clk
		.reset              (reset),              //              reset.reset
		.rx_analogreset     (rx_analogreset),     //     rx_analogreset.rx_analogreset
		.rx_digitalreset    (rx_digitalreset),    //    rx_digitalreset.rx_digitalreset
		.rx_ready           (rx_ready),           //           rx_ready.rx_ready
		.rx_is_lockedtodata (rx_is_lockedtodata), // rx_is_lockedtodata.rx_is_lockedtodata
		.rx_cal_busy        (rx_cal_busy),        //        rx_cal_busy.rx_cal_busy
		.pll_powerdown      (),                   //        (terminated)
		.tx_analogreset     (),                   //        (terminated)
		.tx_digitalreset    (),                   //        (terminated)
		.tx_ready           (),                   //        (terminated)
		.pll_locked         (1'b0),               //        (terminated)
		.pll_select         (1'b0),               //        (terminated)
		.tx_cal_busy        (2'b00),              //        (terminated)
		.pll_cal_busy       (1'b0),               //        (terminated)
		.tx_manual          (2'b00),              //        (terminated)
		.rx_manual          (2'b00),              //        (terminated)
		.tx_digitalreset_or (2'b00),              //        (terminated)
		.rx_digitalreset_or (2'b00)               //        (terminated)
	);

endmodule
