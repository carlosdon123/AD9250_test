// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:22 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fEy0M8Z/gufr/tN1UHcr9ywsS5jRbLBSe198RQaq5FM2KfCYzKo2KGRbFKrx9Kb7
Vbt3Tpytkh5KSy+XVHvfcdwUWISGC71wJFmwzfYOmOlubCCDeycaGAQc+x93UvJ5
tyJsuTvHVBMAn84WLcLROOpyQjYLLPoYPWS+RscGWBA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32160)
U2A1ZUJxNtr4PGDZ1OZiCA1xnSvtwvzHvbfXUpboCIy6WPBIGHnVQa6vKTa9fo84
Wokqr1iX8bHETthjXt9W8Lu/wmrOuKJokCTnGs7Y+fCr/LeEcZ2TIW3uhJk1HQKc
Hs2lDulkX0NKBJz8rENXeu/Vjj5UCarcKKQyO1IUlaestvfhNLu8d7vFtas3XUB+
rhxQA7iKUP2lYPU5kg9jtaPWfVJ1a7wLZw7cMAzrSDaHj+q3DjxdNlOATYc6EcK8
lvhIzwPl/OfJmPAPHW3nosTpRkp+Su01qtm583cTS19oXNMegtDy0zKxqfo+aPH1
DL5ANCjze3YZsQ5QSirJPFQDER2vPgqzAY4jd8hTXPHb+SYy8BZdJhbPEHP/K7L5
ELrjY7Z1YkDmi0N/QzBaO5UQjab30/5RMSBPBoVPCXIEOWonqUzAEmEtQnCasrzp
qr9t5bfbt37GAVi0AF5ZYG7lYIe8FzncazO8D5jMFZZTNB25PTgXAFxYMEgHQRCj
0pI5CZms3IMZI1dgpsCdxH5GsveeRIebVmA0IMuQehE5yhEnjShRl0Z9aX3T3D57
/xhyLizm8tjq5hfi7qQoF+pWCHxADuR+rAfq0WtSqjaQOS9YAhD0MjxiRMHtMJyU
Rvyb28Bt3ZQMmXShUCj3E6TMZteLvx3eYAkr/8mRi6cwNTFQdfoK5YPGRK+y4KIi
CR90uHtMbED/tV8Vs3mpuESIjDRsVfaYEcn2pUe6jEUgFlYcMyHSMwCjH1YwVDwV
V2FPdvNklvw4s1PckQvF2BdmTw641Lqf6R0//sBVAvbOXxGoUacsnsBFKYCWkr4x
imDkapJbyVuD0gOk8vpKBxth+Lrp8QnfKJC7obkmBMbLKwJckrmpX4sz7smQvnRf
5GaDNwmvlYrXzuUcBA0OJG2SfATEazvjL1Q3yGKkuuQ9ZaVjA5vLMphCL6kKkj2y
D+WakSFIv1DZZTxLHW3LgkG764HnzMBlPUKdeaEwI4WTROIwcsbBxbcgsKN7xGZ0
QPNVAlx3+KyYzwMnnu1S5aGClK5ZQ8N92xge0XHp+iYxz0hSNAE2tuS2iN+yYOtL
puDc8tyVOGZj5fxjXaaEUeH3DOKGir/W0vLvNetP5TTY6FYH+bTCXXmZ5lz9FvsK
qzZCF9w00OJ4dl4wcTODNBrEOnaexJaGtGDyphp47KHVwNnHZfq7QtN5VCVgaatv
xmRYF0H+Lqbolx/2KJ4X3Zevt+ct1YcJciW0R6ZPzSuazpf+EnlAhTKhcfhqgUtw
MVtCOFYUFi5L2sigH8amxBk1+hk6dzH5FYp14Bwq4rt77lSmKLdZjV/mBnTs87o8
WA0mbMqyeOcw6OMLbJU7555s2Y349TTPcm6yDER8eco8v4YfMLhSY4m1I14Z6AXO
cILKRM9F41v+kwprIvu1AVmChBApzhbCL+GITO9kqyJNb9chBYHSgzrX/VubfktB
JXEl+wHN4hYOud80wICwJjRlhBqN09g5lXKeyTwVmqFZ5xmey9I4dpXwMPQIAI0z
BlYiC8G+inanMNxvMDe1Lj1ls9xwdPWk3llCaDpv2ppvFPtK1tLVRMfIl664SFoZ
g9HDiLz9jLI4NzARxck+3ge1qI6lSTeO8+7CzeRZYZlLIm2ueCclgMVlXppcbrqo
BfrgcdAN82u7rZ4gvj7DTZdm2GPtaORkRMvQnXFlvdF9/CXQr8PIEScJjVz7QBFV
Y8VNAXV1ESaUYqu3AlAwRkQNfxQhPWFiiCFjcIDOTc5x4DzO3qvUlvIDxKpObvhz
i02PzqLR5QkRhn4i+0HnMydNmRMTnFnhEjSt8ciE2Q9OABSltHpgkFzKV5Vb6L/a
L7mGfYXSG0Gsz+ZzMlixbtbi80JyP+Kl552Gtv6kevvN7H1TEq9OpC4HQkIjNNIV
HqFoVTJOnpckBWOsHbmBIE5ePxlKh2Ll2Spl8W4EZhz2sTcaHgc/hEyRDMheehX1
AI1y+STfraVl8Iwo1xMwNUAnGPVOp63o0lm2yfcYPVMX50rtfdckOnsAb6bE54qF
/s7MUosKs1NAk7a4mVqIUPufycYEm6I/HEfuZjIxILI3Aw0aUWT1jGNOeWyMLte3
3kw8OOFoT4Jcl+rnGUIGd2H8LMwRUwybf5AgB43bktI9EKo3nW3OpSWDFPEf1p3r
E9ZNOV1AoNPloYjGpZE/jNK67usjRs9HgMtgyasLXxItNC9zdfRshNBReXQjr6kF
BFUQcn+eKfWzOMc4VPuVCds2ao+5m2EhSY12gqbPu/+ZrY7nWNFmHl/NHzBHRG7L
6hh+hRE7Bc90WOnbIJWXUq0/W5cNmysBuz3g99zQJ0kFik+76j568zlzBQ81mlob
vnq2rjww+RYkpnmvppIzjpHAml8DkJRaL2a9gX47JOMABCzuHiFWbCCJi7FursBd
rW0lKpECQugK8NUzmnFEDYBBTFvS9xynqkYXLCoWAD4B6XYZwdSCtC+hVgJwYYAV
4gztxW43SF/VE4sNzJmK8wgK56C9droX6F9T+2UC3KvA3F9XsN8QC+qrjEmi2UeX
PHFztli/UhdyKsUZhN7wBUVoIKX2ZP1f+0slDA2bOh+Ad/WzDdrmxijDBv7cDah3
l9W5L+acPjbOahaYMIf8wxzmeO4LjTKPQtUoKRnK3y5T73oyqqsomYur7rmcszyu
mvyfW7Ulml47k5GDWm7G+v9vX8G/l/7fefsk2iCBja9FAkScPwCYmFxj7UzOFUqy
r6sFMnRvKz1wDhapTxP22Rkdnd58urxVRFqQKD8s6kVKUXrinzf43YX31QP0GNy0
uhv72izsI9Jl/3e3qnd0oUwL2xH1GGVp5VKRMLg1mSKv0BYgjmzJmsOWk3ultA1n
0MZCHOh8E/ch0VI7E9P9geqxSmdOY1W24x6gW74NJ0MUeC9ctGaM7Dc0qpFEkEjL
Meltvfocp4M3uNyd2dlooqO/2MiXtop33KoHlJNEoGIoWE534vlSAAc45zNJYknm
NfUJPByL/uFF2BZFc+m+RowhAzEw18D4c9mCKAXJU6m+svVovqWyu99SIeqxhN2h
hAPHsaBy/nJ/mYF6mXnpiD5NDeMZofqhBRr2z1wEG4uNOLSqqjXlpxZ1dOAE8g9F
rWRNau2kpGOB3C5mlJ6lLP4kbacxKsek8UlyjNEZbFztxBko+a7MLerBbROrBkkp
x9keMNEl4VlZM5inrCx2YLQddfxzTtL5LEv4OlAEN5UY2eri/2KEAzRUWikbmRIv
mVesg5XRK0PFNMnNvDbhzgaAZTHHjcBK517TOWHfKz+XZQIGeJOsQSBtntz/vHaR
vEPcUGZ/Luf2A5B5kqU8qxVwMXhym/r0yX8acw+HFXQkeIrbitCA2DKK1Cq5tEBG
O84loMPBsG7KAmAZ7hJCGiD0c5vvEGrb2BxdNouwrlx7C4LXAuqcXbkajTqv7SE1
KZPaRKrLQ9H63l02NE7mnTSAl4Qg5svoxq4Iteg0u2Pf8DJCjjjYfGEb54efHDbl
0YaccMW2OxO2iWkTTzzNlApXMTh2V+Ltt+FN0lNrfv9OlR16BmYt1sdkFEKIkSVb
XWICwHqm5+D/jEyfkFKw4Ze427qwUQc+EmP7NSp1fThtJ4O+rZKj0g/kfmg0TDb9
2Yzf55sCa44TBdRV/MfvY+Rt9ugU+2C+dAQo+4VsIQOlSx6jotkk1J3HSs8e/Hwd
p+cRSbixK8BOWSjYvPKgcZ70A+cuwWKQwhiEHb2sm1uoxnTZae8K96nK0aZewuNq
KIewPTQ8BgiIWO5A9EU1qqU8M4FQrsOaZwDUS4PvLp7VGKQ9Acv9ZmKRaKN9Slxf
6XY7dJueNL4zC+6GD8bQhH0szId1povWnNlNFr08760XvlKx0OSh4gRZFr+UX1rb
7eq1sZphVbYQBClX7LYEDwEV0atBVuFap5Hc6C3RieKN17GBEFfLQv/mw3n5AzXQ
ceQOBkf5ynforjVQ1OOwI5qO6wcX17piUqamOuDcN8OUWeS9cZl+Vtm3dEOmijMn
FIzs8J//DXu/OKVD96OGGAjNht7WnfqmtcLLc4/jhXwADnRuCtzDcWibORDSsJFq
mx8WjybOuUZCen6LGFjZX+kvAg1avW0SiSPY9QinnzrOGhnspEhnmmoh3rRAb8OV
0hEaRYCCPPnAsVtNY8SBsDtzh2kWM1gHDDsbozC6ZzvX06IrpFYWvUV6LvTR81df
pjaOLBHC6hYbZkqskEo2gr3lisVW8Zhb61QXprymnlq8b0BQp7qcSbgcyov90VOu
g64oDqILC/CDbU+j6+2hKwKfv5h4HFKL2IyMpnjDcTNaZXxTt5yx8Rfe0sbaxX2l
kFbni/xNWhkOYL3jBwo19G2jWgSPprnBNC+QS1nJKy1+eVdK7YHLoP4oeckoGWBN
XkbQwPlKyI7AzGDx9UytsHU/UoU05RG07Zo0/SuM1coJ1AXd41ptLL0B2YepoPup
5f+wGLwURCJDVeiaHcHJ2Lt2OPlS08q8p3+M2nuGNitt6HELr8QC8AZqnbSxdiQX
KUBukjuKISLvhNJaUH7JgSx9GTsC5OceSYVrb5gXRv0HCmEWv2ezaKnxP+BlJn5U
CHMEanUST0vULhnMN2iqldxBgNY5mLifqbXF5PLgpFh0eGWWZUeNi2pvrDqgdwFC
x+Nxiqco5UAXpbne+SpPGFuftrCriA0rYN/ZGLXgbg083d8bzPv6CEED4dqb4DWJ
DUIKWsWuKIaTr0KYaBei9JIydtVBulM2lVJUEm5JWk+NHc7NNWCKb/N9v6183W6t
hNyareMhNFjaCCt3EDEFR3VkKKMwTZWMNwnWdAtOPQADLBM5wWh2fQgEagPqbbpv
f7VyHZt5houu1tHPKBgwOQaNlyflvDtF8lZwxQ/JKw1+U8AAfdQHxIwtdqT/pRxM
QHQW61FHLyq7MA7JyxDdWeGcOLmcFfV10SnmpCidseMqJDfBtidoNgbtHvJ4CCbM
PEe9GakFu/TTz3h9LJ7Dt8kgBMz7I3xODHHloFljawD4D4iIbyU5y+cPz/txTXjx
Xc7cZsyik8zXnU1SPrJWDTVI1UjRuAoBylHeVoCa9NHrdG1K07qZg5dqpwN61wC2
+YL4WIZ9haZkrspU/CKa3iWfbtNachcBaDoN7vc8pAVgiuUkpOSD/gkxyGYCfxhq
nCGXJEKWpkRTOKowS33ILbjrNe63Pw3D33SjKajgHrEpzcF+GAcLXXKM/Nq78MET
dnSkTIFmEbKiPGw+3CcRFcoV2a4k7XdMkl1AcxecIa05ZeQtHu3qhT1aEtQ8WeRl
JzgpPfHpTleSEAsIDroOFNi2r26N388OCzbKhX4uBDf9gx9YkTRnJmSKD5g7O5/h
qnRG0+v1WYhDrlrCYGV5jhKDSN9Hus+dOxsp/1hUfIF6hARl2I57XIJnQeIbHs3s
yrvGGmLi3XI+lLPhkc4Qpx5nbOiNUBdiR1X2Xy1KwG+fxgK/+aungQ7pt0TxKAbb
l9+68YlaAH75/7ryjgmRQpUzBYE/KZdqg//PgnVnPbp5shWX9K4yzqjn7jeSxfdl
JZJUSQYYWUv9D2aFYjI3qTQW5/NQUTS9nDxyObmT6qZjCZz3HKdxYOpgeCxhjrSm
Q6HwEGF5mLF8m+snxrE/dXWmy3Bml6vbWz3xjpGHV7K9XVkIT8Xbp4UcteS3JR5Q
68spfuiFJVtPUg4ZPuvLpYgGAolMPTedyINhJCSbH631t0KHZDQ70pYaWl/Sp0zc
MWda7BAtFnUSuy69KXJ+VIq+zxkeOzUSihK6oMa8q1io6uq1x0r9SP6zwbTsVQoi
5J8J8fahuGxfAm2USmf7UKMAl2rTH/gGWUgldmoL+vteOyWxeXQGM3/qUauKy3VN
uYM8cAjCdiaFEWZJ+C4LbxvZqs1wHkzoboG/FhQRak2cl5bhvQX6BnJ4eaasUhM8
Zh+fsGX6f1cQpeX/MlgI/N5FDyvGsleTF2LNph1SsUX4Y5aljCR7FHjoS4ukWirI
NttjciMCO92URnqzf6RJHxDdLjduufeZw5jjAQBVTPn9i8s8Pd3ZJn8Y5fnt/78E
w3lPs71KaDplZ1ttWEAqsAgFrvdoEvATsF5VbYMRQSPmCJUYLfRMI3nugQTplXkc
PLEN13ePNdGFymcernRuXRXj321ulz7qC09inwJXXvFp3c8hnt7hDTItq+WXvnOD
fWiaeN1KYC+lZ9zA7yXFF+o0yeU/G3tvKXuAxL1CJxh2JptA4v/gn/+YQJgUTrDV
gyudhujWX7CL9pt3Q+XyZ1LMlLsapd0DYEbbqdlBznfZHzMLmSjSV27eQSHTc8sC
X9VBF98Y+7Ilc3YBWkf9OGiIYJiY5+7E7DICSLqgCluItTZGtQoF+1NmxxmhhJa+
cbC/48YoNyxaMKcWwHB4Y6AQHXQ6hPxxM/yBGMxlFRQiGKRCijELSzf8XD8cWjfc
th+QUs3oMHcq7F0qMvlodpNhHbUIgLx63ZcaAmuWlk2zDxcTPM4atqSTkdPtFOmr
HE4Ixcsx0OyBRdZXAZ5QE6wnDTCBfzc4REVKlOvn0Kb//7gIQUV1Htu9HPqb3NRw
wIrez9vkfQFw3PirBnTw5/ZKToUAsFeCtC5pkya4gYsZ4wSET4f3PwrFffA67XAk
XUeqPFCrRqg/O7Ht7hHewH9o8rmEKa22A0HuU4aOWjjKlsVOc8LDILnAJaG3W5U9
CbQV6Qj8jinqFsozvWDQe0cMFgsYX9xARiUlUS52QW/e/37YFR314w5mU46U5h/q
nMafO8AV60tX4rdY+spTGgR3Ydh84wNoLXOrzAGNVLFDrJJFk37Ln3FDPOjCEeEA
pOH7IN/dTsgMJDVF4QNv6adgTPuqR7EhZ+GDULVIUHDLRMLKk59MqOrsSmOdFHlL
1arnrO6L4qSZ+J89r+MwKcbffP6osrWg2Zx218fWBgkW3Bfyfn38MSd2cObPuo8S
CBeLaNi62IxijXPXnaGSdk2cTrHl68HU9ge/mpUXlBrZScI0eizv2QAMOELb2G8f
S2j2rbXFsrxClntf8x1HbaLIbZ41zbtErsMBPEfk7P7tZjHs4cYErg9gwbJXA5fP
wWYYJRS1j9ppj8K+x3BNuUJqwcyvmfaeNcxAVHyTLkfGKqpsEav5nfdtSDMjTvaa
6x/KPQsSknCRpDwpQoDG98EiqQZpDZlEDJYeEdRj3BFx4A5IRhNye0J3WOeivjC3
1VJYRoYSP4kIqg1LZZT/G1HucQsIk5EY+dwdjIJqs8rPUyIqbcR1FCC9Ho4e7zNI
K2+o3vyMw5KaioyiVXHZqoIpwOafUMSB5I+53joxCdwwKaTB+awwwbEs/CaYNmMm
o2YQBxCSNwBu1pAfsGjtvGC8JFeUhXeTYDGEpN5wHIkNwi0kOT0/1OGuj0lhGRY2
SJby9EBOOETbnw2Xg4bcFCqIsBfIFcEp3pSItG7T2yFlcZpab3pBNnnRZUv3P4kL
a2nZ18VmjMSnzq/wLqIc36fhLsFlmxRfMUbiskivfYOGiY1vvsXlevY5uLNFO8nz
VYE07gf/I8r4kpHAeedRh9efqVmxuin9v4jtHlHKvGyjlIF2A4o8b8gS4Y6BG7OI
ZZnmmua+zvIA6FTUXFmInVmTEEgZSylGrCnZR0eixHsbngDb0fzDF1BTK64J41XP
WXeM0/f8qNzhhYPCdXmwSWTIfFpt6TPa0bGfcre7GGAxGTFBTt3hs/0RUxBQiDaj
bNhhpexc3WYZRAJLgjk+rud/rQEhbj+6OeWPWb5+j79FcXUv2OIpTvlJi9Pkx+rE
2zke6QWS3NM5ZN2VIriinLTPaCYi9V2mgocnIG/T9Sl9KChiVWLCDF019BZKGNDO
ChOVjrImGFEj+zcG4BHitYgByNOM0KL9pg4iebMNQkpu1bEw1f/nabEl1QlALRjd
3KZPrIjshgcP12vQWk3bGp6WY+khXmh4gvhnDT1KroJoCt1CAT6qaLy7a9MQjCbm
DNhL33/rhYbW/g6XK6FAytZN9Yl88XmLr50IHzm0iYChPuYF6ruHN2AwoNN+sj68
Z4jwOQzrgDOnD3Kb2KdzJ9L6vVViiIIwi7zI1ZrT9MvdB12k9XN+Ghmc9JDFUobA
ClhjSiyEp4qe/5k9P74lUPVrP4064gStfBkyMtDy+VAki0hnASrmecM6dtAe4xgg
x4wukFe1OO27RgWtft90CBvsl72OmJ56dtN5OQUznMpMzEdbdsnJ4gfgi/Idz6by
bhNIYItT955Z339Qsd9YQuYsXsjBYe4hzsnP47w2GloayHk7puEmzj653F8RoGx/
5ZEgBFkMz2+EgVz/nRdJjJnWqFKMURd9EXXE86M8rj5avx2uRAacIcLMs8KLzT77
53CPG0RAYefn5DSZlXs120E2l2Ohp/y2BBJkmMT/DIDe9jBxa6fzvVV+tCJ41idX
ZDa2GdxBHIfIM7BKJQR31jYuJtjraUc1kZKK6xeo3UjSMRWlOPSX+vZckR0Mm0WN
iQ8B/57VBxVf3AjNUR0P2BD+TL0xmbK8oMT4GyDukqNR+7AMrZcdb3HZJxXlkrac
qRhfo9ci2VuQbs9e8GR+/5QSRb1jRj4Ppq8AmZzZ+PagEGtpEHBUUjNlZZHdgEeV
ou+IjRImnevVsHCYhIr5UmQBmBDvHCT4CD1Ajz2nE5NSJo9KtV2CuYVZ/wc8qQJO
PhRVKzNFqSIfys12RlkVM8XutdiGmrK1h+3jEYexVgS3Bd9caLQnwhmF5VUZfnb/
S9wjObwn27pPYhc7MFyQp9Jax+hDVLJOBhbGQLXo3QV7ABYsFFGrThYAlBDvLxPo
AFKiJtegsX2ye3R92eQvtXs9WD6vH70J7/yFjJChfikvx1yLftUHcBqrIGVl7cGY
EjVDfss1jJGR7Wp4KtWjVq3hU24iGeNICKr6Ta5Wka+VXu9emFy0p8Gw3eaKs5HB
XxRauMU9By3pKx1KrVDybloVrgQM7fGBDzlhSVyNtsNDTnveHD8W8OnBLMccbbJD
E/02sjPo4hJ2vJqt2zzTaBBOhI70bip3F9tnY3I4XKydxnqt0T/P9NTv4dv3zSTx
5bNS3uiBWTw0tCoYju14d+F+Ym7d0DAWr5pJiWTDbZF7MucxHENgOimrLRtx89pW
d6meHof09kuQezZ3hKtj4YM5eizT+DbdvIo0K208bmstTRf0dSLWwWU1B7OWs58a
3wSkX3BJ3fKNNmZJamavz/sVNqrNo/5VPgwh+xk+Z+poRl4E1AqJHQZnQXkAEgRo
oi08Bcf5uejab4UbT6GNs5Dq9Njz2xM5yg+KLXLQJvumfZ1czkiMTKzghR82Y7Ky
h78Mne0HhoMH/WgGwpIhkCoaH67We01zyMcV9tUCD0/jt6GtVRMwzG7kcNDkeJSD
MasfUhWgY48majqdsOlljMCYF/hDaIW0HfuGDA261Si+8/qMWW548e4RftkI6sjn
OA3GRaO8UYifZC5SCDFYS+KQ2Uie4jOU5k23vWm3Ghz8vJ1T0mf4CcyIkkwL12Bx
/bcS1JFJQoXCyhi+MjcdHzAYQhHpzmbOHk9H0A5Ix2Rqenr94lWrFBlGALDQjp/n
ug7ze0cKtAbASgJfeWVOI/swku4RKKO6F98nPTeNSOUw48cG2hSpZqXEfliXxLnb
AomTCqWYySBjgYgrEoHbe78VD7palWZqZAnCe3BYQk1SFl2K8WUMGK3TNMl0hL+d
I3tGLj0pbBzIUAhRTORN7Yk8buD+/gMJEzuKorqgheWh0WU+IYreJHXZwHlGQ8RM
7t+2I/l4+VGDcwY/rrYLNASav0UE5MpKYC0pDoEoJnyTY9XqJhnA813R3CqXgwpi
uChvvMVo7A7ZJfVN7z0Q08aq3tws9iclROplw7u3gAUHVGxnjUv9cTvRSQoUHDNY
yYyui81Ky9Zf/J4epaJYaxZ1hG7cW732bw0pBifOREvzspxHlAOMAw5kIVbmSOB6
HP2Jm313C8RqMYZErnZ7vSjNiIV6/CFiQl4Dz2lvMNPkFPlwwiUjJbyas+wjE8rn
4xoZDVRA78YuBvJKyYfYfKHNMsLIOy/X+/hnzkAdKbGHZPyZD0bvBeJ73OGj/RRJ
DTW4PvLt12sY3u2LSDyevoSB6FvX6j+rO/cdX/ciUj74dowgJRNBgRIjfMuaIh1Y
mjs15PRtX0XiUz7TznQjM17rllv93bBrhOZrAcrsxL/OiJmKeh0hW3FkMpqn2DyF
SM65ZrpSSaichDWR66hBDSs0RP6Qr1n85E8c/2yH3iknIkKpQHIVmGll6ibLZIo2
57rWaKWy0ARhpKSpHRngBU6SEDrwYhPCW67Kvy41EPL1DfqBGXSkBLBm5lnHFgF+
OcTQWUp56d7sc5uAF8BY/2M84eMza/8Va5fJ6Bp5s3vcyopKZD2YIiId89jFzcfw
eLjT4H0+Iu+WWSaxInw9z7qr79QUzRISyRszRMGHOAplFAlwq2/4i+3qcIi41Np4
I+ZRO8L7pUxHL3t24P2I5Ui7/90uL3BjyhMtkjD0HgTZZ4pgIKVdAMhU/UEzmbP/
IqXBeAMjDOvbp1CtHOcLlvf0abAbRZ9vc4w75joWzXEh/l9+gu6SyuddXxFo5QHD
YZO3UcoArl9d7UuQD9hGB17yc3Ft/MpIrH7eAee4bDXhkknJUjLtvC65wgK7tFDi
YLbedaPnJMbNjjlB2bxXKrE5TdJ89tBNdI+IWC9C7U8/8OBbfyPV4PCUs5QiSRKu
1au7uWT3kbjmxrk0wNfRq9UBDl4eJzkbRzHI31k4N2FWZnTaGrZnt9vzUyPrEsW6
AVHGKu/Jz1vr0aTmWq2jdU4qgjiEzmH/F0Qpg/2ZdVZExSzdvRJ9PLZugiTXKOJD
1rptLNIvP/XeIX27S1373fsw3LEDbWuKU11B+LUNWI8YnpDkHpdRu3TzNP4Og/3R
DPpg02q9jXNDt99NiUXd05VhBH6D4TMHp4u/v4x9GJ2V804lb9ua/CNW9G728A5R
MmHiasnqwzzi8xZkMAIZhiz0caeChSl8r1KQdCYJhXwJVifrTO8gsasO07erDA7i
7HYZLK62EA/9nEx1V0hYIyKK4WNogS1/P3A2cl2Ke+MVdUazkY61D5p3ghsYVf7U
kbSPx2QRetXuMzsI/9CgvI9G9LjoyCSecaofOQvrYa3/8RR+NSH2Jc8pKVmEQON9
EybeRcbh8AkRtQ9btTPaCWz7CddVuycsde+gCOiwxjsRmR8uC+h+ciY3d/L7ZZYT
x8kbBpuAi98jn/BJb87dryVFfhlaHNxHO1z5b+yDWdhF7dB1QQRJeNrH+ESVIhHC
WtlxBqbVInsRG2OSGuOlWykYWPQ78t0xP/lqNyJPKswDDF/KPJWMO7R0Bl6c943I
B2Hs521xIOx6dK9WQiGsgPUD3dPJ8wB5D+mivnWM/H0Pm7XKZMyLIPO2SVijZ3hQ
rZ4yq5pPQmyWLsvZQFCSkO2f/Ank2g23X+i+CcLv+ebGJkIbdieJLwaAsZuBBTVj
8e5BWhUOCKhYuK4WkRfEQH7S9pnNJR3E4pSGGfOUzIVx49b8Ma94dE9sS+79UfT2
F0y72zVNCzofNgGDbYxW5U7VeBL4TKmhtZlmr3d0zxSstPSBEZwGeUvkl5/iroVV
+HXssMOATykF5NXZd+ZSV9+bKBT4uVKE/0eciT9p8XCxJD76GPjghg5VuPZTW4Qu
evF8ZxOgvDOA75do7CvqUPaW85JyNLouUGmDfKEN8w+mJHkWBNLLhptFT+3Y40rU
OzMOuRtpkZ/8OURDnIAdy2j1PDMGuChGVM6tFJQNdOCF2WOO6PDaVEV2KRX4RbQR
lh6Gmlun37u2dI0k49MlpqTtCsCjOHFW5Yjh9kFnwGDKHkKAfPSLqE1FrmgX1rQC
6g6dMDdNdKvmojkZ6BgypZZZ0Ni31Gqq/OMQqPf3lzBnpUitShE0pqZ1K6j7l35e
6+0xsq3FJZc3TOxrF4z3Rn3RPQ9kMcHyPcynW6+fnSojVk46hKkx9rktbr6JrQFX
YVEyNYiWKveyq5ue1wspizrexFtFyPq/PjRGU1KJT+IvA6GVTNtPFxfco/3Z7FXR
qSyDPbJnaBYT4rstQR+zWhW73tGJkXFW3gN7+Ob0SDpcKe61XEDGxz8OdrqLACqg
niar8YoUhAJTmmgRsWBlDIDzGLsMIGYIUOfPXsJT1Y4PlnJHO2+kmnX/PoUc/o2V
7E5q81iKIKw+lPThS1L7GBeSznnc8tXF0ipecJIs9N/ORu1mH2qnGldFm2F5Cyxc
9p3WkY4UOchEJn1Naom4urZGthHTcXj8uFvEhQwbVlxRmGBWzxDxaxgTLjbfRqtV
icdVckP/csJOthsDBt7Gv5lOwKmAt1ECSXqcD4K7b7o6d8ERLynxsW5LVWVhMjL+
xcGLXz1O9yyYbGM1RD7CTreRPSCYxWxQEqDYTRwf/65UNCs4S7gKnjp7wUDuDyII
UCufyzLuV15dQpj8JoK7YxHSLACTlVnnoNdYX7ccnk554abwFM1fxJzXyKYcis1i
AbPQxG2KDKaoricjzaa45BhEZ+snStImm+fyVJ8AXGdSJlNcVHH9iRMGN1b64+eo
NoUFLBDomq1+XoAOrPF9IEkIOUmgzo7Pt07o/iipymDoXnPl5JS99iTi9snoriMt
64GRCdsjm4h9zGbakzwdLXPzm7WOiN86QDSOActyjJEUgaGjIrsLZ0mdbX0sSgYP
D1ZvXxXhFXHbYeTS8qdYqcxd4V1Onxu2ST2BG0Qps5rK0ibhaCde7PWK0v47802m
IHzH4ABDo8lT/Zjk6UKVraEQG6qBMjnNBh3XfzusKy/qZ+zZ+kzwcXr8X/N6ep18
jY7Nx8zKII1JkMiKbCqOvy52OgK90UwHqSYe69sm0pQWSauRBVF7O3roPGP0JUSw
vamZuXYb5lfazKjqSiJw7NYdA+x90ju4A2z9h3uQCnGEOl2/2Cs3SoGOSqB1VkuY
dUpCuD/PJFhGEWU+vnM9TVa1Lrmphm5vmmqI9y+vJkibsh2tHf0DAqlGfRMHV19J
sgXtQt6jcMoNIsS7KvSyptFhtkFZjQcwUxK0ufPtxSxuvvbw4UVR6GmC/bP8RTPn
LViFMDDnabeBvnvnClJf29oMQ991BdL7e80gY8xgmoGlxALTZL/newj8QEd3SnSc
cohiTSCZjccU3YxPnpoGgVZn1GQG/FkK6hodnai4xgi51oCpHs27memc0In1mXc7
j3+hjmVli4FMg9+TaSHE055C9VpWTWMSHLxf+EjItpSB5Pg7ATfZRZ8CxWLPIiHT
WauUZur+SaQLKYPtHsdRyT1QhOTcPt7LRvL7EesiDIzVJVf3nzcv5xbjTwng5LR6
Noyr0nwQzGr9vMmAE1Y4qmEXNwO+QD/1iqXfpXzW5f3CDNYBVzsGnY3Bj57ItHjW
gk7G6UUgC8o1yVPiQmMSf3Vcx5C5rs6R9DmzheDayKC/5rb3jqNn0KrJoUwCQ+vk
TSWYwF3C0gNN9qy3h94Xp/m48NgNhnO931y8AB0Ak1BzBCFYOj50dF9pnq+8DrNd
Q1Zq/sb0WfsLyHhq4aPE/0kUjXZ1adosu01rRnV3Rm2iPr4R3hmQ4acG1OFx1eid
VNF3TtNmcrRYzQPhAKxl9/SnkBPIHIAJWvkFujWBp4SdDkZyRYTjWMPSxjCBl8Mz
v6n0KOTH5MfH10Ut4Bp2HJSrKGPdqBQTJ3IW1EdfU2vN5LQvLo74Lvhi+EFfboeL
HmDTlZpNMRA23A52MXMxzpnGq0KeRSYIGcYg8EbsOxQoZS0sdLJkqf5v1FwC9YoR
KQaFXiWV/RydLwPJLaSP1V2f6MZmhzFRwXTrz9oEVrVBL2y7g+BhczG3K2NKxVaw
1qe0IEighwn2ouM8EqnGnGCEbsnIBvdE0dOCSgfsimwsNi9iAExnd/wjvJusGUQg
0+7Bvwa5Q6h1twY9m5HyKVbkCkDdmcdRDyY5LlSYiA0Tg46GXya30YtrZpbgEfPz
YPOondO2zuy9nZJdfMg3JIBt/Rds9I4MK2USb0Z3yKaXUDH/j6M0QrAWMsTw27Nh
gXbGM38tYO9xoVaUIYDzsE77E0sJk0x7r8rAicVV33kkEvTR+/rABl2s9XcxgKXk
teg9BpFcUFJJxzXkx/sYRI1rDEm/6Cy0aOZJS06lvn0mmZIqJCmYx31ZZdewQh3z
hqcgTttRypMWqWSstGErQsk+JfSU5A3tQFwFzpTNLYqEuMKZuWBpYqxr55GjFtLp
79vnEJ4ye63wMg7eBxL+QTO6Mxc6hd1NwTh/VcC66KQGsklSi1xXQj3TKJz3+AQX
6V8+U8+QUMvU7yH83oDLer46V1Eg0HsRL1RfuD4WEsKHN4wIaAfJ1m5VmgWX8DPh
aBvIPZY5LKNEMUmbE9Xe3mxYv09WObrC6f2AAzb5h0l9N16cgh+0TeJlyObo6XAQ
UBZwP0VW25ojGb10yusiWOsaUG6n1tlDzErdXkGOdOg0cv2mitkLtMEpMPnHexgZ
T/vqwPi9mXOxB87zLShTBEORDF0+5rC91i5ARDBDSb0KRbBJnKFaQLFRIW6E27ph
B4FG/gTnD8b1jXBV8s1QbpW9ASCHM26JnjmjMsK+yBdEzWlyYC6yY0YN8/QX6SH/
CeDXxotndU40gro7Waky2lihGYn9bB8MSi391CglLBuIz9Grdqk4aEnHo8QCrzju
DqJ/sDnttEO502li7KkzNZ2NlkoE5tp4CYAq2FRp3ZjYW0Ak/VGA9XWNZkxWBXYi
hX2rBSGmnd46C3OdfY/Fab8pdqVa0s1jdncPplsCfXGAVHn7F0DR7vbgh9L+wOdn
lR85qoUtuxqoXvGUroui9LGc2NreLxEUtyHVY/XIdhdofCXU7ISLyqMvslcSsnBk
IpRTP1fW0CLEhqfuWUGfkZORus3EpoUr9BD/XID9t+FZFGpXY11xkbI/rm6TVOGm
huKjlZ0r0ssQ7B/tTDbKnCbskDy3Zkn38WZ35gblWjAacsjkf1Qt8Pa5BItOaVm0
sGb9bU3dhyLdsa81mgPmeavT8MiUh7sfWpdPGHud28VIOjCSuSJrvA4mZ6XIGgz9
hdAcXFTgYOydwaQ7yV79BV7AtOYQ5Z5zGj6GMQUop58X0ycjiZvWC5cDRQU2ZRPy
Sj40gQ6oLF3vAKvb8r6C/e0b6o4cjVtPpynJoWeocWB+Aj4P5crC3RyXi55W9TJR
V5YeC4p1nNmJ3+u9dYAySBbFXIxQsp6NLQVVSUbGewjAOGEKjT4BPKuo1xm/eB2U
Y2ib/K9j6CHaSNBYUgTiaJbnjlSc/xOc9+XyQ81FqIevEFzzyVjrugf6KPDcPHQh
LD/JRFgDlDlNABggEGpwW03dUjGXrx+xjH6LdOAkZfjC1m3WK7Zig/GHfj7zcPMT
Z1PfajnTokC62NlRwI8CVal5EApxUQ63+9JTXOS4rRzWmJNh2lw1bCGhFPxW/phh
ps4AnHXng+4kiYGJMq3y8nUHlaNYwgd0ydppDTS4IRjfGZZztqXYRIcpKQFO0MSS
sD0McHpJZr3zDC3nqlrZAHs93JeiHpHXZrgs8NIJttGUdYKBKys7O5O2SiJbxuWl
9+/xaeEWllR+bBycBpHXPc0NBqwbQiG2hYxJzR3QxmdyXSBUv5rLz5M3JVdxsc92
YXiECEoulTqmlRO0az8i6AzSiP69Hu47chz0qKZFgndx+98ejSWNxylJki99Uwuy
NDdYwZAzzL1xU6ttZOQ/SImw7eVeAMH8DoGU6qAAEfBK+VBH6zCy6No4iU7VrW0i
dB/rsZz3H53R5BULtdwOLs/dmV94ALHbI24zoJaQSuizPJs8XytMInPcH+146Xgd
wPgXZt3Kg5/hd2C5evacVSMhpCFH23PKlLwX8OXOQ9XTW6vxmw/+WMh0lzvpovb2
3k52xaUN+trxH2kh6vu96FEokyycM7J9/VJyPm9GATO/iWad6Afkz47LvOgxcSvc
P2WnFUXlwkV2OPF1tZ/+N3ciVl8Lt8PGzcPGRslU6KF9Hpt2MXJXtAfshEkL3RoR
8RjPm0DjQKM72GLeRTV9OGqkE66L35+qZ9ZuDUXs8FvH1VJRF76kZTbaQF3KUl9o
rb3LR9BKf49xGJJnbOqD4Dll/0rADog3CqOmAGqI1aMv9aAmhyv7rQSx9uNndH62
r2ZVbpHD0tok1vTkx1s5uQ3sx9AkdLN7ObS+JdOxWZmj1Pwe5+10nKwYIgf6Y9ib
QR7kBhmCYmsHUUGTM/srC6gHCccQlVJf/djBLTz2zYdGbw5ly56ZZIrz+9ez7PdE
U0LfeX49ZlnjshUvRRXZq+jWXOPw9KD3Tr1nN2ysXmPQX5nmI1NLKJQgSsJkfnNQ
ZdO8lAfthfOUUdy/gHWNHaRxk+xOmydobOpGoDhMQubSRB5HKq8+aKBEnxLtT6OK
LzaW/bTcFWNkBQiaJ4ygglw0hdfKPoe4xlm9RrhcBKkoGU43O5m4/wPSR39Jb7wS
KOPKhQEABsUPVV+lyw/+IvvPzdnAyWTUC6hLb1CKK34kuIKF0+f9PbE/Kt+n3l6a
sGKdufpz/lbXkIySBPuDjnNCIe6sITp8FwTtOUHA+IpHe4qWhZBoeF2Mfy/EfoNO
bhZNLNCh+QSlDZDanmeO8DwSFqkEkxTEi23wQCY03R1GW8ZZbS3JjYptbHjnMlM1
Nyo3VxSCsdMmOypDb3/QtOy9C8TxG9VXHinNOsmnrtR8+0FoO4eAJa6/2a9RBA2z
5OlzyoFAXjc/qHVfnRSs5nk6iVpBj4sR+J7GVIeVdF9eJN9H2FrQhph5a/f/GsYu
GcR/f08laWt52Vmm9S0NedchA69+FFelqE/7RqSJvkf5GUUdVR16Jst81/qTtG4r
f0enhHPrYCxm3Pmy9/iPAiweU9P8/yev8bXPyG3tY3LQPrdE8qEMmlTcy981ZxEw
j4QXNELJiI5NYfLOa2wSICWGc8+Uvzxvrh1CsEVuJzMGCwIvkbaifHpF/g3BGpnr
aws2GIGwJwxNdpL+gLotXbQqqrQB5yeuz0ivAk2yVhYQRUQh1mDObt07dmh0OL0X
/pN5FgVY3qabt5OB9LBgjFKRDh1VHmC9myudQEcWBupvvRk2VtK8FeIDLCz+PyrQ
l6lLrWD5UsDDMP2aI2CJv8SZ1FtSMazVcVlNTznSv16bZDO7ZTX99y32uF+wt83U
OOviXYpNj9sQYaewyYssf2IA9iuG7wZiTCj5Q4DB3iyWtWmBOy5dJLidmETji/ak
StWXjvdAQ0SajUBYLZgFu0hM04UHsUCgj+XC5RdRPqn9xBSI0ZzCWLsT4fFXrzbo
NC0fvKexKX4aLiHT1e2HbmhzUqmx5jhKxekQyf5ZihnlvLZaIeoiPx+9ENsQx7ko
Ky29DV79Ohw/y2VRT2UUNj6ufjGNl8oBB0Cbqv8d1/hBvH7Ewj14BLzy5Ut+2DZl
HB+TxzGZn2TRm2n+Sleq4jvUmD2CfkA8UR4Qo8sp1R1Sn29Wq1RsAIiYL9y7o4dS
mMFJ1ZmDieJ4mRSeAl338XKfyv0WMRNPk1gwn5OcOWhVPQfEpNO52s1liO/YJkGN
VAj/UuNch3xvUIbuy/PMLk3tfPb0ZhTGvrU2EInAuY2seDvtTxY5TZn/jBgHUmFl
Hit6HyHlNUd1qNtldloRNL8gJFe9yOju0K4fA0KmG7fSzMogYT8R/jZLBTQKRN6b
n5Di8V62FWk7UYIwZ3Z4keuO7wJN9sPmBQP1YUDWy8q6eqiqapDiO1lDNkM4rfX5
sw4Zf1sfO7RJr5SLeRCxHFAbRQ2/rbeQ32Q3FsqoHLyeT6+6cyVxCdSb2u6eC6iI
3H4Bw8B1O4E6vTcnRcah3goxg3/kWZr7AgGVCjNWDDdXxT+CaE828ZWQAlTEJHPW
caQtPIvUxCMl/Qg/rvfhmhyUeOnOaCV8w3GArwmMkf5gVQ/RT2P2jZfyz9M04GNp
bpMfL484IUOAQ6GnQFh24MW9qwf/mdq5iGkUtv/CAo1Dv6zgsiwZXvA7GUJlhLmF
waZatsT4+PKIIRjsYTWniVK70+wTzf5cAAktQYsbXSlI8GkMbxWQDZ0mt7Cqz4yN
aXn+kKSukSBTSwnj+V7bL4gJb4fLhnCExO+vaoiYSWEEiCid02XACvQRxL5bJnXi
lP4sn5gtaQYU65bQL1c7wqQHUPgPUoBItRUryw6qtx8RlgFy+T84VSzusv/traLd
PIQ4UiRlyz10E39ApntV4g6OLJVnnvhfig7ozYScNEaQAxT+JcNndSTqbIr60P9B
Gu0Rre4D1ob34aQ6bFeqC2rzWc83LphSNughLbNPV/YDyF2i4fEtdAVW9yXwNmH8
4lsD0I4EVPAsh7sHYntqjsE0QH6i4dZqIe9OEEDE0jMYS1PBoVVh5ywXhOQCSh7E
qTKqQtoK5lob2GtQoPaPtq1sgSfNidPErArCgxbV3ICmYjRhDkxVI3ZVzwIpNg0Y
o1nJ2JuJridkeUuUNV8pv2CRYiNkGZ/JbVGfyT45pxMXh5OiAV++mLJC121iiRLb
zWkdwF/0KWjPkshQbHvYrJRMPy7qtzhg8CWNwMUFmCsBvVZbYCPf4GBhnv7LEcsn
DD9MHUkM1IWgQEtJ11bLa2wllP+QjMB7F6ZIHnKwFP4P9xLHdXEzJodIihbdgqXH
RsC4sqxsv/V6wAWUgQk8XuznqdqtTxm1s1kSwROhCWFFUIeVEujyuhKRJT7CjtXI
XQd0VHnpBXJ9DwzKazLmUA5mkhOUKiq099EyHPh229oMcyZlc/h0bbnEsMv1F6do
F9E5X5YSq5ESMS5FAa+Rit+AjqHO3FlE5lw4Exk7vFANbty7EenajzljgEOcc6W+
kwhjZ0Pl+RDaoippRhPEJlEguo6xmGf6RbsT6AtQlcDWCOUXV4u1NBHQzJNd6iuW
smFw/eypfvRR48rkQFnNgk03myVQxB7svCKmUPkgSEWb/HuVC+gudj9HN+A8Hd4w
omlDOPV5K3O9HpbqXgIpgQdVJ+YOK+J4rKPzwMCtzpoUFAvCvoIesXDfX80Sa5sa
1MyK4BuSyO+nwpq/JkBX6zbrci3YLc7f8Awq/TQi/r+50SE8NWqRfYf7CEeMvNsJ
gpXgGhs9GfWOrorSBmrNz/Mj3uLdDp4ohajva4PKivYk4MkrDLJtBqADPhTQKfr8
6AT3Q6yHpiCAYKDU7QToqbU43sr73AR8E/C5KGnsxLtMDO6vMPegOAJjihbWEYFN
5yRp2zPHHA5CqX5Ndh6BEIIB6QaP54TCm6QkHXQEXmHHZEeEHoBAtQEhvKHYRgOz
bOra/I2Hz5K7gT+qYs3q6bablVjNz+rwys5Oq7+W2Z9Rih83f1JtuA/VfdLe8aXK
7E1MOOgWFViHdZDBPRs9VZqz+2cYqsvYme53XOPG/r2Sq/P4l/BoIKZb/Vg+mG/K
8H8hNeuRYTJaaU24SOMVJOaay4LeOvZIFQWyxTRu45wir8td2YNfU5hK57FHxyVh
FqZmGY7fJ1lblE+fTn0Kpb+YhrQb6vZ436PkHk+0HcHdEEN1U6J2ty1Kdf33eHai
kDbMqVC9DzM+XpspFN+OqcFLom43TvFwUiEDk2+VrHE2qEM6i/rgwkJaEG5iYaUr
o4oOliaMvYxLgD8DukjpiaGdT5ygjX0qeX4XT9HrnZEZMiZst0cclZgBJNcAKixa
RCs40Q6ardRqcB3ZW8eCHE204cczVCNZl0Vmn2pJyYTCzAsq3XG1txQ1F/XkqXl3
4uzG5XqURwbWBQVECU6BiFL5iEEpN/OARIxCZmVrJ9ZTwucBwrT6+SPMT0r40zQT
RSxewfNPBJQ5OmRCDybwNNP5gPoAhGV15TYMadZo+f+hyD/URGdulVzBUH1dodYR
nrNdL9wjmIxML9Nk54Z8Yo/0LcscmwZxEiQKpieJQEzj18o/JLJC8XDC+S6qDaqW
LceV4dtXyoJRm3tcV4pHw1nL0VWnhmukS3ejfW01Beohhu2IIdWyxT2ixgOBGxcn
8OlfQ0vbNbPRr76LPwDbuRF1CHLHZ9DWVUrw9fCVtPBFVbh7yfMrWwbQ60ns8+2n
GSFpH/a6ztgv6aizQxOrRVIVRw6Cb0wJdV7SUjzfsYrxNi/onHcUCCoBYkfgv4bm
OFS+4CZDrWYvNlYW5Wam/bSqs94LSrHhS15WWkt+M2lXGag/oTSgVypWUj6EdbIf
MD06lY79Fi97fCftaLNZqXe9pivKtqnSK5rGpB9Gamd1785LGcfUTWKA8gN9GwP4
SGsmMXAmcr8h4AsoNtrE3Wt/5OZhSgY7Z8h4zBU91AhbsxaW/c8u87ak+Re8wPC6
6MJaukWwIpMn/sq7jDk1wSWXLrZF/yP+zZLsInIW1S5lRzs2fGOblT5lFM9AKjGj
884XBq1BDik8Ci2gW0d1Js4bXvwNIuwlmaHdvqMCboM2ztybXuq8lO2jDJVP2Cnv
yyUHGz9rd7QQ0YsEKKKx3xK6c+gnQQtNyuKUaoaKFKJw6p9+E4CaFx11CQmXOHut
M0DKIMyIWV8j/qq9A7cFtZlXhcTmDRScmmr1wo6k3q1GmntJkWnxoMEjRHBP3k+B
VaTuyCQi7iOgOicKVi+Z68tTDtNf8EqsMhFL2navNPX1VrPBwHMbDzQ90U5gvoi1
oeTRsoVzJBX+4ZYO/GFURH+GPYU1U0RyH5GbgsjFdQRaoSbO5JaG6paCzza3SDyZ
pSYsMs5QHxN8ZYfW5CRGC+LPf954g3J4DM+Qedd/RTfggSr+p5sf/gNYAS1YUWO9
IegTRoKuiaxzC3AZw/PpCqnyY3J3ltfsBKLA04TmwZSB6obPobfjp1L4y49rPffV
VNEbAGt5XUOdp51MMRhakZcGH776IR9dZPLb5XD4Wej7kAGx2cn0HiLUH/g9PDZK
EsmsQoMFwNOAlu6aNl9SPldoZlICR3x/Te1TYGkfnbNT7mMTZ60Sy2cGvgHR6rrZ
vHn/XWsPBCz1MVo8yeNX66T6onzL8lbMrXtZz0d94SInK5oGI/JJtzJ3o4i3anQp
1EohcKIbt7ndb4Y2LV6VtJG5LcZCIsPNZuKXlVrJNh+Xwa0/i0GAar88SqcL0+P4
BwBYf6QE3RzYGAuN8ndbYV+LjYaxVuUmoye7F8j/G+6qKFx0GiY3x4tzxzWfF8Cz
/oLM9tLG9fla7WicGvA18C0rFTQ2bflh4PzQYVs61Nr9dhAAMB9Q0aNECMn91c2g
ztTJXux3yDuXx2fs1uEqdcq1m0rxDEKEroKxKWR4wrnPi+mBcNvFbi2scgJKW0QM
Gz47TDHXebJxpgw8hsamhPsoE0J0GeEKBB8edn/XznJDE0+UhSUwgjeCPChY3RO8
kaIckhQ8hgei5ie840DCkuV9BWexUKub38F4uafteUxE5tdKPfKeQApVf7U3PzC7
mfBt2u2uxK6B7LckxYF0vlyyJcpUBCxFhxYzkM3YYFawoZ2PkplpnvbQWcLMIqV9
+nKsn73bYKdUJvI7TI5jFAqvE32gT1C5jznbvFyoY6MvSzO7Vj7QVUglELvOjWjV
1KjKql8gtwDbaDBxLilrG85GhrpSpvYItTSkFEyVCXNXiEgU+EtHi5k/NxAFwAFy
HN2c2fEyozFU0yx+2lkkb18REVPHfwUPZ44JxLVfw4Emthncozq+++M8ZCIDm6gW
H26ZB6Z3wRDlMUCDGTG6DPXAeQz0bJyzmHhhyst77K+E1BhuCOsavEnbjRKlqnn3
jOYYhxOWWaRXV0XhLEinM4Lsjpo4+yzPYlpxD58P5AlCpA1qDzL07SG3p3y/8jBq
d06jRRLD+GLcoHeAHjqSAUvaWwJ1mcKMvfUkmSqcxYU59iLtI8VOWiIs8VgEZFtG
ETVNcon04maFNr20aaFlOV0emPhdP2p0ZtrAjSZpgJpS24x1H7QeBa6DOyGnrZi5
F0oPQdbH7pwPHnxGlJoevFg/zCl0pd0nCjq/QcEfZI7hDirIvKG2eZHKVNhRjh93
NFHYm8ZZoAyRe/F5sj/lO48lyTEijuFzuGclth3K0jV2JZYVb0pWDuAuaFZTJt28
9x1QWkBoR/l1jwUv4ZuzMNyK+P+vZ1V8/4M2UFTP3ky/NTPQ/qJbWiaHE/u4xPup
86I6Uyx4I1FfuDgWbHWRRleuc4fMfdMOdgHPfOXN3+roctJBexdc9BL3MUh3L7Z9
R8dDi76r6etYrd/pbrEDzNARNkHiXOmEpybejsuSpcj0RFyH2yYrFTuTbac8/zao
wKsqqEgkvum/MsW5ntlyjBMgNV3T2ALu7PdIKu4C4noJ71vISGSt8QHYIUVZnM+g
H172d390wrKhNoRLlwrXdKzZ+5BeNLoz0S6PGdRrZAPBInfb1TekCL3IzCf75WSr
xNbmkGOJW6/QnQ2sEqTcp3hYrQTo5FkGzX5vF42UbvEg9A1f0TgrJxMK6ZKUo1+f
wmT/0l2PMWyUZmaycsYAoU5ZmCCoKPK1hvCacoOplOjWLV3wIjWPt605lI7bfsXd
Ifjg3pP00isHXrg8L7ZJTlBz0cEuQXhRTyKPw+R5FWj7QWDeLrIj1Bh45hqaP+au
/34xpDTowLwQR6gJjVdI74nUlczkHy4CpFhSC5mkMkJrwIoGNkq0EXBDp1uHVyaX
T1Lb7enLkLl7djogUnj8dYz3tQkzMwdOYYSyl+Q6LebQXQlplxNx7NM8cWNHl/lz
0NLgkmuGVf3RdPEsTqVutKrCouqlC62gelzuxgajEjtxnQShUvuuW8q7TeCOf901
9lO8t5zKGop7Z1NH4PNTjvjIKUbsf5yGOYvoZKf0ARTPCwfFY8qnqUXyOhxtDg5h
gVzngjq6wnsVfW9ooZBZsNUEvHMPsDXjzpk5xhLIdcvcNC6CmMyy/Yik5/80hQAh
tTf1yURIY9nXmqU2hnLBIV3+TOubj9L9526QXY190sij6iuIbEslMprhoPh51RZF
sKk1HV08PVTYHzrBOlEMjSKHaumVGknUCQSs0Jb7zP+9BwIhjHdTBY8ZzRXqfiY2
Beq3+G0/eG9PfF1kHXfUr5GWBW5B8YdjdDuOGjNSWeMbY6EbKViKFBxl25W3nj0H
c9r0djTMBzCUy5LFThdO7sSQAMD8W+W6R4G9Oc9th+VVX4zCN9g/GoBbm528G2Zs
O74Gn61lGShr7noB5B1zncEUZ16YNFqypy5RE3uw9hmUKSz/zNS8DtCFZt/gZqV/
2ueEIPPsP1Uh+wOPjzkGmmpSAq5JI7YBAa720kS3f3ojsX5i9YdTX/Lu5NAd1izE
HRfod/jomK4ZucgKQ+9Qtm3Zo4cWqKUQ1yA4OLkH57OYeP3kOsDRbPgI7RKEE0+4
5IIvguZj//8QocWqnp3JyG/u0nSzCycgs0ketYk1eaQ4I/jlR3lcZYF2TlJZmxiZ
Ngs1D2aX7nIIiCWU2qkcMKHLYK0boDkKpviRusH7C1cTJlfpUKdDE77Kv97bcZWF
f329/nqd3hP5XNsL/Xg+4UmRQ68LCuALT2tP9hb7aZrdfEz63xZhBmi1/ynFZYkA
dDc87yNKSwtAfdfyPyGb/lLezimjk8Kb8WWbmVtjF7li3DBn2gnt3chD5mG4Absi
ZxSrGn0E0njHNCdCqdnDrHsu9d8TuxRCbiefN/w4aNJoDOo+aPOSrxamm1druPa1
0pQ7o+RIzXlFekzYj33E6Jo8T0jXtTtzQ+zZreUcxbQN295y41aWYmJsirUEUAzM
AXHF4TeMgqLdalUxfMdHkm6ROJwA48qVsLvCJkcRBKuRpTsIm58k1V8NDNQOcTyw
bmQoA3PQH9KvYz6OWfJ+YuIc2A8JhnaGtfOBbLlpewedZddbpvOAoK9pbYBdQPdi
R5K9AEzDsLOaN0UlxQUn3tdSjairc+NcfD/AJeXax4w6ix1yXn6x8ugzVdCLmsfa
j3cFtUNw4vB2gGq3RRGEIc0qwd6BUP3YIfs980AD9Y7ISFoVBLyT4zf2/9Wgzw09
nwjrLPL43SqugEoDMdVp7jQaI/RjAO7Qn/1og0n5U4yf+NM/hR4JFQz27oB77dEX
WqO9GM36HzNfVs04U33r3BT2bhaoEedQJCHDJqySv6ykanqJ7+PJBW3ETr5tGZex
zp5zhUAWcF0UwUl00+CBxkkHj5SGJU0tjseoxjbNyDtSEtBKH/GAxG9lCOUSjQxE
j3MSWbfIT5l87NUCixVr4nUEdyGwOXbXzGZflRgGW0ytdSMNBsp6k5YnXsPPoTkJ
qKwO3moeCcUXyDGvGXJ83OvKqkm6ukQL1bdLsM7+quByhDJbN995y9i5/IsWZOwP
Ex/yJY1i9BHeEfSTjGA86mT5hIEYnGZIkWOWPC7UJfMcotB9YdJ33vQlwfSEOFmo
1yeQdsYjj7doTIzMDuUAFI5A0M4Uc6esmP05KcgcmLUYd4taX8URuTMnVqUWJRuS
Su2ebsznuqEXFNSiZfi1KNvnHa/K980wnmj2dTKXfWcuM7O48NvJCR+X+IFL6JB2
2zn1c3thALxuqqoHHbrzdxAsgJT76x6Nq1yNdqbi2dXiq4wNRKy8F89RwuKicRIu
ZK31ltezhlG5T68LK6a8vnQPCu9HDTFElNnrGX/Q9sI82dsm0VgaQtbQRTFalM00
xfbjJ7YBvKgSed0yoytjnV9rClETctAecdZOfsu1YQKVB6JDQNWhFEhMgtQSXsSp
HImG/eIAdv1CQtlkE7lvpsGXl2MzBtxoAuLXtx1Cp/6jeusT7cjLZ51kV2ukb2nN
eh40u59wg8UA9Yp34OPMLFr6w9m37kBJxhUoEPf/TDROwZP2f5oCSmeP7o1khyZh
n5XutWtIOYRttO6omz82lH1hvOiyifTSSNvuoMQQVT6l1mV5puBDKx7DmcQfMs4Q
zzZcjfNOoz/zr9IGmB1KygnIjlLlLCe8tK2QTM6dWzNkmErAoS7GFCYJ1pgJW/Vi
PVyPgqref299Pts/3ZEttRvSsr/OBj8pszYITzBGso03Ox5PTGyDVlQQCVAbZmzN
iMOZt/Syy82v/qhSTcN+1C/rM/jhr1LFnPx8y07+slpJJSw24QONRnm159kMovVV
0OLBCeX2vKhjSPGO3HNT5caXPpscY6G5TY6U1NjdMeqCFi5AEmpupUHhObOfvP+h
vDBy60yqscdh8MtJN7E+iF4ZBt98DQifQJxdfeOIyXawVPS5fTeg0+23DITzr2BB
5Kdnvkt81xYK5nD5CK5Ql234A5A4VYqJrmKEhsVI4ojanXv3D1hMO/JAzKHVMJjy
vPNrYr/3x9LeK4dBgRnOwLanejJJ5IEuGj+HQr05Wuk3lCs/Ehy2DomN3HLhGb3d
U74dlNraEnnG5w2jWl89m4uqCbb/eaqI0GuKiiOOpa+FYoE273dtFo88uaPJRtMc
u1R5A5rD9VjQi8FX74+3dRKmksVLHERPyne1MhPzwRfwvUynQ/5B1Elb1AJdWac6
UJo2aLpXsHJ1ru7KdQ1nYr5do6jVStuF+qHJEfe/8NQVJ0AlSHLvAHmcfK3NsTPg
HO7Q52pl+pXQeI3Sajw4xRjhzMXCB6xLHgN3pg9311lp8QfqN8A2RD0rJEIQfg5Y
YHieW1RJu7+eEztKXCh1MO2bcqFTyYp3xEmwjh4Ci2i5pA6IOb2KKhTcc/7TS5r9
eyS/CCRuaUMzRzDv9zUTcj1QUzwLivgx1U7YQNKU21/EsKPZBOBJMi2eMi1ZFq2q
CLU+Bx+8L+nNr59dIVQ2jquSpbNa1e1yiHZA2TRgXJF3ymMNAzItYEcMIw8WZ9wT
Jw37tzANrF++FnOktiFghax/L4xaO4K/JXEq2k8VU/KCBbAmgIdRV/mqdUiCo9LK
PorlVp5MnmAs7Z6DITwrM84zRoINZjbXoF0XpunQG7ClMrd5ECkjs+D0Uws1KSeE
Q991CoQEamsSq3to2+aKkZfoD7CnNcEBBwyHE5aH7x2vQitok6BKT3L/dBA8jlNK
Q7i3PKL73Frrx1sd0zmeIL1O+Nc9WyCH/uu/oAdzLRURJi1r37Pjvsl/nZS2THOk
+7EpLsWotlCjSzFGZJfb9QYRtBbEHul4XP657cdr0q2cjDaSLLKZ0cdaTN3WFv/H
8OlryxOQJLRVz/69HnjLdIsUZ83jE3Jj7YISjXuRYHpfMD/aX4N2VepSDzZGnyXq
/R/2+vpTUnWK/zvZDSQAs1cnayOasfSjvPao/0aTtC+v/zxgO5fcITV521m+I3JH
BdktDDdsWJWH8w+wPPro8fQ4uQ9CcQt+0Sl0KV7NoB8SZmmmTCLYG4BKd6FI0IYN
2eSGpx5CiNImoUNn94FKcz8PlxKtLo8hyFV4AlwTczqyFSuQcZ0WswpXuOXaVg+M
/IFl4LpPxbiSTKufSc43RJwx5nFndCVkW0RpugrjmZnIwiKThQgbb32GOY8brONZ
KGIhNhK7e/TezpOLRhJpAqnHxLl8gD4/IHfC17Ga+fWIsXwturVqUYQ9GhstYirr
QmipoSZ2nDthyBNxUupB7aQ3O+rW8625KbDouITSU33dac5wlQ/5BnsEnPbnbP0t
zHBsn6fxqGCR+PF0SmZo1+0wvwF++RUSnlABN4ckt510juSKKkBAPFsUdB2hO2/T
vyY5C67dE1NT61D8zB6FyjQj6SdcoKuSjpz/3H7uc6nGUUCIbQh0UlD0ypaegkq4
0S3igTC+RlZ6LVyVkZ01IWbESC90F8ReouArJAY9tYzmTsA0fjBSfjnDdM3gzSgQ
rysNbOkUzSluys9JbRmK11LC1OOHfjyan+JqLJZkCmdvxvu7CjiKdG30ehtoUfWT
i3KsDdK0K/dspYS7XT6QEEWdX19JaHVLf+4/MP7YmC+wa0S80gg+HXsHLTubB/CX
gjVMR7unjM0j6fH11s7APb2Wm+rTQa7hlvGFmjwgJJy+sQS9/FuhIICYLFcfwNDs
aNt5uQGc/cupbDzc19EVTRmzTFM7NTJKZsbIRW+yV5fbm4D2CSxtBflBn7jfNsq7
Mb3DBBTfAhyZ4ctSJQ8TI1e7d/xyhNhcXG2jffTkIonWmEYU+h5XpuKnmha4MuRA
89sxgATDLw1cqNM0YgjGJJEJcz07K86kL7xW0d/ce3ckdy/O7WDDeEy8pl5fj3Kh
Z6JZ2qwRybvYFHygBuDKDU0mNXWHqruW3rC6Z/Izv/TYqFvx0YDd2R8CA/oVhKaZ
nytLbvWU2Am3XLcT/a/oQe8nUN+6npaa1DBzqnSLT6PJWC0pIbDjhsMm3xShkC4O
dzB5BJwJEnlFGD/uTXQJOr2ERDIXT7Yf78X1oKzVyeDb2i/GJqGU5xewDwTH4V/q
oTC51yqBo6PqIwSEmZ4BIWUBwR8oa6tdwR0DFoFilyav7SYvry5KRrIGVnY0M9Dc
/ja1GUjZ+Sf7JvLggot7prGLMIy2OC83a7zhwyP6EAR4lmYPDcf7bqDMttK1gVsm
73YGmug9AQxEDjpEogzq5nDY1YWI56nj+TTfRFpRj8h0H/6+9aSUDTyO5v+9LJqs
on//tO1+OCu2iAXs07eENylwhUDNAj3zcybMQeQpMKXht0KzVyYm/v4uvC8Eh+mz
2rv5+SCyuNJIRAZATQ5yg22xX1e1ggmmH7MRjUvMxXagqaihmRHCTG9ZRdTg816P
XU4W/p+kdJjAdF2B8DUP5gLt5UAoBbd4RgpQp9XcDZzcS+e5L2czYtkfGZPa3qtn
rLyF63pAvKMCunHWBQ+KuO03D2jsyXkb1nw+6V3Qpwu+uZQMeJQGOiDKj1RtTWVA
wX2HpmaRiJvwyysDw3jq3s3kMCSf+wLsZOv0oeg9Eba/iFhoGWaNt782TeSQ5ZMB
CqhubgcoMC9JPfgQUVrAvNrDaeSHSaJOKel8rReqMej9a7hDsqv2v5cziIwstoQD
iDxgnlnsgT89FFMxJnSBXq2aoPkzEdmqfm3OdUN3QQ1rnne5mF4EE96jtZ3LkjW8
NALbXxEUWHx2b7AoW5Z7BmVSWVuzYh9b/ytbOBSNtXPJ6uZYSRZDcz6DzqKwaCnV
z3pNOQhK/22XaXUmOu2gjuzFhp+K/2/kEwDxMEOB1TTQ6oYvPRO+L6zg0KJp6W81
flaue4xuzARxvAwoHdg3IFGnYmuHMMW3BD5DBQQCp6W9hfZESyX2iuCQ0B64wqWs
Ex9IDdLqQW9UicNgeOJqaASZvI4zzC0f42W9NF4RnhVhmLlRCFvZ3ijPVaojSGPv
l66fAW8El21VL+grDeTICHwm2yYjC/Zz/p+s7Vbb/KVhuFrK2cipJrJySd8My9rv
V7KQR9LrrHyiL1ix0k2rjiCP/C225/pLSAU39jcOQlAkPPwHMQEVb+kB3tAWXbed
u8y+h+0bfeFWpQPB6kA0RMgU0N/XOhzpkr/vpeetix9MZTzPExXEBvCNT0VBSOPe
Z14Jj92HoHavfRnKMpzbvB6KWtRbGfvULUe8tZSxsOcoKiUSk5xd7e3XqkFEaQWS
V51m3tQ72N4yebBeOMxpiGkP7WnsaC7N7FkGFeWDCvx/ODRUo7aOvems/Eq+4KZr
vXzoPVYWC3uT4TsFSJVcA67QOR+F+M9+tUrBUFGcEvVveeBGvCKPg3WOcv/1Rzxl
hTRcu27HQTKmKt+2PbOTgs7ukQdKZ1rJDL9c3uwBFBa47RYvPyzixDFdVSohgNKS
nsZ099ONHGBUsEftFYMBPukKITEDjdg5Dz/7Vw0Fsckky5oHHBgH1KX5SFDRAEwn
lXUPk4Fp6wX3mXIveVToV3S9gyHhT1RBKO7M7tEJLKYsyQ4Dh1p1ztLK1NB2UHQz
kwB+XPj/NOfMMpzVUkuQBmkbby6fYWcBcOs2FZVovPayV6DzHeb5vVLex8Hz+Xjm
8busQn7CBSCGlCu8839U7BJGBNCYHtAfNFT4Y72F5wTtIV8YZsNNsFUx8v893r0z
5Mn64VAsp863HleOpUFnseKZ7th427H3MVtTxIcTP+syjgR66prlz+33AbcXpbvN
bZwFGIlbvzOH3G+6l1qT7fM2FbQmI20o7IV1tXQPc6w1F03hry4h9vT6BL4Uz9Tk
ihxKs48W9y0mQeT0knT+pxhMsMC+RJnzxTXV+wkllg9YD3CwmiM0xAjyotHCzQJq
IIojmXPkMHZLmKdFEhQQ0qUQTAvCv1FpVyzIeRpQB6VQmEpKiIPfPgSX+nSXw7MX
uV4VCV8nqcWmJm33GoClkgvK+8JpxA/SSLZs47tRGh1N7swcxKrxngu0YLCCBf5h
KPd9RsyLPeIgkAWh1fO6+gEy9fh/8Qu3pchhdGzgt59TX4PsXIQAxxyCRD+H/4Au
UHkPO5UghIjpaQBOVpqQ8rweMUEgaP4uO3HlFF7Rcp2M2Tu303+mRVL6OAyl386/
SxnGWe/aweHI8A18uJJY5AMbtEKmV/qx+lm1xl3hocN3gnMXRYvIEi52FFvI0Ws3
gLlicviCoYkoNpEqaXQMg0AG6NnSFcum26fbOhrkJ6g56shftyuL6FvKPshmzIYZ
m8Tor8pXr40pVV4aUdLyuC8hb10GhNOzw7eB/DlJYXA5ZlI8B92zMIFO8JRFP60p
ioGV830mlT+CIM/Qv93V0AxQSwO11wzKMXnC+vNL40louQkAWw6zaPihdjpQtKc+
Z7b9vHoH6c1watz25GGKRYWN1ppU4Neszo+5tFeBjuFwK/tAYPXN4V01hilYrAzV
H4UVYa6BujLl7CxOC9nGq3RmGabctMll+rvuwwl67oXHRIAx04YaSeozl3p9l+9C
+2sFZqfrkhLukGl9x7mb8iAm4ffjv7xUvZ5KTCRYERbiWVJrDBW8uQ6ed8lM/Lag
3+R9bTM5HWgGQvHqf8OmQCcMHkXNdhme5f4ah5OzFnaMzTtU5+jfjSGYrSvMqhOd
xzlEwVG0IK5VJkyGsgkaZJ4ZB9BTaTKD9lkdua6qECMUh7dL0N0Hvw4FBBEsrWu2
f3rKOJPJcTg4zS223QcS44Z5xFMsr2zYtwUMAE7ZvlguZyFYfxjv6Pzod0nzLUGh
pKBDCcSKazfWPt4OZhcFI3CNM5E0H6NdiTvEFFYFhB7VhDHgq4oGQ446KTujFPpP
71O+DKg72OBpAS4JrXVe8g44ANogQYAQOBD30GR1MGrnUkx1Uc7dsI7snrWuP51N
ZYqjrxT3TbGz8RJZ2hLCI1Gey8CfPc2YOPkD5QLGbw8Da4N+48VmwmT8cWjBxaMT
iAgI6TNpY26LWBQ4cUUMoRenfTbVLCZu0otwowncMjL8Au0tN0iNzwPvji5TIoY8
cXug8aedjs1bVfVWXHlDoxEhHQiia1StNEIar0Rci9DG9nlxlbR1R8bm4zXlu6oc
/GX3ea2uC0b0Nxkd7l3GY5ym27ejyvXg2+NE6+aehQNkiBfhMIWdBd0euEGYdIB+
whj7rHUK7QhhfsQIxTNtkZC0Y1KogaH0yL/KTYk7AJ6YLO++BVESoFWJdBDruyql
zb2oyP+GMJva0+gAoX7RNTkCIdnFd/RiJZwBIpJVHHjXj0r+5sTQ2DDXoGKPu3lH
w3SVU+v1jDcq/A/utLbxw1O0sveVXxn6BONg/SqJ206qggXvLuK1oHDroMsHAg/e
VIx7x3ORcBrmMpdXcYaWBlXVHIpa62FIXhpAivgIcMqodsI5/Ki8PBUUDpa3UgRF
GymJTV8SsOTaFhOoc8LchjgkJBAzLq1FePQVL1tm1dC+nZxoC2nCc1rKyTLBKoCZ
yOuqGCyAjidhwWW1i9FB0xZdaaaaOfRUqvweqP9UgGtEjWYE2FD3hDGrT7ozwpNC
YW/m0XJpHbVDLc92cp2J1X5/Tp1BGpUbgmx0+R9wBhj/1yaDwokeGKbx/Olqg1nL
ZMvhxxdkN2Yp7rv/zaLUqgAldG9vxOh7Y/CUHWwKNXvvcfNv3dFEpR+nP9O18+3T
PejRo0I2e3fYPs01+YiEH04fvC9/iP35i01Xgzo1W0gGhzFNpHeslHo8C4v/79LW
r56X1NM7kHBJgcp23dJOebHLQIYoSSvuKaAJk4s6+mfYc6KZbiibIw3+lCWMGIRq
MUVx3ks1/tCxU8KaGNOv+gsGw7YmL/1ezEdsL3q09tD8kUuzt6NgZkklU5Ykbw94
GdT62a16jL6NxXc5WOOO2SKx3VNG8LzZi9Tp0P+OmLRsrvpjG3cSoHuh/nilm1ZD
zuHoSnDYEx7FDTwTVClItdmMpIzutYNtYl+eY/IrffAAX0tqptCZtW8FEmEVHUML
64oRPgHwfStkNPBPS8+x9VX4oKtuTOoYzXX/rdUSez58h3DkvJLSmDl47/+bndbu
XnOdiAE8p3mLh6SltCpJyrFDr7BLFjoUpBFmr+qdH3/HXBdr1kYnr40rWWHlcBv8
PkdSk5HAi/kxWZn5Sc2rIy0B0+nl7SGXB9Jjh6NCSiDjxFN7F4rzUWJsWlgD0WmC
10GMkwEHi6+GWFmqqulDrRGo+b+uRn5VqYqb9jrqOfMmdR8tSDfqMF4UD0mZ4JlI
fuf9f54Djf3+EihuKpx6/QHQ9xnctE394JHtPEw64oK5/fcK4FHjRmEpnhBh05dC
j5Qsdw43qoWvOWEJdIxAfcZQr6OnrruIrcSrWeVK+SzGn+VUZxfHxbRc8R5ZRl02
LEtzuXVdmPayjUNab+uEHUa8tcBssOxZbYgszPZrE2BW7UM1ilX/AFuWGc+QnKmA
y7A8qjwzvWIpZUHsAoHoOOQZcyJ35PFnwxbc2jqVDNgRZ2jZDR1Fw6YPYQ/3yix3
MAhzCuDJGXECQbcLwOupdqY9i1h2QuKH3wKqTlLRZ0Rqu7zXp9S99IPfLFvRJi5L
z56FYAvuiICZ0G9tjROwvWk6+nz9LUnjoa+X/xEDmPprTWQAClWu3Xpk2lrviN5p
+cqW+Gr5nz9pf3NfX7vNLjPrfZrTfcOIiM1Q5n2yILrz4DhAjAOxXO2e5wr38qFj
s+TbEan8Dp76fnfORN+mmdzHbmuc/7dJIqdsKyw3vH3DMluxIsvYf5AW4n1e7WXJ
iKX0EBhJeXhTxbQT0LDI3M1jJzmlz5s2FjAFfZ6z6CgYlnz+yu8YeXKaD42933aC
m9SA6D23Db87DpupmuupSaCmIyZ4/QLBrkh2GCbJCJJSJUPyVmSM1VR13lJmkTya
qGPn2zMym8dGvKZwdukILqWbJ85nbRmfXaXN8wOypYgvI0Uyrz/CfrTk6VGmIQaH
M/hdH637BiK1fHQEngcOHjmV2PMmSKJy2i+4Hxqm41uC2LnybMMlgMBtICrgLuyA
TgbPvi8xc7xw09Jr1duME65gdFib2R6lQEedelyIHJztxuV7fp7hXd3HK4wLqbOV
gNbZMRRwkRH7kBCHDlksBEKiGWrLYT6l+M1ExBTPNJdilMDSQAWr8CDUkOmYVt4y
+Qeg4+XHpGglsQpTVDQ4sbC0jJExNFqx6oABj4kmJJ1e0GFoPL2hZsut/Yf8ysJn
3ju43urI6JsHZIetbJW1YMMc15vyf8UST4p+s4PR4Zvrbuo8u1zs7LWCjU86gp6Q
or2HajcCj7QSGycVuDMu3MuZlP/Fn62cEmHs45t6tjGEzWwEubKXRVmtLAsO200a
/NP2NWl6A0NwTWvTgxpHrUneWEfCVw0Ye36VlIRJmwRYhzYG5UJlmFyJpwaa29hA
HiEmX5Mn1pibauHzJ66HVub2m05ObTHoI6rnRZymSuuD+imxyJAArjPImlB4xhRL
meGrfGr+uMfBrPOhmyOuaBNwnwcOrjy2AVup8ayq8Mc28FzdcUEfrhH1Tg2yUqM3
8ZFVu4EF+FYofjSxzD4iuEPM78nRtzOwlQbtur8YmniWBeXOyotZjTK32FzcYcVN
rpT3SCfgy6HVkCz0OnYl9aPRFuOuFFsNVO023kAr+On/ER2pItgvZPxyScvJcFfp
z8GtpfV+8tbQQgCPbGcczpLauCo9wlJyUqxuiBeNLcqJ1PQqwgPvxWd8nnRd8eNI
NWCCjKUlQgn0Shbh9IEJ3rgWH7Fa+FQqcRahUZbt7UIZ2GmcJAniYQ2DvRpKtmsG
4h8/yFJdNUEsaduBnq6bLA+fwHIwVDawUFEEp2wQImwBwQKv6Sn1SE8an5ugHYzD
Mdp3KzPIaPfgRdvhN7JWup8YR4G+tOqErwlNEDrc/Rr1Kr41QueGoMgm8A6Vin7n
TaLnGsnnh7RiTuXTZxIT+mKRY62+7LVn6AReX9rpSiUY1f8KIxvRjkVj1c5dE+qt
CeXNA4yA/p013xP+AwpjfOyUO4FHdH5SPs5+CI93mms58EddlbrgKaGZk0+VY8Ri
q3J/hCrkhsg5iXvtUlw0fu3IUUlCIhfT7t57gkHFgEOLT5L3kU4DULcTZT4x7JbX
shloWa77ONHLFqVjG4Nyu3v0Du2X2heQqV1wB/fOw0m/RhtdNbmDjed4W8G3s0j8
Hft0Pw9iO8+U+nlcI1cCtFAZNO7ZVNe6+UaBjumLjmFwxsQLD2e3ymLQt9NKfCkf
RheISEJMRZxJumm09Cp31NYex4DK6W2XEa7UB90Vazd3hj5+vSPm5Cvyr3GjvUtf
WYXoMnnOkoqUpgxoM93WDENJ/Q2CagF6d6ok9fKgqjK/nlpBOFpPsGNzur+5bmZp
Mt5CMNZAre+rtj2jTmINJjjSsAm6ecAQWasFiIkzah1ppjr/jimnea5VFgaYX5yi
Rw5Yz5p7mR5gXsSPdcppgh+Mp7RJWmbxR7kBS7eoB82TgjGU4p3WjEpFVUdWvObU
gYQxEQsfE+p9g4ZVfLjR3FUDnAwlT4pLNbIy1Qe8ZMzn5oar7NGeexMzsWtihbdU
hNv0y3sz83BH6o36KftzfwgyCmPK+C1wtSRK/h7vji1taskKW/4ROof7oFGo20Ky
USP77Kjdg/XKXrGHs1xe1Et9aEEvCrQix8rQQlNf+eW6VltMcdTtPZ7bnKjKLRzs
MRMY/FQCMpg80QNHyIVdgySkszd7Hx4OnMOn5UWymwCoLTnbcevZTzugvaG1cvuY
iWaV6EprPKOcgnyqodu92jchDe09lCKCuSSvldQ3dchnZZqx1vWoiKdqlcpFUmKA
SLVhMbSzATiq7YxHzz7ghDDR/2/oaLSANwtWImFoYNxOZPlJkbhUuY5hDSSFeiYw
QkYIl0UT3zWvIqjrZum9wSVtIeehw/ZaMTxz5+K0mSCKSBG2gmwo3ZqnnRY1kD3X
f/s/i3uypDHyyJrOQ3GCBRrjjD8cYka4sf5XfhBsqYp2cGbaZ9VWA6SFliGgiKYw
/M+IXL9O6jJSW33WZ0LxAsDPaJfdNV7kjBBYR9nqlM8jhThoANTZbJCM8acyKnEL
aSQnZxzRZa48UChDwGEiO8X1SZUdxnaJyXSqcQTZnbs0H3mTWH6HwAsvvgyy/B8z
XMPWhSwVve+EFg22QGAfmfTFBCnWwPaqS8ygrHzZOq0osodlspXHdL3kVwy7EXWD
HD511I2Pc4DF7chNRcdYRayfQZvRDEiHdN0oDHjdoE7mTQw6wFbIs2QSAzjzLDQy
4UxGBXVDFJ1wNXwjqMzpytuZAoFtsquVv6XocdXqMnmAS+m/YK6kM6LWhgn6d+Z7
GdTENUJqQ6zm9nyDhZXkGGJQwlaIkKMUPNzIc5vmW12/HNT58wPrQtrgRSleCQYc
UCSsVCssvKggGAww69RnfIIxEeOgUZSH7NJyQY65aJzJCM2LGgyyydLWsIzPXAnU
xTOvG+K/TTYUqdGBSbwHlQKCwEwY5ROQ0HOhrZa6bfZxTUneEfUixJ/ibdnIz/s/
r+84/WuqaGgwUdD+F5d0EFPbBHVMyPmCfn8uShGCYL0DCBmv553G7kU5Sh52v4io
V7Va3ybtXXJfWEEHQJzAR0pQ3kfQo35GZyPu8W332sz4oF/lHUGclsuIXyl3Lcky
aYgFRnMhZErkZ8KDFx+i960X4+EheiyGYmeNZC3JYZNya/cIDxUPK/MUuRdA/sx4
wGm58MS8foHHh8JVEq+VDwRSPf7rk5fadBaLjm+Yp09Pj3XGZgYAlbpNiTABkBfS
sCTJTvn5JZZnaGmwPLIPRPDzBgqyb6xueli7MP3NNGh1XH11bBfMQOb6RdJuA+pE
m1y67gbiKwJOXY16lPMIoDiJqB0tmEzUQroqPM5K5sJdc0aDDvic28kzf2MClUNY
q0llqo51L4iI8EQCkDUO2UqLySX4DodvQZ43Rzn5JjrL3+QsgOmJFV/alFnyJyW+
ke1l1ao0KSF9obrM8SBIBxrCh1qq10BWgqw0gXIDtdxsD/VyMZqP8aquPUxXtPcG
mXI8UBBpXDvGLlRp0wGBI19KVjElx8oBDUktEs4ya8d6BX4RHMm3NhK63y0N+e3C
PgSjokIlVES635w7KrddThgUZbvIrOlmFazk9i0lDeBQlyRK6OdiXRK1pdX/XH/I
zVa3blKDC5mirO8Pbi8xIhdD7pDduylayQ7uG2ltG4l/5xImbUZtzTB2O/W0pzeD
eu5T9DPMDiJtxGfJGPWYrZEnKFlZSziZEfqQW2wmDP9YLmAJWTlwo/0BEXEhhfQR
jQbytai+IXtveqpMQkPqKntZT0QSDUVD6kxMAQHhMuuDSbbmjrsyCY9/OOHWEuG+
c+KNq/iBxwmObzJv7IJ3mCLyxSMCuYNkDZ7VBAhj4FoMBW815eInttkdHC7NV+UV
fB27hixornwjPKqkdk/zqta3bqEAm/0YBq8FjiRvZmli/5oP8acFsbHvig5W+Kjj
HOnza8PiS5CiQCh8B7zs08qC08Pk1WVbAfbSRpHgm8Idr8y7AfJkPmIuuudwUxvR
b1SJSOXoo7kPlwBXkZPXKljrywXH2JuONyMcoFIVKzJWEHx2teRqaQaLyPuVvzU7
JpAkp+mW3+A2DCJuZ7o8r57rqzbgNAqrlzpOiXN1u8YfxwjCPdh8GgZu/Dw3cxVv
zQol7k9mcqSQLkkkM/9VO/Pf07NzVwhPqChSr7efBkN/+Del87lL4h/iHAmaSXwA
6bATxF4y1SCL81IFAGBxi9zbZvuEIzy7USvtSaMPmvhhjDeXGzFvrr6LcVH8WzbP
qR3/530EOmLkiJoc89SDLbTKThBlp7Z11ZZkirh2mIx3e+HTx//3XYZlt2j+4q8f
jFs8QXgwfBNM5kFEwrneBHP8ytisLlaoFUxk8InI/1tFZeytfCcaa7QpRC5wZBid
acJrOYo9FvYoJAJTrOoi24q0x8RBYtFFQJph8PMta6SrKQbq3lmDQHdTO6sSarsz
c4Cu04DdzM36OdJVo5tdgpgMjZ0byogy4ZWCsylkOBvlcx1i4PRXnP7fLlnP1wu0
n95HwNcB/p1sUiJTRFSQ5Mjsu1GJVQ0MOPPHL494EvUkypw13F0oDqVkNxqEgzhY
CSgeGeN2o6XH9Yt2MAbmCzwtolf67MVTipGF5N2T3ATU3j4kA5yykJbGZvU31t27
SRnN49S5Wiz6Aa2ryhZ3jo5RRrqxx8zIbJMFw/rSDZdtsBb68hPMNVGwXI+QhXF4
teKIPh7CcZOwN5mUPzy/QP9E8kkmH1EJOcUfSl7kG+jS2N2Y5uIF5MslTctRYNvr
1Y/wYb8h5g0J56JU+uwNUDfP7qnjYa7UA9i7dfMRgUGL1fWoq7WWsMG/YC69qCkl
uwr2v/4fvu4S2X1Q2m/xJY0UBzfA5NDsDxfRRx2WeBU4mnPqDqFItODuYKMzVr2b
49oGUpaPe8NBmQHjtamRCbLTkOriwb496OFTOghxQMLBsTZrzucSe2aq4ZAxBKMC
SQhbYz3/H+2rFctkZECraeER3NnUT3s19ohx6zPyChxrDZDGauesDgZT356skAaI
pkMivSDsSH6HF5UyNQNnkjwjrvfiFrjkLfC7E+iHKFl6O/IEl7d/6wpfm7roH488
ozFnwJ/tK7gCmyz7jdVrpwISb6c0U4mjx5tYPv2B34MdMv7YJ7Z9LYeYZQne5Oc/
Q5geLzDrg/LLmlNaT7GBMLo+pPYya9JmjE+NyGeAofeGK86tNpinS8002/zSMrHy
kWA4QpUXWlvLZ/3MlJhCOVHmgclIhGH23Cm/XO9xFxwjpqcvIRFmODQoSpzueiJM
uQomMrsVW7TW4PjofV6bJDsb3wbpYJC3D1Imn7kpfzQZZHMRhB7ufxzQNo1rfnjY
q5OJrd5eSkjPo5sw6RStQ5o4zjlqgNgsoxlOgffFXNKvCktNM29nXE84/qTALqUJ
Dv2B9SQaLwSg3gBDvDraUrgUTtzBpfopSK70Sc4SRjjwFCAvt69X/It0/ZI9v41p
oGz6chG1Oy1OiNPaI2lRUe37f5qYwcBZPNo/icZszcU2CeeMFTFWslqzroJz1e9g
aUCtLnyHyQnB8x0hjqLHsezoL2O1EccIXoCSzLF4foeQLI/t+D1R51SbLQS15Yzd
KDOOMLd6KR3lOIPSbxfTC51//gJO+43kiAyZpCJ/6hHW6DHAtGTmkmlwqmv9upZQ
kwnyVI38WZqraecnN0Gzx69SWvaAAb4MtIQr7DjK8GIRuDxs2IlNVnhnlMZEiQsJ
jx6bJuODfbpvJMdyLkzDI0Z6Qjh62YyorKJ2TJmZwv73czRessKWkrVgGwWV5pqX
HDOxllf7+641rYu0CoqvdbiaspUtfUjiScpttY4PTNWOnoYYnfXGxa2p+zjBZhcq
yxSsiL8x7E9eo8ymuWdVQEyMANsiVd++wpRjd+Wn8NIFbBDpvFTv0zpXxKe6IGWO
zHT7O+SZlokrc3wKHMQjgaER0ROeiwj9reZxQJnqxpRyQ9L6QgRTEGZjDJrSf2D2
eHS0k44IKyVklOGCpRCuj+C4lATR6oK0E2zw3A/fNojBcIStw9jnmG4qR8Sdc5p2
A6/dWw5DSbSmbNuoFdxU6YVH5k9XuE6IYviFJzBQ1bVQPXv3nLpdqDaDgAX0kfmD
2OXhv+uWncFKulQ2zlRvmesM1LgMes9Rc0Jo2zWBSGeYWfUnx6g6+WG7MxAsqJUW
DROtUwpmRabcX3f+9vxcFthco8Y+fNOPkrj+zKgR3Bwzkz1FK/6iQSL0qMeAo3F+
2JdYKrSSWUxpNFgDZml2/8pzv/l23GZPXxxsh0wXPWSVmZ5s1ue54Wak6VSfw2m0
tNp3anQxVXqQ5tfXgWWRxfJavu6WuWs2cdhS9/BRaxas1djn5nNvMB8mujmwQ0yE
15ngNXK/Dm1CDP/ChJqzhohfZwq6+0d3smLm3ggisPTi8B76jchQzu9En1ShQfC1
rBEFF6swYUGFUDHTUDbSi4Z0UJ6uKiHbyoCuD0wIwMn84nL6z8kCi0s+7GbVYbz1
JXsyoYthTXPYgCpele/y8LL2HJa5oOYkrvLuAn2LfXANFm8BMfN9LhzEqZg+8Jro
yYdU0HPHG/UCv7RcoiZYHsAQMAN0ossrGSpwUufep5hJwdsjuoak/VtgOwQvOOpt
WeHIs3luDDVygLspjMkkqDKTAyqWz4/3qrRH8T6XnRTwSk07aGtrrqklHq8POND4
/lM+ajuqNLwdYE3v/UT8SFejdiGF44mrwGICOVTyHRmcBSrkAid8yN/FkOfq/UUE
/OPUdZad3kjd9GOF2K47SQOAxgpcMnT4FatQjkmMmYVo+JpnZjzxWUdSReaqOjet
E057Lwod4C68CdCis9BGjdCQscf1SmqfzBqdJ0ryhLQIb8dfjfasuJEZUAuaiboY
QX9XqfqwEcUivABmnOd1oJHCllWPvrkL4KTs+Y+hLUbR7ZteJCGMbkK+/K0OlP6a
vwBz/39uHGvsrSyK3oqs1iaIEqWnnTDjAV9MgFiGyJQ2bcRI4KESxCTkFhLUAz+X
SDRC7yQlXf5r6JMfkhyNUKgIFT8YsH5oYM8QQ9R3tkqDmSsZ5RzZ/46fvXr/1NMW
UnHj9KptBKiiNvEpOXIQbyEfIlRI8vKiQm3pBh2lLXd1mXO3EpJKXfbCUF6bRCT6
/+SxlHvbh5j7pwohDRZoMHcFGPsmxmWSm4F8FFjcX8n1+TAyRWsOJqt1FSriMVmV
ENTrZouAGB4gvo1C/0RkrqenSnPuPaZKlDJY6VoM7cxA7oEAfwo5kwqu1Nnah3d7
MkO1jnUk5CfzL3fvuPBll4flmcxZsjKh2JFrnzRROcUXYaf/o2YpnzzfuYp0dVyU
ymwi5xOc6TXrJ9B4268oPdkFxYzZk7GkYXHEZNXXWr38OAu8Scmx1cdXoeGtGrBZ
o/kxNfzHTXTBd03YSKkTJFhTAhSA0/Ji7f/G1T+2w3R3goertX96/0AOcEyvxsut
MOhh0DGBhTasTnyf99jYe9S6g1RIOQmBUjKaU3GMA9CecAzFS16iL8tRIe3y3/5d
h1BVgRmtOrm9r9LM3DCbzAA71VjlBwRzQ8EeAVrvX3ctxdoL37FT4NVflgDuqsOV
Zr+Ev+PS5A+P038giX4a3h+g/5ntWgfeVI+xbCtf9NUSC9VZoL8hVcNe/Eb55kDS
dBXNsanuOvrWhNVAPE7oLpWKvIXysvv0yzguqHJ3KzAZBt48itWsiudz6jH5YHK4
ebPAH71HZ3sIPJvdEXkkdFD+c/KcVP8/DO86IO387XzR/JWFWS3kGofvJVZNgSo+
PFHCvVbQTYd5+nQWHyc5de6ci6FUijssBo1bCNfmnUsbjJvR5657NOqc6cKg1/Xs
RUI73lIO9BmvOFMj2Ueby76i5HNVdGVw93v/tqLHkBq8h2FatwWwJ9GlANJGLUOl
+vh5sisOdNUGjDuWWmGX7nmQYjCIZLotP3bxJtpUglpCQxpyEIToBb4aIG2P4/72
zvDX49FWhXjAapL+MtQFi/jNpB4QwMlW15IszfulsIs7bVBdf0wVvp+Uf+q2ESn+
JZozW1MotEpYRQWWaqy1WeAHRUOCnbKXZGRadgwVo6t60s2T8KMqBt1/pr0yndR1
ricN4vBdOC91ZSRFt43p+TByzBq6KipeedymMtVcr0dUZjc4s+cGSiCtyqBGhw8a
Xzm0/roIcheKZo2KBtS7WZ4eAErkDuUSpUOf6nuUnWc6G1cWbYpB6Db5E7+1ftAM
hjGGSRRGsnXp9ZleYxR3rVh/+vxDm2LILpQRKNnc/HE4eesfNapFdQRFXmP6WnXS
f7uDVOiFbO6bHG22zKVtqTHaViIk0Qmxb97iqSNG5q/8JaqsyuQ4J9qt1p+csqqG
x9Pee2+hlJo+rdIx9gtgD3E86AvyKwF3VKIzOh30/C/JHfM0u+4t2OCcQ0u1rBRm
rbtYdAvmv6aLXy2AfC5t0YNyYbHvymHPaUb0htRQ8aALsaFDTKrxIpGp25APojEj
QxF28wDrkRlyLbE+Zs/Hd6XD4TR6SAb5nYKTV8VM/jUrCkGCqwl6Vwf9b93j5w1K
t3y8qyIHljrC3zy9nhMDpqBhiGLSeOTrATicDK9F+gLXa6P1G8KleP9dHOlIQchW
okzmEu+QNqgs/C73qN4G7TXIioMCmkv726pSmMxzjxty12vK9bAc+wEmorkvngKE
Cn3MChsQOT7jQdHUqxdFbP79go6BVS1ncHjlRho3C1EoTX5KWeq5XjGBk5jyQPCZ
6CIIjPV3C6tJe9QhZcQEJRIuI7+S0nPpBrV0VWMIhlGlfK+MCIY9zSde07ik5aWO
D/hOgFxHnWd8FaX5OdFnsG8CUcUgNAM4q9Z42WdQTcrjSs6bisRoVwbNaNrC08no
rcpXYAmP1ADPWJOES8WOgRoJvy2i+womfqHZx9PTSEm3VqW2p4RC3jcERSSzfFZJ
DbYt3CLm0aTavjPjx7WhI9ePHX8L//kO5TrtS55KAJUZc1NbtYfx8qygrhOVRNo2
8BFIvrF8BG4TCjLXlBls24fQphvZgEpMyl9LFU717bcHLyJEZpCTf/fFACcM0nFZ
uzFnDlOn6v03ruPMhf9iDFPRe589U7Q9qZDVjYOuIWrmh/ZSVuDJML2v5hSCvFSd
LbPCXE0Hn1tZnz1H33T0edYkO8wpQ7Nk3jZkwj2O4So5BBW4xcAiJVgVTcxs6i0S
rmBI68AHYS9wzbr0XMAGJWKS5tmTJSsDwvadEMsmygY04kiCB0jsTv9c7SBk0AAW
NPqTUOQ/Dr5FealccivUQEXBamxwPBkVP9tiEv9g2Y8fgzpgQKa/UjoinvmmPguz
52k+PlZTKL4+DhESnwxCVPKMu3W+UjPdRR2k+5ElWkYhxOCxNOzgmrp6fyALh4ER
Gk1AI0VAeiKFuIm5mh6H8zoOX24V7UVX4X08zVbeowKHWxxRQ3a42aUrl4F4gWfQ
MyVrLVehzJ9Lxpa7S7iOfTFbxiZptiGcJ7SHbvdPdYNot47zzModpJU0KnIaoIR3
9/PpZr21zDd9CALTWBB2wJcsiB/7Tqod/mm5S1KWZjgCVqlmIZw8dDoOe/NN8bW4
5Go20O4yFMt2mfMO1Vb8/CupQ0UWQx0ErQtiXBg+n0u8cg/6vjBhb2Q5fBkZiySB
xIkbjneddO3cVpfsmDCWi1u3ebzzTpXDcqaXbPlsoLQ3WsL3X76zoySTXCqC6M5C
z7tcOewECD6aFxnECgEKw+V6DNvJERuroM7BZdYJJDKw13UJdbLQVpF0XhtdTO40
CtzRHak0AQxNkjJP0WD+kx4E9W5uHbnBsKCuHYT9SW8z1Je7Wp95lKgGXlCgvsS6
E8ZfzCdQ06d7b10pzT25Jetas00Sn147kmLS4lN4DuFghPIc1pRKMYO7D3db7QK9
xMTXwHq5L2K1bFSU95KGcrdOE28Ho3zMKeS5T/HnEpKRhVTLCPYRVOfrXmuysjtX
2JwQedgBgGQFBnvbyYH8LDHABGIJVftcdVkeezsFu13EJaFWH44/fu1XrrzIfFUR
HHYNyHSkJ/S854WFl75VJ6o/SHB2quW5kPktnq0/QfyC7uhL6KpYaU/YYuI8useE
IgezaXpbc6/9A3OEFbb7UCBPs5FAHc+ZyefBy0xFvhXmg0QoaN3Czdmm7JJiV733
ZK0NklVXVYKNR3FrfhnfFrPX7TuBzohBMlkv/24X7/WWXPotIUJE0LWU4qRpWkFF
LJqmDmSpZsTNpVbSoqvllL7JjEcvbZTnq45NSzKDCmq8DYieci81J8tQDmQCoA5E
30neEtAeIgyKzSOWPmWbPtvD5VEKaARJIu5wcXUde5n+ugJ4DcXOAuImRTZCiM9h
Q7lDMRoo8v2gDl2urQF1ibkKiUYPp02iIsbzOn/IzQtciM2V4VWaxktfPpzLBuLt
4/7RMt7gNX+QLoMHwfGG5jS3YIBrRGlCC1R+PualhSTdrPD7k/0BXeFeTWUIRBXs
HxHd202XckBcV7/BU2999LrB60IwTPM5qPJmrAWFEztwD0m8E0cWXCFkOvvVpWJF
8g0/Tqu48DcbmhVk17sykHtSqwzkuv00d/VPkyM892s9Tsk3vxdsSJcD+LJfPnN4
NgsTmEKSS11zbqkFdqgWeQDBisU9Ck5ukTmqCglZGtgMBEfYlcXUqCiGmWQf88ej
BIT0ylfHya90Ht3biD3TOsdzcj+uTOevES360/MrBIB+/S3Y74bZN/w0ehZQF9rA
iViTJ+CDZxjKjvWlABFXb2AWcnPekuN3gsdMmUovYa3cI1S6gZYewHDRnLVrekYU
U52EuPgxmXgrXOKeIF+DWykAiMj4THQyrPoRyndL2GZOxDiSghpWz75ukbbevJcm
Dv3WoG0jXZw/j4uhng/GFHnjYX9j9s2VXf14KBJbgCtRSsJ064hDrukmV/Jsuu0M
VV4uOTlMn1nvXZhBkq6wY7wobX3MDjRCLf2AAYp6tsPdSEQDkmvOo9qrDvNo5KNx
4NWujzjrm19Cf1Te8ifqItcd5kehKqskEBKDG+afOmArXcFmiHBI3lNwjbuRYu4u
iCWWT5bRkSZGb4rgJaWViObAwY6KlfyfvvFtu6aCFpW6YbhpzyjSdL/CUsVmkBJ8
`pragma protect end_protected
