// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:22 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JUwt78uYXs5y3ub+EOIUxLt1ndC9yzxghFlaNlMKufJ81gVcUEAsSRLmMtBJfUip
ozmwA13d2DtMnuyV8vkYRRRYYz8+9wiEleiVAmOMEA4qzWwU14OLC41LwSXTUTOA
UiyDvmnn3Nw8oScIJ6RE1JK70pFgdckyXCVm60uzlXQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2836880)
NyxpagWFb+AQA8quDR0ax2uYUvEArHqEdYrfCrM28uYN4DaJDhmObvHIG7kJ0kFB
RqqcjKH1um5PsGXPIi/strq4CJM0piLyEaCnePCxBg63FEkFz1qqCKgk5h8Dabp2
56u0z19YW+P1hMlbnKST1tgDVmj7ikzUXVndHhI6HUHJJqPc4cEQ5y4h3h2xYfus
xAD4PDpZLBztKqPA1tyUrUPqeikUJU/X77WWSp+C5OlYTG6e3ACJNytZshMmQMpo
35KzacxjiPURWbLFL5nReL1e26lkxugZn95Cyw1wrGskOEF1XWf4x6vvFaL4uM87
fFjtzOZdEXA4oEEFljobgTnPSD03hUqHEx8QviSHzZzG4Hz9IbOh9N0lqMAuEB+S
TAa5FZms6qBIjDCVrQXkKFnR7/WL9rlOud0w4EOHKWMWvmh8ZJdSFrR/ktQQskf8
SbAZ00jCQlTAw3wNsG7vG8/7B4mruN372fLPqkYOGPJYj19OsjuQcV+oj87f3AEF
mw3c7eSaoneG5Bit1GCziJ6RaQ+d+wyg7N+U+ugVrISdFFCLCbqfaVMIX888s54x
TudV1ZNAxeR/sHMGLFP/u6uRgp7pyio346biz+KuKIsY7QvMYtzWuLUn0wSx9RJg
cVSQ3qDLBNMuESIWJ4jeL5B6I5BPIw2UPPOi8j71paSaVA5tI0b/54AkrO6ny3Iz
k60zQwGPr1Y0CW+/lwmGdU7QbJgelkdgxSqbZoMxHgIdH7xl/7h7+Y2QMd3PMlvs
u+Lozm3Uc780fYN/lahAP3nDw+t4mF5xJKALs4zqUOQRSd5o6Kx8JZ9DLZxntOpR
0zTEESO/aNtxOcnyld667B3Urh66yQborDQYiPaof0fhxEXhwdrLAwlZ/ONIBeSf
FzQOtVyZMXEFinWkR3cg+lP2PKGfjPJV16qT00UGIwvt4mS82GPtvtwfa0YL8LTG
tDbjF+Uoy5uYsgVfFjKgRBN9Yj2F6+OkMrqZCk1h38d+Yi6u6XrSdUjXPP8xptuX
b1lucF4asJ7kKQOfM6XQWtofmktPEjJJLzi5u8v7Eq692t9Q62J7ddVTMnopPbMN
IUFWd3LeTPUCcIggRZqnLWFj8koMHwaDpw4WXDwFtFt6vZ/6zEI86JERYFGfVjXA
fA6EUd8gobzR4+x7AzGv2oMAq3GZTysUnmuuMUIAxBczfK37/dKg4UkMaSNukkKw
pQPm65bQ3O5DRAJtuLKLwgakpk4pFdzx7Lf3dzZc/T23q9HcIEcVKOlN9Xm8kJuB
0kIzrQG/p0Ac3OONficTTxFUie+vnLX1GH97ePQTYZYvRoLK/pKWzGEy02msXjK0
gFJeX3lCuJwMeheWTxE8mIEwL6BCH1ukCR/HOlOi2fCcRMTneXSqOE4s39M6Lte+
FjRopY7vq2vPGmiVJzv4ALzDunDRY3aPuCvWdrugkBXWFbAxsLk8sgHJqGWVS5rQ
ux8VoKU5tmkcVrL5Wve8jIq4MqyY4I5/dO6ikeo/jJexkzGvZVejPWvlyEZaqn6+
QRzLS+XxKsQAORgXXchRJMnV3K1oNXADik7XxGxhw81Bwz9qBWeePL+HLWWa9180
eNRkKvqQyk/+0iL4QUbP+QHZJn/gdYZR6jna9QWeOBTqsLbo4Lwl/zekuLYt1JbW
a44NowEe7ZL7wl5y70w84yq3fcth2+g/KissSrypxWXqIcjszQxI3Rb0RlCp1LS3
MM17c6ki2pSevtOmj9VyxAZxof17Q1Jm8AsjwUoBf0ZyNCkq1xXA1J+LytUl8buf
MDSOHusqKlX1fAjlvjBGZuLzu6xATrA3ZzwGrj7MJgr7S4Npe8hj66ssloCLpnAM
8bd/9RbmzFQT01MNxoLk5DMkJuhkRDgOm1K5sCm79cJbjZMAkA7F3lbTYFEY439P
j9htKb7MjIhn6kqfG+SRPDBcCZANiXotv6U0mYNbOmAaY99DNCh1KvsN7MaxxWpN
ZKduIOjVXVnQsJfnDM9i7Ovym6lpe2GhYL6oJk0gY79WkKGG5KinKNj3DmBKXsrD
WhLd1NpSYhX5tGKdndJfKg4yRvmVrzRxcNNEdu703KnSHcY4gTRvqxjCKvf72ieE
6/bOm+GflhrIxIgWI5OqzBa/Js61I9x+uSbxefdW3v3FQOT5kN22zRR995lEzRJN
lTJLCaLM5Y/JgKY2zmsAE3sI4Pz7bnGIfEgnVlq96Xbduuuh0vFfTAlQKu930RO1
C0aN4jAfKiXubYJXYdjzc8rHJ8c0sDDmkH7huPLXwdCxdtIdK7lxEpUmG1XW5VlG
UCqzQoOk99WDoIYDXxH+T1VuZCw4HUNl7fKiAy5ZjyaRsTu4Y/ID0iOHLC6Gwj45
vwmuVaaaDfJx/SJ3eySjJDnCFZUx7dsJ+EU5qfVBdGRCJKxVEd362pJUEiYWCGk+
JAtrvJm00VA+Nd6m6oB7u95cNNf91eybxybMMOa+bJbe/CiH3c5iAIgVgjXhFebn
Rqwr+wGg20L47rWysTOKeAkRTtV7z7N/ttCsLw8eFkhfv/HLWPjbTBx6KS3jwcKP
LJZTh3hfyOORkRxchXirUAWoGYrBXL08Bci+gBvWWffdiIJC4FU3tNr3Y7KOpytQ
x4yHzNQr34tcmwgt6m8EXqPoEbXUllSfLZ8TKF//URvZlHWhMQ5mLx9lrz/Zs8vs
tZrWcNu52O4qqfYtfFVb1ZCHccoOu3ffK2RAk7br0pdhlV8OgCePIUxYGoTYszLV
w+ld6asem2j7JBhIALjKu3HCMXQNCbqlTD9T4unG1IEkLibhjWRD8AILanfdQ/Pk
HiOQMsvsnuULjfoqd87PCPWah08RsKk9yHTs2KYttGNtMgKXxgdSsuBAGX+dl3Sg
OyFFlxpBrCBebajlNCZgxTn1u9kValXaZ2uXPVgO9pxppgTXgVRaZkf0ZOZFT40D
Q42QeuQKL1mHES478RDXTbQtqFpfmuq1TbjCSN7MIN2k9KgwYUiH0JJvzhdNboPD
ocIrjqZObX+K+AJZJzQaVdpOb8rnU6n7rWlNwKCYJqpO3x0wW+g+ynIPuEMmqlxx
s+ih23z1bsI8MZzFvZOPFBBwkyNQLnVDZPVBI3kT8iL8Pp1Hqtz6Fdi83YIZLQ4q
IzKWa/dX0V3KaJF+jBRGYrcznnICY0AU6sQjAcxcfCrE3uMKvloNKkCByuUPqpR/
Rhn1wIBYlhd9oDiFtKGSgpKCGyb26DERCxArTVMczik03c4fh2f9wwa3p7acZ29O
8W6bpQnf+m2xqhumhTGdp4h52Ou7hQlJfPmy62w8OhlhmVkGU3aaB+0UrwDKGmmK
lin0Vn/EihBsw02IZvg0tzfKt14Q9kZhDEhBsdCmqeN949TqS0TM9WjGZx8SQJ+/
N5TbmI/RsqPWTssuRNk8ME8GjDN3bebfc6GRn79Fi4eCqEbU/yFI471sH+FPk8kc
S+vIW/8RvtDzBCDCnfe1qUGKVKat1AYgd/X9sSdNXTBhyLPszjOExrIwM89wrtfD
gNnaa8h0F1VVCeR/JYL9XMLkVr2lTgSyxVBvrfebN0+P7Be74kMojA3QWrKCmYY6
+6FP+55LUBPQmKfUPZD7/iTQKaXbvgS3//YThjG/aqZAiHRaRCLNTKRZgLDFPTFJ
Y1kAa9q6YRsgg/AHqeyNI3WuqQYb3BBzPgqs5j4hDDXjbxKdOFeAkALlFPjUcnQE
bwTs9ULgLSPAHIcpDl9kLzdIZ/fi0fTXhl8UoxE8OmpC9wxjXku+dzl2NYu1+JiQ
NCHwzVyzRT5iYCi6LoTojnf9UONjg72yYLUaiyMhrspU3JgHfr1PJDfTgjVJAQRt
ogDrqnpqLw2oLnaEJdVH1zgJpqvyAQesl2ItsVQZyboyLvyfPx00odXWVUFigqDC
qPpbkcfrI/9/+MYTWePq/ni0AXTxf/sOZZVBKiP0tAdJUNBYF2+4TIl/fEH5eXOb
Q8Z1qs9tBqVTeR9sfDVVDwydwOV3L+I/wcT3uA2ej4ZDwVxfjS6sFT7FTclwpbyO
oZSEn6VeyqWNNx+c8SzqsZDoR/iGj3tMvf4fF69kfgX1TwrNqbcsDi6qbQLwrHQs
HcGiRu4zbL5PJC+WmqmE8t8FBT1IS/bkBdPtPGXMEfiWwIJCY9e0EGuTOJuZ1Qqv
baggV3RpZTGilJwV5fpyWahCtfGjEWP23G3YHrZnUAjPUMeiLnFSTBJepFMwozgB
GHxqa0BDfTdSyWroZ+Tua4dInJgSJJC36O+aTT0GHpsaE6dGzmy0lc4ZHgt336HY
lpIv/LUsrpFjVx24RX0/QG1wtVevCU49V3XKlKAtWEzz3o+OvNLX5v7qPJPJdxeq
tXZaTDyOizkkWglNFdgZ2AFKoxOXQnrJAinYUeCObR3R2FW/kUuawcEVUVlVCtxO
/5/WHBS32mNJ1qLMOpJUQ1R9yf9r/p48jLGalXp6dzXaLceJPv5dl0q6jL3LC0Qc
o0ZnA5J9BNAD2ZfDXr5qLxdTtaN6WTy9CeorhE6cQTRsnJ3/f3GuvZOpDOfk1EU5
3d7j1n4xRauXwocRik2H9sdevdsQt8MeDioxJMvlX88MPxNXXpYpvLiaCqE683sl
GhbT+wG6lGEx1j8sdFI+FRecOQdqwFqgkWbxwBtK3pe2gcCXB0OkeztebVk+3IAb
ILLvxRU9NEq4UTyAz+CRLu5U9ZRmS5fZbK7Fnafo0ur4NapZy8VPXWs9inNZXYN8
J1+tcvLrYbq4RtbbF/0tn5OGP9crn8aWw2xfnE6gmUXHc7l4VlIvQhL/HMAb0phf
upErD/6MAfey3Pvw0YruO5WBgRlF0I1w76gHpi5UvVEwf9v6+4jbDDE1tPg9m82/
PadNSAGiW9FyZimDPJXjkl9rVcjLg57Hgpc9TqgO1A2JScKZsf4Yzkv+GuDMoZ6y
mEknqUUbLz1n2FlRM9rSfiFodZU5JiYWf5QckdfzIF3OoLVJLBqiGh+SgYReZd+U
AG8ZyBKq7EyTDy35l3BAQq/9ndd84z6dv/83IRJ0xSldAsxYzT2hsiVsxOqmoL/G
z7AJB+HOq0DPwWuxmDFAkVySVSIXTH8pTf0DeLzhqB7JjVF3R2imyMmGZ7V2gAZ6
lUNepKdPrGYFVeD356GbuxCWLGXzJj+nbaxLYqsi4qg/8Kn78W1lNdgPDQsAP2g2
lVk0UW5fIagQZu/mE+fT9h6HnavJNjzYzQHd9tDjm6Fd5zkyEY2WIsSa1EhAiLPs
qR4u4oNsdIblygNVAQxckXe/wS0C5dhI7ES3/+9yYXj4eQnJV3J28x4K76iKBUn3
AitE/WtPMRMZO2mjIJiYYrCGqZjzYxb6zCDh94XzfE8N50NMqD1SAiJ5mPKYGHi4
JUhGjDV5axDG6MbDsERWOtx+RvCT5cJ2bBGKESGbC4a4VvmfrHacj2mIPKRvWcZZ
XSdsLYI7O4Cxu9B4lMtGlHOxAjE0q00qEn1p4wPJu2O+eDcCgyqJoSnRDasTM/NG
NbElqUCJoWnwc/8goHqWIaM/e9KRUWbr7zMlv84bypAB+7Na/Gp3bdoH7nInH/WJ
FcKWqTFhWD5eT+vV4bQoFuV9Z/7nyx4SW21105V432iQU7ZsZ5uuqwFEHV9MQfb/
oDy6l55Pri16tJHBSaTjtU13iOfCBBCawDMQpaJj6Df47CvLVChDMh1vMtKvOjMJ
L8Hg3+h/ZaPIFhOVE/1YscqwtmFWBjd6tljjhvbcOLF+KpwGKCrdVsen5hghdxP+
RRZ+oAmQhMzXavqHLHe9P+G49YuVmWhyPy0CvO70oqczCSvH9CkoCcCPva061UOf
Ied2lYGjM4tCeEv4xyqjy2ReF5rW6/jyJcWpuFdybn39UYnrxWqG3D326B5PP//2
wUWFjXxphzrsa9yrLgp+4SLXWcNH0vq5/n87z/qEm741Tqg6rHNlmCmJhwlr4lza
RgxbQyH4uTUYZHTzuQv6BFzgQVToA/FBp4YG2Eo7gsDuX60Ql+tDr5E4Z01iw5ED
VkrX8vLFYhp9j23UY1YZGd4roby2nrNnazc0xSmHEOSTXhlhPXU+eSnCgcdhVEFb
P4CGTcu04RFF/NgsqRv9CCsW9W+xPBGvSyzm4Eof6+sFKGmZ0n4PNBPXiTY+e6IV
yMZ8K0pgOKnhCmIwDbTnDhY2RQg+C3V9s/d/zOJ6dn10kk24Gi+WxKlEbSpeXc0Y
UVLaACdUHG5/rTZpsixr5378rrqnYVG6Pcy7DRxW4ndrhyGXDYB8jn/Zdfhk3l+q
QGr6MRsJGFJD7ec5/kVoMj5wsb9rwDU/acgBspbYz1mcLkGgNBaZWwR7EnoCKxr1
JQCN8qaGRQ8QXfyzfovgTqny7ysEYbg+bMQ2osAj7zZXUYl6zLhNWAA3apbMzKaB
060qXwRYaNtefVoSAgtWbQ60NmQjOqp9FKuzPcpdEu7WcY4RXL+v5yIBYjArpsoE
qz4r4jD5sxr9o3JKN7A7m4BA4e8Pn20lJ8wwhbhzlFkUZzzOciKK6IBkXC3RjrCo
n6+OzX7k4s0hVedSuyQXxbULeOabuBMiaopJ8LxycdL6EiDMeA/100fCJswglrJz
msK2b1FB3ADQj8S4wI2pS6EsdCIsvlCOqtIxCjVh6tjz6Wa4f+AJSywfXnSuEtoY
uuBxfONUm8C/okfQcIZ6vn6gyQYUcsTpPQ4PpKDQs4wUqxuVZyvKOoPHsNoOCIfN
E/B2iIXqm5ntp0bu/B4Uh2Sqzz+TL02D/DJo3PeUUMjuhNFG0WqnQoopavlSQF74
IxGvOoxyKyUvfK2AFe7g9Re0iGj7//eFoHyV+Sq7S2Z5B1Vo6W+lpGEvvtVUD1fv
PlTQtogwxwKHQF81wm5fzlqlboyVh15OQV4k47rQx3EYD6yWRdsEgFslhhiD3dd7
WUmojgY+OpW7joUxM6PEIHDNq3KzXDQ7l5x94RlEdqYA9XUA3lrzzuzRubEl2bKs
lYErGuoP1RsZRYc2y9vWrBO7JP4mFHBCSoiKb0lPQz6rgJbKr5u/1Qbx6MormwtM
iuuYaX5H06306HgZJd0hdcwDAF8WkhXW9QuUJNLQewOXRWujqy5Ie1s0gA3PK+/6
GEyYibKxryymY+qbD1mMET7PvwWLiej8Pgih91wmGSJHL+6Pd69aEJQFCTOturE+
EUx+bLWqr7I52t/dvzVEWTRYKn7j+EFsNSwy9QBYE0nrewAnZvRzxURSUj69ZYU/
vkqEvHlIa10Tp9OfcDJC7pg2vBgnh4XqGMHhXnDjOBRmtqTOYLCnMOF0ffbMw8Du
UpBGQTLOLhBqWX2qePotR3NhH4wIuz8aHfRmpwNO2BdYUSdmtMyDCOtGBrZ2IhzE
DnP2Fy5ilXEV1egyw856hHJMmgU3P76Zz1cgtPKlp3nEWAvo28UYQT276+Gl64Bd
ejlxDho7FVF0DyRhx6YcCdZReyvC+BfKA0LFuuF2pkTlDAIC/QFXtHap/NL9mL2B
vO6LjU/KEYRlZc4pZK32l17i7jb1RMbvQwbMqjjoyNkLLzFRaq1TE/pvfy1eBXE5
IhuB3JQVEZ4MmDtdYiK3gIjxj4oWgIDYhgjNPAvKzGhRxx0TKmzU7X4rRutmNlSL
AgEime7v6mdzaUfyGWJZecIR7gJkG2/Y1Fz6PyAgxAopa+xL9NYPRAwBGdaWzODg
18YA6M54d6x7Wr6hC5yQerZsuOJZIy6NH7awDpoHhS0vrAaXFrP2k+0LlrDbhU1C
oVLgzYO9cYLIG07X2yMnbdJx2kJeYwQT92CyZP2ZvQQmd/bkDyCYhANmFXNvZ+lb
tiPtKO7YZcgAHmN9KiIa05msakbXaS9/p5bLVIQZQ8OgTNPvKzDAhiShxd5fNup0
DRl3L0hYmBfXRPnLB5tTb2rj4lC54PaeHWKnkR7VrGipmEfdpfEQko0OkZ39LwJy
WlD2T4MkVwDp82KiIohIU23lpp1WFZxsAeVoB+7SL2a7tB08MWUC4uWUVCGB+lmi
XoEa/x8bi77BCUlLQXXLdirQo/KvtBmDFqxztybyDpNhcwlJ8sFCt+kxQRlpblpm
PaODFRaClAaUes1yNe0oYMbDV4G9BhmCUFUiX1JKe8EIm5CX9LVpfGNvci+pTaFv
MMnQQjzpMYy3R9W9bEmNjUX84YnLYVTgUSD2uKAoy8omcMwqrLRYlKYgRHP5WU0l
ry9hW03NgRL+oXZj1i1azoUe2qlnrvXGyrNSjqbs42vKs6IveoTo0bKaMHbs0BA4
+oPgS3oBNIdNgaZtUadtJxL88EwI9mUAgc6DC5+Ko4SU4tI0oNIa8iNlMwQ9c86P
1MqG29T7in3REC2Cq2uRuJRzP2l0cp1cu1+0ASlLLzhWLH+wZcph2oNl+bTaofoW
gB0kZaUZDV5MqUd4C5B3fAgWvcxlF0wHUrQicdbIewqRsSJxkUyvs86ZA89fGlfZ
2edAcTcoNofOFzaZmYuI6As41Q3BV+ZWhiu1vsy5GV54Bpvq5Y2dGM/I8KgPIRgD
7CNYPFOPpxR4qcKAja9ixuf1PN68mHdurS6/lvdB4i8ULME6MSe1I/3BfLJ2Wudm
7ZiN37pv0JNmmbRGWkyb/mJwgiOUyzOxe7QVdHKhKo9TgPTi1npFy0v25gWC1AxV
Ug4ROP4gUaU4GpPvHvrwhuJ+MYplXrXpoy1Y6gJMe3qDcP5c8V0QogiB3n4GOGq2
a76Qaz7P/f+Vy9vjKn+W09KonS+QwsJW5Su3plhpWYeXVPIYVaRiYLlnGCnMk5N1
iVquXz5U4EA58azDJgXWiCYGkqtSYZpmiB6HpNm3KHQc8gD5/Xp7x9boVAhNkRL4
FRnOs8uorGoGUsC+qw1ZjwTlr4XI+uk2trsED4dMcktgUWqnqA9AkKdMLH5tWK5T
CFpnLvF129qre9YRSi58MZIsifhO6y0GKu0C32JQ06du5IHt/Uxch7I0ekb0ezQp
G32xvEAJ358k5LMbhmpcDye6qyqn2cF5uXnhreWIdJr4Er5jgyej/9aATaQmgdCk
gFjENNLhf0e9JsG754fMyZTNS7r64Q2lkxdBUi6YdBXAb0tNHryRvSaPM1lJMPsd
PyspGgmdRy3zbE2ZcmH2FyPIuheoivCx17VdAnZlGyDKmD7Z41fuwFg80lwKPMco
ErDs3vtGCATwg4IvH91IzpuZ5dtaG0w4MC8sgBP9GWfNT5Mr0eJPYrc/5KDVjQFW
JhmGQgurduj/FS1RqkoRkpfjIBGtKfyn1mRmu8Jzw1YOqOFU2WzoDFrwU3eTWEU/
RiQ9NkKC3jii6/JdygHpI2WHGJzMHAeVCJTn1dmh6hjUZxtUyAdfFGjkJ39cpVYB
BU6jaiMO+ZuCcaS7YhdTtbjG8x2327yOeBGnK4g20fgXd8Mk6LjtDWLMFtPHZESk
wUT+LsDhHJsS4Elu4ou0nbaVxmrQVmkEB+pebxL8yhAH1dVY9qkyQ6RXzoxpE34z
v47uaz3zTGzcH23sluJ2I/uEw/RMLLrR1Hq/xVGhAZrOf47pqmeJZAEW1n7BWzrh
n3iHkJhYIrf76NyPcmn+vjP81uhJHSA/6pXiFLjOcF+XdvF59XcDEBaciVuJ7rYF
Rrot8ydbBSLSXw4xasCNJGYfFemg3r/4A6lXw96o0qmeeih9cEkZhM+Qcy8VEfGN
h2xXWAS/Y0NiOAGT3UxQDQIXc2Lip5rKsh9nh9kyftiA/ATCU3QWazHbYvKo3E+/
mP+OL3GX90L1FgiooXdIUeJOmPmaY0aX3bZLsOYMdBMkbSckasG8NDycJcuPkD4l
E+MwtDVI+j5gnwwvj5HynCDNozFg2FR7jEqZclDEKMKHGMWVDApPHqNBR+9hVk5C
emeT2E4+S/jqxZIaylYCce/kzlZXazHmEuN/GMyy2D8uNL1OkoJYrpuybS2JKUPi
ykTAJ/K78nGCI5NfkvYYgOThsmtl3SM/n9XPjQTQHR4Ff+qcZhsFcwiMa+i/jeKa
2vom3qC9ObN0M4orn9h9GrNZuN0W6r9XaYA4GPvvr45yhTixCVApe6MrOBMBX5uo
lEWBEReBatERUtM7r7/fxlXMLl0Z56wkAcIUkl1fjD+D4iap9IIGry6w+/BrIlS3
+9vFPDMueOJdgjk4dliMGs4Ldb1vGpadTaPCdxc6jyyNXPauijUnutpuslcoe6rI
9REZ4EI3bmeUzk2p9NZqdb2fKgjaUptQrsSsZ8dgFbIUmDub4slTJBwPUMx0L1pj
DVPPSOuLHxXSosGzxurUW3xNIUrvyZKlIco3cqscc6CQ7Z4qrgHhsWxgk0XooO2E
bGWwPdxjsNx8XNMZOL7K7aLFhVGRJ7VxOIVieNVPsGN+3nyM5pV/eQexzjThNw31
FhWqzrn9jjOM6mS0E7Es4lOfLODwuUoW1+EVKgK7ISkRjDxsouDyVyIDvp7boARk
HCNgTReFwXptVckvFZbWSz5H1mHOiKYf6sjfExhe2TM+Umup+h75MWrCfhj+Mjb9
je/pgkCddC//W3l0SXt/rNNp5ux+U8Ave3AJmPck3UAKXO4UXyStebS6PgEnEw0/
cjzyZNJi3uqS9qt9wa0FyhTYtboOM8WXOv3lpr4HPf6yLErDe9sZFfFZeHhUofnU
lBz5qX3NbnCATrUhd3HS5NZXhT9DTkOX9M9W9ttkAO4RccCXGjzkIbR4KQ7DddpI
fUNDKFcSabZEYTbvBKxo3omeENjccKUsLkV8eQrhO9XFuJNrgps94heXpS+XRkYG
8lOh2D52ENKh5nXu6rpTMhQ9fS3QE3ZrqlsNcSvbsFiMgkjxgpE09KAzfYj6AlLA
fPLsHyFx3YD2YlilsSyDCsvlGQ+T1ocM8+qUjpq6cKUT0wdN7kiPvW7mha9c7/jA
RKeHr3nTEhNnAh7hjKhBX7yJvWmNot8pQee6lbyB3gZmb/EY8MAwEsg6FSqCtrx4
p59zJFjHLqWv9Iiqt6l1j7yba2KH1P71SOwdPQ+aB1V/HOmL391HZ//n5AdAsSCs
ajRUy8lK3ZQl09pea1AL5KTMlfAxwIo0253p49vEVU3Y7DhE/mUiZuKCQ0Ff1P2V
/4g5sCyNNn99aW2i8wSfMkMrj6p6V9CKQTUeEwhBcNuZuCo8U7DQ4Uv5gciu9KN7
0KwYVBDnWKFrjwxq+x7vnPMtAl6P8lv7V8prlJPbXUMd/l/jh40JffIkZGbOw2IT
O6RJqkNlizVt/1634fRSE0NHGlITzmR7WPHrAHd/I7adysawy/8WZeZDowrLRh3n
sFgy6if2/MLxoMRvP8B0KZhQz+565RIpTsIs698FTVKvpvQBknHF97KtL8wMVoSq
ZtOWoJlq/NAOhJjwZ1SnNFLe/9iSF5U0vSLTPM8LF2iGFHWPBYHfbhFe5l32oA+d
tARzFItCgIamc0qJO3/5hZxvyTm/RJ5LwjhgPkyNAEvNT0DMesIdAxq1gjlKD5wN
QEPKJHWJc8l0AjUfaecpzHsN115SOBWDJVYlHuAfVvM4O06dBomnDGAOrpl59ijK
aDmBBwbQOqIighOsHUWRsLjrQtUVfUp086rIyGsRxuqDqCRM6cAFysWOcmiIDsb8
k2pZ0VvNgyt9/+oTgR1bLY2F4AXXK8/3sCAJh8FXWlRYHTxJJ7c0ra1dyZ4r2p5E
RC9Pdyu/pn+hNO6MSOcPe6kT4xqlB9bufUq+HG6wzXWz2ohYcLbQ/q55etUjnj5H
av3mzB0a0fS3RDbsk7lY5rcTL07jNn/gy8SN0W9sPIb28kf5QE2DGheLk26dp/aU
MaBUfU7se77pCi6mnuk7zvWyqQDR3llhxMV9Q9sHw4QLifHzytWpyuhiBEPJS+Oc
EoZXo4TDuwKlMvvLDWRZdQYC2813lGAafucXqj+mC4sqB7NBkuQIAs50UsYoVoTq
E4YkuaY7E+M0KB68nFqYjeOLuTucZF3iR8w00dP5rIAUDphNguumtpr3RHo4hzWF
kSV2jjRlaoNmWFytuOpsi77Q0P35QbWsTfPkjnc1e0IAm1BBQgfsnOrUoVioK9kq
6wma/NEoCm0cn4ejilRCDbmj/MCnXqBDY477CX1T5MwUti8FtA1Ou5MdQ7A3f9t9
HbYFhQXNNHuybim0O0iB4bwAppdki2G1m8w1J+MWWHq57j/VeD/thsIFEdDMDtuQ
3iktnsW9hcmine/VvNSoRXs318ZBGHK25CVPEYNAoUQydJKZkSSy/GD2oWvnTKes
rG0N1NfgGkAPKmU9ovyNjr6osUradzXCusMAeym/htt1S3llFKm20XTfT5OkePCF
456kJoK/fYMxiwEMUnyz4rqEIWAamFIwQ4WHuh6MxsC5v4YFfLEiejBgwwhl6xok
don8TL5yNHvHEIg97zkjkUAuXmRhF63VhiFmVm2WXpZqSw7dx/J0caoi+qpDSJVe
lGs4fyzsXZjhs0X2fKKgLaub9JPCVWffq5mGTY3H55/7lTVyj+ic8klo14Y6BtTZ
I5HRoCS4g3dBMYKdiavDncC0N46Jo0zGqRBHg8DiFrO5reNlbkb+UHTGmUZav3pl
PKV218sv1V7wxsnbEZGPOTBf8jx95SnDTl89nB10CmoU6+13JsSxAFB/XQRYd2dM
jL4EqynqZmU2S/VqjPGbBev34ZtZLpOe/SeNs/8HIzvLWiv1Efa2mZVEGJjAqpCA
BYmnem46mMY1lBVvrbh01nCm7YyUdYN7tVthrDk676t9U+uyAKzNmqSZyJQ+30dn
iiP6Hs0LDOIXJ6oR0ls2MCqExcby3UfBq6hBRyn0YjU9x+rrzOzju++HljWmXSzs
AyFh5Ezh2K8eHeJMBIVtmMFMFdBY2mV+UUfMMUKhrn8on8hyhRujF/hvUlcwv85V
c9Y0a4uByhlpzb9Slz0RjmR8ew07Vjr02NGXWc/1VnrqXMMGRritnwiT2UmtTsbC
c8/I1tYVjj/u6p2PYJgqzbTPxYnuRYPFw9ceiA7gKzNhe43xCOE1u9A7cBPMD0mR
WQk1IME4hRoifd49jQ9Mi8A16TxWxkSfEkmOVxEgGqOpElr3thyynbvrCqSGreLl
PVSxI3YmKB2W19oL9TxVa6RUn8F9UAy9gZKudSVZBA5l9iCq3mfNSsYiKONT6Jea
sTJLqPRD6gaBLfLrcKScyRC6FLYj4wNqeaJPw3Yr2ik5LUdkExwXWJ4qJcqe1JeW
TyjAc9M+BqOCYH+Gyn5e3hN6besrdhN3DAM9iOWGWyZjOTW/OemM5tAYqnJwXB/U
X5on4yYuoMW/6fV2YskKE8CxrpOdCuDxVXL9aIPjeMOSFQPKCo5M23Sb6jBmz9rM
qYmsrrRG/VXmW6W9sD8jGSbpPEO2h25XTjg12/eb84C3iJSeF6eZzCsB1DHdU4ee
NiNFZTmDKULFSLD0C44SDXbuVcIfmoRAq6qjDLecqp6ncpSs9TNrxvNj2nF6Y5eI
u0jQFvnNlwE0jF9XIULXLR+NMS5Co3IoakQ5+beBoOvidCPlihtR5M5lHzy6qg/N
BEgfvrRbL+ZZLzbOM+LxQtAMlOmAurdEZ1ENWKF26kDtI3kGzUAQexOQuOjD+eMN
O5P4EbHt3SgYMhHMTGrnAbNiRSB7aCAVLLhwomSxMh7+D8O99dRNeISGpmuCoGo7
9d0pDlt+3+3/8iU0iEZ4OfrMN4dIXUDDnHfhfxKgBOv+ADiW2ymX8i84t8aKGL7+
kYaGnZop++BXw5Yqs0zoSbt6rY28C7Ik3pG+ssX7GQTrQBqIyGVya34xpunwpC9P
e6kVi+cMlGcAIW8uveLMMwqPqoqRa/cPuSwpH4QLqkMqGwn+scPt/JdXGZtOgbGD
v1BK7+eoEj3qCDe9tM+qiuW/bt2vlOTjEyx7rw/62UvKnE5ALvwr8oXrs0wQeYId
axWTVZxsNWl+xlkflvVgiHj+Z1zRRXcNCSgARqd/HdRHv0vpd/mYtzlMZb4UN+KK
j3J5CM7CBYAdj90iUiVGNxma4XdwsYQxl2A6HVGLWcBU3sOQuo02RVwKL9A7YQxZ
VqsW7UjCxzmwKJzggbHE2CMBkZTl5VJz9gTAfR02OX7CXPNgq+JwzEu/xGscqQ31
xCTx/Vy8QUNITi2ogWV3bvPuHESrN8Zoqavw3AALwnAt+ccnmR6BK+Yr2QN9m8SF
t7kJU831Fcxd+niqsgZvBceeoJrLtShmJJ16boa8oG5p7Lh1AhA3+GCoKhOyGZBt
TnOPoWu8at77PXWamKSrNkdy0QMwF5QwH1fRel95DvSMwZePP9Ibii/WBJFs4bLN
rpzE41gzBr7YeH6qbKNnD9L13kcUg9xdLCLUClNPBZfHrE/QlaYHdON6Frb27N2+
zNwQDq4d+AIajpkJ+jOwP6OS8M2/9J8TJ2yBi13uewpB55lWw16ualdqer9MqDDL
rCq1C0Z4qBoq6VbbYW6CwQtal/YliCs73ZuQ5J8tyKilx+/1X0R/tVhvWqNW4CB3
bdR84QgCf6tbOf+FCcLnAKvbJp5yPd/zx6yXYYQHpdO7F69LNxCuhGBRiNxw8S1F
SLweF5nqBTWsFF1ImslpM+pOjsN0hJzlbUTuSq97s/IJOEARGQQo/ZNaa2duiA0n
qT5IZ4wlAvFWOeMDmLE9D4P+NgX5S4CbAKkuNm09Ts0NG1x7G9AP2F73LZ0Mdm8R
ao4YgxjT3MD99HIaVSReFlTMJdgpELrQFFmVW5k8yOPeWrA6X+O6vlyIfDIZZKsp
MpvCaY7I5V2gwH1+5kvbr5qBuQp35A8FEe8ZsKkNT2GUZ0K4J0BLFH5klRuvtXKm
nsRnzBorGu2ej2eUq9dDE3dhgamA1y7TT3QOQjA4LONrMqAA7SNZF7Ow59zvxWNs
gZByi/CM5YjCUwOr39IReupcxoRAfpnVvqwU0pInuDiP1xK0LXHG5SwckqEbXOPb
qwMhTD0pH64q5Kkqs+iLc8PFWG7YzaHsnmlYeWoPITMpVbgklZt7axj671zwblax
Dia6otF3I/s0qGl6YGxYIkTPdUOnf20pRQ3NCcxBHQVBfxjOnI3TvIcMFIzpDcqe
+ALYEqUyEv7WfqrNEgSocVMiOEqLFW7rJPw5fgGtm28CsZOr5dYsvN+nbfh32PaM
hl4blPbdd1367WLiy7o0ZjetdnQxdpwlrea4moyd7CzzP2N5Thu+R5T3QHuZ+RSx
ql17nESwgtDEXECuU6w36zZwBVt2ls3ZVUjaOGlo/06YJuUxE7xJeBRDpEhQY5e2
TtKmFQoq4ZsZzJgBlYF4LmxVPZo/73xltdMdzfCx9ZDClcCBMPXHuNdC50Feci9O
yKDAf9qJ6X0ZbQ0pyj34Z4LrfDjQNwMA+TKGRPWtD84VI9YtMgTikqrLym//rsRp
tFKvIXPLF2N9gzmANrdZT2zNAXKDMm43EP6B9t6nY2Rxxh0dNq5oYubwNWRdBsRN
mZub6RRFbReQx74xlmqI+9hyq3S8HvUBcNVUkp1uM94PcySiqHMTedkJcSwTuBlQ
FcncTCxVeCbee79KJR4u4nmtxMNjlAAuxQ2mhG6tdl+G9R5DLt+u1hr7WhItq7+d
d60AJr+pNPN5hQIBnoWPRqAsuFIknqQ+BrI/roeAYm5kecEOhGmT0ocZ/FNBvuL2
J9ES+Nd7NxxkNyK06mLTmoH2m5IjTHIND7YTtiIUeBiHu9FoqGcvzh0XTOw8/ncb
XAToN4qk4TVTAA4EZX4e/yidJHDiPzC85lie9gj7Aj1rm4X+BpR6BTtl8RGZ2NrB
49T9u0ztyRISMAxPt+VqgnOJm65LyVBcqX1RMKPbNTgZsQx+RlFJ3rrAxP+qPO3P
AY3L4xAl9C4N23A6PTXwga5C5CaZ9ShG9E33L42+43dAd5X4nCv44tDxjurbQy5Y
J1cSBLyTTr7XygzhgxhnkVtfSiFdj02vdLLBVAEO1QCZUT2MF5FCpP5Aw5hUItt0
Tb2PJOF/UyMz12IvNGkx7cMZqBcWH/O3l38FqDg+XHjNuB0X/hfnatTr31cpNxum
/nsjN6xmG0YW51thJyJb3nRReuIvjYgAIBufKAH4uYyygUvnIA8nax1BDumVBaRt
bD5Ml3nvRd6XpsUgOOAkH6cMpG38X8rtEi/OqS2JuhOEDI7s0gOKRuGGKymZ/yxy
OLAlhRf0VSEnRxzFeVSsd62cmEJyCQ69nesj0DJH8ogEVd/lGnM9P1DAHCijh6S2
gZ7IeXomYQMnoYPdo4yCaZNJRf8tHV9c4byTn6HZUBSBiD9JOXlcrI4iU7UzGTWf
egJH+WNhYDoG3dkJ7eIHxWjCyXF+D7w8JTQrN1UWMBwFBkeElDMDqTm+8E28mahW
vr9X9zJ7vrShxY57728c3GDBTAKJLTznrU2HV6y4Gymu+HedGhT4dfwl+CiD/az/
DuMK/zaETeBAcBGQrTdZ6usu8N1qJ+K7Tp63xppr6naAB69Py8SqyoWgeHrnC0jW
k7CpyyuTP6ctLK6e6cfB8Bk7iTVrmyNeSr2VNeoxNYW77+xHZu6S+iAvdMmDd+Fq
9KbuYvYntymaGFzAMrMxJ9y7mtZpLhiawSHnRyZbWYo2DWFK42Ns5c5VC/4OX7PB
JYD/8m8w7csmNg49ArCMRe3Mn03O4osiHFIndXk6HV8acW/dJl5yBQgrbVVfuzOj
6jMw8xgB5IAUWRbED9FYciWSdBqGAtFS1aNvwIijfjY78H8oN8J9Nhb0WtnYFNvt
qpXnJyiOgof0g5qLUyT9TJxLT6SYUPGWPwtkUJBNv0gG/Vpj/zHsycPCjHqkflhG
zZj+KKFdrhl0lrdoChjBN3mf2J7JK4N+mAfmA5vkSoeqiRt1Y8zlxHqgg6zoQEVs
at7dXm6p+NFOnMTPrqLEvvrAJNofrljiT8c/UwDbDsziyhYxqJRYezjqp2eu/z5n
P+uPcdQz2XI8ldVmVatz4dEu46LmJX3IBh4zmxVDNrJn6rPWFTjh3hfEFPKMHnaX
QLC9NVDa778SsNkig6sLO77UdBkjgAdINkt8inHSLwmthIGO9DSYWT5Q3xepxKTi
ON2ogqcxPHeCnLY09wQex5AB7cXAG4sc/TEXHekQzbBoyuAaYh/B6aWyD7rpcMB3
fDq8ltQTnoV1qMXo5xsJQZypQ6BYHuYIqxmMDkjnx0/z001ssdkK8+iZvlwT5Isu
9mBrDO3BzPKnq6EA92viRy7iiz/ALupVZ7c7CSdrMafZarbu45X9t7WV192wlE4E
kTaNehGJFPz7qgsYiun5euJVaVebJymYoJkul/tvtobmStP0+6+Hx5l+XTPNMMF2
Y+4HuW9fPggW734XGU81y3A36GNjWEQrHOQkI1HJH5iC2dhlscx/eRX60X79f5Ld
nlnqyMBlDNHbYftMxwUyEEkfuGTQWGbvdq7TW2vEL1IefVAElFlyLCt9Xx8SMSyW
7H3lvfWgila4jZvIi+mAn9ZjFN7f8IEKixXj8gbpbCipN9dC3MPp1+nspAnpIja4
43fO1DDD4WP5E69IXJeLqqhmKkEHAwojFs0G02LoZ9IN3nAf9jvEv+zDpIVm1KEN
WyKtCCDTglzzABq9YeDLn6ozaLhKLOetQ/GH/HGPr4ebKm2G6Gcp4JrpXmPcDZi2
73EVKRPuBKZmz0Z3eKHslnYUZBGCwp31skgETMdYxJ3XPfa/l/bKv6HPBjGhDSBE
5GUv1fJNhPE+hSj9lsEnNx9hWz8McURGqgsKCPfhouDbt3lJrtwnG3Raoz2uafSu
58YH1F/GqthxGgQgbEUPVHU5h5r6G4f+DzqMaP1d7iAGh+5+l+PszJlO7jWAsQgI
i8/C83uFn8N67at06KnNqWt18z8i8zyA/jjJWqk+9/LiYnnXb6b6Cmmu7+dpnxbc
I3ZHbz3V0LpJepAm16IFjzihIv9RcVCdDfZVbmAhKvGVlJGOAMCrl/v1bi2QK0+w
MBu6QYhocwetiyXIxv/rwyMKRSAtCttd9zJ7GISTSuaODbLbwzRg5exEMn35J3px
UkK8V/P0+noHp2QQuat0UCAHCo0hdZjLlhLSG4PHXhd16Lo/DjXxacl6A+P/JKnG
Q9CO6CHN+QIOn2yqWyddmZm+/RwzxyAqZN//ENJVzzFft8n+1kzm0Zsh1w1eqrHr
SrcrYUhhWGUtKB9kMTUpsgP/QCfDkmP8/AhquRpukbnRBzKVkC29CErhE/TvoNUp
VsK14q1pebrO4cYfQHqx/ax0UUcM3qwbKt4xEScMGFtfXiscMTfyAYSuB6qw54hD
J+n67X11JExSxlXBJtfCM5CRCp8Y8RcPDz7k1y+QY9IH7nScA06z1l4qC5UlgBuv
IiHikCdUJkg1Wyv6oBe/ElScZFAWnNGuPZXNZIFTn4Vkfr5aA8TsBlX9Lt1yGfEc
PFbsIRphtIl86PemwjCEXhdIQ37YQ6mfcUl6mq3UF7gpBBpyT5b9kInD3pMdaxS4
gH9NntIe34U2bJYBRHBJFszZBcyNYgQX7zegmyz5JdvYre+EeJRweK2jwQXfoLiR
yNHf6abkveZc045WdwGZdsET1jUTeKBHgMOp0NGf4Jibqrkt9gACzaGrXxOrJYZY
zVeuQp60fgOv3Oq5e75XHVRezmm4e84pM6T9VyQxh5TkJZ1cb+HrNo1AtiijVcvo
zUhaRyonzWiRffGGV9RkAMzu1fQmvkqAkiLRs1Hlugb01J5OXiSw+y0UT6BVTOMp
yryLZoRUcjWbZsxN77nLSEVUkP5MQrD+OTg+EDyLEWnohI5e8/2TsRwhIesUcVZz
GA33imPB6c+BwnXOkghKy57utvT8ge3EAlpd02LTuRreZfkUumr+fKxZEFBw1E7G
vmjXmERmACv97rWxqDmGtXbuVQpSN4ym6aHHz1ld0WKm3en7HEEPtSz6lZ+8Siah
YGyNZ2Mo5PCGrEeg264lFt9acm1+8G2/bdVguiREVO4FM2OBDWR8dFixJbpko6TX
Fh1M2F5S9dlDSnILbX56TvF9ig6+O71Wb/72XRuxjevER0CPZArmhQnXsdRlsq3R
z0xI0VmmgzQ4jBMC40kurREcEG3lEv05Ou7+OSeyrVUd2yTMBaU5FVfYualx11JS
TvBZ5CE7x6Z/72EHpIBp1Py2cSMYJ4/PJLAUzRUEkuvvlpm9LLGIjwegp2Xg0A8R
UjeutxU95lT80nFcN6x/QrVB4Eu5fkjhYQ2mnX1v6CVyq4uHKYAwCGwZBlq+Lfb6
xTKL7Bj0VgfE+IgygrZofi4ELgMIeJ0Eo06fcv4amURmv43UDFfSqPK4o5E4EGSU
KLAZvg9UZl+Bn+w3S+FeYwgzwB15Q2Ku8oJh5/FxOuumuuFy3Z7ABXhbewtHZITZ
h+V+6dFYGytQ2cxgf36/5ONNhXPA0evEWYkDg3TSj8oUFsRKht7tQTRT+hhN84vj
s/T7ZwfO7Bk6BYwJO76NZMGvCiPkBS1AoT22An/AoCMNmZkbGMg9zaAtl0LTB8b2
wTiLhRxUGTxLqPBVEEYZd/MmFOEaP5UvZ1M/Kwr6ehsYK4AfRwgm+cnp8lXiS5Ng
68GngQFk1pk7lgLDtlRmUk0fLnkQI4lovzxfMdaYFWJzYVatO39+2t7n0maN2UUd
uEZhWILY8FPitbsjrkNeZ969LJK/OiTyTmkxTM11aUiMzQjTvklGB0kAiDHVVRYR
v+FdkQ7loF3JwtjzosSM5gE5zzueBc6yHuXInjrdGagZrOslG02+xy96I00Z/tTM
pUxisq56gYpdyBvQ+wF6kURIoDKo8eSh1CVReRnDveVIQ++M6Os4yXhR14EUsGU0
c0bHzLb15tcExsaHcd1ijzeF0MMEKTjMEYbmsjnIeiqv+s83bQxo5g7D1blbUFqQ
Ob7/fbp9Px/9Up56gybNUw4zzJ3E04686fOxi3iUvD16hKp9Ly7M46zbb8h7QGan
HHV56QYDUajdY+4frae1fVScMHftQfFL2k/uEGwAuIlVv5VmbTrRURuN8tvFt0sm
yZXmss3aUnQ055MHiZCa17VfjyJOMUZb59CTWJk8geE09oqY/61t5CurtY+D5XFu
WOevzyS8qYX5vWi4XsFbp5OPkqk9wG8CefP+ROwUQiOH05gPPOkZQ2GeLr/scFri
gnejvsROFGN4AUafTa99xikdKx2cUroxzkksykbxdfI+06ov8Evn3S8fILsO5Qtx
dE3UKaKCHfWEQzj1wJz//jIhUjUxQMN6p+vVX1/LT5qOOfhaycEQLuNkzZVcvs6F
kSE8tIK4tv3IexCv/5jyiG5ufKZv6vKvEvIunI1csE8a8a0XUBNgZ23/4mETRKUr
/be4RxzLoE07zwF1hFjod36Za23puGOiBDC0cFlvAwsu/SpMLhwlyXFrD7ZywZIH
dbnBMyl/9wGrOctvFh5nNC+hVlD1CHiIbzY1Lu0e2CKPGbvFPdpJQ5kMTIvi238j
M8rTEXeOItNU3INtkOiX7VXALq/tGsCvACUOi/eTWVjsrNIbu/HR/Jkxws5i+XEl
nB/FDwwga8f+z1maIo9yTIT4NBHMHPwenXaUP63891wdgjOcl1P2uEPChMYyz2Mj
XaLm5NNImdf8H5gEd4rc5QSyagkRsRgHboZD8MRokah+b7MMDhm7AzsNefRtmtBl
xGu74un09qfHNQWcU5ZKIYx7clWBrQ54DUG9Wr9agLmo4lqE4yrUJ8F0/GaIdvHj
Ii/L5Xluhndp9mRh0VtcKzQQWyCRiNryI7XAkuQqQAXNlPeppwj2S8IqGQf1lV4I
QL6IrhIeWI0B+o5TSm9KD6Olzxg7BHuTEglheFRB1ubirHqVYofUnfnnLfc/+aop
kbFou/stGKVSxaZDlZ2H+MugMy0zkdnzWPvCCjF2MCzYGfP4jw2G3qhZ49rAetMM
X+PVWCQMXp8XQUc1xJoTF3+yYvI2K56gBswjSHNzF29dWenZAqx/nrc2HSmCyhKX
d1PjPuXkAGNfa3rp3GTd4Bp77StUA8rSj3nx19unqpdsuzJ1g41FL+zAVfDNOdBe
kz64UU68vLz03f/NCN2+3LFnYGbd0reh3WpN6UtXJ7WA1xxxVr0KqIqmwq1FZwOt
4Ztu+MU8IqWvrDo6mADHdduXkwMhyLwS1O0KrBmfE9HxCXM1ckU9UyL/P0UbGZGF
Eszrie3rGrmbZGU4TsRNHkHsXLB+NLmMC/1fUSwp6PQGOt29XWG7KayX8Nmsg+1v
ZxR3LA7M0j+07QI7wSLHhjOmL0LABo+Pc7Kw091inB0UqbLm0od3/1z/k0pK7Lnf
BNbCwzg6W1rI33KXUbS/X3RYVxzUd2V5NHWZ0b3+TEitA/NUK8J1TUMfEoV3Rp5f
/VqvyHHWG6Lx1LohdOgmkpkvXUKMsF/T+04OZtqjTBpxisRhyoikGUHh80kRYtD+
dlIQmBDN97peEez6D9WK16bV/xsJd2S5JtjiuYjFJDxHTRrbdbCG6NWmikhfZXK/
NxW42nv8O64TBkC8AHpl7sTCW4CX4phDaZMUXrM/b9xSA+CPuhsuNCadUSZj3VRv
mPepEyMpI0yLGpwRDjJJF+zB6gnk5OlbMTC3McdzyecZsNpCRPVRSR/aU3eGWkF1
fkXiwk7lTBtlV/ArhI1ClnJE5XazDJikhkN9fDoUNw2ydJb7dZzs9Ubk1mbxl5gL
LZmenHhQsEybOm8dWgl2BhiFtUSQ4NfwWa0Ki4gVZvKNcx69jrM+mgOWOAXMy7Md
xLlRX4YyU4yxdJi9Z5yihy7gxhlFudgInzlnpMPwk+UywCzCyTemVdUOki9x86xW
qm3NfGscFJvoO2XplelB7202YjtkSfO6BAkS2cxHLIG3EVy127LcDMtWh/1yZj1a
9F2UnnkartwscqPi3FbUAXRuwGJTNlSAFDdyHFg1i3QXIOyRxehR6BjWWo88ZJNy
dj/DqHb0aGNFjGlWV0p46l/Pujq3FfAv7LEbMkUcxihDheJlDS5pGExYxcxL09aQ
6E/fQnF+BLzOQHa8Ha83oaIijPso0Nx6TRMtKbfC3Pm9abhL411ZyW8fWJf9p9lt
OGOA3j++YREEYmPcjIXUcko3zF4N/7dfz1Dv03laa7zCuoS1KeLYeNJF3EhBfyvE
XKx28Yo0Z7Xrw7Nkiwnnq7D2ucNw95MjNJ1Es/D6sKGyVLGZcRNQrj3o4rDKp4gy
DdvuRcV2iktSiEPrhdeN18e27cbbcVUkaRKoPYXYoi1JZOUWcjx8F8Z3gtxRx3fH
KSTuyrogSQIbZ2gt1S8SEQ3n3c2BCHF/6B4HYnO1o9La3aN1kDXMenkdP64dnYAY
MpbiKU0Ew93HhGJwlxePhi+XFR0sKUc5FdVFmRUtUhKPRSBCbzAFqF1jKudmMW4j
0NjOgWSpcW/2zE1B+Aa/vbg+UWEGjiyMfocbBEcm69aQFiZ1if3LvufnftSdyC/A
mbkplx/KqrQ42JsLDmgXoRa/xPqYKU1sCJ9xrzm/vAUhDKX6ru6cU4W8Z3eD3P26
ix7dqbV6ZZfxbP1JJ9ELswCR0TtGOfQ78oM904M3ey7b7tut1IjmU6hsXkrpBunF
bG9siKzPyVFMcN1qDZIs59qBlmy0UD51++jsVScMYAWK6HrIgxwS5okP0gdw+8w+
uZDeq5VozQ5m81Ud2z/rzUkBKjSAVKvVV0gfV8xvN3Y8y9IK+mARKfDQi1HB0Qpb
NhysNLW0okRd1N/nRdH95DDMkMs0/U24V6FI0bbRW5IXVaViBzX4TIWmS4rcJJjo
l+fnoa6YNNs0QDMCJGpxAhG1albnxXhWwvuXeoFC9T24BEteqXRaQcT/JxxCxT4/
Jmt4B2SjGOOlZfi9MjFywH68eAIYeQD3YRMqgAfFw2RAThYhL7fAt1amLHXJLwZb
LKypv9InsTq9o3wt3v10C7P0Ly5ovaBJjBCPAojWfphca61K33PatJVtS1V8AWr6
8Xb7KdeKEHsSMm59zMNNqQv1RRiPxO7DJVcR+SeV+NUmICj7GBk25+ZvCMDqawRi
Z2OzpLuoEI2QbncUKgOnravGfF5eo9CGyGTXG1m1DyMX78D4PPUuJ8S+WLYniCkC
oz/veq2EppCREu+gBRFltP2VJWJJq7Oa2BQZJJCIciv4Os6ip4JaqB2dKgWjlvDc
FWHzayKCgNfy1CwHPWPqrSk3YXPksk+bOsUjS1OeAJXIqshoIrZ/jhmNVMEglRtS
S4o8xeLT1eY7PQ792EW/LC0kezH/B4mJQCDaZtbv4sZEL9ZnuUKr4iNFk/VnfcBf
TP/txiuo/EY7DzHxSBOmrA7v/OvYV5tSfZAEbPRcifuZJeTLO7vzef4KpkTLEOsr
2LvYdIh6ioqRocD0Y6ouVVJMZJxQoEWqtI6lidDMMWUB8nqNLx614pRJ/xQIfP8h
3hwYyj0Ja5iys5Re0GJYluNFHF6qlxVyxe6RSgznrQAAdl06IfL9DdWoc/5+ucpM
wNP/yIVaZPQYTwoDFtoBCL7N5+MHQsIvIYDyXxC8K/1DJq1NnHYtJyB3QdyIIXwG
Gh60EpT2jdKCruANaUrfImmM8yQgsv+KwNrz7k1D5xx+l7Vvj5jlBUnaCiOeIXnZ
dq+5IUQYmwynITPCUJt5fFr/UHI5svviczRXQoewPOD2vtq5nZkdq163b41UKJLF
n6+wHwHqlhhQKjHkzw6tBfgk7Mt97sMC7rywaT3zCDVCOyLkX2krNrZ5SfdKvIRW
GTvQAEWRRn4e8+LXADnuxq6Gv7M+ZDTWqURIDehSm/l9MITA7dtfHsDVPZawYsrq
ZZ6GoxE6g5EXX7ZXCKFttI5nxS/RQgmxmvSqKKe60y8OaT4wgO7YDmBllhaUpUVq
ewLo3u0dk0LU+08ew3U67uFchl7cKubTaSU4WFyui4lfalM8iZk3FD9T0YkuCoJ6
/tYqsFgGs6qVNu+uT6HtCvO6rgOnbTzE2zEvQYzhBwR3sLwcqCu/4m2SnERJTDXE
xZPvLlFacnKCL1ow6D7gdIY+2JT215mvA4BEeEAbdHYgOK/LDDSXPSMcxAIkxt60
B1m0w8GhsMSC7YYdftyfDjjEyiO8C0ZvYS1l5TDv5R0vrezWlrLmjf1c25uRv+La
/To7KZRdyTe/C5a0if4DrHQ3ujqHJD1PY4vOf0SzEgJMKDtNf9mQB5ouDhOQTTkr
qkuxBftHG8kQyx8Fb33DHIsiQ12wcFiTW1bzW/G8s3BylBffLzJ0GBGsrn22i11s
eV1BL4Yp4TjLO5K4da1Xi3p74CkT1dzuHhjKLym4+OFiRc3VF/bxbj6c5OYcbtlS
L7SJ83O78olz6idWykQz0fdiNuuR6ZXDpLdDVstArBUEKiGBZXPjWbfHZBgbQj9X
KyQRvvVUIrtvra5Pg7sbZW8BPn0eT6arSt8uLONYHAB1Zx8mclNATSHcC0cR+7Xa
S8jseCdU0N5AVmqlKGBeDbSMDt/HDsXagxxx/F+IFyC9ei/qW4FcH2IfBzyGSfg+
zPiKNmLp3v8BpB9l+7QVnXGHG9jptBYU3ICg5UaAAXZayFi3LZQNj4iaBaa1JVQY
Irk+y2asUqlByT45wam9xudE4fD+ZwjUmltxO2t+jMfn2OTz0tNz3iKIvkOlcUO/
4OHClgg+w9d8CR5zy7eIfg1cPb7NIl4j/IBu1m+T/6NECePawBlSONKCRlFpcBZu
ZVD1eydTziQ916iGWScvE0SKex8vz2L1HjNh1cHIp07gEb5vWvQWbf65d2h61BP5
PgnYzwKS35VJSbxMk7I8q4iX4/VufITZaaMynfL+G9HitGtGrl3E4Iv7QUVxOhLD
41RNhfp8TO4TIo/x6+Z9UJqS5UfsMjisIPGl7Y3VLWFWQJIKLQJocQxVKQ6a4Vme
d4dOJLj+P/lJu3gT9oUyVc3hg+RkPXKFHk/mm+nkDXEmAmmg+pPH+yG0WLYMbHWK
Gx9Ya4PKcw6G9PRm95AFHXp4SO65ay7FW9QvlEgW6SCW1pgk5fLjEutmobis8Axm
1+L5yr/xZtb+xovLOQl3A4YHZSkWY/w/Btxg+SPTqbSavXSWkdIvYeEzNKp3E4Nh
g+2RsGCbc2j2HQV02Bv4A5KWMXjueNV12nVxiMf+JHFcISmu8VPDSaviJYy6sPNy
X44NOXh2q9u1/hYED2F8k7JKYE8PWlOBhPcWDG5+PRBlJbopQBYl00b29T3vg+nc
5r4ysYkru1VHiViKmFwJaKiVnVUsDFJus3gdSmhWiPiAEO980rLO16YEHrc5LWqT
fLfSnnSr5ZbvosL96TRN9Fh9cw4a0NgRSfYK5FEpQtxHqB+rFxSOYFjMyzhyMmw0
vxLbKxm4oFS7IiduxZ6UoneeTE1wpAnjtl67VpIVeRie+YcLQfgwP9jRY9VLK1j3
UykNGHgZSpsoNQuoiSnRv2XrphDOEvehTig2+4Rw3PUVYBJv+h9AHe5nQBpBcQZG
qynvZk4yWZHgzY7GdVdW8W9VOuZ5lXCgvYCJwghFD5rO35LfyNAdcNySoMGsLXji
im0LJFD8Zh3cA/gBW3XqKrWzm2CfpxzssJ+NWSh8lhlWnU+tWKo5Ibm57hXyQpfn
dQgLaamn96bEorDIdJHPGeu4xtINzD2Q3tb/T0n+m4RPJP/obeMOVOZzZBEQ8KYt
JyY4L1LhjblfWfFG9h6nANbnX/GdUcFL4/hGB0fA6/+qFZ3aXdTHZ9Vb5GsLR9ii
BzrTeel35G+oC/G0WJtdaHxrLDqr8++pU0gdMw4JUhcdIJ+liR3fsgdOMWIBeUXg
msiKmGh8EmLmoywALymtREs+cUqHxgsK8fYWeId6CwFN/svsN3FjBkEEQj8D3Wwj
3+0rQLnGB6OlpTeIVYp6Ydz4AWey+mhAcHGBcYhNLLHTAg91T6R35DhDWuzHBb8S
7JMFrBPfm0Ci4mgI+at2WWtGh6Ki/tej0Q7l8DbOZ+S99IfceT/xVkCjWKKsznf/
MTBqub/aMt3aq3A6cVPffAsQ3ZMB7dHMWihzSagDAGsH2jCo35m1w1NcqYbMPz7s
kPXuqUp3KHK7rfLK7qykhHqsoXg8tLmASAkouyIWGBx+vuunBZGjLO5sg0bIJTCC
QVsbT5XLeiCqW0ppty+zbBwDxMOpKHiA67Gvxe7pCWnxMP+ftEBwG2qtrGv0NqOz
wkWpf4H1Zk0IKDMSPCR1xATbZWQawFdnwn6PT9k089arPLQbGp2eS7ZUz08XerN9
5rVM/3a+SoJx2t546L5jyb8xuCpGXGLvfY3UjklM5mLj0UWzafdOsBc6Kclg8X/S
ebNBYVPbzgFzkqzZMwVqgW7gEMape98ogEMNio4kC2p5JwtfqcYWOdmt9huWWRCs
MvddkP2Rzd27Bsd3xHLdCb/oxp9BYI/WQjxnAZ8L1xP5A5zxJJlGH1FFF2wlQ+6x
UhTLrer3xpTLUoVDvZJG0gHzJPvHrMJpdFYc5jMnFC1i4BPcP/9Un6MwXORQpSPV
IOE4Oynf5Dd8TxDiRjMOsSeBV6b/n7k/ZBkuxLA5uDIxXB5TMLeM3VxIEGJqAsuZ
PiqndGaCvMCmpFI59tJ59iQ7j51xUhlaqUA4wNcGXHdFWUKKBZm1flPpFG5s6+FO
rh5cmIsU4IAtj5UdwW6S6JItp5Qhkiip5s5erId/l2uC6s9vX1D7ety4LOmUcCop
OaDudmCYkClOjAfdFxIJlddQ0YhIT12+W5Q+m1mrHoqGRAy8cotB+c87/v1WF0SS
DW3+am0EcQY9gGzbVGp/+a/G0tRcNVsiTC1CzVbafHySc8sWl/KLgM5naj8Ei1Pt
XNvVYEr5BYQd4iesly693twpNv9h/nJGfXPZVR6x8OukfCUBr8wXsjQ58UvDONiA
T2M+NNoFK68ktgihvzvtYClvllLyuq12ci5rtX2QLhrX93WColG7dcy4JYHmA1CJ
uMPn3Cq4GcF9U+mUWmI5CmGXZON0O+UCMZi3hTLJFMaqYVO6IE+HJdDetg+ETxMs
deHPQrYXzPkTSgIAh3JT17OLnq7ctRFjS4e9fF6pUyWDj+FP5V1xcJah7konMMJz
SFJBWwvKW+AwVm5iR+as+0hhD3KJbnHz9M1MCXPwuHRdKYlwhXrlYKp2fLa04wZI
RkSB3Py85iBdGD+F0oA+M1hnJAgljl+hM7YPeDk/gQA3KMW6L/oiVYAR5XMNuK07
KV7vBGTJ57TGYqgKoMNBjymNInMzUztcMblsV/Lr3jxUJV0diGHJoQwRqILdnqU0
KREgNeOWijEQazf0VxwU9nGR/O83J5ZLGfo+ZfHga8exP+JeS5+QWKc/d0bEL3k+
SqUXpACaeNpGu6hQDmmeaFrnV5U03K1BC6jmHxJbVJ23t73cfhFHYD58QRgq1Cws
uCoGGgaYNyFb4z5oSJg+hFwMSCOnJW85dL5B41/2kLDXmdR08mJQpRYlHEBXTdpi
74GVUYrBoWKmOHwU8kEhoDHfQBdM5c6KldNxmwPI5wNXVAaVj2vQHLqvDfF9ERTA
PWS+MN4flW7YAtXCSv4XbgLHIrVY03y7Ow46eS2LCSyagcEDBjfHLUWtoSa1VbTv
kfgWyQPoH5i07sSLVbJA9chaTMvTf3yTadVI1pJiQaiPGuerqDjzNFcglpRWGr9K
SCAEBz/NlIJRRRtswMI0DrolI/xb2oylla/9bvbpDnHheEBIEWUTTIDoOPoc0VxT
6SlOgEy/enNRGRppygQNiAr+alHbsamwighT+HSAD1kWLI46I9FUPqUbH6OeGpPL
7Bie9Ggy3DVl/cIdt9VoUKgn9flLitfGNT3wWWoTAmQQ68NfY0M/I2TZE+XZIXKM
WHf0iRTRELe4Z87HF9fdsTi5L3wJjvfKI4NlZ3z3dBrb3W/1ZpWSloBCWyDgUJBq
YR1Rlv1Vb/VPJ+3tbZDCvs0hpVeTVmXVwmEv2my/Yn2xHmv4p+ne3Whhr1VLHdAU
SgYCyGH+9spzVBU6/kCkIKVn54xAmzbZz1ol1IBbdMUNuL1PNGwah/4ecuJnVB/Z
zcErNaJh+pUCCqvx7lDKkNn+MhoGgpzyC7G91ktzJn5KqBT+p2l8SylmFOeNXFT4
GqQ2JhI+isvv7Macxk4K7S3Ab3GsEdYPR4xeBTTLkYPpQBGbX2Zha5yyHN21FmIz
tOV4+MD+FY3xg5mQ5qvUA60d5VwKUcOJ/Prql/dY3GFqMsZWLyLtZJAR2bLTA48n
SRx+QJk8m3jNTmM/Iu1xGoRW0aLKzu6HNc1oNTey16gMYkjFrNIx5P+eABVLqi/j
sjyWwxYrgRswq1jZAA/8sq8JVoX7OWxEQb+NolCbwLe3cu8EW/ZHP9OylmAe3YVO
1ia6CS/Hh/qbcAKqujzFDUGvXCMsSdJDMi/nIpk5voHf+YEfPYC8goPSiscfkvUu
4dyPQU8btcN4MD0VfsrW+yWSDxJcePzoJ7rkuJcTSshn5/SxUflaM2cgv53Ygvkp
qa1VmNkZeNJrjqs68g3VVImdedl62vDVclqZqNWPhagNmefPMdyPHmYVhhQ0qxy7
7Li0r10igWNygaMkyL2K/KglYM0KkKVvb3fae6/WAfXJQP/lInHjdN9SXWpyiqKV
1h5X9K+zqvsWSNP/VWI0Zg+TIvNCfJPeWt35E5kmsdnTe7g4H6lqGmzHcaP39WS3
yvz4bdoTrhxE0PVcA/eBwcwjePmjLpUmnCbLZp1WaZKjaU9qUdRb3ClJm5PQPmQY
LU8Q6KvJQ6UXc58vUzkrOGCJ5xrosFcgS1lmibofErHUEr1bXBErVs/ieBvAA2PE
zwcWgpDfrjl+d1IhOkF3KpcNOAPIWOKIVZTifF05RgBTyWfpozjw1q0Shmw+VqRX
tuNWtVTfCDfA91uuoql43Op8v23oRK2qsOnzOmZwrtUuXzI5Gad8yTSL+KKaAAR3
uBclWXe3qjrvWn7yQOfFeCbk1DT1mhXdkNor2nKNDGhzdjA9H2oIHbH/wx4DKhRJ
l/akwxy8yehMTpvKbN9h32OEwg57WIC0sy3pZWwq6GP9/dhfwdFAThauOAooMNsR
j7SDDTcH/pHzd1hA0lnkh1znwSVr2r3AUG0nDmAwTowf21w2Lj4gKxA3iWEfXNT1
zWY/uf8yg+UhIZJXuE9+c0/suvYS0OkAT9DaX5FxZidXKzezEj7Mwlvkbaep9tUV
cn7civ8EzUwB3iz4HZ6xrOTCPod2TAowAnO3SFyseOeo1UgZv3bn3MiON8NdIUYd
S9n0A1Csp1zAsLm48n8+Eb5Jrihmze2LkH4dEA10JtuqlhcflWR2h3Y/QuU8qRpB
qB9iT/Z5pWoQoq5pgI6T5FAB3J5xd06RHVrSPq3bvAdXA3mzrgDAxIQzSwGnTfFY
A4xjpNMH0xJpelAdVaz0qP23Wth77/Q6sSwMvtwQpapRxL3NClDg5rzlM9OOPnHA
9UhnrC3lZYYuOvZGksyOabDREulOMMtwp44WcbBbHeiKSXElyviaeveFVLUs6vhf
Tfq+0FppDfdkwxqLF+71qs//cUNyi2ykGUrjqmz8DB9Au+7XJw14gNcSyCBEZQVT
NmB4v415MsUhG1xbxUG5ebSzHN4s8//PP/dy3ALMtP0eePn59vY4TpY72f8vTUUd
CVNWH0awL0fTNR79Yx7ddxkoB+uS+1mKS9d3/W/hSSq8eenGfhjt/dD9mSBm3JW2
yAVp10fec12mV6wxApUHk3Iw95DGfo/AZbtwyBVNd+x8YTh+3iScGurMo3szHO0/
lWUVl+pZjYp7Z/3HjCng+KAwdt0W+gKfgvEPIC/+W9/74QoYHGfntDCUnGcLy3ps
Qo88ri45zMEAhPIb8Z3KY6wc2EDfO4gkc+aGE/SYsaYzoqjFo1kPXO0Kw7qF4oSU
1Y8+GnU+AjJ2mJkURmqzobHsDMLoQrzMEaqt7R9gQBZaYUFoPjYdWAGS8f/j/gff
kLAciRywmLIunbJ01pTYa/4Q30UFQ/3E6POoU3QRXfUSw0t8uro8WsQSWiiV29qK
NTzZIbL5yX+73K0rw30b74gg/tL6YoUB82nNBV5hRsBYFI9+1o0zNR+nOS/ob3bb
wsHVtHnTfGoKfmpGDBuXCLWAKCa73Lmi/0Z0B6i208SCXbN5O03UeHwWzhmC+LbX
+ZNNlr/cz5xKhsaWN+zbDpQdDLoiHGcW+XM39q1yCIcf3TCf3zdFIV4HVBJl11xp
jRvjnOkF0HBftYyFYcxiPHyPyb2SQW2RCwO+AHjj+gCOZIk28IWEdiofCy2yS3n5
FQTSF1Z26Cn4zYWz9iYytm8wmAdrITQ3Y4SmcTtnIqq/jp0/E+rOPCVFYGuLSNvZ
c84iwFI9ull+Y83Q/NRicX3WLAIyeRp9+KivjNWlbmrZ1f/T6oRThLNBIGFBbajF
fTbzaN3o9/wq95B3DB4CU3Pl47qavK8nmol/SiA00Mq3bBT7bExQWjNsoTqUSPUh
pAVPUbyhO8dHzlUqQKPPvcVGn8isjHQtrDgcwXSJP15RKHMWbv8gJRY8RFIGUHYx
uFLdgadXId/y2MLj25TUv72L/17U3Uweeb0uQ6QkPUCGTV57vhvIMz2Uk6p2nDPf
3BNLSF01+6SPudaHv0H0f1bfo8dkrxVW16hlpPpfTuY5MezylnLPmqLxOh9v/cqa
qJTOzkrRf60EBdebNHbWo9pQtwTBOoCN1ZR3cIaITA2Eyn8cCrSfINDQMfu/b8FH
V9FnTwlvmYDAqg5v+Dh2w/yCTOx6TpJxkOWHl0wDgM4ZpiZDXcTdQL8AN9dVwPF+
V3IZvhRAfkQVFE+6E0fnJHhmg6U7Ffk8si1mCQBpCYJG0OWE+Dyswp4yJJQBKxh1
UB6zekJjc5emuVi6YIUdjS9c77KQlg+aK+XNwPfpHQb/TRfoKS3YXet4rrmqmqJO
RwOp7/2s1WH5/tq4OlMVtBCzuxYqO/6jsZK219k8FXYFT9p+Dxag0LeLOvq0myFk
HndJl1bi4H9Lr1S7MuIt79ycFKPPRoOqKfWlggF5uB5EZVdu2gsGftvS/chef0LM
vJrSzB/iHzIevYKqdVmDdp68uKRMmpMkBfSIoGgVffTmy/EFVbaec62/lXlsKrH/
DUynPljI3GKrk6emMfrwsucn8qjuCKSLBfRX205/2Fb+Xkp148LGoZpmn73nwpyg
CozQWV4Z/pvj2iFXSglVsK+MIvcUvrvj+h4KOjLz4SftW2VGHIvLPqHcOUnnu7hD
nKAh4uzc9jCxaRaBcurAkWzKT7BMhKZ99KKfHnQ8QbhqMQQNg479K2n0b0mSq2IP
GxbVJoKDd4rSJugLSlWjXJzMBju2rLvu4+ubFf3vRmFYxHSphP0N9/SrggmIsiJQ
GJ0PSaHRn2uqc9892kEnB8rpJsDXCr+qfRqGN7yemU0wehZvhC1rYrr7cEgY7GaH
jEVikHmeIc93tLaT6dXzMnZ4xSjx0YGICpqRZSrwyUkG9GdgfJ0E2iJtRI+3OJa1
6k6pY9YNLntgDe8uTf5KSzkfLJVSF0kH5OZcFQUpNhgr4pptAVpGMeknrIDy9JH5
1EyG1hH1G67/w05De93FDIKEIkJ/Xu5NEUvuU0SHnyp2ORnz1x4h5Oi+NXzVican
xeJaW2vB2Th7fXOYTJH3urpYhoJv1gLlEk2WBXGDbsMZwLYKxWx5e8KPJsLXDtvc
gYBmvd+aA4CU3lox5zrX62D1DbWbjvoe2IFBcVerESbeoIlHWFsmTPz4TMpp2aYs
SHOUa/VGv+ORpuBsO1zUfmIQ9IRztacIbE/EVJixCGaeG9sTQavNisX3lDW64U96
Z3CtovYx4L5aTZ63fdrCdjpQVyCOPOrbcuGkyA5d+4aYkCK8ok/r6ixqwSU04Izu
DSiH0x+V8DdbY+WNjJ/Grc6TkMXSDr92j+bhd5N8yojz6zTK6mHl980/q53kwgUz
ZGzkn0SqsJsActULtQzF0fhtfpbfo08uw63+rvzS0PucCXA+T5kbJeWXa+ObbqOV
wPoC9mZai9vkCa5sAvcDBkoikoOQFrhIEbXSdXrTJryrBKpS0rDtKLz5RzrEdUK7
9lQFXne3Iju3BASA6C8plFDDA9wNi2RBKkZf3/sINz9X/LcXmnPsrUjauM7ggZWl
5/qzAP5ctmVWFyaPrURZmMaLiL8rj4vaLn7iFM6hL7E+iSxp7VAMChFT1y8N4BAT
r5sDmbZCYWcPMx7A0xqWD31+KY9sOqB/HBqjFsBHYR+QyHR4yxLXP2cJni6cetUX
pahYWG8v11LNP9q8arg6DdzYyWmYBilKe/Ht8ZosA1SWXykwXD3tKPJmP0ttWm5x
wQRD3Nc63fDPHbLUM96EIgIbIKQpoXHIwuSMEoXm2eCMaBqmRKTCvjfvL0bSG7rF
mNFI1o2xT/o2lL9zpHT8pDUXa5itoiQo+ocHMw35F4Mv2iIA5EMMpnATXVV74baD
mn+OSYqU4mKcB1ampi8fIMIY/hDFQI0ga3M5DgZC04nx3bDDe2qXKgvhIlXbw+BG
qNetczGi4dx3HJqUmOI/TUapGVoQP7ehKu7Y1Cyt/WSA8VRZoDVrjrGsGNeXTc1C
T1h0kaCuUOu78Uip/fZuWfkoNrIpmTZJg6WYLNNw4mM9s5cd9J+woEN4TA3td9oS
BFShQCMlw8dhj+IlJicP8Ze9+nd9CfQRFSbFi2wOGE+6pe7xyoMogX8Mi+4q38i9
AkYl57MtmRvYda3wQI8DnYb++cNOG7QFDQpVKlHNvZu/fiebz+xnaqH2YT31GlY6
psG1vwkptmArfjAc3ZvI2nb2NVx9A5dJ6vOauZIznTOMM2ToYjh8iwM1vmopg5LA
tB/mQOYN/fOhvwnZtlkxIH7IsGsSx2yI5t6QTTQ3qKbja6zPQIYylGCyKwESE/wA
BWZ1zRGvwxBNt16Hgv/mJfttFGoz0TMTha7TrEUaN9kbD+f8QgacAZ+o3EWSW9z5
fM3BzdQFJRZjCVMjOP5Vb39u+EfV9ssPpYjkVwHP1wAmDsPAHk3P9dGyIiGZ1fWO
kOasPKUwxHTpAvoGAqB9+vAapgDjx4qp/44UZd9Fv1XfxU6vKJHvhU4UwAEDIGwy
hKkmayWLTuEcz2XMdh+lBfY5kFpH0nFGjwYXGpU+ryMu6rwjK19ffZxXmufwXxmb
sTyLEzdFGUQlm/X17Ly0pg+Z6QofiAkZzxEuI8/VH5UUnGotefX3mToK6Zk4ogNk
QtMdTIhLPCo7pP8vQuiUNjXlPPVS0zfakbbwzvlihcYWk7v+rPTSbLGthBW73hv6
EVWC7iuA4oGjLGofvrGwQHgC4yjxdizuyTz037HNNQEKkLNjGsIU+f6bKy7NwN5h
QEIuj0YdcwxQ+/6oc72RT1iddsKOI3uKt14WG/J+r/vkqsUJtyD3T5cxy7nmQ5fv
98ENeMYqQmOIhn5wV9Zq9KqU92FVI9UktrjvMJYiIWVzwZrQunupzZ3QIoiFE9qT
BmKEkMQ5eC3Mp7uwA6TUbIe1D+Ka4mxpE88rjPkTgPN3wjpFvGBQv/pWhVp75CCz
X1NhR/UBODpDLtBEorw57eiCNCearkOBLEoOkIr2D6HTvVaPFgeE/kPL01awGHAD
VuKJroFvEfjobdpFIHPeUhF09XhgkI6s1QUU3ioKUkz3D6NqPwMlPCvkyA8W+upq
/YDO9IXT21VIDW5Bomj7ReIg6BuGdqto6Mk5gZWSUTMmx9KRXjGvP/yKp/ta4+yt
zZKsrpifCktWpXlepADhMvdvedpUl0ItdXy9PMitO+Q8+uG41lSbhAUTgN0pp027
VvPf5UhpjXthdiry5O5eAuCBZK2MN6nzj+LAbhERRqI5SJ75zJKVDdsI/r7Kn0Fb
eYioiBp98+CCqp16KkqGVZH3SSgYqcpB8YAzxW398NeWT+9PBH4trm7ktFcYPDaz
ba9/WgAcxqSJthK/Y9QBybFCfM8bjAL9Iijb147mlbQXFyj9Sxo9dDOQJ1zRoK6o
1snNF945dWPgjSMgTkq3YzBBRz3mxY2RhsnJAu1Y6iTOJ+P7W/KX0K9XS91XmPAg
IUsgvy/m6IBkgFOIG1du7ZeWGQEnQYIajPt/DW+5sMBlKIa7YbnSgBbXUrNJZUWN
mbnn05mby2YP6/q6fApJT1uDTrzcRf32WQBA5IdhtxssH9YUWEnYcEhBshmFMf1/
9zp+T9EYi1Cs3ds7TsJXWfH+B48wAQ5f3QBvrE2p1ADTMMFDXjLU0An7rL1+6jPE
RWQxac0Iy1SPHvycJd9DBVsyfa1NdhIctFPg/ncyi6173k8LcufFTsupyt3zeF/W
C5YtUrmPKYzZs/0oos3hH7wRw0eJplwiE/HsQUCmoTNYrQQe3p6UEtdpZzPm6Jqb
V+Kv//Qs8kW7ChjiJkCouWtm81Bs5vS76HTtltxfjCMj+a33P6DD63gT8e8Cq7Oe
87DiornVVEId8nVWGGN6hmsvadNozApnzc/6YxlOLwQm8gnVC/6z2iZILJGnZ5Qe
sOAAzTBvrCNrE9fwnE9uAgKURiqNpi4OBv9VvvzyDDIQ0bMiyhsCpjzjI34axjZr
1RC46TuXryTMsJ7zY9sm/kG+y0h3JzYvtMF+n9Ci9/QTDyYuFFfT21voAUHVJ4JR
mZRYEeRrKEPP0hS9zmmyOSY6y5mN+UWHZonrYg1lKd912ayDFY46HMHW40v7m53j
geVq+DKWarMqpZi/aVRhUtpaa3w2zly+L1+gITEcxHwRzztQqk9iRKPI87oUNw46
1a1/w2VF2dDMoApoQ1lUIgDkCYa7Kr+usMBU/OqKVZCnHblHBqMS4JuRfT1I45cb
M3zgrrc0zSSLEKTHQutHG/Wu/wB7o6tR1tRJCeQ1HhGyLU0wt2l/Me8mNH29GueI
nRUciss1mJEr+OjqYv6ocX29FSi/J1wZdGw5K7uGVUOgsIiD03sxwsLFw+gIa8sK
Crtt969aj43TAhqHy3kFNX91T8ccdL96Epws7uut5j+5EQ6yCJLNh/8VHGacBY5/
CUlpGrR76Xh7onCacYiDIImrauvDfybd2iRekf49YWjRz9Hl/ZV8a0YyRqxDwzVz
+Y3BwiPGXB/Q5N9prSqvEt13lu1OdbuIZZylgxcPyrey4pihpdMObn6Csi0o9/sg
X4NntXgRN4fd/doAZR4LJ+IgybLPxL7hEI16NNREKMcpO8VkEH6rdh2VBzLSYlHc
uub30URELGheTZsygluX0EN3Wi/nTlv02qlo0vYzwCGfOfirqVPFUjOM28peE3pa
S9SLmhBlT8aPjY7Zmub5Jcfo3/B5ewmZV/M/SEBiyApw/DMdfj5HEiI2UvZ371Np
DXRjxCPxFpI7ckP+bhB1Od6+9kMesbzsVGfsjAqOtN6qQLfrGyQzasAg1XJDNfQL
/3hRh3a89VVnOpBEzGFVxdZ1wJJuj9jFVD4u4RuZ73iDCfBFIbMhb0+ODcw+I+b/
RFxKFQpOcog5ktPKhx/+s2EK+E/SGQAoU1oR4p9y7a6BnI7z7H1AmBeuD3DaLas6
IdWJ2Hv0nGzpWadO73b0Qf9jdlXiTRss6W9/6Us/ZWziBoH8XT6x0NL4H9ORY07Q
/jJcr0z37eWaDxPk3TtbGSfnOkuOqntlrUguOP7t9lXu//rNnGjUcjXPPSZi6gxG
pWeUX4leWyZbPzI5eIKSHggpxADVHStCQZHXSQ3kCNZmCznwuU1E5ibNMIpGPNJs
fW8oOmEKC+ecQwWNG0SH7Sx3Unq0lsrEScmtqfmWyBRpnCbytMlVbwtiLSEL99M2
KijlUFzuT5DK6vZbP1epDYNltpfIhDCJpo88/puQWVqeyQinDeouzCMNXqSES4lR
U9Z/Es6E2DFr4VfUEWfCQ6s2hCDwWhil+sO+yuppwIgcOUg8f+MtQklLWBAv3mLp
3bj9rC8T+E20ZmNvfAZbVrIQOj+7GXjtvUj/29V/8lbRXUijySa9CRz9k9p9WCu4
CKG8t+VX9E/Hnj7WT2HB0glILO3a2Curs705HgogG/0z6dJBC6rmpKvPJkfNpGHO
B8npmXpG1OYqD2QxcraemmIjm0j3PUnPcw367JorRiIH/2TRrkwRlxZ4u2OmZUFS
MMtQP8huVkFG7z89OqbHUKnWMK0ycAzbV9EOe9fjk17iufzEXjq6Fy2aPIKrDpxI
Kth/HWVdpOZONODh7GklGHj09r+yqaQuUXAfu/X0w4kjDF6SRMJ4PEaHZnWy3PvW
aHUqi8q4U51gx7QwoSts2HsgcqdHfcW9iP8fECT37Jwnt+BrNbAdOeNuAkZzg4fl
MVxWBY9vxBxcobFbK7IajMO3pIkwUAw3z4ZIeRxwcIxmTq/uwOEn29G8LnORVugu
SH6Qx886uPAhmRHPnycN/wlMV15fMuN6WQiW5Si7b0wlMSKCS5SM5l4VLZErhY4b
VBQXVv7Yr1mA2EGB83j68JPoUgMGVx+znjW26yu3p7NyXzPLXQvWJPXS6FPpBNZT
KtQ7W2yRdAxISSajhnQnKXQpbbJWWPcJvJX8OOe7S4sGesBdM5UMsPBS5DG+tUH7
2wcoRas0rCsdx2ttzVFFPhfZB1WnAST3AP3hRB5Qi3UGv96F1cS3GGAlyOTFxPoo
6b0pCleadCm0YJRRjcWXU0ytAkOB4O7XZpJrsJxYFrDz7ckvP1nLeWEGO81Ba0Vb
CVSVVqA6jWFai2Fl9n+c72ARzoaW9JIrcqTKJ/VJbGfIjuQZpqW4IiGhxgpSNHqK
1QOS1GtnbPL9rDUuTAJuxpOHIVfp+ytK5QCLVnxn4ex6Ze8HSifdp91XyrjQ+fNp
dpAkTFpnUpzjt0SR0WC68OxuvADOtnjyIPxRufW4WjfT638qjZpF8ncBiH9hdOgw
gLKHVQpB5psMHuXGwOZw6J1M0dQMCnAAlTFivrWWyMBg9MaMMIeiOQA+hhUkm73N
5+97KVxvMVi2gol17OmFxYKVlK29EFbRwFI8Sbf7u/Ihsuvrz2AAdbhE1fTF1yZ6
bMhSmxzflEAaxpjJz0JfH9Wz+zE4dPnRnkdJ2QsxdHJuDDlqOcb6phcAmbCnVmAx
j9uJcuaQ+L1mUOnv7zz/M5xQKg5JIqoyueeACVwhaOXHmhFdhcmTsQvXZi429hdU
8KJXeQd7L98FyBn13Hj2KyU+P52urG91jwS+sJi5qNylZpIFe9yoqw30gCfJnl9e
KuigglOjc6XFMKWe+5l0lF72CvlRtO5WxBeJR7xuofBbBsYmiPK41mgUGrKrIyya
lvOJqLs/9r9aHqpJxY/tEKcKORUDqS7DrgeE5sOPoBZgfRKnOh5hlMFIwJIqbJIW
ZQGDy5d4mpAWeAh1dv/smnXtZ1DFwrBGEzwxf1i4nuZPMyymgo6jjZN3UE6oESmg
MFlbTVtWnknAch8H7XMX6/lVFdt/FFVN4AQv1g97EqE0Wy12Kqiy2XWEHzI7yBpx
i/yQtvfMlK0UZJliceKBblh06gdY5vxkMj3mGrbv7Co5xo0ZB2HtWhUNtTvb//Y/
eig8cnEr4JlaF1OeH3cJODaXqOn060EMYDLt6WwgS8jgQsI3led0ZNavLTVOC87V
2TJST6i/k0DZfGstZnJ6GK001e0tN+/7InBsXwqWbb6C/8QIqozLLRoOctEr/H8M
UwYHtbuoNgCVPfWCFVXehDWBmMKI7krX7iPo78+0Q4E+wphawbdmG2cH6tt/oF6+
uLgrJITAdDCiqV6jLm2BJPVJzoB4n1GRraYFoVxTzaa4FJzD60RKc5SUQmR17/WB
A7ynEtur8zTELJR0MdfYlna98rNxp2xbTOoGR9Y7EpBT9Q0s51/HO3MMIHAJLw5f
Ka29e/SAL8e1P8al/d1rxwezpSXTql8/D2CqMltdffsDHliKGIhisM0Em9pRiE8z
BJweqaA8R6ASls1cNNvNROJzBcubqHIGaqyi6SFlPh51BYhqi67hVmLgV8dHkOid
tGFnuBsV8P7KQfgLdCXGjnY+c5cZY6RZP66fH+HW7590YKNXAEYnuDdXw25SMleK
vXh4wgzB/ojEJgAJ8fBLxhVCt7K5zX+WQYzAaK1CwAB5qP6vl6k73J0ClWgPMi26
liLXMxHyIPtI5mbGVsNEi0F6Ko+25MPrdClQJsUXGzE4OmmEeNGiq8rF2oBPUOeA
FIoXM+bFhPOGszsxNkl10oAyDai9N7h8AScm0NExkJLD+Nfaf+Gbzj2ZVMgAktrr
2yH2dmiq+GMccCxBvIYSXDGHinLOoiHboX94ttv0s0bQqdp2XRmgxQW2pBNrthad
dcce4DdcRtvNCgWM/ViVKjRTVBEX/c350tUmGj1VbCdHP9JCYYK7Dd8fInl52bqH
oOlGHDT4slNCHNdL+jLEx+f4rEiQ2VSe2C851/nU5WgRhgxbRHAMA2u7gpo66VyB
q7SrMNyJTgoyh1aXyHfvgHjqBIXS+RJHDLLNuyLWn009WXcCwHaaYWdCcf/3nZC4
RLf+TeKygRuFJm5hDqDLpujXYgOcmQJmeWwcRj1zqDHOnVkWfzxKVtTpuiiD5yWD
5de044QdBJbYGhwOOyGGiat4aN7Z2f7WGf9iS7nV4CumhbQs+9fiSEB3BLrtLcS/
0rZoZNaY3GwRgTOHwXbBnAetQfITTntsOWBM1x8e5ij63VGi0cF6oxCwaLuUmDE9
fBdrRIhv3fJWCgENRN6misQeECEwmwo6uMhlYOoookj5YgzfUOTqfx0VS6h7PKN0
Hgp85lN6lSd3RFCiWErCD33MZ6Uw8V4hWbUEQ/H+W5S82Q0REJLbTa9LK3lvuUh0
UxCmIgd8LZldqllScvCmPR26Sec5pgjeA9ISqZ53Mnae62Qy+xSMGKZMcPf3BZ51
At3e6yNCHKn5hwLnXCvaWF0C5d9InlSD3GQVfiFUe2K4L88Y8oPZv2rvcrCT5YOe
S85G2ywO6tiE3DfmK7iMZvoLIFHW4I2kZEgbjg4MSRCWiDwYChdoeiAkhVrLorvX
W2ww8OkbFpOkxO4BMPacyf7LSk0fIRB/Yrjt+ONZODcBWWfBJwEZC3tKgX0Dn7W+
ipKh1b+9JjWj7xe9Aol1DeJexpgWwvMcGFpOwBazDZh3Ys6rxnhsJ7IpTqZmTxeD
iI0m8d9URqxCl6LW/Wu8gglPX3Rp1BIbnusm8guyzXgghLqdW0Pki32rvMJVHwom
OAMtDQJQyXEZT77m60SWu0npcPuoMGU3DnECdKKq7gSu+H3wS3CZG1mnKm2LPaR3
pztY/5yMwk3zKbKpxKTa91cjSLQdH8Blz72BqfMsLOm5cRtP/vlqJU4gsRzEThTy
4jqUDGyunprMUCA5ba6M+mB0fQsty/KGrl30TXj1r3QMJ+I4I756a0b46JkelXm/
0MsW2ZDn8VmKtlujrpvpaGyoDoRysO+IczNb24971+UmXrAOxI87KCPqmIxrgD9h
LPK72X2Pq9yPFkCgS/s7IgYdVjaHOwJKEp3PH9i+VpAFgfnQmGxYfMxccT66/JtS
RIlHue+BmgRqTu0uVow4tY4Hz0u3BeKPihTtUL3wVGxVYVs2QnPixRs10/C5juE1
aIpZSEWt5OpNhhLXoPcA/XqbVznFQ+HXjBHKMRPvxv4pE9tNUsbnEEr2Fr0o87bB
xh0LXoajSEm/WcifvDyq8uggsmVV7kZAGIbOFKaT1k8nFbhQx/6DjVjxKtwq8RyE
Bs8uhEKOL7XqnLXqbFF4z7LpgEV8/zCAr9/0qsfa7d9RYWtbfJ1GupwbccL/ZSY/
erO0a7MNBg0HdZYhNunW9chgsJgIACfs/2aT65P2Uo5+Mr6NkmOiu3uw4BcmpdbP
2IZVJiV1jYAXGnbd2PJOGp/zpm8MR0DxnaGxEj+RbEIK0eLtYn6aXnvLLvTIjwn2
FKnbiuFisXUwx4Jz0qyD5Qe8FIfSEJNTE1XjE3Q2APahx+FKMXF/zP/Tr8Sm83HE
9r5tcZAtzoAV6yVC6KRV8YQYzeeGywZEgoi8o4PHZ5Nf0YTpZs0orvrzT8qzoMFZ
plyr+09zGbS90Oedz9Y/NsoPGhYtbhEDBm9QJDZoyKsvKigdzL0zIwLjy6g+rKSR
h5wwSqOHoQje/pKLoniWKtshHK0a19a4u4K/tVV4GsFq5qnrBCT9G8sgmZaagPpV
LOlDqtnDHyJzFDGlwXCfzBAXZMuadE5D+ElTTNSBJfwyiIAH+yo7p/Lc32WIt6qx
I37XADhfhtP+BpAT21/yGfkLd+bQMy+8nuvd1FhUWs2SyWli9ftCxVpiDp0zKh21
qnD+tVSop9Mta1ZPWCkENatPMrF8Sn9uzHqgOV4fZWqt1hhgTkdQ9UuMm6qRfzvu
KhY2BiAKrnpA16Xw+mOYQv+tWUyZAsXmfmOZ3am39tCbh/tNi+/zJEm68LXWhfoP
Kh0Mn8p38ZgUdOCpty1Ch8u09ESK0rK60v+evIkNG/byQ8TQEoglBKUd+vFRFy7p
V8h3Svwe1YW3zbr0YmUC6l06ScwSRE/3oEkt8oIuaQLN+PjCJ2qN4wk4yslzFTsO
ZAYndv7A2sjeJFdqHg0PVd2TUOeZtP7TjRFXqg/twKEPB0955BLU7IxBQa9+Yjc7
RzwzPdUhrb1km7UMRRh+Rdxun8lztEOkaNQRuH6hK+yzGQAqnCsaYyXCgoccLUvc
1Y6LnU4vdKa5O5PapD7fEpaAhoBD1ggoO4CYV2+OelM7cPYo9djtbtm7DDA7+KbH
2jzeAIiXp38Wvw5BrvkWqvs9grhNtS3Ft1QtSGQW8y01wLC1SYzyvTRJg3KZKcY7
JQnE1+gbv5Cvi69w/XAg3pSftdsMlex/+r/LL52MgFrjY4bYema4/2VPKx27ARVc
dLCizPJuokf/dNH4VOAWJ+nkR7nI8y3PxM5NdxaJCR9iyuguwWZXrrmfsGNqWWYf
yotyYtdNf0ut0cwxVEFV3lGUxTrgYnhV7X9YEF6KkFDiA/V0kwfz9fP1bDo+zh8K
PkjUQ5PzBNIrqgGxkHx/cYmk8DvM9Ap7OHACYSD1HVK/wJIhVnwSiju8qIcip12p
g2IiJWV1XlZuLE3fFpb0wwcfoVkj5BuqkNwJEphes4gUUH/yR8V5YZ33uwz3RrfQ
viDgMLGHNF/5taLOTTar0LtwDBVsswgpqusqviTYB9fJC2uqnBlyu8FczOGts9tt
md68aRRfqIMGfuijMGNoHduWJc6n5rFdXRqdvj1Tz3yxNF2CaedCmylhzeuHGssS
9gJDJakQkZEDfIycYfsxvWQ2NoY0UeYfVvaaCb+IGg9dVJn/2Qr7qhN2KBfRy9WG
RZ6JqGYF0r/u1807aiaNtwCsoVYCfgbm7PosEEuaajeo6PyrzJ4PRJ0orHKekf+a
CD+A1ijzJTBbINujn+ggAw0wySooJZYKJLIQg8GLSFsBcLTIUnjJd9RX2y46aMPj
PEJc/lIFiiC8q7+R2lp46i7CLDEpyfdpIkCYak7O7RpJXMHJ3zfhRMM8UW8TZUYp
8cBm8HaNx873/H5RluonAPk9/gE10WzhEVeVGXXcQ7NJPa5R6/szdy7LfXQAfrcf
k+wnW9v9EbZsbEGUKZokXwASpnmymwJQEVGQyodNtXO9QlpXic6MPDN2p+oDcQvk
aiuSSU9Iz57HHSk9Q+fXdOc8bHJM1viZAjNqzPNYyuMFmHsPEhxMGGTqnrmtuZDI
kkeeeWaoIGAzJ2olA9Vsr8Lao1K/xsM2kR7tq1zkJFYfqW7NZEV/jFjMh1/s1Smr
UzoQIeOvMDIKKRGVW9BrMaql4EjdItqqoGfeGV7/8E9xIuQhqlQNo5ODWMcQ1gjy
JEHNGoKDWjmmMlbyQGe/BVJh7KfVbDk4MVMmR/d6K3E7ewKcVAedc96s+TEDfGZy
b592yfCjy3j3ROX6h1u1Lw4b34Y4M+pMh7X8anwVG+WshZf4vgsxf7g1m498O5sN
295SRq+/DWlo7uw6tD3V5ilpUowFk8DepPbfK9N5Xml/woBIRJa5NxX6o/0d4FCL
TSMIlqfVoUDB5dhcK6noJR25ayQ+YVjIOwLbIiF+qXUj5kJYqrIo0IrMOTSl2xAX
BEj0LuCyB8Z4N+vsQxav+H8GPBCwZHQnXzPGk63JL6pRWOCW74m8YIR5RtksK3Vp
hy8uXcRpVGRn/yR9/462p8oK38PX3vUjUndyITVazretkRSm6Vvojxcf0NkwOwDO
/IcM+O7/2VclHnWtIPIDB3CMJ5RYNFA/jVpqBqIPuXXAf9l4sXf9R0PYayMJGCbA
+guubbvw0SCY6iG5DWzJkd92qX9vfGPBFP3dBhkc23evIUJKJm4FliZO/aXqjFXm
L47Fd2ZB61q+ssi+BXVzTJJh1z9oDld/9x9UhrjaAebskahefWkZFh9iKpHNdtL/
eZkKaWhW/tMBt4owJHvDaHrqTwFM4gXCgS8WvbzfStSyvEkL/4JyQXor9bkD8Mqv
khtMVF6mUU3f5WNBn8ZKgpLB12Q+Wz+quGMwiRlUa5+rdo2a5P0SYc7mOi9VI0Sp
9tCtjrZHVGrfdT1g8fQ4BuXATfS/1YYeZD3at+XaeQL8+GrU3Jj+c4vg5l0U1WBc
Q6SEGaYZrmEK3TTS7HFKoZklOiCtkr1Kwmv4379FnuHbfjsds+M7N6BecNmN1fB6
u7FV36kyg0qEHXS55OaD8DD+jojAJ9clIMwM/tr5SVHGRg2YIqJdiclJxpOVUFZ4
WXFbnnVvyVUF/4xLzOtaI1fo4UkM/4zBu5IU8WkYOo08qXqSFi0byJADTa0jH7c9
Luad1nNXutYA+I4XTGhinyb4J+TLkTIn5V32fD6S2naHmw9HdBaR0bDDW44as+x0
ytZTg/tmRI0hJtsPCTELpZdnEFdmTM+s2oc6vQKJgzjyOmzEaHWOUzChGBpzQ8Nw
u2YwyffUkik1tbBvepewrnDptoKDq7SeXLrEclSoFr4qvmtZgTe9z96YspgIAfcy
JjhHM/7lSuuuJP+ZvJOkaujc3pZC64KtMOWlUIv6Cv089ToH04z/SY1Y+blDud+T
wrS0905n891sWJr4+DI0YIeOz7fQNwcTUGewdM9VgHiaIQjtnt4LffMYNj/ND+iB
vn8hFZRfW58hUliKmxNky9ZcNpCHYZTZYx8KruWDsA0Om0pt9skpCGUstxDVTsGm
Y19ut6uY3Y8YpqzPrNbZvkjEr7PeOJHN9LaM1Oauw/j/PRyi+ECcdUkVyPe59jOT
kfGgO2o7ddFk+gGjTo3VyW+pRFpi+d29skJxFRapCKLA2Fo/7Hw8xSHuCHK0X2CC
9FZAaKe52aKjKoRLfmpwrUB+DGQOm9awe47LnZbSh7Wu25TbytzxoruM7LGS2iSh
Dy+km1u4zFMz/5GfcpLvCb3UESEHsBnB5FMixRwmONS8Vu/A5YLY5702vLvhyhA0
wkj7YhBJgwK64LYVOTuq3bIfSJK5HHbgtYqcsUryvNbApV2Sv4kodp/6gTnWP3v4
ZZryHpR1WwD1wxwcaHZaAbQpguL100x7E3AQyDpwbLju2Ia0So1pHFV1/BC5azU6
N+nf2ybpNHcwZtArPZC1l+O6qZAhGaaSg46G+zE8Xrs+a7OoDqGerwpkklEY03Y1
k1Laj0cRWURc/Fj/8RZNaZShDJNZhBleAiNCozk23qSiZlxzBta0IeWEPBiOPQLT
fTV3x1Km96Nge0l6nJ02RZZvx8NRRC9dOUnZJ1Y17cTY1+6cCSyALX57dOeFULGj
jdmTYlt+gXuoIWUQf+vPDKO15gW+vqx5ywOD0ltmPe9lvL9V4I7i4s2LzTrmCJEE
NlUnXeljsoS7qNXz/mQCPJ0Rnf4tzKsmQHOucnsSJOsP/qnINuuo53inLcWpWzfE
1cwgJnkwTR2+mGg/9lukc0MvlkNIQLQ7Q4x9NaOCabOr6FZ36Y7zdxvzQ9KGlErm
eKJsWD5twzBF7/jEHcQmtq9RCntO72LEicrvudyJDLefXcc+R2R/YTYPjbElJNSG
q2sVrGb1Ukrb9OQvzN4HLF8NwMVzTxIRqwHnfG5pnEd5ZXDbI6Vvwt1eq0Bdq/Ur
pqUKinQul2dOsmfqved7slaVCuXDsja5r04Mif9d66TlaaK/8nOwXEG7IfPZ4JPz
u2bPdu20/vDPL9UDlbjBsTyCMtWx6avZOt/Up9O4bCmWx6kC2IrvdQW5qlxi252n
GmCVYCitkdyU6HzxbUFYnw4jrfArB6HTQAJrdy/YMVH60syuixUtONCjEmEXHRau
OChJlwiPIVJM7yT2M469GLbO9sL3rWafEGfFqoTNOj0DlCOnr5v+EuR4Lswn5Tui
LixE9+Hbt9HUjnkJM9uzNmMd+iz8eJORUzLFH44Tz8+t8IYvpsgMQwU9/GueXUGF
Y6OZjhzzU7ZcScIwmMFT5jF4B3QvqAidrb353O0Rt1ZwdbjqtTJJnjRO2gXFBHcA
XuRgHT8wmTEwUQ9X0xcvm7QKkSh8RdyeSvrVbe3pCN6siH5mJInEV/xiJn/TysHM
xwDEDdg0rXWECiHid70Fal6XDlFsQDE0dGhY8udSt+SLBtnh/HDwN7MXOp2z/1Ef
2TExMoSZMp3Tz+DysTugTiFg+jtugYI3iteSvsXtfOMZNR59N6da4PKXwxRra5o6
0vvmz811xg/BuYsMfW/acRQVCgwa4Des446YOGhNxA9VuxZUh20agfMNP1spy+vV
nAEMers4RsJIqSc26F9dKG/tvSY9VjI+5G04MCqUqXOI+quaHNGp7QFh8HYSJSaa
1uq6QXeIoSV+AsZ/K9yLXAw4Rb7+h7NIKOBfyEbjEDQLeTMGgsEszhK3KLVGONSY
z0kF+eMwCOF2onEcc85imIB5Hfl1T8jL1Udv5N01ACwGsHZRXnWvOqsokyKHz9iN
vpIS+T5onZv3kUx/uI8ta+dHbL6EDh2ffh2+WJ2/mL+umqjvnBakssGuzBPLs7xk
7r+qth+mnkbC9pzwJVX5q7CHH6V5VYcAff2Z8hqSm1c4xdi2vC5sPDoxhE154i7v
8HPJjAYKk927evrMflFbEwWNzvhOkoEz0qNi89IbEEJxzeq42ptKcmG6SRMGkNXp
wKUxHIrL0Lb2lYKbYsg5t0QoityKxCwQVAYssPTAZdoGf0wtrCsq0WHwHKD/H8Vf
8LNG9VZqLVKAFPjBfOcHDrpZCXt17TB+hP/z4AsWtKNZrhR5X/cyoFftFnAXljPc
dzztN7iR5nLl0ysCTBTvXr3bVBn0Cpq6go8uhiGUDW852jrkm/0YxUqmBTxRadxr
ySVqUi15k+M+5Asg6X/3STwBs/DRZMr+84wj3at1IuyzWKEVmua5UhLd5RkB2+Yw
2+L4QhReNgQsOfmDQ0bFd+00pzaxxiKTOcrEp6jgmBh0xzFBEJiB1wOtYab4Xv/a
MC/5BrYOulLh3VPbOU93qMNXVJsqhfE1aPVGLPlSvSctcORgWeOWcTknDbwXZfud
93STMQ+PoP4x7i+684QFmEnXvKMhRBWJ1806XojQ9fbTaAauOpukdNXkmMyKgyrQ
VO9G7K87JzpfAHasIJLyVkdTvNpM5eMCDIlWEeeiqhz3zEPeieocbElfSInLLsFi
TaV6i5tmJMxrKEs7xTT+1FQZ5TeGQjD0fpA54McvTbzbOZ/3KX7bNdqSd10O43yr
YpF1cAb1nPstMf5HLAi+Bz8yR7LTA0HAS0tA9ySI83zv1qrXZsPoU9cD6EXMnkuo
vTU4Ys10+keftsq/IG2Xy4gRIqgupnBFXvH6reQ7cOoVkK7dQt/nlM3G3XK5esm2
yKdxg77dGluTuwjOPRByeif3ljY67qe3i1p8dIzdYCCZkgeygQ2HT32MZmYnDEY2
8KSozDcd0oHq1JkVVyVVO9qxCSHfqtkZclY92X5W3DYACTQ1+NGcGZk7DnWhkK/4
uRmcdE0K8ajAlwlcLfsB3fJHc93nKVQRXUNNVfWk3qlW2QQUar4xJV6TSgDYZlwg
90sGA0ot0InXlg/AUyK2USi5l31gxnWoOTMjZpBLl3Ij6kSOnXbhm8T6kmF1TMka
kdU4V19AveHtN0XCKh3fAX062TjHIOyWNpaMz3zRl9A0nloZdlc61/V4Nm8FlA6D
2rosbpZmC8bI30S8UqsnckOUV5Dvq4EUoS1VrnJZm5mRAFEeKlcil3MNq7fDk1dD
HhrzvAL/FcTz9gDZXlqTmi83g1s8up4mO40smtd7Vtj07Pg8OoaHtqyW0HA7flir
R0kuDU1lcow3aX8epCwt8XEmUiyB9oSpWh8wIvZsCSFql/saqQ+xWg9hxjDotWRc
ed7+QlcGFM0DZLWA7AYz41lkkcmPslE50d0WM7VB4GlMhJXbz+7Jgv9Ylv/NORHi
CA8y/BTlxfqswmkWVOxlqkA34hS/iHmv8g330nckRgwN2wMCQUz4wNkwGOFih6Ot
J2Q+pICYJOlU50wW1nt2iQmOSEmehE6x11sbirIVGQyztay5oejekNN5UzIQCyHV
Vqk6HzHj4gcb5+KtipL/PvWJxy4ajTl/Y5tUj9/xA8WH4AacK18+Ws55cFgG2gJ3
j0xvdkAviReVZOo6hUXP2rAkfiSTdPnFQd3dr6+3wRK5mPY4A+n0zAj/xbCyWUwb
9Qm3B1mlBNgyYm6QcLQ/JrJ+RnFyWwcEFTMDmqJ5nAwkNZ0JW1TkOfUbB/dNuYEM
2sjujVhleRy1MJ41f+/pb/CUzvKnwo+vVMUuNrW63XFVb2lb1sucycwtryz4tsjh
yBQWX+hQef1r5SV/+Jm91BcyQrkxeYgzIcDAo6pmYHEjgzlZ2cmbJW1aHZHACFzw
Z9D624+h3EFffI1/pQjQ6ThGu4oTpKgQRFhaHLhQEV+aTyXHXm0ou7LGisKoX5CS
A1hDy5mTW7XQ700ic0TZcW17j09yH/jEBWyzD9k38ctCsCy11m16Q3aPEHlxQcN4
eLDn/SkBIRYXjtV9Xgkzzr8gLBfvqABolmkKAWM96N1dyhpqXHtiZH5fu/yvfzRO
AGcrTO66SvirViJrKd96HQsyhKoAavm+QQMOWj+Yz5QitAaLK1NiwAO2ed5e3R/p
3XqkPXkDvu600imjWSDvV5J2d4MxS2H4schdEr9j7LsIqyzvtLyYaZtTX0hJE3h8
H4ighTfIVourprtr1DAZB8euvRZN3Agzb8Waf8BQfpAWOHn/ZsT4jSEK9CiJFRpR
+GQw6mXVl9pb5YOC03MjKvcRaPIy1z28PWtz7Nx4wZJiF9fWdKGEN8tp2fPFROFz
a0/mZHW+3shV5b/h+9qRasea0eqCVrG1CUXJCJN1GMHb3avDsSCirySf+H+Stxzp
p2crBx+i72FBDFj9jpMAPKDyjvgRRn/ft91ubNjYfcH4A7nxsPOH9+DNrddMZPSh
vS/kxpUW5jR0+E4wIiR5p/SmM3zvFD3XgzWzunJDBir0SuaAM5X5JmmUqDqR8M+P
yBNicrHYlvKGUZOqh50BRLBrWyqDqQxEiz0n8/c1ysZrUim+XTmgZ9RgsWuw1JaZ
b/EL7dcunPW31EMChhjBsLHXYoCp34TWNpxI8CoFSgrryr1MxMXlO85u9OIC/K6V
mBqAoSaiqqDj/OeRo8G8tdmfcGE+8VHj4JozciL9T3prI0EKirHEaG8Q2tLF3o+G
OpU/LpDhN/v13NfyiVOd2XVwg/GA4fCDK/ONRqnjkZvLEnZMC7BoMyc+0R22Aioz
+A6kNqNGksW4Fn1CWGOtrjExPHI3U9GKFEKtulKHGbmnds7H9dEUB4NLvoYqNI9d
rjk4t9nucLl7GOroADXZ1DaGoELTOJBLTSwq9h5qVpQlHrHx81d7wtxza4BNjeic
J0uGX5Bx76FJaN7aiczZ8tvg3W1pjWcdWuhT8VidLZGipJXyjD3o03LVvmrtQ68a
4NzAs2NobyIO/fwQ3jNL9iGxr2Tpx6LWfKQkzCYB9kJLev2bmRiqoGmPXiNHf+pB
U9+EN7qylbGktbuO589qF3tXIAnzSUfNeN++oqP6yH9Do0YrpzQs13CC0jt53hXs
JMFHesZygq6P2bv3BeK4OZjqOU+cHVBpMJq8i2OCCs6SOYRhOv/qnKSp4Uo9V89O
si8tkCnwH3grpHQofqlsa4WMaDKFv+M36s23o+eZ3ZIehGvPlM5nzt8R2FYIIyYQ
eNJyyyUyjcPUT3EM43fCQ/C9jMHYpBC9uIew/YaDxi5t+nK/73Dvwi4K9SsjWS6J
3NurGsErIwGHnaJBSrwnR3Lv3prGNNtq+rRxPpzcGJ1w62QlRog/q0E4Rnku0auF
3gDVJ1HVO18YcxxpwrOXTIFaxUQhyId9x5Dcpf4eeogalqdeM+i0kzC9VDUJJ+FS
JWfeiqHTZi27QVLrNDGzKflrlCIt5HcIybHbrTEbvnvhn9yVeAZ+nz6EG7CDJb7L
pRFhoNPuMtKTR04PcwPcpRg1zpHaCyNFdgiTz7EmiqqCLwpDLYSzxPCxi+X/Erc8
emaMLL1gPTw6Yt1sL+eZSTXxtlgOALDJVlazMQ+eVqA3CJkPPUk5LWjFbZMEPzlr
09XKmHo5iItWVYuVXyY2lM2uv5ppUs7Jr4vUXRcNOb+QjLpfB8CfLg1NcKIAai9C
HlDIa7FTDgvw1I7b9HwVCA4zQdCisTXVeom4SIVbzeKgnbl6SaU9rgG39y6UDbV+
WikZTd0NpFXALsp8XCdWyTGpEQR3dbU7P31qjF+bvIjjwoGEE+g0mtlg223rj3BT
Vtd2ftwWVzbESLtf2Dteerqh8BHttQCkN74p7gnpgiXxM7TJ1QcfB2ZdzFEDI+VH
PXM/jcoAZBDrK9/N7T8nDsSHBHaDvK7kUC5ipIzyge4urUcdljAbPXubmoulPSVh
augh+BSYLo/QyTzgeqDLi5Ax+a9anJYvJPcV9hZKnQjoLG1rHdD/6rv0GoXGy+sf
OWMatYMgKeFAXW1K0geUj2Ae3K4Nzh/a5SHeq1rV9rvb8OTtZTG5hY/rQUzYMnZm
8JGTQatvNsfu0B3kplmD8w3oAIhDRLSB41QfLIChVT2OpSqUEnkS48Kwci3Cdzwg
KTwr2JLB1x886eYCA9jmRLDeVNV7IMGUs60lwoUW13u3MJL8LP6m+REMgnBvaNym
TfOClusLMYThDQCQ90hzxu3CAC+DEy20dbqyEmsWuIJ2PJgWIleStIyRlOaPSEU2
O7b6pRqVGjZjI1LAkEz+XR2xTVw+euKo+OnaDJFXF/8YJH0W//G9O7MZjOltsZIX
bG2Px1v9zIEIvSLiKnbJZ3l03EAEFmAvpajo7cAuENBlSCV+t1xgUcaIYpvUEA3B
25EICsbDuAheB6B88hK+XMdhR7xzxPnsXv7DR0vY+Qfur2uq0x7ZGmHIKkVO6Ddm
5LALTURYGWjZjWOZ/t2/TGsOxKv8OYy+K1+M3VUOeK4CWmpSN81Kj/9qr9U9aKDz
mpDF1AdtlJoa4B1p7SVjQz4dJWe5A0hxinDpevVuo4+1GDq5XTmg62SWVb7+7+B7
uV7/MAUsKTAfIlDzqtFfc6OLDtqXXpEWYVcxCh/odhyWNgDWFERXKFXh6ddu90Xk
0RyKd5mIpO3gB9l1d/6Aq1XV+Ofnsix9ME+ork8GNn3E1EG2Ycr50dOePPWjXtEd
HLgMNShJiBnFQp6crdNsU5UFtTcK4zZEG52D4kPQyHdC2sl/Fq2bgS7OLL+auiz3
ZRf4smSTiikKrx70T6KL76esdmiUkS5huaD+z5v9k7hkw/h/mXH0+Z20D3+JGKUT
ZlH0ac43N3BF9kbp/DvcKkkLuB+vA5V8BZq/U7/QkdOnTjJ0z1WNwWCIAOroHzD/
gKsKQDRbO54z9KVSIsHMLfoswxEIzwGVdUDgBCz42ZuroP2GRUrEU/FK2Ecou0jN
RxYhPFZH6ZEx82aSnwNaoh+MdpvvNGNPG3o+jGtfm5SVyrE3a/JY2EQ5HM+gkt/B
PxALVBOXIf9iXlejXMox4X2xnWRmwnxfI03JFhhO2fQsYCeIvnA07ubGc/w4ZPW6
nBIBUkgkwnrJSXGHr6qqm8EMfhG1vZe87Yb3TfQI2Demon/sZ8qFO8QUqk2TjnHA
luxYZPlMv54Lg+hSs+koxHl3n6MjYXGf7yZzIqzcwHwyW0xOcUphQXKXrTcSQhWl
sthvMGx53CIFmH626HsNOaLukOgstvxkKz00FgPUa7fe0RgG107x0+PrTA50yV3q
8Y8Ypxz7NhWO+wOiWwlflhQsZS0WcdvDYU7wH0jv4jYjHlT4fHOGjsoezEwM1Bqi
jfTQFxPc1Y/yvmAAFOK5xX56/8D4KcxNcq2U1ZFPlgcBy/oAtAqViBIw6JLGz2+l
n9m2pM7Mld/a/rEi9pnWccV+2EAQTzIUyNddiBR/R5DXcZopCZeidKRMoWPO5Luc
nT/HLi1TJY2k5bKuSsBrqyb+lapWsb/3qcGGjP4AtX9rPvIqMPGpLV4Xd3/yPj80
o//2g7+GY5D9AxTeISaxnSDwR4Ydk0JHE/zVR7EkWqP1d4sNJPPUkSYSNtNBdam7
3fFoKXOEs+XVpVXLhE1WTTcKmN7q1hmb2MBLBZyT37BFYQ1m18/QhNjn7yDAU+Uq
GoG2iWqyiPAf0SricHbE8Wi9YrJpegQrvwG4hG950OHrhNg7mLmjlyjzaTiwwRRF
+QMPkyS6IseQLzWOVToERGXi142jBYLsdAPdVBC22WQTphK2oQAUKsH+Jugpktem
0X4/a3ZigQ6TAgdEsrVRJKRxLiFajojBdkmg6iDfSF8hkpwSQ/uKWm2jR3U8aKLy
5bioLQ1xTXwGvW/2m4dA27yJVtklxxl0PcvrM+ifH/pTWuOrrbYsvmLHxUiJlhe8
1NHDyKFC4vQsePliMaPR27YscLSSOd5OxSM6BMh1G+XfLCSirGE2mlwbCaWuh3Mo
ZAcTv6W0k1GW0t1ZASC5rSXJGzONczglNqEA45OZ3AhDl3l51c2loVs3ZsnRytsD
aHQdMrJ8+QAecw6kuDOJiRBX6EtsM8sYlM76CJHYr36xwoHWFWY1Cjw3XmlsgnIs
G7aiQ96DOxhjHi/DU4Ylrg2zzDBemmvlPiXVMHrehToDeLr8KdlYyqHqfZzueWkZ
oQ6LkTl5b6bGnvbn/HZ2gMXcuqpW0laSoejvbXKf+Pl6jiKBBQoR10H6HA/wz5sF
sYL+/gV4U/fJAsDHDWi8JFlyUoSAnPMY4qxh2ThJgobG1AdhCoie2K+jJyecafxc
ueK1eFUWfx8kZZsXyio6eYEs0T87uF5MtU4/lqGIexWacQLkN/s+DVTfKR/snvoi
R7I+nMdRiDArhSwzdA4ij8wRiynEbGgtweQFRHfNZp1HbHRsE8HygBu+GpGw1lsp
DEHUEpRHCLV/ShwiX9lBhxIrkyF0bLg0C2hIRKhpnU/648rwlQUU+fGI86eT7ciz
mdum5xl1S71mmgJ1iGzld8EoocQi2WU8HRbw9ug/CvbnodZmXSchFT2QwBrxTBhc
/x0yVAUPzNipt5MOr9/3ifpv9MxafuLk7eCuQN2BD8v+a8anhTSBn2LOu5lHIvz8
h3eZ1RgHl9kQx5ZDdpNM5lIs2pci7vys8ULsu3QP6XMGBhM3eueI7+gVI+FoUaZn
hS9YdAwf8bnpxWA/pnfnuNJt3O5ztuu0yX/wS2BpCegBfjL07LEF9k4jXD/SQdMQ
ahPHY8mm4dRHXCqEjmZSj25BhdXppsMaPI4Z7PZSy1VDPgBUfelfwBgUmi4ZoASt
9dTbp9pwBXyE6rwTb1o+I1dbXH8SbZ/DA73dBlXN/ZlFRDNBDwxXED439hNBLxql
3J/ZJp6XjYMLfgeGzUyLQ2kvjoPq2/Uz5TU1NHGB5Xe39RpZu6GPv12AUwUE85hz
rwla4Q616hITDwsb+1ZX+skESFmtvctFZXIAUjqXzMWvZwa7si3j0B6FhbKRJomQ
3dYvdj5EVvtu8HVVx4gFdTx++WaiHGxrfEVrF0d5I/cxqs8shgs2xZ8ur2pVQJSR
vBTyZt0450XfGeApk0F3nvLOIAbOARPlu3U2bwyG9Mz5Mn49cyYUbv3cHXkLn91x
rmf6caWokSUdjJTmSLL0slYXGeQ+YcvXyAQ45ETrmEk/f/lhoibrsHe/9ZXRgiVw
KzxKI6UA4i2aGdjtPS2R8nh+5wDAWZoDTTi98BMaB1s37mnYIAaaV/kXP7rF4UU5
0/KKurdaMVBLwswVr/lUgXxe9e/FoSNAM4VVhRFV9nqDHUv8lJJQCer4XWnxGBGA
aM9LvU/QQLLJvOxxczRt6yH+E1Q6cv2RxDcwKKRJUSnj4LfKzIPdWDWGI8jqiAtr
+asBhaf9lsVluzrV3LnzotIZksq15+U3LPVfd2F4vxpcg48a3tfa21hAC504C3cO
4/ZsKY6l/uLLNQZctK44qJjiSZ58Fp80FuuYc52cI8nldwFpPK0wh8A04O0pfllw
VyV5UI8bV6W6YOQvoeLI4SojSjZuOVTpNwGgK5pMSO+eSaUDjtonZz5bSp05/PFg
TTEOQsz2EOEzSgJWiREGlOfefKznWLcATpRYuTC88HV5fCQohYQaNikcB9aG7GoR
fuqA1CnL4dtr14iz/u0tOrHS3hB0uwDnIwxf5+DLBxNqC5P7nN0r6wmVO3oneOKN
a0hJQqC6rInQ6MamyDo+pxJoGH3Y+ZO7AR5gojvWQ+CDihIl9RD+RW5/ApqJE9fV
K8WxLB6wkKYaCEtG4w2krUYtoB9cgFH+xZkWLRxV8E5MjOGYUuKMxkTz4L/8Xikt
+YtpLIvOcIaKXacf2UerEFNgIcamhMie3ZTlTQ7iwniHh3vc3tD1U+evx3dWTxxG
W12MpOx+ihVlBjbG8fA0Zl2iw6rfN+Y0s8VRc1JeQS9W0qANUhQAxOqKn9oa8Zyj
XDEOvw/Q5Q9g/dSvG2lUHN+ChA9N1bQ5buzX2gfFRXkowAgjVi44L8YlnAjBQzYJ
mhDOrNzcJd4tdrWgK+2ygXYBu9any5SIUFJMvkXuF0KyPzePeZXng1l4i6t27vKX
Xm33d6UbMMVbt6j8Ql6uhFSsONRl3p1Gksy1p1qfIxzwo5BdGQrtupL+iRRCeNM8
bDZYHFV4Net8IJY+aHVf5NXHCVEbme0zPRmhepuHn+JCqFz6F3u1WCecMhRfqi8F
HzGmIH1pjGSIa2+wMjRtraFuIcglo1+qdhqjeUM7iKoEUZzK/77wl0jX9bGvTnn0
BJWTVwZDe5ntMwGFrN27UhHUMtqPBl2zyxjV5tSrzcFWAr27WQUQS6bo0UWSKVwD
wJTmPt/jJ3p7YHljtFsx9IzHey4sC+M4KCWotj+ecWfNwyl0kY8zN1rBVHfKdyT2
5YZgbif4XDnem8EnogU13LAvDd3dLo8DQLqfCiX1k8m0oBr1IugTJ2wRtZHY/5JN
mveqWVn2VRGRGqi6rDDEYLNRNueqBuUR5O90zwFybg92cWI85zl81iX3HrzVqK0e
cpv97CGqFx62Y0Jj3EOubsb38ZPuH67iaX1nwu7B+dWVT0yB7+FJx3xtexOCu1jn
mwhufj5GYZl7AITbr6vBouyjFDY5WnRbVmCzDCDedySI1rJUjl2ia6Arj7QfMg5A
HJiaugkCcLvzwThacv79/r55QsxqQWVkanCUL+/MAZdRM5KfN3r2S1LlG5iVR2Ir
bWsY8ulkcEBHtcNcVC5izAOdGGgk+sA6fO+zIExbxBi9XRT/uHgInsiY4Bfn9qLV
xyo+I0bR55CYKiCLFeMaSXUWkHJsrQlS3pWzmiTqMmeZHEZksXOViHJKGHsznJ5S
uojQUT4TXUKz61H6295y1mU7YyJZkm9KZuD2Vk0pMCC9aN/Ber8lcP+KSji3J4EE
IDEu5lYPxFm+x4BqMYkFadne8/RivOwNK25AG5Zwc7gpX0C6PfMFyWxna0bfQwvy
P8IGUWF82rIh/MfLzvTOOOf7jN+kbrp9w8q8fPy76aH6bMDgBLKoVIuHt5bUMUIA
ZeDcNa5WXA7iLFgFrN3FejkIcWEUULD2a/hzAW64s8GLQWyit1dU0sj4b5gl+LNw
JeODQVbnUMn3FWniQAwp1ue2q8NSRgZZReP+mWla/5txNYt1h+vjsl+k8DoE9Rzb
wpzbFnYGODbBV3DPVLMTtZX4DfNKOshzflV5Y1SISzkaUovhoNM1/KUCNAiX4uhK
IAF/IR3ZfS7V4+CsSxbY9LJKdA+qIDvqPBMYE/bQwfEKr7ktBpxuAnu46/6Q/AsH
2YrX+dkswwngIaFDx3sWB8L6+IfVFCpuY0xSf6Wm94aUqc5gSOT6HrcwxQZLGUiP
EtDiHTh5VKyL72giWt1TdjBTRChGD14Ko2SohRFSzdowNnPq08YhIJAq+ruTeDcv
23RW9uBmlOo8jHeFdgej2a1ZbeP+PJeQ69wgRCBq7QKSMlJd0sdJnaYel+8O6/2Z
o9gtVpz/8rMUTM+eG//9J2T2cq2LRtlRSZ9msccvX8VyZVKSLeku8atWv036nwXp
fxG/nC3Rn5I/kWEZj4ztrx79oq2B1O9D/thE+lqo90xNVKQz0VA42YZuEsjkl88n
UiIB2ST5QnTD4FEKa/Yssf2Dnd3KjuZ8rxMmJ7G/ZznqoCthXz+MWaCOdN1Eaqlb
1aOtv8Y8P2agtAdF0Zf6RKexpIfFXFRvh0nypxqDa90yl/KNYHV1eJgXwFry6Ugu
UMIlnqtVkZsMfybhwudh3li1S23V6j1mKHfHELS5W7ggUZ/OibcSbpl4lKpsLrky
HtwDjQea8HyxoZ3xiOfPfaaXK2AhTlZfY2f5aHzdGAu09SYS5qkSb+RQPybxM3LR
0BfxFjpdpzAZS7wF0dYM5/FPSjQVeLUV3qJs4A6mVGnxC7YzLcvChyR35qMhU2X9
NoAhgSb8yvsoYfPKQl9NJIXr+GNTK1698eePXtNGb2fIfc8NYftiRhoLEaLbQUQC
MDoK+aEmZm6oQRogpa1t7Zwuju0Y9Xx2XiTsQZe8AVj/06Tk97cERLSOorIsDRQe
5/ffip5cOs7w6RN5e/4AozqZmstubuVWUWtttnvesItXcwgYxZCQqVSTVekmOtUE
CxKns1u6ZK8w+JkBzdaChzlZPXotU+8458KI1JUVYXirRfxz+EkYBTbUBIIvofd5
Ptb9fpetAGnocabkojJzqhfErzGWxHHjP4ZpMV5jAQCGp0V0ENuxk/HIOsxDGEqa
gFisAUPmsiucYQFl5l5SSAmqIWtaAHSB4r1buRl5kkuU21A37YhzvMWn0V3SZgxU
A/qfs9oQV3ZQppNGMegYuz6lkLtDpKF4u0PnXwKanEEDfn3xypCRyRJwp516SJJE
Pn+FWTlDUh7GIsLYFqczjEq7N06TeqmRKnJKHeDv73HPWpnS2GuzxLUWelQvJrf4
6t7bO5WnpWK8hEe0Lo0lap8g8kxh0oNQ0EFs9lcv4MK9t0fiD84zkDTsTAeczBZA
4tNUSy+jBDCBmPn9wFmFeRoJIEY4EILTCQZGupPNDn//YB2UxBoWMB3PFPFszc0I
c16Nv2xs0kNDg5aOR5prjW/uuCmV1cxiedL7LKGE31xH1+YE3Ksz/wL2fbsalehD
fNv0CuCqmtKlYLZmK7qUZfnerrbGwA7SYhzDABwzKbsjHA9JQu9E5V9cxOKCC4Y6
GSQr0CjuutMRMx2T7suTRFXEfUXh/Gyn/5XpYmSz85MRKKccIUP1Mh4aNO5Dc5AJ
8tSMEn5RCH1L057/QbTQwDZIO4Y4VhoW8JAap69EHgo8H3f83nxGnchW2eDNSmx4
SAMNTuHmr/KcFWD7IcThOYI2BM+EK8TC1qMNCMFzkhPLdOzMPKDOUIMiOvqyQ7w/
LulDgCdXmxVeSCgD2Y1C0Y5w0T1/zapyjypqahXYyA6oNoixcuD4mONg6KZ8Vfup
hwAsFLJcxNQQH1V3GRVDh2GC8Ya4WEVttlS66YM1vxGHH6ykzACtJv1d0R86zca9
6RY02wQ2+1VBC7bCJ3Yk7/ByNX9uLMKXZr45A4eucCx4OPTx936JbDf/tFCmx2KG
rLxAWTIIVSN61NaTdZwZULfJwlGP0MfMI5xuYZZkCfFWKXIFqMser9zINym8bhHD
LN/I7Xl79ucYlIy78LFFaxaR3d5c5zjk5exTl6wt63vH/m8NVahQyifX9Kq1U+K4
8W3uDOaKp2hM32lSPEpxCtsKMHic1DQKRQrjbnMhV7tCSY9qqWllFxhlD8MmjCJJ
45kfDqBz8M8cR+41EsUPItrxt9WE2MsH+vTIAJy8+mEugjFnwyKdzqSntmdU7EdA
z08u9PKdK+S2kj7O85bTkKCRKF+gQV/S5nkrECtCDoVKzc7uDrsDZLWye/Cepl3S
sczT0yeAaAuWvLq3njMYcRizFWsiEIuFITtQv3hUBGKbbiOHjrQ/kglWDf9oPqY0
eIimIK+CZfQ1osPeg+7jT1w2/RAmvO8fB9N0QliXUMzs31bbiIxgkKYrWIVu+rDv
GkEunmyiLhL6l3G1Hm0vT94Ze/7l69HjhT6ChmM+c7fHZXWXdzap4vKDG86Ikohl
YokchovZrhx4Pq5kxPdGAxUHoNh6NJz+IeMHmhPdGnIR9LhO4i048VU3koXbMdpg
fSpBCrgiCAMfc16H84eOf4Qv11mpLV6usaCHTsxMBGeAr57U2L4jS8O997xPuJ1n
Q87ZMLJS4AVGZmTVSZyP+YQTRh7SfYh7xuOhAc4w89GhhkrTWo61RL6IX8miN9mO
UdQfRJgYEsU4PRMjxmHKyfTLwAnm6zUYVQrq5DP1hT6fJY11ASlfypxf0laDOvNz
qY0hM/b/egXiJDhD2n/8ji0QtijmWmWx9pOJva/OhLUo4quIFq1NRiJjOW9MNDnz
nSGzqla/srGDtvYdjTfyDV4r3r1MlfqWGisbxhOVr3wz7JF1HPexg7x+5lxn3Aek
JH9awzb6DOww4yNA8pWQsYdtGniJAxgpwv1hKoXruVJ3Q8aV9fSGwQytUNyGQgXt
48TsSmZVCbztHtOa82hJlqvbFz2IRRTTxe/61Np9Kr6uUHIUM3Eat4k45cpHDxjR
jjq6dZXGMTm7La51JszNXwCo92gNyA0btkkvwT2YlKNQEeOuPMB6f7L1k8ZbbyIA
idQwlb4wq1bWqM8jDqy6JZlTNYXdLLWllwhUy0KcIFFq9jFPJtxRmwhEj7qb04RP
kBibK4gcqUsSA/5FUIhCtuAPIE400byUB3tUVWOt3m6C+JwdEB28eL7i7UW4/9eU
2okADKlQ8J6hVsbOGCSjw0hXCnxm7+vlHEPu7SQpKJZ8J37Q40FQ71bJlhWtzelO
2cKeGOCarNXiciygXw+lYAN3d9FDdSFQrUzr6FaxLF6oizeBPtZcnlE4papEKmuI
EZjESB2x4zALxIpT1Xu3RmylU6HaTR6g2lXJQwH8BZJUonJ+BoGzC/9OFNiu4Kwp
O3TVdVS5efgsLaiZxqTNVNXlRvO3Zx6n4QQb8RL1A7mcaij5bLTw8wVZxzTPtmMM
frpyTx/8VD97jz2mkHOmYxsw5R5ohXEnBL6kjz7uvDUAzwnYgIOO4zPOV3IlrlzY
6fiLdD6TNJ4nOqvruQfkYtvtWA6SKxA2kMFrLCpevC4KUZr1hukFUPWYke9JCDLf
AkwW3V8gXeSSfHXh14ouEzpzRXtpEmCD38ftKf8gDtuxHd9BWevFBMQGkH+4P+38
BtUq1fLqpaf0iqefw/IuYliwTEFHHRyxHNhYCsyuEc/UmNji05P/Oq2QETLZHpXa
81jfiBZZYOtp6RYBlGWDKIOUtzm/O2qPPyCp3Am+qowXVIMcjwj4SdQi/ys4Bc9D
+ISkpmhZRwp0cQQm7bbXEjywIe2ScYdb/stGg2FdhDr9Y7Fu0NQVIgEBXT/5ZHk+
19+Kxelevskv1RwDCv+6gwBZ2mBZryRgJN8hgqgIf+bb4rtOmJehPspMBooj7Cyc
/OmaxmJmY0y65DwA6QSa9kghU/9gtJ+B7YYUNHMvvz8VtPXCdTqDU1Xu7UwIUewn
M/7/WPN/417+nAe9hyRSlwzDcCEK+GTZCCQ4gzdbHmc3AGNxgTLTaAW9saUmMcpD
7oMIrGQZCvlspU/azx3VIo1Xe4uEcQq8KQVBBQjpJBiYgaFiDEbZRlVtlQ1dH3LP
9FbRGNiDPyZINBN2imlsYip5Zoef3YSY1527fb6TX5JUFS5qB2RMWXdCT9B0osm2
b2GIIaFxcCCekrstpQAZikYgJyPEPmlTGa5+4oJAPQAKOKMpOdoQwA4p0JB2+8H1
9BediaKhHaJ+zCsHyJ+K5DPqkDKSWGL87bTrX8ga17bSlo2yXKcP7Ntnt14xdXG6
4EJryXuP6la/3VMM+S9zbat8F81PYQGyym3aYN/Eq8pNnrnoIBBHI9b60+1qqYDV
bfzrfUzD6sjHlb0ftMtyNaha2raECXTvu5MagCdX91jXOxWSEQsV47FLkudMUncF
gKOq8lybibMSbRIwxtL5Bc70TQhMw4hEnshB1T+9HWHpf1jTz719qiKkVxWnJRWx
JZaCbbGDoALX0xQYthBk93T0yoQxzQHoP0qwj5h68dOW0HEH1bnCouPmaZp8xMmm
BwMkImWSvIDxZ1I2K0vJqPLgMwY4iIIgzwjKiaIwfM9Y0/mEGWhaDAak1vvpi8zm
qic7hST+5+1YoZ9mOSeCnNSbK/MKlPThCAoGesvfwT3kPF1qhuWbz0uLcRLRvQ7z
wVWlkAdSnuElr34VZl2rBW2F9XnU5yJJbm2wqL4xQYp/hnvuZxeItGrw1f2yHObG
xJpSjVw4330X6WF5ahxgzpOOG0s3HkGuSzyHe7RBTBhU8VDQv8MF7kTazybEL/6R
x/YYhIpL3LH6q9+kV58ZIz2CP4HuFCSP/0cGtr84nZzjuMohAusBQWzPNHIup2Mz
r1c3wp51IXqJxhnH5wPiXvQmbm+q/WKvxkW4RmT58G5cVRlYQgYHAXa/PWfmz+Y6
8NK7CVYYj5Kqx31UKru5mAnnP0B0hd92aEl0kG+cocVibrSh/4LhI56cyLkL11rl
dCGABs+QzBdsqxrKT/3mrA7oiis3pGKUifjgqw0vL3TTcZhf7ARKOFgD1NF+mW+m
EjefvfvL+DmSA9vKrlqOWIDjanyBctqEMj1ANlBh8cVVEcEi8VEVeAlfgrAlH9mF
kRM+zpuD8lPqLBbVOk58KrVP1ibvxWnjGIe7Dj1E71lWxH1A5FdNtoKERyLIS4aj
wu2SPx20zBpOZ7ZU6pP/zYadzyMnRRv/2XC5CCxlHfwtzxUUa/X7BSDcvACB+aRm
HCPlRwSFFhR2FwHDf7uZEY2TDIykSkOgrE78t4siP66NfYOUMImyy9qykwQqQLWi
0nfEvNrrZyljIsXHGyPOGZJj0uEx3FB1yaiDRU2rpmIUN9xK0L2QmHXDQi9uxwSW
JHC1GDvGnjgjo/qVR7meZNNQRHyTzcOICiWEMJKda/u19Y7v8YnJLTL96C6xM00u
A3g34WUtfni6j4aaDdkLCIYVf0JE8W1aSbxoppabuNCohx2JCFJftee9Icb+VCKc
FyWCAq8Y10WrU3e9T1pf8sSL/pj+dWyYaS3HWgDlpGoKXJqwYbuBzp6LqH+OmX8r
jsaEJ57/bU8NowgAcjTbrZI0LKTBWMJcwLVOhkZV9oAlvaScl2nt9pe/0roIFmZI
qlY/gHS7+QY9RYCbzQp3Wl9wZj8R8x7YTZ3LQAVIw30rkLorjI0gMMLOTK0IC+VG
kIEbvnWkBRjhCWoV95mM5Vpa8zZMt5Ha5SM83GEhd6L3vgaMJ8rk5eYt22Cmnfhh
AntiJpPwt6Tamq6Wa34Sam/xFXTZPJCayOnzVrufbJZxmjr7ZkM5u+QfWa4us6fn
PNMEo5yVTtJfB/lYZjekapK4SgY6q8vdoJe+5BtVizkdTOB0mVisuc7uVTajqoF5
Y67C1ECFm1VSLpL6+01C+elgrHBquZ4zvN6pEQLrWRHU2vsLyRAX1IK5YLhh9vlz
at13DsgEKJnUKhcWYC6+cRf0coORx5KGs/JVSvBv+dxlTdZuDf6WyC3pbqiDS7pr
aQyuUZVUt6Pco3No9Kf+1foESwtYOAuUZS/je3S7nJ5tgVI0exMHd5mO6uRdW0mU
EEYs5Lf37hjLXSfk5SnpGoi4qyaW45ncT0R0WYV/U6jr2r1LmjAoGlzbckoWibsc
Y8bP+cfGqSm7x/t0s4tyV9U5m+Vt9uEsP+tliuQNSfWVTxdFK1TXEK5SN9o3HTHF
7devjkBitv6VKe6xQJSJjLJa3H/BvE2bHZ13VLs5QTgeIEZh4z48Bu28sSMCpm/k
kZpuvu5Nteb2LYqYy6qUHy4oJxbMeoO0u3ylv1Tkzw3yox1uJzOTtEjnnfKfEvRT
JLkIKKguBSBBnbCuA/x83HsXqnMLCciedGnS2vcvCE6IXpV/lDFf2cvugs8+EuVs
k2iFYLjJiaLaoc5zkAa3/Q6nWbKLHvlQ4WpJNiZGCGzE3bEzTETtH7tGpkAGWjpA
+FaZ5Nmf3GoUNh2oWLjXEJ4e+BhyRDlRBpJWQ4yNYsynm8Ozc1GQQpTT/S8mVWr8
dOabbE43T358v4bv/3uFGUs3dqG00KUX2/+j55VVdzFbDWqiVtA+fdjJW1uVssWD
jfdLBmapr8ZY9FI/BFnE/RMUScu0KtpWaWEVhHh0URG6pKzW4APR3zIqexnVXzyo
iioouMVpv/b8zfXMlRuGkLoJjECh2qkTRrgT7lJXQaZhlvkF2oDWcDbJiLIqV//K
XuPVviOuxtyvEQSHPRapR5QclfcKVGZWpuDcLCbga1e0M0MMlkm3jNXCBhHqxdV1
+kTb0eWfxo64vL1TNO2Ew0QDTRJG3kOMNyUSRPdhgG3/GRIdfgflrslXaRBTsKXR
6JqtSnqeDFjdTMLkJmANm2aD51eBdCI+h2tHxVW/kSFMxuPNylDDrDX3k8V63iXb
MfCHKiO6jbG/NX42/0hPVY5uUh+mswO9p6CYnh7TunU6K/bvauOLhz4sJ1kBzlam
mrB2Z252x/xJQJpw7rmMzPDduC9EWDe4TYkYx/DjfBjHrEAOxY2Df/FdEguCAGEp
oE2jsf0DXMhzaATWQD9z8ousyjDhtn3ag4KyGPINTL3obC+GlAsLHzv+7hABCb3k
MIFZ5x3cDWYVBaMP1BevvGLtqQX2SEWvzzKzfozs/UuVR5eOhlw9exKyumleW+Ac
nzhMM5CiJpnvi08UU9Ibthq0d6ulmkQw0GRzKRuVOepBgHKgUnxJWvMh17UOmpag
Tmpvyn2sXuRNeyktyepHPXYc2Z5yle9guDr8toTCKecxBwpoJKH4gy4TDnc/FpQ6
zjEx4GCjaC8kYvlRAOQbwakVekcFSxAzRtC7gdkzB4z2Cwbbw0GIqgNxZXlanUaY
VOliP5E/d/YsT6sHza8cyHKm2mYtUlozy2RYOmA1HGPIYSSAOMAW+mat02CzVfL9
SeQctJbxTNjmWTtWh5kTI1xZm5vfAL9EQgQC+qfFwU6LDZF3dQPaXA86OfETGnbq
nu8rNaC7JFCcF0PIJaY3tMJp2pTLIlufio40XptLTxrOuNcycd4kCeWauU98cqed
24SrKVs9aUmHyHH9vaUgknQxB4X5zB3YN/tF08lJ+VdHiHyCKloyZKcquGPw9ydP
qA8Y6hlzuNygQZWxkFoTt02HcOI7w9+n7v25omKdZWPRHWaxabc5HUmetoZ4WraO
mbG6ktNXyEgX+1TtwI5d73rcFA5QhLPUmt1r80QfiUraJ4hGp18VZZFpIKhei7V4
maUPnINkw91jPVs/f4FQhKCm8A1yqpslNkmjN8lJn2Zf+qKjvoMfqOsx3FQtoxvD
ELe/VQxQePb1cO6oEY3rIl9NPYBOWx+r7bUcsawRuyTsXpFZzG8AieOnt0C6PTyc
NHBeYqbiVjnotA7QI5oYMvuZlsFukPzb6QQLLRTCSMbssTatrXWuVI3u2z/pa36F
j5EiScTYg+mc61EDegHtxwbTks+fvM5IZ3P4xaq7GqsNtK+eY65IAZXZpdb87T1U
X4ToZvbu6OUkW2dplGNdqXviikEucF6VBGtgqnNOMD1G726cN0eLzMc51Ycy6x3x
DW+LOJISEn5qwqwQMSmV4veeuzTDqpbCdG61LUiNwstO6m8YDwjD6Il/4bBXi29/
0V/IV4+7k2IPeq4fGuOofFKuil9tZ9f5EXgtUZdnE3NGKD/drbHZGk/7p5O8pzL0
z8pVHwNUDqo4kt+GZ5LcEzMY0URxOyNJApp3V1OTxrcsUlykXZDFhFDCdZ4tTLyP
4JgbHEPp4AE6cLq7vForwW1JO+u16GildKuFYuwj2OjoEzrEa72oHX1MEKAenF54
0N5hrxpQt/BTO/uvGS+1qR+thvSERLP9IvkWzMc1YQn9nZc3Y9ZphKt4n52iiX01
LU7ImFT8JKQa/Oaj5LX3eJiZUX42+3oleXTPV0OXyJE4OUf4jaul50MJaiDJNmE+
2O51oANZjwJAh+rpK0Ebl8J9N8ysqgbCrurU5+vNrdVOSxQAbr5xawn0/fBTFrzg
3mjve38ATBh5BBAP4jxsIsBZO8Sr/WwmBPNIjcV4xMH6R/hUbzE1sG3VzJ/J0tgi
Lh79SHS1LovYy9ZD1RvgSpr2k0h5zGO4jiSXDMZ3xuTL9umahqIMp3disFuMzGke
N1l/EvJpODcxhBY8gq8I0tPNi1dgQTz3s5lXk18ovKVd/bEv2hDR7pMOzsXhnhak
4KXaTPTvseKpCS3lqKNVKsUp5OyYXwZYIIufdRjlROj2e8Vxc7IbTMq/LklAzeQH
3woL//4wNnkGkkog8GIxRQ3DcR4VByuqwN9T2eESGcGvTsko9hqa/+i69GTyqgjI
RNfPyDGj+CQrrf/AfK1VS+URll1PXoAlFMSZhzFXc+xPFaSRQQ8QMqF16rgDQ3M9
N/B74RXOGzqi+AooN2dcK3qRs8KAORwBlHdwgS5LNuAuNWJE59IzuX87yG7Kq9zA
CaH1BtfU7F52ff70Qqsakvk1/srkK22aIlk4Z89pdWNSYIeYMBceqmAWiTAhkkt9
ONYWGiraQY/tdVeFBaDkw+QvGCiYwxMXQE8O65a97DPIz+dhIOvAtdiWLFOgYaBG
rOE13uyMUW2v0+SI+iTzSyPv7j4V3kJtgYYNgu6xZP7Ek/dz5eOlk3PoyTdxiEkI
7ziPoC0zgpdRRs+4wXodnBXyP/3KorS9WYTvydERz6T7yE/FGr4gNYXTx3ZINVZo
9pYJ+6yr5DumF2sEZxjKNswdc/vOIBhAvztPLFyf/2iMwWOtaEnczpiwv2bZR1kM
/8eghJuURc3f1wVx/R7GZbrVLRKwSZ8+uwSvA3zgMfAA+mId/niZsImLJmjjI0s3
O6oB7qFaHER01aJUoRInugrBVCZlsfTHXYeM3U1MBBpdJre7Q6SiFEMjPF6b23LB
91VOt5LF+piGjOQz1Hnt+/4QRrZn3XjGPiOCW6nUfrqONcAUfyvVO3RqWB6e4mEk
6OtOGfofBeJoL7eSxEzUVeHA/fgRmYagnYX7pvyK8XRS5SvetUeIrYF2xfRVx3Km
N/MAbf+Ux4FzqEO0ValQmj5sbBfwaVXg+5PghMmIR6vFxfbyjmabAiJNxIMOqigI
tgDm55W2WeeMD5jlaUtcgL1qT8GGSNWYjcGu83M0yADqLk5MaacqCHRGi3CsMeqe
D85HV8UWpe0MJXfIPptxmjT7cwcpG7uNtvKbVDdEjIUioW751orFjEf5/aE1Dq97
0pZDBJbS0zBtBoj9kf9/4DewFKxSVZ1uSl/6PAGRD0NvtdTDmZuv9YY4+rGgJIP4
mbQNI8rONkojDjkGAoiDINq1pUH2YwW3cnAQ8jsdNcD3izhQq+1ZAaPKCAV0GMww
fL8tW8czPxyUml+7awR68fbjAS87a3DUVWl2mXr8BPzrHeRk37JpMEbrLSdGVudD
n19HUo5eOKBYU0j2cmzYuoV+SsJgIzoPFNW6DfdbBPPYY4MNgz4X+JOWOBWjKuEy
J/C+S6dN36fSjaAwCx9Q95eLv5ZTzbz4gFhrs4cKDWUXFyKJTZAed0lbY1IvGTTD
MHxiZL8k8ZmR7eWvrL9LlvF9nTk4JJHZh5eNkPQunJGuCwBF0hrsR39cMaVkVWjw
P/vLa0Tbqw9Q2koIdFSQF8SNLQ6uWn2ag168v2b8Fbz2+IiOmt0KOkG+eZ5p9vwW
m7b2V1veatHUDzC4JLsrSgw/YQFBKV/zh7yQZKc+xXkMkk7jgkKRV5+Xjebx3Iyp
/MGWuJlh5g/tRy36jSy7vXDvNG275E3ehu/mN2Lie3f+xjI/RV4ch21G87dB7D2f
jVJJY3kE2di9Ih4rzCe06nJKQOcXc6E4djhIWUkfyXqBYS3vxLPvxVv3unOdkO5x
5YemSHTtdPYoKqt0CkmAycMeHd2UZklolV0SYYKI/yZlzqQqaVAeWR0+JB+sF6dN
lSpb8bYh5hPWsvFMCj+BQt/5WDWh54sJi2QlwV4Hu1OYd9FPq8vdHC3y+kxOOVMV
cTYelQYxZGwy4rpLtnTVRGiyXBUhZTP1J3/m8G0Ij4fh871HRPE6uNvVrKAoLWjT
ktrLz23QHvK39xdb2vegrMKgk8bHPu0ihOsEfZTrJyXQjXTn9sYnYYmKDTUtAAJ7
ri7hAe0iDMQ8OnK1kEaQshdUYaajzywbEJyODQfPHFdKeCeRDP7urMLZl+hk9ZAS
FNZKZbt5SuBVV8Pjv3436Z0eugXDqing+/w5fmaQbtTvVnq0Qkn7NcIrS5y+4c8q
P1uKPWy8HhV8w67sMA9nBtJfYXeJrx8Pc73rSYxA/6hgGiypFSpFqof51E1I00WX
Iqj+ncGt0BjUqgM27SQmrDFXfjp0kQx/p8oN5u9vs3xqBDl+ijy7Z7019Shs939R
yNxsAwpfGBHqbxJorpQ/s2552lcw1ikssJQAzEaar4+5MVBYlprKd2UsJRj/hx/q
tO3Tl7WVOMDrjVR8Noju7hBO48tXT+JxOjKk53+MwUfwf1m32UssNs20I+vW20Rd
Qej/W29llH7ICGu9vDOpJR0gv0HhWQIrRDmLazsCw80TfdkIfoj5f7ZpIrgbeaM/
0nNhLnKGwZBCnSEpSaDZwOsPW9pJxrf+n5Rvnez46pnCMOg143WyhRLs23jpCOAX
NZHtt2IKT+VIEQSHAu/aZ4+UFwAWmh5dIU2e7r6AcS4kxto0e+LzI6X5yvbFeIqi
hVxFjjzW6nQr/MEiQazLUrr8XlnGZKdLhULH8cAFXht0kVZ1B/0bpyk6EvhA3qyX
fnIgVvSevjlkm1VQ9ZuTqmO6Pi1PPLmsSAVcOG5RrnOn6dwLueZeQ0Qo4GBRa4MN
R+5pVaqE3hV9nPkYxbUWSJhksP0fa28e6mFgQNzurQQufucSMSPArcPgDtW0qAAz
K+4qLfElBJzeGbRd8PcvlOLptL4mer2EgrHvfpWSvjBIdczn/+xs7jX9WtZdHlq7
e6mzzOwZuC7pVfC8PhfRjI6TW/N8kyrG3l1RjyWMf1t+hXC14jqd9wbQqskxO3LF
6RC6r5O/QlN6qhnAYo7d3wePjls9YMMVnNtQTd1i/sX/VHclUu2v9oD6ImBxE23x
CjZmpwchfQoxqiAcirNPtIYuOi4fFm3gds3UGcCWFBX32BIt/uWufKGoug2kM7x6
VGtQjrmJp4f3+skIMv/nEsncdnqhtF6yrXtVUS0Sx5RxIh4Yy8Hwo5cspUy6fl8F
ggXBC9e0f3g0jX6nGf6l1B3/UrAqS78uNYxf2vlQOEma0bfG+WtOSvh+LA0PiPNZ
ROr9oFVtecBjxiua/K9/fM1lkV6p6IX6lo0jEoNg1FuWUPldtLOhOjVorMGi7TeU
q9i73G8WYwRiQ9JEns0uZA54NHDCKh7UP1PeI/Jk/90UZiRSzI+z4OP1w33C3IU/
Lm/hnJCGvicLPa2Y1rityM8rWe7mfPXArRBcuhgqibdShtKfUlDxzFsEadycyIgZ
dxTMeE704bU3gxdWgtLqhq7Q889xr60Wn4iL0miH33zrvzussE3JgxhV8ydlR5m5
554SEqKW6yXsDpJCo/7w60mVC8wFR+AKSolVcMZkzosq83Se+jQIFzIf2HY2g5qY
MOOS+7cFaISWS0PEqpkSRjR7+McKMZVTdPo40NgHxPUQKJyFD4gsqnABNPXKYh8B
SWHsKXosacyP5kqEMW5TUDgUOYiwXdezG1wcQxoaGOp1MxWb08lh2QYmACIgk97I
x1iQMEuN/q4Tdy6YZ99lG7YoSuHyHRS9c80anWEqrVXVxn1MfehfK82LbAc3h5mS
esehXIv3XsYLcjJZUodm9yiCl3Ltlzn4U77nv6e9HOOXTcWn0sngO08/LbaoQx2N
BtmTuE+PksIBy2fpN/bH1+uxylxua9+KDPBzoInIwwFrA5kCjJ5IDHQ+b8c3soKe
JVnj0vKjx9W0Y+CJ3lx7MW95RjyirfFsfKb+3OORd5Asde/6NpDe0WOB3hNZbdL8
qAOSTiYBT4utzfOdffz5/NSh/U2yA8WjRpr1aKOKfNWigHIbLoYQpnyeMlxzpeJu
Sq8KEsDqd7gFskw3TS5Ol12oo8Ezg9MGkjg35NBn1c/vOYji8Rj1lYrx9rSFRw9d
zPD4gu76myzt30R60iovAUsf4mFc8bPMFwaWn4ms4gU5QWNyZvPZAvthnwHPe86r
Bib2ehzlgOXgA2TxELS6T01y90l4Uj7qbtYVTTbel6NiO1XcS2ZtscF3Om7TcJ6W
fqyZoOGSSKBx0OODPCC6441KQTrJvEN7H5cQK2UPjurJ30xHESXQA2rGYO1nrzHP
25UhDnF/jRVarJo7+s2qu4V0UnmQ1QV8t2xKvjd+n76N3EBjMINzmzMoKGgVQ6zh
GMQjNyjC0ilJZiWd7ta6W2tbde6fqjzHmo5Zy9/XkceJcZR64g6BUirl3FuVksGB
qb29KselTzJ1lQyFAjpMZdW/1S3oNtRJYE2jFdU0yLH7fx2rBNYd3twXHoAdr74g
TiLUnWv0pdBVU6dOoNM+3AYa6AFjaz82lhQnmWcaP5enWibd3jqK53qCoT8Pjzng
g53fdufQCdAMJZT+o61QL7DCU8Dn2dr8r9js1/ejrRJtgTLy/IC1JwcLQO9ao7AI
5glDbIXnmtcwCy4gLL7qU5OEkeFlEK4oJ0DXSQeK6YksfaBPauCofawCzO47nmB6
7ULWdtvm5x1sAmssigMZ8EM0NMZfrremg6LxllpR6HnwGiBp+VNNDdHnu8Pz5aob
UHHUE1RjVYZXMxsg50TRbHyzbTRjGzYfzxqKk69KDmGE2tDP7qalxNOyzKp9ujd1
YHB5uzwNqtisV4P828wa8eidFZwXws0rWQfvBFQOrpyF4u+7v5yipVLL+hLNJV74
xjEbB3Q/AK2TyVWZTiOBPSC/eAAAEoGkGMGsTzjvoKZfOwpSkDIbuLlhWzTGxj0a
adCg2Rt7vFiLQgI371q0lkURLMbBC+pyo0gCPRppAm2IL09XXUCWEjgv8+U6Xwyc
HZZ6qd6GvBGPfQ0vWvpY7bS+I2C4D1qzJytulgJL+H/1uurrr7Sgt+YZpUiReWXI
b8PQADeZQbAnRSrIh0TmJNu8FED3W4UBO6fLNouGagnaLbSLWwBpRulkQNEwqbO9
rn86jmlwXwoqTFXD9NOZm0vAuy41XnRUHxgbfzrMJSLlJrsNLfe6bKh5BQtAZyks
CA7nm8XyPHGb1cShH1iRMyRSz9jB68vW0HYbhoDaHYza1ILsy1uyhh1P1OpfgNsU
4fKBjoR/wkvdBaYP5+jNV/wCDapqNJeomUFe97Y4E8r7iW7h0atNrkSzYu5ete2O
HKF4HziPSgsvM2Wj2qzu2PBx2U0JvHBnDRLQBfM9y1bgCXd2qyeRRDkMAFjoL4JL
v5ia2NmZdV70OFFfyLmuFTH/+ArtwD/ovge1xKmu2xBN4wTiDcSBBJ+ywzEpkTRa
1PnIZa490EHiEcUq186JKYcmDAUnlWAHmUY8oZx/gFSy/FCsL5ReHo//dTSsmYEY
N32P4y+x/K4S7CFPKSqhApdrYToLnOuRCb3HR3ynh3699mCzXJLHS07KiEPN/11H
qSCHQQ5+oCyBHrVEAoeKPYOc8+YNvPCDlYTgXlp1xW7yrgoXd/66iWpkxZQpUEYe
4iNTdiu9DfL66/yw0x7VV3vQdw/CNVdrC92+vD/0mE5EuvCjafpTy5I6+kVBEo4R
baphxEXbuW/hDgSOec7/QfoueeuS7SSPqmy124MxgACqsbsNGZ/OzEHeXjawvbqr
DNR0tzWcvahrMEWw7tfsgHWXfcDs9cH5tCG9JLPkO/W9UzDT4+pKqTKWk2dEcPYV
YYpQKMrl04e6d4x3zlPQZG23jn3RVDnxaQtuMquejk/fXvQFmXEZ9geGktgVhmKZ
IF1lBCsFrqRHvvHHtnFUK8tW6ll1lBC6ujpMnAIPHJCLpBPK4dQMpbr5jOrxn7KF
MhX9i9dMqoj1G4NTfGuk8B/tlzxlxm+o0aelafbaAh5I2hsSBeKnGmFmzpPYwKjI
FmMTf+1FDCaia5QZuAv8xpQ5YE+SOre06Zva1TwabNPcpz02LTcMUnFpTpcns+0p
IJscb0sv8I9coZhfKrzRTD0WEuuLlFGmiZX10mgBaVgZ/wtRJInmRM6SIbrLTTZg
4BAfLN3Uk+yIwonC4AMaMdk6rogTD1D4l4iLOknVtBWECjtsFK0QAodfxCZW7K5g
SPrr491wsAbADea2y3F5IyhR6JHvqYlUtwt3sRBzigoXBcuJw5yhMm5w7GOpCJTH
/2HE+pFi8ni17h5bJ0YkR1N9Khsm/iBEcVWFWOwpgFp0keBuhXHr1Q2oysZox7+L
nuxUKCi7PwvrCsfzcW2FxWs1mckSTYTAxssdoH29aQRkvFwjmrh4sMxbfnPf++F0
JEkllcgIxM7JgZBlzTyuFxNmEK909kF/+L314ogveL5FAyQxI4gRI3x860ooPXqf
K5m3MaRV/I9Qqd1eegKlGvJcZa6aRWb+PkLWHgkg+W8qvub2uKGsi2aX3t154Lyr
V+LNtih/oTyCHiAcEGR58EYTVq7TAbbVPToWGBz7TNp7mJhzp7HNQGW6bKJfFB1g
jEFF34Dph2xWjJnfNIPUtbi4ycq+jpWEqFDHmxjjHFlWnK6uzAsGN/H0O/Zzy7zp
aCWd2+5hE7uVZhfPmYhLhdXJNYGGiYdCq3ofFcD6dvlVawbMv7hqPKfocBlZD6HO
rt798jW2rGBfnWMjEUhWKv8HD4Up5Dfto0mqORUsD0wQgqbKP3tieUz107OV7ZG8
ku+jqyQ78/HXVTjNgWp3GmJCxRCG1IdeUqJDCYsJ4MV+9qwT8fJOM9LNJAzXJEAh
t0SoGGBFfEkSTtAW7Ttv9E4/BjmtmaNjQh60hT/AZ0nRbXgB0X1TCZ4InhsJPe0g
rW9/nJat9lSusPGtN86AbwfPW0POuj4+PFAtAMOFPZFvCR5ZF316HOD5W0TWjwzr
pSQhC9tV8ypHC5D86y9FOVA+ygs9ro+muwi3anzCvdu4x7ZceddG75/K/MTuWdJ1
ZTWsKPkGHxz7JwIvQTidyppvqaDOswIoK50muwYcvR+QISnOUXx3FWbqYtZiLKNk
bhXneFdAoQYegCmDdJArSMTYaD1Un1Qba3ZtjPCwc2U48rbRPoqEIZ81upxT2sSX
4XieGvnJezsd7BeJAltGhxsUj/K3XypWjnZWSOqVKsPVqwr2FQxnfTu/oWhYnFN5
deGYM/w5fl4izoGgVFv72UVT7DP894gypy6FomyvavbzCKIpC5EMvzhx+yBZTuR1
npk8bPFC5NY5e0e906VnqmQU/sNaNgwkw7ZpHpUGrxBDcGUUVcVOyeiIyyaB4QF1
1NSpERqvemKsArDvEfPtAMZlb+peSknGwcrUUhXpjf9AXcobhOIUJQNUtzBdGzLI
pR0jRsRXqh9/0djtPkvMIAgWw2DMoxtaC5hbrWwwvOqW61UXtZaf85HM+DILYfBz
iIvD98nwY3QXp7d8OEuSkRw2wGxQW01e4/WyCcs7P4s4PcTZDMpNLVoHO91zuGX5
zWPH05CXuP+YNffSOfbUHbj1dus0s2lFP9sWY/yFClVbiXByfbvlWyNwmzMiwr67
x3NsQcZJBBBNDqD25W2A6YRy6BNIZs8+bYSpj2eUMjTCaRpHvQ24/WEJvmV0NVUR
KKPaNKs8kOZaa4Tchlov/g/pXux7DTLWyiymTPlq0hreMn8IZ+x0Leu7n6Eq5hmV
3/A/bXQstCCerxqUlJfeibxtElbcUNVafRUufuiUQb2O8UXXD+hsGrHBJl79qh61
rViEv96+5lmDhl3ubo7MZkM1GQvhLOl4ojS6e1KrHGu6s9d5ccSt9V6eUfw7939m
56D/Ct8jNfZ6phLSRWQHMdrPTvpICTZNBb4DLEd65/lH6mC4JabLm2E+zSmwZAX0
yGqSbS26YQVs06xlD+U+wDRVnkMiCMwsH8oP9YNQQ4xCVyBuedC2I62JzZ4uxU19
FkohLhrDtzkodLuPLaqoT1DVyVN4K1G99tIcU2x8niudvjDQsq72tFiFUBy4/BOI
biSNpXxFsJaqkB/nqrkeQfcPtXLjTCmuJOIGs/GiXogjuwHPAXovBK5g1v3vldTx
w/P3CEiwd051+V/IfB6AOdGOc2IHzV+xZULpZXMhlKLykzebWhV1+TuP5hWzNqjA
pqM3AgyZo6MwmsKgS3QR5NCrPb9hcu5b+xtQd3UW3MNPUWZL58FKstA16UcyIl5W
rBWcOq1XjUxhfO/jqIEnvWmsNTqCAgnZ5sPVNhbHPzqb726rs8znmuxpiLJQAPc8
PL00k+82jT6r2tDZfvvyjZCzXZ6WJKCf1AQRkLqrlPiLDqPmWgnnzwvnX0Ukzg81
lOqPJqaFF45cPycujaRCUd0xOUxT8B8Z3I86IH9054kYzczJmyBlnyyhjdVD9prE
6FOnUBrKBSJ1wzvyaebHUxceHrrAVG9RuZdXWjEJ53SHj7HVGXIPHQmYqJrqj4C+
gA4EB0DjZgL3pUSHFKP/P5dcYoau4mp2w0KvJSXKlXbm7ZYwCLG1IYlgy5jNgc3s
pcBJaC0qzl3oP6aO/pV5Rwt2uV/oIoglA85nlNW7eW+rYnanEOJwD/V2lzR0mMRE
h9Ryd+uRqezKEcZx3EOqVn04lyBk3Bc242+FSZB5Q21yFMKeMXrfOdWteU+SFoeM
0rJETXYHHmUbtcx0aU2O4F4Q/bjEuwUyTEvB7L2gyGHi2Vna1NUmteSFR5LrZtou
xt5+HycYX2bok0ETLLZnB6Pz8MELKMMfYZ2MncxlVSOx1t7oeeU27UdQFI7J2BoN
2Pdp5CYmpNwyk0s7MKcii7V4laN1vef+c3ovol//JJCj5CpT2oarYgajxC98TilS
D6GzwV3c3qSCgaC2zWDGWXNsdLGTdKe7qjD47E1PLLPFnZAcy387O8fei1OLK2Tt
I5l1kx75nE8+OLiArxz4wwP63ixeE/IdUGf2vuzqnwglUv3l2V19e0eiY/lx1YqL
XgHvy+Fx7ityer+ZCWLL6Mhh0a0mri+80YuI3zmuQOJHrbzhqU2Y6fyXt72aTHuA
1F7QKmnMTJZ/J3IIpsAX88sdywjNEVss4/KgjOAxI3kRnVnMZQqfXlo8smcyZNoN
ey84pqKo8vkhVuNNpXogHYvheuQtcZq5yHYufFNCcVJvoT9v/z1aohX6klNMOFkK
9e23cJAnHgKfl4rIbMVPlZMrvkol3A734sI8HlfOXk5RTyxeoT9gz0dXxQqLEba3
U1jRng5hXBj0Z2/HZ64CjdQxAr/C9Rjmxa2ElUqNYOiipHwVhxRfhKG4UUZGE5D+
v4AgozqYvK2zPjB5a9rpnqhtP5WcRxRenhoSYbXGE0Qy8GukozHIzrx7f4Sq4fvq
4u+6pK5NlkhMdDgcpgPBGss/sAd1EvxYjp9eKlVkRgahfdeqMfVJko0KG7kXRTO3
PBz+4RRkcz2Si4sMhYxcCqdLUOV5CgCAkOlr7kwXdAPROm2PJ9Y5sbho17R2ytqM
SGUIM1VyobhfF15Nk5oZa8VZ13UgzdZqXbe3B2f+DQvIOBrkzy+noXENK0d+KF1/
uAEycdcpOMxPvNAopQvbuddPdGlj19m/Tpw3G4WGipqD4RfyfLqgHbmytLGraQ5R
LpnEdzND8g16kteHooL7Q1mcUcHTxvMnxxCC1gzh/0Gkc2hIto9gJGAdZEaq6MqJ
7er0ZlA/e5jItfPU/+GqWKOGGvkAKR/25xCg5b+00peAMHWAicnwPt07cgpIejdD
7iRw5KKYRi4AAGRAOPZJJSgE43NOFgSmEfVIBoyflLm4w3qu24xTlB5oK+asIbhx
JcD3sOZzVgxL3kM2DgbpwXQzCwLAbv7jvgAyYP8A4t2Lbv/VKSpddRgfCQttUNTg
7s8EpAfMb+U808l5zCt2fREcU/hwFuF4MGPGSI3pGbwKWgD2YjvN6ct/CaQ09BXD
0Akq9bNB27VBOFAiOj+qNx6X5vfNS1aZfp+WJs6nndCEshbJlQsWWdRsVlfSiFrD
ewohUevcGzE8hE35EH3ekFD+jQLNAuskb1Uc0nSyIq7jM505UUh1ohs+dU20s0Pd
qBGgiuhsBI/tFzb8XSjyj6IzIsPTAQvsvwychNQZHr30X2HjnqNVCJkA1rrlVNz/
ZLh6jWS+ea5xxgQtcAAXgzorcAr8iBYDXIjqvfQ1xcJ6HvG3EX6yqwb/qMCNDERG
P1a9n1yZ1889+SEApKQM8zoT3HqyLHKrURdfIB/ImHLG2KqDdMtmYF5ieJTTWnUk
1u9V5vEaWo/nTi7v9GHMH/A2XVL99B6KnREwo8CEe8G1N36J0KZxq0HeP/ir6pw1
bnWKIGwITDtjqJT6WRggcXgOnw8L89LIJudn59UBiBZ7rHjtSkGkpm5L8C8TWz5z
r+2UuLTEZbwtGQhSgF/jqe7MN2EfqlRLQYYQQpWqj132eF7JvULKg0H+Hrg0IXsF
tQIe3c5JbaBrjLjyzYXdX3gIvgmjz835ze4smQu0XmCKZn8m+r9CSUMtPP7M2V44
9OyY0STIUZ0c01BwAALhlMpPLau3jv724veinK6soJ+g3tjtNStu2z7lt0tM6b7t
rwRpaLR/QKlIbspibK/WAU79U7CQS5C+LYcWvHfM5dM7/WW64xg7oN6UBZCh00Kh
p+oGrvZh39TDpGp1AvryE8S1Wc64NvnE8fy8cZ2N79ohpR1lP2tcmNhy+MA3O8W5
esNnIqRX1YjSWAFF3WdgPAES3xDxFOMf+Yw67u/u5/mGujD2tRzBJesUKSL3Kh4K
qBvaVNYWb2G1T6ekUhzK2iBK9hHVjBdjh+QRcVVNZ0jAZ4pB+lkv5mPY5dI79EzJ
n2M6hDFep3vhAMP+EFs/39y9ZUZzZudNv9AxfA5qVDnylgOahP5IAc/WLXg5KmTH
eogbtjfsbY4dtodj2E2YKJ8C5VP4G5IXSPttIIaQGgnKI4/UHiGCf59K7LWMS/8K
9mFRMus7ADyMik1yibs6kiPYsRM/T7Z7UYObKr+1yduy5LvYwqbzuj28f4S7ylKN
IEn7Aq6WeR35RwsRKqV0fTplOu2IsujO1cNjNIsN4RgDkNncw+Y9f8Fj4zsmY/J6
LDL0V72nBtSLYb/mgfcVb21VqEGPSS92P0iN3PbEtMz37/tXj6ce1d1Z79K1PsNU
S8BEOTq26xM85dcD2s13OHEHmnpwirvR/eCp/KYzZtaU95I1iNWfpskG/aTDOv0I
D6BuoX1U2jkXuhakEJvAZ3GICjvKj4DUacbPeZC4+bf1aPMIpN/+6JqCIoyFKSqF
SXc56M8XY12Z7+gxNiqScW2bMTpixqqijIjuFDr1H8d2Bk0mv39jHdAaChupc3OY
fMKVXRFuaUh0y7hBLDsuUNgbhGR98tEPzn1Rl7BN6DRx++LARzUAyHRaNRr0LMfl
jid314MVZLv4ucgohLQFJO+NFBewRz9DCoBGy5b/bSeo46QuSok8ECmWMY2NfOyf
N5O+UI8+azpc4BI5vOfDp2ivWEvhCHQpzEurXXZEKKSX6cnkuTGjyu3RCVUQMMJQ
7tZcneEXd7wtPxFxfRoR0OLtERSSWglNrzU1ybmKd7V0DPqRZS6B0b/z7T/88rDN
pnWp/uoZUlRjeggSBZW2gvk5N6eErLJ9Zwvw9ilSCZvYb48743gLgB4tQ17eXPbp
Prkh9M5ZmWUvbAKwVhGm3amdiw35Qi+1PajkfV+PE9Z5fjDCaUiOIxRWl9YgEryY
zUE6foXdpv9HhEDWsi4C9pp4BADKvNzy+aXGDnFq3N5wXlTtqkMO2HksHrliQMAY
GyQjIYPERXkp22+0F5sh+Pz8zucWcVMSxUl90E4plElu03ulzA2ngE82cixPP3pD
SirE7zu+iObM+nUCxhHSBzATTqzB5f3PqjtnnxvajW4Q18Zbvhy8pkOjIBJlRk/G
BnESz/rTXGDz4dVXD48R6MTgii54kVHFobCW81RBjxDWko80ir+MrFYtWOj7tPNI
6Fr5wWg4mSC6A13JUoVZ42GtYMYfw1LOGhvNc6jLYgVcha6ZBz9dqLueL5uUvgf2
7jALgmJ0+wyUXV+9EBuE3S4mi/Bvfn4pAQ70MYt32MX1CbU6bkKEKFqlxf7/flXI
wJWGcBWo41JPBoVeLgdZuX3eRI/dXZ+cz29gW4VEUxfDYmuXwzE27Qy07qcX5Rg5
VpXCelgn4H+MWVfpAeIvtAwW/9p1efwK0YjGOcIcwl2nf8NeiFjNQVREE8fhd4IW
nDjeV2YHzbYWNw1Lo4CErjazF8FQ7Nw7bBHhJ8uEto2P3pj1iLvQihvtIhFg4Ykz
KEEvynN/DQHUnxPkW2gRjUVeOZj2lF29f1HNACuMDFkok1ueyp4HGZfHRm+DS7q/
UkKpo2TWFs+l3jX2Bk6AQ0DU6BLn9Zku06jpsVHlgGjmGOkZULHGemvrq2FjDDlc
5LBFyNoIPHbGRwBOsGo/LzyP9UfPZEF3tsBBssJjnVAXyDr37JMgbGpKwmRRlY4O
0I0xkGSHYN9CJWFBqx8rXfVbT4JWHNpPL19GzSFauXHVLJ1aPJsVTIHqybLXYZ0I
EbWx9rb2Qav3PsmEF/0ADo/8a5V5xffSOsAYXZKrtOhDNh9e6l3GGLN4Rkf1livQ
43rCqPx40fBqrm2BbBzFlm/K0Mh4fhqH/OKrXpmXGzGWnaJwb0/7nfV+TGng7xZ5
/2ISgpgQ59kB+HnZm196XKh53tcEwkJBx36/gLbjqDQNTxQDPbUNMZKgoGmsYw9M
2Jl9+lGT9TqTnRQh+iJBIvMW43QfmpaqzfvflYY0bBSVeoe7j0GksuWIt4UOrCir
zrz3gD8EEo7Q0HLGHkkjjk0+96ny44p5AYA0OOdkgcWELDMcU65ot2nReeqLsl/s
/khMqsHBKtbzOI3OEF3tgjZOdPiXN1vynrMcaKrfPXvASxwbCcdcCTj1iDX6cfWL
VUnif6vKLvFCKkmnQn0miezsXUc/B0whQD7jgewfg/NbJieP7g3tAPhkt5z7EqSa
sc9HuNCXSf4LPfb316CDGRcEFMeox5cSYpyT4umGe0ijVUY20wCayBj3+RoB3Biq
jsRgComF9VcUv7o/twjlI3JXIk+B+2svt1L+snOAHW/Rl6+hQOfVyNG0/o1fTr9T
0zW+TVb8BE8vLXhHok2PWn4Fr/1NBoOZUN1frkZ8g54PbDM1n6oEz2pz2u6t0edl
SuQ7ItEU2RkhBpJUFy9jx7IF55PvHfkZ9pCkxJgqGJK4JQ+hCAcEVbDS/KwMCOEo
pTVuhyW8ltrXTBbh+B9gZ6eEHtT+Qtmq9fQaODUYQwKmtEttCHjBdWQC33bkOQTs
qc4EezJRg3vUO13Qa+gsZt0t5wXf5WyFI4R8IbFW0NaUyNTeXBNgMYpYMm4KUz/F
Oq1WU03reEz6/Px8Swz0oD+GI6TLP2edaMq7x5O8W6hgfHXUVLoAtZh0DCUKBDEn
ngvl9RSybUpZA9V1HhFLxWRIVnpAh8l8uvdCeJ/WzP6U82TTtNxiiy9JsEV4QM9k
pt6M7hXmM3geE4uf4HHMPZJli08G0bkd3kGK6hcVUeOpC9Euq19/+AK7Oj5l9it/
h5/HydXxw7twLb2/NLeFLU/v8wp5GaMvosSok1tDMln7m34gGOkm41nHsu77BV/4
E76h08v3SwPbIWZNdzTUKrOmL6UXzlyX0IHkQwSjgYa3rjXszmlHwpiPk6REhxas
2NUOABMiJttsJ8L5I2CAfIQp95JSld9tfyUbMicoQIrQEbhIRl9TGQDMngHblo+T
vUD/k8POkPgvoFLTsl1NIT63p6pVZEiQTVZULef/6FuhF0DVd4hcVyIg/8u2sEmd
d1q3/Q1CoUO6K4vN81DQ7Ezx7WWwiXkrNsMp7Z7dpCQ5juvlPcq6Fmw/gjgqwckz
YnyYamKNVq7uf1QuMHWBGHhJUwWNILmEbV3BzuLOlh3H9ucZ87zCN1qJHtAD3QRl
ORQmk+BpQCFAO8wH5upX8uxfM1xDWVbEFyhS2feo64BNUB9SdQujXo6uuayFU9kh
sk5Hx9XunUst/o8fWDzREHQF4LsfjsRgTGMJR9Z/mTUVqFbM5mxgtRAsJTzVnYQx
bEfeLwwMkJzuFnFYhPCsMvOlIBr3h0LUCOsQiPmIGLzAe51CPGgdCwlVcLzsGd3U
+k3WBavbWuz9pwfd3F9p7p8HTxHpshMa3jl36HXOZdLejOsaL08OXWW1EVb8p/WQ
CyWJYAYtgB5V8/QryN+hLIIqy9a7nDejr+sppToMEnH0UZVM6POfD+sPpK4LVj8w
lIg7dueuL6wcse57cpK+MJZRo2wNrClYxfPsZkFrAqzee7I5zSz2OeYPaJ068HmM
gSvxy2AgvzDJqssTrPN6X/fBoklVQ2yAI3Omou/0EgvRYftiIIpH23uNrquwnqHf
VubZTlFtX7qQ2TuKKsUTO/Yj0RqONDNbkAQD3b9SUiJbLc+za1WR8/lb5aj7tGXq
lUObYMucUGsCs1XIx+ulvHXFyRYvfk3+Y/FGRBPOvzR5BTggcjRWWJw/PAiMHPkF
BJA3agv7K8W09ZMkynn/H4S3jR6i8mq/TAtKuoLlDSEbWqQTctaU+2SUf8zUO7BE
IGgKevvcbXbZpDlAUNBD7HIv3x9f7PBoMVMqalUJ3NRjF3eXaE7buWkqex5Tyw86
rR5TsCfsYZiSWJqutvpAq8330OnMR21ARz3PrSBPA+EP+NDLK9dVlkDl21eF7a2b
Ls2FPK9IKhZ/TfWJ2tT7srp6U03efU6GzI8VSnl7g9ipbeOHNqS2st0l6AopfcjR
xy4n6nfg5e6vQxg3v2o9LCMUFji7a7Nlgt7+ET8e/6UyThwk3gTu9pkrMknz1dNn
PzubhmJ50Quw9pawA3rvDRxW1LlvqliZz37sn3KcJkHlgqXbomTTVeALIGAGH55P
c0TYs+T04goO+c1BI2tOS85Syn892VpOLy/EPs/Pu53Lq0LPu1XRa6uMzvLOsAD2
VFdmDBYNMZxy9X61NLV+xnHoBHFGTl1sA+YFrHj98qU3L+q4oiyfhM7xaqiEwF6X
GyIgpAHU6u3LgmuOTRTIFb6huxZtEcxlL3GbDSVVlsg+r/Vu2b/Njw4910Hd9Caw
Sh10/dhjTgrTDNAd3W/aWPkfGMYVOw0/QRfiRLuAvtrPdfTPzGjOAFZ0XRH6UQF9
TRNIv0A0zxkg2/4Q1iMVrjhJGl/Fop1FHFbcFBm2yJfmPDEwD0KkWefOk+VXV2ID
1GHAOPvOeKL//R/wBPmuTeMWmWVnPYw7fh1rLPD/kGPP+f/1nK9bR1PRb9QbFDbn
SOLPhY1PX9ulL+8MvXqEXoT63nPpVu/MKZt2OTxJo+62G5Qo9AuwKs2BqBnidn7q
EK71hDQ2NZvlr3F6n3PofW2N6bzqR6BXStkELlrM0EkwQiKtxj2wX/WFt4PDlIF5
3NnC+OfVsF9G4TvYjyVnM+rSNk+Fjb7TbXKHN2uf/UetA8yCLnlZ6H8f8r5/bez0
3c05boomWbUxvM9cnfhaGUjmbXQx/FfbKn11sEHg4QYxSg9afs7QNUYC3Co3d8pK
RydqByTZnVdIibUozoi9zk9Dxj3wCMNzIgBreEw/gQNYw9XDgWtETExL44qSB8hZ
3c8dJOln/w6GwjN51mWtPgkW5mvWLHVyqlLTkQwx9RCIefWeLtFYmp9tQ66ibgGx
CotJkSDFx6hy1jV/F6i0Mgqsz46WeNMaHAJUwcn5lw5wkDTT+75MnIMKn0Qzhjbl
OqxPjPibjjhKig1JKUb6ZOQP+F9lwNwn7vc75r6OUF2Gm0LyxFsIbjbSdOwBA3VG
c5zy9uo4usU2c1VR/ZkQOf5K9VTGAHBU5//pM2GNYQsSGewH7VC4snWolB6ZL8KL
MlsAZXnSrwfJX+hhCMcX5E2CHIaGcepEVzt8HRLQarM2O+w1XA5grXE8j1FdKfFB
jlwdO3YHN137sBRmDkVJYIz8C6dHbLfzhO6WbcfyYuIrBoMKwnwsgWpClQOeTHjN
Fdl4v4FVQ8j3c7jDQ1k1w+WG0jFSdqT4M+WELemKpP4YD+tL3RFk/RY/eVMzcq+p
RxVRjZgd/FbifVMuCnktGbOJVY+WxhafyF+IvwYXbokymTZneAmcoFvjPhTjCcQF
kDtiUPD6IzMcSs4C6+qlHlRVApw/pl2A1aAKRqcLuInJjuNBzs68g6XSDbrqkuiG
D/2JUQBwaqOApxEa8AY8pIONKMIf3maXIQkAekdB/ExSRZc7IFJC8m/EC16UnkWt
4bymY8Xt5KkyxJpGhWqC0XYWJIy9m5AGol15eofJWTmPDCwt9vDZnwlZjlArfI+9
81Ja1eLwCrfIB28/tKAAp2Sunyf/E8MDS/mODy7yIgCoSeD3G9V/MscvScyfI/kV
jzHRjutfc8uwSysYLMHOKIkvvogf+uFw2NxhDliA6rbT33uoTA4CVg2JHVgjt8dT
EUlsEtO8xpeAgSBBu3CvpeX6uukPX3FoKPPlP80D7nWFirUr3h9LBS6nDMZDY2Ax
1++VMWeBWOf6sMfrvYlLKEWZHKsvty5L/86l1dO8+Tq6VMdqMKdSWEUQDBBz71k+
BjL3FcIW7UFS2Z33zDtFhblEx0yjOxn+vwW9JesxjWsO+rE3Ge17leNvm++4vfCy
GkVEo7ZoTqG1GsXy9ionC9n6mpb+P59XdzQtVK+gU8vZg6iTICUZ/D214bqyjudT
SKu5VCfTOklWzLGvErsQsh6xEH2rXBFRa9WP/Nbi4ELW3zoqGSJ5Hu3636+CqL+Q
iSv2Ct+oocPTfj1RhoChu2zMLqjhZOh18rdj9qAFnC4ih5fe4EzgAY1LYgWn1DsK
7xwVs21GjrfxoIvi1IPlbyo1wZnjAyP0MJIJqKjnszX2thBG86lmNh3OOhVYZeTR
lRvXDFSXQyA3s6mWIAEBTEiWRsy517BO9EGqD0XcyPrpeZMmsYcixVaIDVQAkd44
Oa8+PHJyZs0Ijwtc0TpYAm8JiE/4dPRAwxuhevlK8+lzZN5MJ+4DtzUhWG4+c2vY
rdvpKN4sbhBQSeNxwin+dhGUVXpwBxndbWY0dJEtRRsx6vtJKV8rMxQpjE8m2yMx
tU+h3ne7XF3rcg7+6fe4iWDZQsn1b44MijLDTCarmELO2/hBN9hyQHARHQq36G02
9nYVvP/o52B7ONg0g5ABRgUrVFiyyNYJ+rWPVJDCGOva0lO3R6JC7sR43zKrCxPh
uTVzWrRjSozXlhNMCIZLvACByDoFPvRtXOiO2tjYC7RvXXU5cHqu71S+v9PuO8nS
nzyVQrr5bJGZkg7yx4LtE9D4unVQJwStsYj9DzRimt0BWK5/gEsy1HdtPtBhEbC3
D8fXC3Uo4h4LGKUsxSYb8dMVnE/8Ac41rMb5CcZ5oHH5RVXKJ6iZRq1J+ssZe0G7
+Iz5nU6/V+ecWMwJdgJop2dpDNJWO+I6tLwqI05oHK/IAIOVfJeviyj8E4U7aWet
TvguFnTpok8V/xsjxG4ArNLiHMkBgFQKWIrqYJIGdWl7vGHAI3/DjkJi0qFdG4EJ
96yXMA/RrV2RVodlEz8AHF9H4iqVtUNHUeZ7MjZB271r3uUXnD5Ap1HwkHdSX+FW
NGORPl/PmQMWpwX2y26r2kTV1BqwaESKsTDbAaWYcEtn1FdVvBkTypXAbl7LuaMq
tp/bHToDMQBdfEDOdY+yiDe+cd2IgpIh99qIlqrBzRfPMf28K4ffQ73Kw/HfCVTX
tI/0rIhYA9dROpayrvwt3fzwGXzyRNsTzzKASDZWBYvQnaoSbzrxeASaF4wHrMSr
TCrjur8XlneQlzVsx8HwcnT2vzcAU3JeO9jpkvO/e58InPVBFwkLvmerNvqAj2+p
v6ehkEV4IgvaGaxvAxTbrTIpTo4JlFWYPzzA80KHrpPeSsJ2EmR8CdupwWPFcPGJ
eYRm0CKjCl95hC4MxdnrBT5QXpJDTJ8d67M2l1iuIwe9SvrnQsJa+bBcdlZerd7h
Y4InHhrL7DHnJru5fccalKtPEmYVee9gVhGzo1tCEFqgW5rmJiHl8qc5xNyeUKyI
EiqPQgfqbtD06s5MffvIwvv9ArIbOQmWCJ03sxl/4Yhtk7VMHCuntrtWxaUsIX6l
/M9w1t64bIkNIptc7es0iWH8x2YBTt3FKada5TTg8IKfCHChRgRhA9AwCVx57X3X
Pv7yM9kd2oMLvwy2QyYrH5wYlwP6CSl5tGgggg42I55cVb9WTmM2sumduPGG3i02
jkMxQy08mn+eUzveoMSDqon/kf0SkVoajbnlNMGv/8WEcZLbDA7V93536S298F6P
1ZjF8GrjPp1g65LeqHaYfzNLWbjJ6kBLquLSGWCevpXl72OtTGyKQJkNCIr96H+5
6qxpZC/8PEEPRO13M2etUO3J8zYtcTLFH4KE9zaIUZbbWY5YDq+Qwjs5NDZYTCuo
gAlXWk3D5ogj5FAWI+0rr42YDTMbDlg4S6wr1NFuVkc9cYqAR5+zGEyYI6rvQoWu
gmfLNCD2+N1jAcBDe0SXG6pS4SvtR4LuK6jEexh4bYAO7bwK74cuyhA5gevQ3g3V
l0YWPIqRKoBRJ1Hz94jMAay44rTROF/ODtmW8o5dLZS1LwNMwsWrLYeKmN/pTCNq
/mgsk6AlLfLR0CRkDM1ZLsIdVmWYoIkOITJFazyIYCa68UMCuK6MrovD3tRChPjo
+UKrKcvNzSA2gmHjl7Zf2g3NNIHYUNHzETY6UhE3faITILzmcof3ztpbdMJndOZT
MnnH3wq9KqQE3xgwALz6wLjZ7Hb9VIyDHicB+C79dwsC2Px2x/QpjhpsfBscbImZ
txEiin6rBfoHFGCcmTVhXGXJEJMprBYG8doB0q9QrmOHPxrEWTX/F8i4Gd9f2T6k
p2/uABTQEfjlTpU3UvUSNROGkOwNhd9JVTe4u69qRd1nrOj400t3vjNCdCWIclP9
7kH4ApJ46zzuuh4ObOCzp7VgeA16yXbST14qcuZ8NxZ/OXztEt0mSRJqCEO5o84T
x9i33KFfz9OqIY8Bk23fpY1pl3nFAUpTQ8DIH+M3HaeLp7O+mnNmeWMM+ZtCc1LE
Ns+zpgl9YXSkTzN54GtM7bDdLW3/3lyq74bz0NfXliXvyxHKvjDCIOoLYg30mGBO
BLCrVrJI4ApSUmyHSQsnXQoaoOnxBt5jh56Dhz7/sw5tBQ6flkOegXiXGvTFiMVN
70ZSNsFFy8KJ3WJFLfWwOdbWQUYST9j14JeDsWCg+tNgf0Xb5YqupQLjT48QOyyr
9M+Ni4DkrTeVzCG8y6Auja/7mJCOtJ0KfJwLqeXzxhUX0ZL+L8Qc7kvyCHqV3dHa
QtCKB16bl2gkPJW14VkpRafXRx5IUj+dw25GItBAra3yfFFUeq5RPuBX9yFOmjr5
EoUbQjfZQyQGgbg5H54cch6lH4a19chgOqI4kbjMzJVulPa7tWiJNBUzFVmahZ4E
iKvzfSY9rc8jyJzy+kSLyQMIY28/LwXYq+sRRHkd4zMlb286vdCimqyAQsXxtVth
/mT3UJ1oll+szotTxJv64afrerJexopqv+9/3nxoE3Y5xJU1X0F+pUTSUDA4QTaN
uydrjWoDtXV2TEWL7W+fh5LPqJUdh35ifzsYapbOLgaIxkltjk5q7kAU5033I3bp
wS6/x6rBH91xGl/wcLCIfrMp0nBJzTC1v19jgWKADhyoGlXESWIz2d4gZSTSX9fV
2IpyEeUDErO8IFZYp1keIfKBz3jN6B+XVGmw/PM2WxViJdioD8/M5eTKzMXVEB/7
SDCnfUkXZBJ7E/er5RptrEgg+jiQuYkHKT/vu0ZdXpBuFhtDq7/VhIFbhZwGoZt7
anJWBYUhFcxwG40sQXj+PsYcJ9nTBewAhErF35VnV+et47cXDrtbUTBw44jpGqs5
UqsX5tyqguEoKP2B4qIc8W7demCWXnU7toS2Y/KBG0PR0B1RBNyEzJapdG8CWdQj
R+/F+XTT4ue26E8x1EwizB61lY2lpRWp3YzW0km1Mk1kAY/9tBzA14bAIQ12Osm0
XXK8mW5A7Qj9MMCP4HtlFlGIqKL6KH2mJ18fL6Jxnbo0nSC9PtSzEEIVvhTEV5Qj
Vvi2D/h+kL4LQt3jM+DOAUcQ6FuX14mQfrfnLP1AFEIMkZVY3ZfBmYFvnpo+zA3O
cvX2TW5PinLxKSb4J9yYsl74EgdvgwVVzEU9IUaLtDvcJBDJ5sP/c0oR3ICJSCUC
THIF4EemOAyANIu7Umt/sFmS9uey2Q4Qi98/s9elWb7wUBK9XHpFawpqU+E1f0nQ
5h6iiwHhPnJH16DkS6E57o1w8K9gNiLKwv/E40KuhgV4PA/X3ZunegSKTn2CXwAl
rTivVp/wUHLReyMCebNwpUCVRjpj5ScEp724ruheAN+L/N7z3/zVTrKd724NUYMO
giyknG6+bEFq+hh9iJ+3tpb6bB1trcIzqofpWld/hYzFJWGBqdWWd1LLlAVuCH60
qhOxRQBQH2KHLUG2ezNsIPr0+9mqBVmQF3ntULzgJEn2OC9A4KnRLf7Sa9ajIqxp
KD1e3lZvLseXWuJAW55oCJxUFUmwZCEY9WzsmpkOUHPedeh+Z28FHijT9YrbSSVK
AIw3QiFU0NwtZ5RxRDUHJr0vlNELYBy/UTGuhRwcqeyw1ZQyrsj0AU0rjlMeNj/V
qkk0WmZbVYyz6x4cm0vBsFEe9mCzcpzpaKkhNJbqtBuWa1YVHuDJBC/wgVAKFog5
ll1lWMvuGVoLuCkZdJDXG2uiWwEvV5lgzLDVSExeXN7yg4Kfjmy3YGXYyvIe8XCq
xCB7B+gm2IXe4JI3qZ424EbCTFvuwqeLpoBUjYsqGgjGrrpGJpBZV9CFb2tPS6/N
zPpQwzHtfvnMWmLzUO9yuMXKmV+hnm9eMC0BK5SvmlPQ1hxLW5NrNrBbpazNghXU
bbaXXxhPTjXDa3VkRHurPWZ28vgcSPh7GQNcZ3zvSOdqI4RO8ObVGo2CON9SPpZs
qpUHDpgd7RCIJBcR614b3msrjvSGmlnwIEZ/5rLGbS/9m/r3dphIoP0L8vrIoupW
keMfK29qLCdnwBlQh+Pu9wSvIsJsHCEVbQTL9veZqgc3CVjgCDv1PDpuOaevC1C3
ed6dE7Ot0kjusijf15YtaMLtfln+nD4atQk3Q0FvOfiGlk47FpXZbpd3YotV/fp2
84Q55BCXBL+1sTuYqEP5ntlAMA8mItoLRpjBOCBsUYyx9Zs0INNi+F5p8Ei25FBZ
Iiz8OY7MGpH6GEFn15USJcVsAUKBSw9LLonQDcIjWXCiEpcwyojBkjX0MFSV/yh7
PlK+fPMySCwQk2MATOoue9KtW0yxMfGlktu1hCHg7kQUXVrEhsr8CNtX4gqeedkP
fCXf2wIBoPyRd6mKqk2EHy07HdHOz72gVGKNm3oolu/VGS70vIILH18FXZ6xjXMB
liaPG7QphOi0hg6Yng9TOaoWSoT1gaOSTp3XkWP/fV4ugt8a/bgh7HUec4W5mUzH
W7LmP7+W4eCEsqZc0P7rkV8gScTRzV54Pr1UcRpfHuFqDe/8/q4PEckPgFZ9BVed
vHEe0g6uKGzG3kR1A0ztP0/p17SrY/TdGr33/ZHS08KGOhv0PHBckfGZ3g4GRgvg
0tiuNwhKKyxZqJ7xWWiHmsm8w2NQXN5u+Ov3UKDBDBp+9uU9iwT/9+rPaSyJ2Bwq
QynT8CqZ5llBj4/KtA5c4lGxknFZxhZAMLh+3zqy7zkry91ftEDQNGuAnubM1CDu
05QOFOY0+I5zzRJJ24te7p68DFmlML/s+PdDHb4b5pKYYlE2z/kBtrSCJut0OvLX
V7ogiqojNky0MDXW1rVwyl46nawmjTrGcB5bs9SYwdxQRuvKVP7KTZkngWXxcJq9
UPIYvqdJ2xE4r2AgTdmmZe1XvlLiO8RipnyAywGvsA6fBtaGeQ1dE7Vzb4mZESxR
lm9mv4FEYL6YPlquhsgwvGQC1l6aoh04vBmECecIMzD1QNETJRfZ2T7xCOcN3elO
vL5eFPzY4bWNdK836mzFYvFld9dZlOtWww4xbNp86MQLmV7OIcMymGPC7FOQZgd2
1e6xRKsHD15hTwbdPHmMFT8R0vQSKAq/FhlUKqwbIHDStTWj9YrPOLePe72bR9OY
MmIxbGbX6Xz71oHNpOvpj+oSLhyQ/taMaMpvcPTrjonKmMvHKj9iRrIkO83IUiXS
I2128R0+8QmKIA9jnkfowMvNWJn52Z/TiYXB+PvdWMFeljzi6TeEmbnwk/kA02WD
iCBHImx1VR0uiFHV/rXQI3o+B0Vwu8jmlJVfliDJs+4moFJ5TVQ4cfy76jKOH37J
xZvKSlvEfGQ3q9z+SZvC2jYo1+y5HcMZLiQfem477/Ulbgn5SmvSoniXPA/QKI/D
KxlMyvFNdWVDBgwJm10cw/TzyvxNgWqnNiBzXjElswH2bQWN/YCmOhw+M+nzKACh
TXB6s8Rg6qszdAf+FhzhN4Fv9MHk6tnDqYPIvq5pJxEkGsIQAVC/kfY/YWuHVQ/r
V1Jd+TjsKeElELZ4rNcy9XsyuMZtI+5YSK068J5f9kT6r270zeVzvjW8GyuLHR7V
yb6wU+q9wTU9QPAHKWRQDCPo8CReUa+g6LAEddQ3s+bUnhVhg5uWBJK/kdTj4TuH
uqimsq5vSugpdvtjgcXYUTYiKmGKcXAM1Syb3tcJpoytXasQHPxWaM3PUnBwjb++
Ufq63ClkRwx+gDFZQyvSX5pRCVqAvLFVftBzlo9K3ykqdYIRnYchMNx6Se3U/Fvk
uv6ZSsh8406LzmAZh1DfdUloaTEA4rhmz/ZaTMipO9ehvWEOxeZj9b3vkfl3YrUe
EmczKTGLg5O7hhxvoUn8GTAhAF0j+lBkyDOtTBxPeRfXfI/fO1lwOx8rXFnptzpP
RgJ9dETuxCfYjexvvskTAwb7bH30CxY2FswpMLWCufHFQMchhLLMRe9o7q7jItjg
JXBuMZkTv8eNmzEGtNQz+2W47aUhegPqjV4M4b6s58h72jPXgLFpUzj85inxo/X7
Kss60gBEqjhOKKudKXIWvRt5Gk1ep8bYiMUlzwSfCfm4sAT6WSNOZOBkypv+b1dL
bArgYdrm0F08tj2CiuBD+v5bRhGmgwMZykxTtR8HMwTIezQhibnYs74W4yqYLEIx
HI37MDLqZsA8k7RYdfAE3wFAlIWMCx0fxo8GwiMk5S+FL8quBmDpt2MlR5Y4ykTe
3CN/iVOn7E6+TKAuQXJSDHqPDvRAqVwLq+sGqhhysqrBC4FwIKbqunxDSQY07CzR
IRtGkH8EFFxxhAGHmo8YOFt+erPCPITBJUR8ROtOZb6U+0Ki5G2OBHsHdjgZV3te
mJ5883yPZvkdmqDmxj0qHFl9n1tGSs03vVe6pbfl1NDQLwr2wQEFMdAY7NDpVZZV
liQL6JBEHjSMBNl6t6rFBhtYpZ5ool36BLD7CvYAsZgTc+gfYzME3syhBPxxQ0K1
yB7qE5XA1dJOW2FZXuozX71xbPdr0u5LoKoBldxM0iAVFjgkFvENSAwCh+fG6vyd
BvsINiwktjgl4rg+JiT3MXl7PC9Hf6OKL06NtHVHc12mZpv5rJyeurFxDMnBYEaH
IZGaVi1mPaTi+EHcYf/EsodOxmvhciTevx2IlQ1pXmaGqycpZrqBq/vSA7qgUCNA
cAxia/sX2XSHInlDNIAJ4sYUyMOBA7tm/L99IkwOK7HBEunxoUfhI9vCAsgWkBW+
QxhjbysbVs4tcmNt4xbWuCT3QDBXBo8c+QzacjpEilEcKLTEfNRrrEFxkco92M5S
nCEk0JQgLbUUz4KRcpYnsJDxl2Bl+XHL/critrLXsa/15uIVzWPe2+2j6mR7IoDG
qu4mgIxmn+lPEsgpQu/GaPyLnLiaV7YlcXK/mBRVn6fRflr4rulUpiQquYAk+BaI
aSX7ax6b10uNTdGjp2WOMZR3Li5Y5vWjCeqyGjKrbKtKanfIkcryTqtNynnmTkaq
fWFpdhPxkdX5SsqbMsmHXm+l+4oediKSn3wP2uGi1LUcbgrhSVqUG7CkWSpoQQF+
Sm08KWDGWAUuS1VsPq8nigFa/MqPQT4+B2zpxuIEqnsM4IAZwNanDE+bjdiMVqkj
BkMp0vgW/R1asXVagYbLtJg6vZKM1smVjUnHZozVg9bWvAgMhKC9zHR+HJbV7Udh
n/oTc+rY2Xv6fjaCbHP2GulFhbzV5TtHF47ibalxVh6yy1mjq4zZDzHPWIoUsiWQ
SBxwFWgQc0uFISGIt/NNQlIlHhRi80f7mtthrgGwkzqRDDShFScDiSSN8+fjFkRe
5ClCj7tvmgVVj86FYlIOlI/r3hzofLf7Sx0sN+5RqsvjY0hFzVG7AUl3+BjxI2kb
OeHB1/pkDmcXS4vTXbrKbz/7zwCyHiRhLUOJIVeJFJYJV0Q6A/NNrvFckKd+Z01t
mZ3VGSucz2a4lU9ZmxbmGdGTiEZLdQX+/kY89j8uEnLJ0nxKhhCXgNitXDrq9nYU
EDCByeTdiYzk0QtWe4M4le8l4N/1ykqJ3KY5FBmbgu5LFiBJNICy8bL0cVkXCLn+
KS48lpdisBrhz4eouwL+uXsqusPfk8uV1GEVJYDBeV8NzonxBOxK4rNlQtVr5Srr
Fl8faAbG9Tm90D3nwhrN+As8oXoz8qr9squ4jSHEl9cM5D0J35kGAU6bdySmV4RM
+GKFh1o2B8Ilfp7a/5pLSliZy3a2l6VneE0WS8esgVzxSeAxJafoiqdNbDLtbbpR
zJ1QShIcJbfJj/OkIq933X+o3DocyW7GKnWd7S5PSbu1FQWdn+ttDqofmU4tWaka
RooUCuqfEAuK5gEa7bdSpiNs0A+LYB2SrrlYQoo+47eXDzkpQer4f7L6KTAepAQb
Cvm3bUMHFoLGHWQySYHXAOt5+YRlbzm1JzN8kVgPsMU4ADCaDbUqWuOM+CWFkKnp
WUMiwSZvC6FAjgzYVQcKpJLgJO8HlrXEAPo+UQ4EsMMKv+X0ZgFNnVTfY6HgY7v8
0qP2ZlQBK1vG36xMm//LmuF7pdzYZfnFrzHT/dMWtdK+pQzK2onOqV8GabNmFq+H
icf0eL8n6tI4oqVeEkSy5CLNjnBNOSVgt2kVYy4UPBWb6GEGquCU/uhYd/dBR3jK
o66+PrMQJg1vvhW9z/mGi8v1H9fNizEblRuxy0bl76IIDe9TyU04iMunAS+1GHk7
FLBqVV12SLL5+APP9GDdS5uGMX1Yfx9+EiRUoK6ARqEfVuspAgxz0KghmOzeIc1z
LnbwRIHA5vI6lg98Dfpl7AZ0sT5+b5wsTsJjcGlQ+Yuhx0eF2we3LJkYeM8GsZbh
0bN8Tx06lGFLRhyfV41JYa5MXVJq/U7Q6NR+6DjgjUtoM4DarzBtIpPdiag5XYCZ
XBCBzYxgSF6Zesf2UEr1tH2gBxHnxuEjlyrVevcM9g8rc9rr+ZezKItPvdJk8DtP
JmwKIiCJ/IQ40HKc7y9Oha79yNhpVw2280dfIlwJcJjbjw1tL2EXM31PHz26u9+g
DjFpOdJYVylzBhS/KO9YbbqRG5Bmg/8iQ5jyTA1Zx4csHj+XQPlwFcRtf1p+mwyv
qeSnCDkwImkcvPYw3adFOIk+dxwWyQ7+Z02F1imM95/MjpQqYwjjlnEzoOmtXhww
0A4BUZRru2lt4nwmsYhLYz7YARtbqg+UgsemWHTF2iIFdGe0vptj280Mu9WP++YM
cc3wzEzbtTbNrxt+IOh6K+0PXwSmKnq8JnYhCohtCfDZ1QMIn4z80rAJ5FJPo3If
91vykpXv9abJz3ZaDtJEac4fi0oBmv863zD8FBFoFxcUMDSv06ItUicrDqJsDDQ6
av3eJch6tALEpJL7r/b2OhQH9Om8X4BIoNzcvrtmVJWAj3ObjEN4cAYyuye2rsVj
JeARyPAcBulu/HhVa6tfh7+yWdgQUaucHE2uqtZ7amARTEN82kv5HQXmh/gRpbei
ldT1+zGUOJZMyktaKElW4DJB4zEu0ntsi8VyoV22L6QsIedcmjrBxNSotmCL42nS
sPAuEIWkG/dHdM3dmEPc0p64bIuHc7xZrRZOlAtKUa4b5lP6DRGAVnrokRj7kYb1
3FE6QKa0LyX0+tP6iwwXcghob6k0hHISbiA2yV477xetrL4XdapHX1MpgyTN0K7z
Z7V7sdBVsisk9pkfu8Qvw0QTvm0Gjcxm+bVtpgWdLpDdzmG+Jp9beTKpgwxOXqde
oB2Zd3B+w91hQ60LEz/FJr9zZoO8GXREuoosuZSZkPGOT5Vc8W4i8LCCSJ1z4xou
FRGwxS1ulZJzjwfDfINe3psWIRRfq6DYqOsZVjQrFQ4JduHIEIoqETgJDqVpr7Ij
JEBS6kAoqqDmXDX9iZmUvJFpdojF1eI5Qxa4113U4BNGYjVs6BYtPjbm6uoUi0Wx
WLxc3+4ZBye7r/MfRJNJAHkoxYbeLlXVVPTb0DloPrvV4y8rqdnIXD+5eq/mJX5d
gQquxMiGvGIWReohNR+scGfk68qbx1iE9ubDMMhsl6teTftr0w9oRGEfEqcV14qV
D7awpI9zNV+IqvZNe8mHDOH4J5boHieRSQRNAYh3F0WPZXZAp/4UAivCBHLyE3SZ
lfC3HcGTXsMMr3vXv5IkKVV545DhARE7aMhju0Bcksa5k/clgeoEL47YO5vmkarJ
8JAlK76vB7E3SVsyjtKTv+6sKi/UGgBUbpUWvuZY2nEmpCSvx98QAu/zd2GuSLEE
XEGOx9gHCN3rh28PvcVEvVjgbFHrJF+UXm0ZErLY1/hgFkmP/XMgZjBnun+P+lQf
QkPy7COAi92fuSk1EZssJMrmONzTPJvuGTnkFIue3BItlQHkrn5HfkHBwgaLKEF/
VRbxb1ElQqlm4OpdcO5pJHwFPnRi/b6+Vd72FYor/rZwmPt9k7FSnXMMUXlHFgbE
g57NKOyEF2Ujk5IdGRD8Gn52whH3u+vmruMWjiwGD8XocQ6/yRimr7AJ7wWQuURW
3pV9XEoREW1FUIjrKSZhHKODrY1NJ7CLNaRRA4i9FZWWQ/k4WLGM7Zc4+LtPbiqf
UgcZLoJljBSuBBDL4KGK0yA3Wv/Hm5nv/76Qw1ySaQTd5+aMGohpK83AI3IXyiMm
x/s4js+zRTmNrEyd0uCctBSH/OCUy/jDxlNyQTqT7A/aCjvewIuqwcRDsNVWoL0v
FY/qIUyWcvxrNYyjPDWfdwRVCteGwkzJXPW6hf7rEic/5591QX7EaVK9TzJX+zIG
GMxOrnbwhIgIamhuHOq1L1JLkU63rXfKYl0/35b0YatbQNeReGSuLFWJuLDmB1j6
5Uqe77b7kATUay0JYSfslPNpp0/OgAy/N8Pr49wGPUcmMs6SaFnD3slLdFGsG4Sx
bY+Oh0M/UfagnPy2fdqVL+mQ3E7kVreYjlDf4rPKL72hLGQOPzt649OBLYcfo0es
6tc++Hb7pqteAtKUhxLM1oo4Z8D0EiXncBB1hhIOYrJQgYQFsdwLHfoVeNj9SpfE
36WXMfujft+/QNnz3mLG5l02jkBRl6ux+FDlB3RxoCSoQE6CxDE19kxXjW0FqPU2
MI4/R7b4tIipgoxdS/O9sWXGsdBw0efq4kQQhomUYEGKfK+p2K6v4bpQa/CSDBfm
N5QpUPiANw2LCwQEW1y1U9XEkBd79P50BEcGQP7ss7JYy+A5VDUVmqCTYefE1ucK
M/f9Y3oVuK5YjlG2jD1BQtyizAl3XKdaoY1MWJGvH9bdf5eEjjcb5hCMnRFZqRWS
vDF4bDjYjAs7PBjDak3Gl8/h9Nj69lwunA74mFL0Kc1QG/gQ+hhbdaJj+cq4bMsF
NdjUeOGBa5saSftvx20TVZoh2SHwlKjCeuQRnX2AXTgGpXPKq1JCYP4JXkzDhxhQ
uFm5pu+9jrDJfmJe4kuQ8KyQhFM5AGgqbHuGBijJ5tcR/D5nbBVvgwzY5UDVBiGr
rL0vV/bzOqO52A5e6NiIE8DM8pJ+TKsgE096Tz6MVqIGs7H7VIMzeJvBsixY5B4o
YnkpE7hIUWkVsD3+QmYjm0GsYFZabP7wq2t+GeksCMtQvyJ1W1bu7YNFwXWLag++
k/gwt9uGeL0RO+M6W1hwuS8736fKjH12YSpA8bMG8b3AUzFtFzwXfQTqfMed1AsP
nll9qZZyg1TE1urqwtz7Il7AoAU0JqVBSU2Vb/IYueBozFyGF2v7RrN9KAT/7qrL
teqiKRTmmWAlhUG0N+0qf05B4dQR0DPun2tG+C8QuxIDrIDYAvfNHJk+e3K9Qido
gDnDK2ddJ6ASSKC6xGMefE6YEPMcgTme9fd6ST3mo51hUlHzjt+O8ZXwZ1sx7MKM
FbMilWisKti+ambkMiFAqOLqehFeM/Q7xo2s1vbO4N2Ynl0AeZAs4KiquCrbfXT2
AKTl6+bCjfZ+QWDKgAIVJ/L82wUGG3RPrVzv5odp+EkexO3utzsaJP1P5RhyMP4E
9UY+JjtHXgEdmdkkZTHCr50yswSu4K++vZB9s4euZ601e8OgjR2Y0R6ei+nHGI0x
T2iReSDUJkcN64YyHvzx8yVmAH+BZylaxAGJDDeFK7s21yvtwDp/qGEZVLHcbfA3
C0TZO1Anq6eSyS47+90F54LPKZHzaUDCCRlu4JeQ78oqP3GlMPZWoyH8Z8dEgTBw
yMos1hdSIQGUGTph3cLw1NCbBOulNYAt7zsgmesgxaIK6AOiiTIxo8ZmcFOU3t18
4SUQdHC0II6D8IIktB/rchztIhzI2m2viTbNBFxMf8matKMQkMZQlEozNQtuhn5m
nTdGe+S0UboCp+eAjdbJ+3+tmh8KjDgO93aP0xgG3DWj2MpfBMUDfbD6MGb4Vt13
npqg6vzn3f3ayXnjehFn2w+DImczmnSR6YQhp1bmhHbqMgNRsa5s5eoYGNROH10Z
e4NZ51+ZmMWFQXzLlcAegKMCB0irvCUpr2Sulr+sWZB1P4FiN9ug9Y285ajyvnDF
hr/lX4TMxQTpRykeWNtcp24k9tAfOPdyEBhsh/LYeAY6McA07MsYZNrWW46zm66q
uIIiZon++VOF1+baSDCuCbrck4n3/lehE/TtXIzVc4XBiGU3GFhG6zhGi9BefNMx
6z/I9a7ZIfmZvA8aTTQ7DjIq5yciUIXla7GyZKQmE9LmAooYmdTPpu5ZdujTv6ra
Ms1Pj7ZWKMjh5VeAVKFJ2mzEv30A6eESQ6QQsAMa3Zd2XyZHpGDBSbYtygbNcr6D
ZO1NOKib1fBPwR7NGQffNemmtGk2kdN0uCayFcX3L0T/lMLM7F3mu0VVdUZvWHfI
mcsM7aE99UypEVsxf8zQcH7wXLPamMo9LN2C6S31Fjeh6ioDUrMSHwM+Hs35vXpz
tlzZU8DwrUEVamTJWE+42MO9x8vM4f33hr3FsM/76dt0mYsL1diaZRg/aQuWRfjt
ChrFaMAZ0vWLPPk98drqXaCevgWj6tCo4W6RUvgc5qmahMH5rnzrVorisIaDvQSK
lt1eb8fuTC8A0dRgwBZi8IM4TzBHDg0AXRhTjfrNGgMuBfGujlAtsIOnzijQxOAG
vMeh6V0ybiNSPxoeWERFZpWNzecjmTue+WUrJihM9PRppEXIi3Wc8NAdlMKp3MwX
7VYazpB49faivxgCEuSggaTw5ILbGsfKsmHBD6gBzXWTfRfocFofy00s6UIzkbCs
jsbnoaoCiTzCtdwTUxZxbe0m/CY9mkyGdn/F43ykMqgNgxRV7Klo5MVA898ZkwI5
maJyes9KkSUUq+De5W4EiXT5bRBo1YYFHUkLSlMDc0vlJEEhYKlGPSoXuLX1VK0S
yaswR/VKaC65eVOzZNljne5YwvJxmlGkob6L3O2J68pQpAJV7Zz6hoiC34Wmzum0
fqO99tN+6Uh0K/AT4Jf5N7yajX1AQe3TRl8O7eIxPDaXo+w3MyKzqlsmW45J4XO7
vT4QYlkv5jJMkZfElwFte9rQZuelK3Z1AeQPnpxtOY/y32eSdJ510QSAXQAw0dFv
wEt/LC4KqO+OMb+Q3+3ThZQALK42V7E0kqNPlh43gsFb9ZnfWFEdp9o4V/MDmRK9
NFyQubSC2umrNBua0el3Yycvy8CKdQKvL0UoLTduImqbNfGWuujWLQNXSoaklgjt
jlX8bu2Tf8FsIWwvD/ilC4ucywS8Ammt54ixmM7w1lTtyDyEBas8zkzNKXnGyYZB
vF07zBAYbGVZwW+IsjB9p1D+KVNhMOuS2AXrnqtxgKpmYksmXaFKd2QhYAdEDsUb
6EGyHXvS08jkRvL1xuUtCZK+Gh5jWekH1QRQgzd5LCiYFrYp/gk5sZcKZVMFqqp/
cYHJv5nXN78RgUMFA8FV2tKUuY/CvA/aW76yWIYa9nOnqBFYX/v81EjTPi1AhNYy
8nT/bnXSUhW/Wglb9i5YDUT+SK0tinYGMnS0h7NnUqaHY/C4tzOoDcYmeVvx7TNm
AO8sPyH3/sAQwHnSkLf9hY41n5q0C3pd3+8RE6OaYdW+PoEVJ6KikPOz0i0kqYXF
0bQbKupKLkAZ3b1nK1HeS/+eKj7EUKJmA1AziIpeQLJNj8EW4PKy4EreOgHqkM4b
IDw0IWQz0wq3nNdbSBzmy70wOEEiMTXw7XovAF6Ai42yVnp5yvwUt7XjKjcFcVia
dA+vF4I9od7dIpHpG1YRipabHM223+Pbg7JDiI6yiRVDWc5QnYBBCgMtKY3QBsaB
KLCAKZ4reWRM712orDoztfkXSVHspgb5vYK4eyg9jloibGSNcMU4Kfu81z6Ps2xx
NQb0iO+kgd/AMtfAvmZVggJ6755qp/N6sW//E/dxrHBAQEAsbNDuAuvvYeTGchmI
k3F5mdsjv1GNEy7c76o+2A8IrZOj6cjvY72h1VRTsyxl5vpo2YVIGe9fr8kfBIFW
eWPdr2yYM03I/LMST/mkXOoxrCEJqrxo4RUAn4X+bhsC6GCr3FniWFFDRTPNZtor
orY6P2CGXmqSmp+5T++06M3W3PJqsN95xZBiVB9sl6o+oUuiHG3pvDn4b9BUDtBD
0IaU/dKp8wgNH+/2ZK6jgNZRaYN6Q3BMHVQtf/Fi79V6v5l/fcWyduHVfCvv9vxd
7nCl0yDcE4VkEbIpYusXqM6Y0xqz8rxLXMFaZPqyTpnCnccR4uUOHstZZpqn9jD7
CoB7GgOWNAU8cFteBDfBAy2jPG4a/ZAR09kqiqtMifUd97K81la84xCGgTfb+F/7
4HSHokoJmxhBXxQfKL3zmJJ5iAazBqZuaJVE9Ox7vxRK4szni1i/4xCz3EZ0Z0hi
k9xQFZuX+aJQ6lqIKifRjdK4CPllFGMeM8Vy95iqta1t1c2oY3TZUp6AYmm1TdRn
g3K1QikpHiQfG3FWFwKet+uXMRCa0YXJVJERZnYgOMY4bOXjwwAB3wPo355t+3sJ
Mi0KRDh8mhalXj7LpaMUmiORPdMtrbDsCYXnUNyX3OCC0RTgZY41akWcZZmtsyNf
oudbF29i1qa8VRRLlKzxdaOZlF3QPxVKjoU4tI/z8XDcWF53HgTDNuHTzor5ERA2
WH/MImSJEHuqUYwf+NYS0M744ynUmA5HFLUcUH0vfRRZZN2DZjWhvy9bUSXu6pOH
Vmfe/7PxPnvEoVREJ4hqZInDhpbVfKmvu4mKSGrGZWd1zE3quZZYWWFu0L9Ohusl
s+NojTtGuU/q0Q/yoJZ8cKc6kaZMiDlei8ySt8l+8Ter/uZlNPN0qhash05cwcSg
oxQvI8Tp9LF7zec02NIyYMVqgvipEeC48b459ZnOhWUsbNR4UjzSCPXGyEkUC3HH
BG1QWMO3oQJ0VOs4hDb7KIFTAXWfXDAPSafgOqSX27YAtHxR0A5FqlHTBaBkX4lt
ezS6q9cn36bG9sXaC6X952F9rHw6cefq9P3fwENUmuz2P9bfwasEx6pCEvbZFHUL
mdAUZMjwcizvF/WgAchJU/G2JormqKV/KMJd0LRMGms59c2wYFSyakoFlZwXyhJE
AVIdfsPXI7QsIOJixiX478K4V3cVpriMw6ybGXTX3SKlA6l8alBt57T9FQurXjSC
eGtsz0okFOf30+X37eE6SHPrHVM4V+fOYOD6OevcOc39Mn6Yg19Z25o8zZf3QmRr
nviQ+S6HUM95dgYeGzljDOeOZQXhGCMFCIvgN5vQj4IxfpIBazxC5nqK1rO6FFQS
y8m2kaef9ebtj/9J392QCyoU6Pdu4JlIvznIsDZ0VmhwH+RMHAg/KQQwbuF0CAyP
WAJ1y8ExlB015sjHSUltb5siCbHK5GY/oKIbDQcfs6nO2CKlKrwB8r/pe7eKvdsY
BSl+vstxBQX5FffqPHtWrrywfc6BGvZG8cqI2hoWntVdmUA8eq94QRqTgBh1gsJ8
wbJTsigVJ5x6dDtUjm5NXUQ4Ot3psixnZgwzghNwapFirnmko7CX6sWht4AyB3Do
2RUCs+U3QJBmHJ853WyahdZDDjdKe+0MoZglJO13QQx4LIhLpImSzZuFH4fjP29/
YFB/tlXDn/AbInQEgm6THCUoDrktewo5Q/qlOFKPEgUKZV1ukFteeRU6FqPnNcfk
Jjifmwo1im+0LpyIHWTv0HpOFejNVRVITuV7dYiBjeTSeKD+Zm1UIlEnMj+clQ7d
6iuM4OzYIyHsrLcUaMjlNrKK/uLAOMqBPg1Ue9EKCsCJgv3K9XnKAYelLkAS8GAG
T4FrdkhLqY5EdupKFlwLikRNlXCqcToppUyh+GlHFTQgrKkiKY8d1DVCa3dH8rJj
3ZM5OmRg6orAgIy6FOIELydxlqoHPMCFbfqF9WUt8AY849x6DlPZZe+rwNTT15Ev
ayKMTtjek4Tj7NdQt0iewhZowlsvV+i0fXkQID/zb7ouvBTYxEDTZrIuFckTXoGf
tMAB7lKFYOAFax0mAgXL56PsaONU2Rg4n3NxfH/gLyvEsH1nYKPqppNzpCepCLxK
i4FLQaT/UUxrAy9jtOssI1pt0X21ImBXScQz7bhzlsaXmLKW6joIH5lms7vLgeHt
DkGeDpryeAfvHcM3Kq0DzPgEOUvjA2ZoOygqYH1908wArtVIdEHnxEBAy3SfV2+D
D7qYPQwD07OnEMoT/TOhvWWSDFZO7jj9kWQMb0bGMdCV01YzXu7rJcrS0HgGi9+G
SRFI1hnp+kMA3ADCy+y3HyoDPyKEoI/ls2sP/wFug1jbXOMT57hPOooEViBX+r/I
hbdvBB43PA7IR04q5sCp9Gag0tZhp7/CmPyzAVmpVaGnPkBtfxdLYmMJ9Vh7YIY0
MKanT5rZ80V14yMmsZPVTbPNyAdRBBDrgW25NNe8b0uQr8dcHMVbn1kYZplUgijm
M0BPiRa9/BJshQ31FvlEhsmx9jkQaLS9L/WuFS/73TtsyjhTMEm+bCUiGwhct/UY
puHK1LC1s6b/Bt6XBca2j8+Y7E2IDBwV4JrNrrfs7+0j3FgRLBpgglMkuKzze/26
LYfu0psPg6IUpWURLuuxyETJF1MAs3M7uZgcqVeKm2lrBbMcV9nNvax2W82Ed5rY
h50PyU2WK+6LZNXKmwxRGm8yj/ebpGbkwPcI1vW47xzGpM1JAG3EjCNYUvT7PTQs
lWkPoMIdvOfvQXUgDLd56ZrPdWIf1potC06/5bHX+2sJHwz6j3CoB5FW8P6Jp9lS
G9GP1DE2sm+oPqjaUi1Yj9fv0O/DdPmXbeKJtizQBwXmUe5tPNPqtPiiuTSyJUYP
xHB29NRnmAPtOUyR6nsS4Az2zWedHdReZPR7e34J9G0qAAZC859Q0LGno82S/s9x
2NODg69gr5H2m74YfFKTpmtO1TKMvSdfT2+5QkEhW84ZY+IuhzdCsXJ22iRGogRE
KMIfYhCLqgCHbx2E4J/9W9H7coVgSOoqSi1nuvXFXP5BG7fLrSq/tmAHbencY1vY
5YekbvTX2ekBiVyDrZLVxPFIKqNniYITPanyToPAciCTz/tdUKYRvAwMsBGAvVvl
q8t4ryM1YEKltabD5ThYPB67swWzlHyHfQMLMq1zQT/yOHnbiN1TD3vWjAHVBkab
ej+3fBT2ZO0iKeEff+pq7z5GJoxI+hdfVlmoIAPDDUFsdXEhRXyTbon8bgQg1J9d
5nfy+KF5TQ6+ZXYEgYk/DpxNzKA47WKk+hRZrBkLDX0MHldYeVtGrqr0xe7Gv6CJ
OIl6MsmmWQokctsIbtoQqOhP/HkGI3tgtNhtK/xhvi0fFYVpRuSQChGLaXAZySze
5AKuZZkPuKpBHW+PWxL1e4ZZ/11ENfjZ6D9Bv8+PrbW9xloWlQtcwlTdIhSov1Ez
pNUKQMjscOtlF/Y57E6QnOeAucUBjgNHAhcunGJridm1YCRHJ5Vrne2bB3zo0TTw
o5a6+YzOXkKBh1X4IrpJRb/pJv2xEoOMOc5xbKtoK8zkCoM5VKUuJR8gpHEfPts+
Y48yW/PYf5IXrcTY+7fO/dvFvwI2nWm3iYDNcygOtkwACvvr9Ym/lKL9Vp2pszub
w8hcQBmjX8+QWjNDUMM8wFlY83bJi9k4Z6+g/cu43/WSaUM+Ldn2e/z8UdNBfoT5
ylsufXluqcu8kCw6JIk6xfymri+jkkvIIXeNM4ipVZvAXxqlWiETHYPryner6IsU
80bcnPIhnZbdN9aeUCLrbSFKzLdzi5dYQqRZ86Hyd9O5P22hzbX6JfYb+fAbDSTx
Q4DAUVpUt+9ifExuQvmf35U0t3tZ6zeJmiNEFlvnUmp4e+PFISXU0YM/tMEsUa91
HO/9G3fbrcnfO6Hk0T2MUbTfYhqN+gtjCiWUwGMghXgRl8f94Tf+1SNPf4EbCtC3
82FZFxV0hTmwadgJiCFSehWTEZ5dxTK6ZGaed9OFd42y0UJ/7gP1w7ftFyU3kpxx
cq3oU2b6fUJICu/7Pseb8jU+eHR9I6C/ELbwr2c1SABwNsJJipqdhd/dvNG6zR0U
daYYQNyP/38NOvKl30fjDKhyBT9f+m4CJtRjVPZMW3qO28Bdo/Va01HDn++qnHMd
o8YvN+ZBRApIa9FjVPoEF7kWnsHDrTGbn+16SSvddy5FrPPE7g+4dXY8vg7DRNzc
yrxRAk2Pc6Vo+drlPjgKqJGsI+Cfw1F5qb+t8Z4D3YK8OwDPiiC5chx/nWGIgbJ/
rslRcioi3b7bCFnIOFbdRkt+ecg2kX3B3vbL0xTEm2V8kmvTUYte6liYFsBrBB5D
lXyCcooyvMPXYmHqx8NP9cXPP/tCdgWvSstTuRMKh1M83ECXn5joqeiek5u/Vlew
W/2aXqIIMwBy0hV10M5CFT0NdO4vqqcZX5wJqNHitrgVGDRCusE/9aTq6zCPyF2m
I+xy2/3UYhqo5E0QvH0lYzZe+3Cd+nfe1VGE4NI6hXHqORRU427dnqTlp4uXBtYA
WmykKsO6kpHfYZstYc8xJ64SN7ibWgMtNyHeggOD2MGrIJAcJbiw9onx1YOePubu
fpIqQp3R3FeZ5vug9ENashMo2/bOTYcgu8/q31xF+366jN6ZSOxt+3sBDVjtzbVP
B22HIlLzSsHSNIfa0sV4UKHL91WsRqiLnbTChubysHPahufAAmOO0KxW3zvtWfQ2
uNYXwRrFMXo3uB4DhUY0iGf54cS6oSAQbLWnJZ2NQGFHDwgwESETBkVFb+PawCOv
JSefU6JQLelLNhHuOz8IB6URERR8LWyfLxFthBK8iAWbVfLeG0HZlb9ueEQfQQjr
zEauK/4q0rPDUHKhdo8m6O8rclJQ21JoazdAYrUhWiEYe+lrCkNwo5merc0Kj0Xw
78VWoQ/vc/mY/iRproawqjEleMMXnigkcDET+NOLEnZOvEb7rzj4+ImYk6/8BaPe
M4d8sLff+eMHVAQck/mYYU5JkLm2Pgv9p4rUEVza7DkryYkRpJ7gYkZ8m2+BDuR8
gaGRpPERLDguoc/MmZCm5NJgxouOfPXkvYL3l98GwsaZ/MCW3sRxdrQAOHR6PbaV
szIcqzJ2dted6LwbnHJNNvsNH5CyJG9OTfaul7oRcCEZMDGObJ8Jt+8OyT0tDfey
uKBWvEGgZrYvTn2WZHrAnt4Ixbrjb4EGy8g6rTxeCdLyHuJx1CYNnF0x0JxWPWyl
/oVFemJOtPC4nXJlpcoK3TjLkPMqW47H54PdP0ueFpB4EseA1/sFfRono6YNMyAX
W7rizrbjIj1lbRKgtPBFS7rGrJPyKbediQFHoPKGP7mEa85Daywu65w2Wqwi5j6/
4TG8Hi7HzoOhOl2zhoz2t9KUInep1n6Mo6455XIY3hCU2bfYqpFhB/zP29i4MWbb
fbGHFXDz4O5XkAQpMN4F1YDONSGbtHYOojXqcedCX1UjX/vKWR+AZk+y0/LGpxNg
t4ll3E4TgHuTmhbeOzmmYlMLoVzKgD1iJCvB03UYTm1BLWQM1UQZuLMpU4QUAlXL
Z7JDuEYe7invu/DE926OOm0zlLvvygLgHePkVWCpdswAReEtkQ2SJXbBwrAIITa+
fCQ27xiyv+yT2dP6uxJSHmAUgd6kOV35nqdR3Ad4karu27tL6rRNEm4qgyGLkK2V
dTHfs+WKnFpr/A1+x0FGaM67w27Z2YwpEZQ4mmchlJebh6b5HZb71Z59XziDSKwP
G0v5exi7maSYhPp+o3+gq65AfXi1+MlsH/sYKg77sRBHTbGTM+nAnUzUMCQesmC8
59zNvO61+PCFq+xl1my1CEGT8Ked/thT0p4Fv3pVPxYAKWWeKGsM6sUlaxf1ZDJr
chqtAvs6AtE5Yhyca4azqMsu64oblj8itTD2tvONNzbswvjgG5Wwui1m8UTCvPdh
ct89WaHsoDVF2KoaMj2kF93LOLRoB+SRXlD/lUaAxUvBLD98usbLiJ+EWOtVRTIS
b0BVqST+WxaDY5P+KTCt9qqzQ33qdJrssIR2/H8idrIfTh/oRH/qEoIslrttfwn5
fjjAIHIvNdfcan0UhhYZF+FYH9DQlbazF3FwXW8RY7UpmC2IryzGOYD1hH59LsIn
bd4C/zOx8njuhysrbcs6BWzlOD57x+LuKwaKmN815wBqvV2HbuG/lTqu6UPJe8gP
bPnSo5bY0EiCY4WSh3NO0erMxCHxwNOhXCXOdatFSYAkSW5pnuK4BjrdzZewnJch
JvVFTMJU8j9o+vjEv6Yzzi0maLcCHM+Wcm2l9kHXPQyMhUFsTLZNgDVSd2nn2kzO
XETQN7PGpTiZtdkzUM13SAsPlqgYdqFlbU0u4rB1lMaeL66UGBeugxHXUacCc52A
B7m7LoUQDfw2ib8Xf2M1biRD6Z7aXcHi6cFZ0wxTUnVbZzX5dJel09KgUBFMkQ4s
v1Qa4Ul1VU4RRGBerbSzAfVu9i8lyOMjSEa3uHsQbi0oBcc8TufdXmZj8VkXd0nM
/B4ylXV8T1UYYttDeI6QUAwHcbf14P+97de61G5iE0CaNnQ+mLbj1DNvoXMYtEMp
f3rS2aqlCGC0RoIlmlnTGuxbdOJTYPJmgqqINTEcUdaTypuISxg4ljBviPliTWJo
wh6/MRn1xDoHQngXwqL7r5iz62gE9UzgyoIeZ6KEdTIC8paW/ZhGf85jjLNxb8gy
tCKl93qw38KiUIKSo3GoBNYNgu+IdgpYHo7alWs2HU7u1VgOQ73gKsdTDBsKKNWX
ifxK6g4/s4OQryZ6lr/rurnWlIrwo2Bre/7EcgvNgeyGfRtJ4NnmHdMMC60O9Jqb
dZGk55eGt+Z+p34dQ+iY/6U0IgRVl7BoLm3MBZNd+Ep0cCgZd0TI3fM+hQQD63S0
HmVKlFP9ueS75diAvzsmB89KBwop2POaeMtkmoK/sfTDilRV84WY4Kb4k7NOpcAX
s/y0hmkLPQerHIaLJKYJIP8ZLhqPnVs9xJKTSN8LRaA2uEC8GLSONltYkbrsuY/9
wjKA8OLqf99hNK/n62PtDVgSR4HDlr1MRHSME/Pvtjyhi6NagRYYsknUSePulH/7
IOh5Z12S1qdk/PEniqdPtrrfb11iixo6GhgeLAJLL54P+1g2C8LuzX5skRgI+/Cy
07M6JLrmy/nvVY07zd9Y7K9p850Jicc1FMWI4oWzb2wrtKes5IDpjkYKV/YOHxcg
OaWZPRB5+ScUTZLZocn3w6Be/E+Mfm4sPsXBe3u+z49n04oa1aleJwjJRJWWftVp
xKGZ4wBs6XKWVDVQY88YM7zlN6IZYkM6wFkIsg7swNjStmXh3ztA9mnU7InLx0LY
CX0+EGnhCLJpOnv4O4Zi6AVc7PkKy7ea5UYLw2bu9MJPpYEwmMlpDCw16aeEMXOp
nFquRP2hme/UFvXb45/ZsGKU+5tars3fHSkoloKWOr3f+ga6/GXfl2yos064kpMI
SoVp7IhhtyamD3e69eN23cgyHIFoHpPqTzJKBF7g1XYUDAPf05ATneRmhajP3WBh
7aqoDxEQU2sIJB7AU/tWXb04NAcEJE+DmpeH4lBnU5EWErWyke83a05Gn5qxfYcT
Tl9IzDuCr3IfSVAFhPK2JA31N9Uiudc3ZAAW1Q/GJ8RC6FQYxI9ZNaqb8q6pIjFh
qfJ8lnmNqrB9sQ/bLWvdEQfjzJbdRJYRRw4MA2vWASyGv1l/hCp8YUeVWT9zyyWw
h6tP39fBW43Cquo3X5AETLyA8WYVqrCxkJlNMF/J6mpEWq7x7/zAY3j2b/EIs18r
3s57wi4cxNx/xkWHqNBmPw7NDmRTbpzuq/BfwxiRBnY/9A7vK48DbH+D1F6Op6AL
fqzBKJBoLd7k3gaJa2WFd3vKSFc06lyhnHmWh5ttrVg/Wz5NrpTh9Ln84Ddur2/6
1hez5vubRFo9GMAxMJLyVgRa8TRilACdFYh62ZxjQw9ZYLgzWQS13royQlva6yYy
VvZTlvtFld32TcxoU3EpoKRv9YGBsK7HUjprRIDh0qsN4L3IYn+C0cJaPLMzyNAY
98NorhV7KAjEaHSXeUIUt2qwYJESEzUYb19Ve3Q974gYbj07brk/v65VWyPILfhe
suk0nUEh1N2kg/AGdNVZ/DpdOaiBx8DlDB+nX1fseP3GgaCHYMCtcocoLQcK73vw
ZLOIW+AAd1D63Eicl13rPhw00eu2ivPLi2Xt/GYe0aWBRF8rClpNGvbjObQgdM+b
jQMYV+qkBuajP9SG/cC8A61HCPaPwfom1inDk5RUTbENxg7NtqYz1DVMh2gnVXOE
Xp0aDUaGFjdso4PBqRHzZt97SBe39g52wE+8fSzB6lr9V17w4ZlP0qkgqx4Ptf7n
PnLYLsjtsjR5/uIw+PCJassLNuai9hB6nOoCLbMoZRdkA9bQtI7DZKFf1D1N1RA1
Dy1Ux3EuY1WMWPFLFDOQftkzkv8XQSaWqnFHoeZxQXaqYf3+1uIDgmaY/WXyFGP3
x1anOH9CgbfeljdBeFH5chc7jxelTi/QPSrGgSzgVC87kba0LlpQB8aHdy9BhTo0
55P5mfx3AEp9spz4ict6J3jTxgMaO7IXU59pSV5a4wHIe6Rg1O1+4VtOhanQx1Xf
Ra5aiVJn8OyAag/i0Y9ElS5ujwZVHe2BomdD+bdEl1kh+IwMPXmCmlL9bi6/1P0G
mo3SvZVRKaquOkBh7NATXPJBEO2GG3j90wPYoztmIxs5cTmH1bDs+xVGFEZe4B/X
qKWOMspK/PyNTpeiqc74+L7s9FwNn5T79yHUoBUT8CXvJVU5sHLa9rmaST6Bt3D6
FeUG2VEqko4zs9kXMjMoyMFlQEOtCrnhZN8R2NPVWpt4ZojZOy88dT6Ep6xMXC7V
iPhxsPgABV6VRg1zqbA+2MCfCYqzA6Mi6cB6VBBD4Hdz08RFDpSK4L/q/QWx6hh7
rGz710tkP90Cn3OKCJBMMYyjkwWvz54VF3tLnrnZg1zh85CsLOk/LnY7PVU9DmpL
y29eGxDYD/1LCvFCdgMqglCmmO4ZphvGoWSfIUX487roa8NKM/ReCX1K29CzvxeL
REFQdCJGuauU0kWnUPi3ba0n3ZnEb0iuEfYqU7JrCKEUb5NRT67wB1x5/6x9/Uoo
XHUQSfo8oFIH3D3G7SUboCoanejv7a0635qAmKpBH01dwSxgelzUbkc01oSJ9obT
d7TrSFcO/QHNkImVyB7zboTRerze9i6aih7kP8O1HyUEOS1u2bplS7tel91abQuD
PDJj+VNMYbJplwhyoB3tDhYvurPxH1ueROE8BXOmR9qDN7XUjMhj5pHdBRsION91
VFZdjcpAmFSNK2Hg31nm35zFDu6ViIAMr/zSMJasUMbKLF5mLmE27shKYi+AdTqx
F04lHpykUwwaOICaSIEoUx0O4KzWytt7X7f8JWiwRjTYMB12slAyUKikpMNSxaY4
4m1TCYFJBS/FeLZ39PRw1vQMHxZN8SlxH8rJHtEaakBUui0gOLwMC1HFWS3k0nEa
IlorMKVer7DN09qL6wEAjNjHkWbYNn75wX1qEPy5ZFnJKbDtVH7gYRHGPaP1J+qG
/qyiyrmdekrU3nJ97KfQEsXuOfqA1yK4iUab0I8+gdg0G8md4BNM7ZKmzkz8PFcx
+S+xuzfFs2NAfpi4okc6rtqaBVo6pQKxIQtbu7MLY5TLuNW7+7RMvws9iiUyfUGa
FH0lRheEMpUQOFdrdq1wv7LDwzU4e2WyHcXS48vYf91X+DpDCTlQyj1TJ6roMgpx
5IRS9t9Mv6MLotc3I7SIw4XgxTajoOhXvDgeiLjva9oOGpSnYP9GXvL1IlT/MTYl
8XOAdW8kK/UqXfZ3RLUwiwmCNBI431143OnsPBsY9vtlqfFq1RK69QECyYIXXJe2
bNOumUkq7hSNl4o29mgRoip9W0psIpWaDzvKALxlRRX8XdB+OcP4wl10aS9XQbjS
/tR+nu2bV+TSsaCxWr1etRbUk3yu4hIPG3QPoEDNIomCdZxxiIhMa5jbQ6WQgOc+
LqUqduHuf/tMMpiZAZpbL0W7p9wiL4BpaKsYR4mxj8CTSzQdfDSg5EyQ9v3+7yNp
RewhbGOTUiONQ/JnXmqOJcziBjQbxEMmiOA8R8HpuWSwgxTbrkwA3DPxISJalFpO
vV9Ma4POjpeDBBkQ8Cr3/OkxarYaJJOT1tjZ8uqteiwIZ1bDGe7st/8n2aNN+65L
7y5ckdtq2c8y06rL2yl5TBGuuII4ov9xbXZDI6PU6DZaRL9Oc77zIuY+i4Utodcr
ZtO9AUjznVDQbV4ZO4SME8TnMuQdW6PA3BL3zwcvne0OH32w/zgPtMSH/ZGMRr5N
Gh7LmmHeAnFgaHCePo7mfOmpvcEGoh9c9PeGYMj+xS28AxI4/44/yZ3UeMpMAuL0
K+JwBn1++VR+tfioCGDxnBe8kbnR6nQQneSor8YHa6OIFK3J2MwRxCdsZ76pyd4G
EAb+x60WIGvVwOGpYC6G34934MO16damw1TE4clePbAas3/agFEIUUe/IlxL0nBo
wP8GwX5Ziud7HfUpbsniymqe8PMHXhhoOabYKQ4CtXUtBCg6b+xm7WyUkq6hMDmX
/9GgCcMJDIg50rTMm0HrwXkuFKkwoOF3Qqnf5Y5ekdKgBxzDELDu26bfnOMdofb0
gwXgueQyK95VRhZdvEBDm/xBAV7oTCPVkz1nLflNDjRsbWkoTQDcIti473Y39x5b
4g0Z5viBMG1v8X94W/9EN5k9DkT6rHsy29WvKnPgNuWNYY/pJU4TdH6PehI8EZuw
MAWM0clFqBQPv93kDcXTKy4cYB4ZfnIOKc1mO7x7WRFmamcOC0Cm1N0HFsPW1OAV
2ArYxPwYu8D++d7vOHfsUmvNmMp7Q6oEonUOcgCnx+p9ZraG0Ml1bY3mmjo0tUPg
zDzLF4ckK/16co1wUHHyt/Fb2G5p9AD5GjHyXjeONQ6wwAr8avjYFW92TrmMxiJo
Ykkvv6StyKQc77NJnOBBp3zh8y+VWJhp8agQDCFa54PPlIaqU2WnzUy4580naZyc
Sd3IIy3WCm/DgD9kIAkhnVAoxvTslYBhBXRRxpsUcB/aLJjafK8DGfV/OFaHZrKE
65A94f+Y6z5L2rlq0lhM9lHur7qQaN4wRibx6owIE+T/GncarN1+8pI1D04VFHKw
nnFr311bdJn3X1429l67MU+xnH3FVypGaMlJmghZLcY0sN8EjS0mGDEP2h0mgx5M
bXkBLLAjAcK3JAlTbzh2qPrA11V+wO58LTm0DClT8+PWWiqI3Mg+Wcwis4HOfKNE
ALFwH65z7gCkXq1DQJh1PP5YEsSn8Zh2iIpS64RVZERYEwTs/eWylvYIAsfGuYjj
U+U/+1asu+rpu/4q++x6KIq3aYxTsRHVZvMJ93GbF5tefc+EMg4gVql8nIkL0puP
zTm/Obez5Pqbd99yp2295104tajDu0ENxtB3+6Xz1znrUBnv0F52cEtYU98Mlq22
/RRV/UXkSYhtiYYMMAzRuCCtaMNkTV7A40euSeAtCW1f+ik2oHn6mpSv1owhlyto
oNX6xOeLaS//CeDx94rh8KaI3nYvoi3rAcgQbwIXiuip+t1rQNUdN/VnWA3KpgPH
9NeaegC2ZDJY2Us5DUuUbCi7A1XCnC//voV2rbZfuXD5nZ7N/zRptXdOaYPT/Gtl
OO+AhxR2JwsO4zPkJVWt2PMi+aQ18+eBWPBe/5xhPDtKZrz2W0aA+Akyfk4CnVkU
n1qY2IBaCjHX8OPCR5E0dqQNyq+alGjyDFdrHOGh/RNyRABsoC64NeaSVAsRFbLU
kVetbk809KjihsdHscC8JfkqReNyGDZwQt4YhhHJOIwyIJfQ3+GVs7ODKqjNhN9+
bV3xRJ+Q9hdZNyaKVoBLgoago4/xTcYRCNxyaNnXYEca7kI0XgzrM0KJv38v4QsU
SNjLMfVSWouFNtjyYZlG5enpc/yrpxHgQUx1g8GqqoV7rbkbURwtjTmZwbglbrGo
p5uZrNn19K7EOlbQRpuuUT+zIdPeDDJA5hlkxnD1FI/XnDGksAm0qz3yjvsY1aNK
SzyM8UvJxLUPJPoZ5kyFAwlLXmRIu2Hr4cLVGulOuhnkWpNdmdYfij9cgenO5Lr1
G2kVDx8L4JZV/eUGqUhAVz3+1zb9P3b3GIAD/YOi9VpgO6ZjEyYI1khclky0j0Hf
1ElUugjmcy7X9tr+aplQCH0u8Wwiq51y2lekbHmsBQ4rTBPCuN6ilKVMc0WvyIhG
FhyKI6LhNiyOMcL4nZC0uXCjnjOc4BJ0VuVLoNx5p7/TrwoPH6buAWpw5oTlInZI
nwbeAX/QaT8OLgOeja7qwF3LaVlpu3yGeEfmJvLMq3ki3fiPPNsC87nDqAwgO5W5
piwGuZJsJws/s2JSRv2Kpt+f+8DBxIeeUWbT66h5Gn5mlsTtnJQXW02HIZ2S7BwJ
qpSNEkK8RF6BQGkHwBl0ico/o/CV+libMecuFuVBG6g0oj4QOYvnLR86v0PNYGyV
jFk8IvPtZNduYXJqwAjJ/506Yma+788ev51wR+3TxhCLHXDuTgRkAbSLaH2SDUka
JV42oWLprdFP5LgiFVvWEQTVxppd+AC8xoA1Rpkr1UwqeCTUA4BXiksRIQsJ1e/O
C1o3+pB1Bi/LnzPIbBCFvSP9EymP/Z1ztkhcc4yIaEMPPRcKKlzYVX3iHq4cQ7Kf
mLiA2VHMydIaWMQ2mDcQTx8hHcpV4JzPanaa+ohppCntVSQ0c3Eni7sSor6le/yd
vIqknBlV+PHbSsyw4pN+0GvBmvI++p80zvUw21ne1bYPRtxHnoWCR9afID5IQftI
OhZA5vB2c0s8V70+QJd0S/6XYc1/FBiP3isI4BU0gIo+Xt9DaUD3XOnRbIKkZu9O
Nifz/gLw7e/ieyLkAp2jTp0iZ+PwGZ2pp+3FI41ZTmD9FCbubeU2RYcssbakFVuC
zeHV5IDJnH7ha1+dM00DnD0eagP0NLgmidxPhGvEF5SoHN3DIG/we9nC7vIGAd1R
RO0CjqI5xTdO+XjAxbZJps54vjqJ+SOS2MI3ZI6SElt2sbKDnVRXyzLTgi2sfKYD
5HLN5K8BUbgRsGbApOfusHlGo5hiNk9WnHS5bb5quNLCDPBR8PpfroF4XTQ3xN64
CH8Et5jKUpQ/AszxlQxWB2Rg5kMLFXHrK9UeOT3gru618UcAfhgT1DdkiMOzKzyh
/kmhw9hMgmIbG0nngAt5jIH9H/tz18TU+7GlOfTXRXSt9PvfMY89De1uPrQ4QtQb
T/c42tI8PNvsH5vr/vMYXopRraHQcAFYwADnKvPD0cklemN1lv0mgRrjUalbex4l
gtVujyBQK1tImZui660Ski50xi/jJjDIe+qWWVdwAP6gXOa1t/ur+CSlaRVGJECC
rrC6YVKefVEj9m61uQ0RE1mwLqt4s/7TpIVACQ3ljfdkZF5tcjmlRze4+/QoubLU
Xx+LVLpDs+dbaXvSIQ2WYeXj+SY9e5gegseGcCwlF5MG1bLjTTLuavTU9r91tOxB
/cpu9b3l0yvYJLjjOo/MPBfdH9euJS+A1iAjX88AbiquVhuzUKNocEguQPBKwaHH
L3oVLgxsV556nfgoX0SUk41FtiL7WYM8sijpwCLH4EAjefpSNqVApfqVORaX/oeH
i0xkTO5m7fOAgyQGQFYP2qIvuFj6PETm17sFCc7KAR3/fM80EZDic5SAMHATmwou
0cbmyuVTV1WFY6zvNZZ0UbHxMuUmCEHCjKsliHs9gpzdUt0lPX0pKfyOqaDuaedJ
50cHySusyUPIEjAXarl3bqb58HM/hapPSQuTHwvCaJ7EHV574tj2L0YwATskxXxr
OxMjUH6q8Rxt5BBQOTD2XE15j7ZJbkBENv5qlnZ5zHwcSNUE25+4u4NEhp0d+nCC
ItpCnu6tSn6AbcvO21/C3tM1WFrUBYulbkpxjmV4SRCIsxKjQENFVu6pXhJtgulT
tu5125pOlp2YM6Oax5hSbdhgnodt6Z5JJBSDBJfU0Qu+bv78tgCrLAg+GzYpgaSe
3eLDRO9hLdyDxqz2zyF96Gfl3sLf0CRVONoYcJwbQN689cikevaQK23mA8mjEQzu
oA8ZVLGCIOYTz2Uu+EE5ZHAHXLBE9TpYoAm/BhV+n5QE0tRPaySvI29E19H6+sJJ
lpQN2MSmpBHGYQ7ZChy3HfZRoxy39oN/Ki+sQsxb/nxexytHENKGUmAJRa8pkhfp
gNJ9s3zkish4440Z8WQ1g0HVhGFSrSPNemzAqS1LdnnLSWz8s8TiGq9jttuj+i/I
TyPulKARHwMPEn1fBUGce99WN4rGz1FRqEMe2ImeO23ajsJwqV/VOffW3tlWrjbn
L6I9Gf6nPOvA0+SF/MPgVr3Ozo2FO+LAkxoukF6L86C0Ftt/h+vl6vNdlM3evJDW
pISzK8cM4pfptfO0jmL7j68PacZJvyVyJRblohEpxUJpqntCO3wXhoCEiQP9yumQ
BoGC4jipgtJcErBvr9cBPw7pUamoCSg6iIrIbMrW3JxHjgfcNjPWYNjsqDphz4cn
hyXoj3fkc66/3LysdWRPRpkz2buIpS5wib38nNpQIarr1UaB5P9dG2WD3D4gCpnJ
fJb3PhpYYxDjGJJ6orm8/bpT+NRmNrnCvwacfVy8uhhJa4PeNSFagwmHzRNgMRKB
AyFWINKkOh4nM5nP+ihqRbxnHx/64AHtgpqdPakF9kmSJiMjh0CuX++x4OmMD+m6
XJq7FrCxZh8gVho5aZDAfIUNr2+q2haDZ/5ofbuLJac/EI2/uKS0PT8IYXFo2oCY
PWkVBW81g/H0lunDHEzNpjMoKyiSpLp8BXnqz1rPp2N4bAA0Hquw2mLkIiT28knE
4RZgFDhrUn7/jZRg5uoQsILgz+u1u6UoLbAaiPFl41yuqDGljtwkdjB9T88CoCCG
R0acJfqDkypddOM6VP3kLCyO47LT3VrKF32OecudD/fL8loADmvihEtKzG+i/HAO
+XEZ9ijozyzzpl53CNwmkhXX9/1zcu9VEWO2quEqZcy6zlk5weLZiIRNlnr8Y0Cg
0MKBmSiYBWYT5vjwA5pFE6+yh+dj9J9UaCR4MCQ9K6Z5r3fTF8BWEKGvqxSBl17P
6w57+UNtQJ4MiLy/WlbsCoM4u13yo5gamIRi4T/hhd+EaV1/BXz83ET4/4PJkKsw
NdUP1ATi8tGzvqdeIzgujz18GtRBkYOOX44WECJ0y3YcCk8y8DTFxbFVcTtsERHw
nw3+CyPRImqBpM4B9H1ugOz2fB6gBxE9U11mMbXizc3hmWs2l2b13NTIo88vx+5R
RK51kDrFDabM0y+X4Hl+V6kExBWLfqNppJV/hwn8/PnBw4wdIT8sxJSIkvOZJs5t
Z0Z1ff9aE+07U2dAmjgCZfSMxkjWrVaSxIvae3wlsH792HatFhSdoMKPgF6hEd0P
YLrVbRsrP49RpDr860yiGqXT6n54ewx1y8IdQXye+N7WTiP/anK5NmvXrSdt/yRV
7aag+Rkrns21sEsOMzF76KtV8i5lVdxPGnLwaXGoSsVJl6eRIl8l6NSh1YDnI51C
KZvF4cBtAoKqoyTwSP45YoaxazlgnIY0MYfrBWYzEFc6vBO2W2ON3X1CA3i2shqk
eh5vgpPmVYRqFlTCv91GEG8J1tPWpmSqf1r3qgHljpaZn3oCcXzaD9epA8WhWfL/
ASc14rm3UHE/MtTAwi9XNcfJA186UjT2AAb7tfKW8homEKLSXr3qd8otxa7a6OOk
ujt3IxEsoA2AjAWXUxYldhQ8X65QvOdMSelxae0PGB6h0shFWVa0r0YVoYcuikH0
pYEWB8O97i4RacyGoDKsx0VmQtTqzAivl2PkPC3W4zLCZC0mpwfxA2zWyBmOKSTg
T7db3IIxGYXatpA7NkrHnh0fBWvm0REUjksa4xsNyMgSBg98gfZzgS2yPbfW/unP
hROq5n1oKVzQ6PQ7NOsLhRcPE6/+PC+cjVUagP5gZki4XZ2MF8tBFzUtOsrNxidG
+Z62H5e88Xs2ZAouJLFkO3tOWJjaNcmQysAdUGuvlMHezXZKK/L+6moATqUDgJma
KKmRpOcnw4bRTIaxYCAUdUXZWtRJcDUbIBPf+zEBHEDbUdYrqaecgvu/UELOtl9U
ae3RqTketSt08Bd7cpatlDR3tL/oqijO0yA1mrataJya+CKwqyecyEyNKNJuLplJ
QKiJIKICX293SWaJzURQZ5AYvOm5CQ9ub8VFb2FReouqNvuOGI+1pQarx/6IAuYe
5mfT9TFtVnDOc/VwR0TwXXjdOekBnHWknws4I09PwhWCyicCBdM6uFnESFn7cocR
lIkwVp6c+epumikz6moCSOmOU8sYcDN9Qk5HFXREFAy/n7IPFwxdqHUhmTYmvB3z
8SpVYkkZ08agTUmAQb/5kRPaaYYtE2u/kwD1eC8eOKcqWnIQScwk0mQvr7eLy+Ju
H55shvTzx57atPQ3E6LiqoV97p6C8d+luWgrLY9e6xHB9UuQ0R34ZXrly85hbPbJ
QfRedifjw8LWrwg1CwCIYMWJMqlIxZaihBhd2F5XXeLaMZg4aE8UO/ep0uFiaP/z
GPsPR9jUkPA8AB9A2UB8khc5rlv5pAwVXPbHLlQfP4Jpdu9CBOsNFh7XSBOMPhOa
0Yz5oSyeazlZmSAdSa5s2Nd3DPcqOQptF4XH6VGMIiUJrLXer97fXHMF7HGtQzVM
EcrM3x0ZaxR+gU4Rlyiw5TiX1MIeB1ITvK+2czzZ0J5zWX7MV6AEEnwi3YXXytGo
5ssGqMFnhCwBulMydvFVOnzZQOOHjZKAUlILGdQWNcRPbMWXdpZvu/3fDJe3XMFy
DEy2wV+5zG8fyYMD345IVhhTXPn190e/PfPl3lPorp8JI7zCzdCcVfCFzfuQHxUA
vteFzM0JTjSHUYOP9c/ADXawIo+bQOTcGWmXNkiJ2e2V7Cw6Pws1zC7sopTSyQO4
g9wp/75zaRetdTovVf1iXmMetpt/FCq/aE6VrrpPG5PbHI50WL+KKdRR2txh9fiN
fQgzVKoVQ7DoLVQRi3JAeHP+XggMRj5hFFbEoj1+SVkDEmVdeGH4xgpyyUPzqn01
8ph2o7BsN5rsCWGrDhTU8pGk2m2s1VTpaztONPfZjGIGyMvNzkFwZaP8Dtvr04dd
41FzpzhWipvyQVBgivlVQcRuE8bxagGsKMIahL1tUSYKC0hNejJg9KfL28EuALzH
GwHxeatoAGixfM+rq8DG82Pw5O+aJtaR5LbAeup4tRgUp9HIL4AeTcSFPa9ljm6R
SBxuzqVELDgTg8e58t0agmK2O1PJYq1tkqqU3rvGI/vi/SmtVqUORmF+Da2gJk3Z
UozpGUnYMwLqi5R4+bATh4lzKdo+tvBZa+ooUqOyFM8ZB/wiy0W1WBEZakU1OkNX
LQFQPPLGrVUPlACm57ML5gRDJNKkyyztd4Qh1HxKFb5GihzSiWY1m9rt4sLEszUs
9f3Gemz7IdwrX8CpcpfesIKRMjYjF1wfQGuzN9R/HlI9uVShcBVMyVJvQzbxh7bH
7QwJgPof4hcB/dqC5Zllc3AgxQVsGEE7ufOv/xJPNWEuRtOUJFPl6dXakwrwo2O+
+OUWcnIdTBli44VZEQJSjW3rmfdtwwrj4cLJoZt+UYhSviDTBNpV1op/9AHE1SFm
2VIR24boV4hcWEcoqoEG6HkseaJGmHoNz7aZfZj0huGHrDeXhr1mZzfHQ3lxdZuX
mFCdfdFrbjsTyBYCJ8H0sbs9c5PjH8KF6fOHtK3wMcLwllh7CfNrOk53HpfsIVVD
dKt9elfHy47MZaO88bclHipFAS/p5nK3Mp+t/JCMsAOyyR98Vpg6k2ysrPvJHmp4
GFFGUQJiszXjp47VNN1eZ8L7l6Cc7WUmqLBFIdHz/JusCcZ/xOndWoLqB9Eo2hMx
OJoSv1xnOP3N8/0u021qsmq0Z0yX0jmAcJ7GmqzObt0J1arxQsRqdb+hfI6p/idr
AjacbWurm2ZSoYFyulu6/uMs0sCLDgUgbBNmX3GSOMbK3LGOMx2fGb4VBfTEOohG
vL4bhIxSq94gmkvmjwGKuyl3BOGAFLmYK+TFOAkB/9hAbO9EjMNPMy3lbaQtu6Co
oUMPMB8aqrsB37ufk+XByUBVJOpOsNbkXLG/1lTVR7YZyVr+qaLBk5uQvqKc83zB
yZoTAnW4TtZyvWW+wQ5HuVK/4di/Zn0XdhtumNjGeEW1BF12W1FjR2TzE+5rQB9M
tO5kamVS4iWPOnRSxip/UqSER8ZJ/a4SUq5VB705ZIG8VV+gg9iQG2VljZI3ZS83
/Npak0+BQYgIJSKtO14p0tdFpaqY9VDWsdout2Lrag3/pmUhqYc3Y5xcUgxNUrc1
gltIl1flZLKb6y9q41U14nz6mhxnwIw4f/GvwbcTfPwfoSWa3dAQFX0btyCA6+xk
ZC6L1skZgC+esL4et0EIcqGxFCtSID7Zcg7i5bxA/umSBcgSW1r96mX8RTQKwnkK
cuT9wMTqm/sHN9pudX/P4ngD6bZboXM+ER5yD4atQYBguCKjt+5Nf09XgLtH6SZ1
5UwlFwo04YamUsCRYxdZAw/zC5ASEyMRhmREmnOZgQkYebVg4W0touuyM/h/6kXi
YVQRTsz5ggAMzoTUnyFD3Y/UjkZOwqWZkxw5GThdyvR7WNkhPKxnecb5ZtyFfgjM
6no8g1agKjdyFfzJ8tDTJBcA6IJck1chVvnltqOcpqdKhVB/8EDFRE3pxuWUMUoR
uoPVlt/pVEUcGERfeif5TInn6i+O+GPliAz6PqQuAyhzeJdkiuvUDCIYxQ1/Gk4p
9zlAjuBQ0HvKzB0HBT7Z3a1f+2P5NdOeuAueYWadvD6NPXdL5yMex8gJGRerjmOH
MSUr1E7uz9QUf9xr+xqH03gb1mocGLMx60PRzIKIp4PJ0ES9WZVzR4kMmMu049hn
wxOKZ9yqZZn1jJeLsnRN3En+ptWnhyQxS+F5wD7FrQ4B2lW2FoEEsyCHsxPXeuVH
Uzk8Tut3LPhWYJcocaV676IwH45eupaVWDQ5yu1o6ZY2601p00CZ++ewQWMm/x4k
kEVq1jcmV/A497ZtrRx8YFhBS4tLGEn2MwoS098heMxvIy9UZEjL7sV0cDwmS4+9
80l5mYNkYBfZoh2Th0SymhKJCVYLtGYq8AMLI6XKaw34/A9CLycQCgIet4gBc2Tw
aI9Brrdq7+7zweV1UwIY4eRkehymTa+YBU1W0qMGj7hnlO5Pu62V/dyuL50D0kxy
biiQ3FGLh7+YPa+CYI8kKPEfisATuCviE0Adf2M4MzT+RoFBwEL3McY4FDTzZQNB
ZAx1BTo1R6KSYLqT9nIm3hlLO0qZmtnSPuojii1q0UXKqrXVo1wItMyJgorVc100
P2Y9HdaH01774aQ3lEBXr+fWS4pTqofSFJlGH2IvT9/9qe/XmVsUz2xNxCVzl+aZ
zVWWu3qU8amVjldVrZSJBBDpKcff43KnGLkW2coqAVIlFC/urItn9NjQK6pUje5c
qkgQXte+J4tGUGLgbzZC3fmJDlwTeLitZfLC/mO80o5ffxCcNUgzPEr9qVpioK0d
FKmyKbcoxo5dDva+9oX5anQXQtnfdCimPfqx3rjwpQd2oGhfF5pjjjORvRWHbWAv
1ihYipGw11g/iznCYduLgmdD9y1mPHnduKlCkYcOk79l3hNs8n8+/FTEAXxZb2Q9
VT4jX9cePv6FIgPNFIBCRa1873jxhRqNUIXNhsBH+FlGQBFAPir5j+d/PWTrMyKK
X02idUFyPzrGS/zQOjcQmZwgnb7cQRePhUvoNv+A9rPrq2vC3kITC6KmhzJe7XDn
hkRkmgtzefZlML/4sOwBk2eo34PdTzJwSGgMJqUbuOnjpBQ1DM5ipAw0AUE9hUzL
+0JiZs21ZQJ4ChgwT4xJSJWRHDlj1ZNeCkUTUxpcqZr/qpyB5uUeClycWXwBgVxW
BuQd27GREmLizBMoT2Fs2VOXUv3dc+7V6a/Fgrptnu3eP3PFARrsVOSJC97U8wtM
d1OufeSM3PemeJbRX/PQXDZVdmLoJW5KE/Ftn5yjypLIP2ZHRHUKY6n9MHMTTyFV
+9Oyw01dUCOW9kNhQAZk7W5oRaSwJguqh7CTd3YtfpIK9+51LrJb4JBEUkWDjIUt
yP1saWxLsYaRBiMETz6JqfaXAmGxaCaU/IOT1M2QX5VYsBsV/9quDlJv9rnC6ojF
RiGF6EYcQ5X/s3qSZ/HcfYXBt8vl4/4BE15NZvc79OTerGIIwGUr76Avkcj+9Wft
GH6pvoTAOBoQ8YS0r/f34lMCFWyKwfCsx+/gMdSPlwaLv9NEE6+5mE99rlRc1Cl6
DFzbYLmDpaqFZPDz9cFNBTnCdKob5qt3SZ7Wpc9R5Xk10u65uwTC3WSljCS32lO0
wkH/vt9pwH5W1Nj/qb8j9iZBdqYlqiTnattJR8u39xuLy50VV+JwGO3jnh8XSJ3K
RxD0Csd24l1FMdhF4yfYfGUhiABkrfRdrZTNssg0Wkwx+/gK0IVf4amWJqANNFAZ
C6/OW2ksPeHzCaXCc5Pqui6WCd2IbTMN3bPpRt10XUSEIuuDzQcbh7wshwHTICDZ
4thJbLjsCaZ2ZGChU+P5cwZloKKEIoXAQbKkJrKPoGIYup8+EZ8EMNoE3wxRMwFT
q+FRgP4yT8Xtp0BkGS1EArN8/WIkV/bbdjsxpScj/PzOlT39HbnlSuZOkagulJlw
gUWkEBlVVeVY3OGjzIM0y8FX5YY5QwTUDMZRW936FOw6kmAaoWbRU3003fvpzYyN
C3DRujTwDBfevWTTa+tYEpjLz9LIA6RLCc2e1ayqTOO/S1H37TGhV0yJbbDx0yVZ
izQIrGUcr98IYqTqovqJMOQafykqV/3TLmCPuh5jZyj6LkidDd5e6CLqp02szX3d
VYxFARy7jaIN5q4WPFWxyaX+a8SESxVPh+1hnOltAWRrEaXosZV5YK1pDHQPCFIu
ZqJRWTB0QW90Ub4O7BBMXbteaHS1WRzCKEoW4JyZkjSlJghTT1di8tdO4QPIa3PF
aIEsqJNXmf8QR1EpBpNoBMxT7PFaZlEOHhpAbr0wAuhfiz9hVhDc741gxT9Eh+6h
Yjczf8TZnA5zLbUBsGZX/BArQiGKAYu/IL8ZGinss1DYSqAyvt3jkfnUH9HBMej/
yAyiJRgvlVLeOwQAdsc1jLGbJbshml3ovJDg/T77ar34AjZLhD09XsZDQzZ0Chkx
hNZau8ou/Be5XBOhRkAJcbEgulqWKDesZSD0K39wp95x0pZGN1VjMpXMVMZuW5eB
TgPyiOSTE58ZAZdgLfaJWeX1zZpsLO/3zNbR3vAxJCxLd2Le6E70LeI9DLuY6Vc/
+1wnCZYdMsRAG5A4D8uZIPi6FWYwXri5u66dCLnsI9QrpIpZc34WLkpvwfuXaJT3
wRxQEVjZHIfUPIf03+Mowo0svKZ3OilYQ43h+EBDI8VbVQoKjcr58y6vLE7/gECZ
ro+I2bOLnrOyF3LBiHSyGaCc853EVuH0SDrJGeluLgd+9s7IJpQ38b8Da/vqGVHz
UnnX/9pmzSWqPhaoHEanZZkgELMxWi5ND3/ab1WqhEXbXJFD7SRz+czSqXZwM+dQ
xZyCV6mc6yr0taBfFBoNVNhicA7k4IXA3+pQFI64+OwbxozKEmf3XMWfqOWfhY0x
KhmBrFbNodgj1bOse4SOIlub0XCd274GQN8pSRhFQ2nPhYeeHztQFD70RrQqE5fW
oyztxyW9hBIy+bTWeFnvK1MxlsK4UJPZLYUph4C3C/NuisinsNHhbw3qdX2SOUXe
00wu2EDrj+euc/xWmly3KC9HlPh1UKW9+sUuQbGxk7Kon8bIT0Sg86bUWJwkKYCD
zg6VqjzEznS6/JNel6zmwDAA0hOzX0gJDgT7kSZTad93hNxI9m736E7q4DfTveSl
yfq20AOyisJsd8RN43yqCLs8bQhFP1CWJVKiiVKF6FKfgXLxRW9jsVdDxtABgOD9
beujlvhs6N/05N1/xTyFd1wd22Iy/Aj5i8TpPwM5umlhb8v0GHuYrqus7aiiT+9K
QfqlJ40vd/WGY/dqOfIs0np86GZjsjGLgv9i3rrjg53H9C6xRKSvmR6BoSlLXFNG
NYSwqzKeLxyrq57IBenoureJ1OiB+ZiNohu3SI0J3Y3kflCFVAVPUjlZ08qPOFN/
5aXy20y25+/KLKL7U3EtaT0UpCnMgnCS3yEwt2Yqv5DcH0SKPe+om5zHSg2gYuLM
xmIgt0ezlKf0haBJrk6qUnwtVFxDTt8rU0yH/DWOT1Chr6EYoKF2H+zXM00fJdnv
pf5J1zG4Sj6vkdbA09vgH6u9DG4Ml+LmDD533S3DkRqsZuXGEsUq8ClNzRxUZLAE
hvJGKEmGDd8JkVCDGLnZIFGMzDeX1VmggYd96Q0ITJGGA/LuzQqXtOM6mwxvIntb
XjE891zVvr0PmdpJNrrTUFHbVUhZt8gW94aDw8shy4TWQTCzY+50SgazpuJjpap5
+UnSCyu5kiAsyRVDiZPLyLhGnRfoKiTwRPUQZRx4jBOm6xkJegvV3KH6xJ5Me+Jy
jXRHFNw7hSYXvzs2svxh0bzuxET2/WLY7pwGP73MpSwLPrA3erzUkBy6AwKNtQKV
jIDnvxJsL2qcEBKqhtURQq6dGdTZ8nNUa4dlK1EIfftobIyI02YJD7T+6ZlqoPlu
d65m3tAXV4Pp7N7+wV6yZavZo4lM1Zrmq8MJ+okGi3S6dbrQDD0+FukXEMUl4cT2
tQLCBcaHAMHpOsrGXJnr04jV2RDUZvY+8GDCH33cbunf3u94hqjnOQiDXgZ0HzT/
FpyWdJ+aeQpp4/K20H6nkXsDcLErMRm6eKw9s7pFGuhf3rm10LkxSHkzO5olo3Lk
qS5bSmPManZdcdZhuBcj7lXV/T+bN0c80RiUBxvr8gJLZvYneCrOd+J0sJG1RGOq
OBfYMW3ulGp0WFh/12OEfcD9dQS/x7l+5edRJKhrUSaKCdlMf8OfJ5lXFT76Vlor
bFqrgCQHb3S/tSVGFTKCM0hSqXUF/RhOIs1Gu9xwDwqi/DijfkImPXgPWqrXuG24
QDYSvRlqBp44h05AopIEIRxjcqdO89AYS1mv+oX00pYZ5UcJizFlSU6gO6qqyT3t
j2amhTE6iYnEFbFFIvvoxWQyOhDCjRFLpa5iiAwJ9RFRXSUNGe0pMCKbmxNZTP7z
LEegUwHeDOEW0m2VWqI+lsEPNx+veZlLSHYUxoFG9Dk+lWA1wtQj7Ks3Z2EH20OI
l1Q1LFtnwVXsbNKG/6O0CU+Vk1cpt54jbnalb3PkFPtQa5VQj+sMroGt6Ra2oa2m
2WfZgWBVzBeEjfzO2sgigaWAflco9xBj2rgKpHk6aRdVeZMnzUYRDB2QcC/usZhu
Yqy7WdV1OxXyhjhSiMho9GT1RM70Rcv8nEuMN+OtWwz/lAQ0IgVFIQnLv0U3RyBw
4F9fAHMyTr6qkfCz9FRrYXhlhLckhHeNH8Th7eHOpj/o/Tskb+jgHGnvmea1yTLa
HVJsvibTSvxcF7xNZCBSF6UwycvBmCEO+J76TEWKEU4mVTILXux8HhPDmo8YZrVy
bnFlXiKE1zqGXR+13wCfJbkfx24sEPAWsJlcAJu1iaPhigoWDcQDtXWrIu4u0yQA
bCiFcRVHx+xC26Sx7FYfmuiHMuZSaQsq6+hBESO+IysGFlAK+VuqlTBXJwMzZSIg
fMLNYhlX+3HsZP1i31AsgdHfdAY24p068lo9PMJWw8jLPBkEc6B0UWhZVnh67WwQ
QobFKwtjhlSFLNwsJL/e8V+dTwxHFoOim/zXHD3d/4I3OH5orAD/OOlzcaPCMgc0
6bdRwPe7pReVi2NNv7Wh+QuY3gsIFJvcAV70xazWeordPfqzTNu603CxG2jhRTaP
WWKtZRdbblf3zmEpoMpj/wwCAwA9/HTaWkBVkhnaIi0mbF67n35aYiVLaTPu0j6E
jDGTyYE09M8E/n9JHGp1QnO+fuUhVWpApqe77D7g9GquRKwnTmc3C6rWV1ZH1WLO
G7Sx0Jjw2isnfZ1VjdX/z7Sgd5zgFWxSj9DAahAfzcox7RzMgRjIvATrCrwMUbF5
iiISSqcXcb+Oxlvcg3LAQTqxpfEG36z9Q/4tvus0WdisJtv9+7P5Zg7CC3Pus3Sd
4MqMTRLYIwavXzAbGeAuhOoCXpRgBUBOtSDA49GEj4I89IBFypTURhgPg6cffZxv
Ma/miMA2iRpRFZL5ssXPeFZ3sCFqanhaJPO9gbgZ7tY/e9jkIhbqiI1hiYpY0Iqn
I3/UNBlcw6moZTbxhf4vK1EeaPKyXxQFNEf6pf2a/KVMKjCKBeo4r4OOGozHPfKG
Bh1zjZcysvBd2wghFiKcodfmJd5RD6evxTUCOBiPb7gQ0nvV/iBmopjDDiAx1H8J
gvYIQByhCNBxTX7JKEiOO60mv9FYh4KN3WBwD3jIuFVxGKJtHKqBUgk4VyyGgxgf
yDn7kUEasZbTbt3AgDIDlpWkfVMvsvN/0CrW4tgcdvzp6KVx7U3tZ8f/QgKz73YQ
tRKaApV+ZJWA8kW6WEQhqS+AzrS22W+szRBgun0qn2Y8EnDDfy1K9NkI9kA1WYji
qb63RDe25WCUmNsBq027pjpelv5VajKvVkuxI4FWYVgdb7Lf5AC2zBr3a5Rd71a2
ZGE6A3S7wT0liKmexGn1rzzDawKuPbUsWzN8CRyaR+TAOYd53MjLVD0+aE4og0sm
a91zlNRsjPMLttxa1zJ7cIG4YVzia147lRZ5oby5OvpmMZegs9A2N12VJIQNnKvy
4kGCA/bGHa9cs7jab1iiCb6trObJuUUETQ0wgv5OLRX+PfZ3AzkLZHF4rs5oIWe0
BWX39xIf2KlPruNdLDw4vj1WYSltDfpqi1UTFH+GzmeJ/3OyFUmcjB4q+hkt5BYQ
X9aGTZLrNTbhpPXWmW0BW75c7DXqiXsEH+KbL3EQfQ84QfpxACixdcm4RVj1JUBh
7KY323AK6RfG+YefYyPytnbShlYRAkNXmuTpLHt8tstPnj7ctjOm9A2/hbaJx2Yt
/k3rScl2e1H1j0Ng1R1YvyObgsuaaCGooobxhtpII8mN/Aj04Al9GuVv6ZoCVrRE
rBnchAf9sZvl9XKiiMTjVvD4tMR4oPGxx3yTg5LhfC2ERTnqCA/y5pQd2q/ZM0EZ
ZasT1HzGFsw0wsu/oMexc0UzAebgha6zNHTUWJlkuxMVk31eyyyQBIiLci8ydB9k
99l/xWma/2pJrck2O57eGcLFiPvz6Euw8YONaO2KWn+qfLB1IU/0OmAYD6tuMQno
RMUmBP09FwtGP3UMqVttiqH/75j00nbbiDOF7CapG7E8hKa/oHj4gq51u6L9h8fM
dw7+5TpKOkWf4qeLqtHPG9DzOrLTKQM2eXH+6ljmb5AqC3PJu84N4eHIF8YneLMe
dRJjXKSosmthOTbhRMeRLxu4+Cxhf62oO0MhOkscSJyfNkUFsqmjW5pjlDbw0SrF
P60lDq0CClXXCpkp2rgv4Lkr0jTCgXpvFpiNyOI+6XxSRjuzDuibYFsSvnrYyByx
e1BNgOoeEjX9D6660sY6WM1hFMfqgaElwVzKVkn5YcnlTAOFrfuvox/dv84sgllo
0CowOA+PDu1f0W1oexYfAMpPrrWKwLj6ITClgoiKx55WgUfhxWbpeA/wlIt/mSEO
qeORakKkQRST/+HSxJyXwTnASZS9kwZFvUpXFU0PtDkmFz7gKFrSaKRlMPT4y84+
n0anWiaAh6CoA89Wv58pK5g1mqeEQmClc863rEnUzaij6ORONrhG+KH4c8I/crkV
BEyGUx9xnWmndlLwfg2GAn7LZYhd8xh5xT1ycHYo8iGYqLwYjiwGYt+92FCGfvsH
evWD3DF3K/GecJVVRmjIt1TvjMz69mlFRvj/qZmXJ52S3MpxrSkiwP7pRuAzVR6k
vyJJ/0aD9UeRk10JmWVdsTXrcadevxn6mSdTYKwVsm279EnbHzt1bg51zRMDT3vN
zwocLdKKPODdDnwmOgnmk/kRRABVdGlpCkJVztKxVG88Npsb9jPGLKb1SDpRRyje
xksM0QjGa7OxwgrZRuCiEIUu+GB/qSSB0ep3lVxR/G51DB6+sWllhMd6gmGjShGr
/LeOg757khY/SGyxYx7QddFaoT5EPrCFL3+760bGcwSq4c0O3z/qn5GfyF7DCqQB
Ow3knX7KH2zg4bAn3MZ/qqQhWCMJtU1qZ7BTpMt2BicE1MMpSmDR1BcSSeUISXSq
bKwMwpZVYEgbhzl8OqG7gsVmWn74HW3WNQIYPWyWeY8WwtMb2yh/142dRd08FkeY
ucGvKHMi6Xvl9zEXMBPKY2YCHLOM2Qj65vkFJWY9g6KOnWuBRfyJLIUAF+5eLxBH
X7M5cYmVSzI+2lMhshIG96fUypzYOIwXis3gBXn08ltU26kC4X9f+Lz87ZhTKoqK
4LqJq4KeeQFFa+SEGI9n2w153s4pTDM9VVQK/DEoeE2viuO/1/ULV1D58P3V6sBF
MXSbFNFKrEwm1H7CnI6Bb2NJ9NwR6biKZs8R++PaZIUDrlPu4EKZ7VYPEQsb1+KY
GwBrCsnaEG4cpbCDtyH/lI5WeRq1xKfJ4mS7EoVPogK/qdulrBY37LwF4gh34oxf
a6/SsL61GkNUcW2S9akT8NxHA4KmqHEkrL8VFrSFhg0MD0jT6a8uqLWj6SqtR+uA
lnQ/9zsrQfnMt9zyw05OfeS0W0Cto7n8cAXSknumbIF7jZ2LKjmacdgDxidFdFLN
Qq5azYdDYi/JPAGvC2SlRYTwxxk/egSVeXB5nqrMflzfXlyTEN+gNOiICpu35gse
3p5ftmin8Be/rx3oU6rJ/qTb+zJ8+/tr/FdRZL1RuefnPsaYNWeLWmFe2l8DY0+s
h2bOnczsYUY9kol0bS5VqrHWGDmqE08u9nLlUqMILtcRFHpCUrlFK+yK4MrIyO28
Jro0fAe8Yr8jv12/6DKRkdwgb3M0FNIvLCn1tZnVML0DBXeGFp7o8QogMsDJlxYB
WC00eUSpYp54UjycwqXwUMd5pMcLmvKTFzBIihlbKpncBQ8f45wEfsSpUydRolzm
is32qx+72ab4/2DPo89cPDgz5y7XHn+PhPxSe9ltRUP/h7j1ARdGwV4gOU7PIMTs
9pc2yHMQPe5RA4XRIVORhC5FCdb8HRzxZBBHKapEMS4OdDW1dS6wQLm5tbkI+gu7
8AnZWldFQZUBoCdqHIOmlkAib12jLeJn/W3YG1D8HyOp4d8NgPVBkGf5vCUokUu+
mMO2qjeUxX1xTfrkRJKqaeIH4jqkORWVlOq+ag5T3/iEJMFmNhKWknqH0ByAkvB0
HhvPCBX9iNAhihAY4rXa4lyp6yRUtkk7/k0pl+pyy9D38Jd0bnHiuF2NIxoBdl40
bpiQJ+HYj5zsdUTE/n0lXUd1w3dGnWlRGn2DEZgGtk05nnyNr6cOvNZaL2Wg6Y52
FPTF9ob1N9xYFwW8FStwKwR4h69JACNCzVnuqXy+QWJZPikuulZLhMUymZj5UWRA
fDpnQly6fE211x4bZugEA/y2x8nj8xLOsT6V2EMCV5rvNGF2N1oVRvQf8nXaVENg
soy4SglV5qXYmqR2YqBhAagOy6hKITja6KNWAqEZt5xMP+nC/StY9CRPGGrWsFCf
VlhretXsyk0M/3l2gkVHZz6k2sRpiNUnDrJO+SAfcGvlRzoJe8l267g0VYG8UIpp
0CepDCOmaa1f/fcL9B9sRUNWRUBEvGEonqWBcDl8UKkH68ULtiiDN6WffDOT11S9
tk+QRdZe7HTMuEAm9FCe02xgHG5DluCu97ZqRj/URf1N+86dZ3Wp4nRnqVok31Jo
z927wgaDEUD6NAGJTVeI39U72G0uxbalZ28c+UdKukK8Gjdfw+RUCVI8H8ho746a
/EQmHsCeg5mySYTKfu/ER9Kof5z3xNIdqvc4+EGkbhSMV4Pl/jrEBpBU8bi+6Yu1
fDtu2+ai9jJe18EG9jhjMp8IO/y/Z49LOLB6WveUHFJNTtQef7vG4PPBrXVqNQeH
BXCcICa1BYuY7gqmpj0SVC7o+nZz/hRbKkxFbBZmhBOsGqhVKqRvRDH20v5B+Dsp
7Y6NW71LNPXRRXc+vJdWC4IzvF8y2A9ik0IZUUEVRfsqsBaOJAIFCLQsZSvmDlsk
kznUJp+DoIB82UVPx4H2pCBZIbQnM15li1B2lrtopVqUZr7khe1pgzyzOKZwHLen
vXNUNVO3ibgnyuEHOqKwSJ23c4YYsP2qOQQbV/iDytbFMKuugqhsYWMC9CCaW73/
Yos2xGfWZjGjH8VioMKj8ptDTgFQDV/B8KgBcDXoXDewzO5sqZ72Uniot0WvYZx2
xlV60DnhCy8oUIPfAJesB+VRv+iQaWCcKXFmqngxBFOBnwaHhxm7Zqi/Hg+obdqP
tAXm54r0oSciXsdyhcGp1B92B7FykYmHOid5A0qgBbYd46YbSwhzpC0uLVJrbrdQ
T7ouVGO+nC82tMYJ6mFxRhq3wBFrfeste+mh+XScEP44+HqdxfEumYYyo4y2M3KY
YgRcMQtnZQ/XXDL3O2VQ8Ll55Uq2eIL1yNudVTAPI9kMP84IbpSPA+0pXXZvKKY3
6amjHoUGMf2PFapasZpvf47PoU1nqeq0A5viqzHXXeAkHnmRuXs8HvDO640SOkWq
WNOpKO49vAFbuRDY08OlYI9WO0YMCtsn3wCY78UnvyjfVE6qWK0mOUyoZ2oRO9Nz
CUY7cxgqyCTWb/a7QjBGcH9uoW8ytuaTGGyOgUeVl1YcXIe0PAxVYGXF2UhEVbdY
li3Wd7e8jrBwh6XafNlkMt0mk08gkCy2aMaz9m0Mhp7qLxN2Otcv6132oZ/Cxf5G
e/ny1tKMqnH0rjbP7FUMzcEw2VohgOcgO2E2yL/FFanCjk4bbcnN34pok3+odCaX
tQ3LI4SVWFbRm0m6ppHKU18Qy+WofgkIJ24S8wKOI2eKIF42VQp5RM93OqsyH2Hk
LZIMnVexj+t17AZSN4gDIFN2Dx3xRHjo1eWYet1ksQAmIm2FB70foqQHOwZ43FFa
cSmmMgsApfl+oWmjrT98WoYBeLEDNbDbEig7/WAfl3o3Fu6yN9j1hIlvHxPgHLdk
iEuparaUxYUopdocTCNcYf+0xQ398mJwnBs8BaFpAXxtF08frMBbFz9kwM9bvi4l
x+JPj0I+GLAffhrKMlvclX5Q6in0oc2d7cVlh6tbeGEFIdj43HXj9grY9oBQ3KfP
O6BBmBNLjSRajcX7p4XLTEiEfVnS9TtwejOS4CPmyVF/uoJGCxmDawKF5WXHKefL
ak4zur9mfNKBWBJVncm/LDxMyJtZYhGNTdhWJC1wydLRIB4nRt6p67CPm/BZnTMJ
VpkRk9PGJJUFfqfYu663DmwU9W8Xo/7+6vJd5lvIH941pTMw0TGRP1Yp0PnlPoYL
JBv1Ss39/tAFh7LuEwCBWheitEprv07f2pQ283Xa9nveF4lj4TxFl7fmWxZA6BNS
DeRYXJI52uVhwFNhNZwiJlMJPIU/uVH7esefXOBpHFbb+lnLalGSmfUZ/hUji4Ic
FtAckIJSvCzjLQc5r83y1k+JaHAlhS8ocqOGwq0pnhlZDQ2uYi+rTOshoi74bxA/
5cCLktiX/jEj20HRrX3G88iewlXGnUYihLvzDLMAuOhB0IAzQJiOJv1tgagF3gYs
gc2GGDv1WbkLAaf7gaEt0YtXltiXr/auyEiCY6GCM/R2p3AMdDoqn6mvdsusGVN6
NWfgptTULzS8Ddzo5ET3lVxTgOSTrO0UB2atf0NY/lWk3/JvHBlbZ7Ec1qQpI6Bq
0HMFvCG9+JSs8sqdhkwFukSNqspJIwLG9jIt4LcJ2PvJMozg2xgZB7CyEMtPV2af
8PuAGRKqsDoJMVnfec6/X9Vm2afZAxZY14OPtE7VCmlw+jO3y2TRhEb5bkzgl5SJ
0kQ3ks9M5i16054ND59EF1OAOzoHeelad8v5+g5A6ZRlciWljAl7rzSgWnQwLoFR
YKEBAOMLsOEhMq5avb+L16cTiooN7uIu0Dto4fnIO/0WgOfx81CDkpdc9XRp9yxi
vdnEA5dUBdPBdLFpgaaeLUxiMj3e3EzYUGaOdloQtqsY1MsrxXjr+QUSnK41Lg3y
JRmS9N3pz3djqF6cIH3h5qkgbtlXDZNT9S3DtaQRoXYKmKMNahb82LwwMeoRgL9J
ctSB1lk1SXRsGS4tJKl9N6ubUeDVNbj0EwhUQqODkNgxk0UrbYRDK175jTjKCqtY
O9y0jgPf5klPUvfzx6eQyGLhtolUPLRZFs00BmJQHRBg8bkWwnsAvsn+/WeJbzR7
3MkGwvZweKgmx05LmXaoc3/iHRlwSErC84pTUi6yfHtVMX9N2VmJe9nO/go83R/A
8aQQV4mHxgXmIYwfH+HjwCNB0I13VA1pI8PcYo/Qc1KteEPorKe7W23Vi7cbdxRf
rm7KEUEkMOvvBKo2pc5GrT1EbNz39t3C3/TArtp0IsneBtD7uvoDj7178jnjeAJH
0obnImUAxpIZ7pX3rR/qHW2qdluXuIxcmz9+/gkpY5WorNZKS/g6CiMQfHg8mCG9
Hk9g01J2/xjt3oETDQXkYXVhUmxDUs31ZbnglOtSEpM+q652nfw1KB54kadEi8m7
PAsZHzdt0g8F9Mggj72g/arKzirNoL0n7PvLG7KoOncapOpwOb9C9h5cSqVhb6Uf
inMy/r/idFRd+gVFXhA0rsYKk0KNpXhm+fLOZnlluzqKNha/6/Ws/wwcwTICef5N
7u6gxL+71PW9Dj+CXKJt0RR+y4Q6BYxAoptZVMZyWOF2eaXRjRtZ3mqMCMJBeoTG
rkv2/aCt0VBfbMscL9A9JOGspwCwIi0RclgJnk/9nHFyieHw0ZO0zP2dkA/AuftC
nLlVUNozbUPE+1Vc2u+6CIqhWbb0AKwsnpbohBrieD8M/OijXLOWETSAdCCPyMij
qJQ5B2piBg+heO4dO5oQytgjXzjXygWToQMqPGATg0yYPFxuTZPqLWAlE1fijqBm
FZNNkEdaW5Q0EAxsIZE0OGnibfAggHDdBBYFDyi9rb5xDNPD1s4kHvMp3ECvIFlG
iWq4G2wWAuknVwH3RZcndLjmfFlMKneJVh4/BjWEjSNLJLJSrFNdgOXEag/wFrTE
jWWU0Jd3ufyicDUkUoatNRUtdcRfHz3HUiBtEc9DNp4FlPG3sDxhMYPZ051BlotV
kDjae5VOB55nIwitjtse7Ih0taAeqf002sWttFua5rVsr+8Zd772m2iMgQexf12U
lTDByE0J9d66icUqDjtKfbzvJwLtLtaKDDleBR4s/aOAco94SZp6fswMp0Br1qRn
tcs932c5yUXI4DgzqL2JsycGaABl1bZNryiY5I1jPLlDQmHMcjL+ep9NCGzmX2dJ
KLQUXTNUugGkjlA/vNHxqicVC1/0ulAPF8cW6DDaorHUD6dCF1Fyrdh4VAQvBsZ9
1W0PpQINcO3zuqur7x2WNIhJPEQy/s1QfCdYUhoXZwMaP7FkcxHJZVJZJ2DyguUJ
0bnaXir3UmbIWTzCc8SgkSy8MeBwLK4L1wEvN/EsGtnBEcxHFRGFYTA8mBkhrDck
5jwFNGsVTCFGi15FU4AaUtW4IuIJ66KWD0n99OGOqxH85c+a0Qqvd+MJZs7qxAp+
Iq+TSKqkBx8dmwSS4WBFVkMk2zwFfeqGZ1GhoDD4ckiZRxtJiB94GwsHNIBYNnoE
C2HyEINDIJ37CopIwp+1/YdSimBOiaYA9JVjIQdRj0YkNR5zG/5O6Zi8Zayo/NPE
GvQJDc4PDHpOUMfjWYmgEwZC2JAsCr6qtQi+qwpH1pn1RM2MYfQudwu5rqhSyH9F
xJ+FCXFzKNSXaQjkUWyXy7Gz7Q9bd9jc/AanNeMdkcG/tUiGwb4Tthea1DIedoCQ
MbIVx3/7Ql1QDbTzg+h2HLWGH9QUlj2T6o2MPBLlDSraOP/YyGYJD1c+QeN9vLRy
tuNMYNpwQce5jUwszTFDdjVyY8VB1mFmhvlW/u1XL0cNSl2J+b7G3AhvrYE4+VZQ
OzgeVcZ8Z9Cz2vJYUBk7UFhPVaDhixcpYTZ+nbhNMpOYkvwk4KAiqtzTwh9NHJiS
399892azJbWURiLAz6etav8DBRDnPTv8K3QB8/VewIsgNtHnt+930m+lAIlDUTb/
zWofDPxdxo5hCwlhqXmUhpIVyfzTYviw0l0EVKepXn4jzvyJQtF2AKvlO6T0hQmp
ym+lmQy1yUPz+uQl+sP5Q6zAx/FK0CUjlKFQNIvfK8dqbf2tKPkNo0AJZXS7en/E
ZEY3wl0CHAB55+Ze7nMzdksocvbMFbIuoRdLgcdFDG2/3mJuM2H19Yx+8xMRZJ6Q
5/O0UQt0KEepGrODSynJzAdcyWFiQs+36PsHC1OYwTXYWuF8LU/mqHNldSzKDE/e
BggcRepuy5pymmZ5S8sELMCla1YbHDaoWXzmev2SaMGhpLNsE3yMvaHBuJiC9g2N
UpDnx/A5LDd1uWLjjZVD0TV3B7KCGpsKOk15Iq1WBwk63EjLoqY4XtcC8mu49nkA
Sjkx1N27jtoGgtuZqD2EbEEPPCdJ6OtyqzEbYxBEAhCGVVQqrR4MYpFHwYa16SH4
2HmiLnbb/uSo7kWoKNhrTP0DEbOHx1MAJFkpwW0SluM1WQnomEHRtONd3toA2+xC
FkcQ3EtGtij0IwIbE4j7KA1HjXcIo9xWUO/E6PPA/sTQ0L/swQ7RhxV8sJtgVCAu
5WNrYjsdvpTgOgQa3+dey07O1drfxwK9EbOKPahwvFti0QdVGqcXMcnjZHrKbAQY
2jfuPYwjsNiqLxCu94jC0EoleEBaOI/3hK8LyTi66cGDNEz3k09EplovvkzJTixS
KEk306iC7Nxt7HChQrg7Zh2jX5lrIg+5uGszr7RsE6GxJNRu//0VbfG6A8/NbWfM
rMC1lSH9h34nBMRph973i7zMEgK3KZbmr3FEqSxmkGXVkCeWci/XylKV95UQsczA
obbmvtkkbfI6pQnMOL+tX2/9Q49A1WOoZSohArN32H+obLXfOiV21XTQFQzLF9HT
Yazn8iJbROlICc9pUl5dWKMwnsdAlLwZoGDJTb5kGoSCcRgyAfQkL2wkVPCeWI4K
rs+nkYtEti3KiiFxpGPvmlPREQy4UdzA4dwhcVEUOvJ/CYyjyCI7g+CFp9j/pDdk
Dv/6FPJXd8r04wxkghPqHRgpWjdcAk1kr3J+gw5Em01xrtSJbTZSS2bh5U4W6G4D
hSU41NvRLW4yM0A7UoRhVcjisVoGlXL9Pq/ArSU/HMYozHZ12CpNsFuFbPmk1wKv
P/M8NjukLQcohD6gnP1bgAWVQfjIM9ztK6XBYeWzF4Aci72c9cWMcqSAMfCFOrbo
q4YDzkqNBISsNLLrgOGZQA59zM9G+JL3yK15gvdIJbKnHp0NgD1S0aMDAYPkza+Y
zWYAoIDuykj7lhamct44GbzWrntkm8khjIUHUfCop8R49axqVm35IPOSWEXXxB/1
6U9BIJwXSV/lvLwROk3RXEaS23jbJLxYyuHUqD3+9UW5vlHfHcpl1s8gJGb4dy+1
g1R+9bkEf7ldEw/gqPF8jvfXIxcLLOMo2vh8G7zH0mWjIWjdDE/c+HwuN2wF4CLW
yh+lN+QX6RDerX2kI1sh4KoO+ELUpTky9CSJHNHdzcAH2QEhX4YhGFzRchHOz/wX
3e4iYGPcvPAKhlyxX0WXxuC2HFBliONre/75g1KGrp6NXEBQv8qMtN8jxBjiT0ld
Ks2VzDjXh5GxhHGaxSs3iVO6Gsg2TzQgmR1ih6YMDT00m+ZItlOyKTlvgX9pgpot
7BkpMWYs4iVhcX981fXGeVBAdaTRC2CzhMcmO/IOAny3392cYMneuQXTYb/EN5dE
SwA3zLcOYsqlTE0Gb302yOyq5Un8FR2+Fj9ccRLcq2TEFv9TZzcmgi5/GL1xsl7h
y0CxNIDPaoCFWZC/16+pEwWkQ7GdyjPOV8qgyAAXVLbT5OGhGG7TYAqCQ2m/jsZu
CoVhai5HhnGlfRbtBP+TsDtbblCNhKovO6JVvRyiMWMYVCRMnzLB14iJ7/4CVkR2
dVXxIORQ/+FsFE7eWkNZFYcCUX5Yu/+ZFXPC7+S7AOP6AAqhQCuy0Io3MyCIer6h
OBCFFbwz8y0B4dBgT9Sb02D9Tiiq6jAsrO7kbDhl4e96FvbeXmYb8QSgoxLClm5V
hU2woBijjZUCDnFqnywBxyfAPSM5J8GMJVmEJPEwuOe5GZXExMWWnHS4aDkecGfH
E2paD1DHL7kJTFg9Zq0oZFlIIxzMzsVCH3m8sjyW81W2LrXI63If60Ei9abG55bj
g5o2ET9VusqS79ti4+N3i95KbKo+bSZmm0uDHoew29VsmP8PJ+SeZk5jG/tU677Q
P8jhubax2bjtM76C5ZlInYeTEZptvFeWdJN7aTC2qWcWKbmL3m7IhMxYYqq9r8vj
VzP4Cf+FCb/xoPXrSVsmcD1NEFn9g1U48ytB9s/L5GTojV2eaQf4VougAdfyWNM4
kT8Z+1ayjGy0gob4BbSUlZ/VISVbDN7jKLYzchonk0yhLtX3w+uQLy5/QDgGUlQX
HJYrcxFK8yU3i00nQIlICZWSLRR5hNmd4u5Tf980BDlnxOc5SNWf/Or1u12TqTfd
uc4b4Gc5vlI4FdmzqCP8v4bitMHRdaTYh4LSB3vMgW0FIwLGx3Dt5EieZupbsZsY
pKk7CrX3xT4MnBonci+DQk4eKsgy285k3TD4mxhSw/QOnNzynSIpE+BDesu7AjDp
hO9yI7TSHooMU8HEDKCjuJElioeSB1qdv7BWUA/x7qIhstOwa3MPYAcUNgvLuDZK
gxc7CBMRW5BQyIAeirS/PN/pZPfaWsvxnL2DmNXPFlUelXIy3dSCoQG8/7in6ACk
s1KPHwNNEJ/2Imv5NJwqBeWvjmbFLlQN7o3kHPnXjcLI2YaOT3FL+RwUNtCZPFyf
NgxDZPYZ/nEbrbaqAEBAUFmFcOeXu4QGFt5ATDuUbaJwirSQOLDHvitchUrJ51qX
w74fggMfd/es7DDll1CtVUGDTwJ1GrwIOgEI3JtN3sQVQS8/LB2CX6/mXBt6x37g
MW7fwzoZ7VNSXdbU3YV+39CYX2Iz2PQ7solOK3/doVNzXwm2FpUyueTJ9ZGt0iVl
aHZk0idPHPBLuda9zNrIyqjZiynsV79s5FIoQFg6m7MSta20O4KfO63Sb6q0IBL2
Sp91O+RcVMJTv0IKE6DVszUKaCNa1jNTkoCYodo6f5DR5p68D7XWXd1QmUVpOEhg
z7R0bTYqjkFBQOfoyBZS9sB5/GHOOeAFq5B9F4ScIHReyYGWWZ5Mmrt9NiYbAE6T
nx1dvkSEUflNE/HCkAdpQxzilTXkFPQ7PJHojzyCGy0sFmteaiOy8TlScijvKgOJ
EXvLZqIA38t3gsKja4uS5xPM8vpMc8xPKtqRRx5bzqr3aVZynhup2UbxHsffmces
+vKou8Ct/Zg6XK56THM3hkVVXGXr9Hp1Lgwd9X5ex1y8BGJmhV/XXcpxXqlUi2+t
tyOyVJpGf87dxul/pZ/LxkbhAYZbTcmJG37pFK9e3YTPxSlUL5R4krP62IW1nNc3
oqs28rzH3mlJrA+WRIOyd1ky5Bb8oB2ImGKkuS0UxCF+cNQPAvGMcsAA4gfhpQTj
DrrPAL8mzBE4AOH1Um1/zmTFybD2I1Qj5yJbinMIL+m9Qc9ivtvrgFV2JyoTTwhh
JUXk/G36Cy5ykrYdTu+NBqqL+uvFPKaP52oi4syriz1qelvGfVZdtJeJ402HJflV
4Q6eSW4F/WlFAtQRJLAiINdY4uIGFLzRsqTlJgoS2CxHjdlrz9xNrQleRP//aO+i
5bn7NaV8qrM2V6sPz9OfnPrbKRHNEO/pzSvjf5W2gvA5DpSvT2itTI7D+6N5TPpC
/SOi6dQLbHphlAWcfKZ7d+qJJUgps6chafVccL3BFmsXv158Tmw8DFFWCG1moBdF
u5CbqY82LbcktSUBLqos6NsFw3czdLDyH2TxNeArhXOz4FM86eZnasEL6/167X0O
KjYC0T8RG1DPqvbnfg68Hb4+/5UmDhDWdNwCwLaj+yGms4d66pyT5HaGvQlvH8LA
uO2Y3DCowQiABrwmtknH/ASBP5762xms3v2zhBsroT53d4ugLuHDJsJQxrKm/xjS
feND/oLOfPI/qNLBmh0Jx13aY6gIJbN9RVJDNTlfKvD9lALZ76yOFknxbLqha/pw
le780JxZTk4i1r/wa7+VUkB+B6BOYOBNDOE3bZzuPKaGlluDdwak+mr4yjK7SwGz
KH4X0c7owMZ2uQ4o64AEF8LNHtG473JaVwWFnoJSddXJYRr9JcuFSe8LEvDWdh2m
pPQ3nlNZ7Rj+CEGU7JZ9PDNGGVi9HMxy3F3ELgjpkqJ2R6Rcza+NHeyh3PSTZB/J
DZTf9O0N+8yut0u04St+78ledecAK9cJrwVlwVEwNZIF6rh4bWaY1Gd2M2uX5788
7jBh/k54wWeE0IGnBLjGAWwWne5UrBYrFkOLvvng/GICaKYgG4Zu+lGRTJRzy9O6
y1Q9kD/Jf5iPWcQxRQ+yEqf92PByFcVmrEyiCXIzqzWhVMJU/Htm4l9Vsy0wqOb1
KgO2tkGo2U3ucwdNW+RvBlVbjfwXkOESxpQRHOnn36RbCv6o02PsFtnETQ2bf8Uh
Kx5N7kLMS8JuTbdB40rF47dU84lmEz5mBQcWrI7p3jNpUxSQwp2aPDwKG7hGYO7D
oZH2ihNUNKj1gP/LzNBbjbiWirHrtZZB8qA99HqRmuAlL6W2//43mXR+STaRB7aa
9lcw7e3qJaU5ZiNlWWgOtV8nwPUZUS8a8T7qBl8XnywXKs6TYuPDuibi2yF9/Axn
fMBPNH1nGsay+VW0D4gYDOJKOdelJi+nS1int7+lj93BODVJyLGu5qYvYomdzHpJ
jN5Fk9FJOZCjlDPddi/d/pL3gTTdv/P0BTnp1oSxyrVh5Hticco6lCZxX7Yl34Z2
sURRqsAAoAloAs/3+ilmF/10vxxLQq7hvDjXH7yvZrj4L85b35hHfAadFrhiXGnR
PCiAePJmKxWNfJmnY93iwTDGRNijXTjtrYT08MC8toYKPkSWmnjT0+bdsDjIvZn7
pyxhbmrlQ1HdbK5ktsZMxGLQFCBi0wf5bwHpEYGWuxs1QhzuU8PIO3Z9a2jl909k
BczlrFTrUqVNK7i+oFM+/mjnwYLCnredhI07ph9Ej2yDBAnkJX5UdLouPCNHOryN
4UdPtrxeLLzZXLWpMZ5+JPlhHyHJebL8nRQ9IdJhrrV0O+xIbqNcU7tvNF7X+tj9
C86gsmJ/eC87VxLJpS+MkmaOJTdRYdSEOoK0axnmvw8Lp1X2164AQuxuZuNvUlfP
cqrxRY/W8mCd/DSCskaePzuJE9kQp8n5A6tiUmvKkVbqaqoy9PhXC3+ODgAu/xc/
pcM6mn+N1LgDq/LwmMnMDZtVo8a5TSxVuV7Zd9ES66eq9dKBSxAUFuh+bDCi522h
0Vu6JysuUm5nA7ZzVtqCjXTzGZLa2AsNMlMxPtjEqrTKReB83GuKGB+AHfveJfKn
gtKy6JMeOT2e/hz+xOWhL3Af/PDkbM+8TJDrO29erX6fCDpgQZpgSJSma7WkYc6Z
+U/xdPJ4Qp8MW/dXW5V06JzpFRdeyPsF+UqGs4SrwE2miulYvXHVWVKSj8Y2ikkr
BzzjG+dALZDYU9pzEFmWc5p4Fm3CLDqxvv2WDZrcGROUoeGU+pjEt50GxfMQB+aI
FEnYM7YAyV64iDjWNmIqtj+ePjbGAE0K0JI8s6t9h6AjRpja2LSq0lgrHA0mcjZC
X4rwQ4EYbHwpTiNh5IJNlXdPlTjJqchC8SNKwg+JxfAq5v3Sx25fcEuxk5rMLogL
w1anSOMa9EbBkiX6Ow9vO/RA2UKJkw9FIakjCePre8uPD+8OkvlST3r9GSIi02ro
HVXmkbgixBtQv4Ey3u5S9WA5gk/PYCYPe4vU4VcEeJ6JJd8QiHI8s6iNfJtCv8FH
ZbzQuvpJyhDVywJahyi8TUAKmfZ+kVBkCyE9casHFhKMr56eNzJ9r2xDXkSiSu6g
I+vsEC3+71inwCmaVDElYvxaPYzbVC06zzx9sFc8kMG1vOjozW2Dhyh9LxEvKY8t
6Pcf/cG0ZJksq0G/eSMgmsUjEMQSHd61gJ664eWl3fZl5PZJn7egk6D6AaEfAkCG
UFsuuEdY9dybj6dbPZwQJ/SumHwiYZAwcVpZLMHSQmWDNIVcebgkJ62w+7h9UvDu
9Mfnq6Zhbo2ZMRuhTNjOOQaWiuI+62poUjLGfpWPqQztMhmuWCeFOHRa6vgc1dlR
ZXQboUcbYBuBaw0+AsJ4DjoZZAnwFsPJmqop2nlujwanjOx3NIsQUsXeBtBet6yc
u0H0bYDC/hqHu6EUstk/6epyB9Yj3087IX74TfEEdPv7REqiejbghDOKi538ct86
sLVDDq2aqX/0kgi+cZOQOGwsJy09Ua0xzeyH09ndHVd4jP0liWN9zy2DJSvflor1
i6iMtD+PYIBS8+3/YJNlibLKdT+F5ru+YgO2QaNLg/+3YKWnmpxq7IqWRkDPdtwp
MKFIv/snNjVcxeI8IbiSWAfqLmQv4iziovO34UhFErk1pxypUiBA1wyVBdW8+3S8
PD3+nj+FWSMzn7UIFgOtPFEoFq0iiM1PmGsM/SE/jM+9zyks74GO8+GHdUbb33sk
Q3KBozHzmzcTqAjggphizYfsspc6UhPovUA8ygQGdKy5mOfj8gBNY+0HV6hujQ90
DftBIRYlMwUbB4ySjRQfHH9r25hC0L6rwOGrv3jB9jjqJutYGzEmfW6RQOHHjRpW
hGUQiYN1YMalwKbqs6IKEBqkTdTPgWz2Tc3uO1ZdwZflv5rnny2cQ+dXRKXGKmCo
rLuIkai1N3iVEmj5gozb5HhFUf7PLcB61PfzTQ0Dy7TocwCv6MzSMgiBBeipU59z
gPE4O51zmii09Ag7UbdNKnormrVshpwVElrIyJtIuJsePHGVcNh0nYfAU5fut1gG
yB7/h3HuxoYGWcDI/Z1JmqQx7CLqfgpOsA5Oz7qNe1D4GMWF/YMrfthqtfjisrd6
3qeOeNcck5egapPJvaDaMcFLh8fq89pWQm6YizcT3NB+CUqNJkYK3YgZ0Ozs4pCl
QjyR3DZ72A9i6J5wCwgUsw3cFJMzI8GZTpJrh2WE0bHJEZvZZd0o5NK0hYyENboi
PBb3ePc3qeoKpAie5YJju4wdmYzpqoq64znh+FHQomkj4Y9YW//WYR3TFY4HSWix
zif4dmVcvDvrU9QAmt5dJGCg1bOh2S5//qGgxvIP9u5aamvY9z1eSovEn091BFLZ
MFmlHbHQnKQHnCEaCWe0PdOvl6pB4e48nF7XquWtPB0PuSA7K4nQBIkr3nyfLuli
09FI1J3AOF7HCx5Rxa1RnzGDSB30wNzt164jPt9w/3HxDa2zL5nUxh5zcWdNb5sR
kesdmy80G/Q2bMO5jSLJzIvZXqiGpoT42pU3Xiw/GIjMmQeat3ImVLmIYxd0Sliq
0LNng6wt7Hk6BMmbOiRz9JN9/UXfPiUto+2fKqeWQk4KaY6ouj0xSxyJTQh7CXa3
3HDYVFSbdpfZbd2uMHekYuvFoRz7K9CGVRkhZztBGEBvXftwqPcOfop9yrWs4j5a
FlHA9k4T+4E6pK/SNbobO9tb1YM1sKXm6OxhakgvZH+bFS83qcJRwW376KJQvl0k
WrzXunWKfCn4Bbh/SELTzeBbn7zef+oReUPef6W2OdOQlvvXu7Co8XfbyONTLljR
IWsLFey74JbAZlJgrPGv63PjOE39PJiFbLr6fMz4E1lnQPw00clwGGI/NdKNtnLC
H5ofweNfdf8OfxMifjLlBRBHgPD6h8DLbsRD+gq3UhYGaXge79R2sr4z9idZmzR4
24idC0F3nR1DFE1Rib0udk19MumSEB8tok4s1qH1ymuDaLP+fnhbyqSJP1QAOtwK
+1Qn9vrkWhXRrBjp8d65g9M7jByMx+YlnAimD04zQPTubMKbx3vIxJOR0uAefkiT
sD8F6rDAQbvdFVYvYORlFmpYpa4hc7aLm/M+QV3cEtd+fvCFadIT4N2+SX1PhWnv
jLLbVpn8KNDKnrhmRQi2qKoizmMHZr3RXVG0uLDRnO812kQm7PK3uvwmM4Nx0YMx
vjyxRaMef4PEH0sSIKqZ349jNp1P+fg/9UXTHholVAGIGB2pTSr9ZDJQuUIQxGTn
UnzyK8nBo5akytJDeD2/lKeo66NsQsXaJealMkM6Rg4fa1zEukD0j4PmSAcaCuW2
M9zqZJtXofk3+0+lurjhy6b0kjSw1tzYc5FyGNMbrW5JPq1HK0ceiv0RjjOuMaYy
lkYsyo1NfG8IBPUO7pbP/ZE0lbj+PHvCuXyjotJ8A8vmcOHVaYwGpv13va3PJ+kT
uCXUwyJYQ5g2Bl46Wo5Pj0/FSuQhFw/60EjqMMV/twgh+qe2w956RGpOMbAsV2Fh
ee91JdJUqtqJ1g0e/QBnPX00afzvib0IAHhWG9vfbLWgjntyVqO5Ixla36TTkLey
O51m0HOjaLsos9fOypafrxOaT/mp40HMZXVJFxGOLCvH8ngB910P4mCLaqwfp/eI
nVKo6Kq9xDUs9p1bImCLBltVYVNh17CMuCDmwEWsV+iiksj7X47p6FuHYpDzeCKs
wEwP1CGx6Tb+lDD/kP2GoWmyxtNrBl/EQeB91fZU8EXtUN+5EK5ryrxWjOdGuA+/
F0TJK4OFcC1OKZwlGopOEh9tpFu94X0pDsPlJwfyF3DyzY7EQrVWgI29WW/020QM
qoRNsv2B6Vimmo24dk29eP5UsyXoUMisYPgduTdRLE7fz9CK3andBGb3NJetgxpM
ob5QAteq1GwJ67ZACvfBLGfxg8UA1bCPY9SJZZVyDIBNTq7I+GdcNdeyp582Da+y
aFQfae7f8S1l8FbNtnNG9bX75OYft3F1bkubFJV2c6l5ztrPTOEa4m9xXV6AL3pm
wwDIDftaukX1YdT5uPqmSvE1HiZfT7H2puYV9Ho0cLVT9vtVczJtZq0rdcNWsxBq
IkP5WG3i7CMaq1nQq0z7gsZTXcRdXjjQsaeEsSPCjsx6Y5ogSMeayYDJpi5mUnD5
JxXINTuKXdIBgKXt9QLPBe3xR/XrHW5FGdThKKAR0Es8zaeNeoJpE/6g4zxu5s3S
VK9IGZbD7e8QUw1MpvP+Qh6aLtVwwjGS+RMkbEF4S8bZJLq0Ez0j2qVfGxg6QLBy
dhqEwzgXOoAyRvopZBSEu0zHqcL6+uXOFkbqtJpja1gBEaxMVmrMDZmC+9+9Q71c
IvBL1imSc5UrDMs9SYAFpWbamWa6686lxoYlmooMb960mpWm4mU8k7Jfjv4OKQB3
I2CcHiVoETVFkJgfHgyU7lczl6/se+QS1tUuzto4ShflcyCbSQbrlBOMCFRuKRO/
QCRCgacFsBQAts6if426cQapBva/SqusFG6CQ3Y0nhPLGZw2OeApkum9ZT4wZa0H
Cl8qrpf+kpipJUuZsEQ9dh+EqNT0vrFvEWV2NVYugMQWleElLq2c5CdH46FDdo38
KBZ4EEvK23d12gAMPhZcrYyeZ1oGPG398rFsYlJuodSpVYIhMOasnxY2Dk5p8oAS
EnjAQgK35OEU4452/WytD1QB2t/xQQMSDYcb4bIbzJV+9lEQxl5TRwF6A668Maty
hLWioITMNnBJDlNwqib4dPMLV/82tG1Fh0kDDHD3Kh3yueO9n+ya54+0XTPYkCwd
i72m7tB5n3W3d806X6HW/bXpYLTSK/mcKF6F18VTGocDtIDA2VFp8G7K4rPjYQU0
/ZISEddPupKUT72IKqQiInJNUXFTCwXH9GrsMqFm/yR1WqhV2IoV+Mnr7wmsgCXZ
wHOr/NDB1UTb+WPvl+gyC+P/Oia8PDIY92VP5FNojNzALvgOItdu8bBUqwxOilBz
OgGJdKVqLXCLvgpVeYUTVM2hkLjm7PImIDj9CRVQyPYThpgDf32x6XXTt/sbprZ6
TnJwqswXERJg8mae0e/WOktMXlw+3Pf8dWcKbejxvpyZXL8JNeyura68SjaLnSjx
N/73er0UNx/+hfYO4wesG9VkgPZCA2MY9tiju+eqDSM+TtFodSUqMRyDX4Z1nNJw
pRa3baC9N0VP/pXX/Q/eYUxCyarH1iRSXB0SiqUPPA3s89Ipp1ggbF6daHXiaMKe
r6e2ysUhLbgX7382Ou6HYxl+5e2I0XQFborvCoIU5f0PwIbBtVpA72zE1l/c//OH
pogJvc1F+TVh2eL8nLyvPausU11jIAntgV2blLrTAEvm9lTFia8BHQkPUAQULjRO
6tO0Ez7Vktyx+/bmil59owhQa/Mnh+oMyz1Bj6x0590PZH5jxjh5EHeHmk+AsO/k
zWehS//1ob59hx3+2lYsdrMmUEws+PKYLWoP8Rn0ZkQciJuXICR0z7hRyoFxFGC7
fACOhsmg8yJm/aHEOcJOZSCh7aw2bIHhodN07oKbQ0+TTAFt9fLe3tHCsl5ptQT+
4Hj8sYYXXzil6y6Fod8/kMcKhlXeGpMwGOOw+nohFuX6UUzZRXPVcuvvZry/H5TH
x7sQmO7lqGWTkiSIMmfbbDD7KUyPr06oZh9RzYqgOPtoUaSYAuqZ3BfmSYIrv163
W1yQvjdHKcyUD9/k4b9R7EsI0R2XdvrAZxMJodW+piJXU8vtvF1879hHwZ1UuZE2
E91fd2bXdNcHBdIzdDrOX0506oSb16Yq+iJQBmxFUVpDbpXXHYmcImiyWjNLE8eP
KrW2DoU+/O46pt/rV50zQW76I3Axl8ezTZ6URggJEJW6srvIBp0wW2UWq7sIKjVC
8ERWS6cUDyr9G26dIafR1bJ3X/HvimWJ5g+RSK2N0WHnPaaFVl5hxnKrNqb+HAGT
WMo4l5K/j2rg0BZ+EBHRLLL5bRo1vGnBjVMHZMt1JD8BH6/Uh5fxaBSPiuHR4jOQ
7bVYYJzJFgMmaM4IQit+SeoD6cTAppg1t90+0Hvzs89krQZArB4qyE+tmvxHVXY0
Eav77LrrzRh4JJmzKvWimVyaymfFkrSNHPpdPQrhhV9Z+69Gur/RJ+bWrMajrcr/
/21G7EM374uCRBKzd0IjEU2azZf2s/CKTact3RKYx7CFO3aqG5ss/Iyjv4gamAF1
vWPR3WfKgcToDkN8jZ3gAXxe9KKi3bPs+IqjdQqPST1W9rZA3HQA06MfTdgA9uZC
qNfDwUmshIXyVXxmrsi7W8IN0lw1P3cLkgf3VSapFWL5/2pJZJIDfGI3tThystGJ
SJ1vC397ktaSHOGBdziOE8rQIEwHVolN9NOxNCbeXLk2Ky6H9c95k47reS3jWSgR
2qW/KJ9nPOK1N820B4tp/QJZ/R6/L9kVtevE+DpL6TE6th8DaKSTybqGheHyfvap
mJw7fVNHCJLdQPc0G1LC7njmfL3bvx5KFCxKRbPgbIrY+FkFsTY6KFR200TVbuP9
tlIAybo1gqbfaxrsDddFvFHRLOA6RyeDAs82TEOzzUupv9E+pFnu+TdJQ+hcdHAE
OjGMPKEg77O87ErzrJ5MkreAsQRsmQKBwExg953yCu/spYrL7o/5U0pKQL5X/0SA
ur079OuhF6wwpd6Stn1rtUP+z8N8uKJAL52nREETyOD4p9NsQiQAE6XWybsLXIqv
A6qQ3phpBR6DuwwhAaKW023qhOKNmzFtTFreh1pT24UkmEkMYUWM3n3t6SSCjAIx
F9bxcPLoqkkWsVHd6PgmEHumzreAu9OBcJohoOePKIdGRurli8Eh36KaY9tsUtw6
eies/aoRbn9qvXsEDfrzDDDtnef/FFeJ7dtKa7snX4wY7CwYZ428I/evZgjlr/Cr
fMzMj/XDlKWGsN1soJMD8Mxoqz/xmhXU7ZBazT7u8w0lhYJBheGm7eZrP+8OTahk
cN8OVPD4mr8X3vt6w5P8AkBv23j2BVF6XtogbuHkKevLWZtlj1+LO25KytOno2DL
iQSQgOT6MPskzu7GggZRhssHnGru/oDw9RFM2qNS9vfD4Ne2i6QmuUU6S3Yu35lH
yJU8BQJ0GejS9xXuyr7eoyCSoXwS65ubYBYuJbf7XKN55lNQ3Vsj5PX8NZ5h5t+c
783RDm+ag9h0Pd44ijAqrP3PtGijmuUeTpNYGg7W5LnL+ZxyYthGAAc7fQfjYIrS
cJF+LQ9of6vIH5jEdBFWLdxT5fxYm7ieO3wQ9oAEyVXPtRc/Nu52wiVsc12EuNrS
e77ls1ngZcTFxm0cV3JB9jqgn5S7wv+xEjfYVPoMUt+mvXZecBcUSImT3LZrS/64
VcVsEF5ZEoXBnUyCOFI6lzYy2UOvBpwB8qBE0ElsPDT6QbQF9sM56bfglGelzYY4
GdtNgUDdk0Q44uoaN0TW1YZ+mpEO0uP4Dk7EUv2ZO16TnSWb91GY6H2QWB4YzFX5
kPUtRtZ5K2URu5owDPTnsYoGZKecAueo6CmYjNRyUM5WSkObOMU7M50Vr0baml1W
h0tjZcDnstqBFc6+ozj7tRtyhJPykuckQFmmTMhPIF+UtygMoTlBhVnPYGxw612Q
JHj7ylR2e5lVQWTGNwFnCQB/V0Cndh3bhxuQoZBGLuKNw15vN9MTlpgronLuMx+7
wIA7Fwxozh9NqQ+HYYESgUZAoGvwUtPwO8aOLCt2zxMuhMGKZQBrdAMAZn2NyOAL
GqIdAXoXEnVYsyf8TubC3azRR7qoh8geuIAlNFnmMFpaLNj+gAwGxmIe3y8gRldi
TwkxF1r6NsxcR6rwoP7FCx4MWh98JySRBDYrldlYUwuohSbhydWHiyIt6DE/htt9
jLNn22XzGxsJ/fAAZL6GuaE23k0QrOVdibEQW+R8vOP9z5S8Nmy6z9NRo8BOYYF+
8Uvcffa8u+Lcd6uZDNEpI0E1z6CEPdAF7tb+nr2x8CEkw3dUE/FgFabGbfaJ1zVs
LIDPAk6MxtBdlCviYoassEAm780OWEpamAd2iXJX2AFIKDD4mGMsYELzjZqns2jO
+mOElvPj8gN8vDz4pCNvn1I69XYN1/ZnZNIcfmp7WqfY/ybg1RoqyviG8oTnZztf
Kz5DQ95G9kTGvU2iKlgKR+yYAOsyIrsmIU87gpXYsrNX6eawxDhwhg/PPeP495ZH
AdefxqyOuBuq7mZPMfYl9GYc36mfWz+oYbFMutfj2vSCcG9R9oGVZQgc8IFshKc8
QEai+e/DzXRMbKXLy0CIte2MazKxTHTsSkftWkSYEOz6Res8SzK8gwR4UVWjv/eu
6e2WzSB/v5BMHKWZbzVGyzlfCeOGgv3wwgJ3rdpKOuFxLN3dzyQRvQh39ZRf3TL3
ejRWFJsXUXzNa68vZcyx7PvGGJ+MH+GgH5dralx2vyTEHaE09Vg2NPZsQR+Xl4E+
iHkMAuQ2+0nlUCzdBC7kCFReJEGBm8uDd9eP+coshM2SUooqe0WcqdjlEmFXCqo4
XUAvxAlHIEfuO9RpM1tjd5lJcV8ba6TOslQOIF+dIS1B/3KJ16jqUOL4LSBRzHcx
uz9RaW26pm4M4cBydBDBjoN8oJZKC/ZbriPVzmzoNc9QUjrxs2Gzbj2ZIe1q5TVA
V35cqItAP58sFdbgSI/HBr52wbKgWG4/DDXEZA/rdOaXvCbJj+o91G8tztwEa3DU
cwTV/1xsqRGcYuqnwfezNDk7Ater+xf/+ItYrazcIexpL4FvyfzuMd2FxifucBHv
bdFa2bks4e/NLrLfWgNJ7z3eVWQrtSvzBOAM8KtoBygISHTt/slP6gBoSl/EGRSl
wFvxOK+xvZ9R2WnOZNnLQkkO4JHfB/cBBCCjz5yi508yyIfEM0j1wctNrRBSz52B
EPeMqyIl/5A2YM5IWvWq14rrIZD57fAtsECbPPYs9tQHnn0t1oVz8uPskAzCf30+
v5MeMSxnUVt3B1TZVc8rZt7FqgukkwH5VtYCb8421ATrXuyScdA+afl5toU7WeHf
2haUq9G1iYhuzILC+kmvt7JEtKwAY4dpRisl3F6loq1CxA44Y3AIRu7xF39NsDtS
mKgIFxFQ9kCQUamgdVNlpiWtG+1fYjleHplWRe56yOiiLnchEUcF1Km7P2CR5/Dg
jW2qSP1wGlgKNhe/4L7CccdjWXHJbX/KHDFY+iMJyODwDrKyrNO5j79JW0RCdl5t
Jgu2YVk075sxrYMax9Chu5mdL6yIY5L7HRg0SH7220wgo9Z6OSLSV2EoLtOg0KZC
RKIGuQRROB1nUTeFRBb4MwEme1dim4ReehDw/lp2mLrqJuNki/xeZ/DZ0W94sJsG
suuVx4vn1Mdqk5GTPULYleF5vuUYIHBEy7zBJ+QPwpH6KK208InaCVXK38bIbWYI
LJRCDlkpeUbL3lqRTUIirqcC/5wE//FOsGufYvygRltxQBBJbfaa1vfWLm/r4Dtt
d6dXgxcuwiGBeEOnxiHfGmoylxPzRAXPme0S0vc6wTIe82hr2hJC21bUGfHlO5ZA
s7rKjLkvHLv4fi0vidOAixTYd7GucF/l+2Dc4aEKfupU+b3eIHCfn1tUJP2xS9Ca
5i0nTr6Qy126bsoIUqhtPPRmvShGcLOOAnU2ebP4B0ra6zvqxg14lj58nI94j5Di
09CEx5ElleIm9zhwcpHiO02So6QYMMudUKrcUbcvBTo7jl7nuSwo4YZKwlQhfExA
GkD3WIUl433zmcU31HShTDDtchvA/FC2BglUoRuqlfEswJ5DxaatUHhlJovlu9r7
mD9+WXkQfsOb9OTBDLRqhMEx7ZLfHbS2/XN+xu2p2tu2gYPukYhaz6qsLsO3Vy3K
taSAme+YWDZ2IwmQdPT97+R9VtVFywIOCexa+Gwd9IyH42W+CToC2FWkcpG/E2/H
6b61r3W/aOCrKtrPlqUpIlzEGT5qRB6PkkjJJYi9B3/meDkkthx1TUxIVuoNJzLt
Oh3vUzWQ4EPmjnDY2W9t9XN7SSku9V9Ijbv5RDblXUVo5uaQyDMsJt/R4WJbvYp+
MW5ElUyKrQnAn3p3xrpgFMPIecwbgUYRi04PJ8ceaaS+ic+5Bufdo+W9ohw/OePx
5+JyzEvc1PhL8W6qJ5gVMjZh7cTKKDIV/7C+PCiy6YUoCtdN3GS/jld5A8ATxQrI
qiHiTJxMMm9T46MZY3oqQs6cWYWDeskc2NQjkSyRVm5c3XZ2DR6NxAeR9jGhQ/lc
to/y4oVFoOe+dk1Sl7le8AF3WN3pLv+3yp/1hmTfXCL2rH7zvQLiE8iqGqbm7A7T
XPDjku/n7L9Ks2YnnG4kKvKmGyvOpzI4Fz3rkNRJYcBfk1mYwgirAbCmJm1YkR7m
5c2/ma52m0AFVH/zu+BDvr7Pixm+QcIF2aNGEbSk4hlaFa/HzpfK4IJ7SAFqvqI7
Rx3WQumxx1Be+LKy0klhLL/W5zYxO+nBeqRuV4m879rQFug9GjnQ4qE8mQTmoAJz
+ZVuoFO9xXM/Kt9VwUefVLptrL07ohPZMtm9osenp9KpQorMokU6w8v3s+NbaQVA
/96zyFLfXxD7VsaZZ22rT+Uub80aVVm8lMASsM2OqbFURkkI7u5JV44GJDA2N8a0
Fi07EakzfknDiq2BabUtELmpuhDRhSc9MYnqMlyXx10pUWcGI+fu4nO+QEIWgWs3
D74uXBuvU2sB6aU0rc8hTQQ21Qczky3ccSaBSOaswLbOJD2RaaTyVxsf3Zd9vEiS
FRPhHg4i0+4WyuMIcgF5zmPtEUSjCV5VWxLVGwIs08uVaWUy8VZaZm0fPiiml3xn
1JKr+Dj3/YdmIGXuSPfR75AK0CwNu+7llgPRI86GSn06uD5Jw+Ykgam2zdd6TXNr
VR7QkRR2b/1ME/Ye6rQK5F1ENqhHULdTjvHGwXxxquJEF5Fjv8q+UNUyeWD+GiDP
ZIXtHpBc/79P3rM+audztMBc6PaCYAPexEW47/7ZUmzZQF6vzZKOqcFx12eWhnI8
7NRzp2duvF4E+HNBoffi4gwmDDnRGEHVxzb02Dzgdj5cyNB6N+v2WPCvuNa0nzUV
p5RsAcJ8YqoqM0XrYwcHNlRdf7gtQ5pRFlBRfHSv0eN/KntBV4aWnQjk50I4kwWY
gZmrHbBwwocIEdtgsipll7LpPF/a14wFtZfJVTEC/JBln0fzhWauNNF9vV2NhWqZ
H01yduzrgnRAGfa//AnKkKbBMCfwTDGcMDjjxRdYl9rC1Ug1YgFXndGrshHuQQc4
bxU5pTNjAxqLFZjlWA1KWL3iJcBVRS4uQjaow0BUNkdkoCGPyiXCZR/wHYVeLReB
zRiaPnX9xdff65TMzWPui2B1tZh5UWzaz1EE51RGEqZmBzVSSYg+tWab1heqhdp2
gInYEUQWO1L95bLIn92d6C+t/LzXnHy+49p2XMSSyPGyoRfk9n6EZyyyY+XNFrYG
AfIMPRlcLZR3M8OxBejYMwTuxj0o0qFKo0vba7BWv5xDJaYNDU8nIfpxRMeEUlf8
pHkt06LIwyUdfBj+wIyYR07m+g1AMW9WCy7hkBAyl2ODS3BIZPxT5/SGfKgsYxca
cQEmcbbsJXe9yB0jGetZTuyC5WsWXCEGa1QVhJ4cNuh2fInGyT4FkUwF7khY+zym
HP2DG1/Sq5DWFFHYKB53pQFwYuhF286GsWmQ01b5Jgd0ZL8memc7Rpx1CwFq0uRT
pM9MdysQ/u3HAbjWbAJNlOqrvTfvJJ/HIFcJoSM567NdLLuWGrhW8KnH0wCB5CoF
KMYyPZaixUPem5An93eQ8/L1CexDIv4jUtXCLbmNXy1JjyiYAnMMP39DwaEwEfS0
UZIRwrVt5LTl1NGHjDpOyFwLNyxjO98D5TfzCZi/pK3gynUq+vYBTC8szAYXpqGH
enBr8a7SF6/8n1keJ3+IBiCm7/VpSVlQ209Q1UoCgoCQJFbM5kTcoyXHSIldWubO
AJkauZtT6+T2lziLnbqpiUV2u9ZZUv3JKapHhUGPrngwMh7G4ca+LgYyAPHVV0F/
XPPz9sRcHr81A+/06EVHxsiQ+PPNdsFufXhSvjCVaVKPyr5ZNpvLTXhBKp3L+K6E
+CmsgYAxwx0KOQhkGz8bAdK1sT4UlLqqMjGx/C8080P1AC9FEw4qMpDkaxffvCQQ
44p3eCN2pAHAW9k47qEvBAA0iV4btcqSheBPlY1IHF3TVi5Qzey9eYr1YIXpnvkc
1HF9LWpPxx5GsRP3u8xx7x2OnqJcirCx9iqvc5jjeuXGvvcpjlNojgSvqyOZMU0a
p0hk/O7ILlyVlaSKXCWPvcUUyBXeYI+trDhMrc5vgKWXUZGi0NBat/KQqNdSEDBg
j7Nvxg5tpUBSH+WopCoz3okUiyRUYlqtkBmqbU42hPC+0wvRSWLK8J2fqpJUU0JF
JXowVBIUVFA/h+sepi8FB51mkMjZE0LFuJzJxhFq75xtrwupZStr54bLPb5UBp1l
aTsvMWCZ/McGABuvYW2D5A2VCPEAtGQhQ8Vwp3385vt2Xli6wIoloj7sdHpyLlyY
kkoqBPPAuTYDoL3EdiSs87Jdx47UPmPfzqcHGPDxF7FL9GqvVTZPAERj8l2w+QQF
Eke0j+kN0uzitPztQKsHa0h5LVDekdSeJGdocsO1tQkCo3beAII3ZlvAv36sG4Xz
z8QhFOnWotd+vkbY0WiyYCczMEgdP4RT/uyzDYuUAEFcTugv7/He20fRW7ijTAwz
j1gx9GqiR2yWzcUM6FWKZO3MiMDNzcaQ9e3Z0dpjCn1OkCIbehYLLf8eO2iM9w7j
lbgCNSYI6XgHHn5WyXGcffbgnxoQ608hT5f+7zDG+Gk2anL+DbCSMdFmxnZXdEdq
tJeU0X0+33UCVk5WaFh3VuEVPy/aDj5sCb72f/yR09LgMY4jP9WVS5Hqkxj3hNM8
1KAiX/3AKrwhkodCgFpiRxFtICXEo9r4Qpv8gaGhS/jJASTxYQ0zkmq8wGZlXuoq
Cfim555DdoTQ5gSzkvtaWE34rWoIzaoOAq5Lc598w4fXLIggVxPokyBhvFC2wtqC
OpzX44QU4dGGlP8AGRs557sXyNzkrC5kjiJRwuXWFykqOpu7QvdS8bu5PD1T4QTa
NAAzHrXko0b3IpdQ3QhrnWalMIbwCe7B6Tft0MKyKOxIipCtvBzgUaBOBQNxj4Xk
HZq1YRz59kXpnm9K4dkR3+PLXz+bkMNl34zP/3nXwFK0OwVo6n+BxVapZPxBVB1X
hrTx1w578vlOxGDqsJGxc2SoFZYYXjCxtCj8/RvTWaDds06o7B59sA7+SBKyZ9P6
4P0d6bpwbjcg1h/L7a/7NHI84+/DYC0xBfDLPrHd9P+BE1FFmztH0hS8CRIuXNGw
TinI5S2YD8sl8LqYN48YiF86RuKThzQm8vilX2jYDST42hD50O364Z8AOstfl4OD
AWBl5L8M0UXipdOY4c8X6Zn62gRCwSPGypABGBTeTr3kCqoqaC69gpxZxvLymP6G
YIZNf1f0phDQQPXR8ZXJ1PC3K9/fthSIckvHrYyw6pC+DHxooVxxXiA1+e6VdG3L
xbrjJz0fVo6gWiKuEAQc+kNG7PScTrQHDCFanf7qf1RuA/+kPxGAl5cv4MMn8XER
jZmqwZ3eT++YhG/PJ86b7UVj4pLexvymzmZNraDUPg6CoS4RTioWsNPOsZ++Rf2I
ZjtkceyvHIXyxGByuSy7uYiSknYCkOhItQNT2XNgVn9bjOT6q4NGxFZWRvR+jUQ1
e1CZhVK5iffU7jzG3HlwrFhHGQ9ywICen6e2HlWG4jSGEsSRbVMVAN7tcF8eGegi
3LknRvp9/b+wTWyVcyrHultfMN/eTQynQwz0rMITR/s3O2PZxN54c97xenSwelMn
Xi/k62rHL9Q56fzubxL+XXRPajZzODNDHmbhMTlWQGWZ43lBm/qKVShd8gg/J3Fb
rWMKDMtSI2oz58ZRE38C7vve3kTbAude/befNcacjeghaFUdXjNWwlrEO8QWfuYu
BkemXGqG/YYSJ6a72kUcNM1BWXrncLM6Pr774ciZIviz4WWmy942aIcsgTKt6Si1
IICvUlNMZEfFqZkxp+C0tt7nzsmKr2JN2ReGkKPUH6Bc83dyvaGITgUOX3RbNxAT
aD7Z+nTnECv5MBbxeH+JjZTnahkwzKLjsi3TN5kcDUVubutX1jpbbv/EaECsKCz3
2RIQIvO1rCa8/wKa4rBLnyCQO2MxZEK7yg+Ug+moUk/nQAn/xJ0NuzZ+2kVMXeHd
Pwfxq9kbgpne6+M/i5H5oQ0LVqeLeARkQ5laaZBGB+8+4q33cInRnylHluw/IVsV
ajqdXI/GKriMMr4dBK/q95jtoO3JJbioEp8uIQLBN58YsN/3iagw3N2okeuInVMv
ZkcWYeDi2pfaR8AjqRKiLHkEplpSey42vptpGCe+PnyOmqKCQNYOcGw5t0hWEMsA
Ctx3IfWUknQxk7S44gnSxWZfBD11JUgrJEkLBiDs69/W6HQCfLR3sAj1Ve2sNbvB
J+j7EposNTjKBPBxuCmfdu9fBUKAnZrr2ktmDpgVuvIAciikiSg7MdlwfsqWxdGC
Yq7ZYI2MU1dL1UZE7IW4AFaWUoDEsPFQL+rdwVKljYmkZ01SuEOwhpooqao4ZFhd
l7eUAZc2mJF+bosWsMxnLVbRvN2+e+5qenk5PFt5tScKb6dVqvYvfWlAS7AATdul
cAaRX3dAzsV8J11kzyB9rGoTA5QPYtsqJu53HPFCuqxFgtm/ECR1tWjeub07b6bQ
nVy47VJi2zMyfUnFFvyuCN8ZsO6itpePzguy43v7ckxsJCiw6P8NM3A5vK86Fn8y
te5VxaBMnI/y/qvQV5g1Na7EipfzZ25gVZzNAV/p3r/7TdM6ZQI7uy7ExscKTlqQ
Ls3NMylt4EyZ0jTWzQpGJ+FymVQBJL850007U1GLaqzmZyfw+TT8VOY2LvMzKnxs
9oyB9W5jkYeCW1xyxvMdrrlIDg5CfUBChFCZcuauRYXqzGK0BtVQezLZ+w8c5O2b
577iI1e6n6W0gADskpCMoHpMCg9tsR30nKzF7BCSIczMIrjRoI1IeUBJ1xv4GKuE
kZhU4ZF2Wk/5nvj78LmTKbeUgmlZO3/lvp0lzGGuY7ndQ5BNjF99GTYLX3sjqFBX
F1OJJtLaGOCEMn5Eha+A1vi6ZZotlGznoQlVJl6DxfEy/kh7GfSonzHpoCKF6m2y
PfCwj/a/iQWaJlBPzTz+rEkicQks3INKOiwAmhnxb3zatsTI0f4PA3B2FINihKx9
D/nvA8BafSl8N7isrmNWkynA7uAbLkZRIDk3uJWe7jw/neFCcHsV62ieN+ywtaj5
1yubC4muXDXCYztxrbM9xp+AcyzTRtZz1PMx2g1/Md7s8cxitEhhmYI7heBZHYaf
rGU28VR3ij4PmRXR7oezn3EVjhZB5tHhDGDU+391r6W3Ewzncsrfr9+Z+LUH+2Ow
5cQUaGof4yKQ8aZDJhbcG5l3g27HuOzME80yaNIhHPD7AJu1o2S5XDOQbGnARJfE
XN1dSLgw6zlawq5ZbpWR8rS3nQGK4Sw66w3Djr+iZkqJ9SUvsCZykTeWCiJ+Fi3j
TESWJ0rFplb4D/K0tSs6IRt0D/AL2exSZA2p6Q6yqEyQH2NF41fK/hIRUIDCM9vM
QxGdAu4VAbkBAtXQudetKhyl609gTI7iWrAVCAtpiXE+phZjbC0hS/37RHTl3CCg
TUsftS0r41K/qlpNju3mvMKbLUPc3fou+JgB0m6P7PXccD2rcGc/MBgIg+yAVI8b
mrS5Um2UngGRlzfe6dKccwPlpzSAqsgxewZJBs8O4KunP5vQwWsPz5+bePcfvhtg
DFP5tigAUlWj3Ntk9I0RhAiHQI1aOLbAm2MmxTSPHrxYaEC4apd31/wZkP0sd79H
RB0wU0ciC5qfHUaH5dt4B3E+rjSAvupYu176VgMbApn2ywP8oj2m5k+qEZ8ekVS9
ptuRLorzx0QjxocTkbOQoF24INUHtNIQeKqgoL9oLXBlCpo6NrrH33O880wcDN8t
zu+/F1Fn217xKxHALkOlH+5C9gaB2YTsfFxUCBddesdDgufLoDOfh5TGh4MIJRr/
VHHkl7SnNIyTnGj6Lp84H7ZZcgfU9jcYQXOF9J8EDj9vvUed+SlQ4EdOZf8skkV+
J5JMMMMw9PO/l69ezYXYkUeFuWyiyeubyIsaJkqV4Iflnbnfkz7U4FIN/BpUBsVn
6+3v7y4Qbcmke6tVRg1KyfjcYfaXekN3vm9y94pEvVLZ3aNN4t9yMCmsOVzvLPLw
9bf2cDnqVCEhtxqWDF514hDFRGby6Kbt0wnjn6nJvh+Dng5fONrzcRoM41vod5nQ
Ya0G/166fnC+vGssPHxQuwa5Xk6Am69bzxuRl9oimZtOYr5BwOnbwVFz1AgY7POG
kGKffAEvdkzQxOV73x2n8Jv3DImDu+M56jLZkBCcKPvENsSV+hRAke4gf8nSLqIn
VPL7+gH27VuKwQlPhlxN1ggM+8xejljJFvHdl0s9oYTBikvGq75LPLJsPpJDxQiC
6ay4IhpgdDv2YpOXZPMnALkRurHRJtBmoSZ4Ky11Yga8DHgtt6zLNhyjgRfaIweK
+qwb26bez+MIiqWPk+qGnrJqhOZ3zqlF4EuZDV9AJC2viUT+SmO5P4liI1Xn9mnl
OO8u77xkvZpPhauM1OHZki2zNaDv5ieybLuM2Q7cW+ugqafBpPuvbWCZtVfFfXvU
NGX9S0wnZtFyvH/OizjkN9Jzl5LfNqxOroHt26zLfQyXUrDjdcid3jwDzu9sRRO5
0u49Yrfxz+IsGxmtkJuH7UO7jvbvHjlfTEEW1qA/F60aR7XbCWk22qUcvWDagUxB
aFAWCJvLabFkZQWa2Ky12JsK8PKKADsrJOItHVCQzyXNO5ZeJcDRGsxbVhNTQVA4
b1BEdjeDVZv4pBrZrko8U0zKv0k7xUTBN30AgJA8PfCmFOADSeMklvrmYgQ0njwI
1bjaT+KJLY8jZHw3TpQJiEPgLD098uJFW/n9I+nhr6ZSzr02jjkdSy5Pf1eQOVS+
G920A2ruG0acCP7TQ3CfHCryi6t3DLevSA8DSiMciXtDMx1Jis+q86gVWhbLmwr7
t7xznygCXKTQ58qo57+FzERWqgYpj+KS/CDP0oADcUUoZHPtgbX2HbWtUBUyyH1q
+yqs1hOdgu5C0ejUUL8ukRrSIvRBkwR3eAO2QVbtZkcJNwNMb91Mi3R/aDwanL4K
VhwGVGaNK7sCF7zXKJyevmfpIuLog4k0EkKraJMjAiuaDEFF/I5ElYxXsJ+ktyuj
1hyNRHR9x603USQK8UrXDE0lAsfU2rGS/NwG9D4oB71iF/GKlmQ7EJws7WZ7ksEv
6dpTJaCtTgqNqRtR3heEbZHc50Iy2Mr7RageBgYR0Xddmadpr0Wwzns44aRV7LkA
n1/b+oW944bdCxeSlz7c6rVTWhcKM0sxJO85MYYKo95xkXk6xaWGd3u5ATEiHq58
TlXNkyKzqnMEU5K3DGiljRk9O4lSce/KQY8eFTmgaDFT6x1j0ZFFjWtNmTdEX2QO
tkuto4gphYIh3z39O5KyMASUYGwFX4KBvtbpkpAAffytEqPeb/K6qSI+cuBbueSu
LuHMJ7FTS3xggPX6TPtLm0LB//2mMPilGQIvK63GNWrmkT7Gb3URHPuoxGX8ACaJ
SA4UG6xUliY+lz09fQn+ad9q3tOT9SbpL4PH5KKjSNKU60A/4su6eL9l8C1YLY1i
S+JxBhCnk2hnYmlwQjFWyUuPpRdsszZPaSvkZU9t4jTMb5eQ5IzffnG0Qxv12DLn
rd89u9yQg1XRhNGuQpVarQUED9SjVvA/fCh6VEvIHzeH40worXIExDlN0ueCCOJJ
zhBTyxtw6Mvd0QeibY4Uaw9wz/FmBJvMfrGhoRGMmPjfvRuxUdUsRTlNPnTQdqzT
O0mRQp+Cvnvxbv0FUx75VSXkZTcs19bZ829RCykHg78946ixwCRWVTuezDdMU0gp
JT6Y/RsdnUv4M1E8vFV9TfEMySLRla6ZAlrDp5e1cuC7g7JFnIE3jeAnFqP2ubgC
c+7K0lXSpEC0md67z4C5GjO0maHuBRTgLRLomzH51upvLJklcaR77LN85DKb6ntI
oNUoAZ0hHT6u70jfQnZilTB9QDEROpeIIvfa6257WG/RzCT5MVKuZkoG/JG3wvTO
p+LGxoVxWjhlZdbwiN+ct/aQ2+uiKEa+Fs/yrhsPlCR4Se5R8VoP0dI/QyM4AVDb
C7v/+fvaZ+2YSprP2152TpdKuFHzNnldFoQ4my3XrD9QfYPJ/a3TtkNor6tmOmCa
XgTVwhcCr1/duISA/bu4aMAGM/a0LPE3L8i4+mIW8j9rqAvyhbTNYKMyijCUMssm
XpbKm572+y6ldpjQRk/h7JU30ZgNCpe1GS6xGEb/ZOm5CCWNDywnZLOQ8JBAXgrN
S89Y76x2Rwn6608LfpVUPWRi4Nd2xzVcQWBB53GOQeuXSDe8qURU6dKXGLhuv19j
1qEfJkzTpqahS4QnPKNoK23SZOTylpcl2WqQ0R2tyvYscPIvE+1Elx+cFfLpck2d
v8OwpoZqm3NWjzqWbiOA1DwkxDaGjeyEihwSDVUqJ/UVG9YICt/bp5KXozr4WY/P
vSxVFEUqvwArBvmLNVOzgGymEwLaDgdysSzLymfkT+XwNCQfIB8lRE2l18kfv7py
QiDP4sAES0Z+2MJ5Czqt8s2EPQrdZikCrF+5wYdr1IRWRJh3D8Lg6jMkY9rzQ0t6
m5f5Qwv3qZLqTOijfcxGqufiQI3+gikLnOhUXz0x9xxAJiEtrgYEvyf8u9gg0D6F
RMuDN1GVN6bFcPYavQHGbFCcqZAcv+Zgy24PS9bZkiyvofSTx43Vtp7WCEKgaGSj
8LXl53Ud2rDsJHVD0bAzHrCzLIqmdaMKQN5TGXarwsTRhT/j5OHVrFzeE8c9+dmn
jFOZCbCAhyOaQ40Fd5KyOfBqCj/EmLwYVTEFWn9XQ4Pb3oRVUK3wWoLO4BrrZ4DA
1yu+ikue3AEGu4clf9UIi78Vae40/IvDhVEhHv9K13wzvzqBqwIQuk6bJRcskpQC
++Rw74bN3W1avpFtZQA3xEAmAS3BEmA6i2Cy8RZz4ubNoJWOt02kvWyYNrQOd1D6
PyS7DDythu6ve1gqqbga8VyYz9juehxsTlo4dNKnk/axM0wgd2ST+6wPREm63BBI
jWpNmSmX2OGwPvRBm1+BPhsIWimoJ3ghvlGSjc8485M3rP2fz63JJol30T0bG2O7
TZ8i2SavNVG9BsRHMI9Eiow65CXZpsdsLDjBEQCgp8kQdsJfEI/KK98OPz/1eGZ0
n+8ITqe4PhabkDKrm5D/cAboWF+rUV9z1nQwh78WC6ZKAqDKOMjhWAnf3/Odnd4g
9RChVPAqQYgnAiWzOfXqWnF+eA56yPL12d737MEwCx9I/xufGdv+O8w9UZc/yk/9
P6nbxJH5vW74Zdgeho0D+dy573wSF3RGGwwN4ITQESEQVnuKd42LX9HMZ4qPd9jz
OIBtJCJWAhpmUGZ7ykP1oMolHpd7DwVxnwyAdKJ5/Yjp6sYTm+JGhCTLW+XAwyv2
WVVb61SqeDLtE6QYr/sFVJ0DdluU+NuLSIXDpAzpK6VxoArSSMQ+PKoaCL96+sXK
Cd3qW9Jb5j+NhD3R8inIr2Z46YaDpBddnTrElq6r6XKX2pqPLia6bObPeCCPONdG
2ujNtgH13Bp26dpfqAZ99Tm5EKGBMzD/70e9fRbzSf4uR97eF5E2fB4Oo/EQP4zk
2czsfvQTqfh/UmY33sqMWUB7gHpL3VBavrRRtERXPCjIq4jzl/c3UqkgwwG/xQ7z
SE5k0D1DmGKJ55RwQqcU3dD6e9fewtf53BHUu4kIshjBEI/VXDw8dV8TrW4mWkz0
DpCxC9XTULcQWXJXGaIVZLN69idA9VBuaTKvYiOCps+L/B1Rz34zVYpyVEsgbrL2
BCMl/kDt8B7y3COlo45ibLqvZw0wrAxjXKJS3hQi+IyCFPfWktt49LX1595u1EDC
BuyRq+LT/2r1Z8WCSGwV3gon2ssQ/i36OzjlifBtV3t7g6cblYvoXoaL3HLf+JW7
G1ihm9PGIDJ8YC5VxmLZ4b7+vwSyipo2xuMHgVpHijD02aBMBHbSEz/ZUDHOCYK/
crj2T1VSjs4ro5p7Oq+yB9crPTHA4Ka6mR1tdigREl382OqOhAWjTmS1sl7l9rt8
/JDR4kVGWUwRjwOc64E4c9sAMM4Z/RQR6di7PKKpaM3oNzimCXfgHGZBjzdgd+Lf
0VUNp/DUkKyi+IRQTg61t2xfxnn7B6UZmyD2pHF3UuMd4bGGLs6sUwk9Rnt5zbnH
nyan1XDMTkFHkveJr7Psl9mgk3u/8lHWHwhOmEqL2f5lY+hU1ewGchwY65ACbLL4
BuhBayDdBdOcozarCPEghtx7gNheje1hOazM7K+fcZ2VTRflxsyxNNcdZEQ/yApB
mEfFIS49g2Q/xzdVgfxfovoaZjUAKi1wHu5ygloWDBZ83xdtAi15oOH8bUFl7Hsk
AgE+TDLri3noYEtQUsdOd1SO1KWdu9UIM1YqzZPcyWMtouVojuxzvtATAt1yMb37
XUFpB9QA4PIpe8ZbPwjEH0txnZkoOtVZuyXPnDtPSTM5xUIPJpqbj0RK9kWMK1Vg
frkn7qqCVYHk/SArksUFpioVr3qmuRpSPiQERsg9s487mHLqXSYhpeRb+lxvapcm
doHUC8TlImhNDc9yyW63u6Vd4BNgrZHu6/mz2KB5pYOMYm8p/Apfr8ors/10GEy1
zfXQ9jjd2gWDpRAZP7wfMPG66YdyJc57znyny+oDgDNPUyQPFs6QpGPZ+BERIYpH
C1qp3GybcmxOd9z6KutRarSa7qtLq1mciJKPoh18GpRAj2rH9bUreKLY7TjmCL7c
DQ8RNatrSAaKGKT6SR2XWs3A1TOFlfvwaKfVETJAQf2CBOOUD8KzQepqWx1cp0m/
kPX8SLvVhyPeH0Ps2/07oMbu5fRksIyfDB9VhfdeeBzNARCthBO9+0ZZ4UpJP+hv
8qD2mjFSkBGo4IOWE9JMsvw4k/UGU9TD9DWQEAdxBGTNNB4nYhtr1pttwyPAOoCB
D35tUVja34V+qC3yRU+kpqD0Xv0fdEbPFK1AuG9u06wL8+h6MzX5AGfmp6d32a4l
UIlD2WL/ZfLTTKmdKuSUKCvfN1/y+LtbfmFJALmfxkqA8FX+fxSqE/YvrtJqeVi1
I16tj8AcTMQmXpFTzFRu1ZPwNmqkpQ83BR3JfziZ8XDiLbPERnQvtoDxBUPaZ00a
amoCwebUHuSxhoNWJNVI9kyhtym2LM0pg+qL1Jm2iOK4SMNYCFca8RiKx5UTzUFm
koL8SGlbNIfctqm58HfQrtO6un61en31wDrDYNwwfl0L4mjUyE/amBRgjCXuCeih
k1DtHv4Q5d2t4jaGbmYrDDo+c6J7i/Mqn4Ws4610Y6DQ2q5/5Gr4T9aYQSQh+Ugu
3fqHVkjsS/oSc8bZz+gKbK8fCCre/qNyDkObAuOZu0ipVX76KSPgk6L8J385D7zV
8qvZRaPvPKwHcYp3OKmwB0KQ1IbwmscYMaogi1TuJ9e8T4nyTFqgdZjQ9iNyUi1c
CAtT36/dSh0zAebI+nczWpd1ircfKENx6FeyGaA8SuuzWyRuRkDlm7az4xoIG3o/
UmYI1Lwp2rRsYsWm9u+A2615c5pFL806y1JYX3BA67O7raO/JW7PM5NPqCG77XIK
IwFFwLqHvRPh5lgjXtDmQsCRgv+fJMHlGt864bNo1wolu7fCfXW+zrIGptJqL0Om
eq9GLc+BR/lL4Ada80PWk4hWX4q6MTZ41UPnMzq2gVT1qjxkkUlV9lFiveNYTZXX
XypTeJYC8d6u2Ntgju2QLiGfH1x3CE/1XOxuN2nLhZriA9it8q7aHaPBic+tiDPW
0iodY0BokvTmSYyLWslEyuEH2gc7qgnaVMz4/bGcd5+FmvPu7J3Pt0mJHw7SgdDW
ZHVM4QeKD++OZqhqtVi1VY3RdYDsg8JlWEMz/fMX3iuB5z4cTBD4XXB1HAJ2gb7A
5ddMrQeKnYuxIVDCXJy3ogvwQWaYaysngOF04UFz4SVB4GunEcEc28gQHyKCvFKe
L9PjlaCW1DnfqNglt8ZiMu+kL4xJ11joSlq2YRJRVVLQrzQqTkLv1FOd57IA/1lV
jQYigta3zpoQ30loWMcS/Pjc7utjbwVgSt16JWQvdqg4vFFCeTZXYrwpmHsxtIq9
NswcY95XptQRg1vaiD0DUu6jHQLiojTbwI43uyIS2fxw2yHbcVpWErLhu95SUxrj
ARo8CtI9hq9JuMLSvb3qyuDbSMEa/IrcaZMQaEazjeYHMUlBihrwyBUK0Gj+OA0m
8SQL5l+nSrZn3vmOExZD7UptTdAgV3miIrGYyLt214KolaQ7Z/sjzyp4J/H13Ncz
CoUK3i8qMfzlz6T9yBUuIwQMnjbIHOWOrp4EE64u1jtvuteJSO0DEszUe6uPhP2N
Cc2jxUiap5tN5VqGHX+W5uHLgn//ldlrjGcjyp7i1XstelUihlgo0L+raTHkZt8H
kprtnuC5+jRS5gMInZF/T2E4HcefL8ZGvlS6E1f7p8To1HMZzXxjDls3uxt8NUYB
7JHZdaiEYS1MSXYAxJ75P0IzFeJe2aqzI6hyc+7Xx/t1tKPEWEjQ4Amvz8mNWmA4
yARR9u3EB3LWuDc6ChSopVtV65viBObv71HYrUb2FQSIvHHkZKQ4FgqsKUwDJxKC
CqHUAasRfYpTlbuM14jzV0eLr3fPdJFt2ZejiF7xzN7qvKlFS1a41nN4xkit0Nz2
NPaJO7PT5RJqNswxh9XBLOSLT1Ntvp8GmDvZPEH19Wm9HVloBGmISvgnfV1HMLnZ
9ZwpNZ1qJJ+U3o6hgobUp6EhyHxx8n0vfgKhjw4YvSluprhjjwpWn4s1Oxlezw46
ET918N9G8q3cV+yXQrpEAKXhv9shAWHljsPZQOAf/dxZ3uHk2PbgCecyrUepTfwW
dqY9GRbDUYlFioaWmwEjt37X73RA83Z1JdeyYYVdXHzzIS0OFqSo/Tl/FNW4m8Ue
b/DyhNrhJlCUdZt/a8yTT4rEBTHWvNhwSkFSwar9H1H/doS4NdLinWkJHfkolFyZ
9SYyrmBjz63406ppFTb436/f28Jw8vssyiHthNYf+nnVYKqeVTOLarFqquhurD5P
NVGAKxJF+AXrBqmo2N35DVQas3bdDp3deX0+hbygcmRu6A6SACijKrAp0twvKt7x
K5on2JyJWVDixgKuIap91J5qL/2FoMEuTJ9gG6I6wj5yFpbNHWss+YYl4uf2ujs3
rS08kgC65hWbZC2MgNO4LaLwRBdYfNNOL0DLRZnFznCwRcwr0NoGDgvYqkAub7qO
VWJuzvwDzXZ4cBycHTCtJOK+S/jcYq8fSVpq3XjnPbIh0OuOjvvvq/indnhhm1Sl
+pCKlfQRjKADqbqw/goAgRH1D+ye7hlE4istELIDf9EICWXv5Ep0gNeUxg8Flcrh
orgWJgNwQqglYk8zDRszaDhy7NxDJwqc+I/SnNlOR/1G0co/bmbdQt1NGzHvQXAm
bRQ2l0m7Gsm8O/QSBXOjgTpvGqgP2Uvgius3WlUJrdRnJwso0KDj+zwIexFgnXGp
XhC1kGH4C7IlfT3oI64QW1HavilUU2I0Eaf1wCffnJllMSevTrfvyZwG6N+LF32j
+GkzqLzQwEZ2/iQt2njXF50oR0Y5zOn8s1gwlDwkMA7nT/DFkoWrmqbKRvEhVgdP
UqiWmgAk52pLZswQg6TFpiSGHV64rhItNkxld1ztefzLA/ag6vvIiAdXfwyUotQc
JdMgrZV/LxF/xzgtTqN/AjrWtfoIHp1tjRiZJlGavYr63hoQq1uI24GuywkflS/Q
D7p2rQEJbxZNWhUe2gN+1XR9eq7yeqeVomvcZHLIzknmDS6vvDVgrBZ/5hbc74O5
FwsaQReXHZtwr3xu6lW37iROJ+ZI0U0MPc4y6p+NjBTsUnnUqlIKSEiw18rO091s
U9/lM/JFP9sVdbpNbNNuopVpMY2ZXyhNI88SPfqeRxpUhXoDI065ZgzBRDBkHZp+
OLdjxSNrkH/Ir/Cn0luyVdxRvt1/Nmb6Nd7WzbGasNzejiFd9KQ0hGK78jSBmvk1
BnsgA8dxB5SbzYRE4d6TplZP0X6M1RPsWRGRtpsWgI+UgKq0ug6ImrATHt8XXoSJ
hWfmJE/1DBVZRdatFhpMAlJrtXpoqcMsGa/9Y5DK9MRueIsux/ImNt43ZkQJ2vFf
3zwh9RfGBhVuu4jf0bY9N/KcV8wU3k4heogH/WkPix8wXVU2fftC/rEPS0UW+Bw2
EBaL3Q3C+UpbE3sIF4dlDocjgq3Cubi2YIOV3mON5L1wfO53k+2PUJDTlbUq/5gF
F/7kgPilGHDDfN2xZz5Unu9cZYaomvJ8N0B0p29ItErlVDdRK6r+UNa5ADSPtKBd
paWYHARlua26G9ipCm2NWGJEPAxZCUSBBgjyWFMTmJ0GmMbozk3SX9mD19U/3C37
FPdUrWTPRTkySDhHKSF8Ab7RMjZOrS6HqkxBgcLgOOGwtGet2a64KwIAZ5TQCis4
QVhZKwgV6/bOYp/PZ1X0HcQ/99bxK+OvPq2PYHQ997r7dA5Tryj6c9/ntHPMfnWs
294e6n2wePnGadXHbBlnidEJlR1QArl23al4mREZDZ2ewGS5lt7S7BZYz9Ym3XAi
vZDZp5TzqH+xzMCh1MicXdgJNGd+TqBcekafx1wFO91j/DwvHJFhftELX27kGQxw
Ntt/dez0Byt5vuc17UZo7havqXWCKISitF+QaeL7NrbiIBmNqGhmDeZeRtLlTD7S
wXLwRSqUK+PMp3uDRvrzRQ08/8D8QRBrw6qRXptOzLfMWavjexNSVAqUci9O4cOm
GZajeztg39XZXIPFrKLgNxxfsnZXGLh7OlzqbxwBzPV4Q6ayJd/69AHdkGAC8IyO
iAgb33Jd0HVEmK64nHc+DEJJW3EqRgbkiHp2uP+tK1XBBvRA9pe/dRNm1K2yR5bV
EVjPBorDDhHdMf2pOonGp6UJ24pwzI0fIbzPGecUhxLybZjBxqLy32v1Af967MBe
ES0svdASDDyCwmMh8vOK5fTgNv9AnGe0agwaC/RxNKhb408LFgNCF6SLBpZcOD//
SUoMZ9W5SHTitEHYPY8ezBzD9JF42yzPoOVGuPfvDP2zlMDaUMaU4GBvmMFc6Y2V
R7wj9Z6xo9HrKbCHBcnaU/DHE5/eIodST8EyIieBj/6HnO5tjOrnkjWfcK55Clql
W8WJuGlsxEwz2zvTLD9PKVTwJY/RkVhJ0+rA6I1YdJjkSOHesY5qjV9P1bc9TmbS
ZXFNjHTvmsFzxmjuhnVbUg3uVpcQLqV1v3PfdjwGBvuDadbkubQiKwIBbrCYQ9wk
P8fkQZenc19JaZcwRFgcqeRsvlTbjOtacae3wsKWw7QQtnwqzkED9F71Abd3LA+Y
Dv2s6XYbQEyVvo/obj5SgzadVcHiPbmNGsSS1w5lJ8t4qqvAITR03roHJq9Fag3C
5A8VUCeOPOWmD1zRD8tkHTaXu0v4+IXzIsdApVw1DGcHE7hl3YtI/CVZ/mEcWQsK
2rIH5ZD+oA02lzT5/yNWm7e7VNxqAYfUVhIhhYU93hC/+F/Hx/D0G5frvkU0kH9/
ZMPED6j6Ap08tYkAfv5bQ/WgQCFo1Dy2uq2zwKcNuHpjyVjsODa8tFwHHw+9kKpU
1FS5H60rWoqBPYjUD+A1ILV87O60/hBVHCfiegJnRgyxrNWcY+91nxsPdX/6wtVA
MKGswqRZ/tL+CsEnOJfzpdYAcR4RTw5Y6v6ReEdhtHg+/BwDwjEKHtjAOjXHCXJL
VXdIzmUtYW08+EQn1bIYdCPjvYr69YBpp4HmYwZpXbqrh5tJF52AhE+b0FANC3SB
v2JWjE/Kg16rvSQRwJ8OgZEUVe654Are14vB3c+isxbRz672HfDboqvOT1Jfdvm4
O8JiUgGAk7BS2X3O4F/p7yr4AjfW1F/Y+gAVgyqt4s6QW6KkixR1sA1nMVtkGRyo
r+6eR7s/o3qjmfb38A7dAW1KphHHj16bqkvsvIcYLRQqa7auNFmZi2kY4lW2A8Fw
B8Z+Ojb6xJZg9FT+bCfCnQIOeLf31tpAO6gSkRoYB0D0uSalvdguSS3c5zC8kM9m
ZKCXUFf+7jhjr+agX3ED8foTgPdA7fEC48yPrK4bPA5bjGExojOz7c4K6IiikJLI
zjaSkqcFahlZA/YOtnZP28y8xRanm2MLsdl2h/b1tUHwxUn8EJAeNJ9tU6LQxTey
8O6GEcelvx54AwoRAfGvps3Rs/5IjZXZAZu9gr791/LbQcAMiaGQ0Sl37MFyXsoP
LPYL5P0eoXJZqqD/q64lkpnfstfKbQ8kdpnunzcpKvxZ0aqH7SxNQeIoT1yVN7ah
3yVFczgr89RlLtdhVArl+4b0omSUmuHdZKx2HDzGqvAcxkAtSTRNRd6Z9LJDj6fE
qqAE52TzsmySXtu2RBj14rURDV8xE1klI+OYtpkOUvtHHJIQESBLYUPUJUZekJoR
ugyGlaf7KqNcanAt/tu8sInQ+O4Kdt0ej8yBHO8DOmCKd3rY9mzGkShnhVEkcjb8
hrvyp6dgraXpJOsym4JBJizgVDJp6KdVk5ADfwJ4Zr1BYpRrOw6o4OcNv+RNZd1s
SQTia82K6ib0kIo31AKeBLrInEoV4fpMkJqHkhTZcVGe9ns54RzkTvrROl0VUXD7
QrXw8M9SEb8k7AZ6Hk19QxpJidXsv4IimEJLPqa9SecYEkqX5iM+HGCgXiq0PDny
tum7IQ920mcLTZX7pCNJ2cK6ZIrn7soaDV+y03zMzy/5fn94JZuwWdtE2+FzE60f
VsLJ7AU6uupRbjp9PhlKrWwgHg176BoSlb5K+LQ4hirdeowZUo4K5FnJ2/s6A3A2
6sQL2Hgsx4PfggTm95UyWcd1Y9BzQud3Nvl1cPC/5HofJB2dG1szXesk0Io0cYjV
9OAVGkoLW7EZKPj+0DRQbWHvUfgqXR9fFJ/SjebGA/bY+7zsnJ/PYaWeSzHK2ira
0vleUb0M/AqP8lO7G/kuK9TYoP4eTcfAJRBbo8DDW5B/7IN4s99BKkrT5dIpd16k
t82Rtoh4W5BhAyWLbLfkL4OoGnpPk88p+hR5q8sz9QCr3u3Jtuo5TmNg5FjV2fD+
s/YHCk3+CeC8j5H7aCLNe94is1N9sh6e8a//KdYyKp2Om7InhMXq1tzLCJllMAPg
V0fK/iVKwIzEGkZZssDuGyAgWU02F/1NTYnb0fIPsyf4jjVNBIlQxTAt7XWNjfBp
Q9nPKsZUtCH2IPhNbkz94ibhLf9eGt7IIubiPcL3kWT4kBpLHxo/Ia5cZnbAT/rj
txXqqZEezKJM7WnAANnezB/Wm3MSWiXkkY5dqZLhE/Snb+OKMzqa75tPSfTVlKSm
NTKFVzbSzVz8BXe8StivBIjQVZYsXdqecu8uySDNKoMoYXzLHKHd4/LoBzqd2tS1
Ymap8LY+dQvd4HTc19OOnKM5oA4JmsFuOT4mw8j+5Ov5q+JL2Bx+l3cSb/URQLNR
kh9n5xFW7uBUNwPtQckTRfCZ4+26GMs9C7wSqkskyLpsrydLQ0EU+Hled2I2raZW
4OsTl6O5OnhUwJvspWc7KnSqtO/5/6J++0cd0vEVpAcIVA9QqBAmsAyvKf+hUc11
M4GdXK6MPlPe3UI3HSdK73lrabQua3Y6ODtZbOnDDscNGO+duEEnQpRzINsRz/up
1SH939gkguDX9IEOb0S7Q/ciaJRAehL5r2lqbrq5yu7ITA4xvsolLvSFFi+M0lSu
RHzKmVEKMtjrzjiJdeVfIy1Q/BNhgYIZgBt791gnPLCqXMIKvTAzxgP0V9VEiU9/
PmB3Cr2r3p2/1yudCpfBNcEI6zs8i07FJoelbYL3796AAYXpZBptfKyQRR8U5zUL
Uxnty9bUm2WnwDqaJcwnlWSy+3glzQqMBqXhvgOQKPFZ96bOl/v1gcXfEhYPwszc
8k45cQFrnmIXFQHI1ZzazzR5UR3oz0gruH/zcTQ51oWF6x54VA1G4PgPrpggRftM
wlCgsCr2W7FejL7HWdC2uvW6m1gOtWc3pCBaegfUU6LfisYPA8WWGD24Lo8wxZRZ
4GfjK4/jtXOxMm1RmU0ZRfIt1g+8C69bgKhansD2baWkzfHEFg/ijvqQqWpI4PSo
bxiyFRZ3g3GKl4hFHoEEkxHX6kHvCJSj+u6wMnzlVG8aPlmglh03a9pUP9GNiF/p
I3xtrRtzjfilpRCwAz45tACS+/Olt9Cq617dBlZMyd0tCPunVE80tHu6PKUUnHnu
l/dO3yzehUoHqky75cbdOGaVN/oNhh3vc1QqSEbSNydCG3saVVZ9QTd0ELJycmIq
qwI0mKVz3HR1Ld4UwhPOI1I553vu3BxAcHPpwXxI7+vM0E+hJct9G75YpV/RPQKh
/OgxmUrxp+vQAoRzRlyiKLm5cYQMd9IN3qr4J+dLJvCg4cQQcTANKXfwify8LA0a
7G2vVCKGRNWBaZQO/bIFHkmYDa6t6JVOM3pqe3hdaEfLD/5sj/SF9H7IHwzYk9vs
wJk7cQvKcPMv0eh5RQbCIgedmIwyvGZc1Xxun0M0FFuRGDwiVAVxi6QlxGcXljOC
8o4zXLfRP3BcWPkIOYVZAX6Q+1xR5rgr+eEL17oigM2x8o3NvJffC9LzFu4AAzgT
e2Ur6mv8exuY4xGC4Ur/ujMOg/mLt9qmuiIkrifx2u39n1/lTrSccsB/CU5DdKlL
Nemine97mj+bO3LdwkVaB6F4isJ6YMGzmMwMBdmYvRkTsnbxKpt7iYGZmMzEa2uO
rXspi769sQTUI/pm7kLKc+hG0gTOdzarpTVGX+zYZadkKhOISABH+ldX23ruwaoV
r8mFDaG3Jh2cGKOKiPRAUPHhXaIcyg0YBWJac0Y4rFG7CTu9gSoXHGvfMjjAN6EX
gbUg/UQhIw0nj2hAlxCGdRxvfCPE73Pl5gDlXxxHU5rjSQo7yssLMXEXcjcUb0T0
54DBZ91S4JHU8PWFN8Gb2lKUZ6KtqDiVFeE0LJRmEhh6/CBUNkxwL5vHMd/REqtL
J7IPNhmj3I/qWliOKbPNvHUMYXybYeyhaPvDTqy41qlkTW181rnL/5jp0HY/+ik3
5P88O+2gBitvZJW1zMFYxRy3n/DQAIxs1wWdUp8x3iw2NST1ZbnKqgdbMjCE/I0x
B25YPz7Kve8cP0+1+mXru8s5X/i19+fzRl5yAHeDGo66pourAQX5f+pdcUGT2bUS
5/QxHDEF/i/+O1bukazqJoJtvfvFK8j0MsUjV82tU3NTMXjGjXr3cyfZgp3rWXE+
BGIGTj6rv6u2rpbX5XmlAxtcpy34+8jKnSnlVASig248bjy0E2MCaeePKO3BaT78
X5UxIk4XU+hhP9ofVKELTZc0fduqU/GP8zxW5r0zXFbIiCkwyU/j53s4BhiA9qF5
H7/QnjBKEBq9X8IRtLKtzv7uHvikGR6CcUn3BbXCIdIm0WbVs8/y4CCQybn8UnoV
emSp6EiOWU7uBRaFrGfCYp1TBwYApMLABywtZa53NMCjFAF3uv5vrp9TyaXjHkuZ
jySyAME/9V4Kx/hcakVhXXKHD/ifwJWYHv0zCYhu8E28fr7KOxJ/O4UIKKCAb2XQ
P58IpiX1vVSxodaw4XOkiXGgezrCw9dV8CMe0i3IQGqDb6DZf/iTzvcUfC56vtic
s6iyPiX/nIvW7jPv3INFzeKoTUeebqob3BGFX9dI2KyW72yxLJP8DPaMFXqqHeo7
EIf+o65uVCdBHVu7ogtMiVSc3qDBRjuqCaLjQQ5djUu4N5d3Vhnvt+v1wLyGdkDT
INdC82agPs4irp8dzI4a3wYafiR3VXqXJR9BEE+paAnqHyzEZ9KT/sOgZv81DNYj
meZwYqyFrs10VBVhHxvsE6I5vOFHatDroACcc2edWCCueOYdK5P2poDzPdTmD+0b
14kzr/Mu/x1eXAaclxaZ67xi0Cjk+3i4uWaz40Rn/gfuL6/Odh3yicuIH9381WFV
NXuHAxViF6T+rv48m/vLjM9FUmKqvTcU3b8p1+KMwruOq/SB+0PjaVU8rIDD2/uY
zxtwGh696d2mJlaGMHbX93WdUK2OjgvOfDvlLUxyan/Q5f2xQfsnfRz0cvHGytDe
yMDzYwQ84mVXnuLG//JuMslJq/69v6fFzDEssPCGSyvBbD3umt7dNutc4S6xfJTO
/+hkba4ERQTik5OwmANAX/dTdVmWkhuDjc5gS1q5dIfu06sxbGtz/LnSlan0qJRq
uLo7nY7rGco4VwjoLP9CpnDmHFdqVuz/XpTZHay8ssN/2mUkzlm7vl17vTk3EZWL
RCNd2bFLXfSvJdSMUQwl33p1DoVgbjxnxoFG/YTeIYP1OlA4v/ZG8y+foV4yxHwN
aUIrhbMlHRdqdLpHt+q5khJ8zS1ezzJqRNJaEJpyH0/13eclTpEoFcmmTeSxI7yW
8I1uhqIvhX5ifXTjcJ47fWOH287tlOpkhm8RllNYwS3cwiOWfAUcyQGOz6wWgspB
E78VV3iIKgRRS/bglmAXaniNPPSkK2vlBFgYQzW/GUjF2mRasSIivgHkktN6pffd
xVMxji+UcVQ5Y9nvjlyQPo5NWk6lkkXvDuHpcDaY0ibOOydYsstxr2ZsUcpuYTyt
h/0fd4rfIaSe+h7frIyjGv3BGNmYxCpbsRAFBd0RgHYrLWDws3D64Y1RzaJuEIU1
2Y37CmG6JgkpN6auHUvybGxMwRz/QLKSZXzxI1qC1qc2eCrwgp/K9KQsEFiV2z2I
EktkX+u1rvluIFtlxBgW73zSr6vaovjVSlrerr9TTKPKh+Pn56UlfHTKa1BmB4G9
wRfubAYXjf20NCMtk8rXTH9NfF+54D2tnBi4Ozf+FxbMTCSwZZLGYUF44P1ICvPZ
LrajkCs75JQBA+YdTciVmIDlnxHGGPL3Y2b1K4WX8wntsW4QbsQgcqD5mKo3JCSr
ptIyJmq3atEJnhhermybwYbxrP/aaLzjQHJVa1gqbjAOEKeR4XOSss7F0o6uiweT
omMWVNER4SBxH0A4zhtFhtENKxARlAcJEfLg8TxRJPhvarfMMzdSqDFW0GgJvU+/
B/cUwzNJ6GSPZAZy1FnLYAImQtIc3Y7rzwQsHO0UN54EX3foF+l4NnHHyafQ3n4A
GEItMcIxNk+IYSmqe1kJ9dNRyQ4mToCPIhcdg5nsOteHAPkHvsL49k1UrJxlErG5
VH+nObz4FFCxcfT0IxxQ0rCRfhURD9LDCFl7c1lgmo9rfmd8psyw9Invo1NCB0Q0
C3r57SIdm9X6gVgI6zzPxUNErf10yUPcsqCIv6zUHv3rZ+momEsLaPBhpz0L1L/e
EFrE2ahLpis5zfhzHNA7IwNPb9ZuvEWhCaplK3Y+qgOhS2+cNccyjP/w0LvroKwR
DyI6mQ4Xuo9dQe05PiWeHftrnfXuBg+pXa506cXMN20Gx9ecGoTehqB/ySmJfiT9
Uz+wemBddyERmiEbEzVDPw4vOSNg4dVAh+QMG0jP+bKJM8cqFt+Ee64CnzobMLhB
T/HAt7mNVnxWRya7r+t325bCYLyX4lNEQ8nHd2nSWFnV2AzexH/STjSs+kKe7I4/
kGRSZqmb/gZjKotRrAUfOd3+M1cZGau0AXN5dS88JokrvPd6iEYRUEkDPrtIr5BG
bqXGwEEpO7bBpFy/oJmaXybcc+PywWgxweHHpHc3oudJzVs2VDHOG0RxUkvZ/S7g
Yg0rLA19h5EE12GUktBbZxz4eUD1lZuWLE9uQWCMhe5kW+TIWKtJxnpLVPtvbz6F
+Yw2BMbio5XNdld3mFvxhK6/E4M1KrRm7iUj4EJvq3kHObDxQil5qdvjlxqeJkqZ
Z2U14wyCJhTx+eY48PwgwFF3BMObaEGxt0yOiqWVRPNjUf7R70gfv10M8HuqIZL9
CTlKKiGLwsyrHPj2MOmbEwaHMr4NPqxl+H2ejrv6//QoH2QCR9aBEYzWhWpWtxRC
eublTMNVWdHDZg0ClfeqhU+shH8frKdTubYgTzvC79WY8lsZcmJditqLJCdIDMaA
amoPbysafsu3r7HoWmhh/vcP5QhncjWD3j3jrkf2NoVkcK2cb3rO6CKInnLgKBGC
QTVB93xfwl9t7y6jPWRtcxORGihl+JqW7IPXQVWoWB8WWgTZ4/qk43/dG/ccFGU4
ncIYZbIpts1LG/5OE9KGhlGADWd961nwGZp2jSNCQeql2FWQ4pGvasmZxTWwPfP5
Uptwol6LgD70x/Ik6L35WlRuaEaeBit8D5NTDvrEh0xzTFgK3A6tU6AjoSZ8RO5U
KYc6khsaoqt1d9yWcADLeA5Rzd+zlwhYJQFGRig8EzTrEWdTZw4QIRg/QauF1MoG
Igc3CcH8kUPItL2fyx/M1D9nDU8KduQwaLseYEv35Ji4aCAbJkcnQALqXZAYVJIL
HCL5ZMkEwOndj+qSp3DwEKhvgaaYelVhGIWp3Piq8cU/ZLEGkJrOrtywHEwgtSBT
lsrWZNSDXqLCltNJg35/P/cHvBjoGYxtISVx+3J0dq/SbRTxfddCU772IRBn0uLd
WMURJ8g1/OChBTxT1tMxi+Y6/5+0ByrhfOrPujEY4cbgu2CXd0cVuhzSCb7MyK+Y
mizrSNa3xk2R0CaqmvX7BSTlYl5m4E4hd9FOljnYbFOWpb1W27Va/mv4lngqMV1W
hnK//dIHLUklT84szLz0A0Db5HZJVgZjVN+l69CwGHSJf01xweIb4S82QTvqxOth
EmVTH4vcIGlZHN87gbsChkN/H0zogcEDHZ4pmo6By1ZTZlxxn8FG5aBF0i4OUO76
yVgF+SfF9Nj+o/NiT0fkk3dYvYzKNzCfnnH2AXmqm5UuifqgkARpnlgbhxnZgxDW
9y0bf2cXnKPNViU/2wlL99GuJMajuH4injYbkQx3zOKQYmVpHvgxZg3i54vMo+Sf
SVVcnqiNT/fPDAQkx5CDZ+z7QQ9ayaK/euDupFCxq8oLqWTbYv2dm4Ar0dCva+G5
LloxnXjtoog6FzUC2TTmFGrzEooHSLXhNKCavap46ul80930IKo19kceqibgncRR
MyPbDxN/kkzCk5jWigDYj7asdn4sGTB921ADS9NuZpqDRCa+6e/+1tXKI9egePum
XbFoxYD0NLhHLxzH2DO67UK5AvS9pEjDNlPTzRcu1+t6DoIAVdA5dNPpHB26JLTx
sPK9rJ27wnISanawyOBjsbYEjJBhl8bFlIFkLSfZn9KumbeC1Jjt6vKUM3GNb5rJ
LYqBnVm/G5J5B290uDItLvEygq1qLVvjSjR1pkVCfOLs2paZIqnq7bRLEHKKHuXN
5FB2R90UJPVtNklAmlQPpINA18kLUSYvr7yoPg5ETSsv+xf29nfeE5GNAQl0ojhD
srObCAj1GaXdHVHqefLU/++rQKH6cymSBxanca6di9zyydq4IF8KJX+mGqkeV/7O
eGPhgBNorymWH0h+O52pBuonjcmUYjyZfuHaWxpUgQXPkX0DrTVUMMhLw4uzB578
zr3CA3go9VtklqGJtKij23BQkipReit2FnLkKaofWS3I9XMHRXVYMDE7n5N7bGIq
F9crZZd5pQjJgrh5tAB7qQQzDTcZY5zQlHZDBGdIsD5gPwH4d5S1RHe8sPitZa3n
RaPomQU4BRwGlQOSNuAvqETjEZkbXjtWn4mdYHPdjFE5nRa0JbYJtcGzmrFFPQrK
Q+9d02VTwppJ3GX4NUq06ix2Nywj0JgercrUOTUrEDmvJveBRqflQuWxSdD6c9Bv
v2whirIrlnV76kxicEmFQ7QPSllK5M+XFoiRTqL9Kz3zAupkGZ2KgtI09Dut3Hlg
D/ocR9Qr/Ibh9vdB6Vtjh1B3hpyGfZjmSp2agNY1XgVLEedf/0erI6PXWVMFZPdG
Z8g568yjh9laWWF6My4hfV7hN5NvB41qGQRKLPZHkdmgWC0elIuSYV+GBi6QnQ4L
S6ImcksD0Jqsnkg68T/enXt7KLv4HBS8JVPf8fPWRRWsXarjKWFL3qhNM2rio0jh
DN7/9aCNsCTnBKRKMWcOjRf6W4UagD4jO9yFhftLP/2lbnLvqMza99r8id2tOLnC
KAXOLTQ6InM091X2bJZ/Tr+0MzKAt9tIJQTcmy6lDepasRfxuFfKLGOKCnq+A5F4
vM+q+uJBsul8kmo6UtDJ+kPeEh9UNV3+PuIW+AFjBWhJFKzXkNc7NxcTcoffDXsc
SsjIOJUhWStiBDmphJXygyE+CabHUyxJL/RwLMSbTv1x83+m7PLYphfkr4U0n5fC
O3nSn/piv22Aw0lA2xFfh3SrO24J3Equ5yR8lB6WLsIAPZYRJDUGtRV53GLg1UeG
muN/4kKAwROq2ryy1slwUtiR34NVNt9hiAOX0i5z9oeuwnitRmQM94rAPD6kMNWB
FlYxn7kAeynNSPjhdsqVdRbEBKYmcDx2JSk9wOZiR3+Dub5wbOW4Bx4L3hlucdX3
JOaBoHwDg4MkrVEdgu7wYDG/tGtYkPL3e/TJtT1i5cc+YGoykUdjUpqoL7+Z3YVg
KVdYpWX2voKxDBVHLsZPqXqmSquNBDZODMxM+KvnOI7cUge29+2ybAjMnJbXl9M/
FuiRpBIGO5czk8V0wK9HF+BCg0FGJSDTvOROjt7wdOtH23NeyGjJaLrsDzd5yl+k
DtA7g5+7jg8nWLMfUirjHjtRG9LWcv1X6lFLsVAMz0JIRLoc6Z7lP9B0/F73YvYW
7vreC3seXLri1hPD8jE6YRTET/ns03XDX4kNzIZre25YdmYsseaY1rRD3qQwJm9G
eQze7sxSJi1eaPNUSQ4FET8Pnt6ee/BqwdOSxkrhip6Q+XxDJvSP2C3BPissqNbS
Ogmv40o+ZEl9wfFaX3p05upucd+Im14T0DcS53pHOttTlxzTkzHa8jUizYnVugDz
OUfSMHXVmcR0oPTkWgFiAPqGoB0OXhv9AAz/tRQa3eZQcvDHaOptBcNY8A5N478a
GDLMKx9pA4rKuud7b9gN8256AdDHeq/WiIwdxLmTZD1ElImYBO/qlIrKUDi7SzdF
TF8vxcw8bZE/I7+RF3Vu/TnouaDF4FIUZMTqX+q1d8Q3FJ2uJ7ScB1mzPGIInhkc
mz6flZ8j4FsFEjQGV32WWbO++nfJ9nxZ3XFlwYHXuL+5IG3NndTLZLCnsfu+hLXV
wneB1ruXhr599mpnRfzFcI9svnKOSG5tOpnC6zr2FPwe0N+qF9r5nzTemE6JybcS
7TT865bP2aMtCtdHatFAwOnLcQ83IUHtSfiTFUB2ZGrzPjwHpvlZRVti8Sc4zYb9
cDeydcfU+ZN86XLh4g6GxWP0JrX7K/QdEkjIbLYR8ILEbmTS5f3uLXpb98IeiVCc
M1iAWR+Ey0H8wrlZ8mZr/fYqBHTb7m31CQaT6Kh5SpxsmVDyvOT8El0R1R/UKenY
XtBwUsoQhGEHdhA98UbrTrVbEqOil0Wynsi5Ooeu8QsAPkLAEz+M+xN/JcoABT7m
Yy03nwDBWuY+FxSlEzVj1IJyMxyxDx1rRr0kubY9BmudVD2tHYjehxz1o378GQ1a
Cp1vFumyuLlPegoAuwZngx2rmsZ5//CAHA2MpWkj4AYN5/WdvJZf7mFUVSV/qByO
jBLUfhH2jCobH/etOXcLnT4G/yr9EdrEpXBcChDRqaTtzoT9LH+HDZtHfcVjuB2w
tZXORKMHeWSYNvf5ChU9btBBD1R0NLGcW2sDWPg1SWqLvUXtfqqgb3A2o37TZ/Lm
flDyjI6EL1NJfL58LOll9n8qC7ZumhjoG4eJw3BHkF4tjByy11wScnlLb1mFGZ98
HWTB2GOSVUGGznOwLItP4yUXGP9fV/ibYhOadaPDLGRcO3pTS7agSgCsGw0xPPPN
eqMNBUTFAV/HzZsCkcJTRKoxrKUYKCtyXvmU+FGwQZEFfaXON4zUFPOOVsw0cuNr
ZZSG0wqmR4jVs7rit28Q/ZXnj7YIXt6LvCrTKRbYS6syjx+QarcCJVUYaQnh7zHl
+ebqBtudldrRAJCRoCAE9xJ19DNMgohbKCspHRcp/aJdUbmLit1lk7Uz54fclK+H
XmxfZzo/v1ZvqjiTLqPGmoKz5/WwSijCsfALpJ/Coh8WDt6LtYfGcMbomY12hoCV
y56/UE7MJBO9N7nSAqGnkvo7EC/jAUPOLo8Xu6myDq5m03Lpbpe+lOkkMSIZdp6i
wAnQWkuhIn+idCEawhOedU+VKKTXaBLck73SVE11znLQK5ZggX7KhBF7pm2v9ryH
e4X2xQdWezP9EK4doEJt5k/AtCdFCY6EbS1ihBG9hBxPG/PTntcuvLoAfFYVfJVm
JOJaVyurVzqkItqI4wcCYZovXzEkMmjc6tDiMW2Uggw6yEWB9AtfLwVHu+//M8yg
GSFAi5hsKoPlxscH0w1MiiIpKP1oXEJHHma7q+Fj5wLZOxDbn++lUbgm6HqbyZr8
7PEkwautXxE11Vz/7i7ISmxJyjxvl+IpOvpH08Reis86fLPaybCs+/g5MW66fP0n
VRCWEzErczYet3qrBSlJpax7SumfmNxZ6ti/QDzVMOqccByJk1I4hsyk9WeEbMxx
Kz5gzGAjTrwNB1ZgdIhjsvKdjZ6DW05YTzZN2QWFRdT75QjVzKXpy+1PDywCIqUZ
SfS6Xp5JqqTQAE3ja5nQ7AYHJztSdcz8iwCvTCxm3stbFub7MGaiKWI/4cTl9Z+S
a6gtu+DJE8U73BCR9LZmqDH4Wv03I0/1MWtAGRyFdLI64/fIHG2bXXkqQpuKwwHD
9EW9Y/BYIatkc5Nh42mO3MeA0PLG1zoJafmGTP48ZhjG07B3Wipmx2Cpftq/veCW
C/0pSxetyffYmVLrpqFEvdspAGBVcSwZQab6Xf8pLNsJ0VggQVgFcxWJNkxtgoch
00vA/Of6MevGB+IbizArBJttGw45ZuLDdAUrz7ij6fY5GAb3YNfE228CJJZuzEgF
YgI3tLVs22b83ioTXt7nD4ln0/GgZ2pmvn5WH7aSC3G/4E/crg3OGA+s1mrMATM/
hNHLJO+Fyx9tiEEUZsN/Lu017J5d0LXQZ60q07PZtKL74ekugKLQuGYiKL3/HPI9
Ys3o/moPQDXAOzYGSTBD5b2EcK5vNr7wKiU2vvab3WWRBeXt0z3u1jS7KBhALqQC
gLz1pNPNhFWzyfOoNCtw7wGS5vaMPX+x6c7Q8ktirlAAIH84x/zV/xkORvmLl3bj
x/dPsps2Yp6nvMRtZ3eIA3ubTaBG+UMxmTRg9zjBYr3hEEX2kk4MHJnrFR/Ngxe9
hIqf4BHO5dcV9gdAok38m39IlW170NnTX+uK6grbzMJGsWB6nu5sLYoKo4j7R8YT
LHrUqjlcDrVjCQ1v4+smWDqR5Sl4jECAidJmxWOHdduTWyaJHKZ05GnFbuZdN05Z
0MnwS4kdgLmprGn7xb/zeliqKjTurHdUHu6BX6guQy4AdoPEE8FJdq4Kfsl/BzCy
+UQgUCLVUXmBPR73w0ZoGjGH0KMX3uPG+vp7AM9lVXlWlCf6ykHxDl6s9jKCCsJS
LZwTJxJP1cDahCr1qVG5kfP/7HEVo/bC0ngHEGnVpKwstFsTELkaw/N4wBFSQcrH
Lvf8niMvBvwBJKxGgbcd0qWzi3NHysqe7Y/5pIMF6TX+pS1PeohSyxUr52XXIyCj
xPAI+urJzIOjc6yP81rzOpEon8+Fwzd22h4gv9LPRbcN//lcGOm6F93IQgmFAKb5
pERGkwYbOT6eclni+3p1MnTtaeQW2Yp+GCoLnxpwU+dL1G8+6qSqFBd+hOh2iZFD
zsAmphVU+bVwxSKEL/Y8cH+yNZxMpUic5xoKgx2dmxD+CklED0QGcwWgRFigwWt9
rwfYJYQG8IAQADBtsWwAxcNmJnhx6mvbotHJTP6b5jriGS/51nvdN4sT6ylkEbou
6FIdfoSgHeS1dTK8EECnd5DYXsnvjah4B/6VnFrs6trqQoHEPsw9w9qVuOW776r+
tFyZUkhquAZGexxNMhXq51wmIEiQ6OUNhnICMXPXr5Ij4A1V/1c83JN2I/XP3eiy
1Q3qSKT6T9LWw0SqkiKZcUepFIkbDCxljlrlAsxnqCx2LLtL0XJsDnLZO4ytJi9S
OInEBw/tVn7lVFneuCLKT8L55A1B8crIPN97gJZtwsQ2V0MozpYem9C7pnnMV5qm
KP/6jmRslKzBMSJj745ROuWeeIwWebDRh6SMlDd3PGOuOTm7qpsNGE1gEzSr621T
jx7OphQ7AbyNmguIUC9in7d0oLoksXDHobdoNcTGU14froHNuW3Ph0yBqZ7PDKtv
cGFUmGupgn3UTkUaSNFukfAb8PxY6IRT4XANhoefchUub9zgVuf/u1zVYEe8jric
sWY4BKdC1VcKPgZbyZO/kx0+3pg6XBEhwGCdOpHt+qa4HSOIsxNp62oPTf9ehilZ
5TIOK2S8EY7i2gV74/OqlghLg0VNnY0D9FXX6UUKnZ4O6SHKtnlOuJfjhS5hotYC
bH4JkrlHOrLBxXpaT9h5NjALk6AhiD7bR4fOWPpHpHPoiaAWbr5QNdkNL2odMrlP
TR/BhdX1e3xAkjWbCzpGuT7qgsL+CVUzFQ2eeeQabEBWYV+ks0BPw1/WwAda5EWc
qTkb8BR00j2z2P2mcxnnf00ZuBY47wdS02UgYeN1j94BNv/xJRtXWxukdb2lmQPZ
zcoo2trvCzSaGk/HYnUDElGt7lWdhNWK3cak2c5znj/PF5+jBor5pqPNLUwlkOZu
AwaqdXXSKKDCDUVXNaHZzjQF+C0OrJ7+BK2gNjCyJnFL83GnPC9RVoyQ3sAtVRB6
/JTmRqRnlfCMl3jZ1PZAiKvld9GXQ5QrVlkWi3c+HG1i28wolSM6e1Bzvc51Rvp0
Bkkk7pF0H5Lt3HQHAwSNAtSx70LpE/UBvubBK9pv4CFO7jc0gFuTp8l2izmdzVel
BptlmlNu9kyNvCb8dzimXkc8j3nOgmzTxiJh2zIOitf3zoQIumMJWCXgxIpsBgL4
R6YQiEybqPuNNLrKTVEDDAceKmj58n+4WtGe5kDs5Ibt3uDEzcdE+WP4zPe/mGmc
43Im0a61S2az26W2BCK/uMRyJvLrvb6yYGakmsv8aZ54jIa5e3fzXmhPd/3JejaW
49TYmhmmxdiUWRrO2WefXEGnrsED+GNdyY+Qqc9pBSV/oMus0QQtnPcnvL+ccn6e
tFjTmEySiMrB2uRgrMjhZk0dlBi4pG+SMM0t9o10+TbW7nhgt4mF7msVOl//LekH
FY5bWCeLSuu1rt9J2RDbH4ll4ZFtln3dPhL24T8iOa07/z47W5NVeqGoWLvX2UNB
le/gj9W/VAsFwjR9YnTTAWJ6wJhy85yN86xoK9cBL0shuFFD5gjULz0vPpLKhmA5
d310WQIkXkmIJUa9vh2V+YNPOKlVN1eeB983LbePilVx7VjhYJnd7qp85fIkG1WV
Rd2QsEfmfBznwdU9Gm2DQ+EMqqpVxf8AhOS5XhPZCd0wwY0Fc52bAIctf7ZMoWvw
gE7KOTFxlr/Z8387HphUC4mHHXRoOIAzx4CPMUbWitj1yKX0N2yJCvNVZXB73xFj
gxVsKnNA3N2wXgvydArusLgNwqG2B6ab9h65s28P7yXLZgFf+B7bVrCQBSfes+0p
R0ku4qIrPsiX/8INgjpqVPqvt65eT56A7xKOPUv4ek11G4bCjfcPzu2PxP68O8LJ
C8aPGIazdCWLNPEjQ54PukWQtshIhtkaa80JwO+7jIap8QGVO6wBT5nqJ87+y8pr
aHbYc9hNI5h+0VCMxaHaHxhgEgmQbnnEVh9GcG/81l7VTHhZKomMSvBINolT19mI
5dAg+1u/PYRdFkaRT+EUMVTfWbxh3yx/aDDxx8xQH1IedkLbxwW6WRIj84iq2E2r
dYvKVT/cgGZQcOaOQt4wdKizk+RBTwH5DDQKHCDWuTVp2qaCDFTMw5WfZcS/5Mpb
KqD+tn+E46DGG4gfSNkqE7bo/PkFRg199jPeWp7UWqfbESWl1WvXdyItCCO28mli
5v9OrTPSZA52VH99R9WN+P6po/BNrzGNht2SEvt6BYQJuSMNyOv46fFl2hZhuoDy
DxxpxpA4TI9Luk4/5qGDMk0DOjjWxNTn1ex7Vo/ximaLAsEncyMIQvygI0/eSG6L
fX29w5xIPE8LBXAHcQf6Ni9tRwv2spPoVcG22LUJEfk/nBrpIFnHXrk2fnWWxWAn
crBWLsuKXsOkrvNP8UQcW87v2LhE6t6t/DRoGdWSDy6JdzYOQ1rbvstqK7dyOFXZ
P3abqJ9MB3QT6azh+YVWlP7k8HC/RQXowLj1kwTSwbN3nuCtP0hIOtUXCDmFKO8z
FxB9Yg58D8jo6jN2dZ6QvFmtLpVIniNY0qmSGqj7rClhqgLurwmntrldpUqgZBsc
5j8F5dopT5yv0W9n53kO+sv2q11SfuOWCB452MH4NT72yd6cNEo3XwHJnZttWuBF
lw7Xvbxr3hSfbSm7nvfM0P0oDPri/FlUQXnWhh4axwOYhenpgyA6mvvPCpDsWbQE
cr3wCWebEWzevPhM7flgGWqE+Z/l9cPONhJwqmUP4E/OhSneaGsNRY+AbigOhvUF
0842kzMcSrDaX9xrRQ1b7Awzl3ljjKg53a/1yFTfK5lZcRm4vqSoV/UdOeVP01Lp
sdztVmYWkyHcskjq3CT97jtZOzuXlnrVLiU3/cNBJiCD9+z3ixJY7uF9mXeJDyUL
kPhEJSBRbsY4PNw9LWNny+VgD114uYUmmCxO98IDczlyoYl66NW99EvblvU77dV+
NQYqcPD+lZmh7HaXkkGJRmKGmBIULZx/X/XAfdNhkKUUl1FKGeqgzMPKnE55dMjG
AvrEs1nw9OQNz5HvJ8ixpoZSfUu9YzwBuIckjWtqFzy332uAg2oxGOTAV8Jp2zdc
YO10TtcSMAyCac/jutgFdE50BlKtS+Mdqj1y9LOZxiE6/+Yj0x4WLegt9ICqwoIT
uyr5autppzFKDy4Rfknelp6j/C5c64L7Jrs1EKEKAzEl7n19MioqkcDnDC7X9lR8
yQXuNppKFoOfWkSyRd9QjIOCQedtKFIRB5oUQpw0Z2KlV5dViNMtB6+LNZ47ZziQ
8aGgo3juIRKYuj6y6prWpkWDecIAz3KQAYIOvc6aLMZuv9V6EHGBLI9R8nD9MEUT
x8zHfU87tgxi94i6PasZtm7cm5lztVOCg7CG1eN7dRIKnF5w8fovEs/+OXxUWNSP
2ScOb/Z7bLoZts/lrka1CnUIxV/KHE/hWecQsx+b9Q6sxfP7NSInip4xrk6Gb+fK
wBpDbw8+Xg6TXDGH9hGFcmHyGLW0EV64W/V8wooHJsqf8mtQZ91+yPZ3SAl5SlGS
9vR/QssW9k/oj3Il8yl+wpWOgjN2UO9pByeEfcWEoU0TrC7q6xDQV1Tmn9XxSZ90
aSGucNRRVR8df0mW//bdAFMMvm4a85TUV5djjwOqlcWu+buyZkMo4wjvnkSJ0peU
lOwboED353oc0XnYaS1/CpsDLYi65lxVyJCBGVOE0xBvmJNUDBfMD4rgc27hKLsK
/c343B0lx/fFLlViptWBhRXiGZYZn3aaTdXqvI8eBcmDSclEriMMIePh3hGK9PrO
3Hmcy1u0K+RKHR/xrHWeoTw6aA7iwb4hnZswf4aRQueGngjmdspf81+bdEH4FKsS
FrG0BJFt3OEcWdG04biuuPMeA4ANtDzarjpwvfce6drzgxeTVXhfYIG1i7wkJBjJ
MNUp45aNMDqRGz2d8ov30KgXwaYOVq3L5fKq6HE8Nl0BSuo1BJnt8PP3azVCXm9z
6y49k6VMzojmyMPEsbjdbOdH/8N56mDwNNJvTV4Y2hL7rLLCWzm6EUJ6nft39+ak
2pqIWJnkRkysE0S0/6n/1RAtlK9dXs/JS9XdbOOGtCvkgVybTMBWnO4G3dmwGoOt
pu0g8AyBf5gFlmRstWfzXQa0Dx3okYmUEDZZU9Zi57Rec8aHofa7kqWxT4TtuEaC
Q+4vVX8fm31k4HdiI4kDmaIpS8Pn7OmC0ycOjlI7pzan26CDaTZ9PfNX8LTZlnnO
KLdqZ6tW5R+bmVcgLFRrDpcdMlkoRzCjsC+AF/Gv5caNfiOEbxqZ/EuMuZvm8os0
cLC5oflBNv8wPEURccS8hNr9H/0YYNe2ecTKn6iH8KW04aCxCiFJnDoVv+vPVU8S
p/bXRREh9p2ja64BGC2qeLfHrJyGnnNeL/Z0snDIq7Gec7snT7f6RsbuMnnVhJj3
OEY2NB+Z9RrV/3keSYRwW6Twkcx+LHkF8Wcvp7QZjty8kWXh7X2CI3S7zbKG9PtJ
9ps+F/VFDuzo9SgFhfAYggOIzAnJ2llKY1huVljhF1xO8SoxF0IdamxGkwhyWIO/
gBVlZv+UnNhXi4L+rnv8sLVMxT2JGXPILtPOndCrs8LzUawWf/ah7aAsxFD1EInE
UdrUz7TNzbJnIUYRKIPXMtttSA2h6Fa8r42BatBAgcqi1sJiHiaIMFqNmOeYhT25
Nl9grbs57IYYzzg3mA8lc+9BtLdIKTxcyoBA17zQa59fj325+50M1yXOVusUD3OD
X61p43IgFtz26OnRLIe132xAat3CCdH5TEcC9X90Qs8KF0XjA0NTNr/BuiSgLJR8
PP7xjEf0UhrsFnZOBFy6vYbtRAtYc+TpnTLDeOPabbuGE0dwR3PEMIVQaUDK3s8o
ywmqCpgL+GuNx65gzM3d/FtfFO4dHLpnIHQu7JZjq2TWYZlFnW4Ln2U98jkKWXE1
DgqxWhFu3tw9nTtcQ67y/qCodOE1r4TEKJySE0UZhfnxPOAVTUseD0V9dmTk0ZWZ
dK8RQd5hLQsobXvhqIWsWO+yHnRor+Wd16r48aX44n60aVUfbbUeZ+PDbCJMPVP3
7OHvly4u1EbeqRotmV0SbU0fe9FxjLHlyAxEl/MATM4pkKUy05bV2c7pRdSzQZAv
rHKqAKMcQH3jHaC7mmYjLw2Pyr+GB+tcHbHaQyjZIUnNlfU1IFEv7ybY1ho71E7b
HvL9gw9j2YYzRjrNk843NFM9BOa0cHMXiCkS0mavqxMoBNMWyAYHvTqsXKn+f4+/
zd/4R7Fb9KWx77geVQDzxcx5z8DEZdv5QSxB01mKw1QSbjFeWyW5QgclTytgCFdS
f9j9ntyjlh/8qYx9YFLNhFF8v80Flf+a7aEJrhTULfRT2/PSP9/D3KCmFOQptVCz
ny7NO4sIPaYBWQlhrKC8vq24FTeTINHt1N4ALAb7Ere+luC6o7QFCiX4YEFY/SYT
zOBEVnsyfOcj9BnxRxkvLrWyL+TmVOQ/4JLSuNER1vgy7ofjh+NAkRipzOtlkxFv
n+S9vkkDJa6ngBZIzJsK+UrO4nvVycg5Wb3NKd9HXN+soyZA31YOmT5n5f+wMJWh
QXahp9+KA/SJQoEJT4PGoBL87Yv97+l9yzvmXgXrklnAv7XilJLCbzCkM9ETYrE2
m5JuB53uDxppyc4DSqi5ZIGgiEc+TecbFt19m4390Yv39HrJzm/+ELNsj0yTwPnt
KVxkF6qPypuS/ODxvQgVreM11+W1vTIf4vey6ykPKAH4owHTLPptEHwccadtt1hz
ZjnL0FFGaw/qfpoHTkQ1jCtUO+xZUfGWtqSLUJ9rCWKJxK/XDh4WbODstV2FryEr
5uFDcuHvnlWzozC0XbGpEa+QiVH4sAD1+1OYSwgi8f2csz/ah9nbUlTA9Lt4BR/6
K7OiIOH/lhFjQ7KtVH9SsvxnNqVecsCxG55bVGDey3KLdilWqNJuaxG45rqjcZRJ
v1pLJX0kUZC4lxbal4TCQCK6GSCSvoGHoUzlQw6BEX0xK3pfq8Id694LKKuwrxN1
raIWbisjvqZDArEjeH62Yi6lRePE/G1Qf4b/JFw0L8zp93hqKExsY7aI/vYX49p8
FUHt4oqx6pR7C2AG/QQVmPcr5hX+QqXE7DeYDzBQz8u7Dx8Eq0lL0TGEy1nF4Ry7
X37uL6G2ClF7YC9/iiulvsZ//eBlUDBDRoI6kWPBk+xH7kBP88cw8c1q9bTzdgAQ
VjFluofy1MwgC34Ttvg5/8Fx6x4ENbFLs/rzQH432pYcM8vXwFD9ih5CnPcZyNHd
++u8pnw9LRGbrM+iMRcSVDF1Z0oNTT1cI/4922vQuvB82k9pHHwybhD3mrTcGsax
xyi7ZXt0TnGNBm53nvTQd6K1iKiaLh0A8YbwqSTKVMhgtSIrv0/E45u2908IfrHe
DKnx+I0pich550AvLLO5jc/S0Kbu+w7ZBAiJqVsBuC4ACdzbkxyG6PhKdC20Gr7u
Zp9gzRTbFjGeXnVyuHWEZGvVIa1c0FGKvS3gmbbuN5ckNbHf8Y6ScP4tOrKzO46N
zrjcOzHOfhFiWmrUtnR++6v9CFhWdAcGs1pTmhRfIKGr31v+WOld40xt3NGJQrO7
QuSNt9znWpysUds8zQ1xDUQ2OjwCRaqgP9CRLvXHUDneAwoGNx/1FqF/9ndJY9WG
+JFR3NT7UODsLZsfho69ckqUlURbBQY+nHwgI0kcgXhiI36MXaH/chsOjbBgf3lz
Un78iOI5hW7XOuLO4kkPbCRYvsYlopO3L2RZMcPWC7k4lswmkNfnV2cfgTOCJOsB
/jr2BTqyCruTGtuTxLqH2y2SyO8WgzTbVWXQfA9nZycJEWo1UN4f0x3+1fCKD03i
DEIH0hNruzcBKrkw/K73pqpDQod+aQeLDLbZI4/LbjfJEWkrZrhzfR6+i1EmC6Cj
yNaUDUa9MMkZre1rDIsivoaSFulWZ8UgAq+I1315eGzJPP4u6fS3qFxO7K77EwLL
LU/IdUCSzJuLBKw2HMnwI/HhuM/z4j/LqYva/Smf+YSS7e0jGvHx1k5q8ZTEyhte
F7j9aBtxhc6jeYEusOZsZ3k75bxBhX6/y1sbuex0Ym3Rvvu6EmoGPEGcs/nSKR0n
Zxmjz82sbFgiE/k3tUF0ZaT8Wo57f4yNbx17KzZCQESrMesMxCNF4dzwla1b2fs5
Y/tdikel6dccnEPsI4EOAMDTiMW9BrE+nzasml2lN1I55uewnsLuHdeH7eYGzAK0
V3mAjdxQ8M16Yfz1Oq4MPlFM5sLiP56Jzu70PJrLt1tBheSspRmvTqeUXe+w9Y02
m54rtZRKWAuTpIxUaicISPvdBJhGSBO25lIinIdGz9R/jfyRftZTQiwY19VbDsYM
nsmd9Iryp46yNhgXpe2mbD1AcnHSJnQZC4UaYsMRI5IAi6PTHt1V4Qz/ZJAFqc+Y
8aNnph8EyIdIYu0LDWbCao0fLuv0dRxSFwsTN0iG5iibw1fwvY1PO1eKzpDwiSxK
DlANizrlX4yQKo0qzlhS6+88wUi3Jio+hmFvvB+HMfFAP/wyIUyJYSWgDJcZu6w5
EhWlCzx3nDBqxNs2UolHolXc+vHcDueBKqqKwdIUNWEVT6VXkOk5b37rkgyxrgP4
lyPw9UYS8rjbqPiChz3ZhRoC5ueZKmRg4/wi0/X4IW1BGfPhy1VOkpyQ/LupxfkH
VactEL54xa2SG1IHruTa7BS+bJm/RXsmnjKvTJ3rDyEVbUXW7SXuvJYJH0YvAEIv
HCR61uILIsadLlr0nGZHKYUMz62JP/ajJ997IOcLNXX5aBdkkqRbgrgeoeuSCvyu
QH223S1y8pDk5WMIlyynGDdJPokHBdtvIyjbUU62WBx0Q8S+0Y89Ml7c4+uPeZux
7AbPKu0CSAVjNKofhdEgPjMORKw26E8Ve+3j1XGOZD/S/Zv+26QniJdZqnAIFOmT
KaZClwG3+81MDAC0xbwaEiq1VF9sPhJlSMNGYSolHWlRkIvO0RmpSCfgjECbkyeB
KABjNmenSCh4AD2E2AUoDmurC0ef+J0ChenkdtYyJ6orLoy+eAgAqKGlN+0cuzmq
ru7eK2sQR+uxDKBrWQkTvUmhIRTyYDr+2tbKFRSRzzVqzkgLk2G1esoLncA+W9Cz
FVCfCrLapc67Ep54eDdfzskRe0v7/5b3GohK6/s6pW9vA1Cs5iCeD8hB1/gv1VRP
HdHKfWnl40HTUcdofPr6ze5dszDzJBjcW9diEECLM1wgdgvl1iA1Q/YNve+gvL8a
EEi79PFibdOuWIc2Qnn6cSZFRWoTpVDQK+75TU9lS3lJloAcL25EKTsYmO3GcS8m
K1qx1o211iXqGhT75gRiarVUuo4C+v56fgAL8xI/PiGxBl4TtVWaaRrfN8e7TnAZ
Q1ML8jRymH/Q2sSzLP5r18qqF9rgfcabPqHc14FXBcv7UPWCQcS7cLi9WkeV7FS7
iP2deeLvgYNH1RjMJyxAzxkrnFa1FplhEF4svedQT4zmcau52JVnSvGQ4b50BrkB
WLkOjhzYx9lh4MdKKnK9lSUqryH0FTy49Ksg0Yj4uR+QCOb2mWrQQBdbYzqIm4F6
pF80P7YOSLObSn9etDFmJWnbolUkz5cb2s+2lB9vgSGKa1txu2z+amAA+6xkPoYn
GqK87H/FaqsohHMARVyKA4NU7DpfbLYNzGpLWrlrj+7HEz37OgPYyDEws27QIWNp
qzM5847PofIViNScyeC9eX5qmf1Pm0CWnidygBfZoxIFQiiti/5IKEm5nJw43R0M
/n6wTsCTsditoheKR2qZBBHaPO3sLoY+/6nEE8TXv0rDePKtV4/sTtzWpH+KtMIt
luqTzK89ywfveqA1PvIfJFMjjWOilRaB88m1HEGVXJkAPf9NQ8qsQSCeVgebDoVU
xjKWD9OV+2HnJ5pBP4Wbaig/R02974QQORVC1GwSqL9Ku3olHA5GwR+Sw+DNdKfP
YkRgPHzksP0EWrvUqVdlWVDBOxUspexus4MZz3IpZm2vWOQYOxfj2GEQtXLncK/3
lJOhjSljN28x4EsC5MBSKVKc0c29l5zAeijdaoE2XavsqXCIJ6qFN+Ja4oiBQrEn
A3E3olI4UDeoWEX5EnQQIkJDiMgBnjYoiGXZn9HjGLfqbxWuqDxJCD7uviv1aTZQ
8Mi8gYw+Or/ZIrwlrafvXQPrhFAybl7tD/gYE7GIrTh/HksWI398PPdDgz+Jbwgm
cklV+gaFa3G20NVZ43ghGTP0LzFG+xvOpJ20LCGNNd2UO9+qNY5h8ZQT0HRRyTZG
fSXHrCSC0izWgtvyxI4dDfkqTKZ6mpT3GsTQn8+gSzpUT8/u2+PEC3rC950vZ9nM
dTwtp5OHOnEp2jwx/KvGGH4qUPTnK5JKb4mjh7jWYos+LmpIZzGHAJA5p5iVI4Hb
P9LywXlvXu2QrPE459nEXq3WsgmOumHyHdct04nEHd8uVVtot/Mgum24MXY2h6IY
MisuUGIagQtboF3+6xM2nO0NEsDMSV3Fy1KjYRHxwGpg+biNvj8DJezivucLUx6s
qKiTOTMPivNS7/132K3PkvhHXjtuRxFaA0GaWoy5kdOztvB5SJNxeWeCAZ3WWj7b
xkXtogjwZ8Swbb0P6z0ySwUT/XmCNlVVSrbaR6nMQFGGEWQoQJTw/XUTjt5nQbf/
ywFmhuC2TRnLNRRBHw8OdXIxziVxvVq4ztLpRkPREUDksL4lebc0CadfMVjiReNY
xfK7G30lmPjtZIF7vDt3fNja/d6uYNLyqNTilWcdX5PZxRY1xHzQ60MrjdjJgQcv
xyTtYLkhazm1hcupcPEeY/4mm26PpAaAVRoregD/im7JEbNpOwFwMWA8LTxCh5oO
gYjMHeEgWhL0D1iZuwVLZcPESPawO17eTxx1UfP1520QsEag9SgfTFzrfVLWjd4p
eIyZ2Vms+dYrWSvzXnd6C26eKKUZspeNN8JM5RqfvFmp9EdtxRG31G1ehxhAu90L
44tNfMknOnbKQutIvlTnzzkOvJ03n/dp86IGwIORU2Z7F87mUMIi5p21opJJhnxS
ObeoFS5HGuU+i6VjrMV5L7a/F9CXoDNnYJKMjP8z0wnl0nezq43TOPrWlVAiO9wg
k8yd0DIRRQXvjKENaDyl5RbvHbG0SSKDNtrzCNbYm5Re08BLaj3Sf80yOXXPAXKe
tl2TEgPaNgiwaM5Dn0kxiX7K7dk6QnO1ZjRFx2lALo3TE/MNNUJOxFQR1BVHJi01
UVvif55he5d2A0PEBMvHf+bWm93WNE2aQaigrToCYCTe7jEs+pdmYgoITvridrNp
Tq3uuhxGNSm5aquQ6sB8IMF8ktlC7d95AtdQu+Ho2szmj/46Hc1bjYN34t/vRWUk
D3AOrm/fiv8gwKzs8kCiWf6oLaIaP0Erwg7/0I0JSDzVmL876h52ez7jwAQDtIDc
Qi3zrys3dW3u1DPVRTby8LI18BtoInQHLb/9R1ZIna/4Xc8M6Loa6DSZvfMy18Xn
nKApE3xHIw3UwxEc7Pb0rSStMczwCLnHoAuDiB2qAWp7xvIPL7HKHwGqXj3b6KOn
dcaOlNovABNiTJ6RMRAfiQT16RWH5b+CN/YTckrUEEbJtLC1tnrFyZY7+/3h8A69
IgSSBTRfrr/AkcC1VA2EvpoLngkQMkr8yfpXGveosFr6Wx8bMvzCTxQUGz5Srgem
W7RI7IF7R3G3gXMz8TUtpsBhXxX6HYYpiZlLF2y+uGOJR0KT+tLzlVGaXPQpoAuO
6xQTsl5pnskQ+Q0Ir9jKS9CxtOxgdMMLljNWpFDj04fNH8sZFdYN0ZPqqpHYE11K
aanzPPOeOCAQzbZ+7/a7EBza7MRMw9UYZGYibjfcVu3vc1Kyf9Q2NX08AnRtEHqu
/aPpkfrOPxHHCJ0qQzazfGguzx3u7RE7dDMhkpLXcmAJ1kcfpRbtz9iEsC+/n6qN
w1lsRS3YlTosXT40XeZnWfKYsTgl3IrelHFONk5HbwM67b7DV1HnnXw+plRFD9ze
OdwpST4VgptBoru8AsvZ+AC18N0nLpAGRnQH+1JPtrgRxUD/ACUlTcQ/Af4x5SWh
2H6bN9+Rm45hc8yPgFnjiAU3FnuL+ooUOYc3a6OZj1iRPk0d1k6NDWCAW6AYW3Yu
INjcJfgT3TJMwgwRGobV2b/DOw2W+LbwIJAEAgyY6XcQTRMc08k+Vb7wNKG2XFMx
2Izx1jF8r26lN6ynVci5MTkpvE1XWuopqYw+7OdpGZ36YhV056hppIW9p2+RbDhz
wfQnMMx/TwNk2Hy7V8Tq/dfWynXQJWfqUiAgxtLCeEpO1H+lRlb6UBsYk2cHMEUT
Ef4RTC645KOGgwRVAvBYN2mwdYBAs6xUG1idx85fy4qEO98Nz9yXYqwb5FdRbFyv
kCYkVw71kVVGRb42MGh5Wc6ymfEcve6/5fdN9P5HGhDNlZCPmrcKVsqO+t4EHfQN
Hs+CTN5vD8EoWGQxejqJhMxShfKwRpeHWOPksnDwlBg12ocf+WyA6hHzFO9x+l/l
7pdzSSvP29ntrofAPeKxXxlPE3OzM0uR9HXEXJeLDX0HOLtW3kqqGXGNdBRzBRbu
i54evM2H7JrY4KKoju665MTIn7C4J2jKr5pGSIT9olcZL5hwVT4NRY6kjlTee9Qm
5NJy8vmOZQU8HNsu5DpQXhIoWIj7dw6JAXiwQj+/N9GMTJ0mvxVvjEMjD2kKD8gs
S1Qlpf4Yfab9GndNGJ8xWMOVNb03vlbKzRdU/oDOVsQiDjow4xPqluAJwZKjMqom
SFCulXKMeS1kIhwoU5TACYoKq06aYq4ttS1esi/1HZ78I/akt2+cx+XtByZ4qU2V
G8r0BYqCWu2W3HXymmQpADR5ca5BNnl3wX+p/MDqahmINcErjedxajBwv67nYZU7
JjfjYINIQ2avw1S0pE8h8x1/Q02dN6WQ4ge0y42vUknH6cUuEgK8vFsFj5ceGpe7
sZ9Yr2Mc5RRpZE2T0RXR8n2h9AelUs1Xwd90LyHEeW1rGswyqGBTKl+Xl2s6IDjX
3nLxQ3RY5AWm2yIU1GSpBpbxj62BATRFqdBwkDtZ/B53MeMhb+9HIJp7z2Xhx7ix
yo1akOO61LkOPqXgmNX68ghPgl9SuZ4PrWn8PLS7jWZ01iHa5iWA+sDJfoG8o3nP
ZChvQ+QpSvwwmeRPNz8XkT6TH++oBsoEsssgqkBFNj5B7NlmbBG2BvvLDLAGwtOZ
LBZSVib3azlk3Rvv4wYctwufuPNxVP7yoMjIuah3nqs/7RWyzLrUz5UCqwwgCXmV
BliPwQTAgAAAq0zz7m9bP1EBApnMCwSc8nABqY5+K3T2+4oXlM7qx29acM1oKrKr
QwidDCKwRAWoa72/pCPi+GbpFeTATOYY1ClMLuVc4ouYH5nRExCXipT9Ny4ip7R+
7irEv2kS6MM+iRYWX/sJtkyAEBlQGVgdB160ZyMwzYRbuBBFMkjVyxVXnHZrTQjI
WSiXeIp3ac4NAv+e2/6qCP0zAjHZRlvD4KyfFBXnvn15Bh0vMsOC2Na5n5c3H4RJ
CpOdCOGr5lftGp+J37+jeoAcV3kEkzE3nbHsFQS4CU4Jrhr6vaP1nk+LrwuXwGu/
8Bgio8DHdk07PVTj1MVsMc6jRAb4FGkTG1StLTWH4uJCiQSh25nZ+tMXVR+MhYx8
TnVOOPefrKtIM+aHC0FIxZNvleECq/0JAWpD2/rCimn34AKX5fzjM96Jb5gjlYkM
b7epCv0kixAUTVc/RshziM1bm3iOAL7dw9m0QXCvfj+kp0d5cyp72Bbqc1NlxQZ0
SIgPKDtgPiq0RAfnsMndnXDM7CAkr2laXLjpBP3NxXhbDD2q8ghkGWEme8Mh2oEt
mjNTYrBKSZjKMmARLbPNuLGITUA+zkrVcHsTJ53jljHPFA7LVEMl8hkF75KhYu6l
FNgaf2lZojfMhkfUdHGSqOfmpJoitQT7v9R58rNP5G6R69Oy7Fp0Jud0d14/7Eiz
/Dp8HSOTpmd/k8b0yoHVgD2LExbH2YIN/vSI+2XEoQovB7eQyHGbgmO//X8wJYeF
GvRyhDKDebTKvSa5A9/YyJLQ0M8FZzy66e/N0N/+09CZ6p53IJXh92WRUjbwmr4Q
tDrfGqp7WDn3HIlGokvRWg3t/xq3fF5AnAWgUrJR3+5LDK+DWBTWfY/OlYTjBkip
tlz0ScfVPsmCGB3zSX2Rosi6yLXPife8X7uqDhwbHvaKG09gd4GUIfj2fAG1iap8
xmxwjxngu5JI6hLFdleYoPWhh5QIz5tMMNLvCj9yIxQMOofIcdHdQsAO4RFngU/f
VyRII79kj0RGk6uSXB0KU6bIEd/XwYw8zlRaZs7T71ngVxiiGkeezskc+JPobTVQ
bn2zxoFWsjfu+GA2aOXPZFNXu1nR4696mjPqfGwDlpH5ARyxYPxy469Mx/CxzTlw
E64cu98xOkpxq7elV8Q9OhTAiInjut4aHcaVtkOOiMN2DhoLbQPfiDRD1E1uO7M3
9BLi9GNT2TZQuCumV2c6u6yDOn8HPfH65XVyTUuaQnIxeHsZhDpmZqL65/3oqKbk
/fOMYXaFLGXlS+xhGaA5/WnC5dAf4XUsaXs3kyf82CWpJa922Y5tDO0UmE0Ogl31
cfeq6nu+0YtTnuUi95Qx+OATyX4NjOKKwraUhq+kpUBUKfW7hEfY9fmDv23MOG6T
XhP8dhhRSZzDQRFgh32gTHxpHuGp0xWs9CXpw7/YlOQiMNVIyo4PXjUBEoZ1bgxh
0wu1cjBaSuKaFUa8p1d7dryBZ1BBWT+I3nayWMoDgL68mzgVey8JhampkeDwByHI
RbU+5uOvEf50aV8Xcjxzj5VsvypVu85M4XaQosTRp6VBHYa+dq2puYJc21t5lLEL
7Uh3/ihlFyqTS3Tt5KjmNUGtJUoO9LThclBgHafnOdUwdLB1O7Z28QV6pYnorNE8
FE4EKFcIr06CTBAKyESeLFUWaAChqU61wvjiOsR2TdQnCiuOxui3vEuuTvM0EBxZ
QhJRIO2c0XVGkIUwLHtW2ysFHA7iKYlmrWST8W7G8CyhHvn4ne5g/B+uAAO+vd5B
si9rTidNR5CuKYuqkObVotvaiw81yZ58Pch1/JiUp0njQv0YSIMTSUbAXz3IAZRW
0wlunbKwnuFHEQENkMKZtL5bebbZQ7rA+p95WBj/7UzUMDYNgw7Rk3nlveCmu7oK
es9dGKpkHr39Oej1FkRSUJUXN4OxSA1n9xLl9m7z0BNiQ1ws4zDLsy52gXCIY63R
Dn8XugcesZrubb5lxB4Q8SysQoshmrGl2GaabFcDl8cLQhkzyfdIlB9OIX2N5slj
gbzzsQTCR3nug3rM8LR8pxJP5PaB1sGO7X02F+3bQ0AIoS+vu54jvKE8OCb/SWjG
dMdpkRx0EiQCbsFGIKr7XT/aGu8n2SA1t9pcNbbkrcmTxQTMJHInB457/wTfSevt
xaGRCsnhPD4Cs9rSBT5d7iRUNNJyGV09TaWlenlMs32rzGPTqsawyU+iWzwLD9Wo
vtvJW25I6oNz0OqKbwzhlO2CFWpLcn05+Q9FgyFLLrH84FtsXN4Q3UIHFFGAmt1N
wLZXHhmR5AOJ1j7xvgNKka06pJrMVdUQdzo2rhSHIKCORh6y0F2l5Gc0gQBXvgtu
QBOKx242LsI5zhKvB/Z65GJCc12z5MEXtybIyENEFBSy5md1R0bw19+jk9qnMg12
2RWYq0JYIRKnASnG9lMdvoCjnp+GK1TSXfwYjshiePu6FwswIo75Ngod/PdE1/QO
Ko/VJGMPRvuUMxYT1nVEfYU6oxcQN4bS8fhL750b2PiQprFtBXEYBNEt3UrBODcR
PEeY8yRaAqslEICNiUIE/O2GHkTydiJqiATJvXsiAL2filGFQ7ECo/1ILQp9lGCi
6+aLvkzrZW9YqUM+cEVnCnb5scuSW88EC4FwQQU1DkUKAKPip+nbjSpJAFiHDp3R
nQg2rjx35EYq9LK5NhegBm2YPj5hb35OkbzpNXBd+fF5YaHfmYNLMvKfPmfK58x5
l/2QgN3+pPF7QFYgT7Tf4b8vYHMZ4riLc4vy+rveCE2SV2Q8bBptGSDAc/GOzW1y
Eu4fXAknLYpBLE/9vI/IcETJtdfxzQPPzMiFLPIdpysZFpbqHDZ04YQ2Pwgv8iPT
CeriE2NRfsY070eFjvr3jb1wzqwmd1JYpRwZzD/KaW1sh6YuZFAwC57N7zrxdYV+
1zAhWeiD+z2PKm+ZM3/+Q9knk27nRGVSCLEL2pffIALmvEJLB+asyAK6ldqpK56o
PaicNJ9UmfM2Bf/aRJUZLZHPuQyxleRMAWM9X8JUpye6XYtxxx+SF2pSkHW9ZJWb
vvhgazUuuZnhMtkbAF3ecUlKlCjhDs1bLo2er47MpG604cnfcAScq5uKg4GK8kNB
T5Q7iv/vRv5EjY9PRoHlQsAvnkrS8XeCvy1cFduVBASdrazZ3Pzz2gUZ1W28qNuV
YEHgY/sHmqfpdzs+kvn6MCsa9C2f3DFW9zJ8e8KLT9ytlumffqm0AkCGi9sy10Yd
KipFvhTU/2WAm2BU0CoSCLeKxaemC8kt0OfDcsgbiSUx6IR9B9n/cgupX6/BwYwc
2HnI1yfYuy9jqOK2YORukRJXvg+UrDo0u6+T/3gyT5ezXdsEYkWYXPYhvCGVqYCx
SAQMPA+tHdYA9GlYIWy5mUumiBRhbCVpm7En2OAv+B21sOAdagLZUm6WLPl8+62N
fDW4+KVNyK78tS9qcBGkDkAuUfrrndRKJjbAIgvhD1815NV/IW0KNXqSNklaTAYg
w4JQytQI4/bE3/RE4BoWt7lwAfDnQRoKt0V2MeswabW3kvUXvq0rvz7nzIouOVnZ
yzywhrhoX4PWtrTOuhFSCkEdbIx2fczrBl7dCp3lTKhjGw7c77z6X6/CY7iJvVMb
CXZR0IoEP7u5RcQLeWdBxnjTIK1b7XZPBZJiOXSHBDCegIULOH9TuOLP4A87Wf43
cyszq7R08CL19aRrI/4YN1PDZZsY0wFGOkF6zQhl8QSYnrvLAWsp+8hx6Ep7iawI
s6paLLK4sPeTIU7lSaKbXZTGceLGY06XYZ2+nN6BZ82meqsk1g8oFtCTXr2n37BG
fOF1FnbztZESuUFLwed6dZkSkQeem2Hb5w+kgQH1nlunR6fIir5lT8GF/tKqwWy7
0YzyT9URTN6X+eQODFAhpnKlJ3tYS2bQwxa1oe9Sd8G1oBRzC5HyjXGy3MXoYBW6
Qjaiknfw8Ta0P2V0yzIO5qV5eyJYf1Qfs1sHDgvS7qz616/y2hqsmDbdol7G00aI
kIrLWNEeGFpof5Ti3e1C8DY7KOHIAp90vmz44cUMk8LbFjoJTfXeiLRna0cuWWK/
SIaPio59KLwmRrrEFfQcvtELWY9Cx7PL4LQbQT91Oe4yqhD1lRjJkzOu3Wsb+kkP
1YBUBmccZHdS5N2BpP/Ld2MRXebGF14saYufO0kpEcWCdACYBKIVKWUvWVvnxJHf
0BAnmi3s358ogirPAaooNX4KmpA9oLla0gdxFFoWNmeWE3Vu5grbdb7WjaJyvyCB
aq4EtGVH0XJwq7dM5wMmQPsOhScZYQUWHTs/6b9bOmAj6WgEHbLORNIaNgpTLV+y
xVMgJ9ddUGnjhHRA4C3hF6Wt0oOUnYS3UfABpIZrZBszQXhekuslGfGs/XR/KhzP
HWGtpsjBRQ2l3STlGAWMpeUtrI/HUVWSc68+vNIfqPepifhksdxoV7JtTGuQpiQ7
54ai43b8fcLniPfWI+gLh08yy+7K/Vq6aGVfvNA5/Fm/LH6v5Sq8ALgreN7sPANf
HR2EqPXkra3xuQUpWEv4LXkbhX/KRMEkRXdkGqZgy87XBWwSWh7DoZBsbcNKPjT3
whdshIlydHtS+0wJMJRXV8HrrXgtpEPil6IoB+kuEnnSh5ZqZTq0iNr7EQkCQvP4
7PYqfDjHuPaXWIBn8eHDYJSkrlf6d+2DA5kF3aozwmzMIhVZIXGVfHQpJURk7alU
ktiM1HQB/FdXtpR0FeGwwKP3obsYB5Gw4nTyYHPg4DHfy1IzXkqm63TpcmUmA1ee
zKy1aHB5lNR9O08q64wAMwyKyCtFMrGGs3JNZF3dCUpQt7qpJSOgdTwlkVP5FanD
AVrLt6Ab+oTIQICzTxZ5zkZob8A0aCMcZKwGE9ezGXprr2yfLNqT1Yni1/C6jgTY
ksiujFd9LAWDLCarxvfIWxSLLUsnAjEXVZ7WOdmh0eSoKiyWHBJV6GRHl7OoJOvp
2IDKzdRjIkXPiH2E9hddBi4uvaYh73olsLKIRNPJDLQQGAd0MR3QADDCGUW3WAas
Oh72zBmZozXA8VrOexeRmsVhgdIWmRBs3F3/KA5kB8vrOsOLScR0LcT14rvMi7MM
mw2s9jmFfW88ZQ5oiGMLII24gwji057wPalKbvmqyzhaz4iIhcIXtqgWO+jql+K9
VTvkUYJy/iBYB/T42MwhpsSCO6knJeDiUTJkUNkdpcjed1g5/kiz5FpTN8/hnxDQ
CH46M3RiULhqnaDJVegHHG5uqTOPv4mhUCdgj++wKOb8U/mFBPeTeP2td2bCNPoB
KQ1UMtEiV0qJdlqdWYxWD3F470e/ACxxY1g4/y94NeUV6lT8nIMEbj/hGjdgDFA+
X574b5Udxz2zHCZd1jRnKTElJI/8zj/zunLz8n6pdTRIseZPKlfqR2U4YYOrzNfv
BTOTzavV/nquxq+JBgmLhDn1qoFTNzbb0FWfecg1C0+Z+57SSCuMBzwGQ3TgP8p0
Z5rVHs5Y2sL5nCXz85rqrfuy8W5wbTQpx0uYRXYjIuBmLgmAQFnUBKdsBJEP+b8k
rIzoa0yuCnHByKoapkWyF6EIno9wb9vixFf8YY+6awI30N59Uw+8p34plbfvDKWC
ztA9Qj3vtYprtAIYZcuBZu1CB5djKWndzUeiPiXanF4z1nJxxUfYno1kPqQ4r3qN
iqMbvtUWh6zFnm0T7Vi7pDlKw6RIvvZnsWjeaps6SXAFGPdyxUJukJtqDJSM6NdP
5LgeVHzwAN5/EOEF/fb2sgULJNZyQbyJzz4FDFSviISa3YxdtuFhzefYTYS+XAdW
8sUpEe8/Gdz+kE6FZd/U/WZVf6B8GW2DoV7oaQLF5KdqqOraVoUiyHcmfDuaaJm7
1kroTmIP62dQX1f3JoqU4emdy4G0Kjf9xA+OVqAOEmcyn16aZMKWzz6SPz9nGHFg
i30B4MG6rj5lP5Y0N62+K+pp0Kb4o/cdnVTnWanM4Qr5odqBsi/CB7lvRU08v6bV
DQQuzRS98jsLJ67rLIyXnBHMOCS7QSAlHolOpd5fUrjZ0GuMVbsJ/27ZnLfaYOfm
lMb5BjiFbcK2ymrNQNQy9idauxyYqEu5+XZ5oZLI+y7XfrdSguuDZS5uUz5itAFd
WD+JUs8FjgYIWS8CJ0jV5iD75VTrpV0yiF1cT6Zgaj3x97N8AyNmorLvZdnYBCZC
g1KqvqXJu8ZVhTghAyhT/TSypxNOYqsO495jnFYuebbK9xGoGXMtuVNJrOtRUIpH
10q7uurE3ozNZvVeVfTEj6BeHRvL5uFaDTPkZ+cN6z9HS+faFA7gl7DVH8A/RM1N
/ov2JvPKUPov09eUIGg71YPt7WOu60Q7jcHjIX1sIMJ+2JPYYi9xSmHG39++WBIB
PDqLF3SYPIwouNp9Gm/jP9+oIcG9M99a9NedRLc48XNdcGDFkgj50ZT3TMLjFEJY
sV5xXw7nLSKE7Yo8RWbqlbrl/isR1O5d4B9RG+w9qUaAxk8JaEm0JCdoudkzTZPg
0SHHfWK828uLB/rCWaoT4dODKrVV+RDomD27+W56vqTx0QqqAUGUyUdOgjbIi/ic
CUlSuAoMYlTEWshqk8uHM6kAgAKYmjcFvlW302dUabbpoijCQeKIW3QNkPw0m0F1
f235gkJw4pBaoky7ceUzC0gCYQVEZj/xANQi5KgpsWuNw1Wksc4vDRtd9azj5jZz
9uz0KFsPKA2DYAENT611FJORpev8zwJLCuVfbUWLl7kpsBH8Zc2ILbP4r0amPeIe
seGSUS9+Bv3rpcwtwtpvDqQGP5p7/mJUBtaS0fudklmHM/cO7lva2GKpaZ+0OWtO
WDizeN9hhMXjzZgiKkcAGedu2RqVREQnXssihRq/FLEGCkhUs1UrsN/rCx7eBfqh
vgWPHxw19TVynL3v4y933zu8LvMz+uXQ0kpGLR5OkbmmXU0Os2aacdilo/GoYo+9
MFLPOUgXQeyuqqSKTHhNB6B3EftZKgHTdbIjaQ3VUzmfeP72KzcgIhs8reuc0tK0
PDLthWm2PT5pxb/Txz7iZ5HKGLLGIEI4chusJeM6pDQ7ifCKJoWIq8GEzZwwhTXB
F1q1xqNKhCAarYqLyCZbXgmfpXyLL1BlLijIm3pVOd1QE6EGjYMzP1+yWlcGszdg
Hk0unWGS0kw+pvjfNHPlOlVBmruODVV9DLGkrcCwDWGm4FnLWZ8VNopPWobzdDeV
VLLJKojONGl5mTJTm8tYdH5wc/yvGBX4K+lDhS5vPBIHYBbD08wxqx8qJpPufyg+
C0OX618b/r2Wqb6CUPNscJBZAiAcpHU9sarufjHmw8Dx1KmSCS5LsRpJZHL5Fsow
IfEb1dkIopuiKH36Y1yQBAPvDXpkF3MSt1tWobU1cmb8sG5X8QkJLjAbwCiAFfJE
Esk6DQxWulQ1khOEpkMeddahoKHFbkY/9XF0T/3VLpbcP19K/GmvxScXwgOj+cLL
cKTtXnjPPKAJTPuHRJQaU5/DcRRp88YZiJfksMRlu1idJGNOVtvJsCqlMbdNkqRP
2xV2RddH0dZ3/uTs+Xz6bPjWgksXIWD8OwtPlr1tqXWe6aXXn7j+1Jxk6IGMUPpR
UK6YlBOyPeDSstHHy6sbSgSP4VK+9Q4maqS2EdWcRHC6ZueFIQp5VSkP3JoEY1s9
ViwYJ2JTrKHkJ4cXkz954Oc/+6JNgHUIaIejUG0K26lyW0IHcNYhnsOgxHw+w6Cp
TDQmkSAtxONhb9yogBKwiAZsutQfxqkmkhqzh5S//7nOZAcbcWddbclBhTKC4+CI
mzqjRyK04pJs0ZcDHZzdWMHLlwTldDTkhFWb1k2o9i1JoJlCZlWTB4GiXUfZsbgz
SYn8sjXfXt8CMog68Lpsk/lLIA6c0vAE45JPWlMVjfdqw7kmfioLo+XXSYnt1kyO
1rw0gRQcZ+wHgq16XRsq0EjE2w9XBtlfD/PrpJ7VQCOjymU1FUsiQsmEx6fzKXph
aAAGol9ONRLdv38CDr6HO9y+yC0A0/SiypdIFkO1aSGApll8LyiUHSdOvfNjH1jT
ivsH3Sq279hc5kjhp3DW3xS7tNodHI2jzkecjr6Ul80v3G/liXR/oD+i0e5D39UW
DXN4iZdW45NaLNjoazOXk26gxpEYnVA4UhAW38Tn68tp7B5VhM1UFHJJzqHvyoA/
LKgdhZ6riEaFTC9boxuKwQrk0FZ5UPO5ELU8zKvSGI39FR8taCESoC4GHYX2d4xf
ZYkLgc0I9hS0LukU2KHWxaAGM+GZCwHUMDRnzEVJCFGImMqnQYAWbYLHv16/XYUo
raXIfsTg9XCfMFItZQXeGOHq1RtUCgJ94NYJmWyAiqoc4uPLzbLAsE7VDKvetdXP
sR2H4AC/2EN6rj9zulM0mYD6lLwhpfdJ7LLkfH8c8gIiVcXzSL618sUn/P7SaLDL
09p4GllfuPFri5xHdwWTz8j4kx0GT6/q+JOYXdToOuTEIfwVh20/Gu1LOTDTK0ro
+0ekcsVHMEmBTjNgIIAIUyHzJMqYob8aXncArHcSNsUiQ1vyuiKvumJMd2u+SkcF
W5w/BFtU/GwClISiqfG1xJpwAL2M3io58RTMeEMaZJmzOB1MBeu/6URkD4doSQIa
xE6bImOHokIfmUDTitxol8mSNISyNxjp/NTNYfM1PJyxonnz0OnEui2NcIQR+/E5
Sh/z8A7c9oGZhpbnhBNrB4bsX2w+rheLxxAM2KzCmT1FZugvBo2pYFSnFOXu6mXS
UmlAmxcaUCCfWNz2I2OyrDyJxoEoW0db9hx+617iJVcmmvr1TFhDBLmuPCtKb6Uz
mS15elWRSCCsn4d/3xWYzb0oQHEXSLnGMq/wD2kJOt+cKUp50PYXAQi4IbcSjOBh
uFVFTpvUieUCR0wi6QkM3G5A1XFgjdM7AvV3LbLHEqJTNocBZax3EUVn2iXvfQw/
8HARFKJ5HeskKZE5cscoud0zKE1VglqAcGgrETKkwOmpugpRUvieFuKtl0YgjrQq
aKEuWsUZTpSqevZxEjrykM1pbQVMNOBWQRtZ0nuhWpSemRrIRQSmgB3gP2Xwr/03
4CitATt7BIOwMDNtRrhFA7fkDP/GHSGz96M9Hh3RITpHi4Wpf/FW+T7WsEViATza
GJfL0sSVe8LURRj+76iCICYpYxgneGJ5DHiOF2A14ugdtEyBLEz0LgvlohnL7vJx
3TmXaBysI/FX/4oRvbDSnXhUEpv/xvPGq/dNGDbDsU35YW77kfU2enzVV7soZcpr
E2UmWCPSgXwKFKSkZnAXNDlr6pz472KZix9jsgWBJ3Q1NLs1LTBF4sFzKX9mesZ2
ovQzMYmtYY2D6/WW+4ugilhnK8S9q6pORc6OpIO468eXIgiKXWTL6VsR764JK3at
yCpfYiW7DM7tdaKC2oO2buotLi+fXnAn1l/aq2LhGZLBgCZB8K/iN3s+FLU4/toH
j1psmxZ2BY8FxmLVQaeh8JbuSkjegmPHSJ4u7HEQgFtPL23XqY6yV/jNH4J4PkHb
NxYYc9CEP8nZ9m2qtIcYonyZC+6GJ/V+KywUTB4K/ZYPIZGBq1j2VriF7/HJ26zf
MMeTCKa8kUfIKXwpmW8dIlmZLFM/frBoKUQ/DywO3ehsLJhbn/UNl6WecBNqL1vq
GfIq5m44Sx+Gb6l1huulq6b77ZQ9Moc4fjSSFkbHQcfy7ArKDeHK+qCdPP0/k0EK
sDo3VKl4JKP9rsHUajQrhkZrqD79NcDm5UY7s6oHrDPh6J7cpUCzPjM3pizFkrGD
hUk5qlJTkWyM19huXbQGiTHN+u79Im99OHYnJBN2zTCbuIvcgkVAhzgW2qaahwv1
EqRncnoh6UvKEikbDnCFOTqfDJAOl22SNEzQIA/VW+tIn9/g/FJGE7eXhOoRF9L5
g1/8YIvZ/7Aj1hLAdzsOnfXXFGAZBjFv7X2gNTMg2Esn4tKVObLdQZK5pWtOJhUJ
IMpi0P7lGFm3jLRzWVfOfNklg/F/l/XeHTYjMehPybNCzFAfsgCTLZ7P59c7Faom
xW4gHnY+tB/qxu4kCYAe0LKatTO+zc7WJKG7deJJ2cCHh1FiPHmjYgjzjz21QDc2
XmFFbRgGp9wxz86ZC5Uo/+pQ0lUyDpbwBCPZSOlWy/aa2CAZVAhb33utMLnGZz5m
Ks0g1rTFNuhsJTpLymRBKinkjUVFiL7nUR8lWq/UtxU7WymlAsmjuPrTdSfx6Y6K
E+9Twk/eyZ6ktOZIWGQOzeVNJ6iodeVCRGLQSBuSxDHQF8Li92mL2/2wsk4FiOpl
MD4Bxwg2kfnc8ErVv1pR7ZLs5xvyP6la8BZ9YQMusI+7Agmo7rf5yJAnqCtt+1bX
ksEQUtVaspOKUFzWzoiE0FiyCiWHgTDvonEXFrZGPqXNnOtxwDL3cnzY/QNrdRkg
Q5/KMs2HNZOxZAoCt9Dm/n2YunaXwg0TNP6f9hO3QHGCtI5uXz0jsG0INRetiSUU
Y9y5VUlXPCpwocsugFmCLsHRB1KTwywN/rRNZl3GmsNrNZAn8TaLxmhLUTN4ZpFn
aLMz81xneoweDtOcxYPIDg/NzPrXxmI3sjjY79tE1DsMzsRG1eN8FnAOXhm1RsbA
QhrtHH9EJ76kwWIc+yDwig3/woZYZ0SbGISKDEY2eVl8KA/Y0GQCgrjZPFo6GIAw
a8+FLiArTz4ndvPTok2kniHkwG4HuC/8eZrV+2cEHDiFkRVrRrwmnmBn921k7nEk
crl9ELRpejlbCEzrIAxpiffhlzCQed37GIP/LQHHlbVXTYbjAMXKbADkZ74mmhBT
oaaV546FdwOEnf7dP4L8UOjMCHbnELxKWscn2IrSwe8bK8O3LokU8WsPakY8kX2O
VaF/QV5vW5CweDA4KoPtJFB9mLV23RLpc9HL3EXDILkN16pdD6QI/naMDQIYtwuU
m6PXT6emGGTqV9qhprDVAu8hTEH7aVBtud+lNkDLjyan3wy5GJCBFKoloEqC4oMA
j9223hgc1Qx5B9nNZreXXY4rRtY4X6/mvflnOjjHi0D5UAcx5/fJiHIZwFcq/HHi
hF7yMwWlEEG8ziUoykqx6+uiarZmsBm7e1MFdc+pi9qgXbri5b6btKoKjPLiA1yO
lUuihz/uoKa5SIHpN+Rxa++9AYaTODM3asRUNLGtWKScyvDOheMNyyZFd/Thyso1
APvTmWHbxkhsHX4WSG8x8oCLOLFuSjyfcKkD+EofQ9d1hR+WCbXcTzU1DJMpbB9I
OX2gg9vnNIRM7M1fCE7La7KGoWMYkNMYI4qq+JB0BP8jPLn/+uQShzPhL+hiwS9k
GQOQuR0FE0xkmAG9CaN5q7v86f+lGn1r+yIPSjnAW5d+/eGMNF8rdYopE4CoElcM
ttzB//E/xtcvI75OTYGniCEDoPyFrs/hUQB/DZEmqQRDuQkvQoID8vHnQXcraKiS
niaV06ZJMUCCyXdbgjsI7ppJlnlz/FChLwUWxQEo0WMsNe88nlvRON3JHHIYPkFs
X4jon5114n/LgFVuD4qVUHiblT39pV1M4I88/YOHuCWunmYNLvVoNQ/X+9J3oHfT
HOj9THNHr1SevSyxtaRazTGgEnRRPhLhsBtfdd2F7ruspyeMKrwoUtJLTvK2JzK5
3RJiopGPxFNXhuxGvzmlMNR5ouy/njkuMqOWXqW9OsDS00QuYIX6mYFC9+o9x37A
H+OY6IGU3KyALRF1MB7maWaW1Hbho/Ea5042Y8yNhPNCePgO3D9dTwW3xcnzqFcU
RMJH2EgrP4t5SDkuHdC0+HPDHqVhWdfDUTVFo7p/QwGLF2zLWfCtbvyurYKeYhDZ
g1uh4RNa80sPdCwZtMNKzcB1iD4Y5abB20Lft18E+ebkVxqy+uwaL3uD1nv0irrc
Fdha/vzOyOhswNCpmXFBr/0FoY4jwtdMTy+kpyWGneEJJOZZOOhGX+N8KidRDE1j
gpP6I+toDIFgaKA/R844TkQ7Yznc99emc9f8zs4wmJDSlj9Y6mDVf/C3Vw0odW5c
awEz3gltmJpxsfq+Ab6ethTDZsQ9qLSUxf0A9qAl9NB1B91NEH9sL5eNSoAxttgA
LwgMNDr03xd94wlkoUf9jkn1z1E5AOrO1NA8w8Tkwkobz14s6fZGBkLpTX6fLcWb
wr5tkJTqPzJpFVUOy9I6Fr0qGUgPrUynTHfxcsWy08kaJ17b7edBYskHVkCqI2NK
pi4LhwHmY7/BhQmjaE1VtbbkhWQ4vdoEH9u5YfNzZiIGO4pIkjDz5hlNMZCUT0xI
uQvHU9PNgZwG8XzpmhfCWrx9HTeB++6ANHytb9Pwup8wdJKwmSGsQ6d07F8MhfAg
Srokl42oMkGI+ba7FY0JAKtzBNXm1gsRhqpsBGHmidUC+qt+Uu1mpUhD0tUlNQyS
efTC6H2r7kBEQdIR8BgqyBv7pWhF302UUgvsrrpw85klMxUeI8x9sYyhKvxy94eJ
p5G3twwJgH6744jngeZDeF260YQe8u7ik+wO3JRh1Kf2GCo3MI13yfZJfurNSizI
JHSUdFfmlpCLpnOu+9JJylaaZD7SXw5uzDdrbIgJHlD/wPPXTXDpQNGVCTRxBYxp
0IsjDR5HjK/Hwe29M2DqPA9nY2bEu06j8VyroOzKyX1lDm8zfBM0kBuXKB7d9wV9
gwsjv8oIKySMRZoD6jI8WhqkVUEcqDcySqW65PMAG/OGaEvKHSXO+eE8Og0gJc5c
+8GI8OqKbYx2nZp6p5AFSUPcR9zibtPztKsf/NOvreMjfsytUl5nVeukTHRY0t/1
1hFlNQGIFsC/EJksHiYJSPGy8W92TXcgbnit0XoL1ptEtGjEgiC0c2tEWjH+Mzul
6VdTdGH2weUifSd8qI+awhBrfdD4ggspSO11PXQ+n1EsAGPUCj8Q2jXbrWD6o03N
qjs0HdgUldgjH8Cld5wC6baO6jvQs4B29kdVBQX0YeaNg75IL4TydRif2NE43v7v
GsUagCidJ26nxyo+jRU0TvY+bwxJMDuz35Ln/KMrQH+Vr9Cv78FkKJZTlO7P6nHG
gEtdYKLx5RTrReRKqO4N+bpmIbJc7z9Apvhd5Yijn1X1Nd8o5OxCxs58UuVxUqnG
P4frbsIDR5OUOWM7S8rmHR7YYxcGv+UNZG7DiiwJRPiSdcsad6tvRVjTN3LbXoWq
vv6BNXjQWVuucNfEZp7zTXUBK8RH3m3I3XIpRH/u05ekH6cY0hoF++rZ7pbT+xM+
O333FLS0x5PsjsNuNJw9Xb/byiPnaICweAmcJEVbqZPOKZ+OSoyi8K9a8R5IL3Oi
oLPUJcuXTCRCkju6H+lent9qU3E3wRjyiYC+aYSE8Sdzs4JRPu2VlxqOb2uVUv8D
QNa1InHmGsnxRgr9RUuek2Jp3pEB4P0snsHErTZSGfe6xwTHa1ul7ot+DLYf4Klj
Irx8x7Ut7h1SrS3Co1svqlmZDqEnAXQ/dSw7h9hx6jXUYHWqM+As+NZX6bFdiNwd
rC7MGn84cYxjVIC0FLMWTRJulLS2IOeQEmF4RXNkWEYm7Mhh/PTSqrW4vZWwSzOr
g3U5sY6remwpr7zqStn++KZNl1WeAd1Z17WsiQTOpKHkg3tDps2PpATsAWVCNMPd
VrhJEjYv2FkgIc3NcujWToaX7le2PdIuWdHw01RkC9GQEQioJ/fbDGSgOwOfo86q
00okhDLYcdQIwpoNrwXkqlL6lLoJ2fe7Crw7gxaeRC102DQH0RMRg04l0GnjHDNl
Qrh052JbAfn8eJx22eLoLlsvFU3mBlHWxrDIkgX0PIiWtDqn6B4+694xpep252m7
SqThaQkONJ8AjY/T+P6HWv8lBDdxklgETjEQvfXFX6gptByHBGm5gEjeRW+6CPrC
bIurpFpkPdagXlKZqWKDfPFG2DEmeMu7S1eIlTUBJax8+IpSQXxAyHpEeuVCh1pm
D5jXnw+JWjOZv1QAhvfUzSHYGWNwj9n6rJSXLAwuUnpchlXzZzOu4Qdv5Nmy15qX
rFB8NlkcHgSx9Pgs7R0q9ALaisnUWgNNOvhZD2YP4lkdySkBF1OKU01I/VA0eQUO
BEw+3BPioZ58WPHI6roVV4sx6twfHxAnCJLOyL3vsfyHNtIRBREUcW32zDw41YJu
Wefh5lIuxnnKpQVGNt9lT/X4RCouep9zbFR1EurxLfjqE6w539gGVvl3jUwOB24k
thRCyHpwn+v+5WXzzEgqPEVufxjR9Bg9T3SEXBdpmkAiLAzv2X6imHSbjCCHO8mM
LBqQtmG5D0dJQnh/nHkHTb2zjmB2FOXqjLkjntYQMKSPXHoupHpzEcaRNF22+RL1
EdG5sN1x9FD+B5gI4LdIMttwwvC/en13m9Z/SnB8qwy3xTHmmdT1kEcfotLJbHav
QJTtb3smze/Cr4QcC/ObsW7kcKMmPinxZ1ZICL1hhcCbi79+RgsxBOWMgGyqmrST
DWJbXLO+KIY+Q1rDXIP7ZTYtd7cDd0frVme44iADedXmfOOKkDeHmWdAU7XmoPO9
mq5N8Oqb/LOF97hjWME8zK5Sk7CI8f5w9tX/Df2eaBue58Op3kslVNASTaJ44DkE
uf1ga+hPO1GaSebMBmkCM/DulQGUUK232ewiuh2ADqiFR0tWxU/Pzzm42PTSaJOl
TpKoThliv2RoOJ8zvkkqlpRjiod63+zwltuwVdbbiQlVXRjl7OY6W4U24rCnn38a
P99XlGmS5a5FrK5X9O+6DLnlzjLU4z5NRT3TRr5Cuc4KvFpPLZIV4nHVL5f11K9y
lgEmsVsx658pjVJHYKjJn0ow/OLd1PUrh/I9Q0i0J6nQHw7Er04TcpaLOYiglYd2
VdgKcOgqbZ/rNCluC/aHpv0w0JlShEJ7RUu1awGJGdpKfBrp7OdA4DZ/7kk5wDdw
umE/syX8HweD7ceRayFkpqRtgBBg5coug5uUCXBI8Hzwa2jhScGv4OKsFYytoK/9
VG95Iap+JEp+53Fwoz1pb8YPkMbLnii2O0hIcMj/a5wctsjLb+UvGuIZQlnquhDS
DqeUeNg2BHZA1s+Ftk9DADUMTucb4AZ3p91AoOyfBS5T1tVnEh5p3QLG05/Uw9hm
CPB5XCG5bl6ogG1OnAzT/5+z0+uB+BMUxA0B8GFaO5Q3qP6F1BAMq7+sRSEp5BpH
SJGsZF8PGva/EUTTxvGQIC7J0yDWKlBtWV13BHu5oFcZFLQQr91fUy1y52xuydgB
yCRNJscaEo/3MC+/B3D0tIkHWQFFdKZnK3PbCvlGnxJmk/SiADsN2CaTJ/2hfPT7
bk1HvODx1PXKsMaVWbvh05N/1l+C9NpJLLfz2gzOhDs8yL1Yc4aJ+pH3Cv4IrDpk
uQSDzr0gKpWhaHj736RMtQ4ax4cnGPCdJdAQX9kWhDrFUMwS5/HwjkM+y9T5MNtQ
UX6yqPmmmiP3unIs1GvsRwP0DfxlbB8GSANhwrANfU8mDKRVD4k/AA2WdvWRyii/
moWRHnvCqrAGMPvAs9JGwzjwhtPcIEtKvwARvJBQkZj8wPfcMtARaRpQiwPhGe68
S70Z/VobFNPoV9N/1a6XfB9/w5JoTEu5mSZ4CZHLXDevexVpNaxCrU7ujsN2SBYG
1zeAH8yDiLy509XmNEID+7VpFmimXbfxe4KcDT+gMSQCBQSaCw7ePYICwsXTbLcO
eT8TXiH5UaJkp/CY9HxQbFk4Ucwk5QkAZwgMImFDaanCYDweiWDhmPcWkGg30DVM
JNPllb8yGy65PHbGVlif7GWrPe/XxtVI47MftnG8HWyTwZFnbxRtbCeSuIbGGZFK
fRXz4qFTjQPuOpx0F+/y8XWyGmd86NwoVsZshkcbFMrVcDRC0U2rQ/DRcdG/r96h
UafnoiDb6ixUDKZf8swxy6UiJTkHnfiLnQudiY9BTZy8d1YI0b2bSo28fmIsqspT
3CHSDg9/iKDYstrvM0CV967wJuWvZhVIBbV4S0VhAvlZt4AZJdxdMApnSkO+n5kP
zzBlBX32Zei5SYfPmDkRcubM6wMYgN3lhh0ePTK38BX3zlJYXByz+ReyKF1JZUXA
i9tVFbR9Uqw2gVAg1ohZcWUndt1NK3/sd0YtMX0kNMHmGSQroVSY6/gwTGaNqfoj
T9dYqyaD1hq0iKDpUJ9d+QuyNhkiJHBvQid7QzjXEyTTubkbNIKZetBDcE+iHCC/
vD6Tf88skUm2ZbVfXk2HxBVngYJSVAXeZdTzwnescH2yAPozC4Z/xSg7u/LSqDub
TOVZIZs5EquciJO6WJaqP0JuJIWXNJcoS9wQqtBYDp8+Iw15mXrI1fit3R04ZO/f
XIizSxrQorZJRJrdLOIU6AajhF1fyjVxPUN1cNLi/L4g2tNv9s2xwT2HymkCvbAT
/oX9ZLRQBzA2BgD5cc0NWnI6DFjQ0BV2m6w8da5wyk6hW/Wm87D+j07HawytUwOe
W2lHc9ToIccJRKqRWs8gCw22pf1KUo1QqFkKWJZD2p1jR6iyLAidQr+YlCYuwYgd
9ZtgXxIJ0K8vUNGulE3P5jzr1v2euMj6EicJAFXiEcSU+aDZavOTu2zAmuQDgmVV
BGuITagJeqfeo2VcneZYlGrzedN1uZknCRTqLvB7ZH5LhDNlietSp8PEPpNL41NH
OEQ4ff9Zxmexk36bsrT0kVe/jjY1ufdnTx5ABZWMihzZ6MvM2EsurWXHHxDwgQ/q
h0C+kAMUg/KUb2Naf6vStdmdFy7gGn1AvIbn4LNG4ssiNnx+n5fkVo+isqgY9QzA
LHi7qq5IjEu15clUVaCTo1XjhdQIBsCJrALnp7s4toJdVvmqaKNfwpmcNLJ0UJ7c
s09vMLLWHE9Qsf5shhs0oOYIsDfLVhAUOK3fN/wtaEh2YzP+RUo5V7TBG7q4bm/T
YqqG0im5G/NRI1YPhgZQM9AdWKXTxEXVF8Obs2oIWyB3mJKkAOMgJBkYxOCCOdaQ
gab831abvtMUQz0liU5QCw8HbRPwKcCSFTgl4G4oThqw5aFgkCWRP5I0pSC4Cn3f
Ko0/SVsrhZdzX8WegFSTzjbHYCizmykgmOsSSIpS6vht0CdTZxKdQ1vYs/CaZAz5
Y+ZkWj566l9n4OowuZFY+nZPj6CapZLwC7Yaw/Xvw6pqeg101JkyCE0KA4HdKR50
2Xp3hAjpKHWW7QiD03ISK9TNNShoHujpbYyUwm89FS46805X/5W/YILM0O7z+vFQ
NY4vkWdY6SczZcr7313Ahuh2xpDdkERjwNh+aSwtVVuEwzEywmVi42rycLQCpzDz
M886k1K6Yfq4By7AkgdqbUqEyprTaRCtAR+HhXBR1xJrxpOWZ/XaE6vAVjEJHUI9
gh4iOVypm+Q5iLpO925WwVdM9f65rWTxAKvdlMBHlnqtE/HCOeHDb8MSoYiq0o2l
EgSF/qvG3hP5phaplo3IKnsWF4z/pUoCstUxImkoDtje8tPLTu+n9cbKe7i8Y8JA
qgz5CPr/2RStcwGm01EI2ntEXCuFqCzEcEjVlN9wyWhOAk26HcqBqCrXxc9FNZGB
6SA+fdc1lMMq5rQFX4KpoVxIAd+dSWGv3dZlTvN+pl2WRW61I5GLpDWX1rWIP1RG
C4hfS/CiSthBjszgRYU/L/oonkybL1WExuvhYWOmpw3NDMGwYqJmfkg+elmasjjQ
EaJGCo0UsnTvI1fmBxbcuvGFFm6sEv52yRlAZ4bWeGsHUuQOlX1XbPBrlcdvMPoF
8YNVLekQFkkYbCKHyXCtqfETuP4FJC1EtmuAuw1uLnprpQzCm3e85ha/xhD9CGwC
p2pUMLBX2JEghfT5Z0opQGnVeTKE4SdH62cv6YWUsNQ9XDd2COOH+OBg68uhnqky
CGf8rukG7a2jBLRR4tXZUBi6tv37ZM1KwICFEjLxT46B9Fe5jHtFIfDx0acQbdj2
uXbcsWzzJcx0CATD2adb6HdFObiwYEmgsWI2GuvhKd2tD/m6N8FRTu8yxMv1Cd9D
JquaUqO8owEvyBBtZXfWFY79e+m+kAA/gZnT0w2kaFuNt45AnxGASxaRnT7bktzA
uENQfkM/uudoRNk8cGXDiNuiqNnKPKXrQxi9PsoS7MNnsDBkffRgnUoo+B0vLUbJ
q90LsMOulKFSpHQpTu4SfF5U3QG5wbXCPKzXB/hNkGeZNw2mv1YrqfE9SJj+UUWX
g71THv6mqDrwhgPY45cdRxiaXdLOuqSWZCmhCUoRwcHXvH8DKbhBu8Oy0l2b4DLD
i3LPWEHdgeWOdhxntCWe6EedUMJtt9bOebisr0H8MfCd4wkL9Dv0Gq9GDdDqjHFS
bf4LxI9tC6yyLDEM1af3cHKoWqHmk243CqasqaffAtDORXBR8ptdx3Rs/BrKavrP
UmZNXdss5ZAjBOQUnAfB+UKsnU8mTlkz79XeULayevNHKMh/goxXkUU51zlxAuKI
59wpK1rYNHPbj0xg86x90p6nKNpnPihfSzGnCD5FZ9qFJRKbja/tx65+Plp8Fw4j
PKv5yCJzVKr6jWd5RMiN6j0DXi0lMgt02XyGA3jt/v9FUHg4hVFDt5vlDpN8zand
sndjs4r/O03vU1FLnFV56Wtpt3H1y3d069H4zrc/IHcNrAZ2aXzu9prLRJhAeKMn
/gG8k4VAuGz8TcAxsvUOSAG2osWNDApVTUmB13xWIe8kcXAsVVEq0sFqr6SX7Ncz
SEmXzR+G3jm/GpHKa7hfr/AGtTQMx/LXRBt6WAUnnjerhQmqyl69Rc/XqfV382Fq
rudrCS0OZLNycMzS4S/4ZBPqXQ0dBedF6Yos2a+1WrqOFLfAAMRPXfddrrYjp0N+
ZJlsdNoPx9lilqoVZw1wXWamOnn6S9SlNricwL7Qkdd713kP3hgdtIovT0lnCm+x
H8Q7oDHBa8kxuFhTrtDT2VywzR9Qm14hMuqaXT6YQVuklzd82RaXjQsbxnCtiXsg
ljRAT2LV93zZhX0o2Ggn8PXOaWbBJRbTiiEPjKYGbqPy7JzuGz9wAzFPX65PQ8bY
d4dNLSwdPM2MYMYZHvD5bmQCAaJRMdyRScc1C6wPIbxadvlsJ3eWH9NQsJBBmgiW
1PCXeVfcIQur+Wht3oz/dmDP7utwVvfQHDIdCBEpGwZVRTGY/aLsBXUk24hzNnWs
uQx8cCn8w3L+QvJFrmCA3dtcPrahYxa1ByzKlRGauJWdqNzccpW/SAp5YteHK+Zo
pjtIkm9jNISUswQA0/5qxsDbHjVngfzwXfoeOS2OLMdEpQ/2Q7LJrZspq/7+5jZn
xXcLxAbl0aIIltWdSiBdOMPtKVQ6SlN1y7a7VnmyqkWNgDnucAMOtfFGSRt/K3Ln
d/B+E61BFz67dZMPSenvdqE6xYIUh9aFuXdQ2SLjnQfEMxOVHcmaYsJlTr/mxfBQ
azFzy20KhYsrak9uNH+4/m+0+ln2Wtr9oBsSvrA6PetVqP9pa3dn3uNMTFstT1IZ
9CubKO2EURpe0ndkm5zQhiKbkZONrGyzBwsFizzWqw0NPbpZ4KcPBQq08ZSysJpR
QIPnsayTbcxlp7FMFBZPrNwqzX+RAn0U2yKJ/NFFWJB8sgtjtcV2mwRDqAVVKCVa
KG9AzuKv6rS8qU+qlznl6R+8D3CBu09MSO1N6/d20pydwfDAgAnCOGpc37Ad2lw9
2dV8X/wUGApBkIs66MUaJnAvvR/f4Dqn4AZm5Q8z094e+jQ9n4tPHNolTbWs+hGX
RCclevVhwVosKsQmoTo/DxNuUz42YcnbKNOS7h1dcU8y5S7UeATP1U2kkXcETYfP
jub3ET/fWDfqMEDBQ7aeqqk6d/Sm3yBMfjEQv+ABY9H4pTGghGl2WaV4UMySWbNI
agV/foaXobNoICD1NMZ5tmrMLxsvDqmqzCisrwC139pb8WR9cB2nBpUhA2uYgxkE
U/pR1MHKSjZQvusW5flRHYOU8fPiAUXMOCIyPvZgJT3kyNGpK+UdswyKztFrnAL+
2JzrsHgwOQgt0OU4OB8SeCjWp3CEnwDWmj8PZBd+fdSarDbtUqE3z9QmUWkW0Kwi
1i6tBTgYiO8yv5S+pD5axSIRYabYHWvNH6MIXXwjnfwBh/ji3x7gnC4+6R4we1xW
5dhdTY7HGTuy0lsElXCzncuJoVOV1XjOyUK8C/8dhjqbf87NMNg5aW5YNu40dFgY
7kd+6HffhMR7qG7LEUpSHPTKuJ/mhD+6yRoq6ZTE+nrdzZ8fmdKAzY9/sJZ2tTzl
XfolsTO8ywLfUpWGp03nAOuAkPirXCJxHGkj3B15ipBB88rLXzeuLrMRmouwoNvq
12fD8PBhVUXsPpNQM4eJfZ7im7MlyZ3Awq6u42DuFLCyOOSubHZ/eMqKrrvUyJzo
lq2UI/d2ithoxiyJgDYgMPq5U+d6CESrvbV8NnCMcFGc9xh1VxKHVrZRVo+P37CH
8vEelmtca7sPng1jl8qJvLu+bEpIaM83MVmrScHB6s7Pfy3PFIX7KEzsehPj5qr8
6uQPrOkV95c5UX0hWtxu0x8hQi3nio0o3ZoGKB5ywBPdVlB083w+eGiRk56oC/cR
VPwk++AqPwLILf2NrKJWod9Abwkwfer+3hz5UUopp+KZZiMs2jWsePpBFohmcG1G
wcBOSMeB+bWo2YkzNGkBq6wcnn/SsYOT0KJXvKE/yAJ+Zzo9E+gK2N+zpKpehhKa
cT3lmPVV6Og3GXXG9zfsU86ZLPVnBwqrzzu2d4Lczy+QtY92aq7wW7NxyAERYnqD
m/h69WVVAmCMu22RGfRj6k7lFm0GyFghrp9/KLa+2kY28P6YKhJ/q6s7ZpZRpVtO
YrldRht0qgCo6UPnz8AJx6RcUj+8qIj0eKycjhaNe1ms7PxJm7ADvoikxUm2YN0Z
9b2KZIr2DFrBz6MJhafxChVfWQvWuQgJvx7jhR+no/eLTP883COgNJ/O7btdhaYr
oxhV53kLpFanYS8imyFhZVpJHXrQRUGEoTSKJkLruCMuT8/YcecvKaVTVXzPeE1E
s2w/Ef+O9SdAXK2o5H3nkZ+cMw2X/1um76K+PzGjU8s9TFsv64e0pSNxXYxDKfrX
9h2zTKEySOOZdKCAeWySB2wMcstgCaBrlyR7jQh+m3mRpFl9zwQnV0vSeKIDdY6J
YqyAK0nV2GwRBRkpqtsUDNx2Uzt3ea0O7gLpe155OuFPUM107b2tSpYU/Ja/DamN
HismHJsM2ucDH15IdEH49s/ds3e7jPl7jrnqP+Y4+WlAjeRDPZD/kxSbxjfGcxyD
YE6M1atolC+aIWQC4hRXh7Lie10KQBTqs7j4uP8OQLBWQC1Qt5JlqFk5dihw86+y
JxDAUygkm5uG06DCUtrMPwuA6XGVb3oJzMcEbHsgYnOBLSj0rQl+hJGD/Qmc6XSO
Trj1LE2+hwgMbrtykdkQXUS1fsXj9qs35OvNPJGyZ7hloB6LMUT0UHohH2v0+kCN
H+8fFJk5+rIYOTC9CGtt63aP8S/8bqotkyG1iPwbyud0BSTUsjBnVXEoHTQ7TMBI
UDtaAHLfMh2lMzm3mpftrt/L/p1EtFv7W2NHcVXOFYhmGhD+B5CHrtTdvZLwrRtS
GmT6z1q6vGsmgJplSjZh4Cbr/UzkWd9gWul+jUUXfMfpKewyWEkiIxJgFZVxpZrv
sDM46zMCgFR52eZ2sanO9+b/ruFbPw5FX4sxc4Cp2aaNRsuxvzzxOhA4YyYvqOyT
TJu3h4osq+HiCtpiWQEz7gzu1Jyros+8UlgIH6Ds2RiDpj7s718gbuw4Ndq1wE03
ERlsGCVuuYTAG3w8yboMQgCzwN16HEHsb9KDHsep4os6oaqO+Os+TmwgLUqhFRql
ghXOE3AvAy+9/B4TJWmpp/YqL+qSAZsVvHLcgEsGOoe3KcztiU2gN56levlSQ4gs
JisLDd+JuzHorl55V9wCw96VghCf48QUpd8HvTByhSGhYoh/2W/jev8eoBq6Srk5
U7tXcOAAXHqZFJMJFGz90JmqOUi2kUb5tQlsLnJbMgghlQXgOgP2tG2s0eWzkuPs
dooqOrlLrWZKDsGD+R0snlbRy88JyNFbRndWhL4mLWkEufHy471INNFWHEU/8oxw
RrYI/pWvJaBqsNluFI2p0TKvCyMbaxk64kyAvIS+Y264Dq5hOEAR+3kOkqpo4Wmt
TG5AU5xW7dmG9ScHJkRKuAaUpX0jO9+wki4B3Q+AiMKjmCvKWkXW5WRWYdo2d/pD
5Op8pOD8p4hKGfgiSn7sBHEIu1XF/z2NrWSK50WPOiL5xyGZDC3V6iA0PkaxMHoJ
U0BZdt/X3ZyGzzpkR63Vf4fEPzbgqHqx6mIQNhvSNQgZurWFv6pmpqN6Z3JEzk3s
kgb+CxIWuhbP9W71klCB2WhY1Pf/GpaDGqcX5A1ylZILCzRAzslmB0vsYuCb5sfk
wyL3TpZ51obcF1ocmed40JZkac2zkQYPZBc5eVrbVYFvuzxwuhe7muvvpVsULgXB
Y5KD5JG9DVLtI+RPq69CB2YuoKeXTKbe5kaM3AcxG0zpx6/Uwnd4ZSk5WiZL8JW/
MV9ryOBhn9UVcYupcCqQIIXOeTkmdAdI+aFcU2U/n+ppLahZ7hZJbDpdfuEApNzy
OzNQX0Qz8Gguo3ZSFM9mZ0G5P6IIhV4ve3YKCjIkEFUC+zz8iPjEJhGfDiBU60mJ
BEXHjwA883bsVPbkvPf0nsCbSNmrexO1wZzUgjwjnDTnzCq7eHyP5pUdIxYYVyEC
iu5pirGbi5zNERL+GvsKWOHmQSkveD2Ke1onvOq6ddXRXlvBBgz4wA7k7sTzfU8f
XYeI28VYSzX8ee/Dm5qvvPkrsaIrinRl7x8RmOZUo9PnU2DfwWfGlA3CynROIEa9
qkWQEgwoLMR+AmVfLDMvE5Pg1HSqYnBow4Mutn+T2JC9AgAP2lgpoFWJMNQanFj+
xBoBFHAM0Ic6TIytYxkpUCPo1abX7d/IntFxeqn3fMoaW38aQBbhSMT71c+/0LUD
Gl+KcT5AeRy3tRngFCNnJLttSHj673SZbHL8t+2EdUPg6HOCZobdwj40j77uXBsL
VZni5qUoA2XwH3/BhC3mbNXIGfApw3zxTDRQ6LKXe6OCXNhGnWfCM8yJu29LsOib
e4UPnsZ18Nw+7INIO4IMUkjQpTpW2wL/heqRAxLpySrM+n2Z6Ol+0WhDMCWZ+Ujz
tEtkiM7CwtnRPwS6753guuVDu3EzHB8mPd3jZxHOyJLV9BF+A/VycFXKutwZ9wyG
4LNLLswVwpABrr2Qg/uwPvHQTPVMo6nGGa7s9r3JHGGRkMPgny5QIcgiQuX4uFf3
F98/Z0jv+OUbtDRSxCR38BonvKhi106EscB2Hcfp5kAKDQ+in4uZ/Znpo4cqMO+d
ySg4BLqYkugODCTn/7uVa6kN82MymDF0eX1v4ZbJ1iOrs5jgI9a/aHRaQMw1UMIK
t49XFEsZ/eG1/iBvgSLPwOA+zGywHy7lTwfFjf1AuhH64jBmzzKwrSU6dFJW/0m7
yuuCLZCPdJd2oz1e09jYUi68aI8Zj3R20KQtG34pjiLmMRY3RooOe8lbGJj1eSvh
OdhezJrbPSYpL8gq56WnlcxlSpCgCsdL7A7m4KECliOKA3PuevoA9JmFu+wAB48L
8Ac8EFw3vPcvuZ+Q9kyylHgCq5KME/I+DZTH1MD/Zl6r24drKWddYSzYt11QCq0O
70GRtjEzrk0bFLPOum9I3GGAUQZBm2T6G3Z/RuM72WeEL8MYUiPM+6bt48DbuP0q
SUBxNruv8J0JY0WcmFRxQliqDvmjNMpZnVF19xCk89fO+834jETkKOGcFa1yHUb0
m90koTP1w915+fXT5V7oBnEAtM4o+Srk66UhG8NNcfNWYBw+/mk3qhxGFfTyN0ST
gcgf/qV2owcsDhLVpuCceNSOXYPstHvrNxTA5nycZ2RPqPt63lx5ZtT1wrUs/Rg8
lpZJk/YfGyjD1XZuQzpwYcCgAORBMlivphTowhowFV3+WPGWDopWcrSQbT1E3hXM
OYt38rJj/L7nOHNLX+5fPhLqxMDzx0mWHHl35TG1vVBBJfdTmDS2aGUIGMdEQs6B
GUm7aObVDWnUo+fw1TUSNCPWZPFYqrmAub+8JTfmnv36Aoah5Pq/WljAru0XxhxR
+e3BmcsO5raMG69P3OcRG01Fxzb7mP68p8rJLBbP23aRm8J894mUkiOWtzaEP/YL
mpuX4+8PbeDbPzUT7FaTVITKoO36SM2QC8bWSNxdOkB6vXzNbpJJ1LjrqC8yOJc6
r2Q/xCSN33VgTrj2pT8/1NYqDWERIDQaK2fF3/uYixYJHcvUAaSrUAJBAt3z8sZM
2zrH39R5ZEHleEOG8GKe+RAB7y1P+B8jR8BRtndvxIOj1nTmBWeutVdiqxixLXRA
/u7RQjC4GCIZJvwiHbCyCk2gKZNynOF5AbUH9wzcd3ZY2G/uvweaZBUwMmMaPvU3
3IrdPeg/7hS/UcEqb6y91D6BtiCZVnz/pm2ji7gBCWHYUHIi9UVxfZ+FNWVUmPQe
1TD3982S58ReHXu8oNno81SvzsjNrGzUlVCY4FAT6aaAwW9HVc6AcQo3z4X/P9ze
M+HZarC1mmOfPUcjh+7AbQ4Vw+amXPY1/xhlLfleJzgGu7qZ9/W2gIhjOKk8iR0i
9pt2A9LFuutAv6pYHokApHk3mFOy0lTiz5C5v7ZM6ZBu/Ny4ExBA1JLRKPToVmOH
6KOQyuUSC32rtdsSVAMcd+sbidZSVnvWKdveg1wSrAxADOadgZpvEOy7SPWqn2xZ
+BVygQPXfs8I6hbHuqKOgV2Lr27c8pOTWypnrhTFdNhJKQpDQ+hYu2QfM6sPf+Iw
iM5gV4HKAzPk8T55J2NV5rGoLrBm89inS9SUAGVicin9GTIuSj9sK+03zYf4psfo
v6hKm2BylndsKL15I+ZKmcmXDrczUi5U6MbE3UyShhNqFLRqhnSTTDAMeNQiUvMR
hU7TRE1YkMTbFcJ6ZUMczKViETf5RO2P2y/olVASsHXLw7iUpcSB/YVja4kaE24f
zwb5adADqwMHvGViJf6o4OgwfjMpw3Gya4L38RofzlOBohNl4sM8dcZDOYIwR5oH
QcKekMb4CaHudJn+kdLGBmfANrNp6s717vUUcViApRMqNH6Hs+khgvRAj1Z3FKSZ
6kWR7M5w5rSn8O/93QlyzBgzp8g2ZTDu1EI8HkgEDCVyiLtx6e5JSk+TTvL7jk3A
ycLMiv0grI70SVxwjbk8AEEJ17CmJ3+YhsM68+DnBh7lbo7yrn8hfnnwVLKPry7T
GeGSQ9wdkUy3xqxoqTVyYd8ZHPKFqlh/BLCdcI/OROpZIRBaTFDLZicfrE+wcaJQ
DOfkfsLzwXpFdKE+Zs4gz4/KJO5u9RfAvehCoEhCv6mmO0jMKp2h6O1MY7ZDSJAl
9ItMpWBEhZ+X3A/eXdqneZAibx0d/Sn9hfnA4aaqol9N8ixWhsBGKMt1LR2SQQZM
KRHmazEYihCzCExyNPYMBem9+C7qPLeFI7kWLJ061yOuCVNQbjd9ZAtScOl0BqR5
jiHBsRZkj8fQCfXYaegqDEdLiyTNR1I6zpbMgL25u1tjqpEs1V5TJv/PC2zUd0Iy
ncyt+JdDOkAqB6/n2niuHysJDNyEtLWp2F58epbBKdSsIk6EC/WG2FnBRRI9Bvsc
3YHPfjIRUAcWWUjhBSqxPt5OOLosV51QmxF2r0XdZRxgLNKa3/6Ksv7KMWCWHEL1
U6WZbFevDZFrnP9JbOzi1pXa/CzjJNraqCWuMLSBXrX39zWMmvQMTf54L7yYE17G
kJ2rDY536AF3ME98CYrPp7RcEOULggwGcZ6rFYSyjrNpEepRHx9HXifTw52QKccN
6eW/HdjpeaEYy5zgTlnpq6mkYs5qF7urLRoc4towUC3d+R1zTJyGREqCNmeqQ15X
rCEL161EpwL2sHIrc3ssp27u5d1+ETGL+UkT04jWl/MQ8FhjKwRj5CC8J9o36BK2
pBesKqZjAe7hrGb2FRnyH5EuN8/WUvlNz8C0OtG8/1ftiyqz9h9XxQGipr6viaIg
sUtEGTtGLQzeRINGyqG615Zj9pjC5BuC9r31qhf/pqtjqv8faVl5RkIHj3KzsfQF
MRe9khOUwGfEWrDKyjBUSiINVB5gsUbCNQDV6jdIUEmqlOycoKu6q9ryU3PZHesY
ClJ7hV6zjM6rHcs9O21CSqkaAtOBGQAfgLtjXnMg2cuhtwP0PE61mTxd8LunMCTi
5cv4hj2FcuZyCqDIhqIq2Qhsfe7POUPTHQdMV6jvbJ+K1v+deO0mgj7RZFjRARQY
bcp1yX3v2ivdL7BKpBNmdiKfZr4/usI1q4n5foAct7tFMnoFStJUSwT6pWUIF+0o
HQlLsIdLeAYSHRUSNyQ+/ga5fjkeSYQGBps/09OlcAc2E78yNJE50YUZu2ZuFTLv
n+/W/19DIi432WrQ2m53Dv3UQXNOib5QxW8894GJHPPvmy3r+wkjAykRfU3AFSpy
3ZjyADfITF44EX9Z88tGUSxjhIyV2iJUBQ19IJKYMOdjg3Pvph74R9fyEXpAut7a
za+zWmKTylXSN0Zh2SBlrAUMClZ7JomBBDrCVd2tcbAIg2Od9V5K64PEVHdcy2uI
X/Cq3acF0Lst5f7PPNmUggWEc8908VhZ4XQS8w0cDt3pQCkBm7hcc+SQqqAsyPMw
dIG0LnfzAy3wLs/R3K0KaCzy6FwKwExcWMjj78AuPFRkZqoyZ4GiOjgz6JeVbuSJ
VGemwGXVGBZMpHPebB7w00WRxRJK6FCdspw/YlBhbe0MBkgHvlHcwhXcjxdDBthn
OVJgd7NADcHFPQpa5jINLFAKYpmcyiWCort1AdbImZytuHjLe2C8pSxujYeHbDuB
me/X7ubiBagfO7zjGR6fbJ7qkRJ9X9kVHdZvEP/M8hakxOBTScKXFrQsDzr5qpH3
vwPpmfFDHVjoXdh3V8MhIdq0WgiFtk09W4c60jzJ/ot9ndf+XzDJ+CXlROvtSfMS
gmbPb0Q40NaiWHk+H7D8jAHxDT2PNLG6URlU4CGvx9sD//Wk1u75p+HJX3T9guvG
7wYM/WNm6NHaFYLa2nRR2Y2rVB2nV1URTo5XDE761/1o6a76YBuoreFWnfFf7nE7
FQ1gtsYf/OWbgtXVS5dy+KI3N+hI3gIjoQgXTYQr56fb3sPhBbw+LWOMoMoCp3fx
UkfTp+t5g9fCE45ABv1FsBo+Oib5wUnC5tH64rI11Tc/NC+WJAw8YBHXJWcB5fHR
zEreIDCyK7odg+94gUOVxJjo4PN23fQVWRg7/dAh1NjWppSOIMk+emAli35I8ubQ
XlkVM+RThBrzEh9Oxod0Qm5dTWYrIrGXYriLfqUyt7GKYJ35YT+EalVzzzAZoOjz
W6msJ53ujA5iO/URd5i35AGbOlWG+R3KvipJZ+81NDyAuxxooKLqUJXRGMcCn77L
anMbA957Rrpusu9G0loKGZo9UZU+XGPN4O+jNJ85hD2tD+nvssY2TES1ghQpCguY
xSczTZ4inbVATtcKOlmEx4LX6Cqb+AVhk3RQxyPM4yX7gVhu9bXBjkus8JCz9JBE
82IaWaee3WG40azmoRiDdn1r+7twZjQN3wp50J1rsPlPbc4zv+K5YXFFU6ukxfV2
iWhJzQV92KYzhxmiYaC2uegBuOtiGTvAK39l9m2Gm/F783WmxUhGFFHDxjMFkyr3
/7LhwHyk29omedrzX1w4vju/EgRSo7TsiOqx2b+XgLTUFlxIq+TPz3oKpKg4Cpxh
Airi6w8DJH84eC+rfeSeQP0/2mNIkoguKzGaN/p7A5w7UVeDjGTJRpmnm4yee6ks
aQaBV8UodHbmluRjfwl2gKlMmtrDur6ssFDa/kRpOcqyvIyb30XV5hiCTRujsdiP
deOPgDtdnyY4n2xSYgK3jIyhe9CtiVFMImlhbj9iosKfEEZdBGFBHG6NLqVNE4js
VjsP2ky8A9inJrX2Fk1Uayd+8bZBuxtt6yvANxeF1FRLfz0BrRce3pWA6ZAKtEej
qeQlqyV7t0mS8KKuwt2+SLw2SaMHi1bvLruiyxv9H63n/6XUmpRpbl+waYaSZuq+
4Umw/+UtoUNIhf+Ek1jEZpacNhEsVF5lCQLJ6nPHBDd/heYrzfJffnbVSjPhJosc
boPzLDLthF17/AxQuPXapdh5pxbLFajNgeTsncrdICU3CtOfzmTTDmOrRegkpcJS
6owKS0ry++7iAVpFt0ebqxbETIV65iyUW1rrS/RKmizusf11nPDLQHDnkguv12TD
hOsYI4617QE2rZziBVmvOcNfhtnxKStgCYEluqxehxF7Acd1qT+fgwgcBcdL312w
GeBJ8e2Vig+ycWx2yBMf7JyWLOrJ845tCUqe1jEWICYC8+eBcaUyJQcr04McZkLR
dCLQ8O/OUXLdxXVJ+2uPgTWSiQENYOMyEn16BiQwT/owrIWxKhxATqIsd5tJoE4G
qzmACQbZXXKM0+FYEuSmAZXzfa8Lm7AHrj/3MvQ8zw156UA50FDQAl0lT5lvvbvi
E2zn3rgP0xWhh0TXdv4Tez9ltqkCKRVVHA78wqXEGgeU+ncKlbE5/D4voiwXlo66
aRyrlTkdtWIsSJqqt+mKIv50jBURmPitBdndAE+vijNMqUtNDoMIBCcUmWBbAcY+
jG2P0W0NwQyuZ5QrD5bBFd+WR+07R9wCiDtWKWiCQSJxbzC3f9Y/TWlA7F5mzKAU
gP5CkG7IQJY5I23zuphiwdWyydGl8N2QTHGTnaDYCamZg4LIM0tFJ+L2CdtDyzE6
lyi+kvNQfKP17wHd6CE/mLnRiPOVMB3LMMTorYZKVoX2CSjkj/T6GpejYer9Xi6p
bEx2B3vf696b7IdA67/Eezfe855Pinhyods+mAbyMW+LV45LVsn4vZS0iZE89Byd
wn4rSWU0OnvPbxpdhWx5WYqqYpVe0fsogOoBSC7V9qb96NMowtKJdD6tyc9vc/3H
/Vb7Ci/Wjget/irJZigYB30PSu78lOeRMAe+8gUwxK9tAksP3pKl0gCOBDpt7MQs
/eUrcsDHZsTxLlluYRkj4gxJygN/Yz+zSk1wyaDhd2grmQWfyOp77MnLuqR1oTAq
8Ibhy42IlnpnSeuCGsJaWNQJtc3hJ4D5m53GDN2kpC6BpKdH4mVxgqRkVZJLYBNx
eW8zQ7TCH8G6ZodyucSAvd6FGNE38kQDstLdJ9Axx22j+W6xcZVD7YmYP/7L7sO2
8xJu57QXd9xeP8OXEjWGucmyFvFS5LD3XG60ZXYAwtF0qtPg9WeSotCt0Oj3/45M
e+LdquUs7eYOe445uBpEm/KETz1Et7j+JHL8ZURnLPGLx7RUrm56vDBL4iGoj+lu
Wh1S4um6380mO1r16FJWWK5bVsjr3VCZ9mzkdJ/jR6z+C/JpE4CoH9zdMjFlrDw7
iXYYaW81Sd32i/OaJy5vOP2NV4yt8laVWjj+Srsn8EVlXC7Y/ZGYFfs8UEzCYMgu
O96MQ65UNiHAgoAylFJIo9KQ17RbAMHtfObOJDfAYoWTq5dcYNbcWbGOtR+hbHHU
YWrCU1QNbxH0/Wor29MRyW/mWXtMiPrCO/lKLx2lQ5aPnR0YWpwgc7ba5ibdYxaX
GbfyYYkEv2ny+UBO6If6s1QwpFMaDIfJDba5VnYdivBnW98+vKrWh3sislKhida7
q8xig168tU4QkD49Fz2Kc9KsEg0TmvxNyiwsFk3kQp5CBo1qK1gHHmv4LuKlc5wa
ioLWj2hMealWKh47t5l8B/iepz3TyVouReP6i3STHopaeOh+Sq8lroTGcia4ZOcg
gr7lvRJv4bB6ShA6swnfTJROgIpwSfCgOuLRVw7Lom39v1CavnQP30L7IXEjzIg2
wNcBMeu8Xs8/VeQboT8FY5Hm9ZkmPXTMPzSeie+PAAxggUvcCFFhPOLpJvoKYnJp
0nZLzDdaJIZXe03MLgd2cXvWfoItu561pFgJyNU1HZp66O65Lb2Tx7LKOqyW5h+Q
yvebr9NMIRGkQQ2qKua47feMXo0QNbpaAG6QDXzR7iyswfVCE4pW61wb6UpvuBYp
PyDbqscMwM2AySCUd5txs7P/P/8gVPcB/zFdzjvyKfJNQMwrOK9PElTliqeLwKiO
lXI5t4luHQjm1hnWhLyehGEX0FKF0sJanWVdjtatEa/mTNb4bSO3sLmTd27SSh7a
Yxm6whXsk9K6ZNRw/DYzp0qprs1US43/5OB9uM0iz/yPExibHdyzsEzo54jqzgso
+VDSgqva1ZEZr/0Pr55w/BK4ZUW0AT0h57fz8aAJnJdFrbnnpNvy8qlRs8OWuFvO
3qP+OldcWPG+ephCoUiDuHhlgqn6lmb1FPCONLUtO5Otj9Hj/j4Y8Ntsh+zzIbjr
+aN+lfVoybPiNz1lWIN5oJo6KkGapLvvNo++cNtv/49io+CWkGPXpiNBHULiWzrx
N8UlLOEgNVfH+7RavwA/6w6tV981Ox/y7qwd6LAyrt7eCY3XWXeFpjFSxhIJOVGr
UXLYRU7II3JHmEF6Eo7lU3EbEjC7SGjMtsSNpnHiaglQncmztoVpXmiqArSbdlL+
ffR0pTRGtj3Ln/naibvcZ+AeXrM2luksJxIbpw7eJbXQ/0+mdZPtZ2TAc9wrF7v9
zsSnfJ9PXb+RkWEwxIL+0EJBOg+sneUy1Dh8wQ3KuTTDPu7ssqcA9QDz9nt9LVje
SaolkCAVxSIm71UK8nOBClMNlUNSCcxybaZHYsET/gWkYBWvEk+ELymg7aHEzJbn
t4cTCSlbFcvHNnM8s0tNOy8xiVnHKIhBbtA40zpHwqksB415Bswnh0mxz27Xf+sd
/FS5Un7c5MHpLVnanU/STO5IQH1yBzNc0WUHxAd7JAi+iVT/ynhZDrTxyrPW7sJq
yZ/s3mMVSOwbGPBvRh0ex/GT5tv7sLLG2kqehBRGvf7af8KA/sdzp325b39fIjki
Jd2JTo1EbNB350bTItua8B9Nl5RaO+PQyvKQJsM582aeuJ4VnAgE+rvfV0QFQKlL
ubxIFEB1/EcQWMy8tZq/H7wCfNMtjiTqdAUMMCKtNIPp2PHj0H+1RDqhtGpc+d3q
mPVMseVi8R4CkGPUUgHlN0kgbHr76njKIeNhH/pu1gUenu7UB+Bv/nLDXVib1nQh
+7YZnm/dBP21eBK7e1SDSc6GbFFVDaZDBwPwsztv6s6614wl/kqD2PwwhprilCMM
t0qx834C9B6uDpT15Q13gY/Tl+7qeNfOBrmR+BPum1UUDKEUtpJcba0CW95a64vf
CaY3zwM/hBRR2TjYPXkFB/KR5Ig/6tmDDtwnYjYrU18vu0uE7cCnGkPKuG/1hLjE
R8QGrd7IzQDl083293ADXSnxOpm7IWYHuDElTwIH4vSJO5FMB1IWk4Z7aPVwU7HD
iEZBN/PeSnZroc7QOZNe3o8A4GUMfQ5+Qu+QSGERf3AR/XRYiaWBmJLfZ7WwI7WY
OnhrSbjslZivbFhH1VQWSR3Hd9cnc5G2wSyiLiNYEM65Fmp28qANpbtKXR8n92SA
7Uj48bisGtICrGGsNVebvYwHFfiYCWv8C4GUoeRdt/48+NG03YA6rbEwAc6YwxVq
yIzOM1ETsdkJtS6nOvsme4msB+n8m+7OErXPu/amjAJFUzir+O5Xuug1hh2EgSqu
l7cqVlqorK51ewU5TL3Oa8O2FOE8FUxelkuaNSY9VT1VVzRKHUKt6R/5vEBOG+c3
SkJYrACAq6bFAfcjMH0NdVvcsp7jo7iNUyCLK3QCHQGr06BEmWHlF/1MdAenBKL1
aA1dMMYKfPVCbJZq1rhbB/cFqLXIdqffm2lrk7CnPuWXnLnetL+tyY1jhwPqbBBW
v2wkvWAFellTJpdeu66F4nI1BmNnGCjP794SahunRUPINGEbT16wa8RiLT1eOQXs
nExUoSkiOquNVr7jEJG4l+tFOSA/BkIh8JHIKmMjSslFIBF84+IhvSFLiwz3R7P1
167vpqHQ686QeAQ+RalP+AqSVqVHz9Xfebfsxfr78C/Q35XasdQ1nS/b+W+r3KrJ
+NP+CyDqIAAZFjlViy7ZkqEIlXsYjZM2FJs9kJVJFMQhizFdSFf/c1aDpbxiZ3x1
8dPPm8MfWixfPp3SPdUnLK9+QzMxSe3MtkbXcgvFZpsFoRKHJc6cbgQ7grL6tQZb
Ogtbuc8GYIiNcP/b9acTONXS8a1JzYXUUW2LJYXYGJ7jNh+ejmL07XhXMM1NAYNQ
x6XZs3L7/tUDA2P5inOQx8SI6jaVcEtRq5BD2pZdzLgO939YGtGqxGrV2HajcUPA
XU8mhhLMao68AxXo9TsiERoQ4+fZgMcjnODjWq6uQdpaRIWNDKM1lGu7iyaQDXTN
32wLrr44byZ0z//GLQN/777SP5oim7sPd7NglkRVZ2QlcRN1ktO9ibBZLknhUD4+
jjV1+KyY9who8yu+HxH5wRl8YMLh1UnnR1roV8lBI+HjeSiQhBRnqFUCnxtqAdnk
pyP2eIdQac50Ziyn47jJF2ahcsWJGu94eOa4td1JvTit6kiCV4Fa25jdKs7u0Ahx
cr51OBoeI1MSH1ZSzq7pN6X/jNbP/FbAj4vkEwMhaPQfcU00wQgOqXlAmPs4yv+N
xck54Py3D4igPcUK0aGLKNCrWssc5Wudo3nSpv7rZwdeCSTvdbmWOFjq0nJS+yah
yDd7tl+ZzVU65kjcheOsJRBC3gBxFw6qYhh10wq5d2Hr5gjif3GcmEah7vm87dzm
SVABpq6YqIQL0V7RlXr/SH4MqYi/VvqNNe7tspjGdyRLU46B/a4Brdllp2rnNqnu
hn6MON5p1fZ/RxSByftXIQb96F+ge5gxOxmdoskEZMl9olnygTRI4BXqEiAZSUZf
0jyjeoPypnCuY6serHNkAwv2B79imtVBZo6z1mhEHAgIkkC0oLNnOr8BguYRdvWp
xcphxvk9qY8UGX6wSv+fsZDZgyOXKNO3bpI8/qdC14iy15d943y1ZLKzM/F4OZeW
kQMri+lOLCGsR7/Qe/dEMuSkE4ZyRxiG5gUgXdbV617yRIRJ6heH0PjNdwh8hd2t
1kjCtxzcMyD/BfxF3XqKITagHfsaFYw3yAQ3AbWOWBFwZSzzqGKCedlNHFKm/j2a
sGCSQvoN2KZieWgt19Qca/ahQQDOZ0CvLjngzLXmvI44fmmucf+NOYYsX0bxvapc
Lhy42l5VnYlIs5QmVmosHsD+78uBc+AKa4okAxb7ozL5N5bW0tSqKNU9uG8/ZBl+
tUJ9wqAp/Hc9GdR17lr05H1ZYCRgN89jeCycHsP8lT3RrgKr3XkFP0SxsCdg/hbt
0E+Txlseauxj/kYKOxT25PcFYU9ESkuZZIj4nHA1Fjc83NOxMw+HTDfVRIGfQxVQ
4RDZbF7fVvgnBwpbgiNFF2yv0uwj6QVCxPN1svIiFlknV86//pNjneVmrM0FggUX
SoJ1+y7OJqt7FPjVX59ea3nGkkf7rFK+DzFIYGYNGPqRwulak0qSHat7oAIBu+rJ
u2jmuv6y2td6fBnZPXI1S096yiYy5I3qkfP2VxZRkELVeKth2Kh8Fn6GfAB40wN1
uELY4Pi9DnQNn2hrdYB7t9puCIKkj5jLCgSG5vzoemZ3Ik9GlN023lLQ5uFWqE+P
+f6N5fKbyO0u49fpglL3QORq2Un7xBLddyqmS6c0brMMFvC7lOoklqRnFkSSrCo/
MG7AOVC8YSv4aJZ11ZF/ZoqCVtmWF48urvy2vWBazf9/fYzRpRTBk3PKYhCnlA4w
SRZF98oeDY1cE2R5JjDli9r+TW2RgGWJG8++ekifZXm1uz/ahm5NAf+8dvFkFA+S
tqHSni8+c5g9UgAZRqZvktBYXd8fCN9QZgnXCiKS19vxSWlFunXBtd85+DdDb3Hi
N0NILOLSwd03NbhIWTy2aE2o22uwcUtislF36z0p2QyPAJSRZTUPhdDhW3Bct+n1
VXFWb1Kx1QNbx3PgatSDMrKn0lX7PdTTu1a+RjBv60k/mhFRYs35uRpiaUAOZgMZ
0hWOsvA3C/piO/sQQPIKZnPqmPBWIxnklXtn40GezUZs2yCjvFX7++HWCWntkz/C
vMT4ObbG6bCk7QdSdVk/NRWMN11Ole6XKu7Etz0BH6tREer7TNBeQ0h9O26rJTBG
f+nYuxVfqgYkNtNQ8QhjrOn+/79CXugV1usl50tjl3dvFiwtQtJQtGaKq7YyPXsY
mHaSlsnDeghIzPGkpCJUIzZ3jlc9ZCNIzPp+cc2eUruX3ClzLWJdQY3X84UoZpp3
KWowkmX8VuiwYguAtYEIOcKnl1vhkY8S3kz/JCQ4MREcawrwGbMPPfpK/eT5n1mB
WuPkueJa67D7W+DPpsr+vCi8v+OV0dc7zQ7O9C+fffqSSWrxVNs5DMhZ5d1LY0Tk
cZ0EYqfrXuIykQGcvzP027YJXRuI2XLQvpcxPDx5iNnTRLHyDrOn29jRrFlFM8sr
XVuUBSLV2asFsBTS37UJfOpJfZz6htrHoN1ecaze2IHywDLhkk49UbJeZpW5eHik
f0PLjJ3aWy8EG7VJkQ7NOxQ2MuYUkC06oD7kBDupXWvOy3lgJV52fZUjctnBqjhs
rB2HSZjpgHzGLpokIetCBqG9EPM/QiL60c8eY/LgndYtrtVOvfuVDDSKNz0OV8pi
1G+Iq+ETaM+tXnCGKev/d2hVnMcppiLrFq10FxrWaOCyDp5KKHDZHEzOcozzUJTL
277I2OSGuAfnXeK57jWV3znLQ6mJR5T59spesOxhMY5O61/5CfNl/biHtLRPJTIR
4CBI6kRnjyfMJJgZszF+VoctRK0Gu1xx1+2Xle7ClCe2A0NJiX9TdXOsHBzHpoih
OKTzO9FoZSZzDbR8ZqC/SPysahMdgp3zdxZGsmogN40VB11YMotZanvo4KncEv4u
dzpCEF4UBPXH1T2t0Q22mUmamNO9WaNLdOFCE3lRhgiC2Z2p3rWq/+RHkgH8pKvk
FsyzupyPF0GaXPkpct4LMrqLYUxj21sJKmuXD7QQNhH6Wvglb84P0gbV/x5MUzD9
18JCLWeEWiXb8eRWqbgl5QdVht0HkOvEx52juwcPu8IFqSFlIkhNDPInvGxIYpeN
wY81LIt9DDae5XRq0LGz6Y4ddiY0dGRauw98nH3IsUzY6mvZrw/ztZTaIG40WJ1s
OjDD2nqYQ2NeXptz1um7KGQ+an7BIxwvIFv/9ktdm+eKyUHWNcxqHxSRErzEgRyK
nbssmcd5kC1jBOOKeDI5iTJUEtbn1jcnDjhIIciIqfXLpejnunapR0GG4YYwiS82
jKgxPL322crB01L1bWTHuknui0wyqdhWyyuWV1x1cIzgvoRL3ckcTgdltU/gI8qV
ErmfZNRD7JQf3MOpqDoQHSe1jQAOFIZF7Y/GxztQpf251rGrbbEW8aZh+oouF5RN
o9pqeK6lMp0VzeN++leFhNkCgpgsUobbf1/BsjuIFO3m7Ish/FvNeO+tvhxqTF/l
Ld/80bxhH7ETPN2lTqJ6Sk9Nsyqi1yEJmuA8oyYyYXptnsAptZjEYA0Cv455ED0z
v/0jHUtCgCIzYoOly1te3NoWWmW/+od8rST/ZnPJ92ZHjKlt1iw5yCXDfgA+TW/I
UUGkxzYyUF0L+922wt8cXqW+7dzZ3fxrOjWbmXHCVfshlI2GY8IbHqSulX0qfaIH
p4CjuATejiVT0gHUcGVFuvM/sY8ecs9bOOloUeUTcBaxaGJesncwikUck5scdOpJ
Is69vqIjkZzTCrA55kO/eVdqj57BerR81z7iMhNWWofpVui9u9WnuTdDYrgVrRGH
E76ZplraDzQwzUQMvvUkuEhq53iLKqnENWRF9q0DPeoa1igq4eeIZURyeV2qgezy
AE4HgUJvmnwoS+sPihKI8zFRwZRi8MVuiWFjH5BGqckm5cxO97AGMt5WJguLmBPb
2qpazGCYxpYLELQU8fJy+6OdAYEyoAhjr1UzDXvX74dUCAW6TB00rsi3QsmItGGe
SOh+bkqOc9L444fHx+STaqH/pMQD5FjJOhKk3C08Z4D5sS4YUWTR5WPWhZJ18UU/
jRfhB/MDA2izZW9073/Ww1nJ66LdGI6h+cxcdcdxuSP849Ao7j67eQVLgmThe+R2
Hs8MGkLi1qw7bfe/12Mv2k9+eG05h/qLjev8tYUvi7hLyhiw6Ei4YDI2g/FrV90h
bDsyOmOGthaq9o7J2zAUJW7a1tvOj1n+dr1+R7QpmQpwInN2qAIHrfCpuI+Ebqa5
QqoNSHug9QAbMe5/8NdHnbc2RpRCoSiqVNb4/Lq5hGzWhzd+1YJ7bwdEScB9+LMq
RVpz/b2XOTWP26FxtkFMMVW5LiDS5eW8osJOWO7PF06asdQPy1ConUT72gJ9Ac5V
UkXcprPGpncZVx87MBpBpx42YCXHcAn8NA0hVgQmUJrqlh1Sl9hdMVLgduhV0G9Q
jlWrDmnL0CnmDZY8nPAZaxvkSv8VG+ROQqDgUb5xXARFdkFMGli5qutSRHgowAug
im2wzYZXIM3oirLMCY+ZRAdNpsRV/SgQJMyR7uZ+aIA5yBGJEJP5Uy7l1cvT89fw
iwdD6E+7A6gaPyt3qcpNjnd0y1u/LldShD1Q03zhINdxyBkNtOOhwTUwJYnEGTAa
2fyXrNzGKyEtvbCEbeRmMQdNDpL/OmuVJu/5AjaIrKRJpIY0KxoBsWvpffNLthvp
x9N2fWQNjjBFiQK9zwRCN5sSoin1RusGMQ51pr4X+J3EZab4DUN+Q0YdNI5OUIbH
61lsQwG9dQJr9fkjBG7tii0iuEGgjNEMq8F2SMonPvHQ695FXKWhTS/JgeT49Hsu
zEwFp2pFxYEzzU4BtwZx8Y2vFZoCpvw5gy8yxf01h1ptU3wJ7kpRh7S/+L79QvJA
8QS/IBgKOk+2i/LLoVd/1AMfpkhZCl86zcS7o+zAgEOmyDvic9ZcB5phWgSk34VY
K89zxK/0lxOImYP2bFsQZ4IoTXJ7lG5p5u11D1GAYB9Jjic+XldJEl/KW6YvTzRg
blfENe+vgSjMkBK/ObyruoTSz6LJEKTtdCXIH8RU/FUFLkr45XFEI/AKcLoxVCuF
7QCgK/7NG9QBAhlKypjikLBdzmJ7Aj4EppIRu90M+c4gWX7mIsDH1rY3jf6Zvjjf
PqQmIZmXTX2gRmb+FO9MzY2DXVL1XXcrgfb3lqAsGVulSPZHiL42eJL1CrlZAWSr
/134Y3tdhacSxNRQXGKO93+aH763pfmEyBPaw52Lw1UzbUtj0iztil6Q8hkfVoj/
mSsW7Ote+Gtsrt0/LIu3jzRBmgi1bb4k6L7R+nVl+c9WwqmPA8TX8k0zMRZJnqVB
xxxuiHFsD82vhPxPHUCyjS+WQDMIwBllS0oBCOQHYp7Rw1CXaXSinsCYZjsF+qdP
YrPb9EUq+GLz3vtBGTTUOY9rRgLlhvjv6qf+yQCLyfwzinE1s101yPqXux6gh9+u
wxjy1qeiyi+3O7XmDNDyibCU1utWfSytJXiWQFTuh/WTZC42qDyqqD8yWv8NKT8w
1c8NFvLEaaKznwATtq8a1LvJKVMyC2dDJUi4mWlsywkPfJSBYO+rvKUKy+yVarSQ
9gnwBzff49EK8V1gTGAUSlJUw2rydxkfy2pzx/Vb6ZkYndnzEnbdyt0v5Zi6aQWi
g9XUPZD4jc5Ya8kbHGMmR3BA3jln6lM+zqXH0TcLkEFxqaBTskVNQj5NoUA2swuu
ONacfTC3urYUVab6BWjgQ4aaNIv+dZ50sPA8FzA/5MSYJfoky7JsmDyuix6qAQ2P
qNu68kF5pjj2Z3uiolcFqtkxixHpLCXx5YK4PpuSJGQvR8wd7G/tzKxuZhsqsugM
3wLWxXTPFrcNN3nEGE9t5mlNR4Iaolqiik3mIGsVu/ssh8cvVZbR4Yty9RCxCRcm
5QTQnETDpu/QdYI6iHzzE9tJ6c8IHShigFsSMy/2lUenY74t/XNfn3FKK4TT7Lv2
yap/40EQCYOM4unb0ulQTJMTJ2jChWDP3LB2v5vBGg8Dab89qSvYAqTgqka5Dg4p
W9oQWDYOopX/NCyv9Q/9GpM62nAHDhCa2B3TRlbqnI455ZgAJT5cw74oe0Yf6B57
2yKtnZRyCviiwFNc/lhe6RjW/qdPTGil1TvKVSkWikZtxpcORbKGA5N79bmAREky
w0izUGPX2Ioh6usi9LkuaaWZDxXoGuM21l6t05Cf/sgn+nVaiQw6H8c5lJLS5cHB
gxe9YfUIVr+waWlNrRuFECaqAQFJjUiuo5opiKmMMmaqJtHOk/ND54cvOluGhewg
blOaptartc05spQdgBiYwBKhkLBO8a0gXNJWioBaklCbdmq5ivXpqyIQkEa/g31e
wdur9aMyNTszGoSfO4LgZemrqYJCaF8n2hVL3JQcPYV+C948Tt7D3IlivFzOqsZp
ul7IwwJmSzQlUh9lIPMsODDYMkmA5rGjmUQAemw7t0pcTuQzkQATfogkMHQgqAYx
YuFMZgfxKPJTXo0ibXr1tH8dLiwUiBbbOY5sx6Qs7i+7prcg/hno1eRY0v5LDhMl
NgGSdBBCLrqz3lkdyBMVRkbjON+SHTKayIN6K6WpPWyLSj1FgJEoR+oRUH4MEKFJ
2yMky1A1TT8U0oJ6hrXkdWXgm1K5kU+oS60PWnM4ZoTFX9A1wmpUqoUsgBRm1cnE
Y5n2dWGOZP14Fiit1eCWIZ8xVxD93rZhUv2vJ9hFlzN8gXcNrUzrPSROcR1h0RaX
wQLte5Y8icYvN6If4iRkuUobBKQ/NzggzgV5f7sxuSLTtcKbc++ptJtldFZFwkKF
aBW2fwIEqZX6iUnApt9E34o6L6chVcy9GPw63gQ05efaw+GOmqsClwnqGblT7kgK
JeWpiVFHW0AeU7dkkD93lBiTbVqwP3+LwZ3CKBEzAyJZl7ki+r/ylMx/s2JZ/RIn
taLpK+v4jj8VwHHpypumIVpbAswjfxf5N56iBU2QF/ZoigAr6705lzFRsKBR4JlE
TRil2KxHPlHIoO8AnwANYQgVGZcLNvPFPfthdGyw8kPBtKPrAXsj8FsQES8CNbJR
xZjpWA/NozocZleEglD0BcEyZbYd1I/sEMpKKPUPbvQvtT7jGdKuBcGvPdxPQLLC
vUC7bcs3D6x8ryq6SEXbxylw8QNHfz7rzBhrFDuSTTjd/p8PQCh4dHeK9lxdzGNY
RACcV+kznoYQDFcljG6kL9U2QTom7bc4ZUiTfedG1/Rbfjy4DszXpq1uDcyNHUNU
ULbwxRaDUmFJHI5Mjd0HxysNRUN7aSSMTlFYSTXLc9KHfM5FJ3x2sbsDpfBhuwfK
s3vlZy6Mb5euBmqk/zJSdnjalHVfQkmDTVVuy5/v9rROPHcYpUMbjc94+bStopvE
iEZaj7BYm+ab5MXk1LHzrYZvCH3soIkVrlxXqrtM2pz2jlbrY5mmfqhG918+zXso
1mNiXOYbTLHW/v6eEmTBBg/YTxwULDArpuvARv0FsT4THiKGGuWYs3vq6Fodim+M
GcIcOCs7+K6kYu1qCWN1p5YATb6gOfb9oLzuwqhQrX2lA8bcyh46x6Mupr9bHI2v
WH584OTLwrQp9ITPJmytQ7qMh5LBjLph3TRTjUvq9tyPmJ/mM7xXPECKn+U1irlT
67Afpdi2y0yqtA1JY7h+HWtgQ90d7QujzkfNs0UyZ0vPHhyUttETxiEOi7kfvAeI
2i0brHnLArthlbkOWip0kRldDRxDrjXYhH+swW+QfPWftKdEcz4mNPia4xbiVEy1
ybITtGYriGGlJowSC8BbNNYFDkDmDfkB5Nf6smLpKaPM+0GgsrXFJyeQdODVVWKg
9SzKeec06scMg8gnT7qtCcE09MxmyRA78udvNq0RNZTkMme3lY3/aN+7p+qIPJoD
Uke0h0GWcQUlKzu0I/We0JkCh5Vqnum/rfHcJlXnIGc7ypAU+gnY9CV17gX0tNJ0
khFV30TSv/z5UyNGUrE4rVa/3x2cC3I6gXSpChQ4KZfIlgxQdpqgLqNRhv11OH/7
Ov4enQmD0MeGeCJqnbWVyBknKWJf1Hl6PVhHHbhCs1jZmWvy2k5vHtXHZLDj/1Sz
qdViyGsOzqkkw1opz2XQTKfXW/PUmt5h8K39NlwIbdkj2h57qLYlKJPBlXGHQdym
WFSYFLn5/Fen83/jKwQPOrsCofIu3mEMQFwnOT9wkAvpo/re6xLJlcd4q1q9Ntko
wRJXWMtbPxLjWLhg750rNqsBkVqi28Szpz7RgpI/h+R8Qe5BflGVlHoW05wkO3oX
opzw/36jjHxanWnDdqBXGEOCBj+gcDH9M7p1KagWaLGmB9IY2DnUCbykC8sKAAmn
P88Vm9nvvTN5W2/4LkGHBXlqzGWLsBG3nx78/NGJ0Nkd2K2iPLmU1rQLig20+CvF
LdbI5gNF8Ygv55eRG5xfHt8NXNKOyKDxKXFiS+kIJfKEFLI43dHNJPe2oubP9V+Y
BCDH1H/1VOZ6+fuMBMgpQsOjrereStmDBFJccNmA3qd8a3HxYjd6QWSNcStKcYTd
11Y4NhYgLlmRAdVLxOiNN0q28RcW0PfiljANQGpv9UGojCUO+L+Wrr8ieGU7sTkh
BDIRR5w301tUTDrY30N+0vahO9LvULsscdnIjl0dLdb7ZitgZycI1QDzWdWVEmyl
C8s3Iv97bliHDGjf9zfxGDCObRwvG18pLSu3XNyOQkRG1mqmmxXc5Uo+GUpXTrv0
Kuu63p67JGoYIHMJp4UkLGDYnuzgSMcPcr5uhAlTuJlWdb1zh6ru8pfG+c5IWsCW
5IWT3n1O4E1BDggWvYcilK6No0PDO4FrE3oqRCwAOIB8Xo8RpzBpqBUTSpvE2mtE
Ii4N0h4EcaS1tuyxKrlM/DiIBCrD+6US0HJGeX8HJHek4x37n8NdDECBCeoPOK61
t5QjxU54filf5/syAZr/LD7rPDsZsdA9Z+GA1MxXfNS/WVMU3YipZHTYYl2il01Q
Gi4pta30iWnJbYPpuK97K2sLAT6XOg0UYW/tGySw6bsF2bDvnaeM38LY/5dUHh9X
TOWuAVxrAHH+PEloEOIPaFIIFbH7IrePLlyEcVKlMHH3szoux206IpzoF6gpGWlB
0APb/tSqcVAvXMjbVjprA4LKsVujX5C+a1SZ0AYFbYAtOs3GTxNzE+t3PjkfJ+nK
argFaS5u4fno29M+D7ayWjeilYWRpWOeI3DqtZD9PgU9UoLCOIZdIHPvB5QV/a4B
lLEn6rkhh+QCCA2os7hOTDSVoCQB0tJcUtSWeNi8h6e7RK0VvPMSx/F9aXxtxuyv
vz+D3QV7xboQcQwH7DiAGdVZ32LHujk+3xlntwvlkGgkxhRQJYPEGo35QSy3PRmX
ZdSavQhwUitaC3Ns+dtL/nT3H/UZ+xtQXVQsmIvZHUh38VEC9mOyXGv0I8sh1kwE
BOPU3cvLA3a0DANolUoTFJ9GMeUCobXbRehH7LxOmfYFxlkVHUGOnfYwUAyDttqk
8ujyfgpa9Zzc5ZUTPtWm5ByLKN09dYAt3DwrEdgtCtZjsCk8v29ewZneWOsw2WO2
6r44ib0BC9RK/JANABc2tUmMzUB9m/2Ayv1avav1eYxjYykm/e3eIJhbL/lE++46
56LE171+l66qwSizm8k94Keix9kMOu/bfqlgAgeLt1SuMrvRGmyrezmGNEpYM4Us
EUVy000JqIQ/vfYtNxUdn7EqYxbAqYlm6Ko2zL4tigMLbMspf/nOT4+IVXTe3S9L
MqW4S8K9SmKwA6DP8/KkJzvL+wgwe6p67r70k43mL+X61xZYmLEhkmNZwgzw3cQ3
M2+VUqS/7y+qy2mDB2lX/0GUd/D2x3YyrSMFYa2+11QiE59hk73WgBqLfzgW9+QL
GQTyomyGAXAsiJzbkezKv3qt/zy8PJe9CLGoBzg9sHDuEKSzpDZEVJYaODRfdCVy
wsRabXQ+g4OMQrY+/CrFft8k7DeMr+bchSbfHrAF9DxtukI0ZgQToKwhZhRufHua
q5TZSiMqDoPJ2MUh04WxOOucucfz17mNjY3d1F4kIdhyxSrFZnsP2WCLdRYvyg/3
t7XRMUSqvgvfM7Wnj2ifuudn6ccHg6GlKqCeb8hrSixZcqSMdGuqsGZ8Iu44mqF+
W6gETYqMkygmWqul9PBIi1T9t3w3+ebC/1AplP9winxIJ9HUUbAnDvoXRhKO8zls
gokxrR1CIFCzdWSOoUqqo6lyT3k6N7IbRwcLrpbbyMy3kcenUpfQNEuhAAZAfxfY
44ZWo5xrvUSUGvJs5ywTRHg+UgWYuoF9vHSPv83cy5Nr1EGdJZ9X8hRxfoFLcmSE
JRrVbx02gpQOD/+BVxBS9wuOhtM5jXCxmDNgbXNv8ZjNzG+nQpNu4c+wPO7b/KXv
o2pM20qAfZWOEKEx98K2X1dswTzacF449JmhI667CP1I5Trydf4WwMaEyUzFftC2
zDAaE3lSpIVrgZgFYX67zoAVvCgAdZA7PdLWAfqGTPyODsVJDqZSbHNMxAW6JB44
85PU8xzbiRSn0082wjuCO8yENEmYV7KYKRtnNvDH8aQcecdRekd6Gk4Y9isQyAUs
KoFI4qhRU87wS9LrRY/RzT0iTRVCZlRh3pjYDS1cJc/bLjbbiwPPslBHGZJsM6xt
U/3nAW7FweRsIVycH12kJbaBYz7E06g3tAmZtu2SoSFqD2sGOCagkoOD4WPwp5ir
MfnsXkRv7XT82l03sPam/UCn7rqKpegcdAfUWCQj8w/B7YZdXExd62f7Ln2YZBOX
g3O4xnS2QI2JCFnYQKlY81NdvRlg3niD3cfQuvQNWIL/9ea7jBquFAaBUIse9YpO
8nrkCpiXp139Ug7XA9VkXtFDzjtFHwg+Dx7WUu/B4Yw+dlwu/QTI0ehIdT6h0IBJ
UbzQ965ixq3Cvcb/vEDDtcC7MqzpEfoVX9aZNjrvqjawOn7vTdzR4nakuHpvXXXZ
K06a/yL4tvzyUO41bDPtIjvCSVLLN8L4Z/jOC6xvB1HvNJbF/+dR1C1QTnHy91sc
OaBpei8GPSmc3/oWfCwpJ7syQxyClCTv0o96I0r84yqrR2oQ88B1uepPXs4PkiSl
AT90swPd1klRxQsmEgc4skj/GIRkv3PJPSovKDWC5SScRBbX8HGLOqD1up+QvDSt
K/bXuGxMTqWvXgMf9jtc+fMeKORx9/jIAxTX4osonqdcvrGVXtow2A2B8zEEd+LL
9PbONA/1MKzNcNqZyo1vr0yU4be0IQf7FDmowLkRrYEjDnRcVppI8bKgkbgGpC+O
6+OF9wQLLxqpRXIBHW1bpGWfOY7BIsMzfhzH1/b1WKggM7uSXPjOVO+UMv8LN95w
1Kn0OgacwMuE09nMicYgdhc2EA1ODDLxtvZwQ+hQJ9AfBDxvxs2I6LR6yBMYUQrT
yYf35YaeIshiziDU6YwC6DxLoD7YNq0ugSazYhMYwCsOvk24H4YMpO/v4yHbuwCx
K5Gwbg917NXs0WB8maSis4G9qJwATconDJcgdlWIZINc09ILG+DI+nS6ZouwMkET
zvb/Vel6B3s6rUiTF4i34KRCgLtrN2cxd8EtKAy8FDsnIZPm+i2dNwikJpyhZZRr
t4GI/OF5c/reM19dQs8en7wPQzmz0O2lyytXTAjrnkyQvL6wCBtvVVX663XmWBBS
4aMgWM4gnnUEZlWrtc6NhAYMn9UJtwYcwA5/KkvhmUXrZTh5+qdtNVQTlb67YAJW
/UxC8evJoYWuy2+6laATe+KlSjOqtJa/A0FSy2XGY29vYhd1qRI9EkBvHw6vkEXK
eCtUo+QtHS1vtFDJzO39Ed6hX85wXzfgor+KbFzLg70zRikniXiyP4reG6QfOlzz
1oj6ilFjtPGP4roys8Hk54zbRRfcj7z4oSqiCNY+RI5IVgrx2YAsgBBMHy2/hpPs
amb5CyGnjfj0oqeeS+tEQ+VJHPswjJL33nPcB8l7VXbuhnu1c9RzyGfAvwj5rEja
q0Gb9+3xhW8MiupoX9PSzcNx6zQ7l0ifyrP/9ZUzs3VUIa51eVh8vw5Xyv8vYR/e
wQlw9xv35weTX7qP8j1w4m9sxklpoUHqvRg/BqzuUEdBOvoEskQ/J8Mj/lXFFXqW
Az1rUjD3OxFpyNFLTsGEcr3zeh18idpG0/28INBccurAtxW2JQ+ZcpiOPvAliIGU
O5mxHETxIbkWP6n4tPDJ7eRuE8AMS0eHGHjZqv1OOdAfSfSWni/Pw26z7quFKGSL
rarrKAAH/V/Y3VJYrOU9AO5i6Du7OcsA7QyS2jDZh/TuSdFcoAFds+pE1ZDlU7Rc
UrIkNUYgri3n0nDrO2OPwshbImvKeYzHVVUGLSSqENPxCOI/X2DYVbpn1xB+oPxw
UGOAItzr17KGm6EmW63bLbxeqDbjFcZpKfuHpxXNwJ09d/JsKPm9eUWOCrYZZhBP
wodSMszodiVRbZ/OQ7W+MAOCPSMuVmXcF8DkAH86C0R/3Rntg879/UTwZ/wuLhEu
uvRmjJWQRN6BZxJPk3gVtie2Hg5yCx4OK3uswJUvtE2MCket3GnaP6PZ6QGwXvmN
ixu3vxLRKvbAMmFFEl4PziHE2dCnQALmbIU6H57JnHHKhrjZehnoTP9lS4BgDGfQ
DT2ESAaCu0YHtDwXo7hDgSrjOtlGPegtKeab5TsinqD8YSW+ocO3ZAnzIAIRVP87
SpytxiyyGenC5jhXg02+aZeE94VAW999T5U85vv3JxuGI2DseL+x/hyXRaEwpYUM
IGYsVg+vHaiNYPscMi6fPt49cQYu3LBksPdZoSfe+Z4DOM6e9Kq/lCmalTPgsL8H
lHq9HIIE8/+X1UITbvmf4uOXaBTnVpdqsk/T3s4VMPY4+tbVUJgTpAIE/HQjMbMM
S/lDIS1Jn1lZSD0VpMTlxL1XPNy82ddjLJ+KdwF6KTNYYitu7P9bHJ5w4a/6MUBH
E5ubdSerx6szyx4cMF28o9llXiIkMEC8BTmHa1+6D4g30R2zEGbLYKdoBH1TeDSP
DHRyaG17LjBdG5c340XhXFKDML6+yCTSNydw3NJ47yY8huZKwpKqMJfMvJgHNgJe
va5aEb1116uGUnSWvjI/aYc09DfTBSACgbqKEAkPbZtBtxnW1SfnOiJN+uEcbHWd
SUgdkOq5PBWQYbOJqx8Cog5U+49wxf9y5LNeoUh0O7wCPjNFm2b7Ulp0S76YEP6N
j145ukMlhmASW1TbqP70/914r4lc6vOf+dCaE8GcBQpu4M4S0xF/ZIjrekk8dFxA
7qzVthJn1h6t2ilkRVyw0EPMJuxtbBHmJlfqnNJPxkdOP9Fuo8LEiG9wkgcFrhDP
0AhbHY6Hxi5SZbV8qKWKf2bEeUNZ6C+6x7bg9dJK8yWpgFWuqkdUJGoQJ7PL5MGh
UTeGfLFxTGsHMnR4guI3KvOb7D/5b/16eqlX2pCCOxa3jvdA+EVHwSWQCQad4zWA
TaYXLjdMZ0XRqRhlNmPqSVwV4nkHovLjipc8R7swk62/iEnmHjKMAB+MgUZ5aKsA
aIPGTdyCDXzz/LqlMdhAE25iEeVbCw4+dNkYrH0y+evZ4Tt4v2CIRXMS5v26+Wpc
BG1xiqFAOf9L/GMggTV/Ea62wFRdcMRDH8zSgG3ETrG6siu7LkvK21g9PRiPEn77
gyQheRKy0UF+MMg0MGsxCJOJcD6iWj+gRq+MeHJoDE1M6AvhjhGCVLtC8Et03tAL
nunA11c1z2CnHXUldpp4TKnFTLJjZTsyDebNl8poa94M4g+gowVTFBg3lOqTeHTA
dIhNIgPs8SX+6gdUFYCNjeMdYgnPijCVgn+rk33DfsEPaCLczEHE2z+A0854yfmX
MmZdIhi43pL4nX6R66gcaAn+WI+EFOjjMg3F2WKmZarlbRBTPLbrcubCpSz2U7Aq
+h1+0Hg3d3Uk3h8t0KsGZ1H5EyVXlWmbrRDckCUDIwtBam6NYkGB0UcJd5BO0QOU
xTdJP3Puxp4pkrfkq/ag8hW+7omKxIQFJWiAXO/jos2fGnZ53RqOp3osAyNIne4F
W7slSRyfGLuixrL/sfTRaIc3ZnLvEZxvp4J/wXTk2enTP2DY+E8JFw741WvOLJF8
QnpW1IhuX2WLW1t4pjwvgy9hMAvC/hDHT81hx+b6xCrI7odtlolLLD16RcsgIiEY
Kj3WXB1uMhqO86wlXtHPpuZJs9TXzfd69pa/XcX4PcBxI8NQMh9zeQHBVOrzqv3c
feFzcZ2PAnweCz3D6UUeAjxxapm7bYYpix7ywNfaBV7VNJ5RmlAqBP5oQZ0EBKiB
AWSRMiQvLsqwEu1UPG2/iw2IgD1TddT0qFxGeoYRQ6zZ/OsuETiZ5GaJtJhHZ81T
Jprhr8niT3jZgBHkaNWeZ4IjhgNLrL6HM1+eP2bvrwjJwemj5Cv3BRDqPB24H/D/
CRyp1qfXmbJZ6IQvKTAqqrvpIWSX9eUAvJAr0FpUx6Vs6E6FccgFu+7RyXQOWm02
XpRq3/en9YHMwCfyos93UqZdm6dtcBAPdJ3gVuyb8ihxBU8bwDsw+dmOOygJWEJ/
FDnuHbaZLYRoe4yDhF2gtDdDZ/bGZ+gH2c5gACpErYd65b6ek7RJmXUuUMgdgJ8H
TK5dwr3vfgZqthvQ/nkyCk2lqUKtgJBf7ZOCj4NCyv8JCNn4WBPcwYvAZ3DiFFHQ
+1dyoL+4d9xPtzY88xyuCyYkzBv8JK7iy6PV7ZFBMjmNLYDNFP/Xa5RhpoX0i+jf
VHyB0tfRodzXYdHdkZ0K9G7OHoezNuT7pbqYR6gsJEyTEcFMiNNKOfaYIeJ1D3CK
OpDW/jm34brMIGHy2u6A9BQrLQRXX8HxID5TghSgO31mDAUeha1SSa8iuE0Ttx1J
GfWsEEsAPOg03za8pG2gfdrHaBfP17tk9/6LujI2NMCcht9DK9H6RMF+x+uahDk8
bU2LuNDIcKJKUfoJooOAnF4uAQiqIgjVytNyn2fa0MVslu9ugE0ppXyGJhJPducr
a17Nn3UQpQrSeOeTAeP6gowsQItRsqV7uxIFd/NLm8zi0HpQSr/xMX9iJdcnClVy
S3I8xm37AkKJYwLG2agdFMkFOQQ832nvHvLeTp4cil7rtvI2rhcDlJJA+7bPlh2K
X74F5cKJsBk4TvdibAUHWjD4HFu5mLq72ikyCP9CwxZ1IH7VA7H8III8O+N00vp7
H1WQBp68UByBLR4/XFu8cXNRn+9pkUfvJnJFSPXyzf/mWlIaFn7Nx0S6PBow6yYf
nbWwPxgZjZa/JefnKMINWRYvZvpX9p5cJJJ66st60yzu/2Txtv/GzEb1idz+i7yd
cgvlzuXNT9PEUNbVvTizrwM8rh9RSzPccfLs7wxsWyJjrh1+zG9ZmClButhkGKpo
N2I5MhnH9CGjE3coaeJWR9blqN6YxtLIzNIxXZfDnSJZPOpEN8MZHGf0JUb+j58c
vRPqm6pZAxLLlz9H6Fkk1M/vHlpv4iV7HTwA5xzKLWhODAbpZ3gzmLyRRAENp7Sx
Rllk8uvjjaAnMgWO3ZPm4vSv5o1y3+pcq7qkv+pDPA0J2lktQ8t9mo1IUu1TDQXl
JaEJuCZHR6oMEGQfndNcZFMTU2CnOY+Xj0OuK7w9oQ38ZMcUQ+JlDy8I3TDC51np
N3gJm+rbrv3Mebqf4rbPjdkOecjjxW691OB30U2+fwR05CmA/Mvm+J9k/61eld3R
GbIttgNgKwVhqVjJMMwVonJQwDO2SSHkd4xxJ+e8ivR93lCMOou8Vb2fhA4Au1NS
69BwlZmRfOI0cT8zfli4JI8J4A3XPXGMIyA7JRBuyPBtIUpyXCBMi4qHUu/ngKKs
zYvgsdUrvbXQ1STQZXHNTHXuDGuIR7cc1Z96BHcgX6IsLMWa75hF6TRzCN4cDYUR
eEC9Xb7uke3zcmYx0SwCRwzjkvM76U4LIrJz0qTUfTFSJJDZ2fDobGcThyS4gTR4
JhdDLwpPiWdV1/7fUs/mTocqAXDhbS1AVOAUx7uML9BD0WiIbW7KEh6H+ISbuzIV
67YqB7QydxX1sH+c05lXlL96845Bga2Tag93fJ+iPvDsi8mfzDxLzW/ZrrwE6cxl
NAZCBWSs0xmQdEFaPyoTOLujs7nfeLVPBcFXI1GQsmHC7qEr2z32n5LgkxqvOYna
Gpzvl8ldONlSUcLqEYA5lURtWqgGkcMJw2PJX7BcdSM0XLxvZ8Gy3u58axnvd0HH
GZuiWT2pXCqZLFU0NnICPy8cp7e53+pq9tdFURt8PZNmDZ+bsdXJdiqh/X+0ZwO9
aeTsh0M4yw4kCys6xqIgVGDIlVdQ5BzHKGFyBWP5UZKBQBh6sexfE8nKijaCgV1l
0lFdgNpZbwmKF4DxXCJyArknaVlv1KhqvUvQlSf/DvGnyR2OFyYmbAQd/VwlLOsL
JaTtu5ZStNc+DYItvEsKnMaUgqabxAUDnCuOsr8RZpPYGKyr1zHZ4F07vffZFZ4F
UwtnOoo5jkhxWtWt5cwb6OqamYsPOpPCJaOvPm8bjzNsP3uFvU9liT39Jugd88gW
7GcPneckiPgBBafrna1tsgq9CZMcrDLpSvwrFDWX/MpIU+wC7Ym03ucHTj5hI9jM
IfucQZQyj5VxK+Ir8S5FcrL35uFYl9sO1Owg7RjlpKfyyrIYdldKt9D+CV4bFQNg
4udfTxMy8fYDDdbjS0U6fQyXvxpm3INSFC6bKLoiT3OWmTVfNv4/lxWrU+e6Q/gp
btzwxtcmVtdCSlv7BvSl61QvQRcNYVOfVn6M7conEmaIhaJeG9tRFw3GvCBumkrT
iQAHKaH62gy7gDt53fRAADteLIOOLgdvLjaJRQrote6CnYK0FbNQ85exP1bLAC2f
lDcQ6/IVXnzE/Q5qbGlkmgR9obeZiZ48fikStOOUbeml2GsbvNH3ZME6s5tsbWKr
tppVKyjKOmEWDEeDU1zSCNOzM892gDaeK9vb5VAjex6iQfHne7RqosxK+SsnS17x
GFWKCL4OxoLZC355I56X9EEpB5DKdKeXecovNrwHY2Cad0s84UNb1/ZzdPdes5fh
qG/inN6uDoHL2mai5c6hqvKwSC7AqUhw5feRHFgVM5KDFYfDSlWu75rnQ6nuCj+s
cCtNAOLpy8XDT9KObBo1UPjKtJH70ocwiE59bxnbMJ9bv2b3a3grxvTqUBU32Z2J
mZ35jIRc1W5aST+rphJTmQ8oUUz+BfNBMSSHJd8xtk4RD/sE019ef+AWGzJ6/YvM
diGHj6So46wkZlrAgXktTUko24GJ/zn1ijDQTZB21jFpeS0y1A8CkqMU4f89cf7T
QeXN25MQrY43c6ZrJjmTsC8R9DCvgYlz/uOl03xbBE7yeAWCLrVKSflbn60HQXJe
AdH8e5r0u4TJOE+uEgNi6LuK1gzNnPa//NQ9VkRpb3U76tgWL40qS0JaFNTulrEA
wdzev3NLjGCYjuRLNelJ0fU5TqJDAGiROKhLHWLiLiuUqOf0/BMO9HcHDA2GoyD7
OghPAYr/Yuerve0vswLtYDLsF7ktd3F4IBu1SDQyYeNJFzWyqh7hLytFHYlmRV7d
Ust91yGSPF8SHlgtSlYtLYp6/iwVFF6+G6xiTfwDSeuWfMe41ZZVz5foJw5wSlrM
1O27VNLT5bFP7e0Gs4K6nvmyT8Z/YddgdEuRiOiNf31hae0xc1DSaeX1bUIPUG6C
+I2H1xgpggVqWKxZOMefIRiZQx1IPts6+AriY4JGLvxG1efloMe0V6YxhwOmD2cz
YMrHUtQ3ObaCL3+JTYlCTl3HgKRjB+4dMtIkdMT37I8jwFWcWXfbRDKWamGwtKH3
qevryDwQjWpQv84R+BGeMK4rKs/YphRPAACwOE9YfVKPQOzu0zdaAlTypTjYeCa5
Nqu9Eo4lnrTstN+z5f+I2LFTHbhz4t60JhXSWQpIwcF4ow7HzkI876euKKO9T4Vr
1TYNyzfJbSPVlqCkt75/ylXrWzhDS5yV/x0yXaEuAUWJyGpi8a9RHb3F1jVpqL2i
KNfVTMYxMbdTqbY68owCt7jwfJkRBMC2wRnYTDW3SAemRF1dmdr7/KpSaNT5oi6Q
/AtKHzIf9XUz4n1W8V48k7oGxQkOj5XZJMnMIIqtJmL7Gg/+laFz3mjIdH4jhVYV
LHyxGC49SD/LYEsU0EEJ1l1I/rBOaJQrOixrZAsM90sF5jhV9l2Ubhf67ctR057H
9wzyupbexmiE1/3K3DGgjh46M+kncIpzkE8TLNg8oBtTusckdAKEAXN6Ebl/lk30
imse7Dlo56neC+9Uh9rubLIbSPdofF5+cIa6eTZeRJYnJymW0iNalpRCsdcdSqi/
PBhlJAIZJLm0qFx8bVsegxHxLll2lx0IRxcZBdCor+9A5mkFfaoroalJcOQ/w0eB
ysNNCmT6H2XeIlcg9kN9nQSdwsYy3OSSfW+8Jzc5MqN5QJMfNVPi4Og3IkeHS3W6
fDsbt1rx38MKYCbrHamSH9azi16Kne7BBJx4f8d+ThQAybFhAfgNNEejTHZqmfAZ
+IKewH+dRJJaD25K8aAgIO7qf7Tp9YYgj+9ob10oABIQmvSeNWlZ7dQhvnOulSUO
NiF/laoa+nG5Kas1afxCNczzpYtXtD+Aqd7Gkm+uKMAF0z2jy/v05+ojDnMb48kq
z8zWP6bQijy8cjIEgPRMoVBLQNreulZVatOAMz1NN8KVoNWMQ/rHs4UjZ2+Eb+Iq
b0dXWvLfCu4gAW9q4nNUXEJxmplFW4IR8Oj0lO4vvxduyVgG8sP3aWREqeWoAbix
fo6AHz5gJkHxBJK+MjUsZCUWU4SCnU2p5u6YWBMZVaPKUEGRwM+pklybLvQtV6w1
vG0QeVadhCauUv2njVPVsydLpuJtdIHr7hQ+PsbC9SQNq5lyxD0r32OfhlcwAnvU
4z6WA82rO37glMXQcLHqygX4S1IlIh455LJnVjx1IhAIn7VQQIeI9Lk2ki8SJqTY
vrvyE0O6u2KSo8B/M5f0uxYq4pYWk3+x8e9PW84/wa7rho16hdlNxyCHzGIJSJWt
NZuTrwpDVxPx/4CsRUnep+lzsVFB53HmM4PfDP8gTCHWFvZ8m7njClVGw574psxe
o7Zugu6VZsPw81BfG4PFmLhx7dM4Zy4C0mgkmU6aYOXouo0DqZLsmunO9gc7GTNu
1i7aRkbmm54gDPfvA+IyWsEEkrB0PWZOLh+0TdxRtUSAlw4W1M7AHnrzd6XR05sK
8x65sB5F5BhNLWvuRkB8j4LWIHOsT2iHdestG9wVQvCNRu5T8DhGeUOx7P/26eXA
XtdZ122y1fpYArkjh19ZUci63cW7wX/1+HH04SDsXrym8MZyDm9CJfOOsN3rkgNi
nKQXwXgqNXhe9y2JTMCdGcceeyY3Lb/Q/ZoUeEyjRBxywBN1hWNAgoarrm+/h82+
q5wclBWzzdKNZ+zJIVoSwBtwuSU9PJwdnZPpImekud0ud4cT3h+iGCj5mpFoXnfh
iQyfjMtLn4BhSS7cmVm9xMT9dFChmUZxgq4fBxCHxcw+JlzG5YUeSEcURUgUG5oV
EruR4QcuN3MhSYy4X7ns2ijhH/8HeJtvgJCXRcr8FmsZVtlg5sReaq3Sq19Ghfzb
yBhqZDKXV85kVWvNp7n0sZl8kKT75RxWk4Jl3QLnYXtj/JFUlTRsY+aEeGDOin1T
CGkCFvgSNISGFPPfvRalu0NHZpKqy0e3Kl+qWYiGHsYc0nmLLbEIb+FOAyxEOG7d
TCkimKxLKRNJqRENqqvTOz5y39GZCwiqaTcQwQG9VRQKZS1cCO8yKQTq6c5ttzzW
V0SvWnQRbNDIOvXc8m8hbwAjYgZbEHVpSomCdTrHHJY+16Dx/NEXHFXq90eadSH1
i6azhssLOkIEwF05cwHI0jH8jL58xJi7ey2JfBxGUXL/5YJ8afkN2MzTMSgqE8pe
0DUpFcJQz1VTukIzw8AU2KT7PTZMyOlP1DLYwru+0h5r2zEZX3NNg7vsefYy6QC6
PcaY8q5RJbykFwllK4iM5yVUViUo9v8K3u0/C66XrDFQOOVv9LxMpuBK+rxG804s
rMsJ+3n8E/JJ4B0MpYJ010IbnBRvA3hXOVyY7RjD81QNaWoDNeGLIxymLZpkyI4q
iF1rUlC/UlBooZs7qRTb0jW3INtGEbbqTIx4SuBYjv3pr+549XIzbvz+RmAF6e/7
2LewafjTraF4wvDxMam33b0R75iyPhR1JtVV+4caj+gbc7n7nysyNQgFhegY5lHs
f+NFOghy0kOQgTm37wEORitzj6P5E9pBQJTowYe0EnSPT/478dyHztYPqFqx8Br3
9jDLbH+TtLP5hxVfMpI227bbjRVpFV3lVwyTlelAC1bXcDygm+V2ymEqZGOe4z0Q
jS1DE/wVaitAsqpA++EI2mwR7FknhiNpMPvdL17EONaMOwcHXAw4WGjtzyCUt4dt
F42zKq1CYFrrlz3LwZHh5wsugNDCRnx2102cqcoA3GeY0NtEXVof8wXMYFHGPElD
xvseiijTdmEbX9poiDlkPH/21nswSpa9kTPRLkADAzR+bbPriBN/aQ7GjLEXlM6s
tTFu1bJUA8HiICzMyXnf8wc+YudFZTEUPeOGpWtuzegsIo3rjfDUoM8W1SnjdDhL
zqgTSQImgjzKcy5vhNLze7zX/riM70Q0cQ3H2ijVksy8euCqZO0deTT1Ie0SEuFO
XQvIZ/I9Q1go7zhH+G2+NlxTOxrzmoxlDmlZmTFCz7t/MZdXDMOBM95vJ8KvgflL
AF/EedlHeQ5s5PG2PoOtCTHw39Pu2rBYfKB7zgkaaCK/FNULcOz71wR++PHBLIN0
1FFbYWTVjpQOeNLxRSt7BfpVK/BHT6DtPhcLsrkA2pWktG0sj6HLtVWoj5im1ewh
zxSJtWw5gZN3iDsRW37po7H0StXGrSZX66C5Fj11k+73N+pYmMpx+mPiRmAhYOXf
SuWaIejuW0IFZLN0hCHwBmo6GBL0BSvMz8PhvAqMuCpVy/Y4d04nkkpu6b1Ike+O
c2icGYLhhI+CvYVaG+oN+UF6OTwl8IxA0VgdXV6kaAwt2xxsnDPMkZJuUTFodjL6
ToJHh3eG7rlOgjFmaIVG07mQq1kk1LdvJeM367igCQcvq3rGm0YNTQ/FckJkp70O
5D3RAHq8t8Apcy2jWCk7vdUlX1HFnQ8K+3vTpHb3JJ4wiLuX/hEjQvrYPFJZq6Xg
L/DpgXTR6UTtVazetjf/mSYdPP7sRqqfx7VhdMjOfBUzo8cJSDS7EaDLZnXRePdw
yat7EkbaWH1VldCnKBf6q++ynJkSB5x9yxADQl+uLDFvyNO2r/pYuuWz84Ba+qmi
8V2AvvLpB9+hDY/ZlFUPW56T1LxBYG+//W1AogZl5K2oimT9jZMIqrQyaaNgD2Yo
a2qopnhUfNOpz8ID/nujUDmqIG1wK5x1/hYbSsHrpUR58EZXPHYzeLrDEmXKgd/U
uKchWxBhbTZeXJn7c89+243M4LdvfI4IfYDA8vPzRTCzKDE4ZjPcCiMEarKPycsc
1rEZFe7sgszay4PCk6fEP5y/hEqJ0RAb+jWv3sY7E8YHHcV0EITDVLnDx2hJCQHd
dApZVPMfRlEBAK2adcvOuTdx4RqFHkmYbMpolkPQ24qQLlpUhl3LCPZ+05L+SCWT
HLJEWycDnib3GXP5I2jUZ+p/OsNe10h9e84lB/LmVvKds2MXtFVZNuWuDg7eYTh7
WGGhk3Rvy3gDr5Z+uyrNtzd5yiGwxyg/LnvdIyqmoN4GSF5shT4jVjASX6spmwiz
Od+pYAiAd1753jpWroJUUSgsDtbYPdZmTbqRPLlD1CsB3Oed+xLWtbzxPW5IZOhH
6j7574NIBuTJSXya5zSf6wKX5KINfZHXtSwYZJ0n5phpwSQ3or0XS6sTPWQDRLgJ
UDr1nguTLxeC+7mYVyL7kN5+JoR/UPGa2tXXZrD8+fjBfgjdP4joU5ywrLrAK4rJ
x09vvIBFjpRVytTqey1Z6hqJNZ/qgjN4BpqdW/O/B66fLTnK6a4qHPgQIGDZ0b+0
LIufqvb0+M5FJrRsLlev3p+q+/Nbc3p9ogw2J3ko/jJ1GdQuB2cwF++W0Mdf7yCR
yMxeG1giOQHzvyPY02tfdZeHzWTT+oZbvoRU0wbxL8SCsuk9zOrun7bUZN8WEDU2
QFcDz60aPMhzhos1/y+SBude7zfUU6Nk/qGyoYeOwj34kGuqtL7CdRUY6v+cGPgO
myCQvGqKCqx1HwI9Yt1hJ6RwF9ncMSJrvhcupoN3mgPxB2y/E4j5XRPByqzP61eh
H9Z8tItTbRkMaHMPNkzRV0ZHobeJ6zk8ewyWcK5wXGhflJ0KN/LxQIBTD5ZESfFE
mQoYQVPwL0VRa/SvKQz5OTHHGp1A3FUiV30sWQPhmEzqvobiL8JwOKBv0DWuq9fW
UMtj4v8Y4okk9Ud5FJImIxXNUsneCIv2ZKTbaAxiPkcY/NB+zVMOuIgWwFm+glRS
CJF9aCZ8oub+QJ8B8FOI8XqEwKL11mOWctLho2Z/Xgz2Xpm+GAlqPbebGspqozwt
ClBZKUeYHarFcY8z5GM1xuaNN+rWqJcwlUsQD8k6MEErUsw+pD+1ph29IlX4uGsj
4mP3LJTkVzzp4k8Yxxvrvl0M/Hdagv61t0HHgdZn7I7Zdfwdx5RpGCa6CithzUeA
2T+8oNTrhs04dnIXe2umMtpNF+e89W1qX1qs2GRZi+/71RqIpjK3r7wlkvtmQyX/
fum30xfWEpVIbIUi4OpbKVWKuDet0It/m4+smj8raZGAGAtKE9D1EUSLIatw6l7o
ye3XV2yC3QT4iIDTZjLEak2BMprLPtyteM07zhgjsj8n6dVPs1UbPU+Ij8XAdxhO
miZhPPFyCfJhlQWIsoYfmAP80YXjDhIR6abB9ho1kN8IMgxlvU3K5LsIY6ZQxamp
YX8WLuL2GJpw2W58nHqMfzngJcPrzcRkeICUEJvQWFIEr8JwO+c2DKvvpwv3vPvg
tOTz7ETDXLyxQAHh42KP7NAthyOsb1gnRRBSNq5vQBUkLjolXnxm9WGf4L4yCNqO
VG/RsmRvBhCoH0TNUnSBvnsn3r738eEeS3YcN990NdOvnapmjTVsX7hbSu0YLr8c
V72KVi+lXP5y8zE1nkKvXNPqG0v+ya5o/MZUyeheBrad+fjdQqMGsRLK3G6RZP4L
flHqMI/qlSN3hBcT5wQBO+6UaxnZZQ/j/Px9rIlfiBhyTSBOV3HTMWHtiox9SwSF
dFzN8PilnnLP5JXkZ4+5du/9reJ+6syTNiwlPVROZ6S6oMHiqI30FX2EdvJLHsYi
bpcfcpf1yAa8L0v81XujSarbNzWbXnx7CVgL1QNGvbXlF2RIEjOYhOB8wR2mgW+2
6vz6FFbOX96ktUGOSUGRPcMAZUTZoYLbZmDPebszpxcxTju4iJysTeGARp5z67uc
tEKvQaYFwsu5WSJf3xtk/0Xn0SuAsEkRlfhNW61P3DOLhvuvxESu7xheGZH0vqxv
udAzTk2yAxgscqzj2CIOzv4Uhb310V40nURCx5ffGc3SbjQR+zwAh377Rnid/Ozf
NQFfHfXrh3pXSSofcWzEW3TIn70Uv2NhatRksDHFsFa4OyQvm/F3jK49sKsqJ6PD
NI8INwlQFC15njUUT2L4cnbW5mcozps1Q8g3KAi1EHLTzrBGf1cVta/iCkQgEUXN
JOe68ivQ7A92u5dqf7ZufmgUfHwJ/d5A7WGtcDLbJJqHFbiJ/SKf4dTZykptgCOn
Dyzn8iwIn9gVaamiWNmMmshQDcKyKGXKOPNreDzBuhtAcMH5Cux/xteBnBGLqVfX
E5oP9kwBVxhV58bDf7gcimrj84+ci6bbzkayBtLkM8AIBdVOaJmw1a77K5WquGtG
RAi8/3JS8Fm2z6hh2lzXYQTrb8ZKFmwsY9FQ8amA3Zjs+B+RF8SPq95wR3H0i+mb
xIa0YHBLmWD0vaf7rGYyrCKQMYi3ps8piYPgSGYoljM/rGh2d8ftVNA3QQcIHRvb
+Cz4SVzubGbEZ3erKtPopwwZJwkkaSiOtrbgXOpV34qaIl4ZGtSLQLGAv6AKFdSI
Nstj1NhcGNR0UI23PkBlb9W+OlUEaesasqS/XtfO3tldaW6k9RmwOHTPe4ApwyOE
aPr8PAN0PIP+vz6xXCk3IZQGti+gQmHagO6DfSN7dw/oR8mLkXzq7ObYr8P8205U
FCoZ1W0kdnyKszW+jECK4ciTpi6nk5t5rwyklQdR5k2YVaosgmXWiy5aYm3iGRbi
q4hpi5nLE8TEXOEN0EwCGh6xzKkkCy5jV0iRUcKuPV0RxMO7WY3rEzqtmen9kSep
V7omr91pt4GKbf8JgpWXZZ1+tKIXGstc9CUb5sRKKtNdQJD3ZSIF6/mNqZ6ZS0kL
vabNMrZqZnugfrIuKFNpc7Zx8QNaYIb8zQz5+5UEWYmYDzdeDvk0FIZ4rcvELnMF
Pq3TsvdaasaUQ/s/IiD/zFgFDBRwm2Ab5fvYZ/LZNKQ1LOEazH9kqbaCBaOSRx83
0H6UVbYebN54zGBb7g0Tf84X/xJ1v9Z71X/ux+gW1DcLipbtCByn4gSGa7naHP6w
vAxQvFw5iR2oGJE/zDEygbbNTlnzeTWRliDKYbxLzuafZvJ8HPZjfrmqlLkv7hrs
GxacdkhdaE35hGNEcqU0P18nR+pWpyWcr6P2QN80rbDDQU7+MsfLUmJi+WLRqxxI
jiMZCph73gy0xE3TZCxCAYRPgE6iQ7jPJhb53Th9kE3daU03XvWL55Xn7byt03TQ
eyekI4VcC0nWTYFce731tSgwJAMFI4E24ZzRLZfruWIEwetCa3VV+0kORA5O5XhL
OmeqK7LQCCSCOjTCHCUJkW67M3hrOrdx96+q7hIRJBr47wr214YgOx6sQiGok3+t
HvUpLIfB0OwgVAVoVU+xEiB5FRBrlpSiRVISmRw5aGXVJu5vPOqbt1IKfDB6Z0yq
/9+RIJigKLo+VnCdoRprbz5eFilNNvA9rIrbeYTq98ly9zSRZpWd4x1fpBvC7l2h
hIrIUCxhxMOHl+H0vv25Ug8LqCGmgz40jVPOHggY3Ag7WMqBLo3CCcVXh5T3FBGp
fA0adv8WbHTlDJ+36d5SYiIUsrHKLZAwXWf+RYY7RKiIIgR6xZ60+jZTU1BtcoCB
tweKQE0w+IuFTbGzydJ4K+Y37g3bNrShN+P0aghy2larN3QVcR219qyiKuiVIlSO
5fZSHR+kq54r9ABI5mpsgwd2kG9pDtHL1tgNPudV7nGeqItRfuO1DNI6wczjmnZJ
ku0iMcIVtbzLJcksRp3XqhpbXxflNDzn9LiEnyKLd5isipGByIZlOEwnu6BQZ9lD
oDAB3WBG59If8iUEoNIp16+LY0fxE9nDlMaVmxR1n5ggzCMzWIDItW0KPrhQCTkw
azRhjYkVDLXQyjJqK2Jtl8XLfd+3MM6A61sXVK/K+b/zyy+z3zzuZsAru8oLUPDR
mOys81UxvbLmuFkVXrABE/3w7XWnmhSrDAgeo0LavkEZltaZXgSe7tIeBezN4K+Z
Nuf87z0ahR1QosE77SFe8X68LYoRyaUD8VKOSHAQhuhRnuffcaTkZvx6IpFmlMSX
HFanpXZe+pEPaZrsxL7nWL3R3guZ3uq9fbkP1eFCLABd2uJszPmJDWFSVP8aqvos
h6aJGah2mWj1lX8hOwC/ORsA5hqfnjVZ6nnMfiNsuIqWhuKmgBQIP6sTf+Z0W89V
fSS3w0nsSOk5I0hfM/2BPDqRyruTv9YadodllBwK2WcJsS9kbKmje0mBiVFRYhd8
k9Z9pGo36xwaVc5ZMBAQQag0xiUyHy/1Y49S8USG3LHvro9lRRNeiUVKXu/iaCVb
qCxLNNPmLABJjnztuyPuGWHUAui26/K9Gy1LO20i4dZwKKDfdhT1JDf463kszAC0
6Ymhicf2QQsA2zYyvZiHCZL1Hu3M7eQrX3bwEv5cKW4pAh3mw2KtJ0SM9ZON8ImQ
Plh3dkfCOiwpL2a65II1YiZPnHkDYcc2SI/WkjdNtFMlCthsS+9eYgfGYzTXdmoe
R0+IDHb7n5auLIIl4SriINvR6moWoaXvEqFyoXiM1l2e0hMQW6HTrzSS1pf0gVEK
NUSyI61wiDMDdUMZUywBIXLXp7PL1rA0zhAqXOk8hNzc2KD/QIbgn8zpTvKECsRM
wRwoWPzG3tEY9ZDFLfietRqoEddR1UgxTbj1E5lT6QOXVasFTZT3F+TLREDw4cla
98dBYnekdeYgitTzI1s9YKfz/bXGWlxBL0S9wXOz0oYOUOp+6AH0bMNCBzdvnJWV
nLz3BGnUyAgAtEdpdTY5cXbwNF+aGYfkp3ToJrJg+nj/bNjUrAEediyM8nAJjVIm
8C1/haZSiGAipB3ObyzRBogaBZu3aElAhLf0LmHvmONw5qGtEhxUaosG8z74e9Jl
drDZdQo7hmzqxziAoXv5cGa6sfMnZZQNh4dL/OsjE2duoMtrnEo1+MVoDKL9WHhf
ivf1qaHuD2HZk5Cgvc5ooO7gvm7ZGOc0PAo7uSO+9AAYN5q8GFGO/wkKuPFoBl1n
cve/FvJ8y7He2zwHfqDmo6FFf/F/O4MV4034UHhP+SfSYjem8LG4hH6fiiNz89a9
UxUJVIbbSxy7ZOpZkbEC6hS5Q9gVH5/ywQcpS2t0dllXsvzC3scr31sK2tU65AbF
ncu0Oc1toJ+zpGKoulnktTST5uMsox97KSt85NkB+LZ/TXGPVx57LwpiVuMw6CUC
3DHLlKqABw2uBQfmR5EdI6u28UXAEjUJ3KpzLr/jqRuu2StSrgOuWn2UxVnMU+Xm
r2MPaX3y2T5ge9EkuDvsq3lkDvsap0vwniUOI+Vr5p0+Q0NWgWeT+kvCUQm553sl
OpNUloAOgjoO7YwJ2alnDZp160ZOBrSuDSJJZw5g3W0W7bDRG+4oAaniSVp5sQrD
q5JfQonuhpFPQzNb9NN6JIs+ArakNAS3N/qzad1h5CFTIup8uXL3WK6zuZXGFH7Z
fLOm0gV4pba9xWmyxbq7qp2Ck5pxxsqqfIaq/9l33nO3ORqh7yrKF8CpTji7VumI
L8amygrODcIQ6s4sJ7GP2syE262Wowqmpw69ty3kBo3ILM9qP6VDaz8ABG3Znp6i
ku7H5/L1bhcOH9tsmvpwj5T9mDo9LvszztYUmyxG7J+4PdKBl9mWgwCxbSDhpI/k
9CDuMp2S+fQZWbyEELR++1x5JEE6DvQ2lYwILM+VUSHmz3ms7fSEG+LH0qtU4tcj
pxWjZzMeeeHcMrmgbodR2Si9RqXgkeVI5Bw8rhBFy5d90UPZF4JYvaIKHktjRmqx
n68hcgbeRIgZB2n/Ak76rZbd7e2zU1M2IQ4c/1+OJbn+wMOflJk2ZsFRbCimUUaU
Tkf2bypgBzACOR6ryay5Z6jvtfgQZryVE6cAc6X0KBSf7Tv7V31BI0h6rdyjIgAm
wOvecNb59QUXHvuhtVIitKhuqSF47hos9oai0sKnRQZeDzGQdFI2hc+nTWHLQqMW
QAGJpbkGXlkvuRH9NDoi3CFOE7UkEEdWZGfahhsmcMqPuNuKAe0QjWocbtpTAQWF
Ncl3ulm167s/3WhVqf/l2/e4AovdcjSOfqhyuhC5ButspNPpQkWkWbrBl9jMHXwi
eXtrTkYau2cjxo9zYuPcAVhou+su8Dd4Ng1L/GFxzeDKAv/d+tbnnbhnuOteKdVS
YI5h8JMkuFJL+G+E4OYR2VTOeG8kDLpajeAVE9HXosw7kiGmNS/518ttb2FTvbzk
e3hur+ZKN5hY52Kq6nzOEZpGlHDlh6427zmWPGGDMnrAro0PbG7Co4hym0GMjcvN
8/8t6heFX7G5KSBQCQfxcgH+yI2ZLd6hNb3vERdCyc40Eush+Gkgu7AYKRdEXJY5
y66bNv4JE7/DSR0tocT/WUbl+g2c6cJrX+LkkEq3Go65/Atl6BIv6/AYAzqHb7Pt
40OshOoXLgGsM88HGFvawQjvmUs2iJpQUwUKvhx0mx4ljcjogGO2jhP0PBWuY7Ox
QArVSQaff6bPIFfK0vNAqMHTAyvqVgrVsyq/bZWKeaRAnKt/NsbrYIqzYqVkw9Bd
4DYEuFFEamBXOuTRzwr/DZbGixryNjPPOZ1UjjKeFuKID+CUOnznn30o2lNNj35L
E/6S3TjfBFz4zz2tyn5/niWIGpBndXXse80SoeWuvt7iMG6wuSscTSahOw9jQWC5
cNGdW9saITPU5GB4s+Wnq2G+C4s28i6CXlYWMoYbpE/hfmgGcRVssHkdBgKrURmb
cawemtKPAOOlJcvaU+ny2OnHV36aCH2/9wVdoJo34N7k6QwBCQ0ThEqDwjX6hceF
bEQTtfsAtlubMd7v8m5tPhKscsC8lf2lr0ezs1n9uku+brU/RhyOOSOsSwOTugQd
IB3ET7OJMEOvq1XYeZpgPqoOz2z/L2CHvQIWHKwATcuKXV6M4Pnk5/1zDEdk275m
GKndg8lmbEq3fyGcBy/Cp/h5+SWh+pOT1wkTB5YHhPtJusTmbLwQJt1A+78yW51a
pk/mJwxgGdmNfaXHaE9aw1O6Peu56S2X7nEWVB4yDTT0pVErRSw7g97CieIhPf4K
e5I9L8ztiNyKa8ayXhHoFSwOc18a2P7+upgMbYM2J3DhBt2GuiuFZ0LIA41nke13
QFT8IfNeuxflwrsvHUVVNZKCmQ25xH0SPkUS1e7zdfkXA8q0VjZUg0RcW5h97C0q
q8JbdslDn36Wf6xSsGVSbNES2kKY0dSC5wBscaS9wsv3UI2fFmFHVmCKzBgcCzjL
hkBLY0/4wz9QCQm+3Q5eAITXAqy9m59bT5wf6xmUoLj7jQmnNmhWh9/zATIfuCS8
E0F8snNUvMt7GxbhqOuEifdjn5jPaLp5JdqOTttBt9kZf7TuFwZsXJGQJ0x1+ym5
zwvv3LObHRnzX6gGPgTANvV0LwarGq/4iw5VeNa1Jcuikmq3RNq1T3389rPecj6x
H00N/AJQUWBkHSRAJjJxQyHlraIkxQpKG/E03SIUd1BnjUZz09antI+EfmG8alMo
w3CJ8AIXMQi3EPNRLxTQOLRVc+GyipI/JYRlzk1myRU5EzqykiVCev2ImIoKVxBr
LdgRDfoNAp0OiUVWa6IBbsd5BiGyxJ0OugCSNraU+7m8rnQTsu0b8lLMi7iqFMmo
Zd+2gcIBcLNMKMIFZY2pCO83QbTvJptbceM1VEAW/jq4DK14eG9EDNvK30qEkHXN
KeAqwWQRs6fBk1XVp4DVdrnIUIL6D2R6ilUrQ/NtoEmE+QJAXYBDf86otDxmguSk
Wgbwoyy1FeHnODk8a+fXUshH2lnFK2Zybyve1e47EI2HQ32u2JOvVmGHGC2e+kPg
SOmVHd5dEJH1Qicp9YCQXLrcJRixfCVNTDoqmqblnEzEGEkJotYS5eZ9OUUqv64k
1+rxkjlgl6eGUwqpK40Cce1oJGc2/HtNYOWvF/GldUvk3Lgx4K8QdQhd8rzxTTLw
wrD+YtSiI/B1vGJuJ476BN4GyGouAftzvgjxWa8I8hPAbTxio350cpcv4iu6Rgk6
Zjl2aIavSEisjPritwDusOsgEz0uo2TGkDzpGmS3RAdpZSgbsP2n3Nlkp9vIm6A0
H7T+KwrsbgBXlCngK0rO0RKlWNTKTcQdjgKJRxDzjGHbEzVryrX7MhGzRr34AbC3
vT16f9qLVFmdyu5y4Oo4jqTrMTRJT7LSShPOYFOWcYLDRCPVMGkY+bujQJeNO07N
PIqvCJNf1xUgazXqMsQT10ycLCHs0Eh4+eyNHcMD0ahzYrV2oHGLWr6+CIDz5v6X
gPrK2k56a1g3UJ9j5Vei2CLgmse0raJdJOJNjImyt6i4D5VB0rmKGIpRnYbMGGS3
MpaJr5DWG9ygLajsgV4kr+L/iqWLxlLoFXC6PG7hdNiBgITPljOhT0QMSs/LSyTs
ZMUiu7SY5xA4jbnLD2rLlRlDffgN5NkWlFMNwUEvIR0/dzSdyJHk3MODlUsRGfUa
jHI4nL/+8w0kAw27cC0jC43ZlcyNsGg8eebLJbZXtEMf2i4A+goAVXJ+hOy8t1tp
vviWPzDrmmYKB316wfH33iQD2UV765ztxCxHFwgHN16osKhtNb4yDjvmAqiVnSKs
JgBkiWlNOmLedpriGkVdmoM+8LYOoNImsKlCKTkF/Pzm5xRPfa97EpXGlIsAaSOU
hr73+EK60glKlqzS7zTg5jAHSngdC9dyQJrR0+SKk7aEHMIJAsGk1wn0MBQcvNoB
oMA85yeLD4yq8ubxB5ufAiUyFQy6cUX+UNWzVcNfiCQcT0VC9RjxVUpaeDa9KJ94
p2sOH+c9FXKaYqabLH28gawZy+Uwb3jxSV1OtBCs3R5HPmVjLPe0O1opLsgiX+yC
eOzudmmARnHuT6Z7goyPO+/yDS1Vfd2L8JW8O9N7ARYjStWfPr2wdhbZWpP8yuqD
+mksdCb0Z6Gl5O95NhbrSNXyC0NpKSq27DYuu297CpmpFBNr5pOCUdT/PcvUPhMV
sZQYJUqy/4pDPTRaVl3aNkotlvVxSEVBoSQ2CfwkaWfC5EfCwhZCn0yijxg2ayMN
85yaBtL+NWEFLeRKTvwwiz2PSGZy/WKNwLsG6kHAMxDj7SCghW26lb+P63iTmJp7
mWWMaQz7WJ6UR+9JfFc8780idyxhJRL/Nq4KABPHnNugKQ5hxxMAjNFcj7xSa2rK
91kC8OM2CqeY/k9rUnQgoxcx1M5KCOJPLEOwCBTNyJulPuy4XkRH4cbrOZiGGV+k
BCxSfATUp0tSAB9xwxpDS93zZumNV0sFeKO/5f0YrH3t59vBO2aQRazVd6kGX5cu
076Bp1OYrfNa77OXBlxQVL5mkEQA/T1uj2j5SlBXJZgnblYIXuk2EyHnTrxFHJ5t
hMP0Ie59NGq3YtrRkLcyRWYE1svQ7jDNOU7YWxUAl4eR2bvI6hwArUl5p7aL67wk
E8tvWm97UAMy1UQLx7mdw2LzzQGlBlufVKYUKTkFoPhHMelbNRBRD/0zNZ15VU4x
wegYElT8rN/GRQt4daOw+R2EK/Mea2JPkOJ3khY/36lnEl4//tUXGIITSWBcQCFW
ITvm6B2TnBqYYrIUbD4a2ofLq6phfXCRqb3HNdH5vQLDK6SaMt4Qqi8BXc1pKSFy
NbGMDogLDM+FbuUfxeyuDP4XBvZUYYTU/jG+JNJw6fi+CsmcRXZYeZLaTdgm/mCJ
9WYoi5xSUF7d1A+nL/zGioXyHJz2qEMLbQwzuz5jTnhtCyGNHQ5Mz1MXiJ41HWsa
JKMCkEpu0JLG2gTk7ywd31GAL9BpPf+Nosr2JgbMhOiddveVvHo9qmGFKrakeXOS
CgT4zClqeoxu50/kUSd9ce4WbTH/fNt3T11wjCEEIiQv9job1uN/OyJ1i6vh/bZJ
Qkb+el61/32VQ+orkHMxZvQCSx0sCo0aq9hm1HUf19XOfC2mAZFENucS2c+WKv5x
Y3gH1wy7q0nkRwR8rQ7Are05rJmOf0l+AMIk32Lr+Ko3dgAnTNGCdwl+bUBjpmJv
j2s3qtgf3ahWJ1XaxMG+6/AXhFMt9VYs/WreXbse6iDrgFGLs/BvhD5/yicj7Lo2
fM4ae4It/CyXuBWQUPLjNEdwHbcqwXPy2164r/GvmW4kJg6N5/DKyfSQbYSsN0zO
sLq8Dx1EtKAzDQe4Lg8J9lWgbtM+Kn+hLY7TFF32YjBu7eypF3CFWDaSRiDNaRi/
QWIlngZgsBc7XhVT8MQey5Af1uDQPUR1kyZyQufop9dT/GbJAk36p1l6g+mak0tE
5ugCUMqPWphxq3WRFnVOWbue7EBAlR8jX9tTwDd80FOoC/bK+3m002n8/fEqzJuL
eqrSc9k8DLDh16ApuZVHbe6raDIbAFNgeU1Cy9JEXgD4Awgz2nh7wBJyho5gNGN7
3aU7GYQXqc2G7AJ2GyKc23UdtxdZi98lnmS2uWs3avL2VUvuFiQqXoK7CPZ/aTBu
vLho6kNJ9AwKMEDy33smTzfg5Lh3HnWgafRrNCiCcEdRdCC8PjzW4qomQErk+5kj
xXa3vo7H9vZ1WLMvNE4gXbfYhpjR1n6vMDq1TNx0fSC8xKOu5Il5A7thh3HcrgZi
h55CEfRquj0wGnfjkEAwzd37HGf8fJBP8sMfVY4+oq+a75JHeb/AeK6Az1KtTXIk
Zks6ABa02EQexfEGIguXKMTmjb7cXnaREkN2V1aNEevzPSwDE1wa9gTI/d6qVg0r
KWwus5B/LRezAuMoKriH5u8j1Orts+VSPCAFo0sWLx9LM/5vESy/mrBBY4pNbVdx
1zLVRgFbyisKjasx0cXVQeKy5bkP7J2Hp/5Ylzm3vs0Av9qnyoOx5KycvJm6taHK
gUv91VAA/qMHSoHf/or6yBmSCGg2n/RK8Ln3jc5Q1dh6WORDPA+4yOMnHd9zNIV2
W8F8FWeTlvWwcnTXJvbvWcpdD6QWq8/r1+vfn+t3oA/0to8tsXjwpILMr/D7kVRl
kONrNJdulf+lx1W9fbtFiHqidSX9BUwuJZng8gT9pwEgcINPlJCe0LnammR2zws3
NH/IWcVdDh+Jg8Z2NHaS7PTOXsinx4FOYyU2KZRjrc68epsaYJtxz8hEASz69Vx5
DmAQiiOEn/GVmfUP5eOjou6kD9B/dnJZS/zXcUTzKxPmpb3geGF1A/Ww4zXgZMI5
y+ynsZ8D+G67bN3XHGciZ4V2ky3FBD+zQyIULY1SQKeKQyAfUfso0N1jG6dr8Bnj
hgiz9KQRTvJ0pCr1e3+qRDuyKWRsJ2MdDrTfZ7jCkmbLTBekqjHjWZiN/rIdc1EF
E82nxgWUkEAEHElPkhTXAU+NgQz3WutnpiRChD9sr3LAqsmj7C+13spxjVf44vvF
2w5ZlIaINXO6FsFEp2l0J1+GWzrebYNajJRAkD3T5rUvaEJcduFL5pinL5rLKo8a
5n+oVo2G9eIJVY/+8lKXimqBga2FXlzlVdzznNJiiUpRL+zdepzCF1hVnaVMCJ45
usyInhSaeXfofKeIKWU60r2p1DCc06JOLJL6n6V0x5BuZP2uEjMdy0aJhyb3Ll8k
sYjaCT0XPj6JokkVKh+0ipWsUk0PnpLVL/2OWW5Wfrni0EYtwlG+PCiPEAKMqjpu
8Gwfg9BAkgqcftEiPYIbkWtWeWpK0HMTCZPuw24EdWUfn0Jogs1r8N05VwcmPzq6
kFsV2Y9peSBIw5ElO+WB5qQOpsnUn6nAUTOVeL5HZ/aE58kWG8p1/fZZoIZGmNJU
gOweJR6XsTxywG8ZUjgK0QXFpY2QprKcQ8erdueakARF2Nu4QaR+5s3+nUeSKfjQ
mq/Xt27s2aynrYsajWLl0MlBKL7cz+r0RgUhQIwJA9IRpEybip1D/B/M9MLTssLm
OM0vjgZkB8oI1P/hj8TTAYG2+fxfnCZ056I7eTxttHh0A81awxNxkJrE32uxzSPa
2ZmN8UNvwvHNXfvB7Iw7FqHFnFAYPJep7rOs37POZ/kMK/WEhyihkMfc8NGXZrNh
g00+vl2rI9CvEutetxQrAQrl6/13JHNY8C43y0q9p5qcEAXBQSJHGny03wyDvxZN
umMTCSBUQgD4MGQ49rbcGc98Yr36dPBtF6caAfKLDHC8Ve2ydoOmCjmHCm7o+gVE
ofwEwu5C4kGtUk1dN8DMwfcersFUaxCCuAVyqn2sUzN3LdHaNaF9uYnTDpnWtSFE
hjerfA/UTNO5W2/1/tA1y6X5fTW89lWmQ8dmZm0UoCwlg7jxdmJocYT20mDnwoqW
ha5UpBEwBVH0QzZEmTyj8+WesvvcbH5ZkhHAm3AenJmKIH91s3t6ERbnz+yKk83Y
hEJWXdbHHhcrE4Sv5bv7eqcwwroutDa2RjXHM7TFFs9gPwDrtHrVVTcUKAeGyu+l
qzCvR8QMla/UOl+YxrATVeJv3+2N/B4Z21v4VwJwZUPsLlF1N7DkGeNYVaybhiRK
XS9J2w3rCGkSVaoNgEGU/zvpZg+s4ymfUhknI930D9bQ/GzEk9RheSVJ0bWspggg
U5Foid1GzhmEUt1u/fGd9NzydnpY70dPwf+W7CqXSdqdKsukuFRJZJ8t2I2tUgNM
ANr5DlP9qQ3sSH0muPxS1NCKHxKT1/plNTbrWod4JdP27exTqkvssU4GWsyNIC2a
Yqj0TMs7igu+ovBbDMuPz1e+B3tMcVOjvm7zXLBu0+0+5hXQ8CXwmgKUDnuxeqw/
bXqwWVYzOreqe4A5/T4xxzvHqA/5zrYxeYt6QM4SbEmeNUbTbuczZuzNOfQuSGxD
Q01TwnTMeSoSohZfCEjQreC9P735aJn2P9SZMXNNjIb8qhqFzGnraehcI29/rdza
RrYM/AnW94qEeQ59n/MtmykcUF25ZIt8qkyTk8oZVIgs4nsB3ZGhzEC3q85HKGD5
eZpOdpzgqYdhIhu0rb8n9McSLOg1dOPfKVYkRErEXDskfkp/9HW525nVcm6nTnGQ
jkJh7o7Opd25l9bXrqooc3u51aYVRCShzhztJjEpzGUQz/O6AIwJqDOM8Hti6Aoc
KGdFmYeh/rFyN0OAE1AgINqjyIlEVnwXmZkL0iHkpY2AG/R5IOuEF9kTcvGwf7j2
KpD/+C4tvcIHiBS8n/Xp/G2PDeswpFnpwFjIQF3w5s3LVNYtvWvh9NHLNYLOc8js
VYbgfme9mlu6/M9IlE3SKt9YnjxmK++5HUnuILAWwQMIB/wqJlipaiy+3Fmn7Pd7
I7hRSroNVoMlVmVa6vG9lvjyXObxGJ6ro7qyiZif/IDLhrH6+Pbko66LCD/HkHVE
vPZdLvL9lTCrtIicaWtzPCJH7/1NTJtVfiaEKYVpEW45YYE1hHyNA4w6MfodxV53
MRFARRcPP0dTOkRyZL0xUh0AudgxxbdnJxVR9qiPY0TiT8hWnUD2lhOqZeDryFTj
Lxb9uoyNMwUQ0Z8maD/w6ew9RpfNYDeQE+Tc84Mpk6D+iAfd7qEd9v6B+q7GqkNu
pZHkXxDe+dHJpJBttZ1GqvgVumQeXGBYJwrzDk4aTCmH/I2UGVPdh777r+Dybl43
iJ4SzKEycnEtBBKdaPQhUajWnb64PGP3LAqS47a+9+Et9qrbZVJ2pg064TETmfCg
WdgKqLmF0zywsGCTNe55MqSPvghHy5VWb2j5hfrXqN1cXMA6CFnXww6/AIstAJVA
iZWa6aD4Y+WExhgcb/G7gqdodbVY35JHYxi32/JHliYOUO/UsXN0AgP/XDjws8Nj
WVOumDJIfz0NlBJvMS5i9mwMxc0vMmmgj7IO3XU0wYlZpNLhGM/LvpF6GDUinbYw
bt3mCd+2ljmZ+KEHwWSBx3l1HcjCGbiUyPWH6XtWuqHeMJ66GsoNxJwFClQfgbIB
xNd21sLgrCfrOkLkc6TBe7PhHAWL7vPUjybSvbocaP84QO0zeFWpdT945qM9Mnln
tIIhOBoFpqztjyaFNisjP9ERPRhhP4wpkmBXVHT5DCLYYqhjKWu0NmEW2HRsDfLx
qWYy8m4PCpcWNHAWx6d51oHSvo8QyWMxrApgfNE1gMVhw5Jx9xBTgZwKRsMT5usK
oVuPkHpxBuPU5LNjev0OBv2qIaLcpILzEwwcF5MreFUOYLjxmUiCPO9knPtSUbIx
sbOBoDqMXD4VTAHX6+IhxSupBE+kUs7mJh4ifiD9ARQI5tGEXy1vsgKgZ7hhgyoy
7aNXotlxQ6WFlnrrJwkyjjC317Re17fakZyBc70sH9ecz1PPDUKljF+cWKTgpZlr
abOckMn1RNoW0uxH1GhUF04kiqcH/1H2aN6KtJpAEm5cknSkblF4971KFIBssPOH
Joa3vKQYELmY4yk0HkS1LUFRpc4PLDfHqzxtyMWuH8y0rRMaCJKqkmIZE0BloX+T
89xh523t2/Li7ra6AL5DwQaFPOeTqHebzKf1GJWuEAYo8XSqigICbfjP6M7vUjgv
FezzXI5OWc5WpyJzzKTAgpiTlVtJ52AWLV5f/Vbcjwibo2XaWNrYt6b2MDgEwkb9
7suOFQ1TarM4gk5hGBQK6RtS9AtqDgbEjp4G9y7JhrlpwEgpefXAvSBbGhRPlXox
N8y/tgriG+p9ZeewV+zt5Okc69wRuRrWhF5Jwpw72xsizKWuwsOtWV8KMQtOBZxW
bUpXgiP3ZBYBSLDXnvMp+Vdi9PM8YpH1xoYdextwrmklaFsCHoAf0EiSqhTJNXWc
tbqR8ayHVV/Atisx1TFv4vJ6m5X3SKEQyFy9RifUt2SsUPFoHO8Gg/+yy1fSner9
ciSec8fByBeuECJmPgPe8+mWU6TO0mHzEu9DQe3YpEVOcyC9f9WzcxJz5NbFCbJ0
kmHaVTLRr/fiSw+Nnj8TXXuF25Vak8PENdnvvrDf/5vEPjyzm8jQOv96kNJQsDeA
mOdIFuEayAxD7j8F+VUvhPgVqA2QM4sJhAqbXnOpM4fHjYuTJNHRV4CRfKYarg44
rM5pqRI9AvvNoLrZvJ4EXF4X2w+0DtEvdk152wIgA7CuPbrmV/kG/+HFsTWrGsYD
/HOZThJ3hTatXrUHl719OfEhedJTlpopq6MykUYE3RMsp8Aq+g/mqHlrISC3bu7C
fGcrVMertoPPaX0iiQlTDCFukhxJzfC8KKWyqk6ieFCO+f4cH7YVtawfzdvavOuG
2r2QWpStdeXJxcVp3bEDh2obwRAikUklGC0hb1EMw2YiWBmC0RTsS/YtLs5ro1Nk
a//4LKWVOjpet6MTcmFm3yDIV9yL15BMvCTwsRclTLx91+0n1HUuz2mY0Ve1ElaL
jbIbyNx3mHGaIIm5stEQm9bndPMYSIVm9WZx96/EgynI1n1UssgwMAFhD9DMtJvn
7Gfp9qLM8C/+iZ1qhq7BDhcRYjBeANtzfZCtD2OLsvrOdZNqvUA4Zxn9GPh9fpFB
dC5mM42cYUVqKbScDkalpaIqehUtll/Ailztu3BM1nLWuuWL7BVKguA5P2PLNrca
S4mQPR/gps4SJhUULw2V3dJZCwkl8l4+cLSBJ7MHonMMkLVyIAmfCFFdXGQKu8JV
kY2OIen99M/f33jrmhXqtDpRrG0zU+bKW3qrG+iCWRz1FH+YxGG98rjswnRDW2d2
+6J7Vt0dlyfUlLjKVxDyA3kBfQUPDj4BA8kWs8o+jc4nl7b+yW/mgdVZ/NjqwtYa
FQp2+4jhqlqfIzePz95o7YeQbrmXCJVzplQakPEU2WJU5w2b/R1MP2+lsv3pp8Nf
5M46IxTOxv1pSASKsqlHWkfLTdSyyZZpCDoXKWD7jIg1mD47QW+SUsS0r5EavJNQ
7MU7LQrVyCHumoKcqICERyiDjI595q5kYovDdj8FTl9yMsVEpQLklgETKpHZ2RQO
TzR1QdgYn/OrM61Hb6m2+V20wAIhQjw7+1tAApOyRYnUQtf7GO+hJmev5b0RrVR3
aagS/xkbwiKGHnUPdnALLDNG4WGbr0jgp9htslz8VrrZMEIXv2EYt7D4oHepf1j4
dtPfgmBp8NsxBf7ZrEfZxdYv5Wnb1iSlTBs9WHwTgxvLdbksA2V6lCGfFo7XyhYp
saHub9B8f9PrnD4g1+H1VoAwsvfMYgO4VayEwWD2wFMp9lWrGianBZ8qXPoth3Q9
9+nbsGnhrBerIrXLSRTTYuEiwFJGhvUbJ5+rMxYVam4NEcsWRZ/HIjBntZ9S/Gs5
ACMcAuSnKPOtxrjPlDvYUlMWFhPFlMpZPZ9GA/RkHNq8ZN0Vzz7chaosCaIriYo+
7uERtU/O5LsCtWjESTGf0tsr0/kuV8k+ltx4LJ7Kjm4CqFoukdf8hcPjuO5iwYow
vDlaoOKWtb6HczXNeWBdRoSTSI6IdiL7c6UhStjyhDaq4zdMAAQTq+6dRBGEJeW7
PN5YiioaVqAhGkvm5LHKvf9dPhavZQFQKA7F8cWf+bpoyTqTXAppT2kJftAy6dRZ
f+J1mcazF2VPGXZc++gFwS6bh2FQhxEC4e1t/GwwCswOD/nneoiPd+0fId98Bcgd
QwDo3XVIm0cWsbErKpcm0JvA+IoBuVfls21EHQVQr4ae2yOPqgHrQ6HcrdRXQRF1
/mC7D+cdNAuOf7qZEZ+r+9DAyvlPxGVg6WJWHYYIJKWGdCJBHOW+QBUX52n/tm0m
P5RD3+15j6TBafMbtqGZKbvuXU9GSPqzRqpOEhALQjL7YPFPPRqj/LZdEY+6ihGK
KCXwCyO//yixPyKjwngFYWg1dzkjpRItvvkWileHrMO09yCSJuz9vMoiUQvbcqLM
EHNlx6yVMZbZOxim6TlhuMqC5zghx/vYlD9PXoT97AA4eEJJ4G/eXtLv6zahP/+5
L5y3d0zz30V0vkf1pWedJBqhTQPEjfrUBX72zgQQ8tQp7gXpp6yNNgNcFZ2xYa7u
6HzvMuVbY7IyF38BNC7qqZy9bsqC8Yfk7jCoFpHnRC68mLmDLhTd7OB6w7SJQVDG
DYeH/Jf6tDRBl6nCvBMv6Wv5vaova7SAxF+pk/9RYhW36AYf4nDbCV4xlbm6BGsa
cVPaXYYCxVWoyvH6hiSAM8aBEgh89UtPz1s69x7dLGyxp2vWc5H6GhgZkGeFzWIk
LnKp4o/BcP4FCocTQDei3XPivqbnz2ZRjeCX321K7OVhwlF3nTfpbN15ASW/cKe8
lShVVL7fK3so2BNMF/cdDg6a4eIJazrzJzw6tioWSFTPLYUlfWR8cLwvSSp5R8IT
hFaSuXtvSZqxuxfqFA7ef+JYUtbiQxA1DSD9y4L5pydDsLsYhyBwceDvL/izAJiZ
/HIOXJFDuUq+HaTkFNVBLjUOpGtWcz+u28ZJfk+ZffnbTULZwaQGVxXTW8e5muEt
deEylWhMwT8NmjvECcfEwLpVnAXru1z0Rfexs1ENiSnRpQQNKiqkqfUXogZDqNEl
Nw+kCaVHJrqFpHRhFRck0Hgjb7Kk0oC+79Bz7LYVscJDAoDfs88qvYzgd0uvVUg+
8cuodAjgjP1naucMtcMymkUe0XkalteF6dsmk1dlDq5bV2+enVmT97VyIkSfK783
TdCdS/LiNeikBtGBJ3xJCLSDdrFar+6kech7vgO5HX5022L0NRHH3hGqP49tBfuL
EAbqbcKaQdlwnSY8qO93Bs85uqnbw+76Imn/cszJX+9n3YFA659cdAiobw5cafBa
pHlL701ejI/Z3RzY1GCbPB+BPBnnVIjE7RgF0fiRvGs2y4aoF3xHbvhRc0zVshVo
4VuEJlQnDxln7GeeGnZupi86Gl2mMGio9HF7y70lCjpzaswM0lxajOvvg04WUTob
lTdopYGUBEHpcmboVqhanTvOTXy8fq3qYH0eFWZGcGNpAkyv/6Xk4Yabhxacex/c
T9gpCAnqUAhYD9LTDKoTxeAzu7P1Dw7o5l4RVXqAx1s5E8AfjWixyV8AeBoLtJJK
WgcGNjh6vDhlVyhj9VpFPRTBWRLT9O2CYIkaGmZ4D71qejIEHTyFQJw1M0K1Wwgi
Ti7X6qfGnXsv5q4HhZrlfqTFePJ29CQsotJEMLfMStH0QQLXRnRiYQxuQl3TgPoR
exmGuUZKlWK6oaLJddhHRSkltta6PXTZKuBb25xAEmAAD5jlXmYi0N/VZrfEpkHt
QKmpqEmaOPsQrHtGrWDe7h/KXIPxElSTD88cjeY2nNugbGC3SG0yi8tIHanRnG+Z
AELHxB2jSpUOsfo80H/DFbbwds0MWAheVgwgll8Q5qdwTOfY+j+AHha0VknPAz18
Ip9rhbAKxdCPjdGTKriC8TJ8E9O9Qg4v29otWumLfgAShUGYppCWGISqFiKkXJHc
L2wDFfhShyE4hZLO/eKYa3AMk9ZKXD3HU4t/9591DI0dYCQeT7ArGnyRFFyamNZc
i2pbzYZC23X4sBaXwf9QrKb5guQ3v/t4jvuRVYyyHKtkgfG4OpNHl7VHT5xSxCa4
qMLMq+HIZAK5LKjIqbD7mMdcgCfphnLL/56efWyr8Ir37rwN6A+NguZs9YP7RA/j
3f1MCYhPNINnwwFBMXYhCy7GTerIlE2FC+nQoKg2dx1Cn3CU9KyMvzWI3kowySHs
Cdy/gg9lIWunYP30U4Zjtrv6kxFOzw0VIcytSlN2+Nnrrre5h73QJDVC/DDOoJ9o
HVxAbhwi/mPgG4UskShEGUf+2uPqwrj5To4EGX8opu3JceWcN60elqokLEz8e4/2
drV4dbu8bavaiiCrWvBKXeyPbxrxwbC3VvgtCb7OLjTWVViG2s28Rr5ZZc9TgZIS
ljh+eMJoPenEUaMxMXGVLIry9oF0QsIWh6EgXWjNHrQo7oq+NhQvCEI9lnadEQ6S
ifa4daZae7UgTYkvHQrq1YiYECln/WSZ/tqOU1vZZICeoHlnHwNS0PgBpnc3+N41
jEgcUrtuyDHNf78KKukhurfMhpDbQsr6rXvy20MLeBZy/s8t7y+fLVtaj3AY/SQ2
wTDUs661yQAAS5IDitpNVhNU2F9tFMTJuqunoIE58CDGLvyATO6z0NoMQKcO+D7V
vxA15FuH5Qqhq0MIy1+th26RZzqe4RnHKarBiHEPieYYoGW4L0we77B2tdHYcwR3
iTuTu+jk9A/SnrFg1q1TklKJIYi3DJiXguPDCRn5I2FnFIKKuOgA45Yo/r+TgyNE
DJfQ3D63lqZyCLV5ufZD2JN9cymg9+GOrNeWfx2KtnljwjWdwvWCBLyPKJTSada7
myAS87ffxGqdci+ITun6rdSdQmm7rpqcMi0rbhmyYWjiEYukSx3/qxMhIZ3ERUPp
wgRVmIi+zdzvfaBLKzRqemnTFDhw/5QLFdbdiUySdSXa5wmrjo+CQT8VgQ0MVaRH
P894hYBEptt/8plpuQfi96nB1XVZ7Of+f5dS0ar3pjKiAOiC98BWjFBPsz27DtTU
74ORQ1oUQWlcWZa0HqTpcygVSs+WHTm7DxzX09kbokNsnShTL17KbXthXq07pdeL
mUKytnqFalm6+Bxl1Oubs8jCgHD9c3aO4vqPY3Iyefx5W0joMYGVfr5JBdFO1LEu
zjdEttI70IheGhX80G43yegyRENg4P/2xb6abOjPn9sSpyzsqYygQFiMRHnkqN8m
SaTNxIaJt6L6Cx/wqmB60KWOI57M7FE8cNapyuRmCoKWZjlAM9tApcM+o0PPZlUp
vFuGrnKEi/KdtnHfkl3TOniYx77FBpKjFvLxhmAEh1Zyh9622VLzlVFxxVYMaQIb
EFrTqmHJJ5HmYNrryXVvJBDWvUMQrxqe0P+EApvTnXhGDbyX8RI4EeioKybxymmx
KMkQrp+k++A0ctK/Z8ENeWPAArOrTuU9jBJo8+rkPbtx6Fxcbwe9EZTZgm8R9w3K
28k+wN1JI2bxFSOZwYajHjaVzEVr1WBMi0nu2V/3JL5k95lyzh/vdAkd/qhJl+w5
lCyhYd295TssWBNYTDZ9dDFedH89xS2zrCt8IpPvZ909EST4BK7VJxhiYgwCkWFu
PQwf+fulB7NlQXmM5jwR37lRK0C+TiXPgIg+WOeP3TV1toO8xqdHD3xAgUT+HRW+
gYyNsNtOrEB/u2R0Kf3REaCWjnTSOr0RkkvuV6//+GV+6hvAwyTTbuYNJq6RpfwM
I8qqWW+rmVfwGHUtXcERMFWZnRZmdL7GyjxHygGbdmkGR5AAi3XibmTsjp14anm8
QbT8kkE7Bp2qa+Hz2DE2NjFADnky1SV2qbGagOj9xCNUCtkJskusEeuCaX0aH1Xi
m3T5NxSqhEIeydrhDpRmfcDWVqpEwRNd2C47D4prvlmakqgpNixRVbMQEvrCAIkp
HOkwzHJecKw8ES9K+msig8s4aZOAHaAG6VjIV7VKwfHLr9S2ZWeDnpzm/0VARViV
8yWlhzV/ZPlpTcAA5aYB1ZV7hz3VyLfHgb2QdBDREYaHit/gQoC4PzOs6R7rJMRB
qCDZiDdg0WEEv/cWcLSXNOoodzrhF4tksCkfyGYLOvl6NT4fgnJNsSvQX9JNlWzo
Vj9GCAKunx4lz7QoEAjghrkTy9jTD2ZDsQKDVFL9Wla5EhB1RGyhuuVv55b5In3c
geGA3itlMzTK9NlVtSn0bVlKn4UXhaQxyag9RWP3Tdl05DOvG6AOczyfdVMSUCHz
qQtgsBLiFVgWkUGxprmP0cozyhbxJ/RiVEovJi+/RmYik3QRpfWlkD2i88Vz+GbM
TKOTNbCvZoZ/+v8nj5cnAw6c7h9pVEmV+nOPaOPZKJOA7uKAibc55ckqMec6y2mU
iVoNQl9CC78E+uI7hmlCWxEd+ueLTed1klny+XYzHLcorQv5o1nFhafeQU3aWV61
bE6Hj8cxSw8wzeUrDHdGxl7TdB5zCv9rGk0upCg0mmTIAfIPFDqsEQRaNXTkIyla
8gIq5WRcq7LCDTWK+qf1PT0k9fkImFgKTvdVKQ5XDXlDiLMqh62Nx0w3krvs9NUI
EkZKsXSF/ryQBhs1fAQXo8qPoWxb77a8dONe7ZCap5KLMW12jngMnS8wYBT5AfO1
kGi+sxaznKynqK6b89RtKwXQnPLH6Nyk9FGLo0m5fyLBxf80Df4/Ds0bUS3QL9LC
vLBerOUPyz/OtIWBfCA94deWW+n2P8tujeE3QQXTIl0yhsuxYH2C2OXwQd8ejCbb
QDi20DchLGdAtedJABgiIboSRRmUb/XWkACtEjVL9hQfmejxhIlV0riqTCCOX7X8
QfSj2LCb1KxgojOaEiU/Dp0JV2T+gPZ1uhMDmVWA4bnEbqDQapGVDURUaSakYxql
Kuvfu+0TFNjPwuNZwdYYRgPzKhIHS3I+wclSARpTGN58mV1VMhFShh7/B2hcomN9
bcGPQFU+oVRtBobH5DGsRMyoyOY85gBlh6PYXYNifNc+D5/Cay72mwlWkFx6q2Ej
j4xDokntvFCTdjvogfHNKq9zqURIxY1FEFygDumCI1ZOocU+932Al/5IvVgpORCJ
qBEB4+YX4OiMeZYAFJxSIjHlS72FfrJ0b6hQx3apAHKr3NIordMpC18ws22UudTz
w2ryuZIW07yYlZFz7zllbD6ogi2tGxUxdy2bC0zORY9SAGEX/fxecEdFjtjQibzh
93zS4xKjNXlxWh3v8qMMQPZvY6nZjbcBHRFYsPep5Vdq4rkrDfDyD5MvNCEVv/XU
dRcbe+Tm4cMnXnlNUlCGuug0q/oyG6KOplCR7au63nmH55TDPPCTI481wOfnM/N2
/HJ5/EGpO4JaZnRNIyguUMDSm/AV6yyCcPa9wF7zIPMA5fdK3SJj5St5viWAQRvY
bH6nHRNd1mVRapcAzw5vldqV70QaAelDFjStBraMcLPJkzg/iQG/hge0+4em6HxZ
m/5bHlTDCRZ6423slfTaNRcnGRirCEib2kRMkOTa0OtvGiTp679HoOvXd3KbrFcv
SZf9ocHlv+2iBOE+C8Mp8K0PrcnqS6RreHekm/5t0hZlW1+H6ZHqAsCfAZOSLfiN
rtB66PrFG5wixRs0vCKhQZMPdlEqT2qLmJ8ptoUKzGRaZ6ZT/3j7+BZME3iSYeiH
pDDg98Y3nHzGzcvUnQAvKve60aemHUIvTQhtzeFEN6+R0QmMNoQ1AYXdl0U6zrxp
ADWiHqQFeDiQpr8WFRpBEJU4isMJXY2hh8BTKIX5fXz7wx/LLs2NIBjXggaFuiSQ
Zy2Fi1Q6HaJqCo4IMi8rw+DSvySGrb6EERJzfOA5NZ8SZapB1rCjX1DgMajUfvXQ
YjdITL2iPdYy1r0g2PkVfFihv7pZ+tOfacwGTw/gxMwqMWBgeFBpQyzetqCHelZE
b75t4n/1vkN/gldyC8gqzO424TraXpsXtiCTFevPVdERNR6YqsBGNYGYzbYxwMPG
GJfejMZL+pjyoCtVBWV3rmQyh+WGOx4CdjVkMmGRvgl0F/6qtgyDw8SWHsSmVoaQ
oOr8SLIKGW7khR+bVBNHVFFga5Up/TID3ifzk6npmt3eZNPLLDCOkJNQ7qCNNQxx
0MHVYUejYGGLfxQQaOmA44Lud+M+joQbPJOsWpnh6i/ADgl1PRRbJ0/dD1b06t7H
fm2P5F+zDHC/huYxhLB8gYKqV2wGd3Ph0JOtmxBRlXl2Y6fatJCCD0tCJUcOupec
44mKW7cX4vPi2kQjvYjPvA8PKem+h370xIuHwx9pPMSI8EM2dHOO8LOkz2knFJk+
flbRpfiq8tVaXRG6zlcf4g6kvucEcPopOf2gsLzXZ+OosYWIrt0WUXwUlFslqIyF
eiq26WV6LFrTohGZQWNQ2SpTTI0lgAgD09lVHff1/StVhi23AcLjuXSIS+kiaDkQ
dE4BvqwlIOosrmTKMnxxlninZo5ol9JSbgZpt6XGHhCbzyMe+5WvwqyIjvd6JwH8
z/51DVK5nrS17yk67o96Inj0xrl16OkKe8wXLiGkFzEQJkQM2JU3evTIHTEj9BV3
xs2T8Jxocc14jbPi5PzSK8p4tsNwPaO+4Y5JdC2U0NwaS+ysBRpJdcas6Ip2w7Ih
D43yEpcwUXml637tFMhz6j7kSQ8IUPou8BmtWZaEkXu/AXUMdD5gX7/X6wOLXCh+
JOpKee591fu7oD4HO49Zb2UnLOgksGcVO7gCjOGo7fYY2A19tPoWunzno4uK0dCa
/fJM0EtVYwSGrVm9oyI5UjhlMPRe/CZeE6jSrDYMUMl4q1oXPu78MdGKndi6qEyl
pCQRErzcEWdt5stfR8uU66N3lGErrJ/OIMC7UTOYtXUFv6uP1FUATqHtNwZ6akCN
vUwtUO5nVXK+UlDSB0XfXS1LVK2lJZsyTDL9GaMajF16luj5CG8888pj+W3+jroI
rPua6vTTcxbDxLvivMHn7bHZWrkshM3oaIgRz+fdAwGm6L/EyucMb3vno6J5eWoO
TeoSkhLvJF2KYWlBPSg1jkQgrH06HHqW2fLs/uhzc8sWGMfOcPykH7bXti9Gww4V
Pvx2RR31MHzULB0eIO6hox8KxHFt5gjWqQTnjahGexe8xSogJE60F2c8WJaiv9VB
IlIw53fJHfZeqjJa8VKVtfhZizB0MhYpkVvrIk7YvAIfRY9aQ0fdZ53Wjjw6Ol6L
tMMZxeME+DyUgV1oGkaoKeqSojJFvqBR7cx/ZyXhyhaPQQfJkgNQ9rerXHQrIuhd
pu51YUK/k1tM/An46tw0TUITgXAFzZSM+Ej7VOVbCC4X1Nb+WVk3tSH0IZqcjQWb
fKfAXmuZHA8al4zKyAVIj93moDOI6yHc6DtKAFQ1t5CI4A4aWkLdt52ShOyhppO7
tYMyX3nIz6s8PENHd0ZBuZLp4ezKNM0wb/RgiKo0cHFPruB/f97gshuq1fEc8pMh
0B1SBLF6fCYhMBGsIpbz49PQdnObt6t2e9FxEU3bE7+UGoY0Lb7z3dBZr3w/BeYD
Xdx0p/Gnysf6Bwf9rlCpLKhAk2QKyIO4/uzdfONvb+DCVgvr3JxDzGLKFy/OMlkl
ngkjaFwbEFfNHM8OHXOr9ncURYhZzMkQPVUAJvtnC9iLNAm3T0NTPmTvx015lDI7
Wb9KorNxBSV48UPxkCAqY0Gfb3w91aMtvCiI9dsybT4Yt6D3ZrgB/VTZiFS5fP1x
V5PLFkYazTRh1sCUE983mCp0fpSn77b3X1oDzhIZ/EhGr/3BKb24UEup/CRrN5Wp
Fx3eGTUfB0ofEtAFfIBhwCdT430uetqmWIzro7cCYqaPpfOSIc63HJzAYBWxa6J7
NDeEkMAOwm57J7pzhwZ9auzkHisH4mgtkVIiniyAyIlotm2c9ssuFdUwuvjKhwjZ
TQC7T+bhjZ7Tc2b9iOCf8N0AaqS2pIvIULuR3236jz0Jb6MlQXmXU1vpLz3I8huA
xy134I+nk4kNT19LZUnVox88eI/LVXP1MxAQSlwaezF3M41b4yB9bHlGqo9oxW1v
W4YdTRpYtNOv74itig4Zva4TvStrL8xhqsdTBhsKdtgnSVqx1uGqdMgoQiLT1Roe
8FKGAmk/fCSqCj8B0xmagXHubK+kQpWwggqv4EjfyWsXKfVc93Hjr9+sycYTmDB/
Z2iFU334SDg4iMqIVBTzFj4/n4I8j2U3x7rE69Jn7HLmEiEv5MPXgQCMZtdFnS/G
ItXDArHHGAwN9i3N30xm2uHhVzKH6+NKdchetQhNGVav0X5n7JawRyfQPRoXNazq
MdSwJgkPvInlEjEcjHc+BXYH8jD6RswsqAunr7v2LYs/TTbK1bnr4wtrvAciB9BK
VnmiQtA2OUULeqem/LsEXzk9tHM+PyorZX186x7AOg0mN1PQusJMdJYAHbMHSvsy
SvKx8f46zgo8v7CUZP7hW4nM4kf4GH1d+XhTN8OY1pJSia2equqxTIIbE4lfwumZ
bHf3A40Et4TlO8M5Cbc8aYRhhG3y0PKKF+LxWsCJWVyf3rTVcjZBC8SO+KzLpT8T
8LMYMWUns5tWYUN+AUoHqLupe2VQojDKvvLSAUMFBRl2spT+0Be6GZb8E1rPoc8G
Lfomf/SOnTMyi/6/PQ4Z9fvDiHIIVZZermSojFHX6peGsMfzgHal9vUqTBfM4gQl
4N0Ad3wYYO4D8l0Xv2zjLLr6M2A7qnOu6jTJbCE7Zj9GIvIWgZZ/sguV+3q/fYh+
eIE0zTzUGFZeZu9Np/OC7JULclpgNu+oJm/NUtjiE1SvinlCWGXfKzr3dVk2zOmc
xGpdMHMMrWzJ/AkCoIxKqQdeElK8zrBt54zB8FqfwsiF8Yh5dW6c4mNC98tpW2Km
bQZrZXFX0tSjmAvuU2fpxNcxhGve7Gg6N9LewD/XbnIDmGDA7gR4YOhA6M50PVpY
pS680Yg6Ak43eHHj30Sy8IAmA+x+u8oRHtYeypVbdMygFP8ZC4ckkYM2ZvFy5BY1
lcGgP8dUyGjTeSdZ0ILJUs1c/QbXBPFWjVAiRG0rk8b3DqYh+NmGgHxAypwaJBa6
W/rM0gijHnrT/gPmQpdzHZ7Y4p5/VAPhqjRIUOLeuFT0hMjXdqRfNV+P4qhgzYQP
Q8WN8nfkDLJPAPSHHjBMKRVL6S5xx7fL5s7tM2y+G+bl8zxg7Mj1ehwUDQ0oglVs
eT0c959/OiVTvQXqqEUwRog7JFaYQmuzbRb2IXCxcr3HPNFcN9xr4OebUMhR8OGB
EC7LX9yUohiHrz5DneQI5AtOXsaFpFksyx04Yd28jdd9uuTeDsThlrYmDQNGKp1d
jPqNx/j3epsJ/SWLmxgEBqn7kSjDBG/tnnUwaNTQS9iflvReCLXYV1bt791B7oVl
GnWHixeD1CJFzsVN60Em1UccauZH2h4YDV9wrEnGjDQ6uC/lZqqd5ZTwt+dXeFvg
w7knFD/nCmhOkp5tIZ42neR8RADYzwYDhq1hBDDLQ19sXWIuig9GN80YnpAZCu6G
U8CPMDOOBc8bEHD2e0ng+SO21Tj10zD74UzRxYjoXZtbRgtD5IfjTUKl9eUt58mE
LQd6WEMRjNTYv76u571kWjli1ZliL39vJL6ciwQgY6OHxOROQ/7TCK8gXgT2uFMU
Zg6CRpZV9BZCJcNRVInWg7eikx4Cs8/PRQsFHbLOaI3h89HqdQ24z2wtVy+oODYd
6q/4qWvPJZyd4bugUHLeXCI9oizmr4qokOEY9kulaORCAMkkTxMc7W944al/obLz
OrRmh250GlM1ZbJSo5xOfvLb6douu5bPMKtPmwQOvGSOGAlvMQLJe5/yqdSXZnWG
sHhUIlGPTq25TtsygfgD0nx2ikQDA5MlnJik+gQCPUn+89fjkshdqHhDVJhFxoQ+
rpKgKWam7wYKEZxL2bP20ztUEtqUl+6f5Ygq3R4AnbivfzAHei3qjQrY5eI8QImo
Rz2n0fdXlZH9svz08qdz91f70PTwvyPX2qH+JzbU5ZElq2yVHZCXEuqZUWMHoh34
ofC+2AvCgbbf4eCRNkbwwzTTLK8QaNpaoTJ7gWZwU8ydsVNEbdAO2YB3XLIWvUKA
xdjWRtHR2ySiQUAKgIO2pBB0SaXHNiD1QVOxm2EbxqKe82R2CVCWUmqP4rkWc8c4
zWItgYKoTM8bxlK73NaDBEInqKOInVUvbx0wQVA+MGqhtqPfEF1tzmSuMXSNFwFg
04Ab8kFOyQTiHsOqsXwmGBy+N7NSIM7oCkfBt7uWfOPx8VAoSXWQfq1KcS+/L7Ni
mpxboe9f9HXF1AkfSRXxBAfzCHUZPUrhrIrVv4wy6AdCaYlgBMQ73Y1v7iKi+2eZ
yARiUtIs38uvJSFJIbURAtZCdlnIBTqt6bTVP5nOoZ+i+pyz5C9Rlt8R6kufR88a
2Ie9sFhnklTwby1RGpxrrPtfDjkA+mgTiKOH9Y9qcoskDR9wh7uXOn6w/S1km+rB
s96eiYctBNB8beGZvZRHAtfuLgA8q0bqASPUicoaK6nm3vLVFTNrFyXBRkKJTtkA
p/i+5S+Dzj7+gNDWQuyJb8m56177+59HJDPF98IXt6WXXJomH7ZZ6i8bMLJMhb8Q
hrO824ZsPU0CePPojWtqchyIidWcW+rCAAsHs+3HhKoFrNiZBjGuU6OV7kn9y813
8lhj+IdXibwIvUzYwt5AE2MrM+n2M1tAsmFJkx3sRLY/2y+gpKT5Ve4Y4i/eyO3f
K8RQ2vtAZvhCHblZ1Eeal0NwUjbvKcuUlo3DRRVnNFGdeeAgWtX/1CPtW4kFkT8E
QhJKRBeKzWkCpBe4NRl6t5IXj2yHmoq0i8iIBhvYu2R7Yjv1Kt4pOPF2FNMQoiAo
Y9k5OeLs8bU0JoLFkInZOGFEMvQQudZF/Kp69ju9K4A7Xaxefr1uwt6jVF+EM8H8
UjHJdXgCwUj+4OZRfoQqKuflN2uq5SXLzRYxsjbLHsWJlmOcorZXTydFBQT9G/Z4
3bcYd1+qUGGiyYDe40JRrFqPd88qj7x2GPtDCzncWRdNNP8i5PvafoxVJakVReNn
yr7EKYpHfEdWb41K/dznLi5AvBMHj1A9o/Bdo/YxzNNcZT+6Az6jImvGDuvE8WWZ
2W953P33FFIiLEnkOyUrTtgPlWMdGMSVpqjAD0Pij3y4OaGukAbinvQzbfcxJ93v
zEE9t1ntuTt2ubEDzv6tODwtX0HwYoB0uFiecIZqeJ2apKBut2Lj3kT/gElAAFBB
tid869iQBEzXs6lE8WA1zt2GZjHynmFYwlxsTE0Y4hsfZ06uHyn8B3fwc5tClvPl
ZaRnL/zCGrCsn+sDy84ftOvwPV5yCGGIQCoy/LsqTY8ePwyW4oL8xKpNLVczUkc3
x24hA6j0BKJshAVWEdq6s75UDu+OUcgnwPSsfW6ITSXwZZJj6drf2Aea67TaxZ9l
JldgTBlytpf6EEMcwsjZJf/4ICZreB5hsjPpgBzF2DENIEnXS6cdjxMvydQ+y9hu
jrqqUYYZd2tGtGEA88IF4fDS/E0Z3suLubD0ThadUt1JEFW+cZuXB5RsVzMFQ4VB
/eID5kvZPcyNiBwKCaF/tQf5VIbMwbePHT92H19eSRJWt875/z5x+GVaTwpuoxKw
HnmQJt/GV8LnjG9i6olRcs8mFs2RL2dJSa/UULa7aEH1gAHXkMH46Z9c3x/n63LZ
RRC4o7r2eWRgSaSE4RWSWBVZVaETYfTz0OZji0X0PgKpjeHKKDdiV7GbQ6Dfws7J
Y7AuDKWQojFsBStJOJ/8Eg0xmiLNeWhjRlN7Jo3CENqZi5L/Z5Yj9OuhTnyr8H4y
I7i8AqMocxYaVMXDNFdpzTFmBIULMJYd11EbKRA6kj/chl4veB3LGrnafBMD5c7K
9oFuIO0GzfVAmWXovfiFvCXFp8AloMp+E7W+iG6IXkTJzwP46sxGQ5SIRjBrVfjn
qErFkYBucnrCfx231ROTGDTSnfK3Eb6uG9MXZ8Z/KWrHU3DZMmQMy12HSuzDwi0F
35+pE4eE+VZxwigUSFdi3v7FkwHu8MPPr/w+TNfR28gQ2NN55osQm9/0u3Mp8Xjk
KKE3eUK4mF37hANQ+CQ4y+UwEvjq7Z1+K7j52PoJPPOii56HNGAG6BJlN2N+SkQ2
IizZHsFGKPx7YfthCj5SwgXJyACIuPHKtbYuQKfSogVN/hv32tjB3iveBHlz01Hq
bo89U+xOxm1aK8SdnNtcDmnBP7JATzscuahDoXOxQ3uy0JNZqEo5WMxWLYuKUybl
nM5pmQ6l9XwcZ5oq+orwWX7rOZr8pEz4Aw08BF4oB8rzjWx9f0UCIJn9vCA8D+lX
EAXgDvuwvUljE0ReTXkY3JpuZw0Ej15SzIzuC53cnZ5RUHriCX8tftYI6O/i6niU
hxLpFwXXg1tEkhWSOy8CeqbQKRSS+qS+ItAQTyhOIsamwdhGTdB06KO/C2IvWhkG
GqLr/gILnZswz3ToCGw9NpGRfhx+HDx8VyfkydVGbKPLLMpZOAbfShEDWoTmtwFW
QrO2+7iwXK9Y65T5FHwre8zHSatmCjwKejp6lM+Gq164WLCyv2sdTerIs6uKfhYQ
Pf7v8PrHzEv1uZPguzJWHCD+MAmSjydl9MryhnnVelKBlCQCYwjVh1EpkGoKjtLe
W+Iikpk/L4/L6HmMKxpH456fkL6hhb8kLcrNLxU2aABO0snLB88jjYyJnm9A4ynV
toC1JZvQ5BWkZ2/ZeOZkEVgSGqwomQUuHg8QPfh8l+jNtpm9+vUiB6POOxgzYUHG
diu5PZhzsjWsrvKGQ+5XSWVPsZIfKNhJlojGSZBNSh6v+NUrDeuTHGCUFg4Pb1bj
8L0B8XEAl1GxmjxvYbIVd4o/Od0hy6I7+YIBUydVvDpJ58/vXFd4fCt4zxnAYxyl
QukiDYe25Vd2B/Pxle00x4SxP6pIxReNXH/5xYPhecOqbTAOy8kcaHwpjYv682oB
ezmrBPT+nomWkzjlkIg1tcXbL9m0gQfFU0dv5yh4u7RrqfPoM9i+++uTk09MV4Z9
+lQm7H6Ch5jKpmoeG3MvfdWnBp/B11YQUOiM2f4xWeEtY7ZG17vHn0O8XJElRjU9
pSlCKDAr7iugXk9o7ypdiDG4GIo3/wqPeoMF2wWctEw1WO1hr/IpR8je7aJiF2HZ
Lj1DMpRVGZX00fvzjhRx4ZWhlivhKi5gfhR5T31dmgqf7Q/MTUUjd8224rPbjY21
ULfdRxzhWCvGrXTYPI+fS5rkxd1MfSqUUPS7tCuKoJeWBsC4W/lmYqEzpQe7DpxE
CnqT1UNactnSM0oJf5V87Jk0FPKgH2ujL9M718x+wGihjJw+8ibfBHirJynxxdWR
oq+H3u8a/P4z3Ja+VurAVfcZTFU16dwR1TDVeldgFwWqRAOHXbW7+QAVCWGA8kd/
0I4P3ReFey04UbCLbae1hnGMCAXYeWSBVanphYl1cTtiGXniI1qzq4o5aOzsHaRd
sOcOdd7VBA5G4vtA064X2xQm1hx9jD7+OfSO2Tb7haZeLiwVBhgmR8pUZRpsZNPj
mBRkh3i5kFlrtgchAeB9POMbzejYYuA3zyMZNV2ChmzwklpDlbm7DJuh3HiSW+AK
j9Iwc4tLSpPnSBXQHni56faCs+r+CBezSekpfdpQLMa1rdeUejEhMzBa+ciU8qn7
xjvgcQfZ2p4mIzXjWn53iRtk5O413wEN3owYikezONNus0uH8UwluvHTnYMUK/Oh
4hytontp79T0ZiJ40KAd2K4m1tGcRn0myJJCI2rmy5kPuw6wKWnJJdgLJdOxmngx
nrtHBsDbN6sNeTmP468KAfA7HObL2NjqDguaWTx7moogqNQF0XD+Mlwk8msxg85A
33SAhZ7xreSp1cVjgrCndPiLYDxepwMxAamW734uzfMmEElFu9H/41FzC6SVaPRX
rdOj5oSvOResHs94H0DW+dJc4FVAWjqjB8R15oUvkOMOAPo2rTI2h+tujbgZO5Tc
PnFg5bS1B2FkiN5GutJP2Ixl6pGTmP8w51Aq1gd0N6fJIffAdtA2sGTfLK4c/8uZ
9Pc3uTcs73DzdD9qkvNLuqgefTmaoO+WO3ctylqCFGSp9se16XsvkOsemMah4ZB3
RSCFHOKGf22Pv9UJ4Ry/XM3V5kqi9IRh2vRAV3z9apmegso8A8eX798wr23PrBDm
Q9Pti+TA5Orqu1KhfbIcVWO53IC/fCXNyO6xwm8AG1yKXdFjiNILX9+D3CuHu3Il
w6DI2B9et6qHi1FEX3zZ0sQ4RpkP8EuEY0NrR4H0PQe8cGzxtNvqfrKwGns61Y/U
ZFBtxVohFeMSoJSXST2pXr+6FdpMrCiYpr8bVoHWmBrKZDlK8ioOp7ZZF3UR+7ec
iZBbpP05eUbaR/hLbseLqnIGfEnNTy2H4kn92b0GOxCB+x3vvSNjLlICzVbp+mQ4
HIYGbB73/mVw+TozfyoZcgzD973QH4vuMtdyRMaXDDAlV3E+3cHnPkDq+rEFD9p/
rfVSFv2Z/OPQRfsLhxOyq8U0dMbMMeYf1e3hTX1Cg0qusTQRuVtenT6s1fYP8U6O
zsWKEip5bvkdalyLe+LSWgmuLojco+JlElANKVz/8a1+hmiFuJQD0e/aMROh68HY
XeL+se5NSmCDFqRI6VEQT+9wuPXMVWA7mJja3MdzGzumGEDQ2XWFTM+IHqAmBHUg
radxvN0PRPl2yQL4+uA8FrbDOTDbivbp2b2wMW3oqmigW7/x2RqiC5sdBWfeJoJq
8qO0FuoJ+zJkA2/1v1SYdphST9ySjliULsX+O9KH3gF2jSfbpk2lt8VwSPG57R5i
Bc5hQl08n16dINEgE7VXDzai5jk1Lcu8IzpuXtQ4bqy/Huu1qE6k/zliGI5+Skyk
wnJQkuqSVnL6flgxi9ZFqtywOS4x1i79095dFgyZjB0XjS3JH8ixpcDU+bjHhPX0
HlaDCHMqxfh07BybieIzGAvRafXJI/T/NDHkhNT0G11r75ipwqvqrKso5L3+lfgt
XxRiqpDzEZcSI7hFB7lAc5PYbO2igtj1/iI9PQwiET/PyQZ1g7Q7Y2jTkkZoJY9/
yZrfACW4qWhkrvqs14UnNzykM/eW7aAWZNyRDflaS7/5RZGX6RR/b4cK3zuYSk07
BZxrNGhc+6vpvhAk6atDFiN6UjRx89DZDfsZlvDgjjnZtbO75MIEKZd3lqYjcj0w
iPrDQY0y3onr2ZeBuZL+iIdJZ0MuwrZnhSxOTR1A37Fej6eJrjXVrxR9oU9ABoO+
bgPg2OY3vvF4xVlP2pWgNBY8N0gTcbvpU5lRAEApla69YnxW6ZftI9IcrOs523Jl
YRThrYjYQAvFutbfTDFYd5GSLLz67ollHng6i7CE6PIAG7twsnSW7I6GsZ8lK3vF
PmULqxAS90gizpUxNcWY/JoXiMJzPyr5NBPtWNqBD0Lr21T5t7EmPy56FjgzPsVc
6dozdicClaKP6jYoVUPI5B+8bENR676+YdVKpsLcThoYg7zu+OI4/nvkKZ6RdmKC
X8fo4VTUg1ZZWq6Nal9eD7NYneKzHH5jmgnwz+UC0uKeeaMEtOgCPwi0FX2fB4/m
BZCHpesnL1YxVp8v4yFUrKqTACB9KN04Z05z6Iy/GSlPhyqQZXV+uvxDNiW9K0xy
1bUSlERsjmXH064xJTHCJzXdrJEJYU79qPLhEw+KiMTG+Np0v0Tfce9VOkPqqgew
7r+b1IVGCrlRAT/neV9hCQAiFkWYpv5HwOrQ88itPklCAqmuteV20h6U2uad3TEP
mOQVeITV4EoqL+eeVZHAxAQImD/IRAWatWJab4ODAscA4tFhfN30lD0wJ9oKRIiB
kY3ZTqllUkIBz20cdo2QPngBSvUfP51qrALxvIp4R9wTNn//ymYGpRM2XocQMtd+
Iqdp+E69229So4eWp/p5Puvj3K2Q7etMoYTDXljT1KPg+/rZNF1m0dVnXXjbEDgR
0b/tVao3v4KGC5TuTMY54evCJjQfJpjrKQyFOolZedAyPJw5Asu3KvFn3UB42quS
gXbqnXEjyeW3LCcPGZCy/0eIo0sTJXSmffm0VPMNQjEWteHaWaIiJCEg5CtNHHaD
nifJAs6glISi78pGeu7QuGgxXeLg7a+mKHJIKd5CDut4gfpywgZKhryhARjMFd6U
fzLxms8CKp0gb1BntWjpxRfDMDC7rjxDKJh28MIbjAD4uYdTYkx59swWuIowmXZD
5y4B9/KLDof4xS3Erc+XZ7ejhZ7GEggS/E+adboZemTjVGySJe7ZWGaGJce2B809
6ynUag+Ob97swPu5rBsbThJJsTmb0oh3+VpOYUY10dtHxPfc28atxiThFMYBKL/5
RxMGwzzpc1IfsrTTOw7eewFYEs2acgAfEfFUGMS0b6wrfPVjYC/IIe+tzrRiA6bc
II+89eBKknXt+6zbZ8NZChlBBm8MfQdmFOE4rJgP7Ya28ajJkBqRu8l2OS6Itpit
dvG7jT+fFIyB9ZBqZ+oUf81Xg5XHQUJ/EVnaPVEfXb5+Idp3WuZKl+RF54uCrT2l
5QzfZppDz973PiyfRNjONvY2yo7q5DP8Ty9MGgu/7JCTNHvlLLg1qyGGxjUguVVJ
g0YOj+4aVsI6sWhataOhYJI8sp/R9O8T5gx8et3u3eTbTG5iEkk8sp9I6E74hGSI
on7HPdY7ridP9x1/QI4QYMU66ytzYKMLu5TonitilwONq22s0B5FcLsOjYPWKJGI
meAYrad99CaLYac8FXAVVJtoHzqpkbKf2CU5WGJbX266/3duMXISBtgWhLn9iTyX
/5cG7b8iUq1DkmmcdlDieHUHS+Sb0XibVfBFPIQaBhN8kvsVCvKZcDOul+Ituu1b
VscLRr0/SgNkTWPvnZEt/N9h4K9mHHnPggPUurecVjJUq+Am6QakYaZepavpg8+g
WQyn9Z6izK6vyNIj8oAFssm5qhcHwZ1HODSQ/xPVNUr9tsbFVqn+ryoegSw+CF0n
e8CmRX+2YNoIw8rzcNvawqi2ch+k7NQeIl+2gaBORXhpee0vs+BzoO91JFqpcrFN
3Gd6xJXOxVSRUg95TWaU9VY5/OE4upjfTWDyiLAJsT8Nr8AqJL3G8D/YA3UPnEk2
xZr9u31n0rkTlr0dT+tiHo8UiaLv/jzFKls/BBAgTGPkExGv8kE3hQGBs723/Dln
1t6H2akYTjjnEvltEroH8BViDQuco6udk3dLstOKkndk23uz/Gr4k+eY9wbfpAlt
RNQEpdT1fgNM5fuszg5TbBrivcksjybwPmWk1TUCksQAXNlt9NpH83WHMw2w56RP
dMlZSV8VDTOgJSWwzX4IKnHHHY6JTcRwPbK2N/9MrhlE3SlFlwfMYSNTa9htGwEo
O7eiV/Jtjdk/TIhVlSmA91KFVx4UWMjXycde1eLhj9HrfhAyRcpK/fy93LTCcxAK
0QTrUTeKetsR18lh+FkDiSwu14NGf7wA3n2jo4IQLRd9vedte9WRtOmQ3BQu2YHh
GFp3USZNhU7uIVXVe697UiQ4IaMosV4n/vZqYkBiZMbOzl3GxtG2zOLAeMRCxJ3V
PzRRsYlSIL9e9pmXz4gqaiml7+EqKPOeJJX8uids+KhD/9eRKyawbUozoDS7cmyU
Lcx3/Z9IOB0hbDc77oOrgrK2n1VcXW71A6A1dUTNx4tGt+b/U04g9yFRBnQxAtyx
HcRNkdifyKOyO/VQtx7VbGHT/koTmkYv2HrzJhfkE4f3ejSLuTX8HhVE6+sjxVGz
krldYSXSNbaFabcR0e/ag3mm0/sbL/qdNhQznLfOxuCzlu/bZFRQOUy/0+RxP2KK
SwYQsHq+K92NGyFkoaJWki5pFTGaLZ0u74Sv7x+xdALI30MSKIBlGzBe16zx/N/H
gzcylEKTVMVXhP/l4jOfdovDtICWCdyLM3hd/9Dm3m18ifKHraT+SK+qZE3aRwkn
eKvYTbLK1HYcs+nbYnKY5EM5LZ+g1W0nyiS2DN3OgP4Z5lkAIcvF6ipqaRLs304A
XcPFteH6CJmA2a2O06C9q/9AHeBl3rlWSZBrSnGLU3layI5f3gdem7MG1Z/Igq6R
RGR0pLE8e56+fXE7qIIpzCfcefLqYONYAhzmUABL9zeOzcEbsy76Lu7c1TIsQ5J9
YWlAlBnrQ+WX2jj0k7oOy/LiDVbFsINQW/tWf7g6HrFSj6Vgh1OzobgR+awokQQ/
/bsVbUOrcNAI9g9c367a3VL/QiGOAS6ZMc6/ofc26teZxCf4jzLWl4u0TCG6w2oI
IILzpuEUf0cwcKli51WTvearwa4FOHMhIU7utzOXg6HL9CO5jr75AwA+rdLUjgxO
X/XUoaiGzaE23jQ2Zf5DGJGWdPNlrmYNZdr6Aa4w9qZF5vUwqy6Os2GUl+1kmAjt
KjCKiImekG+y5L6JeJxZC08YnBED5nIkjr32faW2TLDnLKG/gY+P58fr31v+HLeh
waEeQV+RvTzy61RXgrK/ucb9/SmFgiuvbOyvW3YNfdCWBc3TY801qBjhTkFeN/yN
yKxo0SZ0neWbV+GGh3HhCLHaMgOY7zYaeYRId2268tLjOMgFr1VfKgi0EIdnd4Jw
0AU5HonLgOVvO4pdRv4yPDWOoSCQTdQKbw8Vn6ddnh/vy30fT7scG5/k02Tiz9K9
jnQhBrfScYLjm8HX7x3buY4d2iX2g9OmsBEGjgCTbarkpMFN9YoEfqYD6b5CLwsw
cukjW7wqlUrQznUALbE+gpkcysIUJ1v+oDwX73x+tCSkocGVUNzLwZfPulspCfTZ
pA2lMeOB+6Bd9pWpu45LeRltHQDRY9s6bAoBdb8YHwAQSUKrR2NfTZ3VnBhWep0p
25JfgwjSlniXSevNq+4068L56mfTkrUnEO9D0bAfp5EsxnMDol7HFo872xgKSHRt
Pahe/q8Ak4GgFHGeNNGZZ9Bn/T9Pfu2LR2wHMVbNRjYpmejZqgESwPtWZlzOYecu
kJW0eRaC24BNMzoHS1lqdipjL9RJ9K2WiLlvts1ExPtN0zb84wv5TQnCx2Gzg8nq
GUJViDe2q7U4Aru715ZdgFRQySTxmoAts70Ql2RWqRg9kR3mEJfLSl3WeMmq9hrj
/OcUq0dVahRm4e7yq59f3fwbuxvDCLH9+L1iUcVmFm1rAAlVei5+4hGqQCPznsEj
xHI8zrCLZxr54eBcY2a/ZnmkHCNsCz/eLZPRUIURRq8R5VkKezXe4KFMruqpZuid
fDcssEaxkA15kztpx2VLu9Bl+vMCywpxfHJ8T+9ydiC3lSGjQF4eFdPPMaNNUbXO
cJeMzQo4S4k4eW3AzYdK8l9vcdiI2gsnkHQvqH+JPWPrkz5zApBcL4FCxT/hhQXT
JMFOZgZDh628rsLtFKRqYb0AGdwSGj/k10GwO9GgZrDCpfyAgpwlXHnvpDdVHRHi
HzpgxydBjUgwcabAzFBf+5TWBhgCaohM+plZA4zdtKXJkX/sKIcOueSmXqBtLaLp
D4kAZ3gtpE7qlMtf0mmOWGYsQjLL3MWznJm5ezc+cI59JwDU3rasL/beLf0038Li
JMkfKOgZPGzRMMy4jfhtmCAiyo7s31EPhZdqVqV+dpj52zetiErJGgLC7lhAbiUp
n5zqcSGjITKgyBY2a9fbtA6XNkLCHv/l20WVB0843J+mpko3pOLGnrbgGZq6EQIS
FzF+tt0WQlRaW0H+E7Lg8auVri4QAfA0Wki//FXZ3WaiUkxuzd/x47rXtt+93zhl
Pjla/keUXCwXeZaDSxazRG2Pv26SGv/AVw4NxATTTW0tPMKJKsY+D75gfkK9H89w
6CeVAAk4WB5D7ZEiaBI0D7hA0g8GS09kt7DC+2XefP9QNF/U9wb3AVF56bLNneZF
jFDj8czS3lCyQDEgdG308sPquDu+viktgsEAOX6G/5JPuBrAxhzL+vqgZ0FJbv5d
zfjzZSLjw5f1YfGbKvcpYPxzS7kuIJaI5/nvfHY3NrHaL/00XPA/xqnhKOOWopie
a3QQft5UIefd4fht9iUL8G/JT+Cc1vw9gQhkDKrn6MnYAAbheumktJzmKYtJYUiA
IUYX4wmWt4KliccHcKRgv1ZEJ0Jh18PhUGTdCd5iRfMrMqpyDKu6vaSAfbGpMOlu
CH6XMcyTUqI4VMMV+txqA/R7B+qREko2B5yzOZ9xc9YOK/B0gv5QsfDDCpNFPIMa
7kz/9JY0fKc3pk5/1vc829Y1FpEzP4wTtWalxSTQiMgJsog6O3Juwt1QGVvgtms3
komzjC+eiP37+o0yG1B8BaScS2sa27pSzyuI7YqD6Y9zUn3DglyjO803PK+Nn+Ib
YJ7P1T4rCLU6w4siZ+9KADQZJ5cc9G+8/8yp+qjBmBY0ElvgbyDueG3KYgrhiXPn
NMUwt5x6UOCMyHBOVk/QHRM8mf03fn57HJ9g/+E0e2cEaxeQBPOWzoCCsk2luBiY
h3Vht93qnWibo1BY8Py5pI1HFqYRGC/cQMjBLPoICfgrbmJ+9LOAbcfObZikUBWP
fXHmHlxE/iYjw2DVVUHSTLBwwTFTiW6UM38cZn6eXMGD2FEGDhvsfVDQf4fh3sMK
O+AKt73ptEPEBt6a8JxHHCJNqS2rnvqE/+IsOWQXLUUGEfwK0DyTgYhuax4gq50z
OqZ9k/T//8LpIjHiYszWX9BGf6xKveHkRncvP0EeIkBrOzzxOiaP2LfblRMb4jXX
4gf/U6ySjwLf4H0UcPyBwvM25ITf9QsP+Ll+lVoZXl5dWtg30Pw27Iq+68etO3M6
jzAtSajRwLObP5urmGPr0SOVhWstaHQB7FlQ+CqYZCkNQ/Y+UO023aikt+PgeJhl
ETR7BzWc/EPoh70E2EeempNVB/bVRAiSz1DR+DI/67hNlaFgIiMHxXelzXFfT1/Y
7tPmDMb5MCd/LaRNBnGoqx2B5TgWYcPpdWx3I16TfhyopalCvNJ4vx+qj8gV9Q29
KpJk3PfQDXL26Ws82EkjtwQc/wRE7E5EUKDhVplCWmzqRcN+iCZLC8P86Vjn/Oaz
DpeKCOuFaVmH+erwvQjTWEabcv9E0XPg+swZ7pHWoG+oIbMfNWmlJTTDT0qZB2wD
hjIOmqJceCifgHb+yhe5rMbWD1lamQv2rHSs3trvT+ZADEcOEOQrfCWz4Pvu1jgG
8dQ6O0AxfD7fSITrQEckYxsn4XrtpyPujRTyLGZTLxP/wBktPEDmDfw73q+Xwil7
e+ljy2cpO1JAcAq3tzgnihpJaCamTTszPOqqsvG86AzAJ1Y+oUOB/a5cWqGdIpSn
xP2cQPEgsnJUftW4/wYVl+tpAh0uS3YSVy2CzHWARQMWNk1gGattBUE9iwd9+DgB
lGp5YAhfTRkA4EB5cQ6mx2tpkUuwLMdGr9okeRdBQMtJ2kx4rKllEA6b1s9Rpz3O
hv9GlgvRmgrEaxMNNgW2cEDHAPs+LYmWjXoV4HuUKLs/NL+ZBoNsT8Lkxug3aOsD
wzybIyWvHXMmChq5xfJ03h6gBO/nWegCGMuB6FaFh+R0ZSGyfvQ0ji4S/rroL6H7
w/4dLrnbldtMeib1RqOvsGXEpJZ/iyPbt05c8SqzEhJMjRfe36ZZh/CPLgoWYqWU
OlgfrEz+SEDY0Oo/jXEUPw7O8MlDBuOyD9R+WLiAcPYIayj2r8wLVHappyQsOV/k
jn+8r5ODSKgM7qon8lhF9/P+yA03TdOoRqytcBTtogEdJcgg6L9nYO0vTWrb7RhN
3QbMg9jH1JHdTq+Rd7BOzBwIl0Sy1CLAZqRkqyN8N9eUMh5lxTYEIMx/lcUDL1uw
FAMfgmgt6r/7nXUqaA4pGSRN6KikHGm3qfaeRYDLa5DfQKf2ICNCBZO76Drm5xK3
wx2htZkMiUaUQAwRg27VRuP0jrFqCKcIKbhrABQo5/UN9ThLNiYvdcfZ13oH4qmH
Jiz+VajTHCA2/iG8V0ZnedvXy2YljhLTHK3Ha1mPn0wmMbH8Hw3YLhbu2qfKEaz0
ppSQ8T4Emx9nVLVDOiDcg31iiOq7PpYXH0WPpVs8vV21JDSw1tVyud8qSkFlMx79
xffo2PDP+rZetRzmwvFNJUoHFLURO024bBgfMldkanrIlFextCcuLhZmULBMEjEL
fxECMR0A/UzDicU4cUjBnpbSFU+Gs0rVJyhdrhbze+BV/FnHXpGBFfVotKgAuNtE
Dckj5MipJfY8kNm9oIJx/0J3d+0V/cluZlbVpDFlTrzp1ho/SNsHkKBVVDbwgTya
QFnPvuDdeckMltl/cMgimE6UViz4oLMHrBp+DxqY+qsKV5pHbxfe2tE6xV8nxKgp
T3P1WBa8zcD0Q55eVtHNb/df4z6MeMRylJOUBfUEPbineQ09SdDQmgLdgXc992h7
GPbYh+gEnIcpaSTFQ1AZTRsXX0tdm8yl5Q7/kPPIJqH1nfFNucackmy9f81yQwao
LYRNL6tjmFOUFlKeWnwQRF9krcPRStq85RUPmAcYp1Hqb2ZcSGGexYragf/uKt04
T3DQL75Wpiw4nZR4ToF8hACsEldA+vWd3e9Ecux9XGez2zjPgN+7+uTUz6ivbUJS
fYFmv8jCsWArk29/7MQ/SuPWLx1MvqwxLU8u5lIE/RFJW7qsMt1127RM33kjLfLw
S+O3nS7YkU3WGtljmBviN4xGT5ZMECdVhwy9jnb3Sl92fejcngIUvGKiqq23UyQO
FAeWGYj+9nFCJeNVSVIzpcY9r90Dn+bu1CZP26Evzuqm2MEtHKavePyozY8PY2lF
MiD88XE6Qf2YPol9oq3dUzBMfjQYOKIt/Hxp7pne0EsRtbAbE3s9EEg5PoejLzOo
6zWRlAARcBLX2ubeooxWVReuDJwkqxGJFJQ5Z7w0fL42qh4jzy04IsRLkbTt9yXv
fTpC4SPwkiHtar0Ht1FbJzu3aLYJ7dr0rGpJhIElCdrZkXXOeajExdeWa9fRklX/
6OgiYw6lbetr59i6asANiJr7qdX8TDUuUSxxahcGPed5DKDgLZe49eNNCQmbzPFK
WulK220kw4HtaB3fT0Z448UEO7WJPryzVSqxXW7rO4UDaVDYZfQCamDXTNgyvkBb
HGJvfSYGKevt5lVN5oMFcQofeoTqjOAIPwsAUR9Tz25VI0VDdWMi5C2eZb+sd6Hp
P6Ca+3YGacboqwetWbncst9dyrxCeRymoPGAkpdUvgRk47h55xiyDmIMMy9+XOV9
lYoMCQWWF1URYIFM79yJYRWWmCfXL35WgOGEawu2Gw+WtKg1LYomViz0FGUqaV+M
4jkfYbIQT7Vg/YuZt27giRuugX52BYAOE7I9FrRVFus+M5QDXtEcu+Ghtg+DLzO1
L137AkrBDZqF/zr79/32xUs1+8DLcuTuWMXQDgIVoLAdPo2vGdDY0xrHavZXk18S
C2s/0RCIzDQtYWsTVyjGRe55J0BRvve+XW2uD8n4/7c3J664KChjdCGrH0n9lRSm
Zf68BqIIxF3J3qWlzrS6MwrMm62ZsNRBQrZCm8LuX2vo8A+yebKCk9RlZl4owVo2
ok6Z0QIzWc0B3sxmMWcrr8sgdb0fIavUW+GZMIFImOIgC3uUkghDU/uBuII0J2/c
nu3gBtBlH958jAvgY0OAJbzZtsOJS+e6yWFe76Zwy6jy8oFYOaQysdgOAV5s6NC4
ivNO9sXcWEXCGVHM1Jbi2fnrVSQgpKd0FHP7ByPYzYNsYl6XiCWpcJgN8hczDFsY
CBg7qufjVE3VBSgPkU1JJqB5DkjSCO6mp2+yxZhmEh3MOUvBqtFHXfdO98PBudZT
7pc/uVChMoYBvFXsGWyw+oovRGMNUZpJTtnO8FSP5srXYCIxabqjKa/ZZgmvOWRj
6tUq9Ghs+qqiLJLLPn0ZXPuRyoJYYJ/5CxKMM60WkAWao9kVrNq0X6yLEjEiiDN6
hDgvtorfYmBhTdTxh4yTdfcvx4V7AQPSAsG3AzRj/GVsZh0KPsfexAPRpiM7Xgk+
9DYHXbXWsW0dShy3AUl4XaTkQ/o848ZBIMJ+SNFqZp8jET890Ztjvj+MkN7K9FRY
J2R2tZfR5eRlgIi8DVDPTbChvleyPolH6c921GU9U+D/cm7dY1zPI9oS3ygpjHRi
zzqb9JWQfEKmkOHkJrSuBzfCHjYNWRuJfnc2jqbiSP4jdXudGjyqRMi/MLCBxxxM
F+mw8V54+fSztsaKvVZfzVNATlaPWrQ9KCe15njQJX8NLeFQ2B47ZjEmXPe56wYX
679mKKC6E68uW2DNLEzS3pk06dlO6RzEQKJ/GorAVPPBXaad4sNBEjqGrJLAYXKu
WYTs2yJolGRNWOjHbMIZMuXb0syUbftv6qxODcRnFSEnuQnxkwKjnvEtqu74NY09
MVTE5pv1s/6PEuu93NEK/j7yHvTesCH+XqABzZBoseT3+yvlPHZLikMEBpc95mGH
xFONK3aFiUrUk1jwNAaT8QNhXslDPZFfu9jT0KTNtQDv32i4KZuGkZpa2fQG/MRz
tKH2IFFBFWnIBtPLIB7IE8oHVYi4hn/NvtN/EWtTCJ0aL1SzTIjAZBIk5yoYw4re
nBRp5/s4skKRQZC9Gzdkjk1W0zfPZeFt7ejJqd/3CdZNmKjboyr/L5LCQDh+Ensr
nxFY+Bffnt9NWCL3sBg9hytN6bk6co9aq18lEk3Go8jCIroyMOMUT9NYDTkTOkIL
DOlDxXXOKhjUvON+38CGq3kBRF1dvRNT89QRCeCuHO+5fO6sUbYxynaV2nAUeDyj
pwAcaXhtzo0yE068L4PFQhdQNMmLEzv0rBb5gxuNunoPEckl787m4xx8Y2wyXNM1
Q+2FuKgrFn6S5sXSeXvmpd+fwEvexeFLXElnezwtZibZIIeeD7fkKiFHFkRdHk6s
uhpuSfp0mSTwYRfQfJs3sm8LsszMs0d0D//gnMtc6mKSs+Yz8zpo3AOgoW6zBjTv
7jp8GOR1gCSG5VoRjRHiMkzrARBVVLJ/55RSvnKf5+h8Av9iLITNJiJFVQ87aHVp
LwUKxi980AMA3dpFbF3F5xmGd51SUYc/pMj9itSo8onhWiRRWK5FD+c6VRMkDgWr
+FUxJ5wyWegj1NgxFCCEIXtSxGlzoC2LmVYz5qK56Bhb2Sh+WY5joF3BPW72pVT9
zV2pkM8d1aD/RozVaEi6W2q8OJ95s4yHVBH0lyKs5rsWfsUuxhUNoreair/NscsH
hp962ifvIHKMrnBekDZhLbRZIGXkfXXw/+dK1O7gRA54KiEAYp2Y83vMenGS11CL
Wz8AbJibxs/y9kxJ0q0xMxQkvsZ42FCAdAmU4poRZKGBiU4YSVqBV4LTp1P8A5uv
AyXIODDb2HJqoyW12DclMTRKrnBi6NfnoQxx4lYsBWtkMvZX3To4rIvYpOpLTns0
5W6OT03bMhm5MHLNsERdDteIbnmmaR3UYCVOXognYueV8N3BbMnwuB5pio9Fy46w
mN1gZkCpkT2qS6Nf5b4C15+y87jiVOS5BydxJ+NG6I8vpDCe1cDmkIBu/cU87oLR
oObN23QXpaR0aW96NvMnV5y48mxj3gAvRYuSqqD2exjKjBCtP5mzv1eDUqvppwsq
tKxCzXgeUfeBYhgh2Yap8SAPOkqvdZWxdURl21ZqOnw/UEqwz1Bgp4Ymixjl06j2
q3C/ClfvxtGVxw91OOHyh5ztVK651AuQYNLlDMWeQafQvg/P2s/1QoAK2KmL2dGV
/WBWl1SqegFYPf3zPxaESC2ouBibMkACyU4xjLlNY0v90MH6g8nHcOWyPNHCtQgC
05f1eZGTxZTL6YtJ5OXOKXgHXv0c3aM+otyLCjc3SAf0EX7y6EiOnrQo/jvc0fMZ
fG6t+xg+tZYmLo7m+OgwvKrmFxiuqh5Cgt5gYZMJosurQwa7LHt0He3pRzENo+F3
cqcFFEAkbST0VgyOU3t1zBpLoHpITDs0Lo7uTSPjnD+j7JFvyiZBhilzJURV7E9w
Tj3FCej2ow5Z10QZ6+fkmFYxrmtZCqP2czI6eFc6Q4WDhtOrld1SYDSDQtYTTUZ4
yE+CdHR7T9r1u7y/xaX8UaW3sTcjFxcwnCFyDmCUBbk+JxmBB2fWfZxldhsgckG2
iDkMqMi0TL6wtXtSL8UZRk1Yw/NT1LFM6ORLAq8MGZSbTZeEqS4UFKHluQh8rbGo
WomrHlSPvRnNbsJTfpQtHiCcn/24ffCiiNBT9XHPoaDuIw+BUJjeX2nA+nTVl727
QKM5dWi3iBB69JNM+kARzQrQhowOqu4qIR3sfcsUyFRbu2HsDMUIO31OlNoTJDFa
9rCMWDD+P+XKnjNsgYsr8mpQUyOOzdlfY9XVQynd70Y6LAUf8n5YCLwrxpExyKDS
137qiuEJ4DShfsIhG4GJAeZzi9SanQ4gVMVFKC9Q8yghPPNQQLuFaALc3mymiTkm
xfvWoNxD5WsZ/sJVUnV4mCAE32NG/LezCGPtkB5xCNt8dlcKbd1Y0n/cND1GnA4N
Q2m4/IWyI9aIyN4qT73v32Kd/6IA6K1QNQDFrPcq6dBleycHbCd4cpJc2lPFZHfT
EExtrhhlQyAW8wHrX41j78fedp5afDfUbhpy2y3EapA3mCJ/OJZtonu4mkhzq6np
p7dnvVhe2etRt2vV15Asqsnr+53UALa0etoAcriac7W79m8djTaQyj19aLKAyMwq
LeUDFg5JWRVcHxy7Kh5zPmYJTQ/AkoVpvhT8x1sQmkxA0yVO5Pdp7qfC/KjRS3VY
IaV5lEkSXRnu3fBzEVMIINWYm4haOHGs01w0LAZIls/enII/95cEKoQ0i4hQBcur
dLRgZ3eqc6+io8+q5/20CSmTiJkl1L9F3gp3gTKj0114cN/jes6hhLtxboNmXCKa
FBG8nW56AV+y+CLNK+drv/RW9wSOk+GCzW1JV6hTdNi31LK5hCS+La3kVPJQyjmL
pA8KnL//CYUCZ2lEPfoZCsjAsCoW3F7AbCJi2/Z7wA/gx6DctPX2KouiRqBFCVKD
rqSSVQBARfuBplAp1SGAg/tsDoEXeDkH4tHmOW9vCD2r6txGZ+8yTuRFiKwZGNYY
QdkHbExR3grzdO+i7JJlgBu01XFSXnZ4f2MgJSsAv0yj2yUeDw5+fUrOBm16XEZv
XfVb/Qe1Lp0e/YotNERqSBT/79PhTf8gHoyiMvJhHso4v+RWr2DDZqIYC168tpf+
CVwCZlEgzzPrPMTaAfI3zujAIFFvbTdfCm1dGzzuPz83UKb4Wcm4Syl8iAorAdp6
7axWkdUVGXSpUeIFNXec1iUlMV7KfQB6yzKQ7qdAv6i4tYpKGNsMHH0NYtgdyeOy
USA9u3DkCCqArw0Y/lhGMjFgi9pLr9Rh7jeCaGDd8cGf6MMRs4+Qw5aOpNsExAXl
GytyfTn0B4a/i45GghPc9Jr/M9+3s6m4FdaGLThWDPmdBVi9o9zoDsMgPAK4FMog
l7zRXNt6Qyf0+KoBaKoIDQgl5Zy1sibxEfvecixv2QcjUTkdCUBy4+kjci1/H/z9
ekGf57ZN+xZthUgO+YLEXrjvoEIZBGV680LzCOY+24XNY4O9DJCrb8QPqY3amakF
Mq6vtENOubD7RGatY1cx8OBxFTZKkkaf0ymMIt4lkXQxBqox8r7YZeA/zjUAb5I1
pdPqspKIlINO9KJvAF0kKmrvwsYtKbAg9krs/JMvSyKjQWAuvY00/ij8reXqjXvK
Jp+Wj0xd6TBO7vSD2c8F1ni8noMyJgsGUcvoCg8d1vslSRMLfvyTC3b2BkOhvlfl
UtvPO84C2SVjsrwW04gAQW4rFrkKDa0PtPcxGas9ecyvMs742XvODE4dqzAHUQWU
3fQlK3sZ7BYQ0e/riY7R3Mm4ye7As/BZDW5fnck2RyjgWzh1t9mGjiGFXwNKZKUd
j8M3TwT/BIh+B+pNs7/YgDZkQd/ceA2oYLP+1CzMwMpl+K7ArU7A2S6ZpmJ0jlSZ
oYd1IR1W3s/H2cCK1ztJ/wGXMoBXZH8hN1Vcz6P7rwOnBG52jr4sGVqmHrXEvgvj
4rmepQD0e6XbCLcKPBjFQ1q/HKI1uiIflcukVOH3N6qgoqlgrAcghdsXG9mdW3EV
npbPsN93H7eg3GNhCVkiMr9w5iNmS4PT7O4NW62Xd42Hv9fngixS0Hi2UhJSoSG/
xJxnTa0X9s25PNqt7P/BsxGchtAO2g83LRZXq27lBSDQxwtdMK61gbIsTMjvwV0P
ODltp9hwgcOtvCmro6htHI2rojK07zoW1xy8/HSsHh6mKxM/WhQIAIFAiNy+skxp
mbeIhGYnhdYXInpDcTMOZM7Iub/yAjvKc9E1szWzHZNy8UV1BJv/ra3B7boJYhZl
4z53dsWtqoa4YBhiYzQTY/uelOQ1baqScE8ufGRM9IA7XWLGaJI3YihKXAGnlguJ
lRbO/v2K5DUf/PHSulm4UatE3rut6yzl9jLFVHwq7RvowTMQAwIPOStvvHGmhGHx
qMkWfNwqLYUUDIcHow3kxY3ifQar9ck4qK2S8MD+PHpQggka+zWVFlXRixKVX24R
2ZRmR2EVpsUxw0fn6CJ7sTDTeYKz3VCivejRa5EeuLGcVPKyDLiTrsJWHiQc1e+D
UQp97tdhBUAUXy+vBh0mZH+xK1N8m+JRT7rqLubDS6ePhUsAFa2rlSxWdagL2GIH
BkJlU7xskFB3rfYU4k1myrnjHPt9pFkfOm4CRk8VxTcDk4g7LdW42c+8WT72zmyD
bJDOMPB51olIipE3UNj49/m0XbISR6Nq8HAS9WrWwmxC5dCTerk+ZiZqvR/CfMQW
vggvA7sHUQX+LwOllCiOtBxVcLnlKR0cdAmq5/gg1lQvl3smxb0M13WU7gh4+lqK
HngqzqQk21joU6aqPNcUhaImYq6QVHEUbye2aNXsrinkweqrHfroP9L+1OgxYlUr
/7wtY5N2STmM5HF0M4QqYJGeLKtERdqtm7k8+qIrIqmOjev+nfxnVOxEYIQ7lz+V
FzEVrBr/q4ZTyK2o2CAGJWEgs4Ip86U5hJMO4iA+z0AKEuQ16SX73lsuJul42yLD
hBfarXa/Fvp+3ME/ixVlNLC3huGk9JnlbtjiAihZD7arVHFpabv2VMbtYO6rH+lc
XuqZHzRn0FGnLt5AAP+3gYxxot17exFSHvdHWM5oxt0jI70TD6hQUWwuyMWhrmI+
xAUbm0OOAdWZ3fZuV/aMSoMOxN40CaEPEkl3brrT00vsE4fYDQTlQd0BzBrE+sE0
MGpmCBdCXvBYJV0iMwkfRgp4Z9d4qDdS5lr3GlgRtMTPDhxOX2uNf6J77OwdHWhz
/GHHTaTxDqfsjy5yVH8oxY00CEtjFWpPuO9nfJFvBh6NpcDKPQBS/uC1bMwxWoYh
G7/WPaQr0HVqb0fsj+IrtjMX+su35sQxAMoR26k6Kp7TjlFQGDqqf7CoHJnSw1Yq
WfoGIhbl+t05A05p/LRvFogV+EwjdNrLqVWebdV11XeqkhZqhk+f4+YwqoNYzqgN
jx9pzHR5Lue/AWvFXg0k6gYKBuhDkLgcQx0YWP30cnMMd/VAM/EJaom5YwV8dmjX
8m8eU0E2WpapewvNByQSVxFXVBuYng95dAN6zg3FCdW+ylrq6a/jse4xMjSwtc6H
GFNBnL6H+1DJj4S7UTGsuNPhnWXkKAap66/Hsw8KoWOiOehxZuScI3/Nxe1igb/G
wmb7/go+n+ZWFfFRrIZ6qU4Tb0ZMVzuNQdA0Nshjc82IDSYqv/zEj9lTlUGSKOkk
jPNV9rM6V7J6iprs+Bu5YWeiYNY6tybVOc0wqi3HY6bvK2y1ql0AM8ricE0ZEoUh
+5E9inU4BbpiKmqmlfVtafNaqDm2FFt1Jqm20wVT2ZyqsE5rMeXMN57jy96U282h
GymkMfcv2bwxvKaN+OoiV9XwFhPx9JpUst4v3GzaIYC9UJNsnI6wHKG3+C0SShO7
YAWPisAkjpLzVyeKn0jCptjOy9egNHZRWdqLUm9T0pmXnilWxGvJ4hCJT0NoP8FC
3HaPgTKva8EAMZ2nd2nflMNRhGn2UYjd/HUqrST/W8N8u+D/j/A6gqkA13y/4Fs3
rPrXXXCM4EYpEGHBAO8pF1FXKtFUNaj0RJWuPFMkl17IcF4AB5z58qmvFkNmYiun
f4+mLZ4PV6EdZAQhC0kKU9AxEp5VCZXVqpzc3/705VzHl90N6e7mvU/S+N2GPB5O
yDy4OIzeKcZikHZ5mx4Ah1qMyfjdxUGYlNFAhmXBpY1EubRGJTJtDq49idIhPAD0
vBn4QjRhYj9g44IrK5KBZDEZIiD5gHyCyFpnko3WQPP+bZDZfh8HmOWSyaQTfdBM
yBgTkxFClwuBubzZ0gt+ZUWh8P7247kT3xx+aRbTdgx/ijIkWKGvb6uP7cjf1EV6
ctl4Wm3DhgKbJDqcTFhlO8/ohCP9CVUJCq1AOrm1o4lNtSJKoGcvy0YfzvIN4D5a
BrtFsPjpPZQoj2RLxfOzsZ1K2CK0QnRSJwP++oqhIrm6y+y8/s7t4GpumWWI9kwB
iAAS4FqyXiEp3+srKeMruWjckjyh3M/APZS51OJ5QPLZFOPR74CXe5NoF9cn8Fsg
4ib1g+b2YfSSuN4qRPo1pT7UmGV68k/qNQlhJMdPs1dpAMLo+xYeH9ZuT+QrfYxu
slXYToEJdHiTC0tEKdLMIG+cOtzPAoCqLjYQWN2F+DAnTUnc/tZrkH86YCTZaN9P
T5ftbbQCovbdiqkjVFJXfgmvT70/22Ioq0GhU1IpW7Wkg/VgZY2y0P0ywx4KaWoM
qbhAX48jJ1KmIHuDFNi1sqUIW+V0JXYj4cM2wfLiPydQGC7T9XxH6ew6Me6Oa/0+
zHGqhqHguv4657n53+mFpS5zlLf512YAKDpJ16wabAGyNkKP7INqLWSpkzUdRK63
+fAxla4NcVuQqJ/8TrJ3b2owiBqIY8OPXrJwzOCqPINsLwnumrj+I7AZQaijWMiQ
NKZL7eidqXLbnqP1oLF80nHuLGQ3Ic4hlPjQ8G9G8UDnYiwKA81skS7AvOAaceT5
n3ZYeOIyK2vtS3J5siNyV1rPCNmP8Ew16WLiNBIB4530ltxcnqoT5l2YZPKPxyG3
yUe4D6XF9fPzvhFyF7n3WOp6WcDSOKtazusvEjlguY0TZ64htq4E1p4Naqp6jx6V
WT0zL64TFMDT8lnI2c/OUjpKLwf0N3qCve3cqLjrTCFq6vIGF3gk6WYs4RtcHz5k
GC18sktIbliPAjyw19N2/4EXPDQd3SW/D/YWORFc9XgZ8TagOVMosF7G1F7eR4r4
zqun5OgJw4sViKzpt3GX/399/bEsqn/M9e8QAXgv5LNBDiFE2dLvqBhW/pEEnEmP
lww4j5Y6s5hG/NhducVnqxXj43p/LDwmUMvszm08I+P5V0QGC8NsJIFhYHwHQrq8
LvY61x2PcPsF7NG3mjG1wpfFt0o8CI1gqqUzhNtonKTCkAS4AdSP/u3Wh6wzvQXa
M7E+0ZiPcm9C7KFQ0ejvZsAchXwPTfb9c5HgqIq3LmilZl5y33AP83zoVhjAXaRd
CxA8LR/PaM27c0Wxtto6ul6iMAMUVHS3rhTLEsS17V3r6+YD9r1G6/gPuphtxiAb
ZSgOG7oAHV8OwwWzCa68Hpbjg+l0imP3e2EANTItzrp2DyF9e2O9LNXRH/kCItqz
N7Gogd5ew0e+ybXuf69InJrwOP1Q73SXpY9qn143JBzX2hEhGNGGKBa54zNnQel2
FOL+BKsyDqAwesdIIXYSs9du4joYF6YLqz2HdEDDxTT+3Rv+C7qEzo+BkNtPONKP
VLu30RyQb4YRG4Zbu6dGZzEbAVrXnPxqnvKC62C40r1Sx2Whw1Fjsw24lvLR1kQE
zTMOncgtLWfdYEhdU7hKX/4yPCZ3sbMStHmQ0cI8ZUPuzjetDOqagb90JTjhCfqZ
66NkNMU0SxgMf09OULP/F5MtW7yOx77qq5lAvxSFe4wddJsWRwemPO7gGahapnHV
8gvFec7NgGnGAttpd6U1YAR4kJ7X160tJklK3zOI5pHkf3ypvJVvPBmy97FIGe2B
jC3jV/3TF0CdOx38uhU/8hh44B7FojLY7KtPJ1VQB5urNpZDwPaaKTlZtUdcH9m1
1vDuFoe4/Ld6z+INmT0yb7/BWQgg5hVz2E0SeKUNYOgHWDN5sMx2hhfKIo+iyo0t
QOiKKTQXOXaoOP8ZDm7J74S/iPUEEF9D/1KrqhaWex2I6xisYhLOHEI59RKDBqvF
2VFCOJcyWgRDo/M+Jz7ExKKoaEmC+PPhxMCWacz2IKNICaiTbUXkZCc38/LefHbH
VWPv3m2/iaAyvBpnjvVfpXO7RR2WAXgkmF2c4cQRygw8UefiZo33spowefgLSXtD
ZnDLTyzY1VamdvdIpNKZPu5RoQd5pgbi+WqVJZzu7vSKy9h2tCZeZ6/qIpv7w17n
TdZRLWYyqW5Bmauu1zSCTjmAgHzOEVYtrklyNis5fnMPRXk+Qg9OkJfbm9datBHu
rjXyBFyHgJx/yRPyeblwoH21nboMM3ogaDUFSFT/ZDOmJoyKGF5qvV5RE1YnOrUs
lQx9OUdQDVvliV1gJlVkBDY16N4S8UQqemFAEWO0q0CPxZuJh0hlOI7B4Q+wNCWI
LHHvt2Us1SMK+wEJUiMX8o6J5+H7h22lo3B0s1HAktLc+Fc0Uk6y2NC3nyXGZQwG
YqaLDkkTJyxDYv+s5b0TbXu84sEm7FSdC0D3zjsXlJlrcCM/x2RZAdhMkw+WwT4W
3YtXMPU2E97VNlzcoG9SNQzC4EUX1Kt9S5hYCowEuIuoFZffJcTKDqyL16xZx8OY
RNBgiMeXr2m2vAI3QeWbytT3P42GKUHm8mSTsKNX4z4eSy++G7vbfXPl7l+1lEiN
jp+4d+1RRpEGRHSGcaWhW1zScfnaphhpLaOh7w+YHKRRcBUWN7+dISTh4gBAqFHg
spihshav8Xy8bCbHyLzA+ORCUIfIrMm/WISrOKV6mUGESMIdQ0Zw34FShT0oS1Hq
oF3hCPVk37Qgx2SZ9ogIyEBgVbWAoVliFxGvNDC07bFifd3pzWOP8ivT/NRcC2B0
oBGsie6w1CKfoAoEH8wrVxKa2jOoi0HVDkjeHj+/I/xOv4bNQR3i4muMZl+pU02Q
Q92/i44J2ZvVpAKPACHGG7A+2CLmwpIB7pgjpN3I07lb7u7py+SocBJ7t/2fSxRX
1/SuDC4eALpVUfM/PN7z+h4W+qClzE+ReJraZBHVIpZn68wMih2yEut3TXIWVmW6
86EptD14aTXMQys8+YfKvcZJIEkS/qXZDq5PeNSN4N7cag/p0mkfP5DMsBgCCCpV
RmFJk/BvWbFNFJ5XEIZAw0ED/wDBF7q0PegYgXa607sLgj7EXqroV1EmnUqU9PuH
IeUKhvCcMAvNuFGz5pI0rsHpYhB7uqiybutavGSmuxvZu/iVFhEWiI7i0UXq27AE
AA7oz1eoxzstSJ1rjcSHUgRhfUtLCMyQJGLPqxUL9ngQOFKOdle9UeV7Z0z2LG07
X+C48lFKPpnrluar6D4BOtrEXq+pL1Qk9N5KR6x0CeR0vj0Oz/qLC0rddtDAxJco
uOA5HlBRZ0IEfUK0cDNHAGEhDcNq3SWP4pVsHx/Rx8BCP65Yc8QRZJHLY7WseVWC
wrAgGdtYJzEu5RkXcA8GfWpYBLK+Dn7vI4QrbyDYmgSJI6R31yTVRntyZgjSvnK/
BjgZ3qGihw4UVWEJvSS0pSe/Qt8Q5toko2ZSmM5CV2BKG+dHpbw8rVpNO6n6HZIG
e0j1TPjlgJ1uyBYkPAc+lSwp/Ge84C2jYPVl78cY0PFbg9Mcpzv5/SYOVTs1zNJ7
KoCGvVOkTFO9eSCn1FRKMakJrpOhA8Bux3BjPzNuob6wQgl2YQKBpq1NGLfrVzqb
G4jTnD97CyQ3FcJkHizXMKtTgiH55vWThGionI4MVDqny4q4MbyrIB+TxmKqAQnM
Cx7BQslaMnfi0R5/aGV8WJSZ2sh39YjnmOq7tDx2GYBLMUfTVOIWjVgFSAmpZi6V
tnXqL76K2RKGeY5azPP7VioWs8M8EaHOr0pqEV42FH2PoQzGHd32Ypyl6Tgd5FTb
WLldQHd2lyP+gyDUjR96bI9hXWlDFkud1lxdNAtZIc/loz6HYoSEBoXwszpuL4JI
jXCGLPPGlyByCSuIzKWd9/FUUIx2rnmraXfZVINDa1u9QQvCzfgYqGQ/E/h9S4d3
JtNG/lvNyali6b93pTaM80t9J4A+cxseI4OJi4QJHVPCNB6k+oherxhzNJ6if+TZ
NVssJ/XRPNd0sqZaCGpoYa5fk2f3kTVH0fUlzIf2atnofjtPRo3pVKmbkyM8BDCV
Hr3mB1rEIQBBksZGTx4rrIYq5oGxlkMf/Tqg+fzJLkzh5ux7MsF8nPl4o3Li5qtN
guvIyIiSzp+6xZZ844HJ/RKwGDcxH1xIxdaDfWmrCSdCPjNWRCuKBLuT9977M+WD
e15noKOEKmza2IpAjbtlSn66r+guL3ZkrZDX3xOK6OnSjfaR2uqJrDOJ/k/3FvnJ
s0VLVWQrQ6HjTu9EgY2H0Afbd1NO7/gVtgRyknL9QCMVMDgQ5pIgfMRUg6ngCqr8
+KLgRhMTyLi2qSXU8A1KgwGMfAk3TUgOOCOYJpi40ov0nvU0WtafSH1JXCmIWf5r
Mo8bWDcgvoK5XULy0+cy8kFugnArSWG0RQ73Q6rsa0pS9MePLX5Rk5mJ9kr0e69E
rF+pBy5GdwPIY7R6nnDhmDXCJSblif2/KbnCj+QppJgX9KfcE6RZY9vfRsSgl/ww
0fLVx7Ltpx0eqP1cBSukVtBPLlNWFyu/HU7XzmWWN/DhJL4wul74jR0UtjwRT0Zj
37xW00oIPXNIC1dsu2DpfaZUUacvVk9XRNs1T+kgACeYwBZLQM3JVLRroLPayrx8
xSoGmlyCZbMzeZ1r0DvwOoFUDq4BsQIU+f44m2fsQ3F20OUqTNm9aLDbrEQ1v05T
5DkRR0ZEQxfCuhJLnkuolhtlRUk3qXt07kPfIiq7834tfKPTehEE2GbO2tKYcmvS
X71cJh+/bj0/RNBOSfgpqGYfyCxe33QafxXZ5JRKp45J+vMhaprLHOYTp0pDxcla
NLIQfVf06nZMFbu3SazjX0TDIAP4h5+r+V+dN/IxOUtaAtmMO6Xp8C+EhQRsFXpA
Pad2ww2/pv5IECfR9FWBKUGJog7/tv/bU7Rqf5ddRALDTYBPgQzhfNqL9uuIsN+o
rTJRDakWbVXk0r9L4c+qhDyqhWnQQV3brpbr3a0EHbKzQ7ovtA8XOeQjtU2Rugr0
WwHfvbYp2kXiKE2uU/pDE2VGgKwIDMDsEs/10KtOf3KBaIAsFF4QYfCPjeTbgJHw
UpbJj4kXed0+1pO1Y7ErDr/9UzL+p+D5DdsYUZVEfnzalIilDhVgS7K/XeFHj2Pn
UDE3TP0e5qgrHCNW9yaUe+hJ+cjerTWwEAsvrTo5jhAv95dMfa1GiwprTRDdZw8k
M8rhcIrqNw83P+b2J1fpgyg6zA3OlzAyCLFuUG2/uWDJS1hFC/pB3EVyph9Rpob+
dAelDVknUsIcvDVJpTGH2QDo2Y6+dtX4MpYRwgyapa88EkzEcUrYeIX0oGFwMp5Z
McRY/7BwCSuoooeNWSkbm4Xr+HHzpxxrc8MD28f4WQEkdVqDZOh4knCLuZdXiWLe
5RI244dc+57Kos8OuC+5fOgBnCADskCLLeAxNeTsk7mYdtbuEljXli17Mo/Gu6+u
hQ+PhW0ECTpiLQva9ufLrchswvmg6jfkp7WvP+T5r2GHO9MQUqaI+LJIPgHGa6Nq
us6yu8+nqP0wW03wIes2/mZQ4ip5VNaV0UE7Bqg1J57hWzFPg0PH9/x+dPzjNNWi
3nXMI5wqUWmfVU347puEen6MwEaX4vW3WIyMI77MtN8lBi1G8p2ZdyPFao9eqtE6
+Rs+0nLSZDREcT6rn+1UU2rrHn91XNUUUO7YOZvX41AeHO56DYl5RGCscYDonxli
LXWkXo6/M7k4PPD0D9MfMzMb5oPM19h8bAQJjuSayVgarjVx9zBlkBg+RfGhVYDH
VVBsrDf6yMKbDOK6wihd79omb1XPu1NX6Xu9qmDoFVF5usGmh7RyPiaHgINXbyvy
0ZEKJOw7i3ZN2TPUuoxYNgg0Cn5jbqzqikE8UVWKLlTGIbL5qbcvae0iIF4vc4ll
j0UhOnznq1of+rMjL9CdwgtPyvJkkjyuqRt5RPAojKssq8Ffqd3ODdLct5R77pqd
6m5plB3lCbTrKDTaASpkVo2NTheuC7AXz40NXPVM4BnFvPgzxZBJUuHajnygpp6g
er3jGlNeniyVKWUUZlnGl9Cav6XTgGarVuZp18czaC4RHuBZfYgLykgNiIMXvj+f
IzAKcmhLxfOibzNPdpTKipqoBBPHmCCE46Pk31zDvWA1X288+USBlN9JbvqwsHjt
j/wcLtPpvfCRM9bh5YfQvtymEXxqVor8iWQt2BFwwBzU91lpK+xVsHYhWceGyECT
hkPlXnNxWDjIuVbeJNdWXzJ7pz2nhFfhiyMd7+D9ODSKRylLYGYKNpa5p8k2uDed
aPI2P/LO/kEm7dqgcHz4UmF1+ohesNcUxheXkQ2DopxzBboQzFTKEwRjVXDtgpTY
58XnEQKmHgPrQpvxeVru2AZGFnXdlkuPrjQ9iMiXqErFvQJXtb48X9KISl+xd/sT
hs769xonwIH5Luq9+yVBU8T0qi0K1g8hYkBecuIL7mFc81YxPoo4X6S72CSdBGCe
s8tb4qqsQ7uSPGIKYurdjzx9jzUJHtPVBSYMSHM9kyI9XuLC+QhroNXd6bthgTqv
nKQv9DeaZozIx65hBzO9xL4V6bYXnkjTXjPoAT6sxzh4AnrXxL0ZUB+YgJrQgnvs
R6uqmK25k+0ON0Lym/vjlUMbNAmnM5x0n+5w6iASaMmAqtn1SWWmYP85NwJVaWTl
8nzoHsotUOrNW4byksEfzberjuFRc+jqU/ZvBXfA/baODqVAc4ze7fmVC6RV5Dy6
ZwIXhnzv4cHtEM8kuJ0LII5fDOBheDdeueVuwAr0+b4hZRaxNwXc8toYY3b1qLPh
fm4vs4oDbkn/MWLun4pyqSfO4ciqEp2apgNXfm8lwIPudy+JbMttfvoZ4NynsIAh
VmTd5WtKXfxRyt9n8sjCNUtYrdhUQAZRAsmy4B/5D3XlUSrH6Lo2oTBXA2OoKeML
3aL+FcWtWF4PA0HBiWm718vz95KDe6iIsNnsPKoL6heyOis9KPaXI0GsWWdnIyLT
bLFCEkg13piHSBZGIkvTDOzlJ1WCsh5vrhj8vQsOs/8plRyAgIc0e5VPmqTjt4e0
DjrmPLevMgMhaNtEMClsgZCVxQPyXSbnjiB0XEoY2m2Zpijiek9b9xoxUsH2JAYj
/duo6GacBSh0TvDd00UXAf09VRizeb5ZD13ugEqQ5kxRcJqClhK+Wo+XImgHJ5PI
JR52S2QfzQ4rKFP7JGuVTDzq/Y0eKjJtzF6xNVgzPfsnXBh2IKfTtnGHIjIDSiuF
bHmgWsbwwWWfu4C9+55kdL3SwPT3Yy0P34Gw0RcKlH2RtO0AQYAod0IfQyt1y9ul
1dUEM4xbCTQtDE4zh2fgGz2a9NJELGeF95Q92VT2wn80ucE+7mglGTYUGn4SacUO
nH2g8XBcMO89ccJOfDZZrSk/CHGVkJWc6hjZgRV2ERHv38axVVzPusG6obGcneTL
BrYxEM41CpCkw8a6s/elXYtP1merbQGBWYXiQixIWR+OHy389i/kwxCP9rYlZXY5
p+N6tdhq7u3DqkVcf4iauPoNMS+kD9svtm9q8kwhSP96SLBKjk25KusRK26NXOoc
dgD+GyzHDQnjdDGpoJL2rp3NnpjNT+Ln5Cvqx3wOT9JkbnROdWYMmYRM5JDSM33h
hewtUvb7I1IOJEnGA7cyxMtjjPfuUP0Ib6a1WccmnZxV+CD2837HhSEJYTxkgHhp
VacQxrxx4on3Vc84zstDdGzSXOJ1DqiOs1LdXJ9Lz6M3MG2rOU91dj0gysJM5E/L
XrP2mUEsP2YTbAY6Xa/g0sQumUefhs48dzyViHbuvOLgABWaikdIjDICb3oSrIoy
4uylyy72q8k2oiVG05WjzF46Rla/tsTjYvR3I6C23S6R7MBlta88QJHNEF1fsZMD
V6p1VlrWYsRF8aJLFCxqwBSnCA10lpx0lWKrRp1BoofRluwGlKxkadg0YKTBZvf6
2pOnQQ5fg9VSNkJVSo0lqSu1t1nR+6/JrbsyMkkH6wPokNuBnVYjGw1wJr+eIBQr
znmWcYB6DodE7pp7fHjOyf/Z1CWfVvhB6J0g6D7dOT70lTH9UHZOrSkBUp/AmT7d
scU4tNt/zY9D/TIiewhdYgqOplA1foXrVUsTsfcpSLw19srWkpphuYx9PnPDQYoo
9BUciFubiEavgWRm24vaQ6gKUTV+Wrnj8UaaGgwO8tDGuQeb1Zb6DLHiaDCWkHi9
Htya8MFq1gX5padJfOOZfK+rLj4MqUgiIa+FXCFW5BotFkFaKb8uG6vxhQk6/3tZ
6T7ipTzEoR04j+jVA+rWW4EdV5zPaTg1D7lEB65fkP84HjY/vgNBnxZgs1BmoKue
59uHFyBi67jl7vNll+WrTPXsDHs6RAX3cHR6CceVx8hRo7liTi8QkVqZEI4JldBs
vdz5kIZewKPoAkaCw5XLiHtjtHxoZFMo95J1ZiF+exp4/3MxNIQnrF4GXDmtg5xn
Va5qTW//J6YxgEyByiXmy2LuQaI7328J1xy2UeUWAmLZrNSRKdIaBxJLqPRNFSKv
lhlXyc3jTBgp1cDY7gfkTEBgEjGi/LtmdA4mEh5aqg/ZDEryW9dFrNWv48gSlSGl
xpemiOauqcb0cB31WG7/WLzP6ejh0nm65noaLhhrX5toYg11bFU4SI39bXQBSLec
26h028aynqSI1GnHmqk3yLbTPKhdXlqDMHGJ0NpHU4xYzkxM58mSCN0vGs4YNKfw
RIRYLNG1nFiMAxFK1IZLl+iMVjf+8gZyYpS1CFPC/eY6N2+qLsNeYklPbk7gUkkD
s3tRsV6EOT7KujILPt6KuMC1QeMBSRxBD3Q/TliQcIr8kfsN8OcePOieY2rwxsgI
quDA8zOQDH6tk1+YgdSEk83apwa+d1c2+eaO2OfeoL/nYELGTL7leyRMo8yba3Sx
hfGMBY8HN2FxZlja1RuDQxWSnVsO2Sp5RIVUjbvh6JJQewNV1pLXN8lb0c07vPYa
DCU0CUSzcvyOuPtQ8hGJmMEmo39sjgW0bh+vU2sh1w6OuG68yV+M1NNIyu7pSmHt
2ZAW4tNC3z5C5Q+XjyoYUwRIC+TbCCPgT4/vOPBDwmHToeWELOfOfZJXwwcaUp+2
CMMLoxxe6to/n3Sy/GgP1sI2RkiIe+6+2pJ492Sbrq5Ao7Jpz+XBs5NQ58dkstz8
h3+zQiyKvwFM3QrjXygpXfdNR2g4J7R+/ef/DMCDlHk7W7OR42ifgeRP9W1EivI6
EPMqHPN9diNLarfu5d76HcITINtXCnPSU18JD0KtV08d4myePD5nU056qbQy/d68
0bJerNiJsuou5mb0Ijf8UsOg7V7FNbcHnmliszaktJkWTAl6rTg2Lcr7BsIn/G6Q
1zuFfOhgcI2eO0cjOsQTI7k5FznvEWDpckvrs/+Hs7kV2X3GzFCgRG1xUqEMTlls
EaND42ZjLo8MApz4PCFNy1CzVV/NfBuKrEolUCbp/UIzh3PAfZh+SJereKNg7kyF
WVIPnQF6ORcaaICjhwehF8U+d1bnj9J2gZfdRoPVwcQIWdUkkI5tqA55Sf4MsM2i
FT/8yb0SdxYeXy8OWw6S47tKQj75x8lfuRmlEkj42DpzrY+JoyEXc2dbtwRKN38F
qjA2loIO8+iAXsYfynsb1lsPlWANsAP72yMEPWUqUSmgzgzHlDRC+mzWWKjhJPby
8h8MeYQQIIzpdcE1g5I+90XGUkpU/73fFAxzpUBqJiZvH+xgw4JZTntBtdafPdyl
9wkVG0IN3TvirpXVT5UI4QZ/HqaFY6ZUTNHlGMftw2F9pE1RTC6GDq/ONuB/JPEu
av2/rHvfMpS8+6S2n/dprtBU4ASY1D/4V262s4kujb1LXTxjgBTEhRwmtbWXtyTY
XiojHzbw/u89HWXDoEpoE0axE0N9MnabMVnB4bwUnzofC3O8JNKr8tFq98cFIJvt
BmZSZvebu4U31+FEpV3phK5+l1VAdfxo6aHaEZARFIdh3HPLgfT7pl7n9N6k3Cti
BrKY3lp/y43MILCWNgr2jv934QXGdDNlISsMeo1GyKIqM8QUsO19RqpcC4p3/dlK
2cAMCjJzmUdLG3+bKJ3ZX4pM5xphDB0vAhf6f0044QTzm9sHThjYQiinBgIOLL7Y
LXsRK+05+rzCQkdkWd8hzpvCaRPZHFuVf+esxhs2UTOnsg6iMooM/XaS/ItlHyfr
Ke505b4mCBtseE2NbIHM65zdAEfsqEPjZfdygPHjc2oKpyauZSNZIyZILQvCIgRj
SH3a3OqrtGNvxSBR/TaNFjThrLHWhb1LpixMQydEDXsL3PBwtnlDG4Q2KN0q/Pyt
CgfyupgBn+z3a54JUVFos7Vj5CtArMycmf8PQhQrIDvSUPy1ln1lGNKBNdrUCiW1
btVC+7VLBfzZ4575iPHyJUz4MQT6T7/WgwBqn/ULh+HE8pgPfJ4d9GrNUif5xSkt
/ErJU0zmBXA3wObVx6lx8awvRbmq0vegqN32KsXZtP8S99Uke4bPouD3HA6vi7Fh
HI5gFJj2urnF+ZbS+hBuJrYj7JaiXY+EAtGE/k/d9A7bWKDKuaGlxYyj2+RsyDdP
/bUkT8QoIxAStm6J6DtyYVLJ6RajJTxl+OVoCF/Vb7Yoggnf5bl86KF4Ly12W9jJ
nMmZHopMhQUMNavelqky749Yu2FCyWJ8DLfICylKG+RmI9hphkjWFu+kLJR2Ec2d
DqIw+eiTSCgf9kHu3cV1TbVtzqrkn1kuDeYnpfWReYujmc20bS3dLcau+7GItREa
kFez0YqXCC99Ywzwb9nWfRDKuT4HT0qB0z+Yl2vDMJT5rUWUeEXJ6W3qE5bG0xwH
OLs/FpuOzByqlgjwu5Y16h8mHYd5LflpENmyeQaeqL0S57HDuhTrNgOFIYzmyIxf
pHzsYZ4c9tR4hcNi/1bo0etKV2sAxETV6go6b9WARxgrZm/Py5gbW06iNMZ6TUo4
t9nOod2uVFNMhn1n4UzMkmRSggFIOCoxKDF69ZhtKTrgBYsfhDLHhcEcFMmfHc4L
v326eobWEBVXl3Mz4PfbytUQvliz1mysmiLEJw2XDFtyU+c9pWsNKqe7sBnyvm1M
1MugvbbbDypd15fBY4XnwqJiW8yUffrqj/Mq73FuSiOz681qwFVjZATJVzcFzFxM
Pdra1w7X+gJmxm6/BIAZoBmM6UKL4DE+qeYWvP3780PjsJqN9GV/6a9gxyj4+JVY
7/TLXAykWxIxHWnL5ai6aGxRp4BLJCJRsGWcvN2SCGXLMarycbeb36T2pvvZCwrD
E+vpJii09+VKoAdTPsEpgCvRWaTo0hMSBMAu42tJp/B7lZqv4xVkoTzdrwNCalMc
KW6N884tmLPoikqBJSav1GgHXGJWEXdjtDQF54TGDqBxO/NABNcUui6ZJhcaKts7
jDTA4bigo0YuRfLFC2C4cDSd2z74Wb229LWiXmK6q5yW/enPrjSuEKSCpDJEFVbP
73SM4n6ODnSGJuqFX3rmpECf38h7NrJddF0PDu4JuNZ6HckGQY5gT3DD9JdjcmqG
uL/0KF1Nb559kJFaa1uxyp0rGX9E+mYQNsRm4LEACVFf7hRHPcOWv43Yi+HE5Ef/
4d6zNDr39BaXRcNAGReKkpHk9E3f7U0AGOWrcafJci2DQU22vCvIUyWNoqbZiF0Z
aO3UBM+Yd3gIu3xHLnQ1J5XsUFTZc5WF5FZciSXCnOQtyZU0VHDpyBdQwlhPYI7w
fk6UV6UfOS3vLRAt/s1MNQWAqV1bk2VVQIjZTFWi/USqYcFk/yifUHiG+TGWil+q
pmFS5pOjcIB4w0+0Dv+KdFTE/7qdosym+niYkbBSl03MMM37iLw4eIFxUqshv4JP
jRIwbvbiAjcI9Ub3S5DSU44qhbY+NpT452EvSyIUKG7EsNaeeCy2JjOtPbJ1NZyn
d56DfmkUpitjeSfiNVQ/hWeCh6raXbBlcib+i4dZIDc/wD1CXpRQYPDHj5UAnJbl
vEcKLTR7OtxAC57Whs+8/ns05njpOxlwwVJoK5qCG5nOzbHnUFvA9T058uqS3PPm
HYhXFVqUb9m3el75GH7n+3ggaQk0InhP48pmrzDDvRwKP62fS8bHugELyt3egK0Z
repJNEgs99VYSYK4QkVQb5hJaZHARfDSq0riuY1m9rYF9D22S70xlADojvww0x/P
XTLH3FNTm6bXsRKgdzbb7wE3gMA6CNxdv7p1AQGAjdSXtw5MISX1ufR5fn6gZ1TJ
5m9aYiaENiIW7xndsx8GUUjyMIMlRaEo8/PlOlxlKO4Q579CHttGAJ0SjuXKuf4l
eJooYVGLM1JIgWBiI07pRx8SFdGDFkaMVrtSf77Ifipm60Cbec7i39f3bhbrTqY0
pRuqmX5Uq3EQe0iCPJNsYtPs2mJduphvSeF20pq4D6smco/5hNroxEKBJLuSfVqf
VxD1SBcZwe8B8PEnAQ3WTdE/F2g2oSTKpc0LTwBt/C0qmh3fa70uKNYAAg1wbGI1
7WkP22gQiFC25qm0FrKw/Nbxfb0HgjECyJagsIK12Vc3MSYOATZTc4gzYYniO/MJ
OBx8T69uezuztdujsMGtu26FkbRfM2M7iFaZ0a8kJsFcydcxTwmXt5r23tk3innF
2uWWewP28+zxzvdEbnzlIYdopdbwoHrpmWke8kdnraiCmg0Eoczw/SEEnqGEiNyP
UtIhKfgezc7wBbAB/W0q7Ub3aGXti0VzG1A3RPX69RW4mzU+vgJehrxGCB55B/3b
FlPVc1vFOf3sr4b8i31yQ6lMXhm/1lfpY+QNjPkbunk2A+p9xcsQv44VxUljRgn0
Ma7E8As1jYKbp5CgOopEckLV0mYCzwNsFvbRWVYzKMiiv1gQkgAD7KF5ZRF85CY+
uxp4FwgK6qLspDnFIuVeKdDBMTcEGGRwWnMYzIYcQD9G+zODUG6q0L2llxEF7VCN
ax0ZZBqK6sLaoGmQ3CzcUf87aLMaULxF9/yCdfbVWfNJ2nEEFG3zDb/LI6deAcmI
C8ccLqt2WlZEefJ7wkUscDydeyDQsAQG8A98w33KM8CMkvtjzvPzReIyPk+9cINd
upGb6P6SK4rkZRHCLxLFMFkd7+v/cHrCk9nfPXY/bgEjNMkt0gR/ZJBJw79nTVGN
h1YT0n22fbeXupGw8l+s+QQlm9YsAS3AGLSIX6AkjDqI8VzoH+g0LE+ODy3PHz94
4UtCd4GVU4gFDm8MazA6OP/aj3r8V4uhjkTb46J0STK8WSQ5uiJ78jg7umCduDM2
1KjfRJtrVTI/N6ayd6jNFrbrZxU27BRdw2esoESZvyQ+4IHPnm/LtOd9GTyO5c8v
bhY4JtQwJGT3/qQCy/OKiOFlvpuZ3XYoDF04VLAsiMiRyt5ZqHmm9o9u2X+KxtKK
0ZVCpXDbBGyG0v/zKKigrqTfKMcYTLYTjR5j2HpNLM0uWETwKV1SsD4grbNNYvNo
biYrosSpK2xmpjuN2y1rHdoh3jTjBDDO8cIJWFgAKunXx0+5HPHJJdCde0zmehrz
feb9UXYoZOId3r18VWbsV6bUdzB1yHfCR8SWhMhuxySDRQoTK+zBaBKKmi3SecFS
EAD9BA0tqxWDtDzJCSRxqPQ4buFotpHzHAF4J63a0CU2LMJdPQQP+Xl2k7wt+a6/
rrEUc7Fe69+FWMk0RcnOWE1Wta08SmHcWRdSnkGRFaGSq/5J0o8yaHQ8rldyUXIw
1CpL6J2U95mMtMvCuVcq5LxYTyVlDRmYxB4Ahlb0ijK5pw8bTDYb/pg5GsqJycK+
tNhx9qcYXHUUFzDT0ZvBVFThILsw6mFWWQwO1u033u5HlCuckjlxdsHnPzVHyFVR
TNcVCPpqUxku4etCa/Xz0vIXIQmBbIaq6mT2NZKS1+fuQq+lQNqKedCIx2WMwLq1
Ls9BImBDG519GgwhhNqk3xieP0PRm2djh/z516/4O0W3SoKt2YDS67APqgNMGDZ8
PMqG5fLGSvGeazwVecQQHa7e/c1DxV6us60C5t22/qXG0ZHIZ4XpC8ohw0rfrHHN
d/P18zhd+GvMSdkrA0Jr9ALbeer5BlIOC6+dm13X2gw797y/ev5e+CZI4NMug0r3
y0uOegEc8bTmoKOV0WscnM4U5KXYA0eDML3jzmn1yr/1yez7rguyYBH2i9Eyz4no
BsPJFGs8/q3zoL+7ILncIDJ+KbUl/64NokPSG3cOP1u8bTnxFbfp6X999PeQH3NX
1Mq6NLb2EyJpxruoklDrcBzvFpiUOXnR+va8e5vKNVkNComeBBhY3aesf+Rvet96
Hpm0C5eveg6I20ul+skZgN0RpWONp+1weM5CoFXOCwPeb7pQ8Cf/14TfcYPS1XtZ
Fp0cqxiHCcfaL/q87Ep6vrksguB4ymsQ6nl4Zg+OsE6Ckbjtm89fcnG19VJzP8cy
8UMQbr/rSgrjCt9SXlxGIyhgln8yjIqPGrjbO+BqUA0jHG1lv/9bQG9LkG0+7vuc
7Ga0Kwrn5rRrJcufS0rx4axOibECDdq4g7qVWINA9pfo2i0YnKqBnMl7nj6XMxIy
43Rte52lOVgJ9/YDxPkJkkbH3hYy6517CrDAw2U2fQE7hET1+PHgX320+diJcqJQ
DDbqmF9R4u7DZ/WJOhfvA0e4t/JYFDeOJt8XA6Mki+9FB/gx+0bs8eChFfKiBQyS
qL4KPM+uZ6rSHg/vFWKuGqQXtZBhIWMOT8FJcOb3U0nF0VrIvBhLJlpNi9pQ5pWU
J6a/VGeoTxMs0Sf/4ensFMMWTaYlqWG1l5ZU6d3vOx3F00kcAy5i0JxQYbpQkHNz
EXEZ1SknJLZQYhIJm2VvW0Ppv0mWq93sDtGV4OhDtw9yslDDSiloXe29UI3hT0Kk
QWm9/i4SwSr2NvSr4cD1uzV/oGrpO8fUAGUJW8K34UBDuphNIoNozt4bVuU9i37V
7ypCWB4xsC769Ow42iz19jYYnz6qnXuzmyAZdCKIvlNTkiLBe2tIXD6ibXYo3G8L
HfFZhJFrJBHvfVRr0x/sp2pV1JFlvsqRMxK6l+SePaTirrjJbyV6WeVbSa9d4gvY
JvJdG7gBrywQbqd0aL4gmPh2YiCpP6GG6PV6zXebX8zNI/hUADoLctOfVDlFXNAJ
89DN/1MvZtkiuYOO/FQ4aticjtPbB3wy+rl0DcBtff5lygNnS1xTD2cIRlBgBxhF
Jnn3v+hU3EYPbLDXLEQzt8FGVCiruTHAZwPZDN4dhWUY9Q+7MfoGMkiQP9kZLNDX
5/qsE7lps0aMtOybbYLCbYJuP6J9RnESgskYc3QaeHHLfBmNYd/7nEFmYB/DlqG1
LAH1GchK1ApFZ8hwB7pC0INONwqgtZaY35XzANNOJdpuee3oOOvfcsRPt0ikE1Ke
wqOhjwxTdNWLk0Fm1b4gF5/5cce9DSZdAFp5Y86bskWzS1t9Oqx/3vcCEFMMLjBr
S1cB9jDzGWboblTSJ1xQfi9HkUB3Of8BwjBhlt9xT/ljdV9fOfnXuVFvO9qnPH2C
xS94ZxI0sduXeu+KVe7XyP3vuGMzLmXLZRkaJIjn5xhd+PTWUbkrhsDWPE3taVjv
HBEANL1t/GVgVOkWrdOmkKWC17GWHCauHVAAQmXboI0aNCMC8sU8McfLmfbXhInv
EAqIhD0uT5ms9WFLUxqanKmcge50CXoRzldv73cGfMMHoL7pK3vL/yGPK81By/s7
vNh1c/9USif2umDwy6Ra8MLtN/Kyf3x4E19BlkCFoe/7SUW5QBoGLwjxKaubf8Ll
BCdiFqncNro6kWvdhu5npiMG3SqB11ruRzN3q/kOb/5WH0RdMpB2THzsMuNBoVaA
xjIH+ips7vZ0hIr4ZVxxWB66rURIYU3NS//viFLeJAyM78Qjp9xg7ZRXJ1tp3zJi
p3IYcVC9cYWRz4v+VPtSX9SRwH3aBY5uC+q4/Xqpd5t/Z6ivTUyyiZDrfkhXT1Or
PwFd3KSnh788y04fl6fu+TSkiw3jNR8NI6KNTJMInJhPujxTmHh47LA3gMczjSqr
COHYPcp/go4cMpPor+rIWPgMA9rWWnv5wE9GbgLpR+DKGYaFia4e1ctFLj6uf6/L
MqLPpkBHWP2R1n7MI5UPyBMJB/c1AyWZAbXFsGpboavJZv8upVryNYDHO4T756hl
L42J4E9gxWvl1hA7ppTCxZcwgPdjPpMfOplPq8KX/Y+5koDYmSftKus1WOQUQooy
WeBlSjCAVAvjw7LRCeYF+OHZMY2qnbk08TWaeKB4cDrmik3Bb5M8AmB7FUeL7+xy
k/7leJ+PaMo/cGQXrGJqY3l2zH1QDjKsDlAYL2PNviT9qHlG46Vk8HFKEVon2nSu
/m21spcPGTd18zoir1qXdfeGqUkYi9OSAJH4mRMGnOsx9bv6pi362WpSl/kw6nTt
lXzHFsrVUzQKQyVNkmBpzx9TjvIq4YKYofZrwApDe1QN7JxaF+l0dygMdTmJGoUu
0U5ohN9lnjoJaGz+QvvxL8/8qyjrhx4oN6o7J4WDjV2j4Qk5EgseMOkDoDWAm0qR
Ir51OyqBlHaZ+9mwmilrXxUg6rRRNXECp+tcOq+Etl/xrtuY7z+6Yj3kXmvcS4qe
94pBTSLcH1r/0mF2PqrOtX1uGU8Bw5ewUFFcuau882TeYmF9GanAoTQkWUCF99oy
qch2ivBVmupiHFPrXWiEPTN/tA+CGkBFv6gM+bcu5kKG2GLXqoBpsaWSHDAi1MNn
eFunZZN6vDicMKEhuYnDyq9xni6DlgHMqQP+nV69d/o3yEWHdQNjBgHRvcw2L29X
x6y25PXv4OtmzMo/KalxMtPEEgwoY3kqkIl9x2ZHznPNTLJlRQWG5K/9QuFZd/rq
S7aWevypgXtNDzmZ/yZX9KSpI31DFglOie6NERLxycQweVFL6VGP7ljHuJP09AsE
kYgx6IGizR2xBE8/xDZM0jaC6+JXjhpdEjuuCye9XuTt9swk9E/CRfcVqpMRjttu
AinNzCEyMW1G0PVhlbRQ0baAcH5Zwc23/VM/IV7VfKyspgIC5yMUymLGdfFSkwoO
Lg3kVt2EZYm5s0dSVTbA1hXFRfbtqGEqr7TiEAKbAPDrbrMlSOPWUjPd0hL2qEYz
1yS6+ZA37Kc/xLBCJ8kbw8h8EPLT/fHaFMVu3WfX5nUGaY94iMUZr7XFb1rLrLhF
dLgTfwNoG0Bmof6lKpIZQ2twuX0PrRoNHyZE5Z4KAcDEc57syXzBV0baU6+SoSDP
3uoYTN6KS2y/AoB1K1xifF9fulUifKHsa53Teky9xPq5bhaCYKjbL9yLXtdn8BRl
vmYwOWgo9opMAZkBJRPAiTxy+VSW7AJKr3R3rAEomHoa9XpgZblHPvQxywLooXFO
GQD5oKuCFhH6lKTkZFMyaRnjPyZ89UQiXw9vIw+sXbbG9Q1N0qOUbqHxpOKRfB61
l6AxN3K94BFq+urRBvxtQmai34cGaJ0f4x7QYxXP3i4SznYkAOx0V8fae8yD58M2
8cm1N2gT3WDq+mdaIWrSRfrdI0xi60H5+Hn9HAEX5l1daKb2tw3WAYdJj4Pksm3i
goE4mxHJ4wKfFVbzf/RNsIQxktgMQbl2/R89+5YYwVnnMswM7poLbCKUnkTtIwIm
pyN0AScujoPVMm0cv2eGrqheeqYu0vXkK8xH3kLyqDCLnGz58VJRDB7NNvgAs6Pw
7CdKOz/N+QHqDeuoN4VgpYMqwQb9bziqsl+zgYlJxODNFVbn4DcT0k4CpXTOW/mA
G57YhsCvY9PITor1bgujdVKiFLTPh1rwRjsspkYh9rj7UEMyGuReEt12qo66fRkO
7hY+Z4516lPEbSpw/Qek1+VkyIRRkUbamx05l7nYPtdWkKj2XWGYuaivROQK5CVZ
7v//4S0mruXPQBJMh7cYWYYQ/FlswluDHfVspVKG+kVpm8/GzII8gFsp49AfuU0P
e3C41jNXO9xAixQozaubbpREIRpJl0NBsGWNleoAyZws9idny6Jb/VQJsO9+PzE/
pjBruzhTjVhFIiahF1jGefPP4/AL8bW/cy4gnK/ZVU/77lMdVtzNjPouepAL/BAF
rLtZEGosC0qERp6RjlnZris2CcBqczM3eVyz5N63B/1gFobCHBLSufCqmSH4XS/2
y3QtXcdmCiN3xl1q2hbHARB90b/thUowML8t+sWXQxhePF2PmhXwxxFumkZ/H4JK
Q4oEmkNGha4tegdwbXXMJEyybSyOh9xJoQEsXa5bvYFAhVX5P0cqlzzq9dst8bMM
+2Nu8Efg/7ydrI3HddmkyjZ/hlV7EBliV1iS1dzHv75ZyzcYQO/m9PF9m18JzYJe
37KmPtjWjBi3cZz2WXhoKJa+qY81ytmo4XbQ+/uzLKafyvgP+F9SfLXik8+j90ow
L1Ro+SfMEVKsmAN3VnN+SQb5sMlqwyJtDRGjbhqFZLs3gRo8dJ7/Nj9CQxJe+xyU
fzyX7cVeoVnsBttUJI1g23rDDzHtEkr8nNTHNgYnHtDPSizAwfUNztKpCV73TV6b
ItAaRmPoYKvOjRjdXw0HHIfJXyHa9TThQgqhajSkkvEEB1qVT4goDs42uVDZ/SqU
NK8WbbMUF4SYhDUbzwJTb6qrEnyVSYeth7KjMQL62FerY1BnELdX8rPZYRUgZZv5
+tNKDdOzM8btPouDxqE+1FujqkSDDOP2EV4EC8wWdH9yjoDgHulS1Cpsh2RD8E2B
8M9mzDys2vSQX+JOYnWZ46hEgEtsxQvGGV05DNnLalFjVUnUkPTo7lu2igfN3WT2
mbTmgtnKYgrVJCNrdpTMSsuJFWpb4A8k6UNOQRQfh7/HVpPqUycJMBmot5aSyMqR
/ugTWJd/Z16H4J13WlxYaS/TiPn9kmFexIS0vZcxtWeVTyLvvuL6ryCqtVb9E+O9
y6MllG9klTLMOp6mHSr582mLIkSs9Q1TIJn4Bn22ZbP6Ayua2U5/oUZjLWwtDCRB
ZpSjk5+lHtMT07bQpAQuEhkUN328Xu5KopRi7aUCyyuQ0abmVyGzvWZSk+e9Qmq6
SibDlW8GaFylZ48r95AzrvpsU8DS1/YiIXCCsHCXqlOnCrw28DiCIABlRzjf+KIR
n3kGXXxcn5lnuvo9yXW/3tU+fZMlBr/Q1QqUMxHcj+592hAihZs4+1rr/9wKpCCk
qON7V+SLB4PwIDeXpTlx+D6kFqgnU308Mb0tZe/+A6t0C8DJJCrJXsrvJdtAwqtE
d+Yr0WL4KQvpYB8VlpW6OEqG0Y/Q6YXaIOjUvPNBggJzVW7+VsonOOIbG6loYw5o
Tkf4o6oUvNbLWNmPQS/sYCCpFHh6h7SGS0IHGc9HNZogm1Xsr0Nk3DcSh+uu2NNZ
9OZnwtZHE/k454C3bgRcbdVKKUd1CmcnIZrb0vRAhaJljxmvn59rRo8q6rjgb4cF
Mty0+u1PEQWHYW9UojVn9nXgG2FXDzyKnm4+v9NJEBTF1A2rv7uufGJ8Z0FfM7by
rHhj1mPflhtyOAb6ts5Mk35m1Kelh/UnwC5FE4pqOD2lxDNTY0yoTvuKNximMneB
pWkHMUWawSKkBrV25/J0X2gJzBopCIQxBvWj3RNLj5iDb2/8eBs/Ah+3DHW/wBes
LluHCI6xoyCecrnlil9kjZEQo98LapzPq8IC6GqScLF2bOsdeR7LtoZyU6dtl86x
ILqOtUQfhcUZAroI8lZMolOu1dIlsUqgspfHH6C/C3UE4QNf1qxbNgvHIaYcFYnV
VTXVz/DkEoIwX5ixJbDeWSEa9qlVi+ow4OpDBEEu2XZ2jIJWRv+wpXquh36/T1DS
jokU3FbMvND5rpdz2nn4oXlxgYuNRbCuDdJxknzvPjb3T9tn+DBkdxefr60Z3b+T
VTlJvuOg4UeHsNv4U9h7n6nfXx8Je+1DLZ/9t+HCeRZ13Emeu4HQOBfLIZvtQSX7
KlkvwBNiyIoi4nHYdW6+ui7oAEtCRga00ivU6k8UNMp0ftIpVJu/87xfLMYBTS4D
g/pmKR4TEUJExtaeqZkbFEf88jFVh8Hp2BMhPynGO+OrohC6c72ZnNfHIygIUabB
gtxxZc1qWbhWlnHGE6VqFuNF2mrp9JOLJ7eyIlf+e55OZzdNZ6T66wE7nbXxtroH
ckl3727nemj9Caepw608bj1m9+qGDTogYkYLeLXyDjYZsgsYAG8KwIhO9qCHuvfi
SBlRez7P04JSSAl+V3iZ9u6ZvhfT2s0BBAPOkVMfMWR8SCAlHBi9WKJR3iarZTZL
myJ49ErgFzNLBPBcWBbsvdkbSU0Jku3Hd5jmh+EU3afeytSvYhHQM0Qv9var448q
EZ0hbBBT7TrN0svvBXSVfv/7CoS7daKw+bCEdYdMw0Y7dgAT3vWbV59iSiluxKV6
CgVqomDGOdfvroFyPaz68Lx6JnaVmEcTaov4yWqXXrFkIb+slvCzV26/HOmtXBwT
HGDLhEFAqeHGkla0Rtz6uK4AN2WIo1rUjNJwxJvr2FqUbeBH8hmYoN28TBi9WYyu
jUYdym6gh13Yd9xqtU1IgOzByU1GGFmMPw9VlWCqh7MU3MUmcqpuhfAEfKvJLCcz
3CeTOh6AkAmgFac5kYWc+HQ0fNT91L4b/R9NFZpgHdGZjB/mjupTf7f5XoCPe+9M
IbTAo3p0g8h5zocvLqdrMPWx6z9h/6K0CL8PCLBqGmD5rAGN1vyPSYtKwAstDU2S
1D77aXrEOn8q8bkQjL75nt4X+WEkavi+jtmUW9wkzqr5+nzXRzXKgOiPRA7wcOn1
4xnKe9YCFBFN2WsGCjxj4NuauroXZ+xtYYYsu3Ca0XwSHUeC6bO5F3jYMSDbIMfp
vD+QIj+PtGuRSKW/PeAeA8qayFKqa3s1muNFijM9U2QnUP1138LR7BaS5E6G8VXX
1NGZjNw1qfK8Ka1uxcL+py+Jw2ITJHU2baKzReZbku+JKcb0hUO2/kAkjppJ4tlU
c8tQHVs/boSGNyeCYVXajSdTLv+ujXvcHIhY5s+49spSfqBt8g+vYQemFxaWnVoO
oKJtLulP7zQJTQIydfErXRrc+PBZ7GN+0XLUofvDvqp3ja3DjX7BZOWMfCurrUiN
kIF2Odq4rTWHzOh/Pd5NuSsp9Y1UN4QGzGSOtGNbh1BZXXcY/zP0EmDGylBzJMoT
nNeW47s14e8PP7U2JWWEovO3Bw4tkyFWGb+97Eb82EYrOkDkvyH81jeqBlyr3RTh
A7fMBkq12E8zcvOzbX71DwJ18QU68S75xoN4qg31Vg5dRvVDglp5eqSFbpTgvwrt
xyPqqT/qbe5qNhg67Kv9++NoIws76iIxBSyyxOosjHbTSaG0IivGt9MLnH637GTE
nxQUp3v8ayKMAxX99CISpeah7qbOXSvd0Dx4kQKfMxMoFrDXwQ4FqM49YyRqYzw0
ewgpNtoVCCKNg/F4U8ghUby9xAwZJn+FePkQI/i6WG+xkjZwwyuNtgwgPGkeHIh1
AFJ4Xg4Lj33rX88h80FdZ8YmSmmMT3xgTcwvU9wamI7MIBfhuQoYWGNHLJeuOAlx
AUfZwDV4iGr3t58SB+YYm2NhWDeH3rY4/zTS1kHsjzrsuHGcoKXYOgqQ+R1fWxXD
HfHpretNwr+v1/nSdQmGUr+nFQYM8mPaSYtlWhMHeNNtLVKtg4ryzRKXViLVkKDD
1uRonqywzC19qMQEtlKUs+HDNazDh9lpbC7/5k56hNe5gfO+4gVZxlHBUP1kuBqx
2dYL6Vy7loQyPu/zJKBrAUbKzyLpkXM56FmWhpKIxjYwxpvkbWsDSGS71K/j4a5r
OeX2DeX12nsp5v3TZX9UIMf3lkybL/DvMrAKapPtd9HHDU1St8ByIKFtkAHQcHSO
q+ktg51iGivT5qk9Z1CuCJwpRwHN0L87t4FRiUGyMH9cT6Hpib9AuSTTFkK/Lpsx
8TkfdUlljQDCS2zk3AhjXXOv4lU0A0blolGkVKBFhtLcZ6jifcKy7M2vWO3Fbzzi
0sZkQfi06LWzQ76ocAqOiRljGZSQeiM3j/Qfg6Xy/i6oJLj0u0qtftVgM6ZP7d/s
IPx1hvZ44hCShnCYMPi5sZLX93MWfBL1mQkuqQS6Twjil1oTrOjcD2xEvwTTS3Z7
6gPs+sThES1pYseOQCPqCZOiGoorSTIg18jRheCLN8qwR54lEAUoz+8QKvMr8vZ8
Pmg4E/OKp8cO+3ioqn0DF5ACNlknFE8Hyi12297eVHziILkx/ux9tN8RF7e5w5iH
n1XLBiUbU8JbAOsyAp9qx3Hg8keRE8qxSzh3ZYHDDc300K3d1DnN1VfeoMUJv/yi
WyZIRCULrNETbOk9Wq8WhDthBcQau9rYhohL4oPPtXhpGAVJNMxeC1Hums2nmjdh
uRgxFMuQcv8B0MPXGz11HUYcubh2kQcTvKp8Pv2xz+Id7Wh31e8VlredQ6uQiLT5
728pg8R14S0QQvQNyg2dVU5146ERBvetiTUkZpTa17f+JDp9egh1ucdL1LgFx+gw
xXc0adS6SFLD/pJE+suGjKhCbMsIpR1YuwnPjrKZrL8pMTlE4ShQWypz8uOJvmMq
+QQreUh5lO7/r9eZfjnLIbOucg95Lom4OMiZfIHZ/NhpBO7GHYRljphX2no9y0Ru
e9Z6jm+AwIg+mgN18YN3zjwNVYYTP90Jxa6eQEsF7o5TaSlm1DvEKvGtFttgMofU
8a33OP3Jm8o7AJopBda/CSBHpbzBRaLytXH4muhKAL35rXekmhfGgvHKySBfPEmx
jzs9CfmbszHbboewBJEBS0wyiQ40ACP8MDN26yLkaVGa0dKe8TVimty0WUNtU1gT
T3Of3Ifsyf017aMf7Od4VpvM1VcgHH0XG7PuZ3EOvvKRONa7dnE0jfKe/NxB4r6K
ViI/7A/8QHNkU3G/KzpZGZNIDAG4uSg8WZTG1IdygU6ac0ntD6r5gOy1c6rFFNhR
yqOHUYoRwOESThn9qe7vpTUP3GFriPaYkeYGGpIuIjfDQBPL+Ys+OW4a6tn5j/Lk
rY5G1weBrkOiU/AzKGNcT0ftvaZH6hg8RVeFu8mU3850fT7FgOsL8WnHY+eSXHjQ
E2hc03X/Mx0ENMnrGOgFpj9zWOXWMT7pGDL7zOsXw9y4F/mzw5dvs6eUWLbmGzea
OfsCnhs7OVAQgLVCkHljAf2ECG65YbtQ4f2Ddkok9Bb4ab5tRFNTToLRhnUt+yod
d4tnJSoSQJ4Kt3DQoTVxBMZvle3zpFA5PogjyF0JRKwO7z6NzJWZXGuW880dQKIh
rmm5+lAeB6hebNaT4ALOPRppJx87ubNd+dEFqdQjXd9/dIo/ZkmIPfhu/xfQbSaN
CtvNC5f5vccc8MOumnAzg+ccOItL2kQQim6UifPtNhCRg8CZtAHE50C8qZul9dVz
ga1UpsReFtFhXsxwVBwnaGSobAqP2ptDUiwhT7mD+2WkAABfh9D7ESE4MywbAlpG
f6cNx2XbHfLcOG4VvrspG06dwz37SAbN0PuHf+TFJQibs5yIltOat2TotDKbzspU
uoa21ClKZGDrPqKN1zhTGHiubLH7Zbn6q9drwjJNS9sQOadsiilutbETYHstW4Gb
SlU0RBk9F5It6TS4zrqe+sq2urhLqwh+Quock9M9g9vj/pC4qkJcHJuqp2b1MJiy
VpBOqsbXH3pr7jXRRP1oZSzfT4szxcdkMBPcgD0+YvSSuLIca7v8nOtEhx+wW4Uz
w/IqhJEuiU8zF/I308yJuSzqVrT4vpM3QXudeMoBz64e47SeV85CuYfd2mxONOCQ
XSGeNs2kc2kGxUpB0qSx839KU6QPwyg5iIjJrHEI9T1YYEGMevTD7KnLvYi3az4G
TNUMF7unWz3pLIGH+YiwJnzeJRy9cAzO0gS6UnaBqLPFvLL/Ck4cBk5T+icHxCen
poyVg491fDZlHISnrRxxxo2/fB2htCupJn0F1vuTP69nQtLTOJRBBeYFiMdI6ZUc
MMVC0tlskUz6q4h4T3HZGF3UvvI6hS5+LiaVjAoYCgKYsVccXD+5zYgQcsw75KPn
0+BxlBhxb8QEinGLnD1laE/oiIPW0pMBi5VrpSH6yKzhStfjFXDgThdLp64sDIjp
opKHkksMVWreVkGPYjrDISkDkEKV36RrKbkB6WgQBiR8S/ZnGKvcNsOJNMELBr8+
HMmljSf5JPPkcJTaL8dPbx+qKJa4nUqH4RKRSFkK6cbJNVLr9dWU5OTvBl4z7qYw
RRaOcRJuVrJQ9ZNgZUcvKq6g47el+P9qRCQ/M64Rcrs8hN/YH4cYUeXEYz1v6zj/
Lci1IH0+B1RNtoEkxOHmK+kvaKuGAcISJfkog+I9MJC00XaIFNYEUmD/WL8IlSfZ
3OoC4KcAYSHx1zJAlWmpCtpyZTcg6zGk9TfQFSMDgKq45mwY5P1Pp64F+eESyn/Q
speGFxYnLVlNma4d7FYhYZN7V6r562Ku39+Z6vU/zNZ2Ajz/UeDXJinwYSJznQmM
4EXu0l6nLRLPBSuprIy0y3qCY2WnFE0DGlOtUSu0MgKnt8hQ2ghsBy7zPwLxtdAu
jeMdZtpFyi7ahOp3ad5LzAptnjKuIuBwProyPxRKKHIOmo32NpEF74tAMWomt4ci
6SJVTf3hzTsZq9Dsia/9FnvzzMzuijrdq7KF/iXs16fokrrW/6UksdxTYo63+qNH
z2rJPzynvnhe38XqRDODPav/D7enxd9WLCqi4HzDnQHPqzKqVHJUwdKoF7woM0aD
YnT7EjdIMQSJ2Jh/7UMLqa3JO25xC7ChGzmOcsWEsSOlfFTExEB69iPK4jl/jkK5
8kYJx2F4uKBLhOGnAunnYvgdVVf0jNSYTD1eDwMspBrKROaFnjOgmTPBkvHRzfvp
3/KljC3i2lY5f1ZZG/SzCCiYZmOC+5E3dn/reRitPc393nYmTWeJrhi6eV6/PGsW
xJ6KmUNfSu7adE5Y9Isf9wl6SCjw2odPRA9M28pZm+fYje57adf/160I6W8TPNJf
RGunYejGGFWhhtpJ7x7CXofXSvZAqjPIxIaC7W7JEQ7qEaKpDqWIBVNmmvqgt8YU
ld5an8lWGl3PswsSqDqJH/i5ViLzy16wJvq0p1ryLZieV2hBzgGh9gtFcsYQCjmN
nwjecRn7/AU9q/OVV2nESiVKH2iWVI/0gdjSOHIrkS1bAhkspg8g0VZaf0T2aq/r
jI9MuLqvbuiZojrMVrD4gIeQjQ9Nrzb3okCCopsUpiEqxpxed8N5D58nM88EWRtk
5v+Z+l3zCdJlgcVj6fcBJ5p0SApC9JxmjTOQjetiU1+s86DarTCzQdz3PZuJ3z13
TiH2GeeeYC3UQW3LltF3Be/o4AeAukcuse6qckEMvu6qp7jswPZESyK/nEOY4R1U
etgEpJN8WxZrg/TYBmIaedK5b/yIgLxkS9/7CXhtlrfKFV5Ur5tTIJbVyYdFZ+8K
uyq0TdVfjsH2t9bsQuB1TjGPwUBRxc9dxWH4KIwt3T4TUG/5DSCe1dfLtVvBrzLF
H4GYoZqtEz1T2KRfQ8d/LptpQOUdfkjZrfHDRAqRlDz23fkRZZf+SyY9toYY81ER
jGBoJAIQymTybro45sctSaVo6owHAi08P7QEflUpui2amxryHjrCohS2NLeEbuaK
z/VxGhB2KAi8F1kv9TUlgmj2LH2ZQNl/LyB2LI1l8zPCrjaDMZHYzfCChLN3SZdU
ubcVyDZ+c5NBg/3N/s9deacb1RpY9+q6N3us9gXVBvFwcZ9RMacf3xEgqZYmxAg5
8Hip6631AFVNmayQmQY+f7agizAn3OaLwXPoPwhwqnOyHoD+JtG7n/+hTNACORfH
pNjAgC7IJ7Hqi0BJZXT1FPVnOOPONN5s6lAW0xlzfFcUFUY+vrMwnkQ82Bsmd7pV
EXqv+ZlZr+e5/feMZdQIAZ5dLFHse84Ghr6rfblIuL76YJW5vFCHKurCE5F4kLSU
oPXFdVQIiLx7KEvyCtxEg1G8my/mP5SZsRYSUeA9ca1TGeKEtQUHG8PtVd7xWG2h
IxSqHNmCM4GzBoA5qL/IFa/ezpfnGAlh+Om9pFp3F9FU/mJ6yE/7oCnT5STWugKZ
SDHHGh6iizLo3sOoOZiSVT50XLhD5MQ4JGb9EKul836dA7uC2sgqaAiF+JZkKArT
iRj1fjeXyeWoAlpWRuqOxHMMYk83qJyCFsWv4J2v5l84RZi7+J8fm/Kl285rZVcX
Ca83xbK8Njj+aQEjmoDPR3iAqpgOzEqtdCzwDk6zS1F8TMbwF9Mt/3GO3EhPpbTP
ng2owIOZ18sEz0ybp5iDudaXBQQvZ5wDCocy3Wy1c/bQ/WlmTcOu+L6N9lVFE30I
rA0opyND1UXHCgQurr1oIloURmom987uBAva2BAlWZArvvAeaKhDx7pZuQyEttou
Ytfp4OANskYuU5sc0x0DUjBW6Wha4IoKJr0sZCqUBQkkiCaeCq88/U4+SvbC4ldK
Y3GznwUbX209qVk99u65lq8mdRG1I/0ONPEVhhDbDiRhwF2Vj0l0BBDEQHmLRQIb
cOjQ9FO88lYq6aRLni2vqSheavtNVHdDmeRK9mzXR2EnHtXXQxjVOrWy9TqaPVfv
9QvHznTYOqwUum0lz64Aa4ttXxIGVM4YjELdM7Vz1RLV0nBw3RY1C3Z5uFMDX0QU
n1NPh/nI3QeytRYu/XFKaF49F/XcvtWupDqvarUu2v3lx3eae8q6qXXYboWzgPxq
aXoKo2g7aGEemoYkmagdzS9M/DhfoKZxKRwj/VNtV1nj2nG0f1P7+MX3I/16H3nt
ICD2aX6PAvlk33wkM6AyBjNHCvBLgVQWAGiYERPqH5hj9wFDaM6eyiy3WmY5QRQj
XlrX1fWsgJ+sWcL/RKenHEhq7UFYC3jJ57ZvhuA2XL9vB3Mrlan+w03uoOR/BqM1
s4i8GvpUsoTfzdb27nlhbVekzqexsQqE1VJMCDRjbliCrdQl45RqYd+u26RfKLv5
XGWd9k1wwNCyIRFZY8Cmqn9Apx4TsidXHoGEbTEmG7sAX1A99f2ZKfUUMhSp0Yme
v6LEsvqrtUYjROvdzjLwdkEoQqEaMpVKtwMw5PTKRIVnb2uficjzzl8lc9lvkRUi
8WhbBFgDhSqe23FwE6vh2QZWbYyVzBEn7Sto6r7GQWt7MRRud0uEIjdqJ+SoqhYS
bnpnP5vMVGk5DSYwxDl78frcDsfLtSWKiipacRdKWxJaV2eklvYzFVGFrdZ4ndiE
L12/DGZpdzrQQgXylsZNDkoj++pJVQ5Q6KtkiLeZfL4WjBvED8V7ux+8B9PW3xsf
m+0Me/Nb3yCAvzo6UEGnYpHcyWRiLnmc38uAyzDtjGZ8gK/Tw+pAMAGVqGrK8/pj
rMyteWURW1bzeZiKgYKyzJyQc/irfxqD+r0qp9c6+krcZ3kRHWaSCP2r666J0fSD
p4rXpVDA7dFInfan4bLI7AsE7rNMnJIQBbvhBOGiQynLdGjJVA0hM7KExOTzryjj
NnDnlteB+gjCFL0SUgD0ZzjyHUw8bQXUMTKG1a5qDNP7olmf39qz5nZ74OM3Y2Ur
x0ls43hE2he58fbpNRNt41VrxiSTgbpBtinkaj4QXnaP6gRscoY+OYYaV2krApQR
euzo5/RX/N8ZAPSkeDYrgbAZv3pgao1rOjZYHt9WA0tPbvDEd2xchT0V3bImvZxv
s/mLxnJNeT0It+pzfA1Pny/mkTMsb6VGriedxT9UdFCkxcb0E3g6xslTjto6ZONW
UYJt6/2AubinkuRfNPvc42nPzPqTI7SWd2nwGGyQo9EHnYmKOx9ZtZ9l1J9RQ5Ty
YWohifNo0viuQOuW4vIi7E4x6o3OeDglzyb9XcN/gddRqUU76RSPrlt0wpjt+mK0
gGHIRb3MBQm5Ym+0aYV1kwAzgzFk186qqRpsRNlWbg+IEgYx6u5xFCsjfXW14fjR
7WT/y12RoN+3g5dtqzgTlOiz/RLjTTm/165uGxt4Qv8PUSvSZtK+3zMm3zZROF5B
sfLYYezuROGpslvAPOt2fm6HcjR76g2Lvvlwl1tgDt5WxC2TWfJNiTtZ+GRlP+q5
aawHZwVwK04215Z9RhdS3PxFDTOb4R0PFrGXmf5h2RllMw9sus5Io3SRYZCCivaI
hcYUfCyax6nm5vJiT4hvwHzSlfdf+KRahdeLHnb2JgUb2yEIxNpuJ6XhfyJWFY9a
HAJilgX5GBRytZ3C3BP37GdM2tqyAywuALsxwTsnBPsUzeoDbjr5QUoFagKfwOt7
DjwAiHX6TLIWgEsLK+fpdRxRICQOVuicbXMuBWrswv4vm/3D47p/VL9o2qOQY9Ia
ZXefCfvF1GlAKELqo6dFJ59C+dHC9ZUywb4sUwxg+fXal6HhSvEncwMH2kpw/5BU
EKS13L0TwLyFatld8W2mm9LpUFng/njhFpI3ty2CXDhGL8OGONyQFiJ+rqp8XOuq
s5x592ZPVpJrMHzP2G8muGFq8sokIfrrLWqmHrN4gw/GPvTueM7mmREixAyi2DDK
QiliWdJ9l7NTSw0gusryI+4XmhIS8RZ5GLAlLsr7fFDXS9CoZhL2zbrFmF66Sqiv
ziYzIexT0YRdF0JCmd+vAIE4QoNFA5mLF0TrjRX6MS052X/Up5s3OG9zec9V7r5c
8+3lgAUnzGOqDHudkGWOiJMKAUAdLsa1d4Gb2Nzt2ZXLxdkpS2ivCOb9BUJ7OWO2
UI0SHn+YakLY2zbQaPiTYqIEbJdV58LDqQmxhZweCsybRbAztPPAxae+JNMmFAwO
l43eVPdOLSk6ASgXJg6CGyM/pXdPyj3pJ65bqgVMtksIiWB2E+NfDJHIIqqMtfxe
YIMA/g5xQTkSe2UOjysu8oZwoIFGDpkYY1sxMX0PWvge2mWYWZbX8wl2e7ZxHE7O
EUgLm8ucMhFoqJ0qJ0W3voHZmQahIa4cG2bidMPcEaucDauqgpoCKEEgC9GdoC43
NBgGXbsRJ0XWQC6moODsZrPjN5zSvKT9A/1lbk7uAqQ0M67n+qptaUN/4IxxzXuQ
6/TBxvFejE24F/qRS6yTkjp8qP2AkufLVNwlauEUwRntW+G98NBmMyEPnaSR6dzS
JVlXXVhVlJnx+WicYPA3VuOAQ93DzXVoyonk1QOqz2EhzkkCQr0vbs7rOJOxLyE1
4jN6i2eDG1eny4g6K0ow2qj6uAYzeEBekGdAlPPqPUKnBsaCfaY9w6PPJ8XlWbje
wrPaE5XNR0FUuFg8jEIInVyvuSq2WAy1yMomhOVYjVe/MWZRdreMdy8mdN1jeBR2
rW+Lv8fsJnSPlv29QmAl1jls+zRiD71fVvOd3gTVSvLsPqpZGeYIii5dpLoL/Iy4
PQdDtQVJvp07XDlhOGlT+fAY1JoVdPnVpClbAAl6xoS6ZwRwLyDiPjUxf5IGF7mX
LbyMACXaXn6GVvqeqC0ywXBgb+1EvPEUMrnZIBsbT3GG0Owkbf4pJFl+CgKhVOH6
YxRF9NsW17pV1s983svtaPrF9KujwBB8eMyzXXTPlEGfjyh/CkjxbvSCbaRuUi1i
IRZ0AHJX+RGLxqxqXK9CQOsQYTBNJfDQTVxWzRJirjxhSEUjN9nSWjQ7zXBGrrx+
q75Yx/uGX4ZJL80mfxjdV9wX0EJmHIzIbCK56UBsr00etc+Q9OCP0CwGoSK8lAUi
1R5ezWwSW+vydpGyWilb3n8/FMEolrdw11J5+jEh278NB0fLR/5uTJf4r+yjJSdr
J0adi6C2bVGGazVGKgEcA5+WQQWnAMEs+QKNOQ+MlPd7OL2Qu0QPKgx9JF7BDFB7
h+8Zvm2K0jxZKrlWfToQEFy6FP1x1t7RqA2nTZqDv682OMuGyG6eCOYdJOepJUaE
lZpaBjXaJf8PRn9k8PP9Gbswy4WNbKkIQAVe8rxvEUiIpmPszE/9og1AxELDRIJu
vNQpbUpXHgDnTE2jATQiha+A3v87GoG+BTohdndvUTuFWQKByrinK4POZIBpO4/r
6MsVAKFhXonMQv/nadoQ1/4Ct69NUR2h6262qhtD/kxNgym5uc+MPN5g6AMH6tyd
oq8gJ6S2akClSNAocZfoam4N2WWyqP/qrSX8PtVdaThc/KwBBhKLxmcqnh+DqNoi
sYe3b2LKjMX3DRDd2K6S7KQfnP0BitgBiHSmdRJL//p2/PQzqVFMRfkUwhq3MUam
Jzi2kgKcHQ/tAe9+ppzpjWYBnls4PEiXEu0V3M+ZdDSnyGrpmzYT2hsrHM0LRhDz
TZNS9jZUrD2seNEcpNzBzX5VrvYZ3GbzFDItzXGeOyQKN/lAmQVGw30qK7DzSCpH
IUTRLWxK4B3pGtmNqnQlOssxY22T2fKH5qpPB9Fzwf6a3Jg2tykIUDqGRoW4nZ94
oHVPpBjiYZIyqN09AJjOEx5elSGTCXkHnbHYUelG6XTwwB4lDx9fpO0NStyw/PBz
JVHwCAe5V8S2TWYKLpJNf18JTijGw0Gsrfl83YL2QcMsz1STiW8G/TMOJ15dAK+x
Hjuh63VOaRycNZ3wuhbDZX5OQubpvjURCB5YdYfJ8Gzk1jWOyJOqOry1Zd55cSuH
LTkbUDqDbG5JQaNxaZMymC3CIU8Hd1PTLoc0zOAUg8k99wRaLZfki1QSuz60lPb1
IsZDtXnJ63puMqYTSwrgAFq8D8kaeigAQ+aMYVM7uUZQvKcIsRs4vmjOmpnRhTXl
Y0lIdZa8bf6j7krQemKxS9bDSAVSiEuv16c+ranYy9gCnmMLs01BUe6J8H4tx36p
L/onPrUY6G3FnTVW6pYkiJrltHwDD2h6QMX4NW/+RO7muM2hF1VwCYusTVlrvapW
cKv8YfP6IHGNAffmm6aK9zKOyNlvORbA+DEedUbvhy3qaEVD1tq/OIU1f4HHY++y
ffY5ixmbCzC5V4+yBLTAEUVGI6BHIqobrhM2bqLjnf6ssjJNn3EuXWPce/JQm7LS
k8F50DERwjl3B6B1ljXFaVCJv6wrRatkkqb0FpkImzU7llfbOdGh498p8AITuiOd
ina2yAgtfuZXBKXoDOExXiqBR2MMYHFnIAYFROYCxaMAairGQLWg5sXIegAWRsCA
/Au2zElWIjzAuVsiMNm3t8xYdfHVEQdoFKpkqUSsToO7F2v6vWZetmarlGdHcCsz
qWdbr5Nf2rQS6bCGQTehTr8LtxSG3fj2tSkroVD30eJW65OUEyrBtBGlOQQKWj8U
ZcXMPn9/mYO/fH7/lN+UIyKZtRImpIhBdKqywCS3QQqyz6aztVsw6ZfRZiwNFadJ
34Wusa90OQPel7KPhyYhhhwJBjbwUNQ6TveEqMfmywUE/7RlEhc+EOUBQeWWlTxf
KlB1o7PfKJ+ayuUaT6wuH2uBB/kiNzDQUGTbFgcdCwjtC6oyeMLhilbz+28bS/9M
K0FwMrwwrQI0FhQ1OZEc0cEbvcl2anvlhV2IitTRurvGic/JVpENEmAjm0a7aT+3
UoE+jAEMhxZrFCNQYxb0IwKQgaYicUgP9SfO+r5iiA6m5pHU6CFrlQ1G5AlKw2ou
3/R0f1UeLmvN/oe25MMy6a6tzXEbXE5QSr2zfNaUTxziQWcgiVsJx7jS5LdrdmE7
oFMVRJqTUltrAUUbN0wTAQjQSZskkqr2mz3N6XWJYtFYPXURUeqQJEUBhxXJ5wqR
/HqWJE2JPriq9SqOZbMWOxLB/XBhSC3pxq8kDFVtq0dmMi7GrhfCM5/BfQr1RNU8
5eCuQMv3S9PKhXKXkWYCj1ctHn92UBJCoUM2pcnuEAvfYu/njnt1wEnmWdoVDfdm
YfDnmaBJqs4PzCX7FVQxUVR8f9lit8R74mEZHT3QU4npIoNtaLvkSI546jq8VFCu
5F872OGL9ZM7qVKuZ9HL3B31UqVGpX3qPfaxcOKi8ZvNWS/cE4+BrBFgbL2bR5ZN
FiO9Hce/lEUAXSFUUGlRk+dDJtCigtax0aVsANgvUftMps8aUwakaOvIuZHWjysr
lpadXnzx2nEs/Dn/lSP2HgOgfsA8omkDeiwaNaRqZykGW0vJgqunAuvg8ChnX5AS
AF8hAH2EMz121IRqepSbED0yZ3ilvMokoLmyqasBiXq7N++YiZJaVkCvWd+cHn5y
rGL9oMidNoPKtP1jRSAl27bxIDnqbzBkKjnXgKc/ut/KICtc6rKC29XbdElSQw9O
GWyhmHBuvDliAf2babOJ9h7d5e6AlJfVN+GjyYa6c1V088pf7rh7YXFZD0lDkzYI
DCa7jMxtwM4xyB63k8M5kpYLVjFZHXPZ6bZyDmTxwXFQWnMtrTx9TZ5hcApNgdXR
/6g2m2p0OEkN8IgJHq5Wk6uA7df0eC0uw89bclYAYv3ifFWtGeJk+uDcd28ETbzs
HqfYP3pZA25u4B4qed7f+BXW1GR2DGKwuu8NQEJkDRK16ncGRUduPZoQrpueyQMA
dhkcNzjjMdMLaque7w0qhnB8uZo1qzscb3jbGSgGGem1i/yv/5sNhZFXMLxLn++O
djLg+ckzGaLkESWKjSxQoJWQu/NYYeKQqFmLjnXDSDjlEmZDSUxefAU5Zq0QtQwT
4KwMPXEWGchTjOCgANqlDQon9MC0l7lNOanWrur5poi1dOKr1Z4pH2fJvKs92/oz
8tZFf66dhvIdfN7FlYw4jbC4Mj6uD7GreIJ/i+xPF0tuBeIeQ4/XPN9gh8JAKT0H
5XkI5CHEJLHbqfgqtUthhymquW+zAzfREHQlCtS7ycGSIzpo786pjzlgMWTeN1bF
QpeaJ1aXxPwEu+dk0nsvkiE5Hv9WgJRW9wQ1tnGgsJa5629jJ4bcMtmPEtVlOuQD
A/azII8u8VIVBtFW7zR3hiAdXSq4CynLl0bGrZzNHHArwlICyBSun8+y79nSV80E
rHhXMUr55en1r4ai+xvIKYYx3EQbKBx0GrFp7mBK8dvYZ+kdePxHnNo3pQiVvFSd
l/gkrYf0/ZFUWiTYlYCACazhYuoiXjHuc+Cxc1eeY0VmEY0LY4p6zTTIN5XeyfNo
A4JvwqyeTMrMrnCbiYwW4YyDhXzsRsJ47N26nP+6KYk1ORNuQjyzO4mwFAgcIk+j
JkLGPybOPCYZPnnxWpRTrfFkKWx2BdNI1AIE9il2sfOxg3hWU4qQX6RN9MmS/VPo
TzGyBYFdY6bNhf+9CZ3hI8QY4O3fKiC+XvB+WlUJeKrYbGqcEG1kvndD7Ca38ohJ
4hsRsVHvSL0UnJ0g2dMcgyrSMNeaidLUWMGqneRBp9UumGUoKBqSsE3d/IDQQ195
r31Z9tjJqBFF/BDuiaqcINZeOSku/kN8u2qTlUJSWR669J5GyqzAi0zBIrOuuA1i
x9uHB/j9WLNXuslXy5+9rZWp5Z+pbo5xW98jWzua9gJSC84RpGuabgalU613kfqG
Gmd10ctt6u3GXw691iudISpOgG/FwkpAAFoEdGcAe1zM7BoAY3M1GLL3p9OvIwew
5MAlzn4ocsSGV61+jZniA5pmcYxT0iHL/FkRuxffzenK3JXiUQ2vKzF9K/2nQgyT
Iu5Fh3e4TqNGMCkMIgz8razwyeXdPIMG5rnGEIV7KKxLNhF/3cAzKedVLEyDdeF3
tv2sARtrEMBhk6s2dP9sdcGacLAOrtcAL5JEuiH9HFfgPGqrjh1CpDVF0gnoiH8l
ZAVZU+Ti7mNvnYoc3AG6e4Etb3XEJUvJ1jdESEi7lxhI9BNiOmPl+SkltsXnuKFm
6xmZGPi2pvwhgCoXSCMxGE1Xm5EpkuYBa/8Rmk+AfhhYskb0pwMHWvveIDhweHWk
eEEkWXTHLbAe7c/5jeXFRoJJe5ogM2lZuZfMVh1moMdsb7WJKK/5BpfGaSfe6R6M
qZUWRwf2E8Ne6oFWCD+lgfRS60BpeZguBfqTpkgt2aglQmL2d3b48ogHp98Oa+uv
F35Ofi4OkBSZCo9oT0HrV+bQDYKHlRr0frHxVIn3qsamBbya2zYan2FMajOmqOUD
dqLofvZZWK8DnmpkuJevrdCfLwZBZCRxTS9tZ+7hcui6eoZ2YmhM/6wLwyssffCY
io0Kj8o3jInYbCf0jokLBcZvsgfaAH1/1R5tGeXdTSFM2ODlt21I3tmIGSTNqnUA
UXS2+Z1lbmGWUQbzuwWsw8gBNV3xPah+/Y3siy1Pbw7bwhFLruU0YJMULYUsfvo3
aNTHPAEIRbOwqIMdATANebUeFty84bJhTFfCv6qarwLELjMES6eRjCNUOjD5iTE4
Q0CNjrVd5kKtJ+R/5znhrQHN2f1QP1mRRprGgy+wNdOQLNHwOBcaNeB1zwojnEnj
rCasfPmxSnQXVIDU5VdGJDpy39DIUE5B/BfB5fEdrcY403bLVR1kOhJ0OSYLzqbm
FPVNcS9NgSIh7QwLI/i/Mrn7y2W7FcYDGQPB7UC5HwMJYe0WM8mOzCIwP1BmZwcb
0U41K4woVsvkAYXaMAjyJYEYvWwRUMzONVge+eEZBnJo0hDN3X4tcEgKQnTjYCyF
IMDXb/kdD6E5f9lkl5IcG3WkLSvSvO8YJ9DHdSc2NaDQbw0S2M9O81kPzm6Ua/eO
2XIZZM1jeIUAmSaj7r/XMABACv10B/5iKBMabnArXmg9idI0XgRQIo4GSvwifVQ4
G70jc0+su5tuBpZAdQBXhaw3Z2lAolXK6wHMaIWI7mLlw6eJgGRZZQwG/i6hOBGr
LE9LkG7wrjT1WIJUJ8rwHX5nzY1W2nnlFL3I6aj+LjOJATLVACYMLEXYPkjCloho
WSqLVRF9ryj+gMyMAMPSstfPla5ILlPsohPbJxqqEOBcuqFoRbtSeDIAOhZ5FrVB
wA9kyyST869d/ZOOqZDtezNoZUPgpyVaucqdZ0vVZfoddk8CnyYwMUbNz0tFQ9kn
tE37TsftVSR17Y+bIIh+OFzAUkmp/mNcWI2CPlsMzVQj5iQfUvWsU/CLzpiR9Atu
4PULWTixTzT5iVy9n5fPSOYAlP0lMMCTYB/Z5OVAupTkCU74ZyD9+U7USZ1p70Te
J+6ZTXBX0mRqBufxw2IxlIT4eFUN7yK/DhqrDDSjl5cNsIx0FMaFKToOwfUK1fmp
dd0/zLdSva6K7h0263JUW9IcO1ync9fNz8kIElWDslRGsTuAqtTTAC3A8mylykM7
7faHyYXxkndSO/7TfKmSlpGwBcNG/6K0SVzvjh3WxKu4pBJXvZnnlA1RXhNN2Oes
HLM00LpXI46DEg2cGSzfmF0rnDYidqXntbKMPpgm2ngsvDwSW9UXdvqRUEzVO5FE
vJNk+8GAwy8CIu+LBkkpcf0XR5SV/BCW4zMnXG/jXwFfTFAmcrt2Q6Gk71LWEQSv
EV/NMfkjahaKthZj2E+w3Ey2SlfYb0eu/UpdFICsLT1oo2n1QUNGhjcChT2KMbRx
IHyXv9DOmm2NYd5ARrEL4OzsCJwly5Vewt7WmttReddOrw7Y4btyW++VMaBbKoeI
GyQ2lglSBN6umsQw9umUNfd4yUiUBzxN4YO+1zrPYJQZZ5kRqusbKRe69OTEc8dV
XARqs/GC7vwbCZyBzBxAVKxXf4onIp3EaM26qPNO3QXrFehMUDWqpozzQmvDIRte
4bHZSROF4r4Rq9vbBcGTKoIUbjWAaLWQEtbTkcBzRIj2FQXwTwGFJ8FpQK0sr4uH
8kpGQKTdM0PBS+Dm53gqSofeCJkbfK7x/n03BVUsOSxP6JhmzmAitbXQlU8YEKei
a9F4CNoNRE0VvugUrNuUmHK6tgYgxVWlxdqgsfPmYoKpfBxEs3u+cmQuLb9BBfgq
6sNdM6QdIFpEZkoUK6VrZUYk6aEK7aZtVMj3oyxQNBD6w6A1ur2UOJhiitRJtU0U
n+WcZVVMGKBwklix2Hvlh1/okMRIG+THm7JIPNSB9W8fJMBPUE19gsmjj1vE6MIP
o39CpAMxy/9+C56g6wEIpzpQuGabMoUEsj3QLIvvI9Ajd2gQ3r2DHC4Fk6AVgTgA
KP3yHaZIGsuexWc7+Pi7/ysIe41nzmq52McgpF5C7fq3unklgcpXpvEkyhQhtgl5
UmNxnoCgh+wWoXNmtxV1logJuKZKN7PhrNyRvCu6j4aLU46W5YKjqen+SfcBtTEK
ZDyN/rdq94Xjag7Yy8TkppK3EeAqNMYNuMZV33jJGhzugkGuhTEKqGF60UQR1Irx
odVIoKSpyy95YQFt9ejJGoskaokDSz1/4yhabNvy+17qcnf1NRi6xjg0bPP4A3qf
2yFUhbTbwOGMIbIegHvnrOEdtLlnFn5e3JpJ2R17nfB7kSV1Wh5bOhv7vEeHzv+I
S8iF1EstedA2s8PVVH5Il655ey6A0sJkeiOYmtNorN3U+XvKb1Y90dsu7y2OzacG
/lEMfEiWFASyNvqlmJRIs6u42QQIYdbx63JGfEu8EmBCUH9YJ5fmRcJbpGh/dHVf
rHc//nLNv+mLcOiCOs7NNm4n5Xnm8MZu3wlMXIGK6N+efCXKpeGiKbuHCZ40Wxz1
MB7Sl7z6jv8CVcbudr16IhnqJMKrd9Uwxb9jfeYtWLCvysbC13LuwRKaKZ9yRoGG
LiPKHZK/AGaTaI5EZ4M8wGrlJLE9N1Ju6V+x67xSZglh51v7XrknsPknyAd/Y8AH
Bmd0D31ePTpcNLgvR5O3MIAKrhDiZ1cCD0L8+9ybTJTe3YBAwM+DB9bEZdl+y2Kh
7Hux6psdEhoUkXJqgJiae5UsB70zHDHLNbZRvtxCjG4i0vXdf81IapdWVjn8cZSf
2NcCb182QxClqhm3cbN1xRCpaihxqdhFlPdKodgZmiJ8QIJmWx08DQeqqoLbb5sD
J8drqY09W3IB1xDDYhKJDirfeiyfIMxooxqXkeKEuvCywiUvmko+WRxcg4yJxP1m
ZgojVzHp8NDVRxdTfBoxfhPks+nlArR6l9FrRpqMRrX2gaR5CoLhl79Ktc3j54/M
HaPcGG0d0tOXqHNWAwU74q60bZ9JDvlOUTJs6e8PsjqKp+Au+F0IumeRA6+rAKe3
RIwydoWJUFK3/wdlFa00pjutmla9PPa3mvglL/jSDMfxR7dl3YywxHEgDGLAySNz
cHHolzPAicOQbX1reNdg1EMZ3gFIfWIT14T3tIaouKEgTOjAMnkbfKrEC1Zgz28S
goVcFdO+ihSr30/fJesrku2MmvTRn4L1W16ifjyUfTDPDoqREkbWT9P4ObeR0kng
HPu+LJhUBspZUC27QzupqFbkEyiX40PNqgJ3m1y6bHz6Xni8c7FUzX3N9bbc8OT0
5fLg5Vy2kR8HMZ8AnJgFgiihfiiexTNilOuhAL3bDhUx1x37ijNQ6mgHEH8zyvt1
8dGonlkCTOcYDQHPaRNc1gnPCCtigNIAUXvrqTl4/tp6GP/FU0GeMh1+J8veHTOu
QoUdsuhnfknFy1qVa8WUqWD/RJOABu4fWhp7z5SNGN9MsWCH9yYEeJWQ06TTtg5t
PXWAJmuVaEzsTniyeuYPW5tJnNjt8+qnfWD0w4xxcxrN72HDJgWXbgCpdrLMwX1Y
EKtCoYgpk4c3aNjP0zyxT7Sy+wUx3kwLJxlkuTjxNLE3muffMSdnC61Nrjbsz1w0
rcwiku9tVfzmcbrwZ74Ci7GW07wV9wT+V8b6vuBRw0KIDYqN8MfplxUJ8SqXH8UP
FOCNEmSGUaKpy4dnlynA7kk37Gs3GLdw6LsDN14rofqtMWl9ep49vIBxQn7pf3JA
T/gv+/QliqxwGwC7R4hiUO6dr+UYtvXbrU1qSiVCaX0QgHMM5FrHCCP9+Ehw8afs
xaZ5gTp7JhSGGZtD19v/2G2a5uZnANMbhrJvRdyEsQTPeOB4DMa6TAbgiZWu+hqL
nBAMxGV8CHjnEbuV9V7lHm/Yn2tbFhuDWvmQmUR6Thx/jQ5J90m8YcXQyU1jHBR/
oYzovXK7pkojNxIti1X/cqWbrfbE2N2maeBgWE/GIMTouyvjwbifjs+aTpLcIwFi
nFgS4RHdxS4iGJlTFFgd4dbiTKzAFOPLTi664uOZcL4MTTFN/sXqEhn3j4yveDEm
lE7ZKtuppCm3EzQBmlqS/tlbe5hpl9/ZMeCsBpyBon9Ww37/GWF80C7EXyOkeDb9
ZLBsalTSdQAtMDJukRuICFqG+07EU/nj8PcxjiNPhvJ192hdlNFGaeQjyP66f/Tp
DehcG9+QnLvJ3+lcTPbgof2m7m5pyBif6vhqKkdmYvB6xqzWVIDWf2p33y7O8lT+
Oi0IGPh0qQcD+bSbf7MyqKwWCj/wZUmL+aKC/bgrrCgBSRWxKbBQfvtux12Ffwkk
JWx+TCMOmFLDsWbocisuzj3XRbIIGsbGE6ESdhzzlROycSIYbBVtMOyJuhnzv/MI
66t9l1pkAm0biBGF2qFBi8j1T5PE0G/fthh7BFX5p/QkWidUCfTVo3i3uqXFAkb8
9uOcXv1Xv1QUhqokudyTWCUJSwqoB4LAmD7VkHbxdxTsC+py91CdEIYDmPA+E/Du
WKzX0zHsa+pM6QycEiEPuqkRoFW9WArHXxyyse63y8htB2MFxE8h0JSELTKeN8Rn
BP87EFgLuHIF0wc8eLfcE6z3fCaSzkE4kztRdSfV6HOACQCZMB/LxFAN9OdWKDed
3PCaqxXnbRX1eKpOBbQdCCQ8ANBLtQA4ZVqC0zx9Mw/gqzCiQkk8b0P529uzTOBL
VqfuH43lUvCswy0Est5zn656OvqtXct+3gm99zUCj1aLewaav9Jge3qiN8qpf0Et
6c9Y9zMBCdTiB6FlLvreGhkBxHNHAdlGmPSK/YmmUD5E6ThObiOxc1iEgAr2FMc8
IUAVzJEli5VeCjShoQQc2ps8veFMstOrsH+zdW4Si5TvLBeotOtVrMU9ddqE9xhd
cYQvfiMqWx3mMKuP9VXnab+I0UNXq3hOdYHfnCx5Cny6bw7f+LCZ6IHnHV/sz8HI
RQrcprr/qVYEUTlxEwCj0QApQbG2Jg98HabmJyIwWp/VVDG8ga4Cd0nFPQc1JK7O
qZY59X4w+wGR0O7xkIpLccQ74ykSjW3dTD0rWee3aFz3S4vyIT5BGUkDn9yYSPag
x0uCtDK1iqPptJC1rPHGOPMFwLTooWcDRpiF/BVi5z8AbK6frNAjvqKEOL8mZZzI
CY7Se7M3OSLQ/YqYUFX9VO2qsa03OFQZPL6jnJUM04frVIL7mTci0Oot9psX4jFD
c3DuZD3ZaEQoT3H3t2BzggjRX/htBjy72ukkLCinC0hkqbAi+H+bCyoXFHvF7B8i
Q0wrFJJU/oxu0fC2tbvwqh4QKqRbshaZvpQIiJ04DzEYKrrTrExWqpAC6iEX7+jN
4k9Q0z8h3dvDR3K7+ibjTb1e/N+o6XAO5TNbnvwzUH03Nv1z7GDo2bZWHuHRyXzR
S6qvUKGjUX1+A61kCmf8kerWHXhC/kJEXutkvl7ZvWn9mN497lK/zAjdyFLzu0ua
9UUHNEZ3iA9cjD1NFh447aRVpdZoRiLkpDDOkg2P6/eiOt9lKiMgEJFmctam5U2f
9LW3xboj0aA38uQYKL7L30X8iFN6qiYLRGnXLMQOZnvsCwBfAJcD2chh4uFa3bQM
SR54yzIpXGZdZ+xaVw+iek3V6mDmY9JaSGDo/7LfjwOPFlQ5qFR7I3e8dqAjI1oa
Af7ITBaRbkZE98g2DhJNo299nfw4xtUGmrR3rjptc0YhoaOXOYcO/DUGq3oxHqfg
nvEOc/ZTMbzVZUR/Y2jAKv/0pJOU3mKpTOdlP8FLWNxkJaxw71HnAIAHkhRK7uhC
VxZLVahn3faEQGJsCqxI7eWPrirDPlUXyKVmTfqZlGLBCOIZbN30XljRaEq6ev+P
pHmTSzhnLDGcNqkHUj3DIHIw8V5W9WV2TQqwMRd7co0wcqkLh8RMjzHIOCebMOO9
Y8/YVi4gAfOSmY0aDkV+n3G4uHHSicaEw3B0mK1fEYIv49YxGDUb3jUI6dOvbj5X
zE+ngKV7rZuik/fgQQXj/vEbC2AL7T1RKJA71+OIMAWXEyJZTCPHZmZAdF4QfSQ0
e7Ff5H0k2BXusqlT9dEk4ur5B4K/WDpHv9D9q8d6R4yTpwv3y4XfhCTjWQZgcoFC
eyBtppcoxlfrTmwyxkmfGqvvvRLbNqBE0sURYHSgdJInKov2rnyTWXXT7dI8A0nV
KkaL1bdGy9p2mIEoO4jmnxjZ6kQ/6qTzuZvcVQfqbnxnQ82GOpCJRZgGXmoNtCUO
JxernKoR6NZ9PuQa1Vqds+linRdCtZ/cXb8i9TIf9dLyhKd7a4ErgcrLoD21r+gZ
zsHut3pz1WGJkHEfoK+O2oj9Dz72VLCRbME5NCZcnDvdmO/u/TWW6SgmdqVNHeWo
zhmtPSsIHlP2sOXVB4bjd5vWE+1I4ke9BJkEXYQvoaFmg+8uzlIzkyXHEygzS7e/
wxRkhEtmhGr/YPD9UjWs0OOrg3H9biQHjytryVqUTLULx4tPHogYUEC5WHVp3Ikh
eH5CffVxFkpc5o9EaL80frqnJhGMQK+U5TGtpKJtm7ABmP4dbKX8FBURhIEVahXM
wu00Zted+ykxFA3o0wVJStBA+qFQleCQ0uS7Ajtclkoym7Jf2S/nn5d2PXLyWaCk
8FA2qpjWSQ9iSQoiqxqNrc1i1wJ4rA78549Mvc+7G2P5UdVYPrlL+p/Ksx581hvz
ianGlhpHcmgN/x0Nz1fnAJW2158xmAje34b92x9QNep8kr0tn4FtXymHGewEUSq+
B57LyEmnvPKkmFIC+NH9WQ7ZAqEyV04UKLZ7f5F2PXiEVyKdQrE/vp1vQp6B6GAl
1GGsLorEPYOBHyOeq31S30umr5dhwMCc1rAx9vG+SkIsc0ZNAXenkuaHodFWZ95E
e8nU3RRHCTRnz1XiWOaCyc8VbLKZ2l/XIQpm7pULHKXOM/VyBDLzyg/uUHAJVbyT
qDWTa4/p4Ydzf/nWhye8eobCw1HB+N78TTGj+tmQxCNNbkJFaDjZxiKRclE59Cpa
CXpqvHIjLKu19knEmorneNz1auuOISl1JiekrYkez/54Kslj4XXFYC+sarDgNzNI
TMGiaT5DbIAgEKDG17ioEuBnNdJHXIdEP6pjT0TNHLrldkT0L0nAqDqM3/gA5561
1MKYa0JS1yzd03ABiXYCdRlczCIMOi9ql2KS4ONRhgqlg0yf+pKhb10LoTpDMnl7
LXF3bZLILwg1+Mkx2kvRHlTNoTRabIgCIA5wDXW9poxwuCbYsiI4Q9S6oyihMNRF
KPKnk/k4WdeEnTds2BEn7O7ldapxWdbK34Be6bSihdaaEdhQJjdeV+4sVZ7Hleeh
zR9/neI+w6h5C3Fgku06NUhnkBbG6WEW90ftT13ijX63I10wYl1tA2DOYL+gprpV
8ZRMKGd4WMOk2JcnAr7zfOFEYJN/gYtixEVgJbHrXIc8JtFkUAGKfspLEtQNJZJ4
dN0Vl4zeAM+/sneA06WwE+W7z0puCbotUS8aAd7z3e5IyDpTzvCLqPTuPhuQ6lML
LPAxImL1+tOBNqc3eRO4NHHBWuk+FD1b+m2+L9Cz1Kzs+O3tDtlHeE9z6isUeMA5
uEsJpbU7ZDj3PzboBuXg7ebcBJUU0LPamRhyszZU6jTQdJV0lu967sRuqDXJor0f
NMcaqpiHEr2VFj7Y+T6ognDpKk9Gju9Cy8ss1MfFSMDhkVVkXwDJ35+Rv40Zn6OO
PNazwIfR13FkdJPPXgHGGkZQAQNwAeHmPnc9/kpygX4qCWrtqs3DYxK7smsbCRmB
wkA7dFdvFiHgGIQJvhaQkg8yNdizfPmRX4+oX4YoAibYZZcPnezdfa1P8JCzKuNN
InF+4QY6Dc7jWofguKk8pCWFVCLs9ElYw8INhpUUB8I6FTCSKyucZj0yYBd5bvAM
pUzYguZReq2VsvjJOzqr+Krlyh8/ezSc67hQl9D0/QGsZAvM3ftwGp4+6ILFoBhl
AraeRrsbCuP0Kw/DWOM3WPzrdsk29SzKXe7T9NaD0oodjHqoK4c5WKye9yuNJv+r
92X81I0xXTpOxPyeMnv3c0bhGoqNEeL7IIPG8NI/ZuYmF2BvBBKxenJZ2JeKaCyv
MHxZpvvb9PzCcfCg+nPilOidWIdqjN3QH3Yf3C+so24gj83uEYOwOLfngH9M2thJ
PtHYov2sCL9sRV5Xmn1P7+wx+14DprkanAa6FmPpjIMx9FBZSDD/PzWoK9ouunvF
eHLW+AO+JdnCf0a996zO9jwHcQok43ZvUShprg79OQXKl1FsLkE5lAnfukDD3rgR
IgiENnY2b0g7kFF7YmHYcrgYc7UgaddVt9vUaFqvyLBLombmuapyIR0J7xen1cOa
k0X/4ptAzemvprRCDJBP07x55C/xHN81RIJIS1JlncPYzMaXjSd9boS8OhdgRwnC
YytDrF6uERJepvVdqVZ6pO+UxC3SO4XGKi1/cLO10tkzxa5eyx+whB2Qw/cYWl8M
zDMSud/OaBDcZ2emAp6s4b55W6P+NeU/RQcIYhUJt+B0peBPA1p2EPLN4X7LeTkq
opn1bN0L4GH8lw2YjNJTswHE9pJwbtaLzhjkhBBh7+mV1kK11p61Ur52eGTV/3tb
AAv9OyXykc9p18SOLgKUb4sqXHSMw52kGYxdbCD7ouf1LBJs9ojdaHM9M1a+bKdt
ipsRpO4A6K71IQ2IeM4vSf08EDor+GzS5b2etRz51J6VwS5b6VQM1DFWPNFBL5Yw
BZMmlirpibaRv8m0kIfdplhgYtJuGbtUXaJMiB55VWMBDQoXO7qOlUmJDnHRj4L4
OoxIW0XWIa++r/S5F31E4mWh5y8AFAC9z5uDTZXIsZ+EnbiitKnr9GtxNrW8YVE7
pc86F4mwRzQPW1kKFPWCOOXdzCcjGl3UrkRYkTVRlndD804ThArzZIrtahpCHm1U
YQ8KiM95k96aj1yX07SAA1RKZ3HwjTLikp6TmO4mPf9VssSkoB3QuuguqQE5FQJz
NgU9KrTVRpODyI58OF8e1J5JvF5q57kLHjhFIQaEMc7eyKJaw7rzDm1lsWsli2Dq
Vb/bCjvZ5G4fSH802uA/Y9aQot8/iBvB4RnbDxzoBfZKGXoPx7+hEHGJFA7G8kUz
A1lGVkbjs2jXklTVquqlvF9QF3hXyzPeiRSPXWA7MGxDami1BwLjWnT3UEed20hb
dCIeVLXwJEWcTou9XqLBkwmcBW93Y4id7QDx0xrMoPJOgrSJV/Q/3A6LlNz02G9G
hCrFry3FJz9K/RXeLLJGXqvFJkKlHdDvxABM7fRHdAO+k8RNllhrAGY1AZnGkGvY
oF0r7URCVwvOyAGPC2y+JO9V4/R2cJJOFMHN8Ujl4Sbqhyor2LjfAMJoIkdT1Emw
2H9nkseWRKxESGZfC0TxqdNLdcIQ0CbTPjbiXodey6x9X92xnX+WfFUPH8KpgVZr
E7t6Ywj6iTqEfLeu2L8dpcgpuLysmeCDuAiMd/WI81CI4wMdBmO4aPgfY0F7Ni2W
b4MKgn6QOL3dEDZWD3FIQgEZWoeEwe4P2k8Mv25W0Hzi6kovEG2orPbyf6t8lUrJ
1HWHsXN1kKJJRPtljyvTukXvrl2py6ANsVLN8/3s2X34VKr+pxRTX7m7AdVlkG4l
gncxkDTa0lImVwvrErKixToLXAIGx5KwM9jFAGJsAl9TgLftR45vus6ddD95CBrD
1uxUdJ+CIGt9BmwYv7wc0HFaBO9d8+3TMAfqy9HDh97dUZ64H8QkSf+OKajL7ulC
bbkjNX6f6ncr26hQvxxSQ6wvhe+6a1TqeASD6zeKxKsT2VJ5elOpNfI08bMWqe+B
nzI5nLlPup4nYHvfjdArQTbJ1Gea3znlnH26q3Mw0qSTpCvbfS3sdSo1MFOBP9JM
M8ujmOGc9nYSu54da2B0QrGOwkG7NZ/2NCNDqGFbMCAsVl8Gvtnpop68QnaCygv8
TszIs0UWWZUDnky6idk5kAQrYK9CRXS37CapiTkAEyVZ42nK9iWAb3rGM/A6O2aa
54C6K0CedslIw+O08FDb3P00JjL/RyN4VBHhLoeJBmh+6Fi+M7Yj4nQqZx1o+Fzn
qJbve0z0owZi7vkyqAkJR9KqECeb0L/OFLsN92sEp+tvbc9Z0E8fmMNLjb2/Fx/f
aLeqvXqfPEA3amt97FxY9ZZtb/65NFsBa6dQ7mptyG42k0gX4wAhTMcSGhWRrb9r
53rMp6BkJK9mKFnr4zoaboMIj12bmVHIVcKwl/Vp5lDKRq/+GYIcj/2QSUlv231P
iqbGEkEFJxSFrFZn78CQwcp3QqaTOHP23BxDoWLG4twPdZI9DbfE3mGytwIst8Tz
D07ovX+OKGMTVQLwAssWxlebDMi3RrXF6nxPgGVj3ewwhC0gumUCS/OSIls2aPck
XxvLLmtwm30cDBvJfY8niUmDHJlm3Q7OjFyu5IzWeZUmq/0jR0h7Db2lrYCSx9FT
pVi2zU9k92pMPnPBu6/Iw3hKR/Yvl9MRusJEUm+m1bO+5SExsa+PnfQD+LwkSdsA
9YOMupMwnTNdJH1eWGz2OwaoyUEIE5VEghrPveU01I60n6k4a6kRf73Gs71pKOL3
TOXnFB9evgZaF/nywi+YY0Ppu/EvvVNffpPnsfkaVlzJ6MDR0FpPGXnBoRj3cruy
8qpF5K6Ybnn/rAY/yc5Scd8uT3nur8pLtyN3Zc7PzyFFq7RHf3vwFd/xn/ARkMOO
VPV302ZrUH2PzTD0yiH+VNtHXNJN/u4OyWh/nQmeXabA6D36GqBj+KuHX99x9Pcc
dZKzL2PH44uFdebixSgjJYxtw79bwcE+HZA6LKWH1QWhoMSQwdor2amaowxuWMc1
FhhtSgxpH9tHC07D3++DWR5gAgq6t5jQ3E2cznqDHtfAWn9rYmwBuFVwk8mhZzlx
GsqoqUNMD+mJ8Pkfqjzx+baob1s0jrFp7HhIfOE/AK0KCuubVQs33aCkQ3qPgd7K
qvcvE5p2OjkhCPbC12Nl8EcfPBIbPc4O2xmSHzTCJr6uBx5/sOZfQ5zvUJLoPiJx
qx5B3XW0mJwV0MGCQsI1Flo0g6v7JotKo0Ao97/t2xbDyuh8D8ftiCbgp98GU7ji
85/YVeLhxAB5ja6I8QlV8xeBX2QuzdsAiJ0o4xtGxwI9mm3YXb04bLAjn491udpR
S4R2o1xylp8UDsA6gIm4qkNrRTFB+VyqmUMiGhkqSH4G6yy1KHFrc0vMnYqXV0sc
AVpRAm0hpW2EdZD+EDf5VKsVZV8V3WiuBTwLPFsf9gXuDKRQVD/JAdOuE4w5i7xd
P+WBLoj9L55QgBec+7kTia7jjglFICy6IyXvBm6mgxuapj/jwXdexu7MTppa94Y+
wlt+oibn0R73J357am76LJvKP1aiC2UZpa0evAzVOowZMKx1bREL/yjzPmxISO+7
W9VPMA/JHWFaApOFrO+r+x7iQM7JZw8KIHbCRNY7PpT1Wq0kj52x5bu5QMH2oyX9
5/g6SJ9wGkqeADoDc1a7HPGf1d7jJBWZyYqgiA7SKaGN+K2IhCP9e+8HdBFjZLDM
TCWTQ/oKjZBSyjA1xda0gACagGWvtGKWlDZ7MFHw7sB5vu6CuUfxP6ewhQSDp9Dd
6syxczFF3jGASc1qBhffdv8KoSVd+4C8lLBfL4/TCPlyzgEcj9d8AoH3u+SoKMZs
YlGZETjm3QewpjOjF1hsb9+WoPRZsVY9QM8naRCU1QbE13O09M6t7SMc87tG2JQh
y7QgI7JfEeEKwJJr4HLkbqT6poLJam0yidUQK3FRALM5SMUrtvXtBC9fgIOeWhYg
G88zrZNMTceEVLLBWbKlypts33XijZYIoTOjluv5j7mZNiQIEhVkunhAgk630yro
z/wHzd0Nk5vF1BC0wBYC5+XgFzOhNTEPy/C5xgcplrWzlJlVWqQ8GhRbahwQbY3L
g5ESApZsEm7PQOkXeCpBt3IbTvguINM7RXcsgaQsyWsQPW+2iU4RU/LFBwpFbjiP
w23UZ0LWPxwddtQQXqTOgkzJdr1mZ3WFRlq+KlkVnL0vgbJ5r5PwQb+qKoTT/4dX
DSotipSS16AMdajg2hIirHcWOK9hHcpL53/u8Kc4qhdehr6CtrxAZXLCtkUUO4nt
xOgYxg8dr1qfOyR3ffaGl2/4hUKADscn5n+QPPRBhoi+tLEonGM1wbK6ipSYPQPI
JVY0GUIz+Ca2axerndT7DpSYuhcYOrpC+DfHQw+dBXFCBAlzQwCVFKgQWG8bauRa
irrMGdLCXvVkwrz3WLYjs6rAjcxMgyzaZ9tUkMvL7XNJ6i73jOrNhm3fL8SiNGHr
xGrtmMWYEd/9I29VmShaziGONMqFtvRbwEj5eS6U+17wQgc5W8uHrQwH2KP9u7fr
6F2Oqemrwq/GCSmAChpgggRMnzmzSIn1++ExGUf1Q/9IVwgU/YreYZjh70zsUzYq
5C3fYnzUvrT7Wu6mySpsHaTX6Nxv7BPtkHo5DOrN7JzTWzCB3uthvfdb2lnbsDJo
fBSbbSq+HpCly873IV2PHd7YY2RCHATkHTtQevi71NRN/qaPCv6fXKNfT0xofOQU
YAWVRHIo5+4P7/Jj2JkpUwHwLVdYHe1z+djTUXTrxEDofROwtT/3nRLVG53qBhIh
SUWtTTxMocVglNU89Cu8iRthwTkOqfx/Dtdnb1VaLXbNdOea7KG5L7Xo3qROWTpe
mFE55oUlYCV355QwYRgfN2l+5jaAloGbqfnWkT/GsvB27y9SRd5esCOPG4txqfC/
cWtXUcaJwd4WK90HsAKv+wY8YGSCkl/cf4m+Eng1TLLBv8NszbgiMq0+UtDtLbVq
sf+0jOP3M+NVwT3iw8A1YDxW2jjxKtVdZPA04jik90V1MQ8tTGZbSiRNAnqymvx2
+C0vISi4x0uJwmnEiqD8Cw058V/0e5p/mvTe8UKsowFT21CGsR7Jmzx/fXfBWciB
monOfD4NfWWLjMHGGhH1m8vJfpOG0bjwdNN5RvBaXalcQI7IXFNR6Np9qZnQyyty
d5DVR5eQm8NaV5wo9T26vHEgIdlwnVGRfxhrcDcpfxMw1Tw5G0JsLQ1mw5aRMYgs
CXjvN3arjOajAUtdv8qTtZOySwCi+lQLqsZDmzCktI0Ib7uRL8FSs0rRDcb6eBE6
xYchAyFwInFq4B+zGnVubP67G6V0cK/EiOOcz5g0WsnJMLKy0v5HDgKdqifIP3kD
jEX5MninupuqjtAOBgVdKS6O6gQ+ayrrSzUvCK+Ss1+WZOs/4spd665piE6uYq/5
0SZ/RYwnkYERvb0sxyj+KKo72/ToxvXzazxV780/G1v32dIUnzZm3SSUrEMFO1Jn
UCTkj3SVa6tLtsNYOZnbJ4GqER1tA0ttR3jTk9KjcEaF6FCL4UFh/jEmVqD0uYjK
AIPENWHih33pn6C+RlhuJYew4QJtxDGerwuAX/hGeLKqj7BpqN/gMi6dT6xulqAG
HT/XFe2w/t7AQ4fUdQoQVcyLM3B7PN6aXTUQRBBxTrWaXZJ+JtixdrrF0zw80q5D
vQnyTMmUo8Hgv9ZTFAhGRioJXTxrTlXh64JUgJyPYytHM8D4TWGTiSthymbOXMIV
99+p+17367QiCoO6dLfIhvqk/rlOrPv46FJnWMd/j3wuGn2QX13d0qN2Cm7CD4dv
wI7x6k1kDuBlsPWmpDvNMLf6Iin/g5nb4SCiE8BCVgiNCIPSIraCQ+PfE7rh6EmE
Z9H0jVmgMDsxGrgsd+XyYmvE3uwH6lS5lfJWFGKySd6AxTspRVZqD5WPUee+xkZs
viWa2Py93ey006n2goLmwJV8xuKd3dLa4Uk/VndT4d8LjKqBLrpWBahX9ZPnn8M4
QllqJX4lZZZoZl25aCr4/5rMld6dpRE5QeB/Qj3m8AKTvESTr27tNMvnH9LTUv7k
fXoZH3IPiNpx8GpwTQrnca9jGqYIVJAycExN5wKZA3bErlujod/rSAghrFPQFlq+
1y8LzIcb3zzCXnAtKkC9SAtPKxsSffzRkW3jX+hyijLEXuCeg9OpFn/99DQ/jgDt
p+n6v9wHKqbnh4zUBzWFidbtci1xB4d4l3uKHqlH4qYxPkbtB0jM8NehtkXvg/SM
jOOESC/gxVbnhgLE03LiT+iOuDGz7njo19Eaunv8n5O06YijA29lqO+7ZIc5H63j
QMbXj8pca8S42H7sKhsLpaY7KW5vx16EI57GPwdlYg+FrbFC3Q9eB41cnp/ey423
sCc+O7I7rbDqHKOSbNBrvSwko39cmFwYWSOy/8NbW6qudacv+0TEH/ed+DSbn85Y
vqT4Mv6mXgsEpEn8InnRgSWxyohwo7JBOwHWuxLI8WXbbTiXoo8izrWfFo8Uji5I
mAeaXNGIMYq/OCCvADZmYAw+cdPxJQcPhlZTR5M1EChJDBlRa19RJp/dvr/kHDft
itfQOsg//6SXub56OW6HqsXR9ToMpPQa0ungjzA0mtq/n0wTYTdUxuD5B4kc7AyR
T8akpPH7t3V0CdBhXZB/8rbJzb5u8vYwaumeoudg8zCMyk2qMB/gAqFs78Wb+D29
ZVUKAf0oe+4eINujOgozKqj6C9beiRK4AhhkNY92T2LSB0awh4XAZDDwFmQ9aDO3
UteDGAEVusEairDXbQDZXIFX7WMKxGvtHhpO8h20eMV9P/QxGtbmgI+SFtCftlnY
j5uZxQJb3+WgFu9Ld6dnGg5k0rpNc2juDDoZiaK8lmaffZho5z8QappmSQhRTlDg
ZLsk0hAGlg6KUEzZoIcqsJkko6TmyNayXWolqYgsLhspLdESONlMDimR9AGQwap6
DAxyiJFJtT/RqkFdaoZilHzybqqmmEAdXXgro7IiMvfNj8mUwoEyQbDIPGKHQKQF
rJA8QWNCYjXVer/mFqEMPafipNFB/9VtvQWEvKdPRMqza3NnAXuWiNx/IJkgnKpc
DP+eLjjQ2lMmitE7cZTg1nrmqW1AiXL5n0VML8ZXmR9LV3LK1Gnm7P/3lRxTgEUD
SBcqdXTfuaLS3+D5Eo2nNIJx5GcXkRrMYyIjUWyX674FGMWyoyBKgQxDNIV91vLT
OCr+fHXat1BbDBH80EhAQ6YqswgjGrIuFOQBN+UVA+E0CQAjj4FW74vBEr4Mw3Mv
47e/dmOE9Jq1kMIDbZZnKbDbmUjT3J2ecPXZtO7IgL+HmOnH0rqLYKQSt5HV2Way
xJeIobMrHyaL7vWGoZ7BENN4syJh2bIRbM7kiUvLmxyK9wgfadGwYGkKdsLHcj39
Gj+5aPHj5dwUXZ5PlrI5e5DpU4tC3YqcauuWwzK3EnbZQkGEboQjB/dn5tHU6/8y
cu9A36p0wYelCLCc9zTQV+buTFA8JVa7nYJkbHPTFtLic/BuUz0yTg0kNwrtlMhO
oAjjomObecuk+rkT7dzSTAAeuJO1nTHNSkKb9MTprmbo1fdugPz4/m6OQwqNT2Qs
WPY1PjdLxCJTfvxLiPsqf4Uy+wd0JFAbDuDhQ3s06N/ixU12/uvYqvkNGVTquKZ/
6tyCEtbMPNKkOnXR/cjxQWEssTfYW2b+iwE+6UsSd41XBTm/fz+t8z6x/tz9lBrU
RYg/oj1krYhumHQt7nyZwq4tpZHMfb0eEm1vodlnpT4r9sgqXAy6IC2Vv+jSWukl
aGm19NzIvVABEuLxXMYLRa6bBPQa+G2wPoz0+1/7XK4dYZ2Nx6VzYfsLlGVMNZUS
innS3enuSZDZXWnzj90bjG0DSF8+3LgJMWaaz3077zc4zFTJOHE/YrB0CtW0f/z8
dUMs8XXs0VFp4+hncfjG+jo+wqvVL8cG4rXgVVrESnSNkRBZqLyCOVASHdypdlTW
i5heyupKWB3QJQS73ytDdOLXCV0NI51a395aTageMywESy6vhrRBWLOwsAB66KUQ
Nbtsa5H5FnsAeuIttaZ5FR5fr/16qo6ogaDHVNao49dQqsIYZe3J387qMhQObldZ
1lmwT/qlk7AUwogDxG0bpJl/4kmrelcUd8nVKOCnia8Vm4FFXaulBYd/D8SoxcgH
aWhGRqss04aPDKLuS6zEbU2Ms7e6ttgm775/HW4JS1SKURCkB4n79S69rhuIZsnr
vKvmciLi9u98f0Dzj7lXfmaD+49jSmk8CJ15zu4jPU4hTESSJVl/alM6pg8jOUKr
ZQNDUhj4aHyBfS3TuiYk3fyj/yUmSgWYrQQeDMib1pBwuhHKk2J3xZmE2YtUfUwU
tWLmSt4WiHoMEFcIQY04gZ+T7Hx3m+r5evqyypaD/K63MZF8wKeOh2nDv3d+ai03
J9ntjPeSWzvBLCCF2MivVKa7sWUOl2k8OhZDCkp2Kqvf5W/gOuACYYJ1H7b4VxXW
LmfUG80HbN/SLbL7mpjRyZa82rJ8cPanbmLyh2/oyuKYhPXbZHLZT7TuCkcH/w9x
/wUOjRygkyWEL4n0EVT0r4fRCf0/iNylAYa7n5MO/KYtv1jVpi0y/ESCvS1oEd+M
mDmz3XYh1yLK0B1n32nBDscfu78/wZqLX5y6NLbC/UtQJ3fGni6oEIXNtsdmJ/0w
jzWjzkFGXQ7+g21Et/9X9RlD/rzyzOGEqfOzgl5uhqRnP8PeP06i98vXhHs10KHK
AW4Gz24B/WZijFK916JSTLR/xmcfCfAbqAsHcU4lKVVZ1+tYMn0J/rvMoGrAVkxk
MRqUmq4tHV8SAlCdXRG/ok7zaRgFDjr6XKRDw4PloglyY+c7lu9qsJt6KbtCTHDN
HggMeP/K78SnbBrtoR0RxYEIEz+WjF+8RVD8qtblq/P1J3bSZ2lqueVOXsPkM/sn
EzvK4jSjDiV6IV8i8/yG1s8GbaLnwJaZLvPp+iqXdXAROeyFew4wLqCm++jUTmpf
xng6nP1xQKjqOTNFoU8Drv+pEZ+jqHZgpMy86VXwZsWPToqXTZwOPcN6rx2ppGCy
IqGSweH6xAdASgMZ1Xy5WDVe6rgNB+UqMel5ilS07TrbHXy/ezBgqeud+M91nTjz
AMl83DoSrW0Qy8wk60mNBHPsBqvH1qX2/RUYaTL4km3hnniFkZaHE3n+YgZ7Xg48
0okSlm+XUPLtSUlKzcdaSicXMv9EJQS3GyN1yUw5MEIRoUAHQCqmcFQHAFQ66wgO
kDitcfppCV+wVsRBzeoRk5evaY7neLIbAbS6hbpNBTzNqimSLiFGv+2gCCvAG7pG
G6s4k2spU6wybierkDv0lM8Jx4CQ3X5dsdaRYzN6pUhN2zeZn921qusvACQOdYfX
vukUyjZHw8sa2aQEZjrZw65mmaLXDMpWfEBPyr3c3Y4kGtEKNWr0n+EcQKobDmv9
zbcMvNFygyQ2m6LJaX/bBDkuABUMImHXTiC+hi6kizd2fJVIj0sCpTV31b/c4kcd
0+S0FxeoSefu6qdr/zbhbwSHhD9JoMFyZZDu/QTYVqa/S2fjhAYAelOv0+EoiX8o
MtOZlCK/N0eCKRUUFCRZJOHXrdTh+da9D8yrQ91+YPEguJgmvgl1fVK2UvuXsKMJ
9I3CkNrTbkyed9n7EdNUy06pq+ANRdB33oGLOjBXJ0PPHn/kzx3CqqfW3/E9se6R
nI1Guw5trnv//r2fsJyZbdYALpl+wTzyk3PD/WVhtJfjBuA1Xa0knbL2PWPEmv+2
MJ04GXWToXQzwyH1dhJvr75Vn4oiDt1U1FCVVg9NwA9rC/6NQtI6ToZemXVjZGNF
rZwGOTI7RPcmg4TowHWoJJI4576rMuP3FkkYk7jAhTzlf46L8Iuky/XSYU4nBskn
6Tboa3gwIo1gWERQ+8YiRz1IIEYwucnQkGqJFKPQDXYkLJJMi63daP0jMzhCC9ct
+zJYn/KwkgLAp+fJbJ+PinXdNEbOx5nonhgKJ31Fprnk7JOjRO+eD05eCaSvrZVH
m5zXUc1hpA1FUHGzmX726xrLA6PpZZCXKSj8l7fE+yRuV8JYzrbi1Y1BKibEm2IQ
2najL8ufVQtna9FW7zRcAStMIhfplLHBJwvU6OAHGNI/4G4R7+t49P5cWeHINaKx
OIQd7DKYsZlSqBTr4Iyj8UEH4uwDjUcadSyLTcpP7Z1azd+mmSZr1DbQqjz7rPn6
oJzx6R5Sop23PyZNdGyfaZQ7vTgkA1LB9L8MF0KXKvaDzqDsYRI2C2GaGNGvDPbc
J1X+QWPvwbL1xNY+K/QY34MtlonrQjh0dTp1lcRUm41twVMimiHMViroRbDlV7Ji
FbvRvuYTG94jnwEqwrC1ooe57tqgnOsJIGihzAX/oGcmv+zZYSF55iqen0Ya1quk
Pp4KyviZEwOVVvhgwYoO0i9yM3M9h/lzSGFFr/RmeHBXwJ5hCXbxbIxDeuTSB3nJ
2dvq60x4uWf1CemTkhrvIixZncWR3ksQVANZz2Z1r+jer1/Hbx6/2xdjLlwUCdPW
cqcTijQEK31bjnDOIDMj3l5YEfBH8SlYNbVKvgYIiwTEEKB/4I0QrEafMtaCmUyX
EROd1hp3WfDkDRnNTHdEJnQFZmj9O/b4BK7vT0evrpMrc+TI8fVNM6ZvohyXgF5L
Ws62U+TKLhYRICDL6iPIwh3/L32PaIkzRhKtJohXNe72kX5+jiQyqFVGTkaiPMl0
Eksi+v4yHsJ+vhQWrE4KnixDHx1klskU6FY+W+FgKBe+vrsPud5K5nwljsCtAW9Y
6EqegOyNMpRW6GwM8ci2ZViiq7HkfW8ABUh7OyF1XZ9F0CRND3QaVfCbCAXzd6QZ
/vmkiogmPn2MLY2g93VHOlxXHjudJT8sW1Vtb9f9f2MTLdlKL58DfTyIAd67SoZy
aahFHAQEaCypNXIoosHkh1GdlvGfilkkucIp7L1JPyc2ZVS09GVGZz3lU6COOXV2
4GCRgZ5sigvHF6KZaOxremxeEsfdD9dl0OP18DzaH1ms0KlM/DH0Qp0XLX6ixbg5
zCHlkO9cz0KaSuegIgT7XkRM084yrmox/NZjtk7IbrxLGf+DOUN4yk8qGo9eaXu7
h2AsI4DVbc0rE9S+zoL4/vmpY8SebZfrDffO8GE68dLGATfHB8hBL2j/aEBslkrR
2Z5m14AH6FnxR2E38U7Hmx0aZxxHDg6QWgMgIeP1/BwpzSZTENrPRofk92lTPK0u
th3Qfn5pGz6eJlyuiemVmbPGbXbMwB6cA1G1P+A6WQazcg4O2i30HIQO8Oq5VryO
08J7Ok32Jw7TldQgG8VA6xg2wcMfTDZ5yTxUg2W6n3D9D46gZdT7mUqR7MUQsuvd
2tfspOhruTuYT1AnNE387UK3ZIRkSNaVhd5qwXCTqgQ7k/06iRqN58NMTeVrI1Ph
2gK6MGa82lr6glciFMYsoBm3MaPwCAFXFepLb55VOsGFF4A8B1lRpobw9QIAP+aU
J/gy+MfVuwkWd1J3mZceGhCDVUsEdXGuNeF1O2SokrfSJgiPJ3kgq5EQnBnEacPj
hS6c6jJ0/Z1MGbvDPXL/Fjsamc6bAF3aszQQaHmoZ0eNaEamVydQ3Luv3vPCKj7u
kemEwxfNCIvBxCmrYH+096ljG3dKFQEyPB3iotsqCfwh2JTkADphFbQON/XuIoVk
ft4BRrBk84xelpKRyGYuCwnUp3yNl4c8aLmlqbZJir/tJGkV25NV1r6b0cuIrdu6
LqYryW4ipxWIgqwLec89sI30t4Nd012zI9F5giuNN60ZEFH7wyy7WZw0/f8cOiGW
Fv+T4Y/Cy43CvUqS1MgiCU2mmK7qZzOWZjtqinK2kgTL7i1lYknwexRHKBDCkAuo
gS/WeaR8VRiV36QOI+nfh+h2RKk4Ovxt2X8FV6DPaJiCx4MaDMh6qYfuiO1wcQMS
lMvcyajPcqO1C57GmdRMQ0+ATZDFaP2+vIJHZl7W440kAg353kFWg6DqfBxFJyGH
LfLaFQkz4g+2PXi2yWokMpmvasSbsJt6jInZMHmYuM6dO2rcJJtBJwclYIxNj1U6
HqnSTp3PIWvKtG8dFGSJ+ExPdXe7Zuk8kAHEw1a9Qc0QXc2qVML96vntKROsJbUE
u1gluhGEB8vZ/ov/WZAr9xP3SlJbpF/R2+9EbkkvPMePMR4Lg0ZyU+v5F81JE9ef
cpzcuFi1S9kpgoqxKB5SC2E0SAcm/n+pQbcxEzEJ0E/9BzS5KY8F27Qli4v6+K89
4y7fdd9n/JL3zqEEbWTVjfKqkMTNHE0irHsqLWiX8uKGyYG7iwcD6X0SBxiQ11tM
5P2yFYr6TnRr0a8Qzz/q4H3DZL1jzP+R5ClTcVuahdH3kvTLNYSM6+PY4mFPFC4W
uEjnpZpjk8OpI+UVUtzbhPS9IgSlnLFeJ5sojX4JDLsD63fG+sfZiz0lJF+T9Jcq
3GI7aVy/9xePY34WEmb6rzdvddQiCvRV7f1YrUwObT5LLUr6+yfpdddFN3RHrMG+
CiY6HUs5Uz9zNNe5CnBmAY0s8YTO0PglgioZcnr9QZo5HKDU+cyH2WpH8Ahjc40P
00YA5F2P396AG9RooYpvGO17aOWuV6mCb/ujQeemAb0HhlupTX2AJPftEO5snKeO
lvh8A93T0XUur9X9eAWf61jS8BVRdkoiewmdHvxfAZzX/0trwGq/X0js8thpUVbE
2bPtwiFTy68Lj/bslDdk1Z3ceEz5yJzi+co6Xe9orUXGZqq9268fvUaJZYGKxWMk
PL4YWPozQ6ETTYTQXNtkkxut5Bs/Uqg11sodKKMlr37ITwI9VqwICootewL0eTUU
iFagGc4H6H4vme0Wj+Nuy5JE4UfNAxiohSp9O5gmOM5Z8B4NI8/o9cRvoUdt2fAl
T3jR/1oQhhPEx2rPdJYVa2/2DGbjPs+HbcR4A+rGv5qV7vK8c+eXPgenRi12gyFU
f3m/bo79GZARCItl2q1bff3nTTNt/k4zb2KmPuyhVF700XPfVCuX7xeeq01fH6Jw
ljDWbkSFBSErwDaDgnTcrFpd/cIQ949p6PRWugarU0ApGmhhlfUA9l4GaNYCP8+0
t/ZVdGxzEjRrhO55Hh9dQxjf1cqVCJIwiEFp6wRx1Yi02ZclPSJUpgwxBAT9iwcW
glDzM4PN+imfjc4LoZTBVAy2KXSEdFY07Ag4Cmm54mh9iCx8myn64CBI+9dl5nv8
R6J1t/Wk8vyx5m+7Xz0/OJGiU1iWVxY9vmuSpjmIt11E7lQMLyiNzKc33iT0T3qP
GMdDR2gSLt9r3R86XFt0mWM+98E0rVNuBE/AeaT3qqivmbQtDsHbLSM22NHC8DEs
tKVOXfDhmyvWHJLniREgN1KubiREUQJXZqrGwPjaRxj8wSJwxC+UwKm93Vo+tNFn
NOAdBBW0QN5ZTF+7S0cvOeQXXb75wgeu1Z9yUeU+QRTUb2QKBtZsTSKHuNDWXfxc
MYO6kILuPLumPqWL/OCdAcFukbwEQ6VntLNL2tTmQsdk4ARGBoapBs0KYaPfDxN/
bLr5N8dSFTtskLgzLx5cBDwgpLvlOLRgf5WmParlmGCbaTyienwXVX4PKo+eqbqp
QcU94kf5Fp23g0Z9HMYFHzI5xpy90umN2XsuZUO8Wbva4wT7PYILOKG3R9sq6XVR
v6ZajNzOpCHZjCZf/QU+4O9jVFx4hiQzFsy5/cszP1ifkGjwKu9fmdXdUpegRC01
aRhUzVmXdsCP2ZNILCCpBrh9yyHO2jhUAg8WIrbJayoqaYpcpCsuiaxk3WsuHmSn
6lISDBOKbWWmBpsa6BU2gga11Hj/zczGiwO7ECgvVz+G3zuqhy2Bp2FHrUy/8Py9
v7eFj6052Tvtnjh7L3MBg17wJj9Zj59oRIxDPYS37L88dqF+zPtaAOvcHd8KIVEd
fqvH7Ws2eCKR7jNuQxy5VYjdHSQiZ+mdd55AWpODRYNWaO9dWbnKmrSRtf38KXt3
zgtGK58WgA2QW+6X4kkbxPKfK48qIP/1Rg4RZ72KvmuoZC+zvjB2Zt3Y7aKqWjjn
MpzSyED2mbpug4pshXaTZbxnSG01JdS7V1oUyneKDybEQr6PuM0SKw4+D+NrZzw7
rkM+jh7ErdrEuSv2AM5v++3Pszsu0vWhD0JPMG6G7Cfk9lGCUU6LHANfh+QRRhBQ
30BfdazkdAu7i7euVAUBCganOmhNHnZa5d604iCUvuU4thwDhVMSWFMTaKCqBsBp
8F8eQ9C0o+lrBM3YxozDMTcyHuMdHiJhhXynZusGI80yGTfs8vSmaoBiQOBBe1HZ
AdIDTgXUm2p2u7QWr/8eHy/5B3nPsITav6Yx9c+PjPC0Es6FHwTgQ/VwraJRcYQw
w9TH7rDi2BednbPRof0kidiydii6Bpvh3p2ObDFq0sR17cgegcsjm1VJtO+ecCmY
tCVte1ysB+EVNCxq7qFwe4eOdgO9H8pY3xTC73fMoE25G+1mYLDY6Mzobk0BlMj+
L1yBFjyizFroi9E7cw8YxJr1vc1KO3b8U83zmb+cd37fXe+Uc+Ccujre4CVzVAzG
BH9hZyxHXV3TKX6vi6aAJHGo0A9B5R0oOOlzXR5RXdeNa4qayrfa5L4JjNI0Iz5R
OijhIuvlHUWFXnUS8WtG7J2Z2kNHkuf2UV1R0Pjv3zti0VusxjLnCfAROL3qjjUQ
KuF1CU9/LRiR2UljNaqBDP9JhY1aXKqHkJQhSfZWGnwaXZVI/ROh2HnZO3NoFQW4
RsMYP5iBMilfZ6c9xZbpXU+GWJHqazNcPJxW2fy+ypofwxJwSvoIfnReDqYY8j5R
pSU/Cr7qJnYonI7Ai1L5exvfIpihGeRHZaWLCxyNS7UHOVn8pQf8L8W1XltF6UYm
9JsdWNhTDYEj3p3UGEa4psVL0b4g99miexyWwZsXcZvbSvplPITAOcTczQz8Lezk
ywSRi3GBB/RCOPkm9afuQQVYQuDI5JcySMDnpxGxYGnXxJNg/yQZmGvGwtRS6nUD
Ukja4N+jU0Z1ddOvAN0w7A9yudcmnc9Ief1r3NJ/CvFQGm0zNfs+OnIYzGMWyw5d
F6MUzIHqJpqP6YXFxR+CYDqNvM00aRIBrGJlYALor44peO5W7DACDoDA1EEArhVN
k3c2GWFoZ9BsSuM/iYb+SgLs8zQalHb1KOzkWCt8v0sudvd+G9sulATjc/SRJl0K
cO+eZ1cYTq1CWAuTM6VwvOHVXBYA4NICD86Wp+u2H78ccSIb4BPKfSi6hWIgDHK+
6nrWFo77zhMR71//7CeVaXBU2VbwCgyShaiDrOJV16uejZ8H2XLj6Ca6vp+2C9s6
uLyBd24ZpbuLfVVik6UoRhOnbfigDHhSeKhUnBuIGUybONXGsuYV0jv3hOTh7VgD
6bzrlaYSHWgZBN99GvWDgPsFOgYOnNlg7W3bMAtYc/FinJl5GK4TwWUTGkXljFce
JAqIuTNGKroDETeTN3NTmbpqu4TQWy1Wiai4sxH9W4H3jelHB8dilivPLeQ8U6Wi
fNll3gUPgisJTUhRBFYjmnXlk2pP6ggf6XSDyDhf2WKGu9egbWNuAF0BNXq5ePO7
ARDraQFkwcPSvETI4+QDsQk5MOZ20noDmaVwCnGhtACekV0ivLKLTKaj7V89We6+
P2dIsv9CpRwgFzepVgQcEZnBblq1PIqWdWX01LfqNegf/B6L+heCC52I2LEasPOO
S6u6Fwlkb8zrKRIuX16cs4GcOAQOJpmA8gT+PwZSzOZA89eCh33jJpJjqp/aJnO5
0ekHe9V1aQvdWhJz7EsBz+WvVLveug5mG3HD2Dgzb5aipzZRNjCb4y2DeJs+C+Dm
Kf7KKZytcnPu/g7dX9wdYxdSdszwVbdkkvUAxTiT/K9bFSDS56mk3mWHFVpemcJE
It33O4i7CfRzROOli70wGsTMcuplT22wNBeQL2WOXcU9HW5T9ibK9BGyGlQ4PhTf
+gqLMFnwpx2QVKxP8kZBsbGgbK5aYYRy0hnbDNdUUBjxYOakO9k9ILEEg9kNLcWZ
Ik/EjbvKUyanmh+iaf1qpKp4u2V0nXzKkGUPgzQOCAuFKsKt2X9KDj0FlmGabB2D
mGLDqELDnH0Mo8Co2LIiL8eY3I/mRf5rcyglMyisWwiB/2RVmLZqdS9gg1r5EfK7
uyO2PZJ4tbzVZuwB7xSQ2f+rcfctpW9cMid7csBKFTZuQsJEuzDuw/wKqGHVY8wj
76lpDv+VnOTji98HPeo12stX5UKbZ8yhgKXgGjKliqybp30Ed3sQzpYwqNgo+Hjt
EyMTj2MMuGrEoNFq9XM73ye2xQFAnAleah4W2OnjC6eAjxDzqq0HlRdGFzfVwzrm
s1vPH6T93zIMtbRSi458R8MeR+pSgsnO4WyvGJ25BcoJT01g/W643Nxi5/e2z8GQ
VYfbz1LHqnpQDVsN6T8lD7Y287+9kicbqJS0rlXPs0kWnVuJmjDpwslERXgjdnGR
s+3biD93g5ZK6S+5muYrJGJtKf/mYMU2FFaBOLZgh9PaqTK3NYJjqD7EXHG9pfLM
JBeZv/SN6zUNYkzxaJFoyTr1PyHr+Dd+4Kv5Sa+EqS2DB8S4gbmXBIYJBFhl7zX+
FsGcKZt6Lc62l0HMtx8bJP/snQLxIvHchiNfIqW/5yJewwTbGw8p/PAPpIkDrV7U
yhA72juP4pNlvIDmHOtiGF61mn+3170FZsEvVRnZemVcRq8TWmb+NMM1tz2X6HwZ
XFCcjuxjJnq06nVtWlhQZ1lkVpOrR9ougtYnSPTaf5H6apLdpjE7XbMgdXCtvAvY
PKVkYw9FIXZ9DcTptWYYOwPkUHeAfCzxHeQUvmd2zen7GodsxrBncNlVh8SWtYfk
/xaetFp4x4OjwdgLm0ExwRkg8XiiJyiJ6PexdL+jVsOmbYHKGM/bwAQZc0Tj/4q2
euaipQtN5EjUzSbf0gKMoeyZVeDhBeW05Bg/smZ/H/PGVGrZ9wd8lhFjljGbFv0T
rb5e8lsSAVBLRslKRrs6F+jF/dd8VuFwToa/XP2ESkKKoEutJgmccM/JlY9X6hWh
7jow8HRhlX00N7Y/lxamfsyzX8EC+hS/JvCeUurZzsiYiUIj4H/gXSU3mG7cZewP
8bGgctpwoylEr7qXpx/Xwo4jOqPPQ/7vTXfrCCXoazd0p/t5t3+KKGpXHUqw2xQ2
Ay8LLlTCD5FuRGHp0CPW7n8ssz0xCTtcja+0qpLTbz1N0TnmMYWlcHKLHiwxsSjh
8MoS8wTtY5mUyVR8k6SG8hsaTYF77sxZc1nSy0F8B3OpvRvW6i6fVQ2N/ZHc8fRA
LbTGS8pHhDBEqXdWNfGT9V/v1//aVs0sSVKTHfBifUuOHeEhXLFb8W8ci/CtCUX0
chGCoXxo6vgjhfVeQl4xVZopqEzUuPebHnnKFo8s2Ge0CETJzKXSOBRycl9ova0U
eNWk38KTkre2Kl1tfNSgRP0xdAIKVPEeAyM21AWiAgiWSOboTh7VSnyqYxsUmIpe
jDKiO/UOckIAKY9rv2P51tVfwMHwJJqh673hQsoWjxAsnjQAwI4oibVc38h8KCZ7
2Lqt3zmcAJ6nBzeNhABGwRp04eshMowk4wuRrowARE/TrXm4lQ1xKth/QYJmMHsi
z5Wik4vDTXN1dk1EPF4kSXRCpJkrGBWLMFcL6MlD9Ed6ccpHBBLdzWgs2bBYuEI2
TZb4E7Rghvnr5GNvK4hJn6MmaXxk0UkzdS7/kFFu+IAL+1xCDZdZIN1jaMkBS8AQ
8YRXFBitqTIVaqIE1JWyQPGNDkYeCRoQwFR/QFAxcBxVzw7kR2EqhY75gemd5y3E
POaeAO5Lpfi7pKwiUBy0GGQ2lDNe8yTR5sctQ3l+9QF11ylnc6gL719uf97gRrL/
zLf6uvBMJmAnxp1+sCwYuiZryHJNTeYMZcaL3TSkXmlhXn3yGGxqYRmopLmMatLv
ISBkCYv6XWJ+JVZEUnzwaqy4p20KHgwcUscAojOZKCheIdTuNJvKlRaDtZgZSjul
EqZomKRiNtuw4afHmNlDjDFdrBM9rEdiWM3glQy3ftbLwXF7dOumcC1/eigQnVlM
dISd7BTl8kHIJQN/HcLvzBpwLZ3bXkRZWZ477d+G6gw+RRngWDIEl4W0bDrAD7wd
h6nqWb4YWiDwBZcdcPHhGhoes4Wp0KQFEI7Si2N618mLAbPSF93Eru8K35pGGFrN
7TRUAa/pXqbsl40ivIZV5wRivG0OiwOgavZE9Tv4t4wnPdJ7WMJeLDlOldQ+bPH8
p20JYfaasL3XrafTg9qK37FaiV+0Sz0rg/8ccbDQyQDVYN4ywN20EaxcEE8yQzfW
G7NL0hB7/bXteOiOlCVkDs1Bh7Yo3qVP/WsOkSH/mFlsoKBoxxuyLZIfyTSdY798
hxSzhCjsZiz4H1y8m2oarKKFZwkzvypJnjEIUzTU0HYtkZdYVV/pAuTcC69odwS6
rK5uulTSIAjr6uEzYjcQJ+hrBCFOSSoNxDn6hISfoTtJAl9StllpphCJrj8Q+Ln/
O/geRGTibdvO89u5Bz09CEN9cQBXvJR/593wLDLYg5+Sh99zVe0JQLXE5ybY39Zu
HZtBwP/IpX0ncq2hpMeX41h/IJpY1jQiO6r1LjXAQZaiP0baYBXY21RbQRn3ohOJ
6Ifj7UIJm0mOGroQU+3wWwBXFcOZdW4l/7WpnNjnUEDaTmdJ6SUNLJQYUrzpnmq8
c8k2xtrfHrhW8ImaMBaXjh7pGCoCmnXKlGsGId5DAvCN34ugBG0WuHl8bJUmMhQM
gJCAl6ecr9S4TqqbX9PnvMC+1caUQHrYr0ADCZSH8cfgiXEFT/U3cJI2SZoa7+p+
TnLrWIDOGyHSd/iP9mdZgQiUfyR2lBWdUhbhgYOK+wz2XFDx6FiHKARZVuBZp4eq
ubDI/SIM2HtKT+mh/JRwLYcWoRJhHyUlu14Q84FDn6mPbPqUEQyx1my1Af49tWmE
h7asMgrM2CGod/VFTX0yTGp8aCEQkf6o+kVM9AdSMtDXW5Z/7cj6qEyorEOBb68C
SqYcgvQC+xdnvQh1ZwuRmz4r614DlPy3orqlogDeyk7glMfwA5yf4zbrkVsKGmOw
z9pJ12OUjgo5aHH+bjxkkcV7UiCDNUW+9wttWST7QYXD0mSjowZ8/XBdpS9oNHxb
/kfbQOHpgfoQMVb9YR0vQ5+me2QiKi4/FVdTDUN2Bz9VSA5tQHBaQCu4dVN65nUi
0kS0EOFtsgKqsjna2rRaJiFsWdmMKxK700JB/xMKBNQZQtng/FL/NIwpMFVHxcjW
aQNcWSCrd0m163aboVPGF0p3UMq68hfXwv1sAMv+HFIUF94VfFbATQ64u0XR9rTl
hSyyLUREs4/t9bK0e9AImCTWJFqBD4F1TPCcnc1yZZBUBXrsfrANvq+5ODQtdiTy
sjJ4BDssMZAAvUy88EXTqoqkYdUTtGWcOr2o7rwB8Geq6I/Rb1VsCAy1xn2PBmvM
MBQZHIZjLukVcyrGZrAvEm2NYwdkJv7EMRSbcsFQ8gT4P//E71VNEEyNDVG9aLeC
hbjiUoeKF8vuQRLpRqEn+uY2O4X50kyb+ZorNxoctcOPhTtJoQ/HqvFn6e0SqkIw
T5L6yOhN3NkvZzqDW4qlyosqsuV5B/RWgxzpJ62bp05XDkwQxhHmAbxeu2Ocl2oe
4LA206ASDKCHB0kEI8uUtCFtNKFO3MrKSZ0BbxjE98mmj93oR5MIfq3eBMaURBvK
nIzU+TbAZ7QQA8mZ94hIbe3oPsFNnyClZIKIxyxMNCMokC13YsEAeqcPRWyJCovU
VnY1oAdribaOyAb+rn4ggeXco30MbCsNcTwBChwZecBB6wL2hptlwdErCuaX6DTP
YhktdcObVRg2nFBaE9mXnGcVCESmMoYaMxxFJcz9wWPUl3ukr9fRzZPOCOA42Xdd
AIzcc31CkEgSIfUqQANfbXtgvKI8iJJ1NjuSVppHRU6oEtKe0+faTtEPiQ/MxRGg
3rOzuHm1qZ6kscWme93VbamHiqInzMQ8HPvzMqoBLK9exDuRlcC3jfAciLiNIFH1
cFYWe/TZSxuqUwWr0ZTBylqSyXJdOmei3lT401uCm+73VDIcTFv8BPTHZRXn1ADC
+VUYAO6VwkbiIf5XxGRIe35/bFUybv0jePPh/9NQgxicHkMeEQHWhmYa6cnqwbam
A1qeL4SnyETA72PkxcyfEGT/TpEQ8QVa7pVlEmG4qOUGAFTsVHXkK2PGsMv5lAy1
XUskQ/wDfNaH8zQDodqQd0ghWGcY3/1esizpLLHxzqumlJBBRq/aFe7I2eS0G+vJ
sJymrmJVkTSPvBIpvXihprVkTb0wp8VKKH0iCV3ThlMCT3Htl2DOZV336tH09GQ1
vctKSpYN38AOTbTRLVcy1xY6kjJMVvtWY8tqe7N6qHH18q/i3q6E7K6JwFImdA9P
1D+o02BfQntvcnB5xkA5bQzYld58b1f9gXrQEsx2hq2zLtXByuZ8chXTpFkOYs0v
SwMjL9hTHYAjNWA96TF2ClIAZjZrvf4Oe7gLs4YDTrnOrEyPbkVD80q+3yC2pJbl
ImwPIe3DUmQvC86tpDbnU+yn/OtLuplFMQyAbxAtB3HcGHB3Kq6LT24I7lKHLXSi
ZMLirREXz+Q2gpx3xAxpiS8Prl+MkUEaxOwolI9kENkeYFDvyZq9OV5G33hcoca8
1J3dKuz5GtWCtOKW/nuhAAK9ANWcYkdqeBney02kaCIegquswx7T9OKYtApTahLS
o6k/1rjV7bPgFtKex8rqAINFZpmXzYHG066izEGYZeED/liVo7xGuHPltLdV2y7j
q3RKHF6qOSr8cTVOfHtnYa4wk5VCq9vB8Xi1AUKaRKxcrrZ4XIToYKu9wGNG9zPC
YEzsQLLlKBvbgHqcLRVjILZsp5Qv4C9YBN0HNeOn4cCxEGGDkaMFu57Gfp4E/xmq
DdvnvzZ74xd8vfnUdsXIjiPpjM2qFdh/4FwKwWbGaXmtcinuDQtkOXMlIrErJr51
byPTcyTWx5QepVQMmmxWo1Nyzq9jVHriugzEpN26KEHot4ipPgvpHe/clkc7+coO
OibYGEF+Q6ajWwOf/IWR9AJ9etP4BzTvmPqaz04y/3KiSF6YDc9eFBxNojZZBO41
5BT+YWFOAv4k1HcwFzNZt+Bp39liOdoRHVnCuq8/LcATT+qEjfg+NgBT7ERZtTXe
i7PRJWtbyO7Ic6tRWa/TYDiFdlKJICC1tUqpMuylhlIIWKJsryeai3Jga7DotOB1
+OYXMuCeHUpz5QUBDGQaDOoesH85mntWmKTLJo34Gg66GHkHOKis+sr8aeFXT2St
9SLvdQ5p8L7EcXjLEiO57uqgMkezG/Orhvm1VgIHC40WDgUf3o7KR1qfuCbAha+P
bCrgW0iZoobfGpR09IcV4MdY0xdHeDV7hHKJW3AKR2i2rvq/bMcPoD893+8GVRBX
2GuKXVPzkYoo630xuYYFtayWkHHbsUIDyqi/4V0neoMW3qvea9kqEhyf38noFXWI
EXlt+qK+dzfHwqzA2qI7nM/DIRrrCfNcmYENThtjIdAV0C+NBU/kdAcAxJmqKWHO
WBXQHlkF9d/Uj8DzFp7GHTyvZmoimQm7AH943gxZlTWphkvPhtt0oGIPrvAsdIq2
SvsSWR+pFwWJw2rDuW8jID5pgNtKFzUm6JxRFx41c4AyBBaCOT6pQTm9NJLqOmKP
+TfVWr2XPLAKMkBCMcfxIzmGO1KITejNfycVbDgOfryd2dT9/oV0AKhsvKxJVt5O
Kn/5gexxb2D2veUuov2Mk6cYqfm8SQa8FJGpiIZ/rxYpKRzUmi5/fpG/XN8JzfSp
yIvRg5pzeZHbIP5u4t/JPz5l8c8WRwNnWbSs3IHqNIKu0W4oVljJTtU4s6ddYbBI
emS2AE2LgaqudcdCRRuy/qDwin0eZt5DZJSbecqIY/T0NuPOiWObP4KqqOwvo6+l
jqvbDoI5b1fcvUVIrAFREWG9xApGzmPXmL4zZZ+nrca/KtppQUZUjIj0eNyyqCDG
6xDUOEwOJUG7DkEzsNuW69vFW8hHgqPwS5tKuEm4Or51Cf3VlRz8jsOqpBEgZ44H
lxpNhpQHfGYTINzvjSSOti1tLcA7ohRsI9n8cJaxom9ZMUNvjtEiv+UuQBpJm6+G
peUtdY7rre4st3l9cJF0NtGiv6aKP3kfNxA7z+DlhBWTrD/BSiRKV3OpxS+IjpW9
//wnpdC2wN4QMy49ntPpzVHV3tOi86+sXkRdncm7Olp03ALU0jKv6YkF+hvYBs2Z
2DuaVTu6jWpjI7epilGmL5PHdF1+LpfmVy+3CkjtGYz1OLwl1uMi2v7209QvdrLK
ltBqYpSVfGfSP/PYk+KJ7Or33eSlnYL1OZDFME7W6mVZ6efsoieKkIRhexFw5PEo
A1Ry8RVggo9kQSeLzILnLJc+p5pH/Yv5kNNmicesr2wB+hGipakuoZInJgK/ugCz
B7omjFhpm9y02e0TGN1FIJpu8AV2os9ErlSBtIpMgvBaHPSxyrLKfsJ68nPVskd0
my/OhRNUznrQFZe7VF2J4On2eR9B37n15MHKu8wyEuhEeN2ypEQeG/fBoi5O1HTU
3OfLjCgUw9KTbX4r56MGePyQmiu8T2AtBd/3qlDXa21kL56/QQl/mNuoNd1+VPE/
uUxmfbfpCXsYMJwoiuFjVqqdEzb4ZY7ra+vHZTdUltQWvWPnDEEP8sGqgark/QzZ
pQUiJax/HvVRD8qmaUA/r5INUNVUuTbAHuGNu1xkbKti++TF+qJNQB1TpP15SmYB
+D3mo3UVlQfm1ycdk5orkuWKsINbj9wzbUNbwfOg7AOm0o4rRDv/mIb5pzScwZDT
jkrv6TocZOM/7pwkJM5DlZXAk8DTWkawats3FAEvXTMqXoOuFbhx7bGZs1qH7TFw
9aTH95LNu6/5I4jWB5NXPs03RI9zy7h0Iu7fYnzEgDyr56V8kle51+2fGsliHk+r
n3Wum9QtgvknURAHh3hOY+WSw/BlR9FzPZHPKgJloXRT26DJQzlfpgGCAk2hH2Ij
TSp1cdCFZ1d2kVU3fcj6+cjjV6rar8vcosKbalfCYtrIrquWseMGV09D4jLZ0lLc
MOf3qlhFnC7dMqA9oflyA9wswzGwqGCNZ/i4MGuTxlcdCmnJSuygbooWxhU7BqLI
ZiAVVmgb6hw1SN7EzCthT/QFpwQLTClK7PP96eR76eu9uQGd4TDY6eApMo2Ry5eW
YOw6esPk4UW5d1SJntVsRlwyyl3K54q08KFDK053erEnjkQoXObWtJHFbVDON0Gg
cs1G30cBBNmjbWo1dVLhmhADmVYAwfrMe7tUZZkNHgvbQEX/3FYJ4bNe1RNeT16o
tImYSit588b35/8sSpwbUgdek3bLSdh9TXAyOLU6EVFVGpIq0T2siiTcoItJs6Iw
jprTrK6H26D+jst2n5WPTUCjA+fSppSBMK4AjRy5mGjlH4HieUy6y3uG8eIts76q
GFzrPLY21RWYlnahVXJp/uGZvgjP981LObYSoa0vICMX8mG0WkvKm4gFPs+aT6Vv
GS5sDV6RKuHTpeHkvS/OnOxEEYLTD8+5BEjKV7odUI2A0qsXFYpwDbUtHP+X19Bj
cs/gUStvvpp/8s5tuqO/z6458niq0QAgjtlBKz8pqA6XP3h3CHwQAnL2QYQh+KKj
7mBEHpkfwvJWeHMGYa4M2+5JbhronbVCD0jeSrt28uNvlcilbPNEsewu/v8yF1Yc
UDOKnuVqe1ZCOXBiDouDFlHLIQJ5jksR9F3mwWh0bUOkLubuTmJPpP9WqbHIcqcp
aj9yD+aUAFBTqtMf1R4q+k9l2QaNcnzvGIr35g+lyBKrW1gyEFySbA1CqbuH56ba
3PNBVpNyLmJ91B9qYeZKaFbAHGm9FYKc92N7ns1EUhIHmeAXGdSH4Bbxg8nQ+ofT
vC5AD7ihV4hb4sEViHQYcJT78svOU4tJVo80jYerJeFoyF2vo0kypehusSH3Y+j0
FptWG0F8G7bmhm5EjJs3/rts7MsdE4t1zmrUMNB1t1xMSLpNFTvt4FKcrv6xuCc5
Xk/oOYqLxSSydqgRr0WCxoCBSfr9gr8j3GcC6KdOOaZevUCNk4Dp5ltjvGHILNTx
sVLUbWmAfJVqer0D3CQfQzePAmFT4gLBVt73lLyt68sm8JfM9xIhHh1t9FWxmQkY
DraIfr0HwkfOEJTt11SIxzBK1YLbv50SBI67Se/jAJtmJGB8Bklz9FQI+VTVFLNR
IsSFDdPBTZOcXGS4GjLK8Lw0BUtVjHoxftQzaWSxNSUa0ZhwtSwuC0P1d9KXzkyo
1PGg0lOkUf7ar6uRAhW4GL325YGWn82YYRFMjLSbXsaEem1H+8IGeXiiCS8A02KF
gjr28uiIrujS/yUpeT6rgpNZYfE5tIkcSsLX8OlN5TPSIjIL4qApb9nUHJIoNAxe
FFXj+Qcq1nVPB6vPqBKYqyDYju1qTblkRE8YvODwf24DUiRV2qnlcdQsTheXmrAU
GTRNfMm9WO+ko7yYtbq/RSHr0HrQ/YO6tCllkOGg1zNIbsRi2NTGPPIQhtYAKEix
GsYCePk6lyzkIBYS8Qp1yHHPlNhhsENCOn46TbTjxvahLKLh5WtlGiJidmET+hIw
Vg1BbvWfdN81lWwgvs7HvmOiEsMpwXU0XyqgIF+1EzFMWmSUOGfrcA6ZWz/j0GFk
4IKjqffkdBspAgRkDpRJx/v0pAVaIX4nh/v2iT6/iP3Usigxd3b3W7GB9xRvzIFQ
4zJfPEzyWz/WH4l5lFfXHdu/0sSkhJO+Si6w/1x5u3uuBR6v20lF6zQ3wwwtkc02
2oi3ap0JwKLhCx2oZGGVZDFumBb3Gxx+yPUjDVvzl56IK5kI52eSfeJr0dRqkPFJ
M8mBqvfXIJ5r8UQ+vNuYrnkcOxEgGAML71Du8/gPAPfTJJLJdko0MnXyXMMLUzBg
SPTAjRhVd7MoNSIXUcDpvBKZZz34TYlHkvH6mX9sqlk72PwTCHKtnEvcCEKliLrT
ARAbFnu8bsmj9H/BDhKpLQk+oMlpxWReSDiIUvyAp7cgg2tRUfwNNIWzm/NEX7mD
+mxS3qbwYBPRUjPk642s/wvy4ia6JnTWQH+9wYqgbpW3KsslMLIfMbuwpAw+zbZ6
2Bc/HyEju0ZIh09r2rLaMWoLi5Exk9tv0aWVvmDo+HEhFNOtSAaN1edmitgXEzoL
r2MzgdKLfOZ/oORLEq146oPPUskSq8jsx9ix0X37RCvWhCqTxIxaZG7SsCd1H0PS
YaODw0aEnUTpISvjjTMemWtz+CvRoubXnK8NqxQUsmCivHBLJJLK8IJKmK/UMUqs
RrdJp08G98H+unQhqGCfCJuHpnG9SdqHGPVlaOUjfYEtnPR8huNtfYU0aBNZxx6G
+dIp+skPQyVPEBnYJzxzf3Fa4j1dFVk58ylSywRGsK0JwJHWx2rsAQ3xsZUZ4bri
RbijSWXbbYcDgiYAKRDydE2mKfV28t091vRP9ktHUONZLlYm9YhYC4J7n2w6YiTn
K/bEdn0e1oXMb1nE9AnJT80fVcEuIsaDGTRINxtZIh/T5c+kQ41sA23C2fYn0eaN
bwHzf5Zoqp1CNiBpwwB+9CMa5ho9cp3uteVYsNP90bbA0tXjdbx2u26OFXs7erWu
TKqHaj3qSZ1KmFY3P9pqF7xofianKeQU5M6EaDknimg4Djg5hvAJQFEBsUeLyFHQ
26UZRmYWMKKyPPrD4p9Wh3yoCLS4ShS88ZsG8XYZh3K0uD2dnspSE4lpORBJ0ht6
xozASY45+tepPusoEPhN/e4Vr4BrZLo3LrWaF54B63mx5/IvtWZwhxX3ztqVa/yT
mzyiSSi+Or3OR+d3VHvIKNg45mFfKlp4vHObvbHRcpME97830Ffle6qzOnx8x1Uy
PH5Z+wgkcgrsfIG10C+tubh0vpElOnp/VoczuzWZGzddv863yyXddt/0H9ERf1fv
2m3FmynnXgMJhobIYwVID2e7X026+NuhsXAqZUFIjPaxBHCFV8Gvn4MWw5vqZzW6
L8PkSSRtSmQxmqbrbcsTPt2FNenfHqmcJ+c3eytqB072tIxDNNv6W8zDkFlgAqdo
tn6/sYEBmeVYJi0K1m9+hqYJRt/J2Ea6fdqVsXjBJ147xs2ly9+4IciFYrFVWPPU
xTMbK219qFgr32Y2se0y1l/vei5sL92JbSfdM+/Tl9rKayQM+Q3lEh3OsR1+uJru
FxWp8Tyk1aCirfdVh47brUqhuO7Y7icOTMHZNi+GmymMt26pKLq7dwZ/e97zJk0r
lPSdQNIRya5ncR0SVW0cuFKPCmjmzV+vmfH4HRiBGLMuYj7YUE/vNIig65T/0i3v
9tC8P3Dr0x+oOdJYwRPy48wPY2BRvd9XiCkZbhRW7IFnovyWNWSOq54xeGjHvi5d
0ukW92sxLgBiVqMei5ow35/8ug/Y4D6ia9CYj2RQrhEV/mW9c547Q3Qc0onqJTyF
78/qf7bcvcPpXg+w69kE969df8GRg7AUXEIXSc/GfAFRKLKfGe/GkKWc8EW/yOj5
KYSv0v/FvQPgLhrwPzN9JBR/o2cZnMabwoDu1C5rK4ZTZQTOcYJdjWt0CDc6dpif
iC+GbNzantenLOXD96xkNZo/MxggYRrURoVKkjjx67lbaYf2aZEAGOWZc2BmsNuX
pJ4vxZ4P+AOIUwV8xhYfCbAK0McalEJeUpu8YQCnT/5Xt6ON9WcjZjBTJQ2blVGS
m//BmhNgUaQGfc9+cz+2KUPns/u/gQJXHxf9VFGMYjVLZOWcx53jVFMoBXqCtVGf
oeqAKVRbgggdPZBgkxKGIubwRNRJZby1Ee8DlQQJKyNqQlyiSfObVqm/BRdZnsd7
vpOwSvsv3GFSMnLMZu6NZfR5aXAO6+75EuyA6Vl5ZX6SgAHWh2GbnpwfehHWBv0j
/uz0RCvCTX/Uy5FnEJxAYNeU5rvPJNFW7L0TDQJr6YsUAhCAAeqVA9BTBG+Ux7sC
Iu1yb2Pq4Sd9eORRSIqLuKVL+RiRXzz74qiWTYIYrluBPqNnXj98HmVkzsAy85G/
on9hV36sjVYcqxZuhIev+P6uJJjt2OY7d+j/t6IOoBToQSi/n+zNgzHK3wCKQXho
kLbtqbAcRP82gDTSMhc1EyCRxXrM3PIVAqNznkQWrF6Sg+UISESFlWEGmjC7QFjs
i9fkzcBfOnehtSazGOAqwnGBfu44XE4KoQ55rBzHGyNkuPMKPBE9lemHpQoWdIst
SEpp3aWhTBfd28a7/2QYehRpMsG9Ri9qV99B6up57LGJCsIEnqqt7fuviOd4YF//
C4HUM4+tLWBvULi2a+vWZeIqxA6OACG+peoxjVzmho9mr3RKF2KbrHno4lk0sPPV
ROcppDppo23RehfVgsFdyrrI+hOaYNy8DY/GLGWGNM68A5HzbTwUk46p60v+1qGf
j0gl72NkFEdJhrWCLlOietUAzv4RiScNli4WZTHQ/ubido10SU5tTxeQxXC+S6Sp
TWLdc23O6OctqUi5ToRPErqv+1hFsEuOxnvstC6hbseRNao17wQYkaXpAbG1ry1b
pJZ3goHvkxeM0SneTPnuFbuvX3HNhIbW8HUt6NSmmuzGnisHlSJivw6Dqss6lrO+
3WYIKn+DVpGVDXs+QrIQc+pNOJGT0qtSAuL+rjsKS/obf8MnMG1SiOaGWB6xd237
IVpd8FEPvks47JGmkO2lmHqiozyfUQVXTnvN5nWJxEp3grRysf19UR7gH/YYTrq5
2DmjPxiYNwfgN4EqUW/In3iq3AmJL+4X9D0hth89Eb4VAaK5ZQiTM8vRKOIkJCAk
M4eHwvl6FZ7LW5EkOYufOZgZHdSa3AXMdaM9K38lZaxJQmTTKVyDOCGYlk0iMHau
jIuVV+pWfhOxSP8VkCvO36y8NVdGcZ7kJWR/X5KsTDc/2JQKP8VhBz018WMb9/ad
noyVbptnluM2fXAbUMu+ZTsYWYUjkOLAFSv2bL/Td9QsUejOBmUo410P7znVHa5k
228XTHFGdCzXXWe6VdvRX4wfSmGIvHgYUNw9mjC887+SXFrjGywhvk/RmBlMtulJ
WJVjNkPG9uXwGEyyUnz+Y8WJlgcXdo4exnqKNgyMT44U1C+VsKSK0ExUIpvflz1g
BbNwf+Bu3ROjp4tbfsVzZTTaoVeTdtQhxJmoGEYoXsgrfhu0ANTBIwKRCSZcTFf7
WXt7/yZwdlQmo1azEvr2jZ9SyR2n0Dj5r45hzS2BBrjiMusNm2MtFKFx1DNzAaS3
vJs3VB1h8bO/OtLg01BRceQGQWz7hFWucMYu3y/ZlT6T+nccF1m7W/5gC0oFLhUR
wxq/bYzjNM7DSc1OC6Vj0josqrYYHX6+fUj/GogWFjBhIjnRASL4XYqeD6HSP6ay
SNjB7Yr1kRI//OZkyTp1cJEk84e+scFXpXfe10utcia8CcSnSxV2Ia42/baryX+x
4FzcTxExRAJApWm6zTlDfYR8u06WKcqdl1mMiLg6dxkupj/FwpEFpuhQAk52qBHk
ykV+reuUSRkEZSUgFZ4igfnF1jvDqCPD18HTxd/dtUn1FaMkZhxQhYAoeCC1+Yy9
I1utGy5cbqysSHOUNW3uaw/mtLpm3E0PcmpeVHED7h9n+/F8KgHtWNLQ6ppHAAvk
+eRwxoyEhL1pU1uw93OJLlzCZjc/frKnn5GwsBfbBA3w/30LpXa5VSsZIabBAjkG
StHRadvMY2DcNgrNMlz/Dxp98t5aFMYJRU28UAI1nkGw9nTL3jxMIVSgZTZcQhto
VBLa023XcyvxTlPyfI++eEl0XNRsVmr1JMLGK0tA55/s3F3SHiFLSimHs0cK2WKC
g/N4EwsdBosZr32mZG4FIz8SLc5gZoznldrsubzyXutXt0juahNwD6Uiia5P2scg
5Z0Iz7q8uuJTW2IIqZa4ALqeDHTatfbIClSo5CA6NoGRE3Ax0nZUF4poatzMbaEs
UunoJ3B1AJwvZbGzCOwZeNR5wIvaB+7bOVbZdCHbp5o5Ps4wVUBGgnVMVPUNFWhZ
tO5/Y3x5ArbKUJJ8fSElVCRkgUuz1vEinjH1afcUr4qpJzzkgwwpH/anSEr609gd
v4vL8rTeox9w2tD7zQDka6WkkkspPHdG3O63CDE+MiITdkQ1IW1s6nAKbMRJURZY
fHRI4zzJ2o9AlnatdGfuSEMapPWwXSyCbL3CN1PdmDYiVOrjxh23HBrU22CV0KfI
Dg1r8xJRqr3RRZwQjUKY37M5z+jTafsxpdMtx9IZbsflAPVxf4LPGbVD7SkAHQDx
lwWwz4d0bMgppU3Wx7b/mQCISJY5bQ4iQRCjn3NO8cUPL7V5dbAnGDOgAIGIIvvF
zIv4CJD/S7thfF9ZQ/vTyJRHsR6XnWYLtqCOx9bXBvKOyP7KZF4rNPdWzNX4KwDH
7bsdMur4igbubu5m50yER1lEilkF9Y9ySiChCUZDsDXDxvIg6EB6uXlwu221yqh7
KowFELz2lWNxdgJfSptL9xQ86YfB4MAjIyUJRTiyyqBY8w3gEgUvMzykwOitsT59
B34b2927KrVnJ5gXb3Td0g+axJmILewGX9PaoFYn8Nfr5mdDkK5zLseOIwwz8Q/C
vFGuHNAKb2Pij3eEDW/bbXvCJSSt0SumVfwnxlpd6KJEgA6KqAGqLfm6KJx64pns
HzC05g0Yv0Pvsv7Nzlg+1zO0H14hqOkJRM0Myoh8r1Ri5463Vm+LmGsPTGRvdX1q
qItxnxFhQ9+TRdjxovwcPhfNcz6J9Wmn7YHtBMjMY2NIgf9rMhO3UWFZw4nU1Rp0
dc5tF48Db+APsxj7A6S6PbkctgBa9OxngBJKT7RhwI9njTNg7DB2AAYNQAYgH2+3
91fb80mj2BmGC7xzKvB/7HeeluQMvS4utuLHUPzeYl6bcJ6FKKIclJeS5R97o2GS
jBymazCUqCdCKFOv88c7inaPfbZihTNlxJWAo290cqHJPI9u7XBlJN9IIccgpCJX
O/cooDgmZ+RS1hdRLM7OGy8If6E6StG2OGiWKrSlqkz7zc2s4PNz4fEWoMN0jBmG
nvdgaFJIkNhxix1G9+vBiB+WOH55Lyimh5rRHZUD4SAXcLzZ+KN0Dg2CKphl7zus
eaXiNUBcyxXo1pSZF/944v1YWBiVJdPEbR+MMfF0FizsVEeLl/rJSzl0jofV8wbh
yinI/XAfxv7BCiubJToDnSf+lXF3fRSV5E4GxTGe3tjm0u0kw1ny0xtUNkxrUYqs
d/vqHJTy6tsw3RaK9rWXdkzlBfIaD7G6OpKWrA0bNj69+Q9okvbMmk0EzWTZalZU
IBGlQb1xPhfzPgDkiOspTHz8a8E6ox/c9u35jSCkzx4o+iuU6ZgOpKwXKHj5VhcM
CTuKAbthlXRwCNBaOuwWnF9mG3PdjQYvWFjUJH5U3kDGEXzfPK66AiP5mhsq/ZzQ
izOthGVektO3Qu3Xgb3IFy0e8cbGIBORn3ls2hxj71QYYboc0gUh4jkoiVE/GVUT
ZYXv6Ped7D6earH8fJYTmbnare5oLlaLqkqL/2N2fndeZtjt/rK97O8hLdyGuRWU
F151YbuvZXwd1D3agY9zsuXNBCR+MxluzCpLEcGk6yQq92u2BNYhvZMVAkvaPXxC
P6qfH/D7qT6gQCyJUDxXlE3FV3iZlew8wu6FvU9CK747rZt+vnpXkOMgGDyAOLD3
Rl+oHwRu05xtjo/UTvP0ECk2dzENRmYzkeJ9IAI6YipqvdxEiPQQk80st4ItucBj
A/KUc3Wn4Q9v3MibHagt9gF4JpzuOE7NKDJVh3EEkp2LQxFdX/sZcvTz/clq3Nlq
zhQs72bS0b2RVeAeRatRhU1PHZUEQ8DWkbC4zSuDXwQwKcWXkZpgIZ2YJzaLy8L7
RHE6PttrKRM/sZowj8Linj0Nxd/VrLBPdToZfV2BWdI4HNfW13yHZwNqk1lrmpXa
hxLoHQCdi3FyGtVy2JtnhnWi7ZXenNQPbXjGuz9ZZn0XbGHuTNcGuzF7QrfNdWXw
rF4K1J0QfI9ANamedSuXSbh+Zc26MsNqCTna8Ivz/j/gQYNt05NAOu8VjItuZzLA
/coc3FZ98topuOg3ziud3OyKPJG7zXZl8S9Koa79ev9XjGLILTVioJ/6BEXVvqmi
+n7lekrvhF/s9nBPiI0oz4+kmpR398sM+c4kjKd+pJIm7o/RsxZT9Y8/JdsV9n/0
gwlRg+OdGcYNtgz8MY9/8aVFynt2abc+x++pr76wqjOhBIO/vudRzUrC3PIVSPOg
KXI59blsL5KtLyD8KMbtFwuW9iQ9U8OK3FLlq6JF87blAv1/69w2u+zjJJ1jZ4ht
nwY21XxR94M3kEFf1n1cMm5/xH56wLkkDIPiKkMNHDG4TrqiN/67EVatBPn5r6gS
ahGLHhVXGP2tnBz68S/zixL/V9GzGsN7B2VOBEGuRJOSw/wqTVdhfustH333hkfi
IuHW4lxBjidSBCYhONQbSkOOLcH8IwN3sTLHy7rFsuraD7T86+ykqsxQQq3Q1M5o
12SAm8pwnG/GiwxCK9LJvanKX+lS+J7ea2sBck5FDaoB4Ql/VHDBZpXZ/g9GnxWA
YLH0Y86CrojKq3tfGPhGb4JMdWjB0rvbwjXQCQAMfN2FET3T8YtTq/WZlzxWudF/
PV1MR85CVS0pJq5F6Wmy85fy+YnY/L7ux62XHjQh2NG5wpmPNzpQ8/hVmUlDAaOX
mWm4XcsW7bs/A85jiqsbyvTzB/vyBFMDDuMoRwdiczqV8JU2KntM1Uu06dbsaNTl
PQimt13jN+b5agGtC4c9c/3iiyNKoM2T1AJJLS0GrNlTdL7kzcVJU0aw0OouE9K7
gq+11uJcvv4DjtBlQLAvvJX1dKn4GD4ENVUzw+sam4gsBnogl44tJyRXuCincv8O
91XwUzYiNTv/LUjDJDmez4myvpLjNzP0R7yPOoTr29RrHDN2Rcie87MAmlJt/dyS
TZxi010Lo8HNjJZy0HIYhInve2O8hY9Q6Kv5C0E6o6kgzVrNQcdi1qrcYjpNw6ks
W3fPhLaS+0i5/RKa0lB9ITXdwdkJgqXoUjgVFbXt5fWG+k2S5aKv0I2F+Ga3Jink
6Gpitl80I/dMC7MhVvkDFsshMo1unndOZho3BNrrlIXyaTAYXVYJZE4UNyBRRNKd
6swJvWi9sOUyLuyrFSuRwd8tQQXVbLB5x/+8l2Fcbvgx88pcWhrK7DHaD9TVSl67
GX2igy5Bg2BX2V9/GUVokl+6Xp3YxwEAUKfOgZGDQKWYMROD8xLlcfrSXHMnye/B
xIpTEPPs76Ch7M2P1VTk51LgbooGTi9/YZSMeIoH7CicUv/Cr6hgwVRyFgrQBcHz
EpJg+Q9n/hbMKB/N6ijI8w5gf+SzL4/nsr54jfB34PFq1h1As61wUFg+MvIylo/J
7HIHy0/KzPv5fLO+glgl8YDjFJ6SEHDASXbkPr3eeglyQtAQgrYpc/n8ihzr9Vby
UJOi0RK3NQjUtH0Rkb8CcL29Bwx92elcjMdVw6NWw8+xZpY6l5QZJs1XD1pe/z/w
VfRMG4AGZ5TllGKK28IxpTErC6DjaYAf8xftk3bI7gAclRQSNBMD5bK+QZdj+itI
mok10aVi4kMl/A326bBx+RqRNOU7nnURhhJ8h/p6UiPpklmaXZaqrU9VPWrm2VJ0
98pZJk7P4GZqyde/0iotG70W/kVzbZG7LosA1tDi4kg+WUK7eQ16V5ybS5ELF1W8
/sunPV9iVs5LqcPpaB6ux5SxEZ8MnV0lXn60qdNKuLKHDcf3uhRajQ+IhbQ+EZyO
hX+6F0KhvNLyI0FQh9i1EMeyRUnb5xedyF9WYp2kvh3UtASsP7qE26hzqOhS40ME
08giySK/EldP/EaUL4baiD28FtjMUGraS1c+V7IDz7zph3/FEiA52zEf51D5QYNU
OI0pFWz1ysgb5yCLHkW7dCD2cA9eck2lKF88RwQAhNbnSqmOtGBiM0VGZJNBFrnm
uvP+PCmkjqn1kBo3KXRYJgG7OEGzuYQyniCh4dc7NjWzSSPtYB4dbEB/Md0Zm7pX
81mSdpxqmR5T5H3LSFjUHzXscbKGOcYNRO2qnOVVH/uDjIy7VoL0v9Jz2NJkwOz8
+UcfgjxQxoqKZuCk5qXun7Mv1yGoUD3eFjvkBDp7e5HfY4PxPUHjPGV6AzCViBOl
gMN2AP+2VY3UkAmRw9LFAdKN4M0RG07pv8vaMnjddfBaxDHBo/JOc0kCHpdtR2SO
KcSXeFpI3QOV1tjhr94Hi3SyfWpYufYdVqPdoj9MNBgo1tYUjwKcJSGZc4EEswq7
vCqfX67LCBmH0E7c/edpYvK/WXvkBk8jUprAcoZsVbcLrDBAxg3aRtqzoPJjh8J/
NemXmfugPxYb/6THcs/YT5uP9dveB5E37jUSgI6/jKByPO+Aw1449JdfUxsjS+xz
8bNRZsErZmnxlwR69th0onuPsQcUIiSdiDJvlJSLFTdKFwvjKJIHVWsNC95wPHLW
+h1UnsvYUekKdWuanxkpd55rxi5QEMFp0JvdUq97JFr2PYjUvqV1HK9oLId+zpVR
XaXByesoPwXUBqgJyEUwbBVDFIBS6stj09Un+jiHtmSNJUy1wTEIbpMqTwSpSTKo
dZ+PjHWMpTAvzcn+hqKbaKCVtLCgqxuhHGwfvonL6xhPnrmkOxLH0rewqeyHpKfX
/xJA73cGTvxPAAIJPXPrUDepakrm3/hqpjiwaVX40m4D/IbG/WsfeOUtkYmg/XO1
grDmNzRvGYJDMeT8XaQkrijjh6r2A1RxMBortJUde4hRJLT2Zx72mP7U5wbuesQN
+wrBk/QTPqEHkM4QK3Tm8fGROZAmKn11L9FZHSmT46KZJtnKhwGaIokwOdVWKvM6
S3K4+YkDYSqEdwI37Y1gKD3/2CEccVFVd8KmseiNVuZaJp2hGnRK1uqt2QaOOZie
+7mZM1Rz+aJ42kZf5Gw/HGXYuHPsW665uyj/FFh3I14T7Y1z3IgYy95lyODL34ba
PBbk4ZB5M55fFd1FZk0g+E/DVdiCAer+xbG0A6PB432ugu+Q7JbBIIksQXXW1Q2E
7rtV4ZoG34mIz2RIQHdOnZ86EVvhLny/lPr93t2PFbeSTxvFPp5i/aqjo/0AEyXA
b/hlSpl9V+Rt3r6Pucep21Mj1sKwjMReNUqfZQRgTt4a+i2P4t84sXGqzA7XcWTg
HCF4VnVwHZfae/SH8h/cfTSA3gYzMje9zxbtxH1NNCdTsTwBnT8pLlbHW6Td93+R
7rCYeqyfrMmG2Sdo2M756aeCsjSt3Nuqibk39hO1SCdiNO7lfUJq/eR+UAFmG6pA
UVDU1Lss+JidN12uqBs2EOQ/pgK4y9TEVV3oOsWfu2aKuTpKU9RJW8aeg9D/j7++
mByadPTc9OiarQico8P8/YeQbr2D10BgEiIUFhNZnJQINc2+bX+wFBkW46Nyp6d7
+7UDgbgH4WfVi5MMZv5n0xCa1tMBwO8KND0vWJGf9qRYjXkdUjs4666IXAYKklD9
72B8vJUxOdJmtpsp1bYgU47iDaTrLLlzd8Lnox/6jpbuyUg5bDaeCK9SLElZeb45
bo8Bq/zrA3ezgfCMdoIGQhKWXezcUGdVQFC6h5ahaCN+C3PhT27ZvN91VHKBESEk
U3e1iO1yPeGFeW89ZMOPP71NrJutVPWk8gGdyx38yw6MPuiXpm2USoNUBJhsgXiQ
LhbtxADePX/jBD/C0VaZRjY4RPtifehPFZLnJ9hVpcndRicgzjE79LI+1iJRksTd
vWsMEhvf2EQZc9XHFLLGrxPprWAhZpu9IPFy8zqYc0HExSkLp6v32y7iZBI0uhr1
YFPbWB9Mhz0kOGvvYUfYgtSqXkRYN9t1RZGRuKaxTDweEGdi4esWkghO6jexi5F1
ANnud33q8wzT2yz5CpAJdTjOATLpjfdhC63Otb1qetmec9CZNA39608kxolIqzgZ
woGvWZJqfd3hB2CfJR9Pvtb86rNhboMzloV+Ax1J82rB0UnOyIToyEZwmnPABwwu
gqPc955Q+OGC3yXAm9bJXf8o8BNZdcn6TJ2G/TJPqSmRvM9DVvs1VIaVNJu+Kp93
fOH6XSBMDaH6uOhkZaxIV+lGolPdfhz6zfqOIOk+7KXYuEfyydMtfbWTEDjoxfE1
1YV8HOMrnbc2rOt2w4DJRW13uUlxvAOEkFZEWyM9ZIKQsjyWoR7+xcF1ek1d8gSj
rN4H8ji0lAP8WmDgvvEY7MFFQoFzwCusm02zbAi8UOLrTtF5Ct00Kgt9tNRgXquN
x/qGrULdV+pIOPaSXU6SDhvQ3nWvrZjVF8a+jyOkF84CLpavnFe8f7oeaIkBa5pC
XzTjVTxIge6vmaiPyTcXmlWJq3Nk0ifTB7qJAM8J/oC8C45LYN817TXt+F3Nkj24
5Gfev3LiJtA3H6mB0Thx380G/2NravfVwqC/rAqdLpD8IQ/rGaxJynOR4w0YlTBo
WoDbAblv79jL06Vqf7OMX59Kh5FPvwv/j5IfKw0o/yyvkIs39pCcizvOEH6PpjYZ
rT2MK3CWh1GnUhdRDwMbmkNfneaLTE1xVJn+SoO1A31A7ShJwUhYECrYmfpUTirg
E2/NlXr8kPIiZMIYGgLcDIh4oMbFYdoQdQSNEmfIvdIJsBsEoMaZu2ojSGZMyg0R
Xn0GBAUp9ByjBkX7evq81ERx7lyAJXCA+pDP1EnEXeWc8jCWL17cO9p8wgv+NSK4
HCs4g7xtQv75+iTIX5B0+n0VN0anCYbrTgjoTi/68n6gILq7eTDzOjtRFW5JeZLg
AsRijxawdX35PJiACtBEdiG2oE4N1rgsZ/IXJITG5+ARY3PyG31UGsJu646lNtBT
FuqaNP3cuIxoF4IBECMT0Wr6eMY8RqvQgrA6i/9ZKTOb4n4pUhyZ12tmStk6ehXa
WwTaXwIX9prqVj49VQpAPjITUxKEe0czecgBhHuCHT+t17pmXhvY8NAoOa+k7vVL
B4oVaI0m3O/UTAkcvhBd3d8mKK7/djhr/mmq4MAw3zA8P9ZzgqPSvDo39mdcWr63
94b+oR1kBgCc9h9NsLSph1vPsAa/Gm5Y2Ltdw7uOaJpEE1KR8ElJJbuH/FvastmR
bG00BUis2DA0HgOf5/J53SCeRp4t/yNVUD96K8b4MBQhRWQl2XmoWeruo2yAbdH1
BC28Fy0ND8MmywmVDVYlykeiiJMZhdLVx8Z2S6l+1remDlfi7cqTSlOCgDE6ExW2
g/+9iB3oMEEzCIHTlEsMI/4r3sqXIDM3Zacn+iyggKVumV9exkDMvndfbUfQt0rg
RjT3aK39IBVX/N9zlQGvko9cXxEUwF0vvmcOG3dy1XwsD/VcGnp4RoSjaH2Iuniw
ssz906GH1vAuyOD0R5FCK2s2/8wXI0RxM0H4F/ketEH996VdC+uQ8ZtzRejxVW7W
fhIVwK8EpL+cPVCIZ0cpsTVbD9//sUh9QmoLWXLeUXQ6wPRMzt1BZfXOfFJzRzhn
CfxUjS1dThgJsngiTQpzYpD7VL05L2XrCF2G0XgUhrOCJar3CMKT4ZYb5k4A7adD
xRdacl+/BRPGsqPNyH4YbC1ZtaPCx/AkXcKlnJ+894KnoIaiVIqM3GNflS/yuREi
mZqBs1dWHLTJgUmJSmmu+EyfwH/YETzlU+S2ez09pbixVR7ewE1DWfEbRlQjr24J
k/3W8KuDfeASCLKnn4CeO1x9oAUA5+djzJjv3SOdNLb+ccwAwBJATjRZVs0VG3yy
NZNuisPKR8tahd+Ea/YOykBV+gMORTieMoewxJgap/1aZSYumgPk8mr0CqcEkYGU
hJcU/r8HnMgk/Qo9/pgWwxpBGsDe9WM3bseXVQKzrh54Rca3VK+a1pWCJvjPYuU0
5zgTQDhiv3sOvwtgDCEfU/6aDLdLCvr02p7GMAPliAAE7nVMYnSxhsDOYhxiV+Ka
RyKqjCo7RXcTMYOAEvK5t0Tz7V72q5XijNG6kGuqgs/Qzw3qjOL128wdVnJI1mX7
W5UX4HugkmIk1m4KpGhs20tsoL4vyqzs+6eC8CaUhB1or12ZUGQ660IKuXA7xgZm
4ndWTaYlVUN/W06iFmSjhhDmNzuDxWwmnqpemqAJxsRgGptRKOMSLtTl9UMYkfs1
I6qicPJNrNLdWA011USDuNxpwxKB4hZB7zYEHgt0+agj4g1/I7Lin7hywopUtolH
28hRRGcl8Ehe+d2E+OxzB95ud3AmtozOFUgEcqVUmGInI/JII70oSrhLQuRDX68F
4naCVZwL+myrCve0wVQrnWwOfMcdtMICvp1tRSirN/jLZZDQr7lwNy2ivuU4cV0I
47af5hcrWy1+p+7P+XHk8zSYHuMDoYezgYENphX5JyVCFjv1SvFV+1Nc91m0Ilfu
cUEBg/iW9Arn5rdOaUI5gPjFFTysELkM1+wmI4qRdCH77of9NzqRu3x1QT2Ftk/y
0HKT6EASkEexi5couRFkNp4HIITvVmuN3DfR7eAVXfGJqRFcAnp8/ooLG9C6udlH
8OxCld/D9lUK0h0c/yeLWxiJl8x5d5xozRX9hxghmGqLFJu0yO+CQ9WHYJpiyZrL
XYUmT+SjaatQb5171y7cILL1g+6IrEKyoUmQLBLuWv4TmxTkYqj9l+4rLGlKJ4m9
C6r3kJRAmUDKqlbHHzrLDNi5qjUg6qD0p3BSNXeZQIIP1whwp1AsUjDqF/6fsqU/
KpNwj1XedyTrZxJBINx/V799NWN19nwUOu4EkinKaVCI9DzUtwBLkpAgMaD6pWxe
o4rg0WA2a0lSCv5kXpbhAqTF+4/isAi9dlGy1oOQbehFkvfLX6QZUellmFsP3hcr
uh31eElLmUB4TmcPc/7r1kRvP6NowFZsGinu8GX76ZQvGAk4Kt+n7QPj9mIvEkgl
POXP9H+maPQf6q1rG/9h8ss/YQmnBH1aGOzTsnIuN+HwBGYbQoYaTiAJU6QIs+cS
NiDrJBlFD2xggD7ym3QYGR/UIrCz5mGImcmTDMOUk3Lf6vaNXZg2dYC3oBfzsDlp
Lh54LahN0eauortYzIOqYWsA0jAeUrvN0Xx2Kf8Mrtswd8vusqP0movJCfpAG6Ou
2cKqeoqSvpO3vPukg9O8tDlUiMywrS/+ffBQoK213+hfDx4kJo/TeCdytH+tnRz7
iWBbu8SgZyuSG7W6m7Q/YW1Nbb5VK2Vr5GzHiY9keJp/J3uREtWGSAwd94Y8TXpW
ToOqPVYtHy+QFOwkck/tog6dHP7mrm6wklt44DnXOKTWGgpVhr0k0ianvCAVqKE7
XU9VPZzgg1meTo+kKX7raLl4uy2zOUUMI0kjis2z2JnIE1kC0lAhmEtSPt5/TFs3
y0HvYS6cYYY2Tzk2hQXX4QiYycbIF/p28EvmA73TyTLRH4oElnX/dKBg9esILxpK
Hh0B0pLPkqfwWNm7oA2RYOOXI0P3WQp0PwGaPE+tsRJ5q1DepYQxmL2tblQgCn1F
ctRNJ5Pl9E0JrE0D7HEjq5rpabJKVjFts9QMCJl52nLOqpS0y32nVnAW2fYfc9+4
02QeUgHHHG4MDT4dXb+TpRA5w8r68t7ldcS4IE9TwbucolvkPuUFnoGh+TYh99BG
eNzSfune29L3niMzGQC4GKvV/iFaXNsyOzeBZkZ7XroJRGHPlog1/NJu+cffLIEc
MX9dkNWihkBQLdH5XIvXlweASqggxIqUkEC6hDwzHEWIEn6FxxjHBT4IJkJmeXv1
j0ruKWa2FSGQpG8Nz8HWAJnd6FG/Z8PY42nFclNxdLbClEej2L64ThYnVPkJHNDY
lhrJhlfUfV71jIwM0y/exLFWvu1g+L7stBaohUZqkPCMk4iFc/eJbRY55MlTawTN
q92d4EQrte133r6AeiaXMGyiHIBlrqgvp2Qnoc48mUQfKPKtQxEsN12nQ2pL5yfD
u6pF7cvXHIwLa01XFL5vfTlvKjS6iRx55AJ/Na0D/nL01Z0S+Q5wHRgW1g3W2AoM
e6VrEvTPkOwO1dEHzraaB+vp7rtyC5OH/swr08uwlTNjQEypk9Z1p1JAY8FTn7Ak
+ByL/gNdtpRTcSWIL/DPJL5qgh4z1JAf/uzE7fNyRgkfS8mnqS6CJMQrGV+XAOnV
bxiI0RsobZe+870ZG2EotIw65VCN2DfktuFcaIUlRh9pU7rHMuJD81jgz8XdYCtc
/gurjJkxKUOWYh2PJenPRNGf892BhB9QSkcTfvatvMrneT5BBqc53txobufTo6b2
MeK69Df1y7LGg+7w7dk00kjIWhvs+XiRupatuKis0JP0yKK0ImDUlOrm4IC9D6CL
C/zuAjcJgv73hzCWxkmFBhHyUwdd9npKaeXn4bo088Htlj77/9OvWWYz+INjupIo
3JDoW82bzMcQYG6tthkI2sSunG7d5LfSqCD1TR1/MesJY9ZNzVl60C1U/LZhR3MT
H2K1GHruMpVZlONAwWScI3bg08c8e5VDZfpsyK4YtsvpLNzw6epIi65z4mn9UOT2
QKfzXtR+jGYTL0929me17QUSqd/yNCKjWSus2Ox5268ZEIdvCaz2maYExIwnmhf9
BANX2PlN9p18lQBQzX/adelit2d41MEHR111skOIxyHz4zGAfM+VtID/T+hqkmxV
z3YZKCPCqKUTAw+pK4UPt6Id1hZ5RGhPTrRjcC0kYciQDc3gjJEiB6uIxz75mKsi
M8kgVTvmhsVHtpGEe7voSlCTmoM9sDOI6BAPn20iy0SK4mmMLNQXqQcGPSESRRLQ
+kLiciDHTvCW+o66SETzOcyWGvekhr7SfDf5CpERaPA8Ck3LiTumKjfnpUDNXqN4
QRR1kXcju8bGqtYbMLaldJYJrWdO5whiefSrqCWYtvtGV4/m2t0lFBcJXLlEFzJR
dky9PsXJHzZcy7FFe9phDmYrGrihXtzT2/aoIQxr+/azgZnG+vTWAzEi2+gxBLpS
/RtAryQGge33doxbeukR0QOeXV3j8bFYLW2rqAqnm2IoeyQQOowEVSbzzZBsrPZU
0w7pN+E/vZETTgPE6+DTJfhSgd5wMV2J21Vfbj6LC5+VJpAj98goLldA152xeuFb
5ZwFHnp6KEgjhXdoKMPUDNY7BRbcVouSlI38vuE6grwRLFyR/lna2IWFyKvddXNh
w6EnwRvu6s1Dg4mCNUMPvgAMOOr3d8WCWYs9zNyDXwwbbuAiORWdvY55VUfdeqwP
StifKDOAvnhIpUxtc6DgiP9WGVptvi9doqTxv4+le4FojUDW9x2hmibJSdK/s7jU
EtrEyuU/dPSwTBkOdVQHXfWsQZ1DhVlpXv+lVzCe1hwB0FWo+NmLlK3SyTA+4LCd
8kq8ZXt6bI9IH6NMJrIw6G3tFrs5lvNxVI5pkzlr/1MLdrmmCzfO1DAiy7RayfGb
E6infvSYRib2ZDxNVWkUX81wxCpY9N3Cht9PoUVXtuHl9oBv+5W4nux0WszJ4AJ6
dLg4Nlqt+NrkFgPAfRo0BPL980QhmKGJtZ+lZaeACofG6oepu++4nmnzNugj1q3C
kkjeR5vCje4lpA5ztqoA9NoBw1dqJRKOWB0t6t5TSVYs0NN6kv9mSXoJ3bFcQ3z8
R8Vvn779TRYmJO0eu7iD1R2MNiGNl450QnhloJKOR4gVEFveU9pV4Y62cmUzwiQn
71npMjog1mzltpBhd6VsK5SbamRdQhmjX0n18Zd2+muJKCYJJ09bD3amgSacx1aO
vZsAGPNUtcwxNKT4VeH91z2LMWkEYRojjDqsNkDV47zqYdVQBaug9K4wOEJGuCgs
X9p/uxO5eacWPauJDAk80bmKHp3D8BB6xiuBAH21qvnnr9eIVcFuP5mH3r62xzkK
uiWELnpBOCH7IqPS01b3kWh1yY+4BRUX2KqBe2nagjm4loX7ryznFBEetIiQbhj2
ACxsa2krwTSMaN+KhIls+8ntBqKy7eFOHY1ZrxqZKd1ht8E07lE76VVcK6S7C5ET
LJUT5N/rmzV2YaREP4Bgy9Oj/oSnJlRVuP/VJ2IOaMSbeSn0jDi6BtkPc+BHF4X5
CZFWdDBWc22GZcJUdBMLOdUGAQ//BE9cSeFdMmKJEnzAE2py//6sonYgrNVCkmlc
deBjz0P4WnNdRiG2KGco65ygKJFy4SgWi2NmXwWUfIdVWYkZkkaOgk7rr87BklEZ
xOkuqCjm3E6KAxepKe19doTpJ+21Rv/MzIJPdXs8C+6+87zWVtLYOHsHzodzd+re
Y86FjwtRdfVBH007WUfh44qVCi0Ccua+LwSV6ruNlCUWjJ661NzYsHzVS3xvC9oC
Y0OO1OXisG9P3WpuGrjeqN3BGCNCAmDH+uDHWZW/h7eAzj40CqUlKRrOP80Z8Wpp
A6bjXDBdwO9a2yLlLTE1VqTifPpg2DaVHp6GyfWr64fnOCi50m3wnUUPiTt5jXgb
90+AAVlKKMf0W4iNjs1J1NWL/PF/XT7ES4l/vjX7ustqLGxmbEbRf0iqZDcoWlar
tnih4YAyx8Pm0m1JZCtcjz8268/IX31PoBaEuVAbDBXcKs5MsGQG5RXZ96Cb0E5J
9GwmT66LOeM/k00pNn0kjutxhPSQPyAUpvXfnHGtkAQZyZTR4lzJBdXjxd8VXtX0
GimK+US4Ez5Friho6mad7BK1NYUV389ZC8dV+H+Paazjr7ao22shi+7k9THmJecQ
fVmXfL0YgBtSG6pmlr9iai0UdNjMTAlRoVsKoGDLRANIFM9gLPh1wHQBQIOpMM2L
6dsD8h0WbWXg7WLg4f9K5TpTIRAGZFmuEi8DYhj1RLeiVolAeutNe7+Vc72JbN99
H8Wv2uU0NWcpAWO+VCR9yU212gsZB6yHhtlmZgX86Q19D3Cejq1xub/YlHSeWgb3
u2aqo7lLU9ngYR5Ogn0DpB5a3IZtxoDJ0tihYstiZrOd9KtTxAsZCcP5I64o/83Y
GwVxujv7Bozt9zNqv7W4rvKoJ0dCqMFcFbRmUksnD+h4VrOrqqRvT5fD7HfUFhB7
2IfVbVT9eaH3FZRiUPFMdPh3vdOjHS1D4lrWr9pgBDWalUNYKF9UtcrXlpfs/uNw
8DJynLq6QUgU7uKab9mtCxhMS64M8ZaWILF+gm7BhT9/s5Uu86RPmEdLDI2jFYga
RiQCGdHOB4JfFR0mkudPzwBA58dh9rxsN5oFZMgvrjDZPIRYf2cW+EANMraFC+iK
pEJH9NFqiBrZ0LAjDHghfT7YWL3ZrzihBRxXjSJVqyTPZku55GesVumNOAMplEBX
B/9u615cnm9bvapd3qF6Uzi121qO6TxRLaZ/x74Kuhh17LFX7znm3204T8OiIStm
gyUZM+6BhXsjOoVDEp9iJyEX9k/9F50oEx/MEAyAQ1goluiTxWpUPtfcsQEWA/26
vzZTf8Bvg0q6aM3S1wmMacanzvOdfSuJyeWxonV8fudnjtfaob7pcIzKaTW3QQ+X
5Vv8VQN4ObgGHlnO3NX+u7JQodRrpaBjbVlASVc+R+BgOnoMSd0ogZWsqU4xci0k
Ebimwbwmw0USKNrT+1hKL3nho7eT1XIj+xGPv3eQ7IVPaam+d7aGpwk/Fuhlebj8
ZV9Ndlh2SIxfrJpdyR2jQEMlWqpsLKiXyUoUjHVlLqx9v4NfkjTDfH4QScvmn/Ar
0ROgGuzKWiWGSwXpmAzgIgcFbkP0ZuxWFJXKVZNWc1jTvrMcbbZrVVuIIxMJF9HL
5SpdMCKNw83KaIZ24kLy6REPVkO2eyBIXm3fgVlFLXOYD9evjcs7cDOKJjh/0spr
bpyQTCQBWv775Tv9V041qNXUQwxpmfb2FAWLYlU/u1JjH1hSD+aI9SmhmJJzFPgR
n9QJDspaShLc2zU6XSI+HQ6Vp2ssixmyEpAb8seqxY13TZHx+fr+ihEVc3k+2Bjc
42SI53OVt6okBjvmpmJ7pkusZ2ly3gWFnJj0p5Pfg45tXOCNNdcRg3mBo8/7Usfp
WlP4yLqgy1RnJnr5dvt1co9o4/E3SNdUXFnLVsj0NlYKyQfF39LueEhB1yv9UCAE
kFX+CizfZ3tTijTQeLSFgKcqa2BFI2dZkBBhgLqKyi+7SZY4DtevGxy5N5nNL/k9
IHs6yjkVl57YHQKikVlgYkLagevFiyjOv5dcoQ1AxpCQ6mvYzMQmhNDu3mwOk+YN
hmN+blMrxpHivxTtdql83JsIYiBnaACxiW8FDRO350rFyXljyPpC8oIaHXbMN3/L
f9mNpjJGsRYaBUViWySNrO27rfcL/csoIgfwU28JEEBa1KFdVqYD8DiLuCMGSnKa
U0GpNtdKHaIcvXGFo2vUJKtCYGc9DKgcVkbOAo7iFWKPP5MWjCZWp1HsH1NwfRC/
rVPFKoeX56eQT7N+rzL7wSi9S1YRzn7FOFMncrF3NTxe/KMmRDesAKPrEphQmbJ9
AvIcCMaMyugDlfvftQhVqqGh13pLZ7cpW9ob6q331DQBafzG2gDobwlAPwLe/8tF
DG+NJRZCknFJurwydc5RqAQBxz4c/7a2RuQaQb3yrVVLm3Q1Aj089CORMW9kaZjl
+QcrMLoa3RnXvjtBRHm0dGxetCKSICW1BE3meqfC48TIrEW13JB5e1/TfjwqqA5b
K64ScMuHcZftQ+GKF4GGJOz02nEnzCZTg1TaVQvwJ6r1ymKFOSSYOesopE4MZNZr
+4GMyrY0OKCk2qLbq268uxtTYLcSD8GZ/j2HQW88zNEPHY56zqcrT/cMnuLlxecz
+u5tu5Nw6WukV4TnMWi31UN+ciAb1bwaHSQT0MpMbBbOcfzdQcuKbCp0dA67aug8
CR4fA/pPtnvhuwNuqHUJ5lto/jVpxp48AcYiaTgKArrnvRkrcNsJBK2AWLVvQed4
9IckigLll7ubfD8RbFI65ve1ir2iTfJNmvO+nUkvAJRT+AJwJjZhb55Qk3VeImnf
WBQNibLzcbFB+D+BpENJlf5GZViAG9ItMAfUsLdpyvGXM7BGH+lwEQNk9qwvWiIM
nZ44BMUbGHiji/xzmJ18H2nQVoqsIGAazFrXLNsv3Bl5GXVViGZQHTO8vw+s+8A4
5h/KCHiIAjMHSUhewzyKUI6PZ9GonmMhqUOlkBRy2AvKGeOX7X7BDRcZtqQyW7T+
bLC0nQGc1C2MwSWmrskg7pEBJzxaauNCrXBBs2Z9ojXwGLkG5itI0tqfKDq59J44
RTbH3+BEnyElo0H3ULVzZAVMbFhlREz51wlN61Cqqo1xf2Y4BN0C1YOWwQoqNqv/
IA3T1HB++VP4eIEoc6oXG8u4bMghts83ETLgpU+4ElQhLHqm8sTkS6cMrfZlkvnq
uis6ydI29vsrC/3Timfnp4w3zRENGJo8cRTHh2oOzR1gSrvL6/XV7epV2Xk3OKDd
P2IKT0advX1TI1rjdN/fkquoVc/DEAzWKez1EH92x0i2fH7UQJmZZzqnDMPQ+ElX
peIZjGjGyLYkMrwknKOQFD5dRsdIinGB4oYcUDbObXdA7iSNNbN/IQQUpMIOrSvJ
mrx1PpuhVcDQvDD1A3DgW4ojXvElSdNvvqVGa8HDQmRWEkP2CX3GJnV4HCqz+AFL
TpiTwicE50YSR06jbXPCLThHY8Cl91cXJOnsFjT5uyeteuW5kM1G0B46K+WUYLgl
F/ZRAP/UKlV9BkoAnLp1kbLxxHNoAWeTHj93lEW6Hagf/61j3x1Z4QreB+ipqLBn
mRzOMa3gdiaMkp5i6VtXbUnxku+E5UhvVVM+z8EnqL8xLvYpG6ZyuwsXCC8YiiRc
fMAJssHBpWPxvOT7/1/87poj7LSfcgIyf6YBh+Z54yhsIlnW9qj34Nci/qGIb0Zh
aFxRlpi9Ht6FihULccfocIM0FSknB/5FcwBCjBr8ACDkIt1/8cajy9rl4lt1luPc
EWi4etFDVxfzZ46E+D6oSmpo7MLjG/MDo+L7UWmary144g1RnFaxOIHyPS7hGRyi
D35MR4jO/zgtE/fhci0cQd0VEQ0DfRKHbiwMU+5C/W7nkdHeWkHAp0f7R7BH1iiJ
gXd8LXcfx9i943rgVLyx8LKsp7rBk4H0x3ES61REScm97EIYJ1mZ1VOspMcVd0uQ
DIaMK3fhAUMq8C8kqC2nxns4CTBWukjJBcOmqx+qtO/LkgR7ghy8r9ds0gdwTXLS
R5Z22WuWLlVzykB0Fl9u+g7MgKaGjX3pwkuf+NB57d5fKoOQodZYvJKc1fCcIfN8
begfcfMXtlkh5jHPyOxf1czPRXznlbKrsRwdiRiWh9ThCgewXN6ROG7ff8oE+pZP
RIOi0w5paBgDCb5fnU6QSoRf+a4lVt/ssCpLjRlPWHiFkNFlZpdPwzfQVQKE3eJa
zH1F0rQzp9RT9qRZzIuLKuJq3fHp74BAdJr6vLVNSZZgE/Uelh5ZY5IudLhAiOGK
SI4r/M+wiK57XsGNyy3LImKtPcRKkDAk8wPMdjTMqR/5zIu2+2E+1n8fBSFpwfcb
CohegGPCoYVxIe1q42qthsFEx2EaXlY2GLM1lYNYlE5zXcHSDJSCcgDMAEwh3bIO
tzq6oAL0IeZK4FL7wlcUHbJnq4f7uECIpYOO8eGurEI2XuqENjjcAiL4OvpTrMVy
IG7+T2LcnkUZLqNDYO6e2vsvxzBiIVGFxMs6h2qaWm8t96jRM5YM7tvH0jYOh7Ug
KVOpEm3Od0MaNAS9/yTvzdatDw8OeZP50y0Cr8qAUKB5cro3ahelnRcVf+mnQDG8
6JU0UioNxum6hLH8/xfnsBnoSWXFxi/RqDpBzjBhuZJHqkuyYn83CeS+xuUqxsnn
XQwH2XOLCdkRUwKJolykA1rq98vtj9mH7H1RKGzPon5UXzmYv985HVgazq3znfn/
k/8AzOepZCvQvB/pno4cRhctreQZ5LeCI68oq6OUbHflK02pe1MYDOkT++epKbY9
fZd67Id5JiEeymhrc53xOtwe1Ax1FhNiQuxDMQrt6V1hIGuJeapHa4CytPYVFcMK
qLW5Vnvd+DeJzKd8yPhIUxWeTgiUNf9hYi8HqFTXLGpLil4zXkf4gMlAwbLCl/z9
1OFM5mbNtsTkFePQ0uc4KjnAmq7PHGmUnDshrFwPjoF0AywnjhafDzUV7q23MG6Y
ehTZMpN8JvUb/B7x1tEGRFkth4TxHX+INynY+5WAmOXkZKfRrgHHAPB9VzkaMwcf
2CvWoGy0MSUQbm/SduEDrEcwN5ftfvPQ6SP4mQVjH988+3v/zVBy7B3HM/sWSgpC
lZA3dV7uNm79y9fQTBU3Xk1yDm9iqTt/UEkgZ+tAaeOdHawHjZTiNUMnC5LtaKaj
f1x+g2p4Wn/Gixo9jaJFrdqmbjgA2wkehr2K+7IAPfRIpqQ5T5s3qqjLpneNlMRD
X6K1bzJK3AKXjSKuo1kJJaPcIvLwnkhL0P19cb/vAm91XlTfKlZ6pHnJXhqWbQTb
a04dOQ1AXVBm5pJwhUm3mDtDRBoSVeJoM4jzhPAIFv7+E6CumEGqwz5DMl8XMaD6
4U88PydsmgoMWQdW81zkce+IqDKh2aaqfTzsbAvdmhVmtHLCmGkzGyX57zIvRKwZ
Fvfhw+dv7743v0I/FTTq+HJSWd7CFcJnXwnOn7BFpL0ZPKji+U/awhaEztg33PKt
HJd8j8nNKD/XPUGCDyXHp0id4suDBAXn6GldVwt4mf1sUGxLOcMKID+eM62ZdIw1
L+nE2Ibz69iqiXzfT1OjNx7WLNPIof9i1UIupsU6EEbBUAFcCqzOz3DXvxeesH11
Kd5vT+00KtRoLqLyMVOW23uTtk9PjFSj0aXLUVUrDX9DMGqzoOXmV3OtGFSjbdtN
aoJ8jUE8Sz+I68Ke/H8R4c4L7k2J55f8MShlx+1M/3ajFAlYDf1y1oRqBTm4dYwz
QwUokXuEVG3u2WrecQZpbczqQ5KuuRhi22F4cEq+kTh1klRMRt+MsGBY5hHykFmZ
fCv0wiyFUmXa+QNqDpDQ7Y+h0Ee1qZ6Jpwy0j+z4ePkzDDfe9GKu5v3BBEh8oh3G
pxCVCYhdYri2tkKzwzhkehSRQqTEHTFYTnFfkiW9WXfxGr8ZOE6owsyuWJgvOBny
9WJD//UuR8U0ma22f5V9uvEW3EhbLBe/zohAmcnw4Ow/4CPnUKWcmUJLsBYgCoaj
7t6Md/jOgk/Q1GEjWZm390Latcr14NbeVvkBtU/G8aqbKEoCvFkhvxkwQNav3bIQ
wtoVc3BF6DgmDCC6MXanHJnOY+K6s/uWW9bwAQ99BB3/mLWplny6KCIDjlMVH/DD
aaqhSPtY4aAwhP0cK9p+et7Dzjl0lIVVpQVvFUaGwo1hs+tXhQCxc6Kcmv7sPUbG
cJ034qxdbRBYdTevlXglq5PR0Yh1ZpVakzXFi9PUzUZMXqbw2VRlUcVkjggMJipJ
BWhHhPi18Z8k1LuPLxkI0SVrTUNVUqB7cnDN3Z9kFWRH3nY5yZTT06uG2TZsSfUv
4egLgw4Ny3oBjQNERGfT8WES8MYhmo3QONmtA5b7+ufYqQb2urs2hAfOL9ijqC1W
FOt1INIUpZLwOnO4D9pN7/3OTGgNqyab5tJP/saRap1xxrH7gu7t0ThWZpDP5YgG
JK7VxEGuoaXjAY90ETh6bl2miLVCj+uIPq2aZQzr3EoNGsW5nj2gXJec6elzf3gO
d6fZye0tBL+ZANBc++qtKwhTEqbuK7ev9P3LHjGUgc57XDkxeajd1N0wS33HAAHN
rgJMps8eYdzzl6fMRqAIg5UqQSvmhV5u7VCa8Z1zCJNLtIG4G5eN9X+WSk+05E94
2PVUBNkqsBpz1J+3b1wXxpu4p1+eTngpOiMzHpjDMwYihcKCCXe/F+2YxMdDa97s
gq6ZS8+POFjdmo7PMDwkUASkeqUP2l2YlQvP5Fyvbw+CHNlDqYakHc5oPFWR7g4H
Ew5mKp356SB7cR65z0vLgFYWzUGJIT3cGFb2D1rWl/BeH1Rcpbk0tcHzgyhy/ujU
8kJZC3nKFJYzZVP9eOgFXIadsA6bNV2S83S8sLebrW1uf7Q7EGIknEHqTQmbd96k
WSU+/lB1ZIzpO3VvjLc++/+4ooWPYzwfYgwDuhls0IqRQQeIzNhsBPydAfh53z9m
tIwoGbJZJ6TtA7Jp1SwM7DcxJYCrwh87pPpSRY1ULeHIfD60APuYYnzzwXIDL0wb
idIjzDvm+cM2mQ8R7C1jOHbs67eHEoVqkFin7dTmX+aHdRAPZ40WtywZO3ifFEcU
72GHaGVq2VPEVJlBefPZN07jKFqFnomGAB+KeOCGkNJKufqbL3UWTy1HKJVzMNOZ
wKyA54b0MsSP/mKfoNhIskq2xx3ZpNQwx6ofJGwXidkrqZlNbn249ALS7XikhC3y
LWHtwtQLkY4l1Fymq6eApSxX/N7WqWIgMD64P3Kbwg7Yj+mZcJct2IL6CA6T3QPO
yPKkZA931gp1S11AjjaJDaGBaEptP/U0LfF/eKRnNfjktr0heScCmz3fop6SUEqI
fUfZZwkQ/m3y2nrPqAzB36xBT4PHAixKTbqx15/wiMr6bcfjnVWRmJj5J9vQe38F
pxvWp/oeVBT8/vxO6dMTBc6rgy9mqGcV4Q3H4lqnCHVZKzlSoSBVVYe66VRGrtCh
c/Ki1G/7CBZc6WH4BxrrEOzGg35yDi6X+VbGzY4QBJmeoTBLbZn9Vwvswa+I4Li+
FuTnB2S2fcM0RZRnk8lDaD1QmMZ9cra/YFuK0E0xLjzLj30NO4ck9/ebPF6R9HuH
NHlJQVkRNy2+I5A3MODmCxu4NgTxLx+9baXwBjsvY2B8I44GdEonJ3K9lXkB9L7q
3xw04VKT2DYvRziwRlNJ8g1f+s7RXFSQtcO9PDp63L9RnAfEk1V/xmn9QcMzrC06
D8nKQ9zjQ4gIOYkBQ4EYz9dz/dCJA2RnFsGlcoUMfCsn6Pu6DYedSA/Itof91kLr
z0gnUiQQrrhmnJ/CmCu0z+EHuzqupXfNDsL9bFjpMNQOGfjh9LSyTNWybHMamU/4
bR92SU24EoPydszpgwb/aUWlmIBYnnBM+r7zO4Eemc/sAXCTW9eN0grHoPKsgAb9
8CMz9xU11j9lBwVRXXu3UDVz17mnlof39hC33AoIaypxRa7ximhxbyPIrSCtnS7P
yadBaC45CyxMCyQliMhvf1no2D8tBXQiEy2x4gxj/ynfU+9JH28GPSy+Q3i8qaF+
Kiet6Q0HYm5eiSPliiuUPy53rZVFymw1oxVnKOhknIGrqGWPHdc4gJrXyKhsL1bq
fThTDAZ9jB5dVkEemxGaeQHp/bOkjwmuAXzwwC2yTeFwZfCxbuPUTlhQLe5acmU7
LMGHT7R6TRBds/G8mdFBWq9toVEPwjPT0quw0UmDntdjlXOLF2LAeJjfS00pjhdR
rmuVZYayz8aFtKw89++VjxIAsiEmQ6qZIgGLlzlODlUnwvJIJr6QPtkmSf88Du+3
F7JoHXt/pQaLf4INSR4WcXCwT1hjy0wmS2SD3arTWGmz1Mh75cWDbQMcbjKKkS4G
qJfGBdSql3jI2ewo65r9+l32AZX8GgLQ9G9We9mGYOhC8GvgRkcNxhtOVpm57L4K
OWfAdDIkslBMMZonFfCb2a4EA5M/i5cbLLn7emZEzJfzXb1sZRBrQXAsWdNYtmJP
hD1iqjxT598o9QCWLrYGx5rVBpMduUSEDjgBh1T0Uk4yEyqQMAr+r/ytd477dh1X
oL+mc5WbX2TCsrgjTwOsRtdf1jLQm1fl7YkJsVXTXJMJVE9dtiFLtsx58gGWutpG
0uhtYQoSeexudacYyUrWoW5ZvVVwKHPfNTEzvn4YrSnyWOmus2apd1sqnsmZ74ea
wD8jIL1ZscStRifjcNSTkqgMX9J8xKWBKwuQ4tePIxzmV97yEaFveyVxlXkAxIGE
hxvIfmdrPYAxOoe1yLuzfEO2cWYMStYhULMdEV5wb52xcRD/h+XbkfukEt8wWtp7
EuiUNgF8C5D+Okylpo8n1/ElEmN8LpALttxKOcF3SUS2CWb/EFu5O3o0cVl9NjOR
Ly0SmxgL5ofgOQwltp/k5wBmfXukRYAKyDBbyJ2S/72gric9+ylOZI9dYIrLHiNY
EKBuRF6Fvr5NAumz0/dtocDn853K+FS78NSo5Iqnbzwc/EDbhLhp98+zobZI89dy
brAPUJAFjeG3x3Xv/pP4kUL7wTwmJB9BbZtvewUx9hp2GppYOJGRYTEXl0pD8ztF
5fdVbGWiGp++rJ09wX3Q2FykMafPkpx+G14RyPTrLmzluACA5r9XBXD0NRujD7G8
Qdr2WQfniOgKFK58oUFsN2nGBqCuGiA3KLy6X6s3tAqSEq2kEMZmEb8I02GsGt8d
z3b0uD14GAAF10duxMQqmp7GS4rOhOTt/FOKVzyZv1opO0+yNO2wFWL8eTFl/8ma
S4CB+7BwIwrMxg2BiVJQyAHwqN9/TFr4Kp91jHh++fNYYuQzcFoFQKYChk0Bx1yD
DYhqor1H/H7uXxB1N2zx3ib1AZAbAouNfXnnFrEYN+Cn+ztYypUJf2LiaNu6xvYV
I6BbozlTtY/k4SEiBzon05QCVyU0/XuAgsqHsOTxKPJR9+6nQQJazjLR81uPBr5m
wOBwia/dazpAvsuVYzV2U9+56TeQaaMhVsZ3EP5ZFuMyRm2RcoqpycTNeHrMPOED
TquWHj8owPjKJXIAK/3Ke5O5XETyM4CV18+kqKKbxKlgoVap2dVfiRsQ4x2NfIqm
Y7Y6L9qey27deDCNusnxDtbxfNLkFM/elfO7TceLI333cRxzyABWGCRjyPwO4x8u
Q4Hcw4OHEjx708c1sg678L6Apf8ZdW9A/4U2dzBnMcR9vfx41zz9nQWq+Sx86emi
V8K+yB8qtpzIZJzRQHJnL0Tnc5uXR2QjfIK60JL27+t3MCk5zaHgQeMsd6bDwZd1
kS5iLkGaQmLdMr/ufOG6F7bgtWgFsaVK1WBbY//qOsc+fEpopgbcWFexVP9emRTG
ihiM/300YEojEnuaGRLMxnbo3o/sY+f7KwFMOlCKu2XyraBp0PpmklOTzEjk4Ej1
mkO5Fb/wmvY/PTaq4tuxGaSRt0e5G+/UpH4qHTTKLRPnV9Pd5E9jmxqzdxthIJYn
q+oTd7KlbFPkwqdDVgffYiLGSzFjynnHy/9KzBtpyGD2lBoqLCQCaBwljQ/hozOh
t8NES1i0SX8/UROz5UjUsKIMJKR7XEtZ/GJQmprCed6Ml0ZcF89dTJtCjlySuAHp
TMJH4XAQ95FbERDwFCxw0Fi1GOYJKHmON8KKDc/2SuZOlen7fJfwqN8At+3tdBx/
AafxUUY4uHAuvS3l25W1PRAAqqmgMjort51kCGngiAEjiJ5Z9CwQJxUSEgj1AQZ8
j7Spsh8VjG/90OsFvq8cXt0BwTUoT6zh3c1Hn5zQpkRjU+9r5ojYT5D/KAMSSU55
knXNoXPyG9guTC0IAtaPaJBGKfREIJSTHVzC8u33KHFrMvLzlHjRTjXUWYenYXQq
t71EoTkniXRDlNPDBZ2iPc+avqyDedXq6IcPRVb31+9o8B4iGM7YEAlNSJR/YUu2
1eTof55Mf4kkS6MbZ07n90ywdlSPVjqQXmxEzIZAA7gLAgyyWrJt+yY2lEfeaCzN
AvWCj+c/AIu+7yArUeAiqJppAXiGaprEuvam4W6LuSRznvIJzXzF13tKjk3GUisr
Sb/zhggqzmJosaS9T3+Q51wFiqfNYgGLxMwyAE4bafCypYs3GDfaH4n6id8DzFQW
rSdhtJvuEH87RLlAKLGHGhN4LzujXXRv/u4tsf5dO50OpImKtfUcRNdy1LppSjHX
uyvl4PwdiwbxsjlwIizYZlfDiDoSGcVN4zF2Xoo0X91pL/WLOgjMrlaCO2xktEi7
59vqw7WsO/GeGvzqxalKyPwxT26NTvZCrJwD8KchgpM7va+pCV7C6eNzAcOwvF6J
09Jj/3BLS9SzGIovAgRAyGHcAH13+emGn3y4BnrAouVENrTy120PP03qdz7ZAg6a
C42/Cs36WOa0p4WH9uw5GkrWVsx6W+0P/yBol+sRQOls9sXOKr9mSgSdECnC1467
6iu1yLKohouxfBH3/48uXLzFSfLDnPQWupezlROQXA7/Yfrc8iSy11BGj4xwTLU8
3d3W0Ckh+082/Vyk6m3cbi75MYNIwhc4FZbDL9ePT6TzO6l9Yr2em9DHkBFIcSEO
TwwuN5TlsARy/bvi9O6JBhB1Y1EkH7PGaV85peVF7eJ/5c9uaNva77xBn+ZtUD1h
rXVeH3ZCDjplZmWhD8PJVDxs3lU4zrsxXU9FnjCqlziNIoYxsf5SquAgehAOwFjI
EnDxPsoMD1aOFQ7fsn2Afl1qjrTFrnk7oOKutJ3b7MjHfxfWCar3zATisYP8UPBz
ga3xt17nU/E9Gsw4AzsN4oIFoGgcFoWgVDVuKRwwrYYstZz7+0RxI9Tgl6nen319
ANWdccN32dtYNq8VqwxzevUWM3ap4WgLxx6FIwD9/8W0ZMI0ql96AvgzZ0b+gjzC
rp1C2Vi7I3wkrQwJhc/9d4vjgjX5sO2ylA9f2nVfYP3l8dTtdS2/5SRCZMGibHHr
BUl70TueWo7FrYecqLazjMu++uIjCY8VNj/xZz+Ad7C2BMI6HMaoAy+2P/oXiQmw
VIYbRJ9tqa+JBQHr+jDknY8zWPtakBzLbOnFqYDfOu6uND4C+nKSFkVRnW3Sfgf5
yH+fWuTLEv/vyoQKZwMFr0TU1R5vY/2jpO4zE9ww8QIWSiV5qcB/HYoV5iqZBUFs
vPy0CD/8f0Sv56JXjsjIxEwzEj+kOdCJjlI/Cr0CUXu5u9xF6ftlR/s/HSh83mzc
s+NLDd2TW/yYtLCdzPgmt6Kd7NR3F4dRrdGHNSGUkQa8ikrAYK8/p/+uvjB6agJ1
pvY8jlXH7KYLFTMXeukA1IhsxQWD6DsRhVrgDXSuLlqlqkANdsrCGIWUXY78Fija
gZ09vhLTnI5oSzKkEB0Ox9MqGmiu5OiZ2CIQnSzLgvYZfNCPWhRLuwPDNfzW+T1M
smHwg5sZfacm2yZem33hR2nz5TQCY99w1oVoUZYcUubWHsAl/B/SL5Ni+f5tHyD9
WEW5tKw6e9kVQARb2AiE7r5/GWrS1RKUMIfsM/DfrDPSM4bEBllw02csgynWRjgk
m5322KCvthL5CLzDUuTYbcBJ//7GqdYplU3BevtdQ3HjpUOyCmfU0kr/01EaBOZZ
yZB8GjqXwLJxQ9GjovNZbP6FCHEAXk7fMNjInr8vhJV077Ogau/tz24KijAh8VOC
4e3/WrFp7j8bp8XqK1iWnRvM0VO3hqH6y8ilTInLIjlc9MSy+lrorCgv9N3mqMOE
saKMXg+aOryRQAawY/GagoqpJWlm6qRkaqhoenrhRZpgKIUblp2oAQubtY02fp5l
/0LUgjNJRq7Q95cWDK21CxO+rosXUUFeAbqMomF81WrPJq6HoxQKOQZ53mgxNE3S
XcdJd12COL5iEWvxgbO9k0xwxD5cZsmdhJ9inNbVHvhmHjTtiPk7IUmfryV2n2dZ
sFFNwheGBwkFccq7GCw7UvZtxCURSH4YByhLDHTNbtyOeDdyGuNGbVXgUFdUf4Qo
s8oi90hqSbB1uIrqI8iYP1yjiRD/YK0VvXn6Cn+GT5/DmUOevRlRAIpM1AMbAmL+
csHgESQ3oj2P1OZJnuxeO/cbAa1MvZjORrrOh7CuQRdI4G9ef+yz5w2H8JysdWXe
CAXKMwaUMiCdtYpFh004ObiQffHSIlbDlyvRWqIOle6XTDu4orQv4ENj7+DP6rcJ
dPlSMpZylnn64Htb2X1nx9l7zJrmJOx8GZmQvcrNk6tWMSSbhJHjAkw4jpYCshMv
GqLfFTyBZRfktcTgNy1IDd/uoWxsvSPxxc0wJve0fiWPd4wt46X/zCBOSiq0gT1K
ln4CS3RGRIRfJdeneeFX29IAzFwSqeNO57suRcHyBYRCD2hI5adhHsWX1giuwG0G
1QvI+PLtt6eiONzzkD7Wk0YJuJbF+JGiVGJDl26vWmx0fEnL4uhcS2u0oV258lCV
w3LN3yOhT+T0vVXTbja3nMgbXv5L1RFA28o+teqyP3T61oxalaxYibIA8VyKld7s
HLjFmg2QJ5dpJ6b5Z4uuWAvpUPEN6pz0GkyAkcUrM9LEgJeKqAkqBgiqF0mWcsqV
0jIk7JHNvpSGXGHOifUa/EXB1027zT8zjcb5aNe5waNps0/IDRExH878gNsC1rfO
RykqoAmWNYkcPoalemeLv5rea/VBknBcbV8OoD9T56yWAsiP2FQoC3CkuWdzuLda
nQs42iDjv4rsUlkN2JSwvEFQQhM0+AtLi5kgs9OfFVHcFOC8BLRoLpUZXeoMM8aP
NTlQVgfKfzzq+ZXvL0Dm+UyH5ssHHFoRi4PgXQYYL+IFDluBaZ8kKfLw45w7evpe
SZ4rAacHo062/odaLmfr6nBMZuytT6/87A1zVpfd7Wv63h1BcrGqO8Aie9tcIdrR
Zhk7d+gz/rQ/KY1MLyw9qlfTdHk6x0NVHaRBP2mQm33sXiVbPgoKTZX+YWPq3Lvm
AwZ21mt1AsBmic7vNxiJeq1VPvEzZHExKoQQdBAu1vPeVjqV/qeHmcKBVXfsIorb
Dc2FzmT67HWZveNDtA1wuPbHzbUvwOb+339+0GDu6G1OoKBBwIkXCUU8ZAWhxo2M
uE4eXIpbJ7XP0/zVF32wSjuPkm0xmNgqg0XZ7i0qjkO336i5Nz0JMe+fsoRgWgD7
JJDupls72VYUziSlnuPobyf7WShtIWkirrqEFn4+LvQWKth8k/RNqbtZ3PFPRK5Z
RJoXNSt4JUnJLN//nMCYh9kAvQrv4oW5H62y3x7qq5PZRqhuggsU+iJD2pb5OATF
OolKtP5+xnxGH3rSZTmm0PMfyqrLxmf0iOm4x+xfjxtQSa69NrlDquxltfozsp2G
1gD5PCt22UeLdpmKM9CB3HwpjEVPsZJXXTFAcvOU3scDB8DuUllVDsJcYHf+AM4I
4RvvIGIqUY3eKYIuPCzp8fHkfcfbkEg3zDi5Ud5jBxBJ4ci3aWvephMmLBBL6oNq
yNKw3K9T1CgCWuMCR5MbavpbFdn6alLP3GbDFLnazg/58KblTZH4vHTUT4HJe/ay
4pt3Mkd0xITvw7DrRNZtHTUhDoJWjXJ8xc01bp4g/igXgvRfmMftRmry8j58Z852
Q3c2qJpV8pwHN7awrMJDzKvKWDIo8TFzzjrjZz8zjwUEIPZHKsCQdmt0WB2SOCNx
QexMJvsAHiVbOkLmEEIeuGy1/IjKKYRFziTJ301RetOcLHgkjzI/e2H+/Es7R5B0
WiLOyy2b6JXNXguxHk20ztbAzI6LE95pC0wjqRwjoCiRkM9SPUFe5WtKqsi462jA
c/unVzfbZjY3PiAfAVmrY8PgSowcwBpWLMGt2TVPZZ+8m0teZWiAEv2YI4Lymdef
MOGLuoeBE17Cn3tZHkmYeh60DDvOR4b24yvddtTNukxIwiCN3yl4M86x7anomsBq
3TIZP6aIOPYSMFvbA8FdmfxnihGvSPwEothrgnK9KzP9RdDArOnRxei0Z3HUqVCl
lfRqDbTLNi7XV4JHIxOdZwKwjgG5Q1bl2ilaBcZH+1ASe7KVRvLwjRV6FnMoTRbg
pIA4cIQqAlOB31tILSrY3yZjWDEGhosfddA2Y7ecJ4QpIKrYXg2+ssjw4HHDAmF9
ukBf58Qc+hV3PjC2JMAv3BXgfarxuF3juwrwMj7dOKh9LIuOn1j7KNgDf4seeYUa
uXFWE7UHTGO1HwWhAHZrLI/eMbc1hJIAkpktQxWBg1UGHMyCeiENCK4QFh7eMNFv
BBWonjB8JbUK0HkrwPdI8pltdntRpzqBk9FmdBRQnPG4+bFdiojH+/Nm1kJlmP5P
mpMf/yi3HljK+aj4KGiBCTq3QRaMd10yd8/uUv2amaj5Ke/SpqcLUBRkVwE3E14Z
1sSbRI5VclkylcSBIj8K97RllTuxF4eeJCGNuPPsVmBFJL2Co16ALKx32tKmpqEN
RmDMNo+rVPJTK7+Jzdp+uBqqPwLi+junpRMXZ5xw9OuQT5bKZOtSmiMOU7v0aErL
MOALBGwrZrquwhMtr2hoMtZIRtAqd6a8UadSzLgKI4q5x4Jj6MJTZlJncPuf+Qrx
UNSmNC/1jdiv3+HA2TeplJ+Ha4dWdYXKC91Jkm0J2bjbl16OBnTjG+UF1mP3Qo93
61OBTjG9c+QoeS4x6EZCTARHN0oNDmklaEHxwnlEo1v1EswfUGYW5GCUhfnsyDvO
gXCtZDIM9ms9nHgD4pTOm/pmJbruBX4Mukwk1viePvyr7xhkiDOhtxnPngklgezB
Sy8gWcR4yTKdwvxdPoIotil2oaFKIXMfrG96Lj/f+2vNyZzp3YGB3QGozoyUZMkE
faR//fcUr3DIRXLMnAmKp+FRy6XurxPqFRTBUS5cNyJo2hnzxtfx0RcPzHI+FyuP
qbfUGgpuqbsbJUjsPuT4cZb8dnbOcbJw6rUK0d7ZWIdFpHXvGlLKBB0X0rqmRNOA
MNexIYnnlyBqzRkmMaCi8Ot0lmOYIurPdy0n1+vEgbmjcW2E5vcCHxKKomaEnKho
joZmWbw98k0DTlZiXhMer4CdARQwbwTTXis3eoC4WUjO1YayvsJEb9YTkTmfm4/D
4JFtK85+tfOsfJ7reBwS+z1K+1GIrTdk4P2vYn2kDdVd1kke+riery+R1EcIXJVW
g3th6C2qqup7FgDVezK2xHDmQbEIQERvJTCPsKaR1TBmvP94ZxGLHQp36hc/bZ9p
VHUuz+jymPeLprmIfiaBBgXGW6GRbfEfG0lhDG1uEye5Tr3VMmJ1qh4ScSBVnhCX
D+80oFvbmDMHgOCEGex47HKOixG3tU/TYmFOE/TPBm5DFiVNQpZSOzmPRLvjrBBo
ecM0SvC9sVyyFOCt7OzP9tSCqrFC8U3WiVR74AmO8qhwlZVjlPRJGKOTeiii/VDK
fkfGZwbgsLRg10rGXlWFRvpWVyxM77JVPsR5/5tJNd8/3Zl0DuzIPpCY9WT7baC2
y+ptylxPRF7JjX/XneinAZjW2m6e9vdqOSK0NLrBZmjpfbC0vx8FsjKxzojR4wwR
OIQfP8AL+EBVMZt1IrZ4fKMTbNBXUnqwr1f9JIUSxuxH9xG41Y3RSiz/d/2qI7To
Leuf1x4f/VaFjvXDNy/ZLQHz5PGiKqfq13tZI+zPkqY2EdxALN3qFGXKZmRx3u3c
BkcJelNoS86FylQ1gcpiprIgMHoJ84Gt+3o78cmdzVzVNwKuVWG4c+3/FDxLaMJs
1egzfCtQladWTNxJSSOCWAtW0f0nqRt4J7cd5kq+OABUHfoRiU5VF8Gi/+g85uad
eJG2BfdpfaDwm4WjoXRlTmE1PDF/N1QyteyrQ5Z6mi+hkG97pV3vhj9W7jGxIdU6
kPT2Vx7xYh7amxX2Kx2U9pYiwCjhbK4ywp9ij7OkdqRU5mHF2evzZe9UAOXWL6IM
89GGR03tT9pT3ZkbBmzxhhf8pniyyL4r4OkBlYnZIUPOdm7SmJtaris37hiQOwtD
arvU7qGVyy1N2HW613JYe9q8isg5qgYMr4glt6VolewkH7yYxBRFzcy7QEWF7oSM
g3Obt6fYbnrQlOzmnKXgRz8ljUCXdku7lumlVNP4OrcjIYuhfF+mRxvXQKKfEPAa
VOU2b3v40fQNQJCZbLKxaxOgrtonQulJw1aeiFdeCdNXRfEYlAnJzwn97n9jNgS2
YaljKki17yoIkTHz3Yh+ulcNN0dgPh+hF+USBzyGh/d6HtmfsJEb2ecllFwDmxtt
DBEMpq7EKQ6BqVsird7FDlJYWJsgK91cwKmDj0Nc7L3ivj9wtRCgI2mCbqgZByfs
x522O3mlWMRGFsoW2TP1s/zQW814RMmdin5IgbZmaeBXGgyqxdXTvMOedXBtBjDT
clcIdzdy4kP6BapXPp8I7fDkgI6ZZS9tSKCjfPERv6HVjPwmx3KcNZkUS2AzSFXp
QTUrUNUUm8kr4/dhPmzOo8LBBW7MIOSSO6TjsB1ZX4iCOHjd+hUEvSPNwiuhZtRT
k055NVfN7Lu+fNFppZdlDAxeZww3Erk6L9di2NAJsU6LGPVDAwUdBbx53KMH+s4x
KxTtbbGgkXquxKJv/QxM91ihr536aROc5qik1EiQ3dh02hypVvNXxCCjHqzF63Xi
b1R44DBpcm10KGMLclImCwVGppwEINOn/MYIQ+xwP9JpK8qToVEMbW+Ww8PwPwGp
6sZddsRRdToqKjYlqR63+DMM/TSx7WUux8kyP9dkKDvm4PFSBHTZ+Elj99eSNdav
/dwGvR9JdzzIwtODLNYVvpKRcBIE3MkzOoG8L84HTTbmqXIpmgiXNJ8fZGgMJ/5z
7shi7V5fdnk1jDIaNjZNb4cnTROn6aHin+4D51aTk+mWXDE/TjaXU0jkm/WZIfwc
XrZK/sxGZp+CCbrLFpbCMc5ILQBxzgRTwCf8E5emQyPr27F7FLMTpf2L61hMk9wM
CeYWEw+XaFhrM3V6HbXhy/Yivct1tiqL1s/mRNLHQjZO0XepLZufpZHodxQy4dQo
JeMaFF2Jfa6p+Zg0zY1BcJwMUONANrignugq5uLbx+gIGPaxSsaCr8jad6QWyoEj
2XL9JRlWKIk0zvux1XaXt3rCQ+w0TLX8lkojRxbUkRcdVBDe2Tbsd8cduvNUpbp9
jECffF0EW7VsxKQLVEaUXnhQ2GOTbiaOTaRScYlYr/9BJ8dL+FExi9EMZAeOeCCK
Ce/COkR/2TFabwuoYhpo8rJiMxrB4sb9ILoNgPG0ZCpQyqubkn7ibUds1yqmGPEc
5PDZYzhXi+Hs5yZRb3EUj1N6Q8WMuNzuCPb7jetjeeFFk36o5Gvh/xnADNfwlZUx
WEbUsTj2rUWk9uSCfSMrUkGRjMIiq6HwBsmVhRCmy617cByNTl8a3KC798t6jQ3l
9VC9O1CpLtH8b97f95Z11eQEGufl3dmfPfC/YpPPt021Su4LbYBf5h9sjWX+Ge8R
ME7t4U3hOPi9wZ8qsRTTGzKH1t7mJc0uAzWR/Wibnq0gFvLrRZw0dsX6/UDx44t6
htiwDfq81GZzBQj0/90PYU35flgs/JwrP0FZRZQX7LOGNbAMB9cxMAC6ELTkx3GE
Eq6MERuqfbcJQRLBvTFGR3dUBwgkJrdeNYqx7yUmV1Pfn/ogG2cZXJm7SskYVGia
J9ue1iNlPdMPRO4Ujr8UvL4vQZF0vfImZCZvTT/aQxrijD0YIZqlMUVSK9Xhqb5L
q3VQz++XobJwddfIkzttMQkQP4zzMUZ8wlAD7GsFPW25yx8RC4FXL41IcCiIgtS5
ojUNCvimeo5FuSm1Q7l13tHCsp3W/qFxbsdz9YoTkdsM9iYNNygswHUXdQlRiXe4
gKUNHIEXRrXNnp1yU6niLKrj8wWlp7P1R6ka7Ak2K/c1q4NTRTp0d5YH6gRxQljC
oB7QjTni36PU+D8/CkSbJgu5VJIvsQIlfZ75CTseQHbZieXlw8THeULDnmgfGLDC
smamhKj5aRqEyUP4MeEC6ipbpZCfh8PyxIziWzrTH6m+a9eKtwnorh1dHtGiYxOR
JDB5GYCPiO7DADlgEEw6awsDQjoWJ6m6xut1eEdD/+n8eikLi7iuDAq01/0NXIzE
QB77icFMgzhIsJL2xeV9B0Fc+iNnwk3DTK241TkDxCz+NH86LQoX2SJJdPiPp9z4
U15Xds3vAOnzLZ4L9bvfoa+26VMnhD8SeQEjjsSUNIpI2WgETf8rUO4S6m0vN4rC
vh771BJtfpclQi97htbaF0gzDdK1zBT0NtzraoJl1tCYzJchhEc1J18BZ+JWnFl1
N1vVsoIyCMEvQRg573JwQl91iKaEZXZAdY8f2kMnTp4NJXuzSe6RMSvsIaTXiGQr
UyPabcGxHhHFij8uWpOfc4+dCKAWonPy9Yv42nrwQVKGpnJGLVwQ34lq0AScg02/
Vr158aW/1ivWFfxIFPWPf3ElvIbRRFW0JED0Zqz3l8qyhteLG9Hxq+Ll6RoO/IUB
xBdGPRKm/ozKi9PRFDnNzaXQYDqNJO8+7bhaXjNlgqKD6tQrupbwxB9z0Uzr2WwI
XCIpM+RMkylLF+ALpccCIHhaH+Wda5XXdGcPDJoYWpVaVa1nUzeLlSLNksAaGTNz
Hwy19lW5iS+kmC9YFO0AVwKkNkgR0FYJWwRbwhcYZxYVD1dUvGFN+AOynMJVBDlT
hxfQtGTpB4E8peqeTjUtOsWHmK1UHFu6HlR/I/m3FjTtSBimU7Jc7vL1XLjAdcZg
Qeqq0iut1aEyoM3RJKBvdkdwtoA5Nz6UUR6UqnItPIrUozfVEI+8HWzWZZuldIQv
bE7EUnyEO62t7lFqIdbgJx0eHSwJAhJYUxtuH93Hj97bwV2z3l3xIs8c9eGDw9B7
KkOTvDOvUeNThvytl8HS2JWTUibuQO+q8IEpHG6MM8w6LwBv1Nl3jHUNRYrK2N2c
w0TejVap+StcUMO9KLurN4cUxqj+nA6t7y5rL9VxDKDPTE4ezmv/L/s7ps8P3IAC
UhaaLG3A4NQUN6TvIH+H4CTEqF+a/BukjkdPJ8Veka3DP6GmHBq4hYoUXAwAFz7f
UmJC8ywcaKRLJ6LUPMC52sa2KFVlLrPYPzx2o+4KLIrXzTvUhGw4kn6ryBdbmZE+
u98wC0TJghwQRwzogX6Hkx+dxmZYZJuWhnrQ9Ym2Cc40OgCG0qQGrBYTrSC6wL65
KR8DcGjfW3DhTUNFFDtJ72TXw/RkobaxAhgHSX5HVbSI5VeR9xLjXfZKqmhV1YUE
n8prhWB1XwFnadlJXfY8AOGHK9TllFF+v2cOJ/eDWFBunucIm2dx9hd23gc+vMiR
OT50xnK89L85EXTjOJvoil5p5fnX2S1HvCuV4zlN8DjJ3U51t62K7GtdjnJOCwTR
RiS82sSBzl7zlVpNs5CI7ldAwHrAONrQHC+zeJ3e0yBd/SAFzyMjjkNDBpFAeDU5
0JGA9sYNxbh0lTjflujxGFFJd3Z8ZPcW+BGhVnSoyu8GpAnBbh0Dpg6LMte/mX0W
ra27okWAgwqkfS1W9p5eRMvmwT/nQnBgZT9+oCduis9Sa9V5AnSCQu8F7o7gwYn1
tJcQNzs0709K3R18/PK3dbTDmvA5CEHvNYWtpmCaRhvKk9z6r8t/bA+ouM1X17lA
zbSDOAR8BDgVLm4fGEqXQY9wEyAhXMFOI/d+ustKRvQg51Za3RWfDIAEVVQIduUT
It8S4dM5nH4mcKMffDpOLewYxBhh71C6mjutNSiM7wIGGW49PN4N8fUwHTxMDoD4
RerBn/uf+Isx1yXzVbmGvSgUtyX8tYaCydx3MBkewRuahj4HIC8wB25+W4yU97Ri
Os3L6hoBKLcCtLZvJPjeouYJUChIp/6K7NshamlpJPalZZOjGEBLnSQ6ZHxsJkgo
qM+PKqV4FUjrG0Nc50t2ftY1DvADFTODp2lGmNALINGi867VT8SIuOz8XzatNXpX
XoS/mtl26d1qfHGxhQQq5sWrrsTUdFa0yt4ZnCrSupOJExJanEln7s7nfAG99SDg
l0HdXR+UYLi3HFg0nQq2GSp0NUgdCjtqiwVkSASRNLs78eN/JLS+mEnSDNxGUyVg
BT5U6RrRaDqxYRWD7HavszDddKXZkrBZk2p1CTuPRhvTWJRiumFYOJLpqmzvQHQ1
26Byiy5Q0ht4WIOpCfl36tS9UuMgvdh4gEdItCyThf6LSas1IPHHXb7OxkilyBMw
/GPjSa0VjmQK/qwOyWxZzcbC02AuFF0iIllbcD46H5HdIfDeCuN0k046ayifCG5y
0Bwta/1ja740fGVPc8AW7+C6U2OGc3cGt5NFfG2F1lN6Ct7lBwCW+xyqM30C46ES
e3U0XBw2KH5QFe0C7Wmt7UCTKmlhyzCYFCy1H+6FtMarl4AgT6W7LntQI4VmLgS3
u1IzyhCJoX4T79mKrWYu9lVPFxm4/jQ6uyePcjezfmDDvD7REX0vkXJ1fvh6CtM4
dLCQPc0xICJ3BhdIe5/Tx40V2oE4Xieh1gDL2+BuOtik5bqgbGX3DoEDMXxVLnt9
Xp9xY/69cPse/NWMH7rI1RnyYktgO/Cn/IhhrO3t995UpEnez/s4uVF/YhGG4pR9
P5230O7fSzyauzF+ZZjb9KyZgLVrn6/5jLJKuCpSO2dnSmB0i+XlXqB9CrJu9vlf
UJLAoEWQVnjE6l+VpYl+1mWZWEwGHvFaDwi/1gZXlXw7d5qjlQmtgg1+QM3zBP9F
8nW3szIbbcW94nniq/POaX5EsbAWvrZWZ9hKXhPR38eMk7fcei1T2rAGPrgk5v1U
ZMgo7rbQ3qXivxRNddMo6krv16h3k/jjL5vSN/6LiS90wmQSgDVE0TidKTATmrmk
wbKGb9p08sykgrh/R87yh99xHU1U1Qo72K1rUpI/gCSxjhVakFXLA3P3rxfUcXhw
YL9D65j6hfSdG28fQYk76rE2yPwel78NZPNY8yhOlzgJmeqw04h4M/JxD6HXBk6C
eB8gwL1kjOjNRb10a2A23LakQlMaeUXL8SnunA4onidhRGClMn/HpOiQe4ABu654
Gku4v647ssA6zoxvRl0O/NXelw5iMfI1GKWK2czLoWigba3jb/bApGtE/6bS6f+a
fOw/zogFJAzvZfaP5hTyDsioftkUhqAQEvttRYwcS9El6AMMj4nUxx0oUJ7lCp5C
SqmXnO1w2/fiHv265zb+o10h6C4/3RogKU66n2KnIgmjT0WJ31euAwcy20CtQApW
lJ5aSSH5ZZv3q/kTn+f6nQDgrp129kCMKHLLftPecUfQy8pEBKzRk0vfWFAZFhGP
x0J9SHGnpmrPCMNj3LVqOZzDEyjVBv4ruFkYVWBgPIucDzSQSRlXkBj6KrFW8EBq
SDUhdi5RFZu5XO8qfSf6sDIgktHflDTGrs4DjbwdQ8Lo5geXNo/2Lo0IFFgaDeS/
aLswBlASukhs+Dp/J4zUPbaYleL+38xpGYgZDLUwkKa+zWxHpbpvSaLhwGVMPAnZ
TonoaKmUo88zvg65RZIyKYCtdJzqZzyGUauy3IJLGYkGr8Xt7zQ2zWYA++tmIc97
xSwZgxDIufe3x7ipBBGIhhpay4CzGJgDIkGc3wUSVcp1Xjsfums1AtH/tpEKGY1T
l+x0uxzRpvCViyqORy8CAruG0h7BwWOW0mrqjmoCuoLl3YvsCbflNIAx6kooraFR
gJYl7gD7dpJmENnoPjTHQN1Xe/bFV2FeEc40cmfhE/T6/6uLcHZUwLVglJ56Y9lx
L2DTyb99mxot6hy+Zth06UaHA8r0wkCty3G3fz/YiRYfJQExjgDUWNSj4sdyNsf7
x7VS1j/E7XEf/4ALhinqvF1mhBLdcw3DgDj37fc4knDxFdENxzvruWtG+sbhttke
dGAO/sTVAZ5amB0joTZuP3I86dIlK/bBN66mH5q3eugg9X3/u6gqk2Qxt5ivm0xg
6UKRr9aPwerCpfJemxw1qxStbLF9E4C6vIy0YGhNNwZAa0LR7Wr8dGnJI/dSorxB
QSsVbtgB1NtM7rDMO6MaKNRfhXp+8p6xA4LbBdvA51L0qhEu7Gu2cum30fgV3EoQ
sH9r/0H+yi6l2uEitWI24OQ9Yom+oWtPp28BNpzfeBIxjzeSRMnIoiggHuekdeZR
W5OqXZousRVMC2ObfOTZVydYMHxUIlEQSfqOT4QQVfobQ1ZzZrupHZaTxGqVJxs6
Zgsp60s4lANqFxK0fOQRUjdCiE1WlBfvI8+8OKkqfV5BWEM0iF7pgZ2Mvx8JImrG
GiZE9p8Rz8pZTLl8PNRlgCi4Wg5JPgE32A6pAiVc0+pJrRIb286E5UCm1cx3Bkky
SQCTyAmQGj+klZLIV3p57CQN5kZMvKER3885Budp/V3yTJlhVpkkgCQD+0uEy0D9
h7ldxGB06Ppgjc1EZr1jZ3aaZy4N3U2hsdDsqzQP0ydADk11KcTROxfbIDEDDv+d
RRSqvd+OVQ4zSEil0xpZTqX/fsWPMoeGMTIf8nhIot7Pdq+1gqU4sU01snesw22h
ZmM9pBz3i//uVnP4bYyZGbdUmBV5vrHRDrtLuMYevEBkVr+/kEoEEdTPE7j2u6XK
uOYD5Zq9TLq9R3xz+ydFVgRpyxgv3Kc7CUJ+R3hD4cbEwg1UnmVSl8d0LqsTsGwW
1Oo6A4Gzoq95aivkt2RjN0e171lXqT9nrjCqrM79rwBu+hvZnnP6jsALPhbPaMuD
JEC8X0lfTIi7cQwkfGm9Dd+1ijEqZOoQ1ZSv9BMC8O50llQ6dSxpwJPul7r3s6Qq
W6AtiR2r0X/4IYRqXKKFRMcOOB78LjW6RNA3ZvTume4E1PbqLz/QiEPTy7DgKfOz
2rNJbSbWsmwVdCoQ0KaVIuRvtbvDgHr3/BRfr0h9GsmQMSYSbsvt6zoREkgjELyu
QsEWGPx+1/IxHiEfcYFWshrAEPbsh911T94sDuUpqyXD+A10VnN6+J28P834zE03
LPvzVV91MBrlcXAUfomOjggdwd15xg7WVLbQ9bS/2y3gfG3aO3qhAh502QQmsAvo
k/sB3ddmmwTZaqpv3Ms1lb5F4d1RFbCuvGIFm9CwqAvugKsMqTfwaYS1eBKvMneV
1LEXQiCatVmRpjU12vpn1cc7iC3oZwhYj6aRsg6xXSgVp+hHnaBGoBLEG5lkh/wL
nLHzsRnM+UWfJHO1wR4lfkpanQtsncPBh9fp7hGJCWXqghHo+DzM7B8EbVWh3h7A
oboSmRMUPkLCkaLR12VAte+Sv6TZTiyP06XKTH4nJrTYHaQ7TmDtWX4PitYQaM4/
1kFOqQRKNM1ddrVVUSaY3mQ+s4+tqN1d8stGLFr70ZK3Ou3YY/ODooOq+bq7s7U+
SsC9xp0luejAVNVLiZfC4Z82CEwT+b+jGkfPsmumpMZhUhPw4Qjjteqe2NjFpPPG
l2P/5nB/b+7xPOJ7FxhFx1IHrg8VBBQZAd6Q4QgfLwq1ml3vqJs229sUdWQqs1pY
D820Vl6KLNZCLukKd7XhS8TdLi0OEY4Q0NZQdQCyHnj3BuRZ7cdsPKZjNNTpU4S0
EoAXiHE752qUIpYl8+XmeN4rtpxgAIz61OI/rGzePugX1Lx5hWVYMva0U6Ar/TWh
UbyrxCxojQolWT1uYVGmosTM6jsnKtNW11pfVIXGsCh09VioFDlm25Z9w/SUzbhY
8VR636trfBrFA4YWy96iu/pCOryOxCp6XTRRRwZXBxLWUAobWwoK2SmXOXO2OqfH
+IrE6jPdcc96DgKsbMzC/DlcZKWGsw/Dm/Hc60By6PGcRFNfO/M1ZMfEIggHZPPf
q3ghiDkpkX3io06caJiNuyr5VO02HyEctqg0DY6EfgdrUwffCCx3LIsT5NYN/cb/
bUNefq8cc0U2RwPX32ANmSZRcMTcnmwlJDz7ssDOi8LC8Z2IzD4FxUcC3WdbVk30
PbLeW6RrdVJQj9Pgs4WhaRLnAzRc7MUz+KBBL+6gPQrfiZAxMerZ/NqtgW072tZU
XwtDhFpMbTnS2fdJH3v+gx0TsZes1AOE3kxT6YGOh/A0zVx4fIAKTgSGl/YMDTrH
iQd196CtgoX5V9Izye80KQXb66riNUUCJLXjlwS5nb8y42+YxcTydBAtxZbJAys0
aZU/zCgHQzw2z7QyhknD3LZj6eX61EGZeVO+tuwNBuLWq4QItCkOJvnxTafboym+
h+JW0DzyqYO8JxU7X2f2+s2oQMw0FBm08N7b+CeGAAdH+c+CHtwFN8JORG3aHEL4
qyfHccXv8OGvizgtdn9Olxa22DXDibnV6Ehgs6BX89CKgtfgl3jKWTAzkGMW+Q7+
U2Axz+fGh5m+UB6nRpYitxndnLxpf9tsm2WEOmbm3zM2PQP2BEvkn3DiXoc9BSwt
0TQR6FuzFSchp1rXbGdlEk19hdH9jccVRYYZlq1xj5jSfAGFUYRfMJa0UVti5Jnq
uP+0yYGKzy2GBtTsyTBKthR/5pKhl6Q1oBYzSy0411SpuKGAgoV5J2iBO/bGfgNx
b4hBygtKSJ5aevZGy24UX9KoNIxrZozXBLiY5SgwjH6sUjpYXvAdGbOLI8HrV/Kk
DEv5VjoV81UeeSWZAk4d5I8yvBdn31RoYbdO1X4eYQQj4d4hRB54ZXU81Qxt+a8E
+60VqpBzyBKIXjXDfy+hYqMOHm2U+bym6rcigOlL31Uh0/xxS2z2sgiuEHZsvP/Q
7NI0aPc1aJPhbdJM5a1/GdGHCOOPVcW4gylSAkQk75nRsqRlB7kj8o3rK1WjcHv8
X9u8r2P1sLfJ2Ln1zZ10LFM/YZAJTCU4sJTYoWeQ4rtUc4NQfRBL+jRZg6cu0Fjz
7qaYTyjkt2M0nc1sk3dNKguyfN/4Ma0jmJFtCoDS6B2Etwb6M2J2hEyqmj5vthpv
rgnrEyfCUe+GcXga4pnyTAIDQwJuBLSfpO6a8xm1a5G/ixcHri1Se0li26X3ie9/
95dEcn62LPhGnZqTJlqdfyWrNtMrogwJcHEfbyQXrH67r2J+R+QF4MPvulU/lk2F
hpGRZ1T8R5srHiSBDUYtAz3CwJXsDIttq1jQEpANAI1d78Hv0sg8KBCPdRmR3xzP
cqMFyPIxAZrMhkwQw40mhGDPbD4C3ojIy4Jjnh1Zz0Vu5cwN587qqdgVc1E564j1
oZckzduNxj51OmB0mV1X2AqhBWOt0CDrhoZiNjRO3yA3WSMoSG1aPxw2jhIqlenS
AbzZKpc1f3sITXkHx+NNMp6FszNxHJbIGBTrHdePepuXdkn+2W6XunrVo5i6tuSw
rc2YK4oBc/asCUyuBY12DHPE3gGtTYMY8+VcLgPFZgm5lvf0SX/KonHlBSyZ2q+N
sES9tDY9Fcd31t+ybJAMKNZdkDidh1PPYVF6enYcp0fksyZn+7gBS/bhzD8DjQS0
Mi3OU5xdMKZCXH0eoGysr59+FRc0rL0d18x6d76S/n+Tn8A7AG+7cAScVO9rk0gb
nfj2LkhmIoy/QrInaiNJw8nHgAKmNR3ph9FhlMHshSCP3EFZfOBzKnBejnAvvLe2
yOSHV8ed1guDl07cKXt0c0puPDgpQQdvJcZDk4zGdUP1Gs3Xdv7FRU7wTZzTxAzY
AjnX4M6/yL6PcuhpTRwQHoJLYtj9EcZx9n5xC+sPeYYkNQjVV/VGTD4zLKe8+Bxe
eZNj2WoV3wUZFssDijhW32LgJ4afiPQ6d44433OXU53FZ7+HDQ48YrqlP/AVMraY
iT/X71GcjaE8rm2qXCLkYyYTI2KBscX2S90+/bpWUKK4YrqtMiZh8Z75qLwcLG4Q
JXFfASBxZdoXrlJSuUW0SPdObtKnhUvMF0pbVIIsrI8i0MhLUZVy1nqDmslxs6V9
3k4QBViGXMp4WCk/Kwd4vmK+5Iv56QiPJSfjuCimFl+EU6iulzGsmEM77YHSSNM0
sWuy0det/iygXKQ6T+OkBCaTAIexRoo2V5CSifybehiuEn3r3vQYG4/fJrEpn1sH
ZcaN5rASjWAzmMvT2JVjNwe483iVs3X9BN8hHtDsZMZuIq66FErCMB/+jgOBNVFg
qqrV50UhVA4JPsIrVprh7J46HfSdIsIkx+PoiTQ1M1VhLhLgWYcjD3OPr5VxXloc
0D+lfV/MDY1PwPz3lkMaEx3El7fdFsUeM0m+pUOQe30vRDqx/xpXs9GlZ4LzERN4
GR/uYOaa5pAilR4aR+bm+4nwthJNzaLIysZouz+sqDg34zEu1sWiQffV8HzDBnT2
FQmpU5aIfNTBAcW3hJvab2qhIYjiPNx6AAqVDRkdERd82gE1FqutJRN25Gev5l5t
Qtn7Ry96VG4xNPBbDbvikuzYAEKtHElGzYAM0271hl9eWYj/C2NKJ4IPCIRPntQY
OGe6u5k5YHLrOkLJQvBi8svq+QnWZixjIGknX3ouCS3kIsvSBCDJKCFL4uGBXqRg
DW+iBlK2mxIRW8caSptzDY7FS0N2BEIClJbYRDIh8sBl1TLjYC0vZIMwtjQEAfXy
H9cfmxOFKExDWIZbEF1G1/uEruXuqwVjTxQtFdc+4b2iX5dTHRwr+L1MnolSmsrr
v9Nm2AANCKXgm2ujYdszvG7bKXRopfJCCUtJFNcvYfQvGCEd/1SOZI238boqPD0J
K9CJDtscIdmjUvbH9fM7Z8eChq8J8yj1Sr4twtGfpwauqOUP8B3/gLutELJ9/QXp
2Pgwb9KDZuDaVdPvXFgQh+jUTcIfzOyOspsUEA4sMeFWh1+Dnn3W9oH2J84yejZn
Z43Ji3RBZ9j2L20+jmrJDreQ0zYxMcVkh/+cbd6qewQoyugEpTqn3K/sGrfOhGWB
onT8ffGC4oD9XmvX4N2c8elnh6xrR+1YTfC7nmLLSIt5vectMxy+q8JyUO3bIb8N
PIlkqUxg4mXlgJBsqwpzlkOCS03zAHG51wQMxPIKucRt+YXwdN1MhHiaZP4QtQlZ
IB0NrSPPY7ZU3OV32CrsQLAuRhcy82+lcp3CHzy11WOzbf9bqaQU/967RBBLJqSB
Tk+HDMLSR4AgcRYZaheQsJUHsvs4t74h3QmYpEtRTwHNIH34xJXYo0TWmHHOO1PF
meRzoiOPCEoVOkvCIYbwuhQ/D7x3jUzMSTVSodsFtaA+sAOJwKswCpuVBkk3UtQH
yxjsrGzxSV2LagJ2ijh1fIyQUsj46Z2OFwVKYUgoz+qXj5GdI61wiMBXbAJB6lI1
zePJ86m/4MwRSD70E83ydjMlxOBYpnu1nbyIdnG1RrpSIdF/TmLFlHlasz97GAfz
c9Ed/u/dcnKyPbrUZESEAqPdcB0O5aB1ehy+pPs+6SGKQ4WQS72VCNVbP2RXW6sD
Q41kAyJLWvJ8w9e2kGMjzT3CuV30J/Id/67tplVOy8pzNfAQ5Erw4/4S6Po6fO+E
J7qnPRe5hU1oN6HEd7WoIY1l+UHu2R3/FX9hZ9MC237kFAOBtSxK7kIdKRxCBl9m
eLZ9qA7GE1uknM9e0vlKnYsNxoPsAVjQu8Z2EEUxyfa+IRbK7zJtNA9wrFIjFaNq
clBIPl4xaOGHsflNFOdjtOn9aYRf2LHVyrw9WMhhj6AULCRkSiesIF14vOlY4mJq
2AK0CFvmCrJY+7LD1gD/SwflmE/mlYqLVjSJlryOaMTk27iGziOrpgF65cxhaLmK
xGbPqOVWr734qIRhjPAWQwScIfWPzzQHlfsoCceMCCo17WJYHQqioM/TZptXyuN6
JxAwUOoNv0WRmhMEAolJDqphSn14RtusSnw1mAlGdz24m20Kbid+YKwV2+31lnh/
mHbOt79RNRBXtdecuPP58ITI0bAFbPs2qoM05xHCGFp6XHmI24GsOvz1tz1SfJUt
scldTM79fudIV3Cx/tgfYjKIZNKY7Xd5gkX6Z1wlMurynxFQgXPFHTF7/0znluqv
cSZA36qSiYhhdk3GNO+udRYl73pI0lZaabj+H7botpatk3aY7S3jO3xrso+Z6m+S
nNtbLTJB9cWcdJa+4w8l+4bPj4rrjhEyqKZb9YpvokTTP6cZwZ2WUEzDPJcEFF66
RjTKE2gL6f/5uwniHu8q1PfvQTk53Xv3n9nmoxYt551kFA08/A2fSP1pahsemxbE
FW+zk0BdoRLVemYrJbnMXVJCmiqddNROjrpw11UKfxLxGXNOfr15vaB55eYyAhFH
AhVmVm61JuK7S+FvyHyTvcDla23Qc7x5/t/CKC55ZQuad66GcGd1jAwrRlk35En9
S+aY3LJNR1UoqfYum9ceewbLskYekTsVoZyhcV47UfiCWyxlMUO1gYh/U58cBCS1
Wa2+DzAlCOkxLVbZmGC75JWLOgS6hQiRc5uWxIgUypyQAwvrIGlVLt+rdhkz82fq
RtcloFvLRHrockC7HKmXnz8IlCV/VB+fKmojzT2kJ11OdLlpuKfKjfRcRY8lkMal
2CIDNEgJkcC1G9qvokA5vXH7cBP2zAeCJ4lke0JTZHGn99pLQId9fQ3RrLgSOHy4
htDdbDOon0doauP8lyxP/TBLdu7vbzwuFPWZwm1oggVjE3ynx2t2B+qno/nUleI9
Sh/OpA6uCa8+Ry0U9B+DyG3c5OTLTjlhjyvvax+m516BxwKpNbwHYM5wV6Jh2Nom
NfS7vmm8bTWOHIB4n1V53mgOO5NNgty9ZPr5bD2Ix+5RdjyYluX0x4/RrDQPiexZ
yyvIsVJxfGRmFH7yca+jX5WvFdls5aVFg0FZqtf42lw5Z4FGnJMGUPVhF0IfwA9y
cwj3FoIoq82XExU4oRB2kbGMhHzlzCw2aCF9dS4oj8eQjF0fG+9hzmliZG9pe37B
Puu9GHs+5335DjijAjLM6uvpoqXSzl9QQuZ+qz9BI3R7lub8LRFx+6SbNkf92egj
mJxnRQR7a3Pm8hnDjjvQIpxJK0KXwHZskBIEwHDOzJJ7tiMhmO4Cr7ZUZ3D8NOVP
Vf4rLfIyVEgJRm6Yf1X724Oi3A1rof9HWbd9Jt906Lo4rXuuCdsf+n21rvpJSpml
suLK5P0j5ufrJFRATBl4hfBLnSknzHVOPtRnZzypMQgA7EnG01KQGQ1OyuNkutHi
KZMYnTjAFE9nB+6DdRufpWIarBKj/txvR+FJYJZvSRcYlCxRHDaFKQMfU3OJv3uY
seT1MgBhx1EYlByvHA0qB2L4ftblgScZ42Ar5xmNVt9Y9dFaf3c6ALkeUQDbxPHw
GY08gTfRw3WVplTTVllDfyqlCK7MmQdkI9fgzJWT/egmd1PljlobMP2xQ7IzRbLz
67OYhvRg5ycyNN53i19In0idrMPx4b9JsvSXkDDqsfDRdsRh9PVfrVZWUE+UFRRx
rouk4BXU5OGhOBGaR4dshYk6U3/teR8crNxmWt8DbJ2bzCbjbf3DUKda0IIEtutx
MvuHc+X3PSVim48TuGrfojjT4l3IvJrbQnDs4lxPC0wJeGFkfZ/wYyNCJ0eK+bCE
e6t3mOXJ7tmiDPDNr7BEekQXjE8Cxje96HUsiDlxHt9Vv6lplnWNGMCkIO8jC+dy
HTlUx+i23KGlHeqVPZY9DSyO1Ff+AL4OulVIKXS1P9aI0gLsWWSbsR+hunQLVROm
As0tSQv9SCS0vMBKmr3gxpvenpCLPDJkt703un+epLod9QaSc3lKiXVmfbzLTf9e
YSrFzWLCOs57RBQOnoYjS5nki2XXp+bosv3EP2A2xfhPx9ESCdF9/Ei1ls5viC+G
1RqRcYT+p+8Ba/91+g1cFHX9bd1NrVFNlFz2eNpadAqhcsUuXqVOAizQa/5+fAAN
eFgNW3SgRalVXqFTySQWGlrxkAoR2LjAGzKA2MsfM08BB3y6WxKta/E/75GG++Z1
aVe5lXNHXn/RPwWPs/MXG/LwnOfCsDHrY9/tzAcL2M5AA+KSzFOSm3NKo8w7MfWK
ERzAAK8muQnVrpNWNqAyOiSHDza1ASVoshIo/QTBDp57cNo/xjWs5TleZAEZ2w0o
s8IywHEIQTdUrefTIc/W0WFIyNdAj6zAfs5K8UA2olauA8e0obK0eBJmJb3HcsES
m1sreTe60hOEK4VBxpYwt06IWKns1AzazQtDSon+lt12TdHWzj/EztkZq/zrLgCH
V7MFe/km+m+10gogO3J1+GPLYnPz3n+S2KUMQ4Vsi8UtbwGpbjBjvT7xL1bqdYXR
Fnre5VIZkIx+9GI6rpDiHYJyPzmca4JokuqH/o+BAz+3hw/l5XaD6rPwzGKRgGh0
AyfhWk4s4vrZwXyOCYHsOWan7zVDD89ou/q2473lx+gDtWut670OJHtAA7LWg5Hr
TiJFoD4pTnoTe6Z3fIhDyh/Sy3CDVqx/8EDcs0TMzCG0dkekpoTUNMU5GARZIeHF
erw01vnJw3KrMn+BO58dzgRgcHmVRxI0+0Cac6kL6yH/kHveVgyeYlddMjL6iMkf
NRIAPpSB/YvVSQE2f3sUpLGbMIv0SCd6e5+i7PdOCIcrKoz90j68yOHyqNu1Lz7m
Oh36bjS32/HAuvtmmYCLtTHbbWv6RYVAqSQGPbPyQ9K/KKpgsI3LVtXZJI/1QFdr
N3qp/AMbj6EHHRoAuNRwiuBO+PPk7lJjHnU42KY3BCy0+wdLrGRcd7yRpGFR6/WC
cIrPsp9nTUXjgMqwl4/jPBlBn0PEQmi4fyr2d6Om2/lpuvjrJoU7yorpcR/eXHqA
DD9IuBld7NBUTqSvLA+O4IUzWLurhD/ZIKrjwRzmLTnXCA/eyeX7VeS7HW4WbRb9
tQt57fd6mkJ2Y/yshfbDnPvCOKwxjvR74U/xVE3gCTrnfG8/MQBnAtPtUOTsumPV
b2r+PSHC8bU/ohkB+NzixIclb+5zvjoTlsoWRg1IG9rqrxTNKB7aJhflY6wEWsGI
zsDZSmDEFvJ/FlQRLTv21lfYrHKPPGMRF2TcSoHYgfj5LjXGxFmzfc3rCaHMSZ/z
QA3G0wdw5gxe/MDGwqm6nJYGyO18e1ZL4SFYlLfk/R/wXSSKt+ZQNPG7+Kq50I+N
8Y7F564jnxJBEq0ITLtG2L/N3ADHHes5Y2/FsTphnLUfXIp0f1M1MO2CO6xcZKBa
BTn/WruFSj4MR2N3rncqbzS95+CANn2UbOkURUQutEPtvaGhB9tB2YsGkUJPBoj1
Rz44rB4t6gLJuG4PIHVG6Iw6AQMEKotFm0c8uiIXOjs+dQn5p48gOqHLd3Thgm6v
hNt1PBLKoS11lW+O8cU5yeTadTR6jwa2UAKy5DzPqjD3FpbuUQ6HAL/2axRtABLH
BNIVT/Zo86a0JeGGlHhOJBjqfuvkEc4uUxxQQYyVVezkBE24h6cWJMgTlwTA0/ax
IqdflqryDH4lgHlASL3Ooyhvr1d1Drn+Z/Lxm9RFQoHgLKgTIkMmyLSzhX6XlSyn
xsBsTL9YDPst81pHZbIFHf7M++XvGZyrvXeK3+c8pA1NAdH91qu39dyEbOZ1nyPo
Jo0U/f7ih4Tv3leaC3N6l/svQ8Rk2wDOErnQNZHUI5ix+T4Ars2/BHKCcEPlvlpc
vs8V/vh/+6RPBluM6W3v53B+MX1iwdJVNcbccDYL2uLEXecEs/RphRCc2yUKknic
f4zuuvatyIKiidm4nAjUE/yEkbyg8aErCckG6dfyQyqU9wn1CXv7qnTVgmQfASuJ
wjpB0NXSBpxqMbYDHqnfBte+6lwQsaQu3pZnHufj7ySfJYzabEzuUTRJ8oAPge9G
tA7TyguJtcepNYY/7uXp9RByTAdq2EGzTdMweLYrmd1SNnrnTESB7AhEV74GcMNC
Kxf0a9jx2HzwDCZt6xJ3FZ30JVlMOXBmp9a6Zee3m98GrthjPKpoXZ3+mmjfMlLH
VUxyy3axrKo/jfEpEOJCWVI++NmH9xS60OKtWKS1UWr0LeuCek97Ma4v7gJ5nWRT
uGGgGkHQG/gFSGRdbG5Tr7voGwBDXyUn6UmhV/AjY0IrUuwNfjoSSohPsAYZVTbZ
u/lNBK+ttw8FfLPMJBX6Nje3bZtBueLASXkSc+nEdB594DoYtfuJ6Rm9WxVH2dx9
cS3i1b9H1Q0DSedZpTRLc9txFGR889CYKXJWAQ2Fvs9B9+uaRHu6zAw3EyeV2mcz
SENhnF6D1WkUwYYxAn49zcbeKAxnwi69ng5Njpya8CiyY3ar9xsCWiJuG2svyDVg
yz5nWO8g450AhvLwYtJZWRB3T/A0B8KT6Jiu5ebp1sq7B37nu7sR8JVSaarOTUfP
srR9d15OgRdzSQp2bzsBOIJLSDaqHIT+LQZW4b8czXno8oK0WmHnAyJl05+Kmxtl
7YGBIQMKuyMFmzifxrX2JzLIjUU5LQ2OztlXZ0HUb/XQs9EmU7A9MW8u5Voc82gc
9w+B6AvQUxymH9DQPjFcnyuV4wcF8DbbKCq04tfzdyBlL9VQup1PCNU2DM3ZWlHk
Hi7lYfpyZiC2CDY2/vkE50QfVwgrNwi14WhGFwSZ5rW4Os2QSfBP/F2dCeHgGPXE
AfTwfJeVMjOp//oqWpMZuWsBHlA8i1BxfrqTh9JSiXRIKfyltXAGMA175S5HnWj3
SQzeHuy5yp9ruVE8fxLOhONmr1Pj3Izh4U6EW3Pj5iSNEdE5tnLSX6ZNZtlcNNE+
bPWzVfUKqexMe1w4nALrjCLbRoymY81y/pabfI6B2WqNnGWtyW+9cguWFYeThvy8
n/BqkWsziC8Q+CDLpSLiCKA0oxTmxt76yQYlY2BWqqDDS3hZu9OxBlIv6WjRK0TW
zFly2SQe5/dViWZPeCkxVUFd+OBEzkQ9dHIgB+vnCYy4qV3p+DMuDZA/x0rrPOGc
aCy5HNI7p6KZbqfcLV8LgHd2ZIfQaExHRUiJ04to3yXr8Ic9kxWOYUqPlSyl5V8G
6EdqAKmjyXT4NDKkYfNPN4Fx/qYUAHHepg/oOUlQrpl0VuIyFXhaERx8aU+jCErY
r7A5oQwdTkh+0u6DkLnxPuQ/RlwhEdcsr/SqPMX45krNoqQDVY2PXj4jd1QJk6se
tb4aq1AWnzyMeRtF3T0IKpEoS6SMEGbptaDUBousnI0u7Qzqzv98zrOugnSjjfV2
m6brGonUwScizuSEIL/F1wGUp+War7ni5R19tHLuEMUSnxG7VhQmWvWGUubjTVzm
+dj+0MPMXtlVeDlho/9bNQyeit4B/upRwJGF6xERbCXHywjMbN5d6zbinvf1Pbx5
dedstiu5Kb0LHULTfPYT5M4gWuNIs7NKs3BmGdXrM+n74G5jh0i7xOvf9hSy4SnW
T/QXOr9NMmCnj3RihzdJvut5LgU+laZCjisHt09Pi9nzJAnuGtthKCKOrXhjI6E1
ZuJKzaNJCprDXjfEiAk/uAMnTG616bdDaUhXk4Qp+Xyuro2OATZr/+ylrVqaFm4W
MxHmU8A8332O7X9psi+7vRlVGMhd/wDd6dfLiLMxh6UbyyOIdjo/EdKvnBU2XdEf
9nhHi9/oa8G9vUm35YCLEHfZepSGCO8dubj+5R5hWilGV19mYweRDACChX7Y6T9s
Nng8BZPM7BOf5Co399p8JqLNepmfBWn/dvYFhzJKQ/ndb5NykV4iw3zZgxP50WFn
BQ9pBikT8HPcdAKjQaKc2NiZwlgLn3A/aCoUH0X70ZSX8gflXkiv+zfqqrjBrpyE
zeTdBfqf9X93ROm2Tico0udVvN+jLU/MH7cwp8iMY1BujDcS06jXsvR8a7260Udk
NpaSJwSJBGQDmOs2x/+SSkYgURiEb7+yAOqlzgBBejeDX5gHl9d3o7VCmmK03Dkv
NrUxLvU+fDAyr7/JLgnfiFK816ajo/b2ZZVBRJn46NUIhLhDLseI6Jk51puSfIBz
YaFOc5+D8NHY1tABrym1uHB2mCmleqoaKYAWNQra8wdCCRnUDu38eHiz46MmSCWw
2T9xSfr8Zu4xjUy1Ts1l7+6YrfQ8CSrPnmRWbgL/pUx+W/Yf7J2tEKAkzuHAVKtD
PB3Odhm0AReoy6UjMF9ckppULBcvIaAhjdBVJsrhS911rE6NyGZNCsARhu32D7Q9
KUhVaXQYNN/919HoJSLmymJDbYgCReuFNJ1mwYkgen+embe6xJjXA+6iVwrzsp5m
5Vug2pWDmOmn1HLXvNgt37mm15vQqcAuf/+7JFepqiTRLeKJ/MGvi4YjxjOUKmvp
yrU3a9uarH3yeDWcbOWvoRwOZM5KAXJTl0YbudAzbtvRf4C9alVPEGPkGcS9P/KB
I96NSijz2OiKdvMFPsSMeP381I1JoEQMlZDVYN8fV75Y8AupRteBmOS9xIqgUkI9
3AprrDa28Kbuce0TpthNV7+7tA1Galw6f7g4yfxGg2mO4yUwSgvVMC48EAivoYtP
kWj942cet/Sb/nrgE+5J4nypBDPLn2rhnk0YhSxPvdRTn9y+MWde9wFG42LZHw/m
JhUtmMCxia77Q/ZHCWJSC9qg4EGThkp2rgc2BMpcvv4yW2+UjkUtiti6evvmyjgN
mcN5XDfgwSlGAeW34qTWI+iiqDePxEHwF47lx4SespFkrY8saJhWgZ8Yj2jNZEg4
NWEpIIpd2gUeTbYDucbCYT5owSf2023JrfZdfdtv9xSoujjOol3vWysCNStosyAk
PDZ2oib6bhyAip/9aqgiHw+rnC8k5SHmXvpuAwpiEXdXZf+gyBtHscSZZ6ke8mHM
QD6BT2/aO31pY5AHXgoSYMxW9eiSjgZUJD/X2cwqf85njwi7z9qyHRARRgEH0zT8
xtL3b/ug1A3kVDYB926AycTnLqSyCri7m+LY7XRo5fWd1z00zw88opqT3jomuDAh
wbT0fd6WPzRqlwR3lTGedFY4kX9Uz0EY0N8QcAQA0iJwJJnwAkuO6+RW5oTSqYbx
JcsieNI2SFl/0meOIk1b5s1AnCH8mZQHO24h80eZt/UDrbYGWPqzWXrie58VQQhk
UzTmh/IHEv62Xve21cyKwSE6m1YamH7ec57JECgOZ1DpV+RoNbqHVkxN/t8kcxRK
CtZmlXvLaMRQHMetiIsPpvKvph1aE6ergt2ZG7VHvsKpoErnQ02YmstBaiJ8EhZ5
b5F/lN67hNSShaAUmrUNZvBSf71rhiBtdo03sHGDrFnmuenzWl0wz3nRmrBQ8Ot5
2gNM4QjUJ4v6DYEUzAN+mEEbrKBQuiDFbOXsS7si/J9RfEZQqqWMPH4Sr/8fkI9e
Yjpnzu9++hM0ZgSfIMk0Y7vyUB25Bo3LQV78D2YHHK03m5zts3EvTXd9FnhSWjiQ
EgMWq8AeCKmeaFS8eguBZx7HkLWUFu+JQjZA9xFaiMB8n+iNs34+NH3xPXLUS/Xk
tvVNhQRvxXN9sC9dTIeXXPHUhLAzlWGCK2Zi8v7HW1n3qV8eynFPVTYvhtbbHk0c
TLz4XbNIfbFSpR5aopqCaDGrKnZv8xHMTxicA0kTPSMJSYppeyvehftsip6YzRy7
ImrS6/nScAbmQaBkMGqx36tGiHKRiRzcGjwRNVycPjYjJsY+f10WUQKhIa6VDr8r
t9yCRzkY1+3GfyejgEMP2MDlxRb+Hq9R9ppxuyOGRXLIfQhgXieBC+J10U9+mtvT
47cYpyapblCXSsdNjqDLQhX6Y64IFBi7Ud0u427k8hIQ8PvOZuDe049fAOOTpjyB
tQ4Worr2lNA7aRhLimylN57/e6T7bM+b/wxbka1eeznX5DC6iwfuTAJgXi433keW
SiQvMSvgwW5WOjom0HNB2vmgpQyKq0TEwBoBInxqD/SjzYNVyf01ohIi3QhfRzk7
+AKMoUDB+uxjt2oSaFyGxmsKyG56s3H7CNURQMpnij+7cwzYGNA0zswkdgoerCZ4
RHMth5h7YyAsH4U3iL3JKfYLvacCVowZzSuQ4gGbv8hYPRXMZyxsuJVUG+lTa/Tw
v6P56C8CN3ON+oPmFSB6E2l3XU4gm81HBDc9sr776/TQjydSHoRC73I8KzIq1X8M
Er5vbf0PTzM6yUd7+EfsC9WT07c4kAX/LHOFDAlXLE+q5fHPBzp9oV43tbDWggDa
+JEDo0t1yUv75X6hu9RcEq/V1wpwcJW/njUP29YfP26QWY7mShlCVOLCgOdxA4O6
tAACl1/az35Gsvrje6gxGnZQIWEnSGvd03RTd1qpAnBAHmoCWStiseDqlnAikl9Z
b4M6u3moCYKCJd9TaTreHU5t6+GvWHUxVvv1v4ZPE8ODSUeNznDyfHxVIpW8OGIR
kNo0NRSg9yT+bhdkbActBy1TIc8fAf2D03d33CxG40Uwty9eGw3vAUXxUjgzCTxx
GWnb7joJOz7S2rwoqdkOKifGe0wLFMkkxneFoti6za6/f4HzeEiEwzWFPZHH8qlb
dKNTO7Vjo6Q6CCSuyT1Shzb6s1fSVL9GtzkOq9iDRMFvr22I/Qqv7lfjnqPwD9UM
HV9LKtxwdQA4NW9t6k3cGrrgM7yac5ueOOMdtjFH1msuw/bbiEDgUG+ApKnXrKZW
lrxbW01PO6jPqGuUCEIuWjDyKgmqIHHxxgFG1YM/4JiE48pJmp+ww4mKpHMRLOT2
oE50EOXF+FeRVB4FdyZHFz+8hqKO7Jc43F8AR4nL+5YOfanDXYI7Rx3avTJNd3MQ
R1A60jgU38Mkl8Ens63trv26jEtE490cdzv4A8PY27L0qb+IziGOBj17g3eyOA4X
TaFiAzFVk6DO6Svj2Iv6WuWLZvDQHquulIi62YPy2cHwbVFtSh8gz3w/zbWsC18G
i8SoMvbK0WQAQPSS/IxrUQKZvEeT/kWkTmGnRdY8J1NzQgHytfSNG+/tGXbfY+2+
+yygqRBfV4mndSLHrrwpSqUDQwqjURYuWaOqQINYEUlhClvqO8wuCqqMkZMwxDMb
utHWNY6UW51nqRgtLENzlsIGyKLFOIJo8Vqup6ltxZER6x8FF2yzO85+ZiNYzNpj
gKQBk96MCtBW9i3LfrBR63ShvJpt+rdulQkhwMpjoUWafnsfpxrguepnclK6oliN
+oApc+UwXoY7tNOO3BIlLMyHw6DJPH1i6xyXUlzY7WgCjeQ3+ESlt2qLVEW3h3kz
Dlpa45KPg2n8S+2vKkGzUxGqHMkPC78jbJDsh0OWv4L2uEAvleIK4BW8KxAzHURn
3XLpdUXx6ywq09KuLaTXETrrPS1YZXKdzATFuLItd99+dt1ncy3MdU6yLXHaNljb
CEsZcvS5F5ZJAOkZNLNzJFeDLMNEMm2iQRzQO9AJvwlonkTAOJvRl+WNZQvmpQzR
aaD+3I3Zq1hSUW5cv90M2mb+OD57O1RtNFRiOR3cwkWjXG4cG+Dc8zGcjrqFzGvP
KYCFINh38uZL4GfKou/Gb2pdPsOshdL5pvdiwnyWu/goN0HeVeu5SWmYR0bp+FSu
KPutXLVmYLZpgDzyuMRE0/N/OHKxC+VS51fKshVGpBZSCnlzoM4e8eHfbgPLnF29
4tgp3tFSBbAEflbYce7K8EY5wILYuK1SdoPnoqp9jQMmVHruC0vNhU9XJ2MHhamz
+cC0taOyERDvy0waTmINpRA7nXc3Xll8HILFAiWxvHsC9+gcklrW+jl0B0EQm17G
GAIkq/EftzSfayrII8fC9G4PTjXAZ/lO8wT5mz6l63GG3s8lXdNDiAbJObtV1lgP
+BgrB86Muti2mWW4ET8XJjm8dHrZFaa7zAw+SH4ijkuRtgCB19LDYiFYHwKnDSzx
Bsb+lRuop7vjCRgTv629q+fI2MzakWPg25c0cuEz4+hEh7s/MACyJs2R0YuFHvuz
2WiRoDIBdQ0ZDlZ+nlm6exBIczgPlBVKTaD9ca6dFhjKBZ2wvLzQGTGkzw2eit7M
AhlZPvxpw0uGva0VfSWqouvUBjObcEWzGYQCCdYivNT7udrdsJEa84K/zL2QIMUK
aIOZdf/zKSCLGshJ0cAPtnVva+ApWq+Ggehofje8mECUKKAxKrcfIjyYkWClfOc+
cEzS76BBRbf3epE3t/RPnchB6pJ+SXKvAa4pNAlNlwggvU0UUe8+Q6AX9/2MTKp0
ycyZIQO/CUFfPHJMFtXL5FtCqAmGm0SuoydGXtub7b3QYlyjshAeL3ThxDPs+tLJ
EBe/wV3ZS+haLn98fZf3NK2dIxm5/z1iYM5d4EKUgxqDzX+gsMzpHG2E6L79zj8b
3oxg8AiAtxRjdTXEoTLZQzLwxR6X9LJ1l6LgXiG/z0novuxeXKl93gtdIAjw3Zih
e6VzkeOiY9kNJP/+FZ2mtY6yhv9MFrt/YgGQIBlR3DJzwdXlpyjL2+W7jBu+8TUl
ikK5uNTFR2Wly8CRKfr97BotRZR2NKWLUGrzVKE/JaOTArvY0IBUrmjGL7hM7B0k
/VAbzbWvEzlDzG7LBXzkohU2czhEMm1q1dXdiOkC5WIjFXK1ejV7UUyMPASr0vBC
TIJRGy0XSddUVDW+H10gZvY7mVoFmCk1ubSHy9qEqTaMElOptkXI0SyDiNn/L2Iv
4vdENwYYNMUZOQJnrMhXRw61H4lYd5s4qHbr9RxyRU5wicUyLCci4llAp2tnTJjB
PRMuHGdouiQZMgG/mTU1L0h2YGdFslcSAQsHDBgh4Yb61MDAgPwYQsi8EM+Ucd/d
YypXeiB/Nnppkxy3GMOQemhMtFMh7AiYyJJxe+gJ0xVW48TT5QTucuWodpVI4dXv
MRyByJkhKid/uKiH1s2LGL2wNkd9sNBcq0+fSnD1xebZcy4Hq24U/jtJPD5WH+As
aXPNP0RbNurpULEaA5+DdffeXAqdJ0ucLGhCNg3mxejzWEKr8pWOaeMSDaPZ54yB
8s8hqsulZfOBD59L7FnM6679NOyftFE22PujNR/wLYgbuthIdona44m89PPNel/Y
wePW41i9tnkEuGOWZfijfXTWnZXfSLKqqEJPXyh/DUCTuLZdeMZSTWKPF93lCEzs
yXMncFePM+it4Lh3wcQ7mQD735zopv2LDVUfXC0zn7p+UYo52utnB/Fi4YOJGO6F
lNbSYpnJDUGY+a7gJQIgzrG/qw/n46n0pPGvKFS8MQ2GHdmFlaScPC5fRGDxqyHi
5Ewtsqecqh05uUCbPiXv7weuz3yL7gWrPUM0oKEnh3dCmVxyI8h0GGiuqDKZMTHq
4USW4rI/uIBfz1Hyt2ebfuBl0MweUObIiQOprTnSCEHItj1L/DYaQbLXAucch4Er
cZi6pNAePznzobkk12U3e23dQk67uIPfUxHanCL+J9vFKrvf5pK2WxxAWyhPUQuO
MUBxKDMO/6L9zF/y9Z3EkpubqO9Ro1UX5w5ykNt2QPStz0R8GdcAibrXnS/FPZqP
nf1wR7IEDWSH5cstPVwa3SL0TF7mPBPnFjVaBKAHJv+AiVkIiDgXseGJfJbClfnE
Llr8LpwNgIP2COc5usX9P3wuDAUtgZIoNhxJxYwwkr9q8xRQAI84ZQdbZmcJJmbJ
91bTN58myCa6FymeAUXLq3q0yZ5HzAWUY64GyGSs7rPOYs0LokAizpHcDBR4dwb4
Jx1aNppH7Yi8SJJ948GN/OtlJpVXUSiTyKVwojr7HHmi9Z2IRVJz0hF8PPXNjl64
eNTVd7u4H7ACiIhSlSDBnA4Gd27ImcuhK7QjEVLgqHi0A8iB+U/kkWHDfw2esG4Y
vzseHYy1fZYCDTlRPP2FrhAsynr8pPoO5Z7/YiD8ljVJgdtTpGuy/wnqFXgqinXG
NVpXhe83PP4Q0f2sJRLuYQtzrqnmsAhlMGNLHA2eQwcd2i35fVwflg4Fp+3gP3tW
aDKyJSLbl3w7Z9ZMPMwdi6zlmnNdlib9Ny21nG9nr005H2NpiJj9hlrLgRewni86
8IDnddAfYepCammxzkDHrPnJg1hrIjOhVx6WjKDNPIVaqAdsj1XZHkTpaKCaozET
tDpAJslnpH16k/aI5wkD+R9Qdivp+UZ3so1ipBVhR8NqeYsRbdm5Rg10RxmnfyYv
LjUVXlK14cBXTKx4gzZU+jAiNa7FrLvUvVOBOYXfV5dXVrBy8UtL3U1MHXG/U20F
Rw4NVw22/qGvYBgniGi7VKvdXEvv1X//aHMgJXswdb2/0j22PeOqoXGQHy2TVmfU
HY/6u70Bo4lumFFh3Sv39zbKNY46jW3NBxb9NF+gnds0Ai1uoO1FF2tzSkcEOvuE
YboEnn3c4XzNhBUFQug1AlDtaVInDd0Ox48oj9ysprkRc70vX700ml93eTYerMPX
p4CBtoKitB4tAEyOUXOVZ2tXWFonA/dSsKMQ5YZWa5Py4+umJJ+i7RfC3PmamfWG
G2EXVSC7G+puNUf+bN0lzIVVKSx/iD+trxuSf3MC9EHfcYFd7rm3ld+lAJ5bUfyz
6tpWsl3CdgBvr+1xNjKF7M7pgAI5na/OpfSlqohACZQIs5ia0kpjbKQd4GJGjnN/
kI6V+2azPh4Y4lYWtkEz367dH9fbqOuXP5LcOA1B8/pinsxqJC7oX416Jxh/5qv5
H4de3TyhesSYDVH79olgUOVs7Bg4Mp4DkeX2oBA56qXkWOOcH78WY9ZeSBFymtgt
XJpltqj2vK1xPxsRDMmfenkjtmht9IT+lMCDvKV7JeyFT1qbOWB4TX3jNlHKV1CO
y7mOLMEQztYBzTYMpRhLBnAkvCSNkuVO8oNqYXFQebnnT+LwZfxqtjub63CBTK7d
tsxZ6Jw2GrCFUq9T8J1a3Z60WualoG9IoOdGl2xStaTXuD7E2MWTkwSf5ixSIISW
gbdXjAL+V6bAwSVuJqERHBUT+jfQtghwz24OYY8QRDdn6LWr7GOKK/csCfFvmNiX
7V+wdpZBpCJ5RLqH7hOjHf9X1t6LTniiSLHrvCLo0Vo/zY3b2bMOtHKlCvhZoqtm
OW2DEw2vBkuXyX5ZDnQC7MgJEM4MmDzAMQWRUa4JByUm5MepRJNuRqxaOLykbpBL
EkcVnCcbG1l07Ev/Qnst/tA3foYuc2O48VgCc1WC8K83Yb7sfMiFrQInsiqRdzNr
D/5qikXeTa+QAiv9yzWE1xj5dWG1sWkgzzADLdMmdqaXgS7XmoZwIHyen/qIb0OW
AdPg6zm+Ae0q+VfVSzVtMHbYtQrdGongBJk1O1WTOor4XHMjOUH0WOfiTmTHBPsX
F2t6NjBRIN3Igi/Kvq5T9Z0xaz7Z4RkBrZI0Vu8oz/UP6fKJ4Ezhlk2ONnGmVk6j
VW0nJmvB6fAgSLNYIn49bgK2Pw3U7xKM0AM+qFQkcqQh9bBJpYrUjcVFMML5CstT
iuQQH9pyjy+LBjtYjVoqVU7Cj8X85x98PSvdEQ5ai9ZnIkkTQzdUcRYQmGAhScjK
opQFXgguB9V2FvtytllxNEulpcH59r071A4jzOboVda2Vp5rTcx7wj9sZBHElv9Y
DkD9Z4LavDUk9GeV+ioSG3BmV2vkkWNwaqQPlypvfgE/PBIHksDEJIyrXeNdZ+O5
/lu8oLYeA98LmFQlg83OsxedBx73Fcxk01CDLzWlENx2NSVzwAqFe/juEvS2Ahlc
KxHleRHrk0Y4seIfC7TvOQeLmBdEWBG5fUY2Bdk20R0HyZ3e0PB4EZY0ta3lm9OC
JyW1p7trHXrz8YerMwrHrqplIl5utiWjqf1BuWMtbGyWRbmSafXxBRGPBLDHX8GA
yanytvSmbJHmBIug51BGMDSmxZKdIBpBgrXMUykpvRnhk6RYvao2+UZ29G2eEC/A
WApQ6xLAfv3kdnK4Maj09vnu3aDhlZZTzNopvmwMlGGSQwRgCI14xi/JoH5WmlLF
EW52/UCExzPC1hEhAHqfth0xTmXZblDX4sqttfEb3OcFfoOMYMNsR/dFiSWLEhhG
iP9wSbfZrL/n55TqY+FW8UBpLRvyqR6/4OeK7xdTwVKQlxXlol9dAMJ4NN8hc5x6
PEX09LAhxzhK4L7TKzUa0SjHPxEvkRlJUlLWq1oHNm8VXY/8RZB+phpWbD/rXR9V
DH4bzKU37MgmL+EVyroDkLmKWyjnkehyVys9mpiGWfCkarMYkjiGsi7psZ5hLFwX
KWXnEzzT0io3mkGZ4wA+BdTxHKOe/VPs+WuB53tHpcbI+VTNrAinp7aSoHi7vEPj
lTkFwdVG4DsuYS/BT2VU3AAH6K8xczNBYTR1dWTQhUVnLRlRqU86tJ03Uj7eVGdv
kUYzxH+Ap5FDUMn1Lkyq5nJ7DjGJ8KRrD+3gtm4CnWzajzZ8KyRXV1xrCLVkRj3t
8+N2gucfbED5Pyg4/Crh4pqY+gu4cdTofHk5ZPf6BF1+iLunpnk1TX7QuoTmrNc3
YNa3YttQJ3GAwRqW2mRv130YKE8KL/dD0RME9XbGIeRZVJnyIELhYBmkAyn2G69R
dquF/DZBVT+QG4pq8cPkTALxFIeCY9XjXqaFcVjv9tdm+gzh3028RGQvADAPxutk
dix721ahVbRvgVCTskeD9xk7U81mHj3CSBNJ3DJHribTmm1ho8n7TTkfJV8BrrPQ
sN2lj1HDkVp1DhUr12C7O//Z2iITyeawnHBXnYj5ALDNY6P+Q4kQ5fIOWJktPgVT
WZ1sYGxXtqsS7rVO1WOAp917POoifUg6E4JC2Z/2CSaSzR25m4VOJiw+4/3mtAvF
RsLGOm5uZBDbSSXe6yYFv5Po4l2+UfU8Qr3oRgFJwobosPmoOqGJEwuUJM1qxxZy
7Al1YPUqJaNMGSfHBSxJ7cGWAKaRlWtrohZP6pyg6lovQZLiHWGndQY+g93FNblN
VtflR4PBsaVeJuM463zLwgqHHYoY8bNi9MCrSmTzxdJTHOJgK99nti0fVFvQ2ufB
NKla+Djid2E8EA+ihXjxgfidoBxAC+Gt4cJKrmkTQWoECjpMRa+CvQ3fG/+HKNOF
lMWn0VtGwxhHwfrwU9tYjTjxZIahmmgn7tM5syu8oEYxtuYdOvd9aCyUSiCt1Rma
IoG4M6oVFuVWcsGgt1BKK1TbtjC9O0WIYi+zi91yhGGUj+StnQPoBgMGkGRvi0u6
eSuYF1Cd2Jfa4frFiH8xpAQp6pZXFhqOkHHYkjKnDI/+DU9qJNr0k1LV72NCOS94
mmPh8KbRh4uGZ0PxlvG0Zmc4rClkzQpumExi9MldAcPTPe2E6QLQxf/EkH9zCab7
r34amqIdbX68gIsUaej3MlZFLCnZl9nneSRUh4xqlZkwg+ItFW85wNa2liGkBQ0w
//katTdBligxuuW1K/NrMumil+OSn619y67QZ+KKb0LBzT+ev+SHdNkHVnGCTFdr
/QAn9GX5Um4gE9PqrJEnH3hPI8gwUvO+juTdtZEQ1Kawjcxxbqm5YFufWfCYIIAe
P49KMWGB7lFqA35eQ8xwyl8dOFNkDGfOk3g86uQZOwxbyt+8uN33X6zNQ6FTgwgK
m8JOKcarl+hnySO1EocR3RL1gSlT6Vr4tZcT9sfNwO41xeV78JH/wYGsEnvdFtz2
rGGUnoAjL668hVqCU2jL3RpzrLps6dlYF/HxjWfIPIBgVDyJrGVGFIz9ppDg9oJz
lUWBiXQlz0Bom/lgBd0TLsgDCYi0Sb+ydwOFfyOjqcTdS2QzO1UEyHhM1VbAcBHr
9BsV4XhYxySx57lCVSqynbjh1Vz8vy8w4E8gNkggTPWfoIzyM2wyo0tj+G9yEcM9
eBUKhOAKa82eUDfMskj5Wq1iH9RPQngh6XA7xHeF53qdk/ZHXj7TTUdD3SxbDTz6
SnRsBqMBnvLISFvDF+dWVje5DGsCL24zqFI9Z4t2wDsy0/bteqvKPY8c//ZPy3TH
eGFWdIso9KE8GCPVfDl7nwMhvzGsyZWznMWvrsJUqAFLmu5C30Swc2mIyqDGJC/2
6D99gU3LUtLZ6qXUanYQJZlV5oMOWvG2Mj6GgD6iIMQCB9AdYl6d4gYU0h55gKId
DAL7jlZMBvuJlxr1IOnqisa3QTQz7Nx8CjkuNyB06ExZaIpWaJiDyAJQtBa7h/ez
aUH5zI7eH9WVSxaETzMd9lbZkGJquaR6XmJ/B139KH1dsNSXpxmvdaGjJnGzC+d/
atMdnVo71OlEpoILZ9HMfyvEwTaKCcwta2gdsXkbMrdYl6rEEP0dOa/mCgKQ8z2a
2SLNBxCY32vdgF/z7qYeLBub2Ia0p3CsBXFELIAzMoEbnhkwUiSGqOf4kCHlDRXs
2xdk3juscTui7Ljv6RlPLYOjq+uKXP95o3mepRjZt5FfQ2TF2EQgFKS0aQXOJUK6
mfra5PdXxyKctz+JTyBGbyJok4COQqJ5AFMNA6Y5troRhu0P79klHQASNACHmP6P
3RbA56+9N1qkQ+k2PRYgD3G1Bo2wZQ5lo+1Yt7GrCRtZCv34AHnlnuczXJNsBRbP
JiDdnhuJuvstOIlHZRvQLnfb7l/hB0PzciFZE0/cY/R2GzXbBpU+90ggoNYGx4Ko
AxKqdkmxAjMYa8Ly/mZyK6NziPdLyjyEC/9TFDoGrdK/h/Jp6NuldHtL4ps+UzaH
Ez5YoxXFj11uRNNvwmk4AvY/gsx5kzSaLo38pSCG3HXALaIdyL6iP16nE4M3Fv2l
6P9tkYoBRQgwwspN1DxF9IQRIcw2ibbiFvBuyfyWd2XJpVxSMXNY2dwGnW7MDEdV
4PG0RZDZHEq+lUw0OTfLfiwL62YREvkzxfoiHR0XJkX6HS5A1kVkLrIFHVaxr4DQ
iHN7WRpE5j6k39u6x14l8V/X7+5tR1qL2hS0UVVT64DZS6xJMAUAcbdCgNZmuNzF
/SypP2tjlW7NMVv5ktEroPFU06tYqRUegxI25/LvJW8pJTm8Mking9UOMXanFXIO
+Ta0hJuClotCfebZH+j8wcBRWsvS7iL2ZBsSnguR2bdRKQoOX+3BZfibyvXDGmuI
Ut11Qexrw6mo+IMgoJyT9be/ikUFUq3wJ98W0tn5yCtngcYEOV0VqwLMAuBbmg7A
7rb/hwhwCVDvX2Mf+2D+BcPHWoHkEZiv4PJ08FMqvesOI7eG67ZsvfOd2dbhEPZ1
GkMF3/Z6ZDoM+QS0I9xZI9yiYkW/kKBptD3gtLhSghewolRm/BRat01uEMca4hI9
9DAW73f15nsZKBSAi/sWcQbD5jcB4H5ZWiv67AKOmRPDOVYOOBD9BULch/bgxAUU
8w8nIph9BXX5PEGkn6vP739Chgi8Jd4hQFwinRGaJj1oZ9rOkBLmz2nDUv0K88dp
tF6uvJ1PqkS1f+K1WBL8Jq3AWA6qTEs700cIRZdWFq0yQ8T43E/NadLnzz+voKUY
hKhW7e8hL1h822xZprLYVI4ZogrHp3q1AN/y5N1IGwZ/llxTCPAtn/gc2VKO7BCf
lDeiQhCDngfDtCXKXShd1H179voXJgntXvCGD+4InROpQU++N7izbz+J1HzimmCh
XYN6mDlAA4WTI6+tzAGFhby4JclgGyEiiGQMFAQBHHuqJwPXRaVJZ3MY0sG3R9md
rDSNiPHK0aCZVFN7WZM+b9R+0/URMmd5yNEGfCUewEQiEM4K8wXdd69ehXqJ7zT5
dq9jqZebAE5iQaGqnrPfcXc0CfajZJdiOthzmkNFa4fOTemafhZ7Qcufn0c8hjFO
T+tjpQwr2g8s3mE78OcJ3lXmJPeLwdsK4uaNFvFauNc/XpC7x7rgwoTWitNdkCmP
m8dDW+nsiD2cuWyLI+tq2t9tD0ecPU1lrJ+JXCKouQOd9pXXG9XOZTlx/CxoRiEZ
NBTlo9WmuxfGXFNO3lnOAPXyjMvHoP9NEsDX8D6Q0glwY6Zv+fBchNsyd6zTcdeW
+gtv3oH3FAltaMovEQeiJ8oCNdwdw5ngFk9RPSZ0Z6qkKa8XirtfMsyZj8FEK3s2
5HzT8EM+SlC7KnEgj5K5o3yCMtZNqrbTDcCyGBtbzaj9GqiKCLSoPAlUBWL/JbGu
+D3q9WWT6q5hnvJuIEmHkgwVMys4sHadEUFeDpQbIXS27Me1fqYktWoUyYNn2UQk
8tD0OSLPtrDfo1AxUD1GNQqBR5tWewe1MGvIHqWFF8KAsbZ2joQdyAmqi+FvHbRF
4DUWJMdTSXT7xR3b2tbJgTbdAirBXwkgxPNhtOXW/okktWbCuU7Ga//Wusmd/BKb
pTi6sjePRcqyywdhpzwgdMtdMu7GlFyuqlB/Yj60XAR0sWwtUijkKxIO2cCC5h3c
DsLgvvi0xtazOqBdSTTxxMvqep3LT1payyCNYv7scC7Wr+JSdxY7G02B0PKuqKtq
sZmYvK0ZtZ0BXPi7IMJgH58kknhhNx7rvLwzmKKD4BCOnMclqmZ//3/nRExP1daj
Nof5DFCNS+BepksyC8sSg+UNftsRKe9LdVWptva3kjFzl1YJ16pP/oPYEesI0T2x
vIB7T5vcGBCeW0Z+aHjrIcpVF2GIuo/za3UNzQLmIA6vvjh0aoktCcrCA26bHZHg
5ZeD8cOKcF4poUfjBE6BgiBGnywoiO4mlvV/vFB8S9bPxkkStjmrxNhcidCWPjjD
P05WlLLvrhCxMjE8QRHXaXIMF4cUMAEncZl0BGm4e4dEPn/6AkfHBKRMNrk27pO6
jUFSuImUXUITUlW4Li3Yv+MTDFAT2yuo5g5P1/5bOSVIK+9qd8LWzCwdHtxi6SMm
ZAJZsWvLriT/+ZnfY+CfZzw1AW0RqHV3aRI4Yv9tioGaNDlKMYCXzuYJp2DgjUde
ZO6IaGRcTOUTHxhQB55gZ3ZCqpGY8N3/eFD5DPVVU6As7WoQx4x1W9/Dd1ZhMelR
2pd8OK3V+tgB1X6b71CabKAC5fURnn5mZIrjNEkKegsaEh168TGAgwEVXMPcI9gY
fcVRlX6rriKkiqF74KLBINoLAJVFNawLbDUPZayYwMyyaCm3Gw5rXqHzf5IRwKUC
nlWPkZJhZRryUqpRl9PhYDVh8/P0mdO2jQbluiUNp+Q2CktcJ9oRBHZSD/hR8nCv
pKbJ0ukEfZZ+Y74KC+XetfGUdH407dAmsclF2g87l0zyf1DjRste3a/I0wOI27Up
LhOvQiLSxGFhVW6EWNmzZENSjqjhhQicfJaUHg6NNzG1Fqs/R78leNak64mgeWxA
NtbaUdDixqOlq46AwHbOcv+M4cG/Ll7UJePYvbchhawuqJR1f73gSpdYc5ND1set
CR3W4IVzK9+kHIoiuWM78yrNk18KLDM8gxwRvgf8GyOVgss/sm2s4urBTdJtabwo
mLWED50aiG82DB+i/4FFgUqYUV6ILinvcUR++V3I74dEqavyAAD4aH/SvSdiB0KW
E7ohX3dkuwi2nbAFDfgkW4Gi+lScMEf+GmnF0Jh2m3MvuGl8XZG56+DJ8VQiLkFa
gIGGd0O4IlyWEHnMPUVh1cx5trKAVytA8r80xvrE7RbjMJY5PzvBSWYr94FHMO1j
gYovVNP7lgYDFe5CzOIjMejL18bxVnTdpRCuhcynSAFo22DHn6qZxF4g+z++42vm
75xbgsxgBARR+lw/U5R+EDGKWvdwy491tLney1E166svPmfr528WTVjEXBfiF9Ql
UYCQ5yrljE9qU4zPhDuAQ5gVBftIRxQ/7SCkrn24uTYnEtAmJylpVqwdN4ItsHwY
Q97R7ELBRr79k4k6G2fKVcFcsYfujCbgtkyd3Y6Ih5hxF1qLcLfEB8Vtfmbs2Ndq
lGwTUHyIswyf7Ktp2zryAHmQ9CBHu9d8+XkYyqXKRWbdv6x2pP4ZfCGxRzPxUxn+
lyla4GkaGrLrKc0MOLXtP88d+UAa7CCzg+UbHvOoVbmxcgtjthv/AfUiFPJU/CDc
QcN82ghLD+KHdrvE/vzJkzBoGlD2xygq3l4gGpCA3gfuI8AbvdLYciH1O7XJoeI5
V8nLUGSE0YQM+vBOO98HcJDs/Zl94EHIFhSiCxZg30nLzP9OnUcGbpVlFmrgK150
qg1WMd3uDsf+OvgBGug7KZYEkgiXY5q6V5zNgro/Leq+1HlPF0agqtQHEqRN7abt
OCvOlU90KytFlN2SXlII+gh4+ho5PRCiMAM9gUsjg9Tlj/mYyS877xL8DtZAjXwN
QEcfoG4Uus8+CxovvQ/MYJWi9ccwjWeIIzpuN8lk0eax1g8ncNmDDZK5LtaPjKmI
9wmD1KWrWAV15PRfXLAEtusqFVbg9eoTVKUVIDIvF92nhyvadOhvQY28dZVtmvYl
6Ibq6+1blFRoy22U5Ty5VzDOYTGfcGYUKGR+oq6fgJBN6aU6lgJDiijvYHIZ5n9S
O4hqLkNFioPiLeWzSgJQotn2TDVGEA3ttrPwtKGE5K2QYJHhpTfy232Am7gv0Dpz
t1jeCNyea0B0tZ5K2okypxR0UAYw2wuQMvCSesUH6/vrpW/rR1uN1sksOy7e1wCc
iIgRe+oMpz6IhCU9Kh6Pr7n/9rsjgGKBIohjfYneU6L4lzO4GQXBaWEjhe0A8nzn
4XAz0bSb+hd0EuQOvHscvBm6SQ48jQy/IQ92esERccmybd65GlzVu8fnLICMBbGY
b2pRh3/o9P6dBTRv4EOKGLXiFsA8WNfm5+k4Std+UAeJ1knrg2PR71Pj3D6JZtXG
nbCJPo3J8a6kDQR2whGH+HVWUdQ/YoN75iUW+DpGGdsD7pQ9IcJVuLE4B/T/hgyp
2UidhSRbmXWxnMIqtVNLOSap/ZMD3K2gEj8yrlha8qEaImqqICs0qfwcqyl3tJ1Q
HZEX9RSW9ThmPaaNjXR0amgHC9ZjnOiYsfHlh6TUx4OGCB0/M6toB9OdZPb06Q+Y
YtnT9ylqE74LVAlEE4gd3VlSYk5xOoJDHickt1Fiq5bm/UrQFIPFjUYt2bAWsnAr
glkrInnU+ggIn7qHlXJjNrPjQNJGenDB06cgzAVkNtRE1dvHG627S/CTVTcuV75l
VLLtzznDWOIzmMFZy5XbnE3bx+0wsXdr5ztjyRIa4Yop4LtMaS977SkrQgxAHNAR
A+fwOep7n7i8tdBmuIKy+NkO9mvZswg+p3VpBYDG1PF1mosj4UUp9+FEn0JmuNXC
DD3V1IK4tMtSiX6TXfk5qm+keqoQhjEliqw26BIXPGySu+TaXWOOjW+8qab75HGX
ToRZicVGxezQCdXER5toQAVO4d2XUA8seK6t9AY0Jo5JuX15LTYIyUAuKSSdH44u
4vUxH7mkNeuncdVdz6xMwqdMUiP2eM7PQyheqerK5okcvvJvIEuTJef1TT0QK5zW
Hm80TiHcUowTGHsVAIF4DLfr+bcy62NtOBseaM43ceNDs4Ku15x2nsLAIoYibOtD
zfC99Rdn+wuFqSQu7EwNksrf4j26RWn/ojcKa9EmXpzIWphZGQmo9azfw3es/Uor
N8Y432F0jCSDwc31lrIXeZZCiXKjbwjsxM+O7wwnuplxrPDMJg+7PRQW+F+lczy6
gnJLKG55RXBcjN4ET9TfJbQ9LOp8VGFC1WZ/PauD0eZTxPB68EU+hcNocv7y4mWC
R3tnFosTLLN8jrXE0zvTNbVyfzTUrWriibgGksJEXEeSx3f1Lcs9njGmGsdT6wcR
iZ1BIUSrIA4VOXjLaxE2FGH1Il0i0Je8B6X4TjbxoT7V2a76Q5Kqfwmmf9A4ng3s
tHkExje3Rrz8EjKTZfn91Nc0YXNa9CqBndWyukB2TrVpvuBWCe0acprAMGPrInzc
PTeqg5rFmU/1WE1R6mQJvbnIunw77uskRljmeGSo/eN1txQCllgXq5D703qhqQhV
3vtM9fq2R1ulhZS25zAp0D+LZ7pfTVRt+kYIuOgDUcD8ss4uHAd2KK1M0XbzjChq
qUlX3JhNDLvpq2VYhC/9ZlEW7Jot6bTnP0uPh6VKbk7B2YceCWUItMJX01X56hiw
Kudonp8+cci6P93wWUjQ5iSh5K9NOZiQclGb7g+QftlikILeLq4nLdVjpLPetWr/
luFG7pLLKVSxEue+/JNZGcp6d3o3eAQKY2ED9YQF1xeLyg4ubIG0+/39is6lqdbS
uRU8Z+pjFLLXBoJ1pACZWGLHG88kTg4wbRdmZ2stLqNDrOyKZ05C5eILJDoWXqcw
OD9yKDrccsvgjgwE3ndStj51PvI0/fJ0SvFIzr/fCK6TowcjzWYmXsCqtEC6aq9s
MnZccG+R6AEDM6q6hrQqRIOQVPyZ1JwusttG8war9ezQ2ve/R+BPEENRcufMUxUn
hIslAG4K5LvDXRSp/D0WMKTnFC91Azxag7XE+sJApC/Hduj03InR0o0mCIsUm/Ol
u3VWBQYlWiPfhpKy8hyQDSiTx+YeqsCwyEhrsIFkZKjYHN3fVLnROI2NaitXg6hD
E1c7O4BKQ+P1sXTz6wwKIXuCmDhNT8C81t1MscuvbeL9UNDRGbxiosCyUv0OEEfI
XvYk5fcwoGslew6xPIi4EJoGwbAOwTL0JiXGbgT0fY9aUkva7jGHds+TCVxDiaXC
UMCiSANgg0eB7ErLsuHdt7qylJ+IzqHYhTSHWMG4h/tZ58j/jhAnF9mbr++tvrXc
rtPxbO6YxJ/AEYd973pCWJkQjYaArAhrZoViGPG2znxicXm6LT/X3kCvECMGyVYH
+MnlEqkmFZFqQTM68vO110eUGt23P5iw6CSq3ns4/6XVtsY7+DMSLNkFuLgUFfxq
x556SYoP9SPn0oGhPnJF1a8Gt9Aia6g0Gq42J2wl8m+YzydxPw+RbvWAdMZLYvxf
VyE7pA/3lph1/Fa2kL+85Xn0VUcEyW7tbNVnYabWwXoGkNml3I4uxPeKdvowMl8B
vumv3YJ5j9OymmxhDcBm2SnyfU9afpdMHUXDCHAxSiQLuv4fCW5GGx+2fZmEheQA
WyY/zFV6Dzo1BdSGXnjwCTsTxagEW89A8YbKfBHUW1Hcm2BUmQSvrJOJkwsbhfd6
cD4YFjMPlazoU+sJA9lZqSLS1JmHtrEl84JgrZXTwI/FVJki78bjF4NCsy7rSd0f
sH5DbkjSAJZryXAbVCTlZ6BIi/+GOf9kZiB0Ny5PTL+aDo4oVoLzzQtB9/H04hYu
zyCFsv9adpPHoJh7q85gfHgR+dDR2XOQ+ntpC8PnYl9y8jtjijHVAqmoH+P4E6SW
nE1T1fQ4DVMBhOdEmR1F62Xo59b7dbzllZ9x/D2O83k0ewBr1a5G8M+QxU3EFltt
Kyh8QByE9ilbBZ01PEMCrYIUt9BYGXSwGlV6HfODB4Xt/UdMyGmRtkZlLGNWL2oA
x6IEHJfY7U3/BTV/FvPrKwtv8pIjXPuJ+yVfHmDbfxbLIRpkRSuJR/q7NEOYOZoL
4Y+M0PuSQnYqZBCoSqWg4CmZmggUfI0U//9GeZvvDO6ZKqqwdL4JyFNpBJ4ZHKev
oJft4Aq+q0ox7PCSTUVnjDE/c9+r15pjDGqt9xlY+Irf52dfMwoNpPUy58eZwiMU
9NIpx9ljw2IoC2G6rNH0djLre+CSfuqcrd48BjjPjEYCwkGBRyzNBmz2RzbepiFs
jjXfDVf85Nfbr9YL0lbbe/Hdfg2RF92P9Tnn8xur5gPnkgGNQ7+aoYMRUh/a3Nhb
t/gxpjl9v85M112x9emWS7SqnXitTgKk6lPEzSBRjtaewZt/UispFgZ49F91ePOa
Sk1JZVyK6ve1SMCDQ9RlbE2qpmc/jgZHODNBPZScNd5msbslJ9v91JQwCIKZyOMV
s5xK99wYHEDm7JC8SqsbT/Z7Vrmoth98upw37r8UUdvRM9Ui/oRYGrWPmg+H6kDJ
6bqBgd503klaFQsyqJstKSsneukm/jNGcjW7HS4JP0d+20wCbqd7D+wf/4hSaBcZ
je72BR4OIQb+NvrXIZN6F/ZG0/TPBG8Ok3rkeSY6JeHQqmZETF+3zsDGBrX+d3H+
uZ4gueqJ80g9CcIa/oKWiRlkgFZRiE38KrcZRCZgGwlbi1uwOAeIvlv/3EMUs0gX
YH4Ulp0iQfNPdSbOQrfjTeK0bVgH+RoHrKasTRqlR4czFVtY9CcwxLAZFRetOY2p
f6PsDx4/FD2f2mcCjo4lHOOR4n8K9na6Ly77BwRGSn8ro3eQyUQcnq0qDAxFdYoS
WP4V6R+JCQESofCOOPGDSeFDZ+UVRKg9guKCDxEBtvmbz3929IT0Joad22/Ybahk
FOtyEX7tfDUdn37F6lknQa0f1rzT/ab/Ba3UBV9ypC8nr47QQNBFM14xJbTdF7e8
sD04DZIxRxEHqegXqgn6JgYBB+6f3AmXo3GlOeAoS1AcrZ+aVLCi61PnLEk21p8K
bYT+6Z9chSN0XTm58F3/yI8KoXQsJZhkq4UY5GODjj+BT21+n2mIrZjv9gjxGwCU
uqJUd+qbg0y1f55TZ+E0kGH3sa1cWEgEpHSC5dajHNBczhmNGg8qPs6ZWl0PcoCm
YPg0h0VzxUTjK30g0SXn3gZDK/Os+0lm0YLfv+d2N17EhLT24OnvlyAchb0oTXEY
QW8gGEX+5xTJ9AzoxmhMSMEaVwBTEbTNyyIxkHfoG2UlfzvxSuCGLtc2aYPHsU2a
ayoM2vOF1bo+q2iZEpHe9YN8EwQuUSbQmwDKfgsUPsZzHTSuKG1M4op+O4ExLaiB
tXFjEoi05n7JegFXn1bXO+vw2yUTIh9QqpDCDuhbtF4p+gT0nelr5j3d2+Hw71Ob
0PZA1pvWAQko0MHo5iJatimglwoZaEtJgxrd6+7vaVxUbS6y1aRTGnG9GlndT9pT
9BBJFL4JaaRaOH/BFmxXHGEizQ3yEItqPO/UoQBmyYPshRApooe8FPH/+VzgqGD3
CsrS10Pgz23nXh8uy16BYSA2uxL5qoPQUQ23H1kjNv7UN8b4+9q9Pc7Fxa0+QTAQ
dFdW/bAePocOdcddAfczPzfxIIDbKJV0l7hQNN0+Sv6FZZRVaij9nkHq3VUdIc58
2mWnlsx9nJx7vuyHr7x4gAi2WXgDg5Ht6qy/O04ILiGiE5aNGX2u9lZB3jQm+KVb
pciXQCxdfzShm3mWBcDB6Cl+YIBwRVmyt0ePbJTUfC2CEXPpnB+csV5FPIbkTYhy
FW3yx9BC5da3Rc2/b0zm82f2Rkxs0VgwAj1+USnIwUeOD0nq6+IZooUlFsJ5OoFb
JSKjTFkBPjvEKWa3uHwNeX6PcEF9OX62mhjNI1UenHJeLUPvVL8jISTMVJ7mdQKb
aMSG8NKDSEFoZsSr7Zw/wiHeKHQFVKvnINT8vckhA2yHgjzDj3oGAWk3YLTdtg/Y
GC6tb6cRRdwET+uJY6YO8OlZJ9pMo0HyI1TE83iLzzdeAeQRecYeaf00RMrCVExL
8VHwjZ+VTOb7ugg/tzvyn+TYxoRqu6TfBAf/+7T6Opspf26izJfNgiWY83eMS5jO
KshWJj1SzDAKMpfMrF4rfUl/euyND33EoRkrGy5oVHaatIOUvB1O9qbjmyfdtdMj
JKAM2Qk41ozyLw2qCRe5YNtohxT7zf5AQtkTc5/Z7nco2JI8ZV+E1mIwnBHZcs4Y
hQkfyk9wNSGYCk6+jL0EaE9WEB9nXqJXhHy1mZGCIzL4mey2YGLw9bDaPTWA+cjM
Vaw4YqOkvSRvElixchrQOgly4OiCCdczdsgrm+8ZHdVF9hlYHnRWLOyA3ko/zvE0
2y7r77IL3zOejOeNQEkovrAhh6CUpHEfTkkej36nTet0TsoDtYU20XLSlhxbFK2P
joddrybwf/gXw1J5t1j0qGhpmgv3zWq8qOPM5D8mE9ZzGMp06wr+vkeyTeRBjbBD
q4mI/Qj0QgqsP5RttjxNhvBNG4wR0cbgg0eDlQujWJeDv1B0JE8JRpNz6Pl2SljM
dwbn0y+RRkPjjen9AF80SUd7D7gz4x/aMseiBL+eayBlDbknEHKl6RxZAHetWc0P
oqRCaLFgkVGu+jnRAlc5lIbARtvCYoP+jLepmoKFhWLObZzajZSdYeCNoIyuTp4A
Pg7huk/MnHdW5CLSX/SoX6dJwEmJXu3RXrOPJWURzGfWKwFjyM/SiHF7Ig6Hm04x
xyWXPDgkh0iZsZGsSaaM3RaWXK+EBIn77PPHOgi08v6/FKezmZq/FbLzVs2Uv535
dQGr/PbEaYQqOKdT2VbluzwLNhBrSHgcvlBmUw6U33X4SERewEc3S3qL5LYH1sAc
DR/oVWlJodJ+gpaq69Jz4CZOKLvGs5JdQ3HjKvbVGfeSGybjDdcX2mnFocAg0JHC
sJ/hwUEzPT4Puk4aTIcAdFMRu3Kx8dnLKjp03zJcpHezaYjNyMBvKTfkcCOZLfy9
QH4gn8sJ742obYGuMs9FsFROeWL2qmrfgVTQUSuyPk/Ps2W7rbfM7b+PW38lRbxu
VjLDJ3AdRIBqiekYFcevmL3fakFm38UyVUw+Y/z3iISsfi4Vf8UbtjyN1/n5V9iS
Jd9wFUmsE3NhKraVPNNklm0wXflzIP72heIldINeXY1yWSf73gLhCnrOcYFoU0Bt
TDrvkY0bK0Xds3R3Rp786wH7SxqYKZBtykAX8ljBs9vMu2549S9I5muWF1gZ19Sy
xVR4ky+Xq2V+5j9NluX2zM187uXQne/FFtXiy88fz7OJo5Zy7U4tai5zVyNzPszM
pjfp8ehchhhlIjsAteNaJACPD9LP+OQTlABW5ARViJGwC2tX3SN/1ruGkCxf0L0t
J7itnF1cYWUgIOfyXtt+lBYKgwKfHih6qjbxrteeIsa+h35JgXYIUSpwMZYhsM/H
mz8Fcbpj2Dd2L/aXnscBlSv88EpIaIYz18pZ5AGOV9Mha+lv1C2AoXH7ZYdbwx+K
qpLneK85XUB/RujPq8LKR/3JAFWV0BfN5IamA2A7fC3RQ50ipPILz3IfrbZmdeEr
YoqxwC0tvxWOCOQL7S/wMy4DBlMMLafmFj/v4ZnHX4Uuyxozuu85d07EhdaPTpNK
yLWZxOxHIhGWgouEG1h7yU5BqGQerTqEogQcB/QbQ5TOtO4J76BKSUgefjQoSuv6
/dPXH9p+k4EmfCG4I1tXPerd7udaODdijp2kv5NWdP4IcDCgd2gLqdtRLFEazhfG
9FfhsMqmOsBGM4vxPEiNV/oA7K5oiSZHBj3Wh9t7qtRraKj3Kcw4SYT8+FhbKEkS
AzwMWyzJVuO/qs6mQu2LIdwF87oJ7RNo1xvVoJQkiYRyxrUXfX80RPpAfFaqR2Xk
6tnOx+VQ0ECNFB5uZq2lJ2La0bL5zhPXmEKPtYYbjDF6Y44EaoIZ93SIfp13PD6T
zDZvTlP62I1r+pgLNf929kmSV/KTPAaAtKOLC6mupikDDheI2dH2PRjMRbNB1rCv
yZz5imgkPiol28qf9X3vbuEDGRZAisPMDsT7Oo5J2XBjdKjZ5n3KbGU0bHAgGJ6b
kOKY+A3THLqO7lGaPM4FEWb8BmrLd5j7cra3Sxg3nB+c5/MWl63VqyI13DBsdHq0
bkI5N0fiB+jVVvi0FHgcOrwOB5JpzCCKDZ+cpzIRtZVCcrlHaiOlLCBKR3gkzuZf
zGlegfYTGA2tCRxF8OVILicUEM+eV809+Jbd13FTllkLWHL4b8KSjXb8hdejRt8J
eP2zA2MCMtEJy/Y7ehyUD5IU8iKuNNotseXXlwRbbvNhNC28jQgtCoZIbglqhEZr
R4dcv7jjCouPd7RaniwKvrHpBQVDKXXDCGN889NcUnQhMitRipltQ8Ow7Cd+5EvY
wqoRnyWk+JXgQsQYuQn7crdJsTSWtDO3iIeUdpj/hAmccgEeZahj8SBZUd34g9My
kj1z/SBhxFLYzLMh1dfzbbGm0M5N/R31tfweAx84MHLwD9Yx12ye2ltsb/tsjOl9
P6GcE9GRyXLrIM996qcHQYFiIwAYy65n8i1Q5ZhCBgLYEWdZgfP/svgHhvEnvvRe
q2Gdl96TD3zZYKy6yuV14T8baPkPU6kK9e3brzfZDPiR53A+80jroRGRv3SKcE0H
H4eWJHlScPheB7UvNLslYe2HjzURBxlhVW2pu3J+HCcJyz0jFlMyC2TnCxhlxGFd
zaIHMu5LRYc1o6b808GPd66IaZ+/jGdLqGsRPVeld4uwKskVTMbSga7yCUcVPYpS
EoDDu0WFNvdOTy1bem/tSVgAiNWNq3cdKPnbpNo/wdsJfjIPaNSzOy03wif9bWtG
Zb+txJcAAKiwN81BL/TobAlrmCbY075uw26hRrrrVA3u0DNyeK80/pMup5XK7y8w
eAAxBrEksoAMgaoCgNZk+a0N6ENBSgb/H7tKmR1p5by7by1sJabSjWiC2s6pmF34
pIJbCbiiZdFbPk/tPLcicR/YIK7NqbzqT8vrdtAXDmp6HcjjErgNr4y4A63osg+Z
gc5uopg0fONdqZ0v8l8H0xFe7sOnSMEZ0uHTzJCRpbKzFFbZeNWhEdVE1N9F1eqM
4ukuEsaW922vNglTc0mnzOi5XYLPU/csBUVWwyR6KXVS+GSwYcZS25/uQjDBEyVp
e3MwnUtcaWq5bb4J1sdrvtMcZppD2T29QFkU+r/nffGKRyMiqZQCMuGZ/lfo8ba4
jGdBA1mJjQIrNCztbKNRXOPPIbFTjCK0y378YyhxygMrqCE1FxyRNFzmEVj+MjBv
P1B2V/2a2PNo18dmeQjPbvQeq/8HYjMnUgbn/E3C3sBgLCN8hvdnTRKNPOi3gFMC
4EPLwv2dOEGuRB/dfOdRnOfxtfNUVtJmFKyJnBAQug9knFLxEQc09twfKNaw89I4
8+pQhFA15WIfvOv0tXbUfYiT90TWwporpXkhcChf/dNHolWDWTuaFvfHoIuQi94Y
Pjz2zbVenQp98CLckNxDvH7Fwv2aBZhWGaKTm37KSQ5TLWfSzUtNoudDWMEEPBjO
IO9QyiIYNNp9uondaNukghf7sVcznJN28a1EvORuZ/T3rFrzaL+Y5HIE3hpJra1x
ZeXsdkFudWd9m/gavEa2J54To4NtHg7vdU+N489m0e90RRuKAR4H6oGu2d1GH/YQ
LcOUIhCh6rvxhDpXuBtTUierceWD8XQwuMeAmPUFnD4wkCgmpqH7BpY1QRypF2fF
BTq6gWu77zb9ch35GJiC0QwjQlQCLFyP84XA7nAxvF38/BCHZtjXQiqF0jX0M6zk
43SME/swlFcf841/SyEN6DiwSXcPj6PEBLgc6X9SVFdBm34QaGPMwbTA1TFcEG73
/u0cVxThU9COFOoNE0KYFn+l98UYnb53WyqgjzDjmUF9zssFC/2zvSpryWkz01cW
9exN59m93wC4YWnLEGHiJ5Rybgf+vWD9Sx4TOtlsi06B483mmy2TPsKeDMC86nKI
zUHMIDs1XeIo5rv6iZcTE/qZKumBFYydLcBWdekzWFeg13a/9I61RB6BgiX3GzK9
HeTjKlEZVGnft2RLutwDUnj3WdqQLbTKjG4DidU+iWx+wnHZCDzwm0OACmlix0/w
yGLvP7iM5Bqk69rgGZY4FtCN9BhOL/HWu3wTQaWQbhxPGK7zrkRZEkdckO1B1y2V
paP5h2PFlAl8/M63e+fnGjjLwe3T30UG8bgaN/S+y7iLsvT2ra9e9K6LYoN/yraH
3CysXgZ43dPGdAEjRYfsPzYbFOkovDRYNSWZ3uXGJAYtj7rulQ6GVQikj1uBfobP
p4uyp5A3opvGV9NzB4AliXaFjCd/fUh2DW0LvNRtrVZzz7rUvO4qZp8OWvGPjWLH
x+r3L9RJ2+j4cnwUgTt2ksKUe0R+aHDEyal82oDX6B2L/sEZ4mlXkaERhP9EB/XA
yxsjoj9VwIvoD61rIF2tL4O9qR1+8PAOCohkdig/tv9mBPHS1t+LV6+ghB+Il7pn
W/7zDab6vmzaytds9BoHXSMnCCVALOEJgFAOr25XGUl4UvY3oHFeI5B/fq7XRDDM
0NudAFGQXEWLPYDXfPsMndwI1SmXH/VXMRQF5+ZLh8OzZNYfdIQEC8yhTmonqoZe
vMYf7StExhGXLb7MkJuntbVf37V4IczI6Y4EZ380Yfp5JO1NuRWURQ90NSpJ6uGM
FxBfc927SMJSZC6EmStxIFbExkEYJu5+FqYH5phMPfOM1a+NHSxlTxu8cACsE2J4
8P0TUd/Wj7rvs9dxTEOkpKuM2dadNWZEh4ZI06oCzhUeMRgDT4hMIgQV/Sx/vvj7
/PqmRcOn0lKz04llDdOen6QILk7VzRKRmKGixNk77H89y+X4vPMnEUiPK2yCbJDE
yhmuXLaZEhuRsmdS2eh7ULFEyyXiu4I8s/yp7Av7Ij40olLzhg1Ac0tBj6JC/Q9f
PYafrpa8xAWE/bXvv5Q5shuoWMMdREneUuhXMTvLHHkV4W7Lb58eNVMTXQLJsdgG
3K5tccqEGPblBH0v+2E6lAsPO5rmtscCVt3mL8/kDw4NZL46fJYN1C7oHYb0QvCl
cNRhACnjRLEnaJviT2XmPQ/+jKkFM6xtyXzkM1CTaF4CrQijyOa1b4jsmL8zIbbH
3sDyi7zDGcuJZxyo4BDqad2KKwzbrOXJrsDt/lyXKHmGkuy8d13cuFRP74WfgtG2
FCOBdJOU6qY6gN3dWua2lmx2ERWqcwiC0QPWGVyL0Ur/tAxVfywzND6lYMrXH6Nw
U5VwZGnFhWbN+JN3Zux3jgDuUZjxmXcdS3uWgf40bAYqpcHCxmYip5fLQs4KxMne
RB+kF85g8H0XPhB9CbtoQZSlTEGeOZqxqdca3CSejIqzn1/wmrZKl6Uxx8XRaKpn
MksJKczQlP6nSs1T+SY0pxj2qgSMiqAOss7wGpjNbVkWzwATfUZo2itWMwdTgHN1
I2uXxx63Zi09+iuuWddhbvpRUsuPYS36s+OAIc3CDCnNL+UqqqLoswu2Sz518VBM
mNoF1Ru4VdNovbaZyN/g4hDGWpZj04B8atmN8StZzM/PY4xGhJ76Ac8Qe8YYjH4g
SChuXH6uIcfYlF9cv+pxJwbaHaH3TuABleDu/9fPPFfAVIQGvEqRjJP/M2YzOs8O
XR9oH1CMRppOmU/7IZ4YJXcqw8xoHevLa0JVKJ+elpEpvB+tVF6J2LKWw2y34tGO
Gvfa8wPMgZTFRybrPP7BVncc+lK8efH67volxgavjvqmJL5aDQ38/5ESWqdtdCSo
1qZIxF/cJpHTD2tjVNUBPGaRCr7B097k/VKJciCMv4/sn/ZZjGkvx50xGF7klQPq
wPimzHJ8PFWiCjCA7BrVo8y9CCa6kWil+Opq3Ys3IHmW0pkat1kteZyFODXX0wGL
nBnZisft4jf9OQqtlrz4l430p1ldgTcO9h92AQoFf+hYJurYiiD0YcikJeC9z/SG
DDWUpx5E3ne3hRv+jhu+XiRZxfkQ0p8E4G8HuoMbSNdHdY9F5TqzqremCgd+O+Qd
vHIz5rveqHNJK48hX6/e1uxMtjuYhP8a5HzFTDZhFAjSCmAvgkklv8+oQC4XA+W2
WTh5KeUwkUl70Usz+7Jhpi8gy9YcUTVxJDkh/uY+c8Y+K8EsC3ErwWigv25YkLR3
RURF3aLX8RHxaMoe7HZI7TGdRIhKikz8E81Ti67b72WbyvIqXc5uq5QKTg1gZzwl
B/w2IykCiLIxZ7kj94dxQ/E/8PEUe3kz7GqacRY0IpahETJnbaagI84M/4qR7xf2
Vnj+V3/dVsrpnbJEiCkzGQMZNGXPYT9BeaKxREt1MgO2WQX872wOhtvtRfSJ1x/i
dCXjKW9Ge3EJ1QYJcY3u9V6y5eELnSsqNskUV+PW/PnTeh6Wx321mA86pgqvMvFd
4ARuwx5ATYcgn0r+jCsPtykXWgVQkQm+NBvm19tzTqyur1nX41+P1ZuTXMGS7+sj
/lWH5bYmJGW8rt2TskppgrG1l8kAbqT4a6DEOuNrASfWn9ZKcCRolrZqPikaEtYe
nJL9lULIbBRazWQpklzESqODqmqwyCEvJaZISlBXECzU0wFe1btQj8qedQFeutbR
8ntwl0zJ3GK7tsS4IX0jmxCKwLqZhrf69MEldHnSVJgWRZHm2DEqRhRn6jnQB0O2
li5yLuMFBvWn6lf+NAOx6DGbwOTweQki17fRK7KiXQtq86fZj4FxuNBIcV3yKuHT
EyRVYZSAvcRbbk0eSzACO06HmUrvdUmnGJ8KW8+ghU+i77E3qzWe5z1TBPEJfwYp
xr7EUk54BcHF9U2LsHEaqflxLw0VAU/xapD5LPqn6jnLjPZ+U71bVCg1rkvOgnor
5oofK9LrEC8Fcc+oWK8z52u5OHXvyZs3owvr8HSTvfayEEwxwyFv7mVnbUFA25nK
5CTTXdHLXVSWkLXuBexSQ8yOvJqQnoy3dkOOL8ey1h7wtObWAC2+Fv1frGJzwN0H
7yz4xkQgWm25DU/Sm0Ui7mp/OxNtYupi/z/beLz0lzP73mR2v2WhGqn02CXimKPs
XsK7EsIVwtvZADWldXAzZqd2kgqaDN971FNy0eiIW7+AwuW2X+N2ySxMhEAm7Tk7
XBo/ukSn7/8bdmvMfnVCg8r/AbLQkN+6PqXDmvmnZAY0WLZe68zkUmvOfwbQ6fE+
+IZZIb8xB46WYwweo8V7jaU50/Gi2ZZz7jg488a/+DbhRivhg36rmgbTpwHPPo4V
vn8I/sbRl/8LDJu7oiP8Z29ytiZfzm5rZYs9in6+0A3c2DeI5w8zEBRm2Zreuqvb
966iw4+CcxImhGKjvCBSsxhu2OdBRAmGwSMiCgl5jT/49HB0lFX8+S6QS2gKyKhw
homtoxONZh2Gb+3jH5zhsZb2ZpP1mrtj88piMP1WILtvnsgBpqoZBDdto83GUXVR
ziOqTZmD1VnFnATMZsM+/RMiQ1rjmmLgvZD9hgIHA/6UtOQHwM9AkGyVRYXLzr5Q
gikxaKywoIOoKjufk7sNOlj5w+++qfcOTIDU3ZuncNNj6Md0gq8Zl3esz1y34PCr
xRKHSkZC4R92rEx3zQiovq63rBryfmIl5N7SMRSLppzpox4GbPC8NOqBkJnJWUXS
JxJtnx3hVDZbST1QREWbQgCLvJ3RqLKhrc9EqnyZpkSmpfi48C+slB64ZPYuMpb9
T6xNwEmtshXVXO7GQLbZ6NolvotJC9fyxdBo+5k6f/gZdAju3IJKES73R0t0ic8v
JWtj71g4MBT8RZCrlMhBVdhlMwgLAtaM80XPEdKCq3IJuzQrknLKcy9Fvwrl4IFT
w8xtOW5g7zOw8VZcAomCDut642x+RjyLFveSRT3wS3HBbfy4deES1rW+vZM02kG7
Rd+8Sp7bI9eETz3sX19Wvaz3Tm8HgYRRcCDU1qPCn94H4elE4O670J8fsSp3aWLS
2d0ecSm1nB6Var3jixa64nt8EThomp2iWZZ+9GYEivNKUU5fpKdAmuTtf5vo63rz
wTrlAECICxIgVKGL/lrM/Na9Qs663iYRrrRNOMBpukffmhU+gPwylzlBdGNfJ5xj
Z1P5ZTI2kZcegzoI4kGk5a66Ms/r5vVrTmhtRLUV4ZscOXXpHHu0GwUOmkwmook6
T5n8rb/gel5Lhn7Gq1QMjs/o6L376zl5DW/m/Bt6+XUoym4hfZzEIzbsl32+BZhe
HtXZdNDwm51uuDpqgrpcYyj5pzG+F9rQWT8TVbny4hMNwRdud559clR1pj2co8e/
BH+TANGt9EjXt4yNB8CR02n7fAUVW9Je1uyZSzmUB3okfGjyL8gV5iolMC4kveNf
voBhINN3dXbHF+gANc75Evss7fqvE5SnriTxWiXo8j3gCbQxy2m1tIwgCkEm7tRB
4cAtruG46hmz71+ermJcYDTYGkvdJ95x4Qg+Yr0x4mUsvZzn5PeGkpA3ptqcbO8X
4KPWaU0icvh9IS1My1pN84H27CCmnXtrjfcxUaRwMHOa24tL++MoqEYhFP26g7od
ukwwJtl70Ht6TN+NbPdkKkHGL1XIDp8LeoIDLuRgKxgBnSAnAe31ncei57209Fk+
jJR6LWauyCOnTP+FalOxK29E9rIA9U4bKLhVlspaKdrfKU7AqILpF3KcRCQwk26K
Lexs0bFfy9dYZx93KevYzY97KghCgFf+W6w1MgG4OQMeEQXX3vgthREPAGcygDzV
Ye2LZzoC1ACskhQhhR2Ze5MWBv6LsQp0okgaubjr8TgD1ym32m7Vjz3EJZ7ksCgC
wKZSFRyoPNrCQxiF+rqSyF+ZFzubYD8/69Qn3Zs5RpmEMY4XoNrzfB1KUP0F/YJ/
Kiu2+sRFlyrXB3qN74j+EQoz83GvSLf+USvEvwKFbN/2DKHyn6lR+0nrk3tc3+4W
wbfgsnKm5XCVWjP2VAYFLN8Gvc2+AAy+QR6+Rp4KNyS3gWaMX3HksQAyBjENjE80
jMbSyQ1V4051Xzr1YD+ATdGFv5oTFqSX0pGXESxRXJb7BLbwzyrcdSuycX0bBs9v
x9kVlvgJz77zlRGY5RBDfrb0Bf6TRcFzU7cWl45Qf9u1W3gEni0PqdtqB94bdoV1
CcrraSrc3Pm6oaSkQ0aFz8iFWiOGskVc4rADwSF3SqHB4iMzBIt3/xPPcNBhnWOY
GLoh3c78Re0yFSCT13zpbzYOyI59v/r133ss+JCGLHxGMPJKeD2CcZZoJU4TOG86
qLmRGya1RC5mhGZFFDzwUXoqjVmpBxToZP+Ua/f+ikZrsFzwNanHf7MyOOAvYoNb
WlUBbg16UmeazMT8C5JTHG1Wb/J4k5nbY4OFV8hPyTHNQ6skHEqCHHqVBzsUe4Ti
BpZAeolkRKZYuBsdGkomX9wzqaR6/FuLF4X7DJCC3D/6Ps5SPugFjshni1WgKDJU
0ocWXjD1A23bTlmh0YuAbBt1xdgg4h92wjEvscxZEevNqnxOwH9pgX7DY1pdhQDl
AZTYSKjqmewkDLR1FTddSBKk5SPl4UuuCA2fx0OJ/uBC/SQGWZF49mWyRMdtx4Bb
p4mNdLZLGfT0td+srOcWJqJqa/FgMeGUYvswtebaCsiZuv2na0y8SvOn8anrZAJ8
zLkFVvXXwMk+2MHH3l3TL7GN+sj1ICfOVFZnQAfQTp9hwqKHe4OqGZD0OZCRWd6b
dVAQIQXwzzdCAg7sjGatTilogINWam2es9PziIfQqx/PptPKlc8I6GKVy9ILQMw6
TG6Q2iAOMqrKFhhaZhzehfvWcsMh6xSYXsz6Y0617pEydTw5N9ejHNLR7O9P1nrJ
+B05AWc1r4Edo61XZOXae65BotVeuXD2+zziB7IqIEdn+8fFS830qc+VurXMn9Gf
7vRLTZ7bCeE/3h8JEda4dh32JlXLupQ5PeA7kp67VcxnzPlxvPfyfDHeveM9sG/K
apy5WiiK3H5v6z8eBpMJLiK1XcS/JA1R0DSK+Og5tWLfYCn+77Z5jkzf0HejDtbX
k/1RhFOisYVq4Jej7dA/Ex+rzgh6pcsF0XBwOFJ/lS9l49nP38cnEpwXWlGBQb1v
3VytxsJLAJWicXVqwyrj1JcwUUVsjpPepF3a27ebhKF1L2wVxVrf3EW6v7iRxbmT
ulQJcYnP0V/+HvpfxcThFhl5HdqqIixQQJyKDyDNqGutbh25mBt8MePKsbmWGrEn
sQMVt6m7E1o57Mh/6KxYho3InMhiOvYgBSqBHM1xWYmacvdM6OXu+G9dYemlQZr/
ojqHvvkK84eznf9rxh+8v/5yFYmLMYsN5TAXsq6a7a2me72LTOH7D3KB6cPcVSLP
OOA+mkVCqccJbyk6RQj76kCt5xYBZWXmyJcSntf3nK2FayTcJqNLm3Rc4Dj8BT/E
Ks7c73Kz0s3n99Vd+5caQw48x0cVFoawvB0xFAWgr6praG8nfwgN+8t4kk1/xQGI
ECCKY5dYu2bJxGoKlKFZjLHvMnk2/2wr81pZMEz8J1K8YKX15bVppwQOXf9zABQT
+OBoKmoFdEpgeb92L0DXTsI1u7j97fui4iKcIuOjN1AOxL7WX5KA2PiG62KwsRxI
exrKxn8ccggR1wZrgl6Puw9sIHCvrerXxqlUKvjk6Te1jY8aFHt/MeVM7kOnCBb0
y1CY2go4QXathw8tFvjQTlvajjTbbif2iEczvrswZ3bRuX4lA8n3ymXpaaGK16br
ywanYRKMTkN2m2K32QW7gq1kuhnUNkHzwIUiPIRV5DYuctR9PTyWMxGY5ZpwPVvV
20iyWGQNw/wlrmf7h9WEVploAYkZOGwrIYnrx0hpEhBAMR/f+H3eWZh8MpGC57+v
/XGNk4XRJqxrVSkXHFMUs2tkfnIWf6/wEEVPaVFXYarwHjW6lfMl0n88SoIwyAm6
WrOCeKgzMqDAqBE0epsF1KfuHwytqjnHRxQB4s3sk0FYhxILASt9mLCx36zNg0wq
n/+aSHQzzl2aut30pBpvFDq4g4IAD4o+jyKyXcbsRYfXUT604cMyBON07dggWQtz
zCxt4z1+G2JWVglWcaE1/X6cJgi93nw9pgHeV8OMEC7g8fIDVBZjWFzy4q+uLULH
uoXSQLprPdmaA8KX4ft8Xi/FAxF6xpj9mI6z4WAUWO6OsWGe9sepqHxEgXkzdmex
w3AhOwqCjuMQM8vekK16s1j6PlU7F+cWY8SNr4rcXdu/vrWFrhDlOoFuvFGBrKZg
AckKtObzL4TDJeuTCSeQYpOtrxkUnxHJ5RbAWebJiZsyBy6xJ9ulF7D327W0IUrf
OC8/e1ejjE1g/X+c3IZ0L3tgpT6OTROQ+iHItuOo9el/lvoezizAtBsBKzGqm30m
vINeN26MRwgRRyaaSCi07pnS8WFLrf7y2y3kImp5fHcjki8hq4sZqlYH9anHGo8a
EM14WsVUnLf3Xe/PaiRYRQk6lz9k/7XScxpssQ23cmrNifagZGirWaX4VN6OV4FX
95lSV6isJcubjGgfVsOBOIlAtqRpijZJDJ/bgiXF5uLnGVkR/ZsQGEr26zJxuezN
XCGrwpwoUk7l0d5WTxDsjMfDjFhZREBcZfvUk/RZgqQZWlBPpB/+aOWRnUTr8wTk
lgC/TnwnlZtquK01vZ3Z+BJAXPQtgYIZFR6OBBfrZ3c76uF/8CyAZZgCqA0wEAme
QxN4Dkpvl0e4sFtGim10oqtTnsWG8esACKwkszSO7WHcMph4eSiFL2UNijZqiI3O
FVjAlqvPrbjlWJzcAw2URT6l2Zpuj4283zQl/G52F2+LrKOc2KFbujUohF6foEMV
++z+8HutNMGuLjSrvtLD/ZQF+g8qO/tzc2/Tr8UG04fsJtncKzMwVW37pcjdz78P
uvc7xlJn6UV0HweZ7x7FEBq93hEJVO8dpLs1IahzvZqmeJKJaLb6lXJwmr9ePzDN
MZh88y0GELi1i/Q2ylw5idlbFp0VcWrsIQ5BsOElsbwRKNS+TMX3dVZhjg4W3Kvx
zBEdoYHNY7aCmgdiISIZRpi/eClEyO8T1JFlzh7Vn+w7LQYcujRuhHFZW1aYCzJQ
jwi3cewQCUyGuld6IWnwR4Senp+3HDV/PDYIbMTTN4FrZKSkcryLD9dKEn+rYCR7
40z0VYuBXS4JAYBkf6xG7FHQT6BNkBqDPwJ3kX3zePBwAjnbhqnr4GylPzX8r6yW
HsRmrn5CF/sRRowTTHGUTsy4aM8KBg9ULII/f1PnVPWqGu7Xb/+MCyzi51k9AJ4V
7LZkqg0+bfCqpvBB4N/KaNNeIhH8GYsZDV5XIJxl3eCqx4FcHSgSLhtxs3VcZCjw
oL+j7bVTUuqJpLB1pIBt9MAhNv0XmDpn/7SZiwsKXH2yjTJwD3E5lOEOcXrMaNB1
V+UZ8boy9UEyqueybkxUaqm00rv3yW1OjWdFbKKII5fQ4iCJqNzL9NN2VGA4+Yhj
ZnLyvab1S4FvNS21KQqLW1FxQQRSde+v4Ljk8NFcjcWFbF25X6/ngG4BqK63HvVK
mu8bV7g5FkrJl32NoHgIWnI9nwP5YDRkCkMES0H0pp/mN8EO1tXih7W7GT1TJ2P8
GAaaLBnXySnuzLrSeRaCck8yUv8eW7zv72O0n4IWV/BA6oa+ZtSkFeFugNEM0Tst
QePCFndCNnrSeQwg3DoUGBzrNKNM3Q2/u6dEiRakr2Sqi7xztM5azg188VkrEVfp
1RyFFOP/8McVolbBdSiXtq70EsIM86pUGuQECqzY5/oOPH+6IpZpAUDTqJ5mzEO9
pbsnXLRYwUFSdnCVbvHHw6dMrIabwKyCSKJKEANDMD4L628kOKNbJdZlLv4Ft7hE
sBmjMlwKGoU+tJfQa7uXe/YU2iASf4GefQAthaoOx8GZNdoORpTdIS0GX2P3qmwV
JZbfiztr9XsORSSp2yxE9FoVQq1fhNHuN40Dr8wm2q93bdI5BivjJ2SyTe8jNg84
bwwSKTVxYMRPD2gG4McDYAImPwNnPRNJ/NDnSWIXE/V8qHNG2T+QwG9wvjAGcn5S
JzvXP8My3fOUzvU+eBydH2kl2umJSGkOHkFRT+vRYnP3yXMb6cxnDbuA9hiy0Oxs
hup5JzrZ6gLgk/bTjps7PMl/v5tiIJFkaJ8nSl/bLuM8BBbA4/WxayqofFlAYvbn
yapd7DYp7PcAV6qj1JY7mRwNirWkst/VVeWsygu4sI9RkqfOCYKgzeqGJ9uTVr/L
7BRUHpW9xhKQ0l5W5nOU0ODe9VvBIOLfQxT4CVMFMb9pMBNuwMoIubbjIE3YOW9I
UDSOMB2+ciPV0JamcCUKfPCzd8VdGkVQIx/f9LkzXC7eCgBABSDVUh+TMo+7BWsh
yCX6UaeuAxaFkSMRVSyW2y4eFdwuXyHmsSS/NAFAK4GA8pjuPy8SN0Fc++B0mHqL
t46tXjIw5wQVJfxq/iz+8tfS+bmympihHD2JnBo8DRDXLFquJ1+zjRM7yJ/wWUPh
f1XUilIDEVLaAML6PkNvNfurED4q6xfDNKK1H9VGOJh/YGniXRjbD95ZKtEiFYOy
x6R0mE4/7dca5GLKNYImOZKn19qnCfyF/lkkx+dcglRjp6qWMhMmVQGwZUhP3NbI
Mz6YraZEuyKiuF5l9ZfV2Lt7ioINKaMCY045xISdHwmq6grcn2H0blgaqjJj317A
hbjCpCIcAA+5sqWA9u6y5uzAIk8CaIoLMAGx7TpoQU162WO3ebhwUkZSuH82mU3o
fp/L/u9WNZOaNnP1X+R4tv4jUFR35fam3qhCWFDCDo+SNuB9HRvYSKcw7MVq9ozM
QlebJe/j6uUES6tFWmZk5KNgGxAk7jOfOauFVS5pMHaaF/Y+/Iv4mRlz7QI/qiid
ToBh86013S77B6rYfztWykkkKSgR4fknUSlIp+/PcgGnIS+Tu48LT/3YoElOLdgn
mGgXaakj4riYJw/b1H9Btd2Qk2rB31/r/zuc2FLAuMe7bqwzC9C95W7gyWKdQ7jn
8k0xLzFdYN/cVbKVTiv/QRDl4evXKtV3CQpVanztIwsa/8TYTHQWkD2jb58hnmbB
AM8dPsP7WHvdPL7PXzvnE9NDDT5Km1fcd5+JSewkie51UYRulBBAhd1kSRwyhAlm
4lyoFj3HQAWrbkjwJxz6rrvTEs1RXR97OVfc+wSJKtU2UkDXcclPB0lH0rFFUJ2f
Xy/dOuteuhRDcGo2qArZGLf57yjdI2jhnRMCXwRC9ASaTZ2B6rhLVpJ6yXojb4Ym
LEsgxXmC+tVMd9LjV4y4A5Mo8iyaGg1GqAoDGuZFdtRECJaIieU0ozksc1YIDD+A
SvTYrALrKfGQfJ+zeY1BZfFhMbe5R+Ij2Vdd5CLZCGHIRiD2d26QN3jlYH8wgpJp
xBITHW5D4q9ozy2v6TyipnuNgn+oGq40SvLLZTHhzIHfuRETXfG2gvJ/NCa1jRbw
4OldTy8usR9eGrHrGRB+OV2uHKikD49wlNubkJzD/58ejZYseDuGGzO2aaJtqvsg
8bNm5o9z8orgLy145Wdqj+CSVARiBm63M+dHY1OZXR1QiYXS4jqbnT6dFWdRrXVz
bFGpCLYihsrlwumlohslW+E8JnpZRmKh7faDpw4A3pvrUg6wf5HQtiFfulxaai8G
eI9uNuRUw8/MA15bBm99EIUQ0taFUhPtpf2mTh9KDY/7rJjVcUW4NjFE72/jmhYM
bfJGJXnjgrZgIjdhDN7vkvDhaCgMsj4wLo0BCQCGcs2Dp3HW7n9vVAo6XAGQT8oE
ZlacwZCO1oao8TowvS/ONvWZvN/F9xXsZw54Au5Op0hz/4WiYU6JcqdiBmS4IJfT
sX5fDP8/tjqZ6TkhdqgwB81IPVJoy3lMiWE3vfS3FIjAuARhYToBgz2D5B8B1RE1
pEzB7DmpEjoXX0Ojtt1ofVmrYh2oCICBXL6JcAMHeDKwvWgFkI2Vg3J/OIDvWbT6
b/ol6j42B2lIMbLe7J7vr5zcJTa5EcAUau0w5NWPdOyBEfM+JRNwDc6OQqVxgmng
SiqhEsn8ybQdSvfnCVaD4AiVLoJIskAJV0/Ai6kvXU7imxi9sKsX1bwmwPqfROfA
FQrcmb0Dyndi3tfssqmRoU0OCGcqHcfRkFUFFAGufquuLbx+PdYEL4m0+Ugc4avZ
IbvAPd13BbmWEAwVlknYsSTtt14aApIX4q/eFLyuHk7mUyxksGxhkvrvGpAmgvdG
19BzRzP2RripdsyHxPkmDo77dB/NmMRxAnj4a0OdqninpPcNtT2mL2I418sFwQLA
/5Tp7tBc0zANi5Oyh42TQntWqWdpEzenBAUl49eHb9Mp4UYMgAbcS5kxsKxi1PG1
eHT0Gpur8Ud/Xyb/QhdbN6LuCx8KVHJbdep+xRIkAehQq0iCi209CPLogg/zsh5L
mOIQhCg8Lf6UaJ/J52pwXsoG/0WKDmJI1++/K59Qs2yGLEcUpkFWZ2iasQvTvpo3
YlRBwlUKtF4EiB7cg62qJ5te8dUY3qvf29SPvbDF9tIMdmj3OCoV6zDMKEvX//m6
H6X1cRGcS5BvTpXQA2/h2PG/m2lstPDegYbFBedAo0q4AC3Tr9tw/LH1JJ+KEQPn
6CYFc3qy95kDnSEwdjjPaXM0g5SOiM/jdwR15RdVonGZ3aq9+JE1Jd7PQr7TX8rf
uSfOJXTbUfsAQHg4ummEh4u+4gNz/GqH4zovPoSRKMIAGFXd6ttFvToqzloJbNFl
oxAyeB+N6OcQh6p17/x3z61gxFwIhWMjZ4At7Ui2OLm5/tTKXfBKzXarzZ5P+9q1
OhAnNFEn+VHDV8FH2nhZg1lFfS152T2WXCTtmAgBlfL4ATf1AzRKIEyw1N1zZsJR
DeUcNjopAN/Rpwciv8nfAufj9R5byfcoLKhwvVeAovb1h6gLkqwpUpT/Votc1kXe
EM1A/wqL7nr2DLCMMhV1Yd0ko+GzE6ZM3WGFqoIvE+y13wrKVabNEcKJXB6w2L4O
7D5wp+DZ0O0+zs24oJdOD2anj5CqVgJICeg5rgN+2HEpzcTUleqRCmN7B2YhWHW/
SFkIHXRycvGuZsCg2gZ+nmD3EIowlyBIXZ7RRfRsn2znbwoX2oEDCoU3ZYMl2MUu
z1IsI2E64FX6hiEt9gnRyXcgCnqCmwZx9yXE1qnFfsSMFB1oRwKpiUFR5aaZ1ggz
O72JNFyQDb+x8+xk92Kes7j0kG+f9UC8/qdibZ8DmI8HPUoPQlAh/9UXWhXq2gr/
bNO5MtD+ichaJc9pI7zgE/fr4/ytWN88l/VBkLnBs5ky4uXx8+ggExpYxarmmOl+
/kufzXL6o+FU9Vh6QgAVkKojv9c9JFBN7skNafU2oykqpI1Jk0kkAWbZsDsR2RfP
jBKALDOTd26OmA1CmSX8qrf81Glg6FINlj8V3Mh+o+GYbrZqtEg4tihdiqe1/zqP
JghP1J2kx5gWa9/EUmsBb0pABIesIqay4avDva3DfDDz3fuLIP/Pfh072GnXPLPb
rMPuyi0EimgQeL9XV9ryyNy3nYoeNvIIXeus98mldtW0f77E1XDN+Cjdd/brEtSM
T0vOe7EORSE6KNN6dx7aRwXTU7J4GhmCVJ/MN+5Ox9OQ5Pas9itwTIDq9Y77YYFM
CO7JjeNIDlGbTPQi0sWDPVwgGrH0yY6imwtmjGWuQv9pPNQAuvgtwIfboZG/IDzA
ztFV40e/jrRi0CSFpgXV708cLN2u0dMz0zsbI3zmHTpzCrMxWbhXHCYgbyqF3AfR
14L9AMtuwKJql+V5V9pTtKsVfozGb3gJtkSgLAkD0rf/gmplOYOVopxzg809iHIW
nXG/pUI5Wm3NUl3iW/1qwrIGQuCkGmWuk4baWEjtVoOZq+9x9Xhgjhyn2rkv9f7v
2FJgS7VBaR4v5Tk/z2g0pAa4p6CbOuXShbRwcV5loIRY1YdqgscAiuuUj2mh92Ad
s8ei41ao+1xKqYd5+1KPGJINlHHgXFLGVnujTPLhxsEvh6nB9bN/87PnFLd5Hx8M
+KK3Rl63zsoUJU8EMp9s0nk+6ITSZroRJTXRbPcre8PJcfFPsnwHRmciC6YTuRUz
bJmeKOdhSciSpAEuJIPbbUfRw9ue+fc68R1TWDNThvl8W5+DgxQucMuet5HDP4ZS
f24i2m46q0Lb1LSz2FeO2rcBfb+VvpX3vD/WrRDPWG3hxPdMKwPE8CEsjSNVGvrp
TXtPG0Gg5+HAePTMeRJzA/fbkYlMfsAUoz9phLBCeGkbq/YbGaur4vTNTxXQZS8U
qpyzk5t+aLvH6UqtaIB9Isu4a4C2RL5PG9/hhCVSXaQJw5ODuFrZjfxBJabMuwvV
V2v0yK1AxcXyc3k/uCCkw/udRSTmmY3c3IDskKldjM5UMNkLCRk2/aaKYdw0edZO
DbcPiA17vr16bVZXI8iXU2IGsyuiPBKqTZ3GNcTidBLNa4gYKbkxJOmnEivFmhh/
lydkS/b+J9GEQvtH4w3MDuY9slhymKYhmgyGr2DMf3JrLdo+HcswkhgbW4lOQSdp
qwes6BkEApBdS8+HkNhvWNQ/A50qg8h0JAC7CBTMVOYRsW/3Jgo+ysOJo5WGHbp9
ibmYE7vysVREra3yDD2Un3cMh+nzKPjvOOUeHVPmsktRFXoBbL4Hbi58NT8MGh6Z
E+glO2xTw//fDhiCfk3bmATzdw3wolDLm81qtRgOO17SICPiVqZ4QMMAD9XhCgB7
VRslk5HNmpr8yeG7+y1Tj/Ml782uCRnJn+/EpOc6oi81TNuphE7Ti/5hatARlxjo
3GPFq4ll+IoDEC71b8lpK6MoWbcWxkS8TJmnPLlnJrzeApXFbbpZKYmS49+AcG8C
8bPz6L8mc3J0F2yy9Vj2iCDYelo4Nsl/jmyZyyJm2DxoRRhaaYL7B6VfHbUJ4Ywx
FHVHkEu97g9OT4BwCozSydZDFyua2bhFz4gpUWWHupnojD94fxNhcPjHhqNb9Ja+
LA/uJr/oFaIb2rSLJ+SrIgaOkLBJ/83h4q/pWUeP2R/QwZ4zLUnRkEcFhIdQFxoT
fPz5WSZLIxS9dwnG8kvk4re1Ru/WltbtlBY3m8Rhr6bEAuD975SNQAyWy43ijXHE
i42e8yYUwjQNVR16Ha4oShR4U/MTUsKTtEN7z79Ti37isFJN2FeQv5Wz9DNqeHqy
Ah87cGffuJqdFlK3dRmDJXBny7ltUbDuT+brqaiRGnMdGBZFhJY5kdfMfoypjGpE
KFhKzWZ9otuE5fEj4eLN37YyjPTMawnHft03qk1GqBk0iHTqRsanzMrvPQ7mhWPR
i+zPnSlXNgR5msKMqlQ+aUTuqjVV9d7vyrL+sUm4DB5H8/UJFvLCfntASFgP/PFg
6UMcwhMdG9scT1fk2p1OdgjVGq2wxheikyLVtaWmK/3U0ggT2tm615O8Z+88JI9Y
qGrpB07Sph6OTbPZ5ei5gAFDl7lCCh+AzrLe77P1fSNMJ/pGe0JAw9tu+4ZsMtMB
W0cSzKejLfwkx1cSMVQRbOls3c3h0tJy5APHiDd2LOLBFe6alI3IT99DkgnE4rgO
Vrg9KFPgUs8lx1FsxFCK3DMbi9sIzhp2RCBiSxRZJB6k65XK0u58TetXWxiuOkKs
NYn4gncZ3ZuecRGckky1SfAqPgyhZ7q9TRe6xVFfJwHkfIb98MIVts4AydaIInHg
Zx4Ijdp14x6V/czZb/gWVRzk63hKSJyFnMtGBYG9bBDnBT/E2VNHBbevBomDBZYX
yUmvv3tTlKdxcY9L4I8seebiuFbgG4DWSXfkRXuN/dQ3HsmetbiDZ7E2mGfmpcP0
zy0z1h5s63H2+5bTFFWIfKxq/i0h+rXwDhXqV4uLR0USP/a8aam+CUmv9c9Gy8+t
yHgduvM8cPTEFWcYXWjYO/L3HeJOhfJwBF0G0TxtfdMsc5/CgPP+kql3PeLosZ69
scf2+4jhD0IKB6NDnGNxN66I4b2tbQW9f1JR+MSU8ADd9Mn9PPlZvbrRXI6O59RG
RThs9gIO9ZdLCneNblnAxo6YQcY6qddWBbZmrCrDOMtfaC9COCDCJhkphoDK7ZwO
9cMZDQ7e3H4t19eVoYdiHeffntwwPfESPRVYGbC05TY+vStSOTY9KscjzNpsz0Ou
4aVICxm3hJ6TRtiiePYA0AyemELLsWeUdvzUvEsLhVosSapRja5B3Hi47IYp7Loi
x8pPOboU4x6KQyVS+lSKA5JvfB+1hGR/3lWDM8xTY0IxlVT/dXMxzQrag7L5WtPP
j9U2XVyujiTdTEg3CIjtnryug9vNnoBKSfX+yCCFO80MJsPZv9JrxYO3Z1Uwrq0k
HumFPTpDtgYvTz3c6JiHeCZ1l4ybneXIEtH0sCO9lqYQLkuTPHNa05YyrYUYPLST
Pm0m+NITczuSZa0M5lV/qmWBbFNKQq4ECwiI32L6QM0NE/aVDWkVWrBCOHYrmjOf
8OP6Py2/eEPLVZNuVwbe2YQgg/M/Z0/4tnL2lfCesNzbXTf7JJQ6xXTTyEdIDpWG
TW3H1ljp9LqK/Fbxjqszv5c3eJ7GEqjsL3mafpfCIzZYgHJYSeOuYCIfc6KNC9NA
PQWQFN1je++7WQ4qw7CbXBNL2Ks61vK71XAidjJeGM5uGST9v0/bUEO+H6ASmauI
rh9ElGfbgC7+tojHtkOMDGXqiXtOtQpdhPaGlxH+DaRh1W/OruA33bTr5t46i3MM
MW4nGpf97S17aoUTqjNnzHlGgpIHWmJcgi5Kfo245CuLSc1bx/1tslsMgO31Xp+Z
YQe+cIuxkJpMqCatWHqpySldZAbVqfdBh/jaHSylk2dlbw+ZejqvatSLOE0iV7sw
TXVBkD/kk6Jii1DVl/6+hAku+yjSXLV/ZnQoZjjqNprk/xDOXpVg+LlUwzQKb15I
MekksZGJKPjVbera2ioOB8nusXx6RYWvowbg9M91ouavImkGWRs7GLl6cCCxMXTm
tcIovd7IH4up8gR2Rearp3YS+1l4nOh2ziDPntqKUuxoQdAJKLT5244fA7YGR9g6
5gQxTDHx38li4sWfixfMmb0PJLALiwPCMQJAuL81Ggz9IVHq0QUyeNFfI9LFq71T
cCczfKCWZq/ce5O+odw1An8Atn1BM0kM0XkPtKPzqNge5/1pD7zKfOuc+dgQHvxM
iF5YHyCTG1LiRHh0cKOVBhRjZb0XWMtcEs88OiHY3db4pTeSmaeTBogAOUFIel9b
SsyXxQoiSp+CV+bG7GKplWfC/AIngVBqDSnEr9kQMoIB59UlwEtIWsdmDVXOZaPw
z3cR5e8yF5JwIZVs0QiSUAyKqhrJN4gMmq/gdHIESitZbYHC+wi+249TxNhZRrnG
B9aIWZ4YnXjvD0pQQTZfQZpOeonS1yk+On7zYJDJlLpmgeecGukveSzRgD1egVEG
rf7BPllUYoePJGNB3Iabc0rRzSZZCIz0uRPKbLQ1x7EEcn3sPcpYuWU59z+VKxcm
tiND97igWOEkPrhLWolpBhVYeYzdnVzo2t5TK1sovUrml3fto+3OlGv3ELG6Ppv5
P8oeYdeAl0sWWVugmWONiSGWki1POMgfN9ALv+mu+SZwXz6SeM6Ba9+jSIskgw75
NIl1W6S4oATgAg2MON9dPrKbL/bzcRdbQkg0evsE06LADmNkVYY58HilH5NRrzkp
g5S8Dx5rEq5TJHdVh/1JPAnAV2xOeoX1SFtHJkWpTS4QpGS+KFVgqXdLp5yR2Cb6
spYPQS3v6Hp1qk4+9Flhxix/hZj476il07RpjKvLrhAlZ752h3T9ggtuVmxBr9/K
gu6GMoBC02XT8rDcUPM4Y99EoeIzmoqOjzkpQbIXjLCJcNDc1sEwAtVomHTzjYoc
dpA3woE481MkOsq0FqT6h6ua8lTzOBV/3u6cPX48YQKmT7qaT1gC+F+p3/wIk+vi
3FiGr38WExfwrRPpDlwDmk5Wf9eQ2LW6aUYRlckXdrNhUL3EtXVLRiZh8rTysmZ3
yvWGHugfXa7nGyt2vkO7s7JzQhf++WZFO0NQzVtv0GTCxOGX+tmYOYc5gxlK6vjS
g57Nz7gPObL8zHI5BABw8pGjyHKGA1xmjWNMfokz7ymLE21ohG579Kh4EIo4FKrf
zNtuTLaR39B2sF3Qezpn7RhdR65tXiIIA4dzWfIsJ0nuyBNbgkmeJ8hlZ/e7q/Yz
YGCnblEg8VNiI+1uABT1iw7cNOT7ZfwvfgwDZWscJyMlnLKYQvKshbt9mbmo24I5
p0puAfZZRccCi3LX8JHjzIRbKneLw3eOWqjJEiWm3c1hPgWziJIQfskUXF4labii
3QDxk7dfJk+yEkV8pOx6+9Ioq+loIvUarmJ7cHwtViX/Fa7R7jb8oSTBB53md/yw
6xJ3ijupVz0qQx6v+/U61olvR8of5HQAt5zrA0doHOEF0seo7zpqrCIBT3oXyoMf
sNWOrc5RU6I5leaDsGcAZg8G+rt0q3UW7cuGtoSmcmwua/qhsevZISlxFhYxbvJw
gn5BJ/2X1UkxLWigluMMnhBtEAFx9gyuLtLTDj8pvkrZ4KtoRwcyr5BV/2SkWVy8
mXenOoSwfiqsJrwrSxk9QvzCq9Plf0RzLDZfpxQJLYzb1slw352QxClK7tYe+y+Y
m6Q/HyqOToDTSNPAjr0snjqBaPphKlKOC8J9mAwpxdMImPvKvT6FcgpXxDxFv4L0
Rv3PuBZR5MY51dfQADZqtKAYklfLIXcBxXxSXeDwRwChVhcgkdhwhVWY0lMW7u9q
RE3wAdIsYith5qzTPY/3Il843e98yRb/RAx3z9v1ImA2XUgQEu/kozqHxTGddoDK
GKbfITOK8n5brxyFSFAdMsEfUWSKikasVKfal0TYfZaI//EeH6teNLJLEGbQp4xB
0xr5aIHeBFj3U8vgFWQ2OtTlyYQIWnwWhi9LYQxcWuCEnd0DZNB+HuIZkhM65Pzu
sl/btT/AksP5eEnEar38rdpva4RcAwB+mcMo96f9jPaX4djOhh/hjxdi54owuUlB
kAwVwr3k/sVJi7WrYs6Dklah2gunF5iLa1sxZQUsbJx37/MuB3EuQSQQdEYdN3ba
gRrNNlMCuVT3AI/T2Vc5PSxXd8+s2KiKsDXF1tNaDsvuegwQYA/miPMNyIKP9TvD
mcoSbNCClnn36LuLupGfmqt1nxfRBLj/jnSFZoK/LJv5yYEHHf5WBnu4zb/MWjlL
zicHNaDujiV8kM+VNwiAoYL5ZvEM8rLxE1eVxJN4nmYu19ZSABdtRqBexWellCh7
dQ7nBPqL2Ww54YEO4ZpcLNWq3uy5JAnruxyTbu63ZXGP4K3vv5nG5tjdlQtpZLWK
SUGhNcV7NzwmicUVwJMwlgu5hgswBOTQm0rkOdqUnHTg3BP3Xvlb2V4VfTntAtQ+
2pFFlPUt00s328U0qzI8apcHI5JhTnGH1stOgFC/gtra5J39JBUePaxWI+2eQJvC
KIVsgX9JwufpyDIWxvF1jpZPzbqt0hyGNgggazLA8HqeF3siEfjKcEfDCVc2sB6y
Z7N/HUO0xuFNfPbsINkU5rQB15D594uGuqKM73g84e2uIKIQ3UA8m1oL5/WI+PXJ
LOC848Ok7lTOTO7MV7XIx3r4SjS9J+Q2hE8suaal3mGsuXq5TIrxT/FoiN2UIRJv
x+jv1X0dhBIw20qEkj0+2ay+rH9p8jJxxyPnq0I7Q0QAsQtZE+3Zh1cU2ZPS7wGz
hi1TuXv4Tz0pjxowa55D7RQzgtk8d2xdpC54ixOXbn9IbNHVJfSoxaHQBQtq+8+5
CbPPoq6Wiebx2TgRTA9VKNnvrQUuJTA+47C7p8ImioQiFqr/i+SDZWZTRt8AQAfp
0n1crmHwOym/yvQgx/XjNkB2fh20uzgMhTMZpVrshHvAHdt5QpI7wyZs7WyYnjbQ
r6b0jDP3NquDXff6VsRagfDkN/blNxh/saY3HCsfQir6jWgsMkjZdI9hVhdGGWyJ
W9zuxzI//e+ASegA4/vq5UqKO1KXPUaDL3vLU9fwAnZH57zsMt24A1OEG2TYeq/6
kaO98gZsosePo7uCefJJ6UiGliMSC6cxr0S1aCPN1k4a1pmr7W9G43E6jHqZlgEM
R5eFpKccuxbrYkqyAtwGSzIjSEwUYgI8WkkzTDx4hsZNn2jvO8oXjH/tDm5TnMi9
sVoCqsENcz7Yb9FuQZ9WkY+ga4ZBavDuhzvM0faVILVAh9Pi0sE7e90aggT1Ys+m
2PtAVg1JpGSfTrgafv07vzpHu6WkIBl+jg5jmzRDAIjd+PVSTRnPYY94uLWyMCy1
VrVwUg6MqbFWksHde9cgGRhn8mrBwuIf73ddkkIGhAVCPNEfqNVfcFXGqBG3n/Op
+w9i1ndCPsv3SqZPFp4NDWecbwewfXbERXcQ9V2SDD7W/Jv2YizLIAbw7v2OjKRh
KltoAkmAylDSVWjU8S7qX11p+sY3g7Y/cUqYidu7AdG203oCLXTS1Zn07M4EPpft
j9nODSf6UDzrzX5H/2bz2oKd7t5AUy3mA/JsLIc9RnBw92mVYJBGVFQPF/lm9i1n
htEKl18xZiZYSvyA9LsjQK/nm3PCBLTnmfw/W3tgC3z0pK67N1+QO34rlePgOj+R
9AB4oFXL0WZ0ZIahe+tP+aWvn8fFoNgM6Jgf+2pbJGvJh0TbSDV3O1gFYvtexRPD
1Qh0u2ONcjBMjNTIn/8oD44gL8D6WcWc6pOpgFHHpe0on5B158J0dVV86IqFFIv+
9MVDAD+MivH4EKyiY8o7fSmku2/k3Jis4mAfZ7T88PbUdyKvqQSHwJ0MmEg4O2/W
43cP3h5d3dEdjNS46+JdET05yChY9sT1AS+bicdcSSAsAXiz+IffsJiEtohK0bLK
ROaLORk2xbXO3X9iZHzQtRfpMQVQftIhIS6bw7/lF6dvArwfBU3mkcZJP8CdQ2yU
yxMZCvGs9uDmUXoMoKNCPbIOxXhvBLpYTaG4oeLBhbTC1Vf49YWt//hhb04acBQu
Ee0ZrLaUTgNGpYBI4dndiRtCpP6h4I4bpe05FC6/0QcTf2l+d3kABQSbwev2vi+j
lweBIycUPH6HM+eLDJs1JVoCSzE3QB9Wa4bn4jTAQG6NF8q+FlMKJ8/v7mencQq6
LcXYjGbyPm66nc5xmaNXgDo0HkMfqyD07k34Ab9JnsFsVA3C2QnvFUYApjqXL9yh
jwnerqwSSCPuSPWlPYnanqtb09VZhPPIMpoi05FaDRa9Xw0eAGKjm3dA4IBlFph6
doRc5DsdmUEqxy8n0scYH9W4muJZWUGFx+MwncgL3dx59cBWG0n0A8mw8jBN/lll
2czM4zaEPzF2CKKMxf8/mdKJQdNVEXIFg6L6bocHxIPs23g1xmOEIH+e7KP4O+3h
+UJVKOCPiRr9dDIkI8GXCWurI5VegwLU+hbGCAVMiTKCjSCCehplsxJzUmGa70pc
eaIpwB8JJV/C80kjCdVwKqiru0cZ8jMJy1+JW57eGkGZIJplz5ThQURrxungoYNd
U358ZUwfnLfuJtW25HnmuhG2/9bYojZTiUbJaC4UT0GnYgA7tgnIvKCXGd221w83
K4m3SM/rdfkKf+Ku/9HQuShVOdM9mWKa6vfo7k3jc6GyuIqZkGYljHbdpG1ZhKcJ
IuQ5pdSw3rXaiWdXY13zanEZwE3cWZigaypPaaCYKVWjr6pWeQiVO9vJXkMFwubK
DpPxseQWl7sWBrTmYrLb7FvVz8esHqvA/nlQS55aI0y8nBmpnFzTBAEpdsnwpghG
10de6y57qhN8qDAd1FSvEBCrM8Lk3TtHyR4pVo/t68rywKsSHgnZ1hQ/8XGz1o8W
mCj5Dr4g28lIcXTKtzN9BI5nh5hEthiBcehbeWk8qervQCM5Bng1MD9hJVuOKkdX
UiLweuCVCOIriRFF5b3O6z/BnC4U6PkYX9iPJ29y1sUaDo8Gyld+nyX7rMFdfRVn
yv6IhtHMnPtblVS+iD4YW9ygcJCAUP8oPaBicoh+MTxQyAZ6mlq3g2CU/ooz8JGR
zy1rIR//zM7QHzPzKX06Uyvv1FmuT8th+is+xoDmEI/9mLiOj8hQmdQM9fYKXDS9
4GMBNaFjQ1XoWsnDVL+ETX2wYJeQcmHiQnm8e2lbpF/3jEeW/mXuKlvBpPI4SrUf
DfjrYQui5lH5ZxWqfINm10JlUAhF1pI06f2m0BTy1O9WaeKkpkxq6Qdx5OrEup1J
E9KAnhXRx5YohRa5hw+ADIL3W/Bj6d+KZQZ8k+F07MHEiRMqPDAbLg/RlexiyqEd
S/R2qatknKYe47smt2hY29cgmNBZk683WJ6txvKKLSfIEB0KwaQcnyilWunAPhX5
DGmO+f74vaycKPQLmuxYIvQ4H4ysgf/67YBMGDk9jJFFUZxxQT+CK7EaD3NOP4HL
spMv2CT+9HpSTeDBxrguOCv76LE8o1Gf6VojN1V8QGqyMY2ZgzUDjIBXS3fhvVhZ
vB2Bi6rXRLJzeTYENgW02QxcRNNZS3WNr8AJdhb8/ZJD5OO13hqNTSlC88Oo/L0O
JljfuK0uL1z3danloK+05rx7ovvMXF7ecMLzYBcphQXI3MEweSaA8Jur1XsTACFI
KechkqYOezbl+j//ZeN5uS5z9ksQ8k4fJ4Lb8oGagSCY5gs+RXWQ0f/z0zT08j06
hgqatRA9fkB473w2o6L6QWE6IgDnwyXzDcQtThBynQTq3bFgM45fEghi3uMir4m9
dB7B/I/Ti40X8/WGwlZ4mQ0wpF4SirtS88rGxDmlLRTApTYFDtD1sgnqnzKnIbcO
HZUsRYR7zceFpHxpUiguA8C3KhdaOKk0KMMKep1lzUyq8V2vne+GEg/cwMp2MoMj
L6TAn+pi05IHERtPSglCc4mLVIyC8C0ucoJayIZNBhpoqZ8iq28oobKJJVRAN+nr
90laJXDyLmaxhBVyy+jNhlXAa9LV6PEFX4oBXqV8aYOrSRNUZk8J0jjhsMtk0Ne+
43wM0d/DkfsTyt/WLq1Xv2cDG2tuetqbt68Ne9iNAtViUX7hSiLD8wUpWy7e9nwF
zKPzcOG06Rfl/imyjH0OpwzOtbMKlJBsStJ6vDzRXdi4y8OxUOZBB8z5o6NjxApL
FaJMd7f98tG7b55ufDiNp3D9ed2lSc8Lo8QTQwJ7KTAChpvv4u1F3u2d4eFxw/Ph
BWqHEIcAKHzeuc9o0Ug1gUBFdllYKzw+mVtneutM5oUXAmGjgNDPHNn9/q70uMoj
Vv4/3pXROQXvdY6asWpw1BmJD+2gxyuT7nbhPJG11Us/h9i1kVtAeEU7uPocFoa8
aU6KSyc2UZHcMoOt/4N9kOG+EiQoKjm0SA7GF0Q+nnec9E8Or+BAEjhVG1kX8IWK
uubHdB/yFIZiG2XNCIBsAf6btQ2M/nPviK819OHcFKDt2W10Du/+v8+3QoFsUwan
XmaZI5K7UBEJg4bzk7RD3wLiAExkxk2Hbs/4J7su8GT1UXhOsOd0mVUwKOwQMHQJ
Szl9/T3SeoZkarr22tyJjzSWFmpM8JiXSnX1ccY4v7TqqN6CARdWeiTkvdy+A+wf
POoc1mSzY4KpRfwTwEMw1miopA8xbVadJq6rsPS7xpR4djSYVm6ojf0/QgrBcpew
MFR4l0hh3h9I3Wm22cje7MT1djuu5/tVs/pWe/zO7JqzRJ65SHoG/XG7FpkRJNJ4
PAnfVMAbPJqmbNp/Wth3PYjk1WhXsZBqOxVOTbJS8m1oQvxak/4V4VecLGyhz3Uq
iLsxNbxnWbLa6ooii98sBh/CxgpmgN5l780WSST7bU0etG/9/1UsDWmX1bpT+qNB
TGNnWnjZ4s9+YESEg5vZHv6T2whzv9bNCCiEPmskgIxAQGnDRvipP+ZSLJabAKIW
5OepVvv3e0BU00SDjrDnVFOK+yOL72kn0z4uaduoMkTQGilWUnfE5fpWJ1svTD6t
OQWB2icVYzmO/np7bjKh/eqrR/77qMgmUhbA39U10Rn/xpV4z4OP00aubCoFwZEe
GLfMUJHmoeW1554Xy0VyltR6wMH5lpjkYtFiSmv8vlHSwhITAPJ7oBoizVT9SBYw
/q2yEAyKPpjNwd761px4z+EyUsXjFa3+oHva6k4FYxJ1Sahj4/ddFOSaYGCNNSiU
Zpci6uaLAg5Kh6buOuGsblddWdSW43uCrJEwvV3T2rQm2TBDZ0j7VhPwYwjU1iBe
TB2FX9L5UK+GqFf5XWWC3aP18nRgaooi5pMV1AWV+ljOV6+U7VV06PYNo5TudCFv
9eOet0QcA+KF/cHY/VfhuzbsxImGK7i7h56YM7oQA7s3OrtyK5mm3CCozcpPsLSd
UcYtrr4hKXVBDOr5tKmFzNR6iUkpGpsq4Imfd2aZIZOJS78jEg3au6+TUjEeXsDI
F1uwjmlGzWewA63He9VV0J9PgOeJsDsa3JVCstVrQ3VeXjjbNIhRyUnVsMWRYGxF
FqKzanNkUdwA47VBSpRSIGD6Okh1Dwb9rcw83hAQ755k3EA5ewSEbXMEPWt3hzJP
bLD1wJrFkfdmH4fK6N7FijVQ/iJEyZxDU/YNe968KJ4poDyesqoEEh+5pglRhV5o
iwRXiWE+/7FoxFloXgo0VLRKoTb7YYcP9no02Y9X9U3wgSRJbtTz87uxmcvo9Sbx
TtwWihbh3wnWi43dzgD8JaI1UMGzQpBvcTCPEKA62SbbxK2Isn7a5DgI8B+/J5CW
S5zX+q6AsDllMvoYfVAlj4r/s7XUZSwqAAHVlU/C8x+Wb77QNPXqVyduYAQbPgyD
I073tlcTZI73n12uyyQowYIqBJMptV/NHcON8MjpsGN/CU7fV7WhFqjOO4pGx9VN
NzZOXdm7SPrFBYvLKtLQeqKChgp/UraMRfEJTD+1o64AzuqOfNChJL7Q+wBSzUV8
NCDdcno6itnVJ/gQ3UpknJvxjk15LTqY5X9ZxzEw8iggqxD9f626mAYI7XUMjJsj
2XqjBQtJFb9lcU/8Hv30kDNqk4tgyNUqQYlNZn7f0Vu+06YXZ0frGLju5K2Vkr7U
gEdqGXeXELlcFvfNLmal2Zm+lJGBDKxXX3isw0Uhiq1uozr+ra/qk7gd5c/lziEp
9u09UmFv3O4ZoPSu3CUc+lUSbMlBwzPKPGHrXahMYXnGnKyjwtBxw0nAM823J5VB
FmbgmcjPMbb5Ca+Urz00KCFvNNniSu1quVAMz/ddOXF/XvUxm7qSuT6YoCquUpiT
UJUaGnkK+J2xLZR8uCZz04T2g6HY9AnEwVDWgULtnrri9ass6dRQJATX/vO8vzoI
Tm9PRaLPawclkLvy2nfwA6QqVVj3qAm6ZxV5iD8r6uRrIaGS+ZYsRC4Lk9clZH7Q
QCXgoR7d/fdffTFa2RmfKGzEZmPE22HeSCKD7sIdTF3BDXbSr6r6rus7Sfb843yY
OcmrJz/MYzjeufEQWAR5vKthehYDsmv8QKiPUhiBD2gOJ4vACR6bJ5/nfQeQ7T1R
Mq1hRzUhQ8tc/v+uM6e29GXF54/NBL+bFSnP1ZyI1VVbaDgtuCuapW/A7JKIn0Sk
1LTyTe3DYqyzxaEwB97XDDKKnpQ3azDJkuwVME6doiFG7xxJOkVP8BpmL9gXzuMB
byB9Ty9KQOdCWVNbLbROnJJBmMwt5qWjpm6AcKngozXJ+6gZwlJ4EixokaFAnG9g
qlMpRJ0GMqh5IbdVSeyBViZ4nJne2MrHkB2phTZi687Vwz7IsDBwp7KqD3dUhJQ5
RCQDQcP9LUuz+moRGpcsRbj2yN+X9wztftGkxyvTZ6QDoLlu0DVu7C6a0XMuwU1J
Bq7TAivs3mhicWCxU9nF/U2FWeXxYVJabkYIT4SteEb6rKpAOmVk5iYkOk3borEu
CAlzQD/ZPIdKju6TgLtd30CTx/DNCmoVSKyiUV2mZ2rpBJnk11D7Qd8AYh8IlmKc
vDOK+OeUgtIndZxB8ux2P/hFnlemxoKTZxPLNARLFvpZ2NfXFbe4DtlfU6E23o4n
5pkwf/Y4e4i2oSQrVAFf6/PZrpLF0FkpENwTNTDece1eSDvt0GBUCeuu40P5GehM
pfqfzzXVf8HBvk+8/klPKJFrkFA3X5DVfHa9QcoM5xf4pO8sGAdaL4fe88GY76Zg
WACyNPiodsjcvl6yUzF9wbnJoU1ug+NH72XLqVy0jxuMGJ9V3bmyi1GzprJZWOm9
fhmGVJuQfCptPeBAP7B1oriiHMLOzXCDWmF3QM5lsJt9Yr2TZosbHtZE1Z9DJXu+
tShqU4ecrWWQ0P8UKj2iFNBWRhMZl6CbK42FR4mb/PqcgAwV4i7dPdQFyjgm09nr
aNImYeJhCaFo5nHmEqCbTuHa+5NhFlbzYCVe5OJQ8LLyaaFFEqqpexmGIp3tmVss
FRAjjsLa5G1cX+pQNf4GzPkctZXRLe8AKxBHPAZFhAOBfYpzSij496l0JqVd0JTn
mMZDWY1UdwgfanfVX51sJi5oeg8JWVAP7ZPXfOkM2dktgC9p3vhvPCMV5aQVqhLs
R1sLvn5FgrJS9zMdUhFE+qewvuMTn8k0xtRxoeiYwKvOrsjXKarAInNGpJo3DnUd
kuHCqVY1A+RSx/kTigyXN1SDaYcY2Az3hyH71zAav9BVJ/dK0+adv9ObAdO0MKco
zbXEFeUba7jRYPYqcf21coBC0qh4dwOxgZBHsMAe/Vh2rcI2J6RBVravZzgD4vYx
CgM8/rWhhrubMTGCrH+qqJwICbrpo0W1Og2BmjzdpVF2pk3Y8lqe09pT9UszZ4xk
6aACxvI/piq5oDQpFKvpX/+L4tDBknGo3ypdH2mR5JSww2bLJ9UkRJlcEeguwzNk
JpFFnaHrH4rXgj5FoWQyk99DonTtAbfq2+M/LiJSx+tAJVzDxh1QqtUBWuCHo0uu
+KN/K2qmwbOftwSaFq6kIOkP9b2Gnwqnj8aVQjPgeoctUZ2GTUzotjQtXK2LsgiV
lzJnlGdjfJ3bA5T8hjKUW4gGE3R4rkPiH5NJtJIztItvzllmMaoKj7YIPRqSNEVB
rj3JXTDY7CMh/hQcKYuhANEfDBStyYxAKwrUrotuAxQtIagWJLfU+9AYvMuxp3Tf
32UevsI0DvPte4MmAFUo2Kkw4Ky067rJ2E0RgWZSC5Fen058FT7ApiTwogkbMt+z
4APKu8DDSxz8ELVtWC4ZBEK6/C7eol9Z+FTZxqn9kr72XomQ4aCA27q2N9dMgOIL
esbLAct7PRqFkq+ci0JKLPGFQhZUsihrv7QDysJL9NjVBHttvCDGSm4Bvx5elYyl
fmFu8sqaYUVBtxdAY4kUKuTf8FK2x2lDHts8V9C1fCWqEbY7AltW9guvL2pjm+Qr
NySRFtsQ0p9GHbhOdaz5GpWl0oQx1Dbc3b6wyozoCjLU0e/4/4I7L3KS4fKUnvTO
AWtwP4yn5IlXOyJwaAXNvEo/KJghsSDO9mmSslqlXwsNiDoEWfReaIoFwG94gNng
VlfT5AlRU06g65QUeks4ndJuzKVvpkhWuti+FmmQAHOi+lLdoidq3SxrqQ1Ks3vo
zTJHoZrWvEZzlRCgGwSNsctjVhjM08P48fvFunbFIxCQokYMRCOtMmn9+IfKbbVW
aUvsIb1zcpcohu/NCHqT9S6jXJpB55JJBoamNGRm+4moclkG0s06pxaSF87KBz+4
Rq4Dh8NrQ6Gqf9OuPp1koOHOq9Py6zBZbEHAEZXrV/ESiMzMjhFJ+sG6Y2fbWfl3
eJHVGd+DkMd5J0CpYgfpFdpNqqmOba5g6h5AfpmHMQpS7qJNLe6GDt0nYPKIfKWF
7uNrly92lfRjDR8PjQoZrv6b0FYX46YND4zStVSmzbdflXSkTSZG2BhsgEw5qW2D
NNrv5XnoJysTBACaMOOBCFfsYk+tUcgxuFZwk83CiaxYgwJ3yY/oB96BhpQr+Yib
dTRyZbT3GYrSzP9t+xHYms7zatPtJ6S7ZW6OmuxS0ko/hY2kibPrLzqMxgmSJRgZ
Sfy5S5KWmidKKd0o/FYD8MVg9yzzzBmwmhQO+HEy9fAZTceeQ+WTywR9kL6QwW3P
sZ8QQqMj8rWllMAE7OgVSUfGbxP1OViwo7D4QAJhajL1iizZHXWsXK0j7lIHvIeA
mFeCsVBnJwnTBcrGZNwCSl66YmH5dpQwsJlw/ZDErG5v7nxFwUlNRUTdFCzhFGmx
7Yvs3hxiHD11XbWRRWsZjES+3zmFqaOuXqXaF5XnRJYtC4T+mWXYsAoCJj9Y4tqP
gzZc9UMs42RRtPS85XlnhpDnCHWm+DmREBlAH0Z9K9iIPnC63t3CyqSIWVtv0rMz
+7yi6cqbMUoAmB19BIAY5/vtFcyzVNe8afBokBiorhWK556rnPJqoTAWbTIz4Jt6
F+FDG0yX9MuEgOUvQ3TKpLcmWYyaY1pvcfhpQNUBSLcO8yQUI9blq0qqpHcW+cau
nCNeBbbGhP9SyU0h2Iy1uLjY2v0OCY98b0vcW6D9rGdpvYO8NKFYdm4GDDrKupPy
MjLtK+fwprMZE3CuNlelq0QC9Lm5jLSkuhf5RPL4Ur5oHhOD+mhsXVmB6to3s1v9
tDwZeHDMKbC/KglvMx1IyjzluYipOhWiiWLmIyzxB78TKabiHZM7SST6lrFuhCFn
4NLwxXxM+Tlspx6s+DxSfFgtmuZQ+dI5igjVmer9vyT2XMzGXfXAaTtowdrzn0VY
NuUpg6ahgccD1sO3MJtmGJgWqaFWIQckIe1+0NZXeLWGYuKUWqzXlW91yL8Jf88Q
06KeWOS1tlEOpLlFD9MagSIZom9NxO+Qn5BVyWvtNZByIAwmuk6jweyhenZdjXGn
ZXCBP361g+m89UNwiNtd665iXO5QVoGzIVwjaWRpM6N2oOCW/+/8+4veyqqkm0Af
gzRVq9Rq2nLR+fFEDhq6VXnVQTShZfqcNOplG3zoC0Z6GRPGtGasrcuGrLnpnssv
mHLqIfegJ1GsSCsmcQAYmkcoaB5ANIEC5kUXsmkyvx9tZ5UtBQyCaXXGV5vOgzNI
ykkE3TJRyd+u7uF8B2InybXJQUsEl7UAVxIyF1kwgmgQBf72yKY7NHwSLrgUnlwg
6WB+ckXHFfcPLeq3D47XVE3s5WRYw3CY+00TW0TlmRj3dEWO7VIPG+YmKPb5o79C
IKmjj71m4xYBsKI7i42HKH2bbUlhx508ne7jhlqLLKtnjIPljP2kPcistqBRc0Ly
wqKHI2g/Bbu4QdNNBavUsWpkdRpiZLQ+vkT1Ndr2nz7dwD5Y0tumYCNdgNfMKkt2
06HbxJyVS3H8OcwmhJh7DUxIjc3SwM5+L1g4pjidyJIFyk2ZL7A6a1NlwCDbxS4f
mosBZIHt2nHgEstDA2QD6/CNljpPKib9L2odwZEyGUhHHdVa2vSYRG0JWAKtwYeT
gZYzFThQtdQoGokz4btH1m9wThebvBBC7DedlZpZ8Tu99KFNvzSYrBLWmdW+Zmnu
wk8cyFMwBjBACpGt9Ju2TKVCDEi+CkzHw9jt4aQpE5kLfYLTya7s0Z4nCU7Vs9At
U7OvofUXt10qnAJCT+810e52zVZrP58PSixzt4v0Z3HxXcONQAlBBiX8S2OwZ9cA
V7ei0XxA2mEREaf9x51n+R7ThVJR1VEF++DDQqY0od6AyDcu1QEjLIvfn5WR7lkG
ccRF0pw3OHtwvqW/TQCvPZUojdL5kQHObcTAMKAdIk1ZY/Oi6lx5mSctxLXXRi05
2FqNsiJuuKwlDSnXZib1RkjzVeXf4aK1aiAGNCle9Ul6kPwPwRvtrClGIdmUlYeV
OoaD2tH09atXGMJHhmmKfXvy/PQEGGOL3fm+W4FezyvhrU9jV+OugsmlP1jnMoAw
96ij2wTrSinq2J8xGadiFXRuxD88/N/QVtaoF1mIYpNF86UaW4alkR+gWVdmQIXB
CFbw35nql8E5Qofe7rf1JeI5PVM3CD7Jl7f2fgepmhs640mQOtKIZVOX/iBvESpX
DgYhE+Hi5oUVzITjwq/atRzeqssLcV22Xscb811PnI0vb2s7fX9T2DUxEsjIhSV9
sjcu5ILHGi2f9FlTY6btnfQ40OwEU7+gtSGtiRhYHWUBv5A3EnuqHiwLKTMg6PQp
YA6f23YpgtCE0xNI8F9reQc1JLvg3UsOOWXmKzNV10BL1Wz2KGJx2gCeBufhEGfP
NBpbkWQh44hJP/+2hd/Bm7e2Hy0AdTHDS05RFPytQNX5rCEddRLTd8NH7mkPinBQ
uHJT1csi26WIJUXPpJkqfwdWqLreX+EHFUJ6ELV3cDInTO4UjVpHlH9NDIFJyayM
3n3R5OqN09HLL+I2Jlay+cZ6PO4w5RQU6O+Si3RY/XZwYjIPsXLSxb80dInQWc+C
hEOzHjETGNcW8LdyMTEzBQX78mEkqdECwW8HQKu2cZGAc4XjnepTrTnwznxfsvcH
a01EsqbFokSoYQZuQrydEttV3p1DwfS2oeyOxPhYlRVfl4g3ynxEEEW43AoV87d6
Sl6emggX+AidyksySNllagzBHvVJxnL+SiemOcToZ5lWf60trILNGNK66jnIzDlL
CJHAbHxMKPwrtbZovB/jol/PCfENaoo++fFDjgjiMZfASdUo3dsQoSXxwtSQKI+4
CCCeEsjc2++Sg3CoOIEvi2dr3BdUWcWmPE2zVxddm8Ty2603qm9DpBtWePhYGmQi
rToMA/KyWoHNVf9og252A2XS07/XEh5an/dN60gMvz7xAdSwjvAyKKLm7K1uJUO9
4YTRfKR+ny84u6HAf/LmvCKb8vgfpwwM2xmzvRU5mryOMvzO6Zx5h7TpxFRXyMnP
3esXlYK7F2FlFVl2+IctrfyRXkKjKdBbNWhSi5CbZ40aYPl8bD364HDS2Fxzjv3b
ISForaqCSN4rA6nodEwwZKUGj8BfQXsqb7bEFGrY9pisHRJ+K4zgZPoomLpNtgZE
z7cwy+uK2UfGEkYOmcg893jPzzG3Bbazfw0by0o0KMRnIEyTjUXuDCKp31gbOnTN
yRtYbXLswhTI6EV69CjLTVAEQLHQRWdgp8RNUPbiVtAJb4IJGKFSqMfikHh7vQlS
iDa3vDuapOxjQ/jotkfYLfSx+t11zzyEFVQ8QPJfV1R+7v76G/OpJgZF6iD0il4E
K5HIdLMeK7jggJEfkSsCg9M0ZwSfbFg0ARZZmdvWCUXXU8s6LcfT2N0OXhncsCMW
wsK6HQTgQzBAeacw3JydVxIkVILnmDZeLAmwJ6+ZaXbFFBrq3JMMgbJpQ4KyGvcw
SYofhbd+DUe5MDMOM4sPugZ+BR5nItI7f8Oaj4FoHnCghYte3AnVVRKjVdLsVmet
gRHn/L2s+F1v86wE6gIea7AGMc5/7HhDTeM5xIo5RH4ACHJdgIkjxyttpEFVfrSX
OXFMSmtZf30+8OkL/VqWIrc03MNWAHIaugXWyMNWmqr0FmwjhY+FuGiIqV+5mI4Q
ghYPuQsatlr0RQs9fEQuK6sOixc46XPpIsi9EtJLaHhUPuFO38CEqCfyKdtUOJ4o
WpLXiUNyw2aqfpyaXj9FGjXLmsCEmnRANw6ZwSUU/stjCULYFwT60/s1LtrrLnI5
kirhmw4xfG1KW1wqzZHKj+IIROVeAYDTtiFLz78NH4/2lmuKiFkM6fBUmm/v3hV7
9bSyhAe9fW1ciWJb/pj9ZxYys/vosolW5ICUoUTA+BE8VWD9+4Eb7JZHlH224vF8
KnjJI4dyVzd4dpnGr2w7Bv9s4h6GrWk+nU0QTRXm5edYnDfWIlItFYfYmtm4IypM
1mPube1C6pPwdm/XIB63cn38bFBAtjUinRs4JQhI1rBG+yEH4yRHL0KZ5BYF1PT1
lfqRaD8zzKzHoDFFvrN5eTXGBkCASoc54gHsNvT3j2waKXKvvrUvPx3ykyvG2MdX
b8pZ0xmS40mSQ6WDM/g9M1/ywJCOhhABM7uM3s7EmSYcjm2ymvmfFI2p003MRexG
myMAnZr7nGocsLQkVxG/dLuphcEMuAVjLIwtCpGaLJotUvagq2+s5r9uIcJ8KsNS
Ox6evUVt9ZRdIjXp+wFBNb5e8iWZ228Xwk3MdcvnG8q0s0fTt6rObho0j8ubkYIM
Z0TaQQLwWL8kevej2xABmqxEjmk7dMDEJu/ezNZ8uXMTbzDcQN+HktJyIe+s/P3N
BkWlDjwODrBtE8cPQ59U2geeD+hSqsiJ8THaTXSKBwfsgTGBYgCiKZ2+qLqEh/g0
iS6rZvj6njprvB7p5MGv+PX3Y4wyWXpBbUIrJEh61dRr+Mz7jfXK0pqvB6RsY84z
po5azquFmrvMvB9GuYPbvOR42YbUP2ZIYnx1s1hkO3sEZe/sefBjFB0MJlZjT5pa
tYymfNr0R0YA2eTsU3tDPEbulm16+KIqWCOYW7BxzSoT+v2Bsmt/lg9ziYPzw3xA
971NZqMT32BlKnD26wcDri9ZGAeHo2XTpekZtkapwg1oYWWKPqy4a5T3ZGjH3hZc
zWdngrk4seGHKWGL4TA1/hbgLDoNZ9iqVnfJpDw4+LapLCEA+KWwyotHL7gQ6NAe
5yoB4khRPlwT1XobUaG3T+YrmlvgB0415EFl7jmLfYor5B9y0e1DwtI4IsR1+f2E
bZAvjgaVydo0TEtTlDFMWZZ7rMjBkw6wSPnv1RY5neBf14KO6lb0/PNppVIJhjvh
m0iQsg6tkiEXKNXplnm/SIfuJ4BxmyGDZAU1x+tolj5sTcj82lYjlYgbOkcU/Isc
UNMMGUpf5GtDgi3aTxyw739vOiZ7Aaza1BziHxiWvVCcCk7dwIcLlKV+AmyH+zLD
YV0GIlzzzOwnVkVfeBFtztRS4bKpv3RiJxx9yRqrT85glbNuXkZdxsm7yEfFC6xJ
PnhiJScYWfta2uAJmpTBEm4UWO2GqoJtZ7suQrYvaKOWHSrzSjnPrErOsVA68l/i
22Go+RlkOdM4mbIMYvph9CVz45bGsGAUqWPHgV9LNkhFcCpDEvKbQ0FpWstqu/VJ
vmjjr81Q2RZKXs01dQz4cCNG5G6w0U+s2yX4OUO0YrUBVo8+c6mIpZ3WIo01lcNQ
7MNTq5r7WKdMg7IbQJ2YIOckP3bpjv91A6nc8RT2v1efvcOivPHwZEacCEOZX5oP
oXEGAkIJ/GfwpscMX9DgtGWTgsPUSb3tM7ZBJ09U2dilA7SaX/RYotUveRUpm2CS
0KLYNvbPHK/CH/ED5ZG1i+MAiVr/ty+l3ptsuJrmRzizUC1ozfjmohVf1gD69kal
x3cMqYvFHjzIxytMN9Cjt2lblldf5D1juD+rmUAAZnoApfbacFoii3Yqxgg0fxNQ
pL0jk2gvgI6E2Ak8i8b2SJgs9dowzy38Fqfg2RwpszHnu6SlIy5Q0j0jruVLkI9N
lYNu/rW6W9fY3+JqRC3erpALA3DQ3pIq/q7aJWLZXaNGUXp3tzqDPEHRxAhH/SJ5
t6UU93mTxtXpEU3Ah1m7z1tgdi3BqmlnP4u6lfnr5rBIvlQMHaJj53gem+CVIP7u
9FTCbhVvoG133C6AQOKCPSd+Aysmb3aEPPqYDJOExXaDwVKQXRwBSY86kPUaCEx9
RW1EPtIofDByKBKl2Sjj7I2+b+LwM5tvdLZ7SNor2bFGWuov6wPoNu4Zc22bEcnH
9g8EqgAL04RKDtBvStbXw67UjJHVMclEui0m0GZiTc2iolN179iGVmMkePSaLuX5
grtNeG7d44uwrqbHZVJIbjXeKVFfa4nkpn2oH5T92/kvqVmOM6SV8Mdt2qRZc0Rf
z0aFHSOYoQP7crhaYCuJMiD1fM6lYmw74RSm/y+bKYN6FBw8gctPX+FW93xW7otA
eNc8mvIHJNu2qKYKp30G1Mng0WL2gVzZhvT0Q78jTypWBvwaw+hjRto9b3YkYeAf
qA0eAvs4EdvxoPWfUun5sz/EqLtEjNYZLXJvVHPZbLXgTcJV+t+1sil5xRAWYcAk
4x0ccQjPAD4xXkXaqMI5n4SJ3PxbKyXm3uxTpKoXAJxbs3tGf6Ycs2bAWogWj2v2
GLDXeJ8aZcMSmnV0vMhFxI7BI/RgNLULzwY8klT+hk8E1OYDOmcObIdw4DbEgOTX
FTRSwJtxVem7SkVeY2qoc5F48kR9I4qZPSd7jDYeaHNC/L/dersIGSROdwSpgIUp
8jwdQMzpqsBC/cf4piueFaxKixktx/tCRuHTTY7Icu7Fo3+RIk0ntlCtjMSAuxB+
SmEUf2DWxNK78D1qv+8s4P+NfE+mAxfYIzXADMNuNoguopW/7gce7CCTlkJ+T4xL
F1volQX5mkyWpZyJ6wZOAWd8Mlj5k7ttOrPBBE8OHFjuzL0EZMR4jsdKwsGcUWZw
e8DcYB2tth/+j92MqfBFWQ63tYXFeEF6naAuBtNAK4ZBote5Bval8OFILqoatkxo
2e2KA3KIBlOfUtdCxsZSwp5jZz9t6Z+w0jxeiS/buRCy0XDO0Ap0NWNYxLM0qrL9
Lfr/aa4lRCR9L+GtO96oLpCLPnGWYeEhsQvE50gkw34eFE7jlfal+Bke64+sw52y
vdduTtMXbemdhDnQhkNC2uD1amcDjZt0uBF3vdoTGH9g+CLFqD4Ap9+bVWQHla6u
5HdHJdsuk+GJzne2MtQRLfoYoNo+yjKzZo+lIRRjSoH7W5PEZ8y5b9ksfDoeR+ez
pW8T6u+GOrIQ7NEUYCyh13+P3dGgaxtizBQSYgyxNTDTYxMXirHBnmPgSNvXaHou
Cz2QHTqIbnk1bUCVQCg1b16FowG6pn64SnftJNGU+6wLh/y/SB/GZwb9SsFB1DI/
64k6p6qDWDteYY7aniXKWdKmSll8PBtahuT1VLAUfawttYd/9n7rsDOMVf9wYZLP
ezMJMnOAEvzp6rntVQBBW9QPuTkGKuig6mrL7YK0yQq3/n160kt3crCG5cnk1VVx
OAb5iMPV7oJb6YCO15jtCe+OIGVcllrlS00EFasN5qgMEcv9ij3qEf4RN/QLt8a0
mlu8AmexQpWaMJvlBsCmkR1m7R+8gRhsh9C/JeUnEJW5G05BSzqPXSLhqT6Dw4F0
DZn5FnarB2IRbMj5rz94Az/VMWXVXLRGOwRg0qJ6rHcTHsZCUP6gVRdofpBYdygx
Vv7Go5KMVW6onAjLZQPR9ejwFLCY3WM+JubYiibxWd7ON1782DfpuzccDo+Ng3yV
LOFr5mmdFfMwFaWrfMfNil7tNYz2kIQ8k1jLe46pCHwDV50IIy2A2yZSEySVovpK
f7lazMNE34qIW/29OE7LwODKEdjqKbkx2QZrD8uYXKHTXQLqHG/u3HTkHBrZvgSd
shFl8d+Xuf4XT60dje/zkv1UY3RZce/EW08f8biG6uJ2osWdPFzSeK5CLSxw3iPs
F2Hzinz2gqB1Vd9tI9dC98scDqioXlDk7N4mbYmJHH1cZcs6IUTAd/GLN97hXuYj
bvWm1ru6VSF0JJVhwV8bjgYnxfrFTn7+DMOhCNYWZiKW1uhYs5i8om854T96+c1L
AIxZ0aBbTTCWNfIV2JZSWORDDhRk6ksC+L9Fl2vHdFHdLHxcnmxE9yOS+Wz+epaq
TGLI0Mxu37UDti5y3qzAKyI+qzUUUc/j0q7hKaklsq8snStFKKbhRaptRXMEo5cu
unI1LYevm9vGQP6+bibBY0Ij2f2rJAzhtt6r6LdAiAIYNFWjC5InsCW5rXSXYSDm
WELDOlth7Rs86pV/xQfLdRttMtaBzKZapTFj9raAmh/VghKLoA5WgK8rqsIOjcI0
d8dmnglbut5ttxOfEvI2s1/OtBdqqHViA85FKS1328tTBcMupeHiLJuX5HVu4VY2
l0Gk6nlSxSL1GKMH5iIBGxdMjyPj57AVX7CUjAeqR27w6r03lxoY6yYs1S3J3s9z
ntA7otkAxWjHJowV/3wSICcafiz8OaNY0HqPN9ul4hVw/Rjq5SY6Y8b86GqTql5O
szDx4lMz2+oSTNRNhxXBS116cLkkszOKgQWooZJ/jBdn8b1fQDBB8bSLKIdiYJ6u
4eyTL6bvZN/jtjVOC3tGYzma3fy+Tw/OMnEo4JrmeU46JTlFPAbN6mU3UPLrfouW
Coto4jJsL8PI3LvOd8lUJXNTYhBPWxssnRhLT5uyK9dQikvgsET2hG2a0XswWM12
GQoTaf5NAj3Pe2z4QPgqgVYq17TnRdbRQRCsi/T3CWntPs73s5AuP19xWRZire79
TQ3X0UFAvSgUoik+Ob5mxgX46b6h6OX4wamUndmG5GsjuwuV509p6wEFOA+ihxLu
d4hgbz/RQxYZgdSwEIPBbeqnuNcGgeF8O2RUFdhFux7gpUmpOIWWMOBbwfEyBwvB
cSkyAZZeAbGKL5qqail6qqa9fuk8o9VzU3HpPoiUFWXo6jaf9smuNDJJJ5ZnPOHT
L5Sz7mUXAbaBBbJX6MhKEaCArwBdkDuMb6tUiNA5qU5h+Wpb+N4EKlw+eBHcbws4
qZWZrFTOWt19Nfw9ueiXXuJ2QLk1Mew/iy5RSlC+V8H8HNUf/k/jHMkFHbDqo7Lv
JNCr5UJ9hwHHCvcJljfXiOUjurOgGmptE29PnbG+8H33YCxAY9pxOJj/7zYhQnc1
mjQ3Xfr7hU+NjHejc+Fe3t5/7Omp6H7naFnSGST+RlqEja5wUzvfj5MaG4cQW5AW
auOH5k/MBElypnTaaI5LtWH1lAXFFMa60QX0dYaCx7VRc6pM1VWVM8PcN+H8Ecox
QNqwbipzPs0gSDCbuok2tm9jGmT/moPnxpjBUdgMSSPBh4KVxFqbqelqmJEp6q+S
dpF/mLvuDoib7L+TkrscnpE9z83aPS0f+2yRF+o0CKd0fbVuXcpl0V+BKC9DCGYP
+7uVO6nUJwlg88zkMEpywHVhcUbAg1x3fN3DFGQB7vO95xj+D7RMODeHk73d31IO
K1txNPxT68Lqst5OysTuz7uI2kWCL/6wCjq2r5ejnU9WLkBBm8R7xf6CzkbNou8Q
9IaRqfnDN6VwNxbr9kN6BzuZAYR9rnXgVHjroCjjQvmEvp1P/C5d84K/Ctb/wf4s
sRS+ubIIDOHeUf2Et+z9vpUkvHOdsrBGB3liF+kCgjI77eymdplKahdeik4mJn18
ScxZ21OSl81kHCARfGe+12FQt8R8OFbAoFF0AvX/qvgz+M8Kf0shSPctKgVITo+F
NL610vORLgB5TOwjC/3le+KDokHmn207XKv0+NbBep2jMPxwOjs/+h+Qy1oPo++h
RDMauIh26t69QarRoU5OqnpQvouLrTpson7NngEF9Uh+cCDfFgWXTBzUNV5C8HM0
x1wMnMH2xxJYdIh+CeyB5ZPvsrg3IUWUu57VTXjXKJlP2ZQx/qYF59duPRL1NQrH
1+oxYL4RDQZARJT1cSjstpMq5SyBHVm6KFzlvZVEPaP0j8VyWghXZSpN369ELnuE
F3sAhp5xfKFWvr1Iez4X2bpQsvWOOvJnobaInVimp4+EJ6D+ajizVgckNxK3LKMz
gf5DA3kEu2YG2MPQDMI7xyhyrVApSIxrQPvbx+RdqPXzDYZmxOHJ9OoUmCisG/tb
ibQTQbA0uJEvpgN5ezMIS54DqoAnqBNWFyx3+MndzOfPHpEeSsWhFvi0cYoliV+g
7tF+DCaX9O9hRdmgcLSPM8EIcLLxSZesMVU6tkCA83jQ3YHLQBOp1KRaqRt58XYP
lfvy9zEyHgXI294CBDISizPTcUfgvJjTaK+h99Qec7YC4Ho2nDyc/oeUhio1kbTt
+7GU52s2bkxyTtdgUhdYQOdiCLoLo/QYXnUy6TcFXo0kVIqkB+IfLSe6U9dySqFp
d3d+xa7ovy8BZIgKU8yu0gYufmIfnGyIryOijQ0mR0pg8VKnqWX4WUopq77e/mBE
OAWuIQMsacGbc6BPMTU1/0OIOrrJ4lGnBQAVxWAlgF6rVyPyCXN77X8UzTXyOtZS
4C76lsCO+h7xjhE4q1EyiFm5HO4ibG1dMXwZ9HEt6GvgUzXNgtFW6KEaHyPmq/DH
4CxR5ZT4DypcVn1+yyLB+E3dbUT+c2DVrpIU1KkKdEtPjWYvg+yKs5uJO3P1igJU
CsrxH6oaIMRP3EDiX8NnElZaPmA3ozQksrgqTH1c/Rr0/VCFHmsZfkYxg7Hw/7qd
eUotV3o4h/uVGSHdfS70PGcf7yGMNepuKotU9dcYGy0i48/yeurc7Zf/n3luAm8A
rKAfG6pHj2+LPIxtu1iEKDR3XieIYh7q0yLyZ2pQT+N99Wi9NShH/PBtW+rgqgW1
nHsNxcleknPRwVnUUsQK61y2Lo+3a1X4k4YyoVqoumwa88oLHyDL+FfXtXPgI56o
iAIuuu6dI0QDiiKMpFr6dF+pbD0DPWm5Q5Y4BLnYeT+nNhU6tV8q7N52lZ6MNnYU
PdLDQUkzVY3b9aY0IjwIBeVLORKazb82Ni/6aJhqu9UAQyUGyg3Y/P/cPci941Z9
GYV+/0j5+s03Knc/dO0EGiHJ8Wdyuv9pgENCfHsv/iSxSiHnwlaPWSvE/nN6mf6o
rutrYQin+MAqNe2CCOQn4ckdcttKDapvkIlN19zPml1BH67V+Osqk6rwnnzBNmuX
esKcb2WW/WF8izSIw807qt67jtkol0eqpYXgUr4L65jjKiPizHecu9C1we7cFKXI
FDHzrDDi+EMM1HEPk+LBmvZ13pznCDEDyQIMvexTYRJJokpu0uJrEIHfR82M617U
WrftVCSCebNmpQm0vmcj58VAXmZRVX7S+HZwiKzWcN2GwaKVYgRlfufgfj958ZgB
7SYziJNdG77Tqa6CT1obA/WVmVzubGrcautpx949+tN4wMf9Sm57hmAy2ZSfAgCB
KxhiOvDVtJJQtP4Q4kb8AB9PRCS90qZLIhVHm6V0fDFTqLn78jIcAMx0HZMqLDdf
JrEcgnlTncJDK43tm5MPFcAmOhdz8Ny5hH0dRjGQwzWA7JdE1FOq/FHD9Os4Ksrx
afazC7JO6A+b3FF+6TH9RltpwsMt6j8ok8pzYcb9sYik8957hAZ1Aj/l16hIxdtV
MLCEPXXu+Fba/oWGQbcGeKOiiLyv8/Fp7Ysx5BI120OEWbAEA1/3kk+sLGKmTIZJ
u4HMPrUQg4bF+N8vHB+jSTHOhUKlW2gz+j1zGmarGlwXQcf5gV1KIJoiO5BCxQeW
TVZiLT0Yo/Gf2iE2VgBZRwJI1/eQMViNcIWnk8cijm7KyCpE0l4yc6U9j/yG4WL8
/DdJsxnS6LWF4LUjeLaJ2LkGMkcxDSaxFfQx6O+RcnmVdkBmFcGQmsu7zIYzd8pm
LGX9C0BSq4MaTgNb73tFRFZ9rlcAn5uHPuH8x62RaYtna6JDuF+FeWMNwcecQd/Q
p7mDKtiEfM+gTLqtdMYQSl7ET63kRysneosd5MfYjxrWQfsi48VtSZT7K6D9ge2K
RrnWj2LQXqOXSCgu7mWpFFowCoYpZrsJzw9LI2ptJKJ6DljagVJ/FbyZUhY+lMhG
pmaWVtO8L85eYXkJAvHFqLiApwUbFrUzgUd/eeEebhl+GLP6WluAqEhbTzbMO2Ue
YrXeFeg557vXPh+CJMlMxA1eC43dgtT70DuaTkfeJ4QSRs61khVtJNtYdl+X144s
9cYqNtxnx88j4uFoLY098g5CTVNyCmK5HTcyrvmF9M5B6zKVMkTtDzvKjfhay65x
AUGnc8lGlpZpjRMfPZB/SYLvVqR4kKd6nplxxunfKpkgFF7A2iUvrT4jpTDdyQXo
Tls63fdEhlOy8kJwIy3I+WY90uzjyg3hQjp+0rMrdM6SsrT0GTB+/hisxtuYITpJ
kwlHj4NpDxcGXcuykUirDGUFlsi1nhrbaabGi5W5o0fnHZuevh5WNV9KSHuM8Tsg
bu3wpXHN3ypMuh6F5IUkOlig6tU2iytHVWdZmubWUrPQZSZcBKsxnmqebY2QZGIp
bc7u9szGpmUbuucinBox0uyr5KCtx90OmlCRplpCk9hcPDAbWGIxwEpDa5p/l9qD
+C4X37UGQePSH0jJhe5M35ihaZFeolagS0qYiGObpNEX6hiYD2YxWKNLtJC4KShN
c/r1HGrbsy5BonALoDJDyzvxTdn51LCY4ibWVJD/tGuKxjmeOEUtbJHYnjW4FGLR
OsKmQAA552XqhS3hD826W3sAuBmadjd6wq0yqKqdHs3+IDstt4QmEG4UvhHYGDPG
mf752K/Lp7YvOhcJ9YEsEExeA6Z6hjQVE9eTNP6IV8VSrvdfn2yOPo8yQkFaymSq
Ygpa5o33I1k3+nLQ3XPkH4TSRiu5cfm0ImGVUQciI8DRBPsxc/s/GiZxAHQlnBM3
yLXfHbPKFpLcCjObS32bZ+SvrMaSvkDhIwCkjH5seKYCqloc5QmVHScTivfy639g
xq3wSwEEe3850XFB145S1+rfFfh+nXDcwtWmjcKr3KOWKImtVUJsm+i9Y++vgJg0
lyYGOiznQr4vDP36zb30FSivNPzzW4Rm2+mzxGdTVhA9TsVYYv87aOWoB+wSLM1o
iHI50nZwACbPU/ybrY+VAtQ8f7hMeP9hrZc9So8hjUGBbDVVcSnCXYeSGsK4KPaV
CnUmv8EskXrVGRsubawt4GaNbBW8GYjntCkyOZr3gfyKA0Zk3pxZxF4yrA4/Q7wA
U6848OEcRp1WhnBo1ULFS+7cHkjLPaC7UFZa7BqILt1hMkWGFlP537Y7nMBfAQWD
CiX5L4fXFqhpJfaCyE0NrXWBrUGWVnlxquM1xleCIiEXyBkMH6DJMKuKSO55mlNm
RwzTuBsUuVuBFc3uYftrEZjpZgx2WczMvWXyC+t+aWf6xRkEYpkAhCp8JuQwCpMs
gHQaJTYN/kirwL+Lr2XWdmhvVmNT1LV+BCr921SEeT3wioD9HH04VFr36/qQA41O
EtW8vMmJsHCvTHXN1H3isIHXrRJpOwVvrfY020to53YLBk0ewmBNfX9AWnZi3Mu0
DNvKrPh7T+KosC3fBORYF78vGFMoSRt/I20mKgtxwSyLJSxK1ImMkc2Db8tUluGd
Pz4AkYGxLlYRTpSZfsDOhLaZT3iw9Bh9cH0BJO4NEnpSDjZOh1qTuMJG0KKKevqZ
FiKpLMzta22N6YkCxIwL7+l2Aey7cWENV0pEvHsVsfCoxh5VcQrWDmTIkomrBsW3
ujwsIeCHz4kpp/pQIOOAhEQ29wzUmELSs5T0O23IzuKg/hRwLxZ9gzJO1UJrJqNQ
0rzPAVkm2d/BS21CbQDYOzNvhKioXPV45q13tJb2mbhO55JZ3pF5KsIs6V8jUwyA
PY3ZBS/VdUyLm0AuBPcAXp3KSTMHkXlEhnQ55F16cxwWA9kj5voyVXfKXqreK2kz
S8jDsNkLt78rO7BlL49UOlK8E+TJ5+gjO0tZpxaC0nVSPnKhUNx9j/bL8ptnahGx
erqP173KEaqx62aHPQr93w0G6nDbqDnNzRVCs40jVlSSt95PfivJDpx/7BOjLZiK
MvU6LoshElL4FTdfKzbvv9A6JIW2JqeaYLTPjaXnV8Px1kvKdzyVS2HCuL689Li3
wmenlKzU4CVEtr2UBUwMQdOoLvdOf7ExONNyNAo/b8mVF8s7ogA0lCLZqmC+qYoA
CLz2ljAD8oXkYVlIiXBiQVMz0RZAtJYfrBrzYDseB2bBufqZNq7W6xRUlNUsOMpC
4khjRHfu06xD8CJiYL3qQHcU0GOmlP82hZzmTYZG9k1QU83ZaYSkAtoStTR0xHJR
vWTyTlGiND5cofdU/9k64S8WOgT4I2xV928RhQI1P8v1kZzIOre0oLjJXhHO7PQg
kzLAFOnE5OKoLuTfqnBAh30u2EwnxhiI1vrhzPd71UJ4UTHCnrC8EtVZ8dmPA/fL
afv24EFpFGfSt6yNW8/Vg3caKri7M0hngP3eNshXyTFKfluJP/WsepR7q0biKYfh
FKQqS4NvBHA3SyrQcP+8ltMileFqXd/E218adw0z9tR4Ju4wo4EDoIDWxGccZa+7
GbBTgjMRlC/SWXUxiOZntCowqm+S2C3pZIPnX5MHfLETA7vUg2EI21RTLteeT1BK
eNSKcjXP4Gzqi/3mjJozajCI3A7IUDnAyNc5+opGQ0pxRRBnvAGyB7BwvbWObod/
nWwVarNfe6H/vzeYj3TZQ7mroOS8Ur8vwDlkBn0kfBJckuIoEJYvy4fzf3wfqVM0
70zcbNqtSB98Wf36bEIj/gz+EI1muZaOMi2lE8Ey/Y0TlpE3PaX1YSBQRU4Xm3oq
MXOEHKpGiTSUtEDHf11Eg6RnQBVVriwISFXU+MbZY0s1VvOtRCZb+ji3RhoTxQge
vcd4SSL5OI/DYwCqN0diuV0T/oXOFElvW8SMwMO0Ih5EgUfrA7pKeUh7PvTedG2+
ZDB6LKPeQBYqIqur8pNZM9vmIMx7BcTUT+C7W8kF7hFMaeQ2+2whGNlmgxKwRR6K
yftwfQlE3pVVyNh5+41dbyHPMMnckHuBMBiumEq5k0Bh3r32Hi2KIwV5ppoJBGjn
3kd4HRt3JV9nqhSveYyt/13q46xkOb7XcniTwK6bPFFOssN7LeZ3Aa5/MiRZWV6J
KILE5Rvricqd2h1tCCzJK0aensEvcIRy+1kDta4wZEEgx3YIukSBxTvP+KsWhybL
0B+1ZN3meg+KFij4YH6NHuUzA+0mEeEYc/ZafNJ84d8nSiYE1T8fiZsGmpxvCNMm
E0l4LX7Ll41Q9N8BLXpNqFxOOZTWYh0lUDLkVccmTbMZsKfAftI5C7GNhQayQRLd
4Ckv9p70CAlCtEKCm9lawSssyAyPG7kqbk6/gIwPqztp+kOGevGJf4Xg/y5Q3yLn
3MqfubwxZQMGLHvppU3b5nJ1j4P11gZj4+58H6QoIrqSb+UG3utHSsANuuQd5Cg3
x5xq7FexVDBqZZKyXdTvKWHnejXrkQxCR37QctzulM00kZzQX9uzhDWzzF+gbDll
ygk4G8sitv8ZQPTOR5xRe27flG2bf6XVrs2Gv8x8PJ+gaEc1D1aIFvG1IpldTi9l
ZMaRE3zQHmYtmawJCx6W7+NKHfRWjjYrBjyOvcoIfaZnjeiDOOxqt5DFlBqVoCE/
b4jGACJ7osQ4F3pX2upWv1wQOmv8DJ1xdt2hdfhUcLarAbHDwI4+tYZoUK1er8Bj
eqZn3lMm/WxSDV/XngOKo3bDKZ+Of2egwMomZmQFlunk9VzeQsdqln2FG+GF4l9w
gQrpGeK9gZNQRUHp//7IxkXxSgypUWuA9MRzUV+c4ut83l1Vu+WlqBc+VsCqpszO
y7rkk6RKXJPs0IIegnydl+0PIuhfpqoMsZ8DodXT2Ab7V6hIT/6a+XnJsrmrnYqA
PIYmgFDWD4AJkbGQ7UXEb4y8q1/qbZpnjQu/tYfP9NYU5w9okpoQdj1KQ+2p1qHw
yOyBsY5YCLS/TyT+tw/Odhj++GQ3LFxuerIs7yCGjOcjTkqI7n/43osTQ9Tjr+X+
7/26qW1Ui1tBaFoGqYTo61Der2K5k0VylKrC8ejs9oOoxVf+CdFlxYBvzCvy/h+M
AgUcDCjOEwSEFN1QHAXpaUIz7kZVkHIbkFvgI+rTvlh75xOAGzT+YeCrC+RUQJdk
jtlo7Azc4xCyQGPu6jDLJsFlPzEvyqJy52J5wimGaw3p3/s1lMU4A7o/h9lWUii0
dXGWAi5H62T7LYt2J1H4ksbolguPkz0+y4laTFf0bj8GBO2qjBWCohJjCJWP8BOm
YHEr9zOH19bNKhZUFK0PGEGKY1oZu9p4Pd3SmAAoaDC5z/xmf9vUvN4PKODTxARl
g4ZphuPsxZUFk2NpjjEBtT8CK655lgJ3G9H7QdoObMWmbtqBjd8818tVAvuI7GB8
aQ2Yz9exDWLhTS//Z7XhmQvbn5EaXWzEKIT8Ux4W2u6V7IhO94opImL2che/xk8x
WUn6nRPLW6HLMLlXplCY7rORAeO3d/Mq0lQGl1bRBT0wjRz2vIrcr3CjWKuA2AIu
YSTlXltOyRF4HFK7w+gEWFcTyHQuj1225wmGsEGle9CIa9tvrpTWUaQcNQ9rugnu
kXxS7Al7VnUzaVV8ihTDQCC6YC66znpXADpskdZNVKKFoXDs4oBi3vJB8jPmQugS
vpRbqph6vD/UmRtWWvmZ8sE/5/CBBEMwXhgC+KUlHZKLrz8uTeTa0Dgi+ZnlTEy7
Kni3LmS8w925w22XWjEImS9MS2qvhDaNz4cu2gPHDJ0XxQbvUq9j76DPEp0ijBci
Ewn+of0KBR4DKRUcCmprm2yxfudgE3XE+gwEpqRqw1FsonjvRw8YFZbprjDdTegg
L1OT6ji9mKEdgMUP9QNt5f0H0cBoJNUJg/AXBICnC52eGtE9j+n6fomcOdtPR15Q
sjY1zzvnIY8tqOcjwsi+Z01al0vVoXfxo4ChPlNkM1rROzga2S+vDXYi3v7khpJl
MjDanQiXreOH7pCKDT47TGKcNzrFtMTJEqX4RnWCZLq0e87UGXqC32G04ZJlBTZO
54nrP6PTIB/hqonElNVsrfpYymchRdYhVHKwyxHfwaU40CujHgVR69zGEzfzB1Sj
H4OT4cDBv8fcB3gYI9NW4sD+ozZjD0dBpxOLgArdhnTGRQX2zkWU5hq4zVTxZ3mz
zMmyQaYK/iETPKEyPkBQ3xA5dsyjfn07hLkGXZEUvaxtY+0Kr8GtejhOrkXmucS+
gr9QV1o+tQbo1Y7ZGNAKiTe9IAVtNlBZn7gNNeFI3okHGAw2rB29XZjGJqcaMyBR
JcBbzIQnnlJEELQooykBN/eBQJ3eW+Zl2jloRuSn8/V4FQi1F6aTh3MkUivXqH7v
eNfu36AdXA3g3kTzqEvWXPP6dqbxMQZjGUPlz1lwygbOYjWkgvjXynnW0KIkZIu+
pnYM3xeEKgPId7eJTMr1nYIhYz7azAsClu2az+ffXgTjnMhHAHqiQsswd8VewNEz
VR9LGE26cd11fXyjiFBa0Dbb8zxpIos/F7vpXb+eLDqoQMSIxNGtnZGnXSztFmZO
cyTwYwQIFu0BeG1Fx9VWWWESAOK8Q8LjiWNaqrbSaA4i6JjrYXgZtumrgaGTn6g3
1qRLjfarjcCGFI9UlpAMfIjxCYti+jUYBx3yfbMS83350U9FcYSZgfSuaXAhgeED
q1kan2F4lyPXJZjS/5Y19cE8K8JaO58u7BgoEGkiYD6ZOKwtGf3UvzFX170f6byM
1DDDaYB/FfOT/+fL8KDjacOKqni9/XzcH3PzOeKRKDxCGfK7FqkdFDFShw2AcEz4
U2AVKzbG1+lpBPRRyprShmCbGBx1/AVOtpSGKnXh3ZNwSSxXSnJAoo+7oFbZpD4l
MOHxafwjvYdMHVh1/iD1W/gJvb5HnzHR864G0SXmr4I9I0nu8olv5U0LilZbYDFZ
Q5fowoZIKjyfMoHzdyzaDl6+uJf1gyn6KMotPwepJqza/SIKwydGvY/VtM/WT7Rf
Bz+c613olVPLdojjnDN7syHu2mcC+n52Aj0VEOoIAtnFJMALWtaEKhJzaQWONG+x
G+kriEaTaRpjaouwWH3og4aQZCjYkB16o+S6t2+Uj5B0Tj4F5QWpLe2m3OBHQuzR
2UQBnck+tEl3BR1olPkA5uRjJdTDORaclB78jclmoc3bn6BWb5zcJlrB+Yi/Nf+V
emKzMYrbt8TbQMUqTA+pM7rfb5YDiZvkaXOGMNdLoU6VL/+Y+k27UByO1Hn3q22X
+IfImsawtKN41gNUAWrGUBSQBbVotV/ycN/c+idHE0JKmVikTJvtgYSdLavYMapr
Tg8mlsmvdzGwZmeKkUHrsVn6fENzpsZPo6i/1kmveKa16ik+it0qap5hYgxrBrFK
yvWcjWA/2zTKMSGTe26p0d/NQP+QjKAkawCrnOM9SsttXTRTafS0fgupPAJHLRtL
WdJTb4UgFbnQEUIEwtYeoCNnJwAM90ep1+JzwjysPGpnH6GZ/CTOlrQpxSTJUj/a
XLTPEcIV8j+NLxFS3R651AGKT05yQScPHRsNGozR1xhgWcxN8y5otyw0vwIDknTX
XeC+qNoGn7FTitIk/j6K6mPUjVXvCGONGeSg6oHp8+sAuJZT7WvRGC6/+hyx7ZpB
N4DG6HMmAp8T2OT9HLEChskuM3L2evJrS7viHBqQRAfJsTYirVCQu9DDltZCpT1H
w9W2ZPNUZPR7bh9NyMOhhWWFIFMmohMvZrDDYOMEcKajfgSdCLANkfyRnx6a9sEV
jRV9CKkQtruZ/opD6Qk3yi4Z10b8eIfhHYlyK6sTYlo1BpCSbLC1kp7JUc35bgXY
okDXgTPIcl886/8HmVk423VGAQc43R9Y6FVwUtz3rWU2R/mEpfdDITnFXStsq8x4
Cp/ru/w+HalnhHrc+poIRmlQWZwQUrsiRXqHeDuIeDImTWiBx4fe0KvUm0mJSKGz
K2bF1nePKiygmt3te+iYYVln6jWXuwzkWzpPWHnyM7KC4tm66E2ZP2poq3MOeXaz
TwEAF3NMgRySObGfhL4kjx6FhYHvKG8zWxIAkTt+xf2fxT3ssPdp10RGiAb5zx19
G5G0MHngK1ntk4FxS3pffYFBakcb2agpObID13Kz4f6F1kh6yUOU4P8hEXKqofyR
2Bc/A7wbGchQoMINijxa7yGMS3zbUs23t0DMswc5+Kg2UTMGz7frF+v0MZdA04rL
RDvAptMWh05tRSqqZ+AlirHc47yJ6TpQT2t9JrT4bti5yV0VpgkKGewK8yohVbDx
0bnmPW95o7VcbDEg/RnYKMfnM2Z3BoUF37HRzeyY3pM9Ww3eXczOxgoKxTPrQmig
hUYUwcD/HfdQ9gd7k+rbs6IF5v4liuReC/UDZcdozbVV+idxA9q+aZ13TBa64S4Y
OKF2dz0pEDh95q7LfFb+iep7em0f8c+aIQPGTHnmeVlvRbXXm3g6QmnS0gUMfbkb
zVHtZ+Erfjjw/TMefhBI6zYBSmG1I84m1wikyh9iieO5zBZ808WXop2nHCtAGpWh
+yOO5QWJ9KnO76KoaLx6A4YMe9m/bsPiaYGqM9IEFgL3MOsVEEqzh6wXQONML562
WQRHZz0zk0F8WcrJFcai0yUZmkaeLX/IYjKvzDdRx/KlR5bsx8MKmucadgrWFICw
JXxkNxAsoi6bVqse8U9+4/lHlq7hsCLVGfayCRb6TDhexleCi4T7C0I3qc6BM899
k0IovdKkPmbkbQcVdhzFixc4OdENcVMf3RygP3BrfQ965YS/7RQ6HbWBVaNKvTk/
YXbkWFdd03wb2ldZIV0oiO0nUiWcoCtV+tHGktqEZyFs70KCiLF8gyg9QC6Sd8/V
m+4t8Tw+i9qZZYyGFmqxmGEuem1QeIW+qkf0STAVds7NFMDNn1dVht8dYDQ19s5r
F4Sy5aGV6usq3MHfGSZHR9OzhO6ImVAVmnXpK09oJ3OaBzPySP/HznDeb6HTTycB
miMI/WoEXuc0UHzj08FklyyPHuLhhXpKA9c7z8jF9XaRbyNwrIRI86L0g6ui9RJ3
9nDro9GsZTGGa8cmC89OY0chWio+GL/tRKo9G43408yDsGSY+Af8P8mQIanSB7gM
RKk3Cj5DPOYrDaGqOCZxEF1kA4sXxAdyuVPiR5S+VSrZYq2WnUwlDnpsvc1iVCPM
5gbfl1FwbDxV8g5/nDw6h3itYyor4ioNBciD15WASc1ksrxH/dpPCNNvMKqt5yW+
nRPVoJkvDC9FSN5yo3BhLsXOvD1yv0pnKNA3tV5WZeBeglSTjB9qWQe2SG9U8WIJ
JnI8DsvfK7xE280BhlG81ejNDtV1RPYdMHeqgx9ze3efLK0D+gzEbQk4gRDh+Yc2
6G3+4JkrbbW9ED9JdwJYPBU0VVNB7uaWALfM8kvlS77wMO7p3bL7wb3wZSXjgoHw
ltDr+FmXvuNHdJwfddPXrR7t8ZQzR24ymQWQmHSx6uXwjq07yjofYd4AMs9vYaIv
x6WjilXiGoOUV4CU2MHeKwzI2gjY+F7Pu4ZdWRsFoblY0nTGEda013HBCAW8zKZG
EKFUiLv74JKxAUzEw2eO7ME0VJEIFC6JXpTQishKLussc5Rj8H5m4mk1y9Cbj/Jv
fPWUG42iGTILpyDoNh5XOuZaxKIHbTP4Z9Ghx8/n+ZVa9me61cpC2RxWmkdj3EOb
WI9Zx95d0gBljqHkNmL+JBFXPkpZ+dG8PLg+nJHssAZaVwezkze7hUCjlJFYagm7
ET20f619ASNsErm0W6vfEOW9Iwb7ryiPFNwxBCpUHsg3wurYe2OY49VF/XFQlEsE
GkzEaQVDgNmhfBEPyPZa0znmCTcQ9PCyDmIdBkGEFET0WdsYmja42yTQmP6cK7sq
2Uzva4WFR8yTtv2Q2HaiP/wvRKdRnejXRFgW8nbklu9oOxsJ8WtFLHA7PceVpkBO
DeyrzIR5t64q3TPlP4Q1//k2oGC6SGkm8RK9a62S9060Fqdt4AWWRl6OolvlBPgP
zp7VEYcFEqRngpHzMdO3jduimY+P5xFpCit6o+UXJByDlRuf1HIvqna6xFJBgWtv
LfUJ/pUibEjgyoLo+ejYBgRhnfXS6IXG7cTT2Vfrvcio1LQiCLZPL3nQrELBKrBa
lilty+stM/qAyK2LqRwHZRm8Fj82b0yNTLwEToOZzUAw2KbWliyJplHnc1HVaXeD
QH/BZe23IYKmXw2arWRASVCcKVqdG4fAC/cSHQ2N3FMoZovZTNTs5W4WJjn3BvsJ
u/v7Xqd0NEPJE5OWyt+bRo+F6T5dK7Pf3GiocDGIRrCm397FMo/I9hU6bLYvCz+l
xHUsvU22/FkXxAU+9apx2ho746w7M9FYjxUNtPeOGIow5Pl+VjzAXVuZDhRmC2kn
15lS31DwAJlY0POzbOD45kPUguogwLWjDg0qWWyaJErd5mIooEfsV1m6ODrGCgsj
W97QU6gz3NNumEn0KpXGwRKvLwa6atsP1oEIF5wzpHiifKmu6shMjuiSu0Q43n4f
2MpBEoX8E3CvNCdcV28jrsrQWYVFhKcPJ/EBq8EfSIgJUjNXyUgqjAFQbCpg+iWD
MWD9DeTVdsTeLhaRMydYlShlSigdH8dBxpA4fAqv9Q0u+n1XVr8HGcwjDFoPoCNf
HiNjzD2lS4OFcjHWxpRu4m/02cvxXfEBXV49wAlqXC0JWpLr8jdak8EY1EP+X1KD
6vOLYYoYBXVn8EWyzLe7Sk5JhwMIuNnGnczBG7CQ9qVY6TvnrSTW8ACA+QRRSSir
OokcG6RdoM/NkmS1A0WbynLrHDRpHB2KXPViGYGeMGhdXYFxxWpBXGRHaBK53Sl2
vVCHNpf5gJbn20F3QwMQdj1g5zbuPz+X6XUrdVBKMkJ5m97iAy/wOIK7tu4xqAGo
ge197HMK4N5BjCPZK/ar9zLWXdMBihwvWkaiAuZmuMPi0qX1ei9cY7a64a/QCRL2
3GHjXV2z88BfZ2V2lhDaJVxvMNGBX3o8igwlcAldQ/4Lmo8ZMLt8COk1AWVRFshV
0dwwvizd3NRl+Mfw6g+1Rtyc6bGqrKzsNufnbnkuqF49Ky280M/ikJeOY3w8DcCX
1WovdbmHlwo5F2NrINrW03c/tMlpAwALXSuCNcwRyKYuYtCcrcF9jSyQ55l4wdkS
jN32QjatywfnicbqYaYMcg82/0qgn+iqV99QfiHviwfDnqZ0X2CGXy3T4ATlTPpi
ZNdFeQYKPGvWjIF3UFWkqJ8nVom2FOaPH2DdtsaSUM78THBJLMiS+YiAcan4DeUP
/WRH7m/oYEi/+lLsknPJ4LL6j55TYq9UmYej1lNRZ57yQXTBTkXz8oO6pwyeSGRy
YCJ4MQo2L48RQ9fyxt9pRMTzc33SnWgJoVypwWxCfBof6MuKE8Tw4FsuO2AmnBvt
nz9jLopVXp+MbQTH6c61/DsD++nuZUE7/lz+f3KhdneRAE7QrWlarGr/pYVyLFE3
wbvDlZOyOvGpIiIpoZYH+YmULA3PL2+O4UnezDjAoMzUWHn1BgampyY0kaCSSwd8
Es3GUmHa+YUYFJfVj5PMLxj7Slp/T84DvLkHc2ERmAUKUsrHwjxpW1a6jRGutiVX
UfaI4RBUzu+dQEy3PVzKl5XG+AmP1NlrNKH/r1EWGlIJx0OTxGZ/OWRg2rdd0oFj
gGTr1sg8XWlrNyUwfDXhc2rEEvu2s9S1F23FIrawzst70RQXy9AEo4bMQi3E3IdS
pcxEnxvgOMd5u6j/kD39Tc/Tn4c8frXRVP+dF6BIjCGk8dT6XMPBmByMcbOFM/zw
1FZ09bSIB8HXJ56iNlNRnf9i7DOTc/ql3chmrHqcyN+9/SqFrd1Q589e+lP5HGcF
xB5AVdPJcyJpUB1vA10Q9HeAuv/FhT/ZPR55x7H7DRzEQz8XQlwjMhwQCc6ekfQm
e4W4DzohwiYxjzKbIxNz50sIZ7BjHkdM+ddrmFs59OAybpvlFoBAK8cq5BYC15vN
a6v2O1GwZmumEK6wjf9sXkYZ0Y+k6C14a3qMUqQqEucirrV/3oeKhjOFfI27wkD2
5nDfKHtVE2KT4WEVfQHA2cSWmRauDG28ZPHe2fRHlZczeHvw+EYwQOT1kioLHxlk
ejVAxohOSjkRRHJAxIS/ypBMJcuFaIRnOr9v+6tRqUpEY9AuOVZDTg/ec++LhTHs
IHL4HFwUMgdtIStgv8OwPYy9ks6IpUt+UoXVQYnkeuG6v7jYJR1Rk7lz+QlbGqOr
ey2xB2Q9IvttaqTdvU3OZxATVxOhvUq9CieX2+zCxEt9lbV3n6WvJCHgMB72yDYm
2frOgveDVMXVKeq8fNaMWB+i0Tuf0pfjFWJm/5uRmPyLDuFTzl1x2ItVjkgJ8wu+
/GOFylOeUFh44Uyj7/nUa853A08k5JulqT7KgFh2YZsKG81q4pRioH2CndsHqZAm
crcL5wR8LfPDkXmahRWfefKBvOwRlRYp5oxMUmujv6eMdT79WtAdkpXnafOxxJlj
Z1vmfylP7C1MAHl8RL7we8+BjvMS1zI9FKGaPbxEnb/DtGN7jFSOSTbyozbq/NsZ
iev5xfH895i6Cy2u4Rm+OGyMboqsvrQpKrrQOaX5ecOt8FsO/GtN5ZJl2Przdr1i
y71NRiAuxyQ7p6+yyNIo+z3UCbWN7pdhVs7kI3rBYrN193qTWFjiIoCj4ZCruWje
Z2uDEuqGdwXu+b8pyTq/LNHBpYZP/sikcMeejxShbU8m7AEIw7eDAFUJS0W63pOI
ojyZVmZHSMA5+Dvszl/QNSTicCmRj7KqgFJk56v7NRNl76ytptcKtl2YLx+oEUFz
l2LD95Xp6UUrzCTFjcz8+HsFJq3xZowJm5O0h9GQ+tOiRA1hEerHlSssMYG0La4A
vCFM2oTLzuHOcnDwuFLiG92eA4h7+zpkdYvDua1AOg3f356FYrxmiG30NM0MV+nT
KK2COwBvZW72WzPobhI2A+uIxWxcfAgNCzSrq0LYUhlw9il+GR7EacJlTqp7pcqF
9isFGNBXS4yFi52Jc0QkYuZm5hZcB4OxljMH9sh/3RqhayNp43/BuCOEyJqByQTN
RFIZhFSOBjN/stvZGG/pCjuSHDB6TkrSO2aOnrwvBOppEebUSLLzkE7QXoZ7V5T4
Yx0hEycQk2689dwGrMO9PtGr5bjkf8ND1KrS5zLFkOER+SoGVNDYkW6vk342XToO
r7XqZ0v/XiWScp63ne7tbQ4e+c8lRrUwQQ2qM8tt4G8fn5tDxJivfsG35G5IW6KU
pIZdRb8TGHbJOGsEjYKL7vRICQzeBh+HT81G1z9bsDSRUuLV+Hia15SximLtENNP
v+UOnSTssenpQeCYJ0I6Qc9ah1NSw8teZ7vaQrAMlGxIWsZZM+AgwnGGptFQkgxy
3W9dXl/hNpjLRPPiv57+KZrR4mRujHNmii2HWGGndSSc+YuDiR+V6o/TZ/USHHi2
NOEAfR9ZrGstIr/E/iLCoHZ1NXgujcGlpnbTaTOfWiXpqKgC65K5WFU7+BZEx3OG
wmEq1YSDNBLBor/ooh0n9/PGbfUC6HFtdIq+MBIgP/UclWNHWBMApABaVAlrDex7
sJ4Eq8dIETYmZw61U9fHTRPv6DfUJoSJ6zDpOMdf6Mbocr/N7SE5JAQPWtvfD5gZ
IDbOyCD1sRoYAJ8nSn5gPG8dcIvFQjTwwn/TDr7uQ1afTlug1o6xyHW07nEVI0PW
ZGzs7AqMSCUbXk0q95G6dp5MyUNzCV66D+QnAlZYtQt0BRXpnNTE61CqYwDK63mQ
swlpO0TscwQ0SoqpnfRAf2Vo1pmTtAAlBds4w7S6ygDA+mu5+ONRROqG1uHpo+2H
t8arZpncFV70h21wsXpBOxOYaZSD4pkVorZp+Ut/4VTYjPO2Zqh+IPapFnp4XlYy
arEtH+rQuLNVFgDtz8Ti5i2NmT/NMiIn31GyjJe1OuWfc4ScsQteEB/zcHlLVpn/
ENeIZ8RRDxUAq74FoVUU0QQmENw3ofKg776UCfabwNRShsIpC9KGKjc7AlXz03XN
/oiwwZonqNbfLer6F+iK+8KDe+NMaychQtJvsXz3Dfin+HpCf/UJI5Lmzizpjy/n
30e3ySJRfcQITWfTeeSaXXuGVtSUd80iaF4B0RoRJkCNnhk1DaSlGePmEJqoiWeL
EjWxm/cnsmhCRUuaHNyjAA79svoG5itXJ0Cpj29Y0s9d6zpmtOAtlBtWsVH/n1f+
pkkUN3kTNag43s+/n8t5XOt+dhp6utinoIsgk0zO3AbMjC3U+KxLFeHvoG1QW5Vc
KDFMqscOyi70Hmzk7ywE5j1L42OxhyHbxMXfU0ZfEg5fLIuo6MLajEUAFfyXpppk
aCSAyjP6u+two7iV3dNYBDYUMMvEWjHpPrWyOqsYXrBHGgd0zbbZaBIuX9UoCHaZ
Qj7+PJQa0ZOQwteYtmBjtyFergrPbL4fJC5fyiwS9nICr62WEokJqwbQz5YOf5o/
iFZZIeSMIZTQMNxAU5TEMsWr6mQngUOz+VayHhcH11XbAAUSWZQ/N5el2Q1ygbzV
81xy+XYRYGeOTD9TJZPXToAzER4zOfWVCxtQCLChFykNqfk5BSbLhd0m+/KsT5zW
QysVFgPIcJpZGR27uijgch7LniiYbAwyzsHGSRtQedO0hf/HahWNlluUYUjKd2cp
HhRRSh6bMep4aSOzc1pRV2vM++RJEsC1VDelS0T2/44LziHCS2ui5cEOD53sV1US
RILpiTwQ6k3u4KoM6fh/9RuYu+Mgug3DlUdTrBxGpXge1TCueCgHDaPVx2IdNS+r
LO84bKGFtCfno4gdXRHRN8o+YE9x9fB3yRSmRLsyYwNFQs1Def7XusdL7gjFN9+/
gKKLwrWfk31F8wk2ztgeAMibuJ+OrG0WGR1mHmAxtOdZeuj/YrqM4JECSAQ05CWZ
Zijiffg94iC+xLFACDNu4Ablc63zB98zHNLAzL0dIhiHMza64093ETm3yYF+ad5R
K1yHOcFg4SjuuEMdBQME7yFSV5AmdelrDHvd52neEhWkxn/Zc+ADic6GGaGjuABl
bVcUNvEiatcShOFaZmpQ5td7pDk5yiw2NDhyXe56Qi8/6AGnQt6tvLNAuqYN+vnA
zAFl35/lLLXKloVnExTvDpbZnpSC8inmxjzXXBuZ/cFdz7Ml6V7wT+D1078jrGV1
LtiZiH7mdkP3fmgHPy0hBhMg/lislPgBQ33sRRB5wSAEAZwXskjqmB36iV4rJPIz
sVF1ZUzLlJDoJUitnxkm+Sb2puWsBVfx2gwZNNc1cJGDsBMm/ZhHwUvE9X8jaHXw
yJ8E4HJkAmK8S0irVkCWZGMRI2NoT+xS6A+WOss9n1MEObrJUD9BWcG33ABi41dU
M2IqAtbPc6tMuDKOdG1mSr990vHShW/YMUdHeNZoBfn/Xw93PrckboU+4W1waN4q
JqOpuPWRsOUa2fvQZ3NUqcdD+1dUsRqCDtrKRIxuzC1HVnkNirdhpn5L7dGNpjhH
9BF4awi7+GcuwHt6X1MBbhJ7YSEz4TmUUzJr8VtRZSNCj3OfJR2ZGhaBpRilLM9d
1zxMrP4wWe9ZT0ZbIZRa46vLw9L8WZJWO6B4wSh/eAMf4Gu5Mxd6JAcBCeKNUIAX
EMkXXeOLq9IDzX1w4tLeAQbDkPqsxxBaE6W6gxbSgYnEzphl5G2dIaKZfgOuZDxn
TMRM2/JuMjbIytABhB1575j8kODQDsjRXgxYVR58sxBZP2228qVk7W0L6w3TRqQB
1Nwy641R6YT74CtjgPro/i36VmJGzQ9jqq04Un5mNo5IIL33zW5tFmBWnksKQnhu
qHBJw3kh6ix3I8ascXSIbQpGlzHpO3FrSLbAhn4tDHDs6UmnC9xuJqN/yQGtHSbH
oq10OnPSvGZT3XYXLBXzzn241ju8rWiAFQIUIzZ3BCvSJFyUNdqQplE7Xyml4lT8
OoDtENEC1CArVL7bERVHw/wSspV0qbZk2K/EfF2iT2G3ClmeQ2pfRFj1nhKvsnlz
ZS5s+p/p36YR8DWYgP0xwhKDfcKcxesC8NXdwG9lwb2j3gEopnk02AI5WNQMvEHb
htNcHe1t3W+jNhV4qy8AuZLY0ek+Pe5TNGMGuQpLLljN/hN8I4fvT5k+QCdlc7R3
eILT2GrGJLvJdHdCvWhfnt2nL6nO4vnsISfKSNr1AyqNHZjQLDeAjTXYr2eU0UXy
zgdvXAaIM5IkuQpbzoWv6hBb/SCkUXk1N7PloA4GVKPOyX72LIaEzwvR1JoRi1y+
CtBX2nCtslXx6ZsahCcLbmiHa7DtQfZuL+rzv7uKdPpME7oMZ88Y3B/dRL4dOMp7
Fhv7rvXwpIszmBE5KL8w+MopNsvd02sN9+DitKAOXW4pmF8L8jCz7zxIe3NRunM8
n+36f3wzXavW3HnqmqbW3Lk0E03KzWukFaV6GflC2Yzuk013P55J+PkRFWQ971KI
VyT2k8yVlwckqZAUNSJj6PmAjM5ZNF3aBQCJgoQ/+2ev8bZJ2erNnk43SPQq6nYy
0oF6kUda1zEiGGobvz8M2LgXfgBJrSqVRjfdMoY6JMMjOh78wbCezuXQLPvl4je3
bio/3YJ5OQoP/TSUcsob2Ql9zBXP/kBnpZf6dQ/HSkY/LrzKM+3kFWmNYIB4Pg2e
3NzaiIc8yuzohVJ8OP1B0789eZgugmvpO9nD3jtMjDFYQFKihIJ4d9994Kr0q7SY
v+9GRBQaGELGiN13nrJT9YGYvupoVBei9DcLZpuz3xUZjJTe40GeWtHYB4Sq97R2
J1MJQmGxsEVggfc0QMRrJThi99tYAo2BvB5mEsHgeh7Vdn66NNYLfLLP1ALiszU2
bZ/4t+54StnZeqpEBY741D5kxPeTz+3gM4LZShebR+MlVlDXKjsHLKPxw9PSHHab
XgyFmsBdiKhTnrloumGrmcd7++rEj5sSOJBjYYeIK57eXY/y3pKJpXwuI0B1nKye
4LGAPwpaorBzDVlEHZASzhEkOZCTmd9JX1EfZk9ECM+6973qtPWgCQD6czbSXMWN
tQUEcIDesfjKK6FY7/PFu2AiXBXc8G0gHWM5JngmzhrYvjncovWrfr0zUDhYRB9p
Qu6w9DlOXQ13HZnJhA08m3dpunzCVP65Wuk4RB6mrqlOrvYeSdn/0jOIyB6AauK7
DnuXgTsKhgXqmm8Mrc2t3R/7HfhaakhHLkxhxDIPXCxYV5kILrYED8m8yOYWbZCX
7xICkFxChmpVKy7mqitLeShy/oKJDAFJip5rP/JTYTnbJvXyTJfF0lOHHAFpS/h+
KTfl+DyAnf9I/zBlmJSOGDOeyDs2HWe16xO/g6AvX6LnDXTR4YtmHefQGouhq+yd
J8Gzqc/j7QQbnBWX+K096a8b2GCqbd/4T5Rk8EGW2Ku4TephPUwZMSoGiySZo82I
kg2GmY1BmeHeXD6ZWqOd8lziOScrISX+Lu7HTu6+SX1Z7o3IYhXJXDzadg3IYmk+
s4OK7J290BN9BJsZCGLpepVMd4GITMxF3G6zR0xpJtvbkJOu5gtkh0qWrJTJZPbb
WRRfcL804+u6KAU9P5jToXDslDxTpOatFMm1c1Hen5w81iAWihA3U180iE6DM+/F
8dxLceYSSS/DPwNM+Uci96T7brcE5EeAuQPHfKxWekB0HTBX2PtqnkgQ7xwP1YEN
QaYplr2U8yq9023xPsyyvpC1lZsME9s/N341bxAhbnYfLEBzj7Y9Jj7shXinIdK8
GNkN/BdfB/z5+gFbAeNl9vzXlXzAKjKzKARZNR8JJXiDJNusIMmS8zaIoJf9R4Xt
c83MhNOau/wUpQBQ3W3gd/dC0cTSwya0MSWFv/hu3/RAE4yQ86MFA9JthNtVsr4L
e16qAKH48TcdYcDX7Ukr0FBEx86fvg7xcr2TepWlWY0rY+iGWGY+Gazc+EGcUQUZ
dJoNQyK55cN2bUAa/MdapCH53wukJcZJ7s9KYCVwXi8Sf4kO5RWtuCNf4y8zzY5Q
CPYs7oKmrHmNEt800wrnoP5Km5r5VnEt2cNEIySxCCN8TS8G5Lr68N1wdSJo2taQ
96Zlxb5JVWXeQu4vnbcC6wNDf+7Guijk71e+XwXQ7eKRbDXSk6dF5uCUAgvrVAqc
a8WFD/yPKr3Q7vSRy6p6R4rtxGInFbBJ9XCSH67aczsc5aZs8nwz58WCIxT9oadj
YHMDrS/0tyni6LsD19rYJPsyGlS7w+RH9Vx0f8eP/u5lFDdZH+cU9kV5JuDWVB/9
vu1p3E/sAaIfzfbLmcD0Z/e3235WP+lDEgQYdGndOpNvZ1cDBqzUJHZivze+Ygvv
ifpQQ9V35F2+jNgXtl/z39I2r8EgRyJZBpbVxGSrwBIRiRvzmv17c8ITOiaC6q6K
OXVaYKqsHwDi9ZJBA7XfDENUwiriTwcbTTYJKg50h3RAFVs7VH03k54Ix6d7M7cj
yuIEFGXMmT7I0cnti64A8uguOVYmTV95zQ+p2ZEc3aSSuAMPJZSjDPLJ+WiVc0/o
zBVEC8HtEj83ShtzwzUYnh5VCV/5afLRRgB25vv+qFPk/T3Ks2NNKwYhem3AR3CJ
M9sJ2bpY+8BodjLRM2zqWKcDCi3ZFNMRE5Ve22WHQaLmzeo9u8uh4L0U+WuwczJJ
P2PotBo0mDrkCjiDx9vafj7A8dTv17YKfebmGruM3VdlPCqg2jwKRKBwQCMH8zEX
8x7sS3poepsgZyL21FxuL4sPDJdAzbYqa9S2Eznt1zkZaJPepp3qv+IfviIc7sn4
4O8FSN0C9ayv/XFCEFokVYLA6oHamC5IdfYV5eiID77JogsLnY6ds6a8UDwGgO3J
ob3OVLXw5VBxyz+XX5mctn4BKYMLIPc1Y5lNMHd9LT72c7ksSTD66tZlil9UZAoF
pzOKVwG/cmEj8p015EpOZ3Z/xiSDHKdJ0ENERIDvfJASpH3A0NmUYIQ3GQWli0s/
DmCTot1gnzHuTPoGBBDYkm7sGRJBPkhXV3czVaHMiBthbAI5sxnrsufPbVHnQJ9G
a215iLBLNFGzbUqvmtQC7n2AQ993oSboCmoarugKo1YMHZ+NInkD4L/sCZZoS6DX
B9Tc4JJp0Ba/YCjoSVECXdzXIKGigdtZU9jEch3PqwdzAjI0EPXg1BIh+jRw4H4N
MW4Ntc/5Q0AKK7vIblbwAUlCnYxUvl8F7RNoHP5KvbR8UuGBx9RNYkB+MsRm5Cl3
AHJafuwsha0KhQTFEs/WNIrHeBM83RZO87NRFKnP9Nx6waWV36RICQ9CnVddw4dH
ztXYrIskskaygL8CEh75UkBaBinW6jdldbtkwy9q8uqjYhJlpxhvy+3bLL3iafmt
50LvE3p17tFGev6e8yMNTpaAYAX1yiVsErerAx+NE3GMz2477t9HzkOtnsO5jXYo
IFe/cBKbJbd1bMjHiU5IW4p8DYdVlAYrNKp4S8x0VxwND1QwdHMtv8zut505qAIV
XxrV5dBotf95c6QTnqHw5ZjNJndg/zdchFolbcPWZbv4cUQEIij+OVWQdZ/DYAcZ
srImgHNJpQvCUrJ9V8iqNnUmUcGNlAak6XuhWWRrt8s9dSyjgI+UhYLp31xjIaFr
iNNzE5YQD1MWLw1ZJQL8Oqmjiujzo+wH63w+tpzApW95XPd3GilW/k50CrR0/VAR
RHohfycCtlINuYeElAq9RFD4ucIP+sEZzsHrLandghErOSSjNyXbKGAKk3Ze1I8M
OuiSXwvmMj6YdiS7oBug4SJsfxpq2wCvUa9K/dumkn3g3sJHXK75qVcB5zMP2eNf
EY2ubnG3OF54XwaUkOFAPMnQB7knj7ryi/dEk1FEs2KmBLUYiLCqvViv0hHVa8OB
tqHqxDXfld/lIDgt9IkW47iefJECsSLFa5bC6rfUnD8eXS1yLHItCO7mTPzKw0eE
ikf1cu6Fahk2GCCq0hnBbTII2R46DqGGAKubIwwo+Xb7skOUzKMmJX1zagAUJ9p9
S7u1GSuw1+QMfezvJSFGGrT+T+3ykAkBHyi3zZELEy8EmkxVd+VQ1SAEHgentK5E
WiIBO2HEGlKCQQ1KDxx0SXluEjWzEkpQSdZTB0VZef0V05C5YOTowoPn6AHOfXvD
TVZ+/pwmSQvN17+xwVySx6ELox/uqAFBrfKVCDgwIVOWMjKCQO5nZIcVpUGamNgc
fAGBmOtsu/B/uLDGMs6zgs5P2+tSy0LMQdwedgMvmu8PmiMwxeTyCqFcO2uGNokD
pRDmLRQ3TxA7HBh8tudfFcED6xSQfelHvGQhgkosKSPg17EfgQgrJAvS0St79OSp
r8JqJG2kFQTQPsxaO+XRuSVJKIFEvbF2vx5MXbOYPyEqtu72gmiMk4PP0VNNx4K+
55nWYJpYfpy6KGjaMTCB1QDKlJBXykJPfxOXpgsr+zZXrhf1X/jKmuNFeUjedjOG
PiIvfkmIOkeAgAYIHVB8uXymW8UlmxZ5jGcf3qE+gmm1S3sFV/wHPu3Zk7LcWtzY
621Ro4r2MLV3oVqEoccBX26iUjPr7Lp+JHsHDxNpm2gGcR4QGPoRgohMQTE/M4WZ
l8XGNfTWVQ5cG5v78/baCfwl2d7PIjaWvmtqFNzXhMcn0+Z6vm9djwm4eoIvaK26
NzC6h7gMV60TxmHAqzHhlDAhCvnmaubLV6HdHed0EPACtpavUjqZh3a+5A1MK2hV
tC1sjQTYT6Iw3Wb+FSR4MqAdZofo5s8+n48k4kOu+qGwQIJzSgmylzg6I0U5i/l+
SVYEMvcS+G89wWhBXvXwFm58qPV5WHIZa6cYrrGFuMEMtjb7Quxbv1ZQSLupKXuF
xp/c3pukOMqEDTLM77k6M3D9D59Ax5OUJTwBsTajAppkCg/k29/bCAKq+WmGhEVO
ZSkMA39z81mQYTnvRI/Wlk6zr3fEKga4cKCOb1OLtL3UrxXuDDiT0ITmronwKiq3
+SMuCZoEZNBENEU6I4ic2giFq+XmIjH7fOJfcnPfOqAz2c/8PdpjatL0OEMHHVQ9
dtRLBaBMc8HWnzk4Rwg8LEQ+B3WXWx9BgK6Xlzhpy6aVRZqD148MnNBQBq6sVAOo
kRe7LgSNrtBnkYRmNvHsFufop7pz1ZcHb9yaQz53GOfZ3BrXZmGb/aGW40XI4ZXn
C2zl2CZR1tTT4/7GBfoP6ruIkQA0zQxIrHvpyhLF6kNrMihDVyTLRivnKeKipZHc
Etm297aIpVLPpUKXnHmWkphMbXy3jr81arjR/8a46yH0d4j5O6ncAYsXTZaa69ar
2Ffgr3p0/40TxDjZC0YgHLOpZBs1w28BlvqKr74+qJgs/HgfhDwNrS3X/eibnRKY
0U2J2W0RyGJ9ulucuNWMAZFOgLYtyhhVnPZEa7xKGQPkXIvqtFtOrSBcC42M9YLY
D2xl4hA/QItpVAT+7rAwgqOUEypA808c42D3uXdREPBvX4EzresFb1gRf219rVzJ
lAJqI3uC3cG5QNrd5+k76PEXcqnHvyiCVXIb3yI+9QIhYVmAcnuQx5aV+18gEQsI
HAWHZaxTHhhMkv6pWfBGhUQ+uBC8AmRLFVAbP2byFFGo6ga74+76VIRvOqRgX6dD
q2tiAMR6VscYKQEmHIDF3ImKdeQMGv4EKk1Xld11W+0HygylkfK5I6evzChJq2Th
8ZiXaLr6i83MZ5t07QOTIKi0E7lJ80If86dtgwi9dqsfY3L8fBmAVeboDqxYByym
Gr8sbg30VYN6k4aVc+cpgPM3fj9guYYFiQLtTdhF/NMMayN9pgG5R+xK/L4OHziL
H0YY15Sx5I44yAm2rCiAkhKyfMNveIC2SdynvqXo1OPsSaAjGlWjQFE6BgxCrgc2
5Motocmdyk2JfghkZk9sy6u6dhfivgbiLpKRtGTMa3JNGboQYV9ut2N1/6I0QcFB
dOrnE3FAbYZuekTPqLzFEUa0DmjsgpLzfOyUODKbU8pKbCt0aZc4KKIlLhzIAB5x
Q2M+dQU9Pc0W96OVbCZtRBX1JBjs6LDv3ancNeVjnvKD62JZSOJela+PCj+crjWZ
5IYYeRYAvWHHNhKZK5C5uGhXUsuvMyFi5Xq11MG82mQmXWGfLuLRi8y7Av+BGpSW
6Ri6Et9Y+3diW7Rh5Ji3jMApaMmSrX3NhVtqB4YF8nDGCrJwPBP899e7oxy+ehjQ
HWitmoB7ySNK9311hM/HwKQoMyG1l6aiUCOXToKLTOI2at+zN2erLwArV5Xl+xWj
hnDScBi4STpLhLyJaV2CofGV7CrWIAzYdyGdIT9TywMnqu1COuK7DogvDpJAZvZE
xjHbk9SzuRKWrFcpBFcffGGwEa5dRqaJa+FHvs82Yb934/LasXbgxADtDbeZzLf1
Vcsif6/iD7sRb4qQ3CtD0x3cAApm2WNxYTxybw19IArA3JEWUjXHFe5wU0PiwrpZ
M9fVgRRZr3zvurL1sJhBB5wzddAMgpJMOeWSXjlr1d/jiKbZxzJCeHmETDBluO+0
oSgj1UyQjs3IyyMFCM/2MOex4iokxXwM/sj+6IMJo7sz1+7lWAJWsmE8V5jUyShJ
jMugFhqJPYFczCIcxw56sBjv0kZ1WhO+4KhRqlb1eRntKL1X8gxyD/O2AErY56Lu
hz2e7Tp7HhvLnwPCjmmcu9EE09+LzIYHbM5zhfMDT61Vki5lE9h7u928j2aVwkFR
nLn0ksShM8qi2DV2OHy640MDX9O/9DSWKVuMJFQD+txEzAgBQo4uR7K6wVZje92X
OdFq1xQwkkI7corhaeGkUllZwA1zty1VYWwDAE/lhaJqOaoQ59JtkjkZVd3a0U2o
tOX5SI6hHBJ5LXUy+c3i4BwEiOlTEaXaPPQyKWD+S+TlWR5RuAzwBUxDfv5CPqS2
5cPYcui1m6c3jaPDKAv61tZ6mu/HQZTbN8c9vIKquvMT5srIaTk0wuTiKMBY2/gt
dVWw3Ib6dkrvScFlEDobBvHGXdaH59RZbHLzJYrsBNP1ZLFPpNAaWgOwNAURELCj
wq0bumwPL+QdrmzZLkxdOs2S9YLAfzN6lRfjm48G8CcBtJ0iLy5Zhsn6z4h/w70s
E2f9tufLg235E+LRhx1NqCiDTZdsIcmMjFQohX1pgq1hg5iBHztYY5+MBkQ+w6bk
cu1XinjIGpSXMVBmjIOAbzSA9o5J5TuesJMoeAEniWBvmyp9x6UYxiyRHRgBfiXU
ydI3bzJvrScp1X1qKF+SULTZUWGZvjXI59iYFsrFwXBI94k+fSlyLl0qfdMt5XHP
+8BI8G4ajYsYFXo65Yz/ed1/LLtGmMQC+4xJYHyXf15cZxdrOtrXx9EbQVxPr9xz
N1e5NYStTa5E+spw0nEdI/Ri4FCY42tckbVT88Jnr4UMT90uSs+Zyxgu523pNycV
T7eQFFVpRDj+fvKaMmAu7GP6NIS+SsZF/6uApx9N/zhdTSQhl9hh0e9l/aU58RJP
N/1ai3yHVtfvsrIHRichxKHc5wmrHDR0w/Tm0jA3JvEXnQ3dUr5V34LRDkfq+JHp
sXC3aOobNd+TxB/uNs64Q/tW8rYQPG1UbvzYr/n2JRl5yy2IWHofYY2wxYMBusyS
OCtZf2ePm+RNxcWvuq1yA302GVe01o6YPwFNXM/vt3ZfjMycNCZqtqKYS414Sbxe
MAoSaCCfm78hsFDB7zURc6zuMNlro/hSeXfaGNHMCaf/aLrnquxUPTaiLpbG/Uy+
NVPoX6M1AuzYQj/LmSYwWt1B3Gn8ZUomNh15twCGn8f6KA0lqhhuSZ1+9UezuwyP
7DvmkL06EX5MX6Q6iNeqHr6z3U9CCzHo8C8E/f5ahwV8lfWTdCcBMebixxA2MDq/
rQdjdDlV7mykoLC1YL2x+Lcrj+6Z5nJcuPddIvh2tL//1YGi3Hs98USh/BySasvf
XV1a8hyGDSlrQhZ30ULoA26QVhhVgR5xmTewmCARQnrfXM/uN6Iq+jpRPuwGj/JS
EuIzrvAEZRHUeL2z+CvpY5AEKgxNc0jqHHYbIrFi8Apa0M2AsyzDnWHuY1/MnNvf
8Kv4hSQC/W7vm8dWNPlFwFDjTMePZyXVhkmXFaK+STI1AVFYjHlUsJ4uAbgvGfDd
Qw0vsFR1wpW5sGS0kCMPEw5p55+9lFN7dBBN/SRnVYHGsxns0yo7btqeaE+MxdHW
E1/xaNHdgEzeQTCwl50drR+Hr0VKrexWHrOVEnk++iVgSayE2qjKZdMaKzzUz9Di
DJMZQzHxFxnw5BPozWwUKax7epJq4PtfFCfeDDrzEe8E3qnl/rr0oGPjXIKZotff
ynFlptj2ojF2GRmMYzRURnf2FshWYpTt8cdkIAlH1fBh+hgWAcT0x401CToeDXk7
JKhiZTBvA/Qw1uZbar+scS2D8yp4yl6QAs8ZKQ32tJqjW6ivU3SKvC528RKgcCsF
hbjasfsbd8eHGRdp30pdUXsXugtGuW7xqIaLrM6okxG7/nJ3OAQD2X/xs2jjbdpU
a+ln9cQb0bg+qS48w4eR0AIBF/wp9+Kj5gVwfjrlqx3if5e9qyES09RpvxzcOLaq
C7mf1LX8RRR69p2E/fLPH0Qd6cIOXLCnJlr/H3n0BXHtEMqIGgu1OlUly4VNVZPy
mA2onpMmJQJEB2sWrEwkVGbnoBh1CfBACLW/51rJzcNy3c5hAUOUj06y+kJN8uRx
Ibd+xucU6214Y0TkMSR/rmBJTgsGU+XvOeITv1YVC28YJSH1pWOVaMoa3v0V6vtz
jF+bzebtl9gIuXp3IMy44+oRiV2W9oUIhwkEXoYGiY+kWqCUgEbFAOCTbOm06PqV
VRLv/n8FHN7IsrARFH9lOi7GgwWt0FutNTrl3Pv5p0YmOvYP85r/EmnEVkZOpqeX
JKMJpH/aC4PpqwdW+oOcHo7itWhbJAS0GyEVXICzUZGRt8USGr9RgNb/4I9Q2VIF
Zg52mKF131g+0hJTqa5fNa+UjlDIE4OL9gnlbipfO19IrVzAYDC7Vz5m1xrWmn9D
SZ8m9N+k8d9iw0LbEUcyOfPKcTufqlF4nNSJ8LsNcYn/OQMgKazu6JEKzpJ9HgLD
MCMvYU0Ii8po91xYffPcPXR723+UDkChEUU/EAJFK0JxgC2LUOEAH83szit7znjw
aTr71ElOgTFzp1kAwL5EsRZJWi5P6evoAAYA/MmGkGCTFpyRyp6/lpb17t9PIc4V
9GByBw7zCd4ywBNppn6HjxpcZr9AZcK0BBVAoXnFh5jabO2WPiIa8PC2EK2NWeyU
+qfOrGuMZwBrbtiS3gJXE2gN+uezBvT8sylQPYLKLviR/XvgDRnEl4Jn1PFYL/b+
qYSsJhvNbWr/kR0bFVNC1LVegXGdGN8ReIt5hIlruTP4evIpbh7cDd3JdljlaicT
tW9+2iTLC1qLy6Ij/UwN3Mngy8asdagoBS3VWQ4sjyj/e7NkDc5peymvNLq3Ukir
gc3878eGsfacyRSPJz10yweyNCCiQlN8GhXUEM+VzkFPDgP13BxVgc+53Ah9htni
Z/Qzh/kMxXZmESo+fEmIRKxJZXvBwCuM9yFD5jL/H+QMgqfj1PRIiAMXKWa9aa3F
2CixzXvLxA3BpUccwD3y/z+TugqrWZOajknPiXYp5Jks7CRDpRmrwsYWNd/5+C3t
NCm2W3ndqYiUHQJt4dTvR9k9F73kLANfvBRc291ggg7okO0UAuT2c3QCSUMyTcnc
yA2f2+diMQuQX1c2z7Cv3Nqgu0IF0LltdYW/ui1bUBk6C+c5GvJsN1TIV135atLP
c6FYkToBNFKgzzC0sQCBsl9ZrZJhmj8YGw4GZTWJCCyJiAjxP3f40ODAHI08cMTD
xtQEra24ydICf+oaho01BhRaks+DmATlxADZoqbWmGRajs/08wVGGGnBs7bAnckm
ksRNQqYlmLm+vs26sxvTTX+b6oRejnFrVbljStwbcRIAOPiag++BpKdUeDJO19O9
Rl66uQ14YWujuXIyBd6P1Rvv17rM9M8CxQ07u47s+6Odd1Ww4x4nWNRFFMbIA4wo
DYGz7HLGibwyD9YnMESuTrIAGojuL6dxnXpeLLzF4lqLJr3XOnmj/uFCkdBw1yK+
iwcw83PjObYblb3ZWDRMnPtCpu/QszRo43EwPy3LJvlOrPqRlUzYjRyOKjzAKxBb
+b+KhE93u9xA/HvKNZPC34O1fbMJh6dHnB+yRPl5qVtQ752WX0Nc0fgxyEJiAh1T
qN6vmZOnkgl43Xs8JHPaW9s3JFcAZhJbwEPbBs23ucJOZyOnTRESG83Bd2qtrUJ8
GKyJd2yjBkSKIJ0vI/K7QqootgZRMDaIicOQgYaoDqIbWO8WQ7D1Ezu4oiydMQMu
jc45ZvXl5Y5jJjabKvGkYyPhf/1zOQo+MyHZhWJ+yB5JuBZfC2u6k/9Ct/048HRa
3FvdW4qxOCma+HvHLOzkuWD/N8+jTL5seC7wg4zd7HPvhTfmWbzRpV2yaffxPONs
bxawuYSRoVpLMqUAWn6fr3KIDBay1S4oxBV0lGVV8MuOUFDVtDTElqVkbUREsxIz
VQU1ctXk4r+2xUtUk+/1rkBSE5WiZyPMTR62sK43GmfQ/IY8zpkwErKDAiGk84qe
3TwZE8GgAgZGw8dVHsw8biHMsSHEgN9ajR8+AdUiG/trhOONE1lGXawXHcn4+ZpI
hHg080aAzL4pst5YdjekoyQ3GjY1r/uqvZMQws6zDqCX+bOjD4V0Kfbmw8bOyZPS
Fkzm1U7b/3NmxC9Pgw21NXNrr6obWESe2E++O4ncAJGOk6ooDIfLev+1+rcErmTM
Q4nJvjpufqWTJNuCwLqDlavm7gVAPYM7nwX8OHrVZ6b11EG4qXlfZ9GY+3GkDez4
uV+3LcTZ8JOj8tY37mMeh10q7/6zmH49m9w1h1Vv2AjpYta8cJeRg25vIGTU9vSU
LC6tPcw/Znd13sOHiobT4G+NotWYgth9po7GOjqtH3e8N0zzS00ARz1VjuVmzET9
+0AsO1IAxcYDm07oKzYx/WPDQEQDjPCnSLNkxMieXABYV2pawL/+gpjAgdccLGMA
N+bDGXFC4kx6Z5okLrpijGMSxyO0dEWK79v7hiSexC7pgfwTSDjqy+QuIQ1jMPaS
FZOjk2R66e7Mlnz8GlpON4IityPfJbTxQg3ml2mtJGqQP92YWkfxjtPxNS3yZ3Pc
WPXuWELNNFGgyeNX+KZEI0Y5NdS7YnMIvmVYS4TJhGYWnKsCWPIzqXPoY3TX7xCO
R6NwdyCCIdtgANBXc2eQe4P7czr/iKt6JSwueSD6XwIevcnb4yEzoGG1UUpEvRQt
iWuqSJ1MgAvyagK0Zo1uhYYOdS+sUkGiDiVu0odELQypOVBUrZvYnHJmc7fRIxJj
yOzZyzJhRs3P8GqximHTohg9qlBdVRHTZvwQ3PnXU08kdli5zsTt1frRhhco5Pv9
E3B0PXtrlbxLxI7GagsAOfOHBlEja3HJbL2jX0WfdvKc/wwFoMdbFkE5r+5mrRPH
d3lHkE4+1tA5JfW7Zgz7qSQ4fzjMf4rN8ZKXNeABGNCgWvVbhe0cQtoUob1LMQ8w
tBNTLsKwt6XcNQS04I+a1S3MRXEZ623u4RukXooVk/QArZQof7V3kmdcnTfH+Vnu
vpajZ5B+2QCfzhsPIygDTMb3bdFBYDGvOu83IWa+I0893l5xk+jL8YP2bE9aRcGZ
9pG3UB4uS2mn6Mg/ql43vOmrVi1iNphyNLIYA7E859kjF/Wm0X9CB0akG0SkAXfg
QM43pWquu4RJj50UJW6UEh1vpJab7w4IsyZMeCu7fLuZqNXeytEO9NaS2BiSo2TR
yfYzb/9bz5S2lyujS2tYrh9nrRo7NZQn4v2TPPJcK+DlOXpnlCyjxp/Vl4grSqbJ
9pmamJyrYj0F0efijmMOwJeX3Dfc4HSa0pipTJUt83Gqtsra3GzQVHDeKZbO8KzG
LBC6PSnAVQDZkjNdLoEhxf1gX4G6oJbYa10Dyydd/oyqdNhwZjNdyn/coHSJq4ct
1HA5y8SoRkFFq6OV2cmMWG0iYKUDFiUlz1jZw6DpqDPJ0pyQJN/fW9aFuZmBYDIo
jtvBZ3HRZajwJgr5bj8fsBh0LN7dE8bXf43c58tcc462YmN7fQU6+yv/fChBjH4o
KuybfKoYfGPlJq6uCpUAlU8tGQh5+mqwz9+DxpcPn5rJCDEx0UxofPJNDiu/upEJ
K2coAYVdLJ+C25xUcD/OfDjAls5mvT3fGCrjg2zKhohnC+kA6NeBws601V00VR4c
An7Sj/y+Gunfis12U9yiMBI2ov7aWlzUa0cXA5jQ3oh6GszpIJaCVTXikM8Cgohs
HYPzsbPzYklGdAg3pBZEK+CJrranBg5H5IC+0hFd5Vq9XgT+/HSHDrnbUEwdsMHy
laWw1NJe1ELYjFoXl0rTyybpF4FDFkGg3x8nGjrYXfHtitud0nWERHWg/t/bc7Vx
V+SKO2rqn0tlGIRi7lYCvFXcMQHO0X5dAnMMUFanYHQIL4COsp/4rCGAPBX+S8Hn
Iyf+min3xkQCLIXxwlvrg0NZ+uAo2K2NQ52+NsILaqO2dgVe7pXEeE4DkJgcQqO4
aNcWF2E91gqdfwD6UdHTI28aqzlfTzlcplBcJoGSCk+uv4WO7AkG/7ejPCeU8dq8
NjEMEQ/WQKhdfH5XvXpr8lUUzin7fDuUVtUTTR1L7j1LRrrZEfOsnzdGY7Oq25aR
CG0XNyY1pdmy4LNfdiXjki4LwLKxBvsz0EMn/0tmIILl2cayD3s4ej/Grv7DwLIq
WEmzWw98z6gX+3g28MJsNJRVnG1UZty6VLpS02D7gxDuhEA8OJVw9+MHK7q5pId+
W5wUT2d5rx1hmGvCnuBabuXH41OO0RTB00KvIRhstomVCOoCudSuNHB1wW9LSGBd
hT75OWskkGALhaDLY5HDQA6vB4OxpIvRe9v1X5tHHa6WOhqfbIbjUkLgNfvzXSMP
WwrDwQkcu64BynoOhGeb4cKubyoeGFJ1FTwTQF6tpsSpBp9bNEu0iEGJEcD0zvbh
3dHsjL7BQVk6jf9tu9vJcLHIUvM9/EfcWQAxSzNjcNO/247gprx3VPr+tjy4/CjO
fRrhWwEw4QJ6vgoGZO83xRhaA4pnaW8tlP7L3yaCgas5rN9sZb8p64PXd51L8bT6
zTqDEb9i/LewU75UZkMrOWF+ZmYGM773GytqIOcWLUxfGn7gsQmeYNYU1gGCj93v
0081dOSzjGcsNNqgJUNFTfeRtt7IvMgjCq2+E8bGZ5YduAzPWJMY+s682lTv13Gj
qCC7PReZm+A+kMJukIwj1CEAXJbTxxk+2Chw3DAKnY7U/z3Mw39sKE4vwecRfgLV
+fSrqo4dONVucisPgerSHpIcTCiuTLjF0ASmlrMhRZLs5NWcZO9sCIK8BfRnD81M
DsKVOVZR7TP71LBqZ2dQIaUWEvQ/uZnLaqGAmuTPa4Au6xmcLgbHkw97Jshej866
CqI1QKBSi6lhqkkQnqbpiov7PoU9Fv9EB4z3CXieM1Hj/vquemHqGUwZNibB0eUk
LhLGisVBT6P9ROBmDzzz9yacrnJI7dhdb428SKsYMrCx1cPBuoY174IEdlMXUFVQ
A32mmtgm9SPnKcIvUfkYgWu+ZVbmd3X3eLwb1zYaEflh7UaN7JqOaNws+XqvYs+e
SVtqQv2OBDqDhbVx261CnzQyRNABTReAt2eETUXiDm9l7zCjcBj5EuhdCZX+GnJN
Jb+OGvcMtDxAcya1ekCW3owRVpM3TTn8UsZwB02DR86IOhaBBtF+EeK2VQaGaOjH
pUuZLajar2yXyA8+AbOBrZl4yxjVkuKdMRZr9P9PCMqflSZ9YpewZdgbE4wAVEcF
FnfutVMoqIzl9EYT+gAVrJ7ij1EcsaBKpHVtWvrhZtK/XaKbrnyeNZmmKeRgxVMW
aOMjXUHQdWqGbMTQ4TVQaH6WYc/sxUsP8v5C/6j1o8veR1nZxHF2syJr55V/l0qd
FHQiGEu8tHiZMAxv+4+L5Pdbx0S//4pvx48pdz9YC3/7XqIXLjkELPB9Jm+CNPL7
q7kgJt2RHLbBBiNXrl9aIaY4H/fLoZjP1AvqSI52ykipE1ABuvTVDEKXl8lc/ALe
o3uhIQOmFScSPYHLdhiMaXODxZKaf6DKbYRSXK+6WeVK+NZAu5UUJKHGDVyLWbiI
9pfnovjuztNJr8QdCpj+0pxG8h7yP/Chs9y60l29Vu45/YDxhcR499hfOGBxqUbI
wPMCVp1eUaI3msL43ECU5GAjz8GGrRXSHWM0QCHZbaiNCxKE1+7qzgAnmPvGTddI
4xRt9EkdNafx+zWPdXsJ+I/jeoVmxL+/BIoWLAfiF2bugKFZ+Y0+Y+PF1I35O/Oq
q9eE+i11q7ufCg0QmKV1s8Ly3jy17kSmGl7kntE2CsLeaB4pr8hPrAYkV4a2qPb+
YdF0AMQGGeZcxjhOl6twsk5sEALgxYAY0EJqS0lJr0qThTdf7abo6aRUBDOKgeW6
1EkRRDUCJqoEJ6rg7GDd/jBoHpH5oMfhIWXiKaimKr2oM2GGQTl27bD7UoG7APW4
Ss1Ue0KdstO1B4w2Fo/nB5v+pBC5YWXbhSi8UiKs9EB0h1h2vXl/ZD+pAyBoFrQ/
9C4oirUArj1jd2H9MCWi7lWfwH6YRsYKITXH2AsmFE9a/B1ZJOf0PSM/lAOVpTcT
vSWrIEV1yVaIpmkI2yy/84Hk6z/z7ggw+SuJhumcYekH+yh1Gpy4YwfdhXnHFKrY
VP8TaSr9Lc7Vu9SIKlp0Iw+O4FDtEpG1sJkDcHLsO5rTRtekb+bcvCYwcIXk3hnc
jAQEvWLMyPoD6m2fsVIiyF64c0s4qWTBT3BcotauyhhMQ+zjZusbgAZBOxcQUVVo
0UD3yEeSs8S/l16KHJ0rCqaKEgB55P9Y4NGpLwgYTFdrGVxFYyuF7kPSR3bLqwRw
tqYZLSBItJJLw8be0TdAE7xBKxXpMo9c7tXT/bTwCHyjUYAtxnx209/0A5Z2YJ/O
PrZIOMGRM6ZzMypGDfTC9lmejz2jln5tEolb0ggNG9amoNF0Cu6F74DX0xPGjT0t
0cfkgWDrBDHvcnWQYgXNe++70CvMNYroOHmG4bg/wh17ahSw8UBfBSaUXJ/FAM6S
th95ptypJ1S35L+uJcQZAUx8oH/GusYfDZoI8bFmRuAsN1sOXBypQ2MAYNpWvaOu
wTbHa+0X3Ouoe6i2pk2COxFWhwxWvFLs87X4cIFEM2msicSn6o/2wOSW2P0Gpz4V
gL3aDfatuMxhuju1s7mPVYpXbr3KDL7TFBAF3gzYPonj9qcT++kU494+yz+w28IA
NX2LI7HeYlQkf/8rZnoXf6i7CrmeA6LalpKlXZEAYrK4wE7ih+oiaGlC3ceVmv8B
2+DzEvH8c+eWbV5J7kkG4eVlsVGYaeRJEG4Rttsjp2WYl/JJci95//9Uz8fIWQQY
f4yUMPbrl2CLv3iMaUmERU+kv/uTQpyG5UE8t2zyfzXJmV5rXbwt9ESHuQyP/6vy
MZ/QyAx6m1WuBWtpsNJFOkbYWVy+/4DdBjnKTEZOrWB7IKwY4ls0DWzH3XE03b57
V5fVVvPWkUuuUC9XuvfFOaB022Y8UU+K5HQhBO7DJI0ZF3r2NIibKy9UVGRgZFcM
kG3lyxA8rKXiO8zX7tFhHUEHgI1MXwvgQY21LPpsBbSYi84YM8TMbr5xJRCXqGPC
7hNzZcEgGbgqW3vW78ylGN3a0+1drep0BBpppXQFEJCdenRXzli+11MLRE+9P1pu
eUtPDZto+WRyCtSpY750LU/Er5C1311eGUjlZBTffyiujv+ScXTMw2MKXu4bc8VP
RhOWAVUF7T+pBEbY56HdhVdSK6EHE7nwaBFQYwiYxS4scKd1VEi6aBla7+ch1YOO
jXteGdlgIVlcbOqPu70st/q/2EZ0rZHRkDPcuM/U9rtMWm+BjfD+RdKMST4Al9cm
hRcRh29Pc5FDweGfm6F89y2xUB5CQzk3yLf4wmDznYHYFnFV4LI0wxgeey6Rxq94
ocNY7gwh5sY0CbHZ0OziBUr10v8GWzG8PIL4kgf6s0z+3j63RkxfV4u+VSxcEmyC
n4dt1kef2vGL+ZnmIMm6SDoDaHS9A20aegrQ3bLufj2DlW0BbILt7PHOJ4+i2aWt
NJacm+kQyJTomE95gfUChPee8EvUxw1/KnZNg52HPrYA+EVroqdfB1NgxTFV2mIq
YLg+Zl7tE/vY7bN0vnpTRMTba27XdWXrAxb1S0q18IVqQBQV5f/dcHMLqjP53Xlh
MTTP9srw+4XSVEldZ1/z9LRk+c9vQZ9wWkX25SjLRPp7nX17ENOlgx52SphZ2d9h
Dls+Sb4x0pafK7vvjF5z6UcHEcEzS9GotCot2K9mfAHHJPkwQ0wBgWMoel4bkze7
GPecydnP4bWzEbScoOWaX/1ik26gMoJVKcXDDcwZ0RVC0Vv12k4Z188fYqeEaJaE
fMBofjF/hxh0jPzInPnSxPKbJ57t4iVzVamJ7mrOGrv7eUywK4fU17YT0OZdwjog
3g3bgBfmoInf53Sx7Gxi/eRJzaKatkv2hmA+SfeSdJU1AYs6snY5qEHS9ACKlxBC
wkSxXn/d5NLaUmKPNAHjz+kxCDp9QbjsWyj6gqIqY+pJeY4L0C/LL/d8XbAGUzG3
RNx4Shfl7Plf+Z2wz+xnFRcc6xMQgCADky0FU/ro/nQD1TSzonF6EBsPsBllJclq
MIEq+J0o6hCHrPEy6+BI6uit+a33vTfPqU2wmZIK0ufHaatDDTiKkjjj1myazQv3
SnT8iY5J2DfDa9hmSU3PocZguDb1LMIzjcAC4vE/YgoI3aIPjLsBNrWBYdjZH/+9
IHoP+mAm94+Lov+BEFtb1z8njaNBdI2dcCuFAtr3yh4iqzJ1Q/hKIsKSTe/ytVDX
byH8YuP1r/A0v1Bwac/uAM9rxK+1GZZEhPK9I1NcodYQs91jGfGwtDabLg5XyeE0
uKdEv03omso/XRDTGdoqWF55n/dfdjj+g9+dmD6BrJMP+ede+tArBFshFda2P5XD
dvojtq/VVbwgm1aGCaBC794YQjWPYnuyFQVpJiBvVv3W6c2thPZr5YIlGJEkbL07
5bJRrmZQ3Y3RPVhKlMLFOsORZtAeF1ybREkJeBDWYHTCK5ITdaXCeBdgFhIZbBVr
erK/XsfTn9W2IgwNSU3EOPFiDDT8N4J96XeRLJ4lvZbRarMwWo5ZBapRg/4OrZmb
1KmfyiZrMZdwOSWlek/K/SHuwYEH2iEuX5UDq+M5wO3BuzDn8bCgUK3l52aVQdBR
Aoy4nKaLoCT0vYZJTYW0yPiwiaWVS1bvSGCkdeqfXzhcAuajx+fVckP8jnVsePeb
QET3qr14kRbkKZy5da+tgUQaCLKaHibXhzAJ+O5SXTPTV1y33rjfj0LFaV7sBP53
lzQrrGtI8mK1mXoYkAv3KiclorULPRSVQU7vVHKIl8Z5iw6ERs/9Jv3oW8Q5IbCF
j6g0CqRQ1xIz48pMomVRCq8Fp1lzRf1UktBb94sA62hl5zBocE7FgvPqy+tKLf61
IDnyKM0kQw/MfDwpYGPzpFsxdot4XLNGoyrYDeHdglb6Z65b9YmceqtN9E2K5DtD
LSiSQWeyLXAGtQGQeBDxJ3EyRQ3lcUAVnb9FTU2CIGNnaLrUi5r/vMVC9V9zVlEi
NTlBTcfRP6bDIHq4t2SGkVkEO4DwkXnr4HIcpqPhZTgC85NWHqNLTfjBZJCQW1I0
FtmxcdC7UQEmbRAaNQwhHP29vKeNHpHwSnICa6mnu+r7f8d9yQZhUgfcOA3AK7oQ
THQIYHsVAAMHppJdlSyIeH+Q0NJUXJUq8ziyW5I7vM0NMXKIkC7894D6KdkGfNfP
xSgQ6z2wJZzAY2rfKReGMx2wE4HUEwX7WahCl9ItLWIr9Fm5Bkm3+oZrPy4avGNl
kpfFB+HnX42Zkg9lkcWjlpbsQHQsDrYiReVDZ4lHvXnm4JdqZN548MzD1kNUB0Ih
fzH5qrNpXbPprov7qCnp2Z+3S07rMSz2KwHEQ5relrzPMmXmOrRZ6DL4rwgBz9U1
clR14pldXjRZ0ygoRYlpgrx7y0lw45qMd70Jr//aplA2vaUa+mJX1HSgj2vC9TI+
v6FL3wuzRK5LqLks9a6qRwG9xcoz3r/qMY26RfATCa1JEwwjNVKXGbtEJULsCdj0
c0ird2RP75XTB7X9bIsfECnbjUM7Fxwk3lNNI1GXsi2/as328srP1xbNcPY6c2dw
gq+P34GdB1CUKZ3genXqMNG0a4ZdbI8QOFbLjr9Vr1VYNXxfJCJd0JwkwTXKTrs3
UNhfBj3JFcSieOsTVdgtiWWykLdxvKt0wNnSXKHV2qBU/DH48G9rx+9dkucq/HrD
85ofoG/dA0dE/iPTjBdIy9BQK2+UUKHXF9ee8020lxqaPjo9sTNPWSW6kXbiaVuS
/A/HIM5Z+YaE03ZleCePsX4NSkeotmqC0orkdj1A7jOA5RrnOUrSueVniGpEg+T+
p9cR1Z7ocTzvyEhC3WrjgAoZZJ1h4FyO31bstBvZ3Bxi5aD9po9UO9vKgxOiGupq
02cY3YD+PzXwf1WDsk+YCkRofhCmCHTAD8lf2DHdSAHxC4dz1UMPh6ZuDDNVF7f1
lRaH/4vP37b01mhC29e4rsTlKJJTehtwsk2ey67XLt5G0wGKDFCADQf7A+eas42T
OnXxovBvJlMQ/Rg1KK3aXpN0MXuF3MERm/JeDNepNaYhRMspxHyK7Hj0zKOPVYAk
W6JLArbZRT4NIw5K9HZs+seYI3J1qLP9wbrkzls1vFSltk+PwFu62Sx6R0aBmCRO
vDCvHXk+7c+RjgwB7yZwuGdC66RyUl+LzkVAHBOHKzUrUJAbMHgoSLnUosOqBCE0
Murv+ADrN3X6IVIXGTw7/BzpXwyf5DBZsW5hR9PldLNwXb6tndEtYLWFUeEJI0WL
IaJDNvayuBU9nSsw/5aDaDGsiR+SkZZyEeTM27XqJeW1nMG6eXOe5P6D/3quSFhu
yUSKyKTcQ5UuFzBVU6zbLZKg7a/VWI9v7tIreLO3hkSwOk/0QLIkBavVzaqg16pJ
8BSIf6YLSjBh7QX14rguJRdBxdlE0in9D9/zS3w4NJuNHYqm+Iav2gE2axwdqnwG
DGVfOBPNN76ixul3geSxMdTFR+PpuiP4cIXmF8U5wZHlN7sZtFf5cEnpblIh1qJC
HVakontOGTMrHiKjt3uUCvwXhzXjhb49cdpG9lEhTmKzX1YZgyQH/gvUCbVVQoB6
5GBYaVYH5m+Fed2EKo4jGcrB62iMzyQ0dh9wszyen7694BW8IsJqCQ8TQd8aVwu/
cpxXXZNIDPZrTEm+btHqmF7XMgteBbkFXbpTvojwGRBJt5uB5EuZpubcQjBNxgt6
tsW77DtUhAyBjHq/4HYGi2Nb9peLoXkiiWAPC5QyF+ItMXmVEBLKArX8xbAbeqhA
9NsCB3rDqnOBZ0qSXEVaWl1KAVou3XaAxXNpGlO0gZ3k8SPqvFCJPqA6zjnzLxLQ
HXcwPM/RvjiwnTLsOtKy9lvH6CGGe9NSEif3BYak6JtBLXiSriGjvYW750D46ClX
bzS+VDlAT26W/2cxchdDEWfVjOUx8oHAN0pbYnFr5El8ceVh5oz2l3PCOQlvMQGU
ZkuafcKM4Yn3yvCyurLUoOpOUjr3ruFyLg9+htoZfdSbq1eNikMcDamVbJq0wZmJ
J8ko2SS+a7H5VmiIrXPv3BwflMuMBKTuDmIAIfhEzfTEegN6yWzTg97nCGMuwMWL
RCmubY5Z5IzfPleYJ4l5BJ6pKhJIl3cC3lRkuYRfKE2/Y+r3ArfCN1ig7ZdE5WtB
v1xxAQ0ymVVPL0DkJ4fUVEZkvElNSHVQPwGaJL7mrs0HRZ6nNPE1NWxM6wg0Qv1e
M43LaWj6RzFQAY4U7D2Vaq1W4VecTHqbggCNNMcDKDcTzAEEH/irOjEWKtxYz/wr
zDvF13Qdt80PLHhUpShDZH720xSvswhKAnM0OwgbmeeZmYvdRAYbokZNrRYSigLQ
n78hGI+qlFymBH3OliMWPhWCQowOgkkAyD1uz7998o3ZvKzel+6FCeqtAh/kdbM2
ljp04lueqqs9z4wdG/0R9UbS7br//+Yj7qSXG85cSukgPD1pyv3uW3bzuu7ggSo/
QPv9GYj7CJlDKhjj25EaXBgY6XtQ3yp/gMLgMypjH7d8tEaCwFaHWe45AM1vLuKR
WEK46bp7PCFf+h8p8Yaj/03T30MAxIN7kjA0lOnYMCV9AJDQllKNzydsyG1Wopfl
6qms1KyZZkAl9JmI2tOW5xdDohMossVlUa1Iugzjf5O+fzVhf6WePvV2dl5rn9Rm
kTGTHs6pVBQpO2PVQ2TPkB/+3NfpVA6hAAwgem1dZTpPPGPfVo1M6cfaqfijzzWd
UtGfA4ADMk1+HFaU+iFADONNaxJ4ol+2ff/PVs8YtzNzVBLcPKrFtF/pb7C5Z77i
LkVOKH+pWWzC0keGnaI4b4OsRLcc5grMh49L30WmbiuPRwRgu3ztpojQzkzx8bVK
qyaGAZ10WusOR4etOjvX/pUZ5PbEH2UyPEZeyL7GdatnavoF4k+o2EZ72BqzrUlW
N4KFVEqIgdOTJM5szeVxR7bf9Pn6s63PGc35OTR+DIqEka4WzqsKbgHtT2f9Ovde
D9nCLbtdQWyZyhE76PwEVkofZ+NAQ3ifPXsovUUtfAzCsxkGkbN3X1agL1KzG3ew
T7uiimhgcqoe06lPzYOwVAUiEbSfKf6EiU3boRv6ARC2MY211OsyyERV8dgQEWlg
ype26WyDwfKQV1TfYHdeOCU86y4Ia48Cqr95wFcVZ7/0nFc7IJVD1yqUJKGZxgzM
l8AcKc8NlQefl92oBz2HFIV0KGnkG+jlk9uMIEis75oGuekI9PweofbHvJEcymxG
CO3j6O/Jg84FvmogwtSrV4yVsNK4wnEmbJ6BtmiBYkdgVdkUM1S13xOIueB0Gct1
KFPiD9LxfMqxjSoGN2hVcY3EfyhKzXmpTKtlL81I1xsWnDQMKOVx5XhewjAQNTR0
JyXxtYDc1Otzz2lPmWRlGmJsQ3hcLTVWRxFHTmxAE1GY85Qmv4Lk6JJDJXJgOxSw
+J4xdhEe7W38bV1UCmBXlBWhFdfC9irjBp3AuZyyrTIGBBbUaGnAWGEQgo4xyi2u
eE8Yup6PKijD++bTAT0DD9N9PAUHzWL/82TUR4wsBug3wlloR+7NKw1vKBX7igm2
pf+0HB4OGtQtr0NMFli9B19gLKR7y3Rl+kCoWcepWUP0aMnaklMGNux14lE2GC1b
wL7uontaNsWx4XQfRfnsMtZkw0eYeorSMKpQbY/BE2pIMTzSzF/5lpafanjoT362
XQ14KS/8B/IQN6mOo1UCIN8LFoMDHS7qWiZTrt+3E7/MvlSb9+WMYCvD2tbC4Ah2
t55XUj1qGXrePphdgrGUO0LReenCKgyJ9Ya7yjv40SCF856Df+T4fWC5r+pyZTSd
OwecNWLOudNo2Yv5m7tmgWCEOAhbdfqfWXp5wVQff77VIfgjFXGGpZRTU8rpuLin
WjZCszjhTrCWVJ0RXOSHRYdsgrN2ivbFsEs8R2uUWnplEikCXrNDmA8EbNB5m61M
r+I9kmKU2a4FJGvi1T2UDPF4/1R7uWXKDH5ZdItN2rTbXnpZMhipMWieljSirMXg
8uxTWzVw2AGCn5gxgDcTlc0Wuj4QxrwmJureRYEawpqhQalWoCljYIqYsJ4l0Xpp
sFm+7UFdUZyhSiAewr8O/BzA6lqvtX3L2ZgF5IoyEXvs/icjMSzTjXbhgsHSLWq3
HzyGwTqyiZZ0kYAXccCP0ouIPkuMvM6IR5OkNND+HYfzFjaf5vL4+tTdXKSlEeCr
YdTimd7jXaiLNfJX78fMdS722Zhk4dPK4LM2o6APuO5YmQRHMKpbsi5D9/51s6sx
kzh0g1FYsVlAKD4qcy4a9aJogOPvvVhQU4M6q+8aiDGrrlUMj1Eheddf3HdOpYY7
se1Fj8KqjhhCgl1xNya7ism6NTCmzNmXTm7LKWrteO0Im7NnVaig51ZuaSiqnX/D
vvX1V9hWEr+NiMRS8MlVMWhGuS0aaVtNg07wPj7UR1MRgevqHcLjrEYq0cMORLzc
J2a35S4RSWDlBbgCaitEtmJJOoxkYlq5vLYsZFWRnasZwaDWmJJF5Js99YJJSNhH
/ZdyA2/zA/PaBGYtOXpTuDMLYHznL245VrBxtWC5qUGTOTWlmW9uFgtvQMaAZ3HH
+3GJKk+cyAhRANO40NoFwYWhg2fzBrUVq+NtsoW8xVhDoP2ecWOJkeq1ZCcoAATT
L5RRb4lmT7NCZw3J6cLJkJtIi8pptoZxWAPssNVyOpi0aARJy6J2pfNbNVlzFEd1
zAvBtFHb8sq85cKm8Fcq4K3wY2PxRW7mCsmRu8RvxODlCU6jJGhHclq0c9DPXPX/
g9Qbhblo30h2IDgVSo1j7FxhH2uyCQlMdPxANaXGaSRLtWSrUpSb6ZN3TZAetqvY
FibGOhQPA53QzhxePBvwob9dqQuDhDamHiomgzIX9Id3sQr7bY74M7ds2mhAtkzh
opHzKuyS7k11EuLw5nw8uHCUkfE4lxT5tnDV54zuACd+h01g9c8wjO56u5lGm7JW
dcrh4zzjWercelV1zn2Aq64Prx1xLXC+e3e1k/6Ut8qfmRo9vpOtxBWnrKrUIemw
4wf9TOAws2SC+ofazdSnAt/6+uInI+cjYAgWOnFqgDEQXTUJBfiWTM5L1C+Dkhhg
kCKu3TJepRhRGRCsG5JnQ1dCXh5z2GyFMdExTO6uWhnzNzbEy2yVV7mQPAnWjpcb
xddaRz2VLozJcQjsNd+2VzoxesVXKExgYlPngvHjda75vOYVbzLnBqolT+UKdEXf
TpA7yIphBwI97xDsGZkdxWNdJ48AdPylUcBAlxSevDBdB6UCXbetv4p4dCC26R+l
ge+QMGcjUcklk/5qFNfIfpFtkNCcm4a0NaEa3z0sMDJPibdUxv/D8GnBys8JlUQt
3YJrkh4O2tbTTSWqAwfZAJDf/WJcXBHlmqJTfMF5tIZi/dVf0Kv+fn6hjku/B4fZ
F5eHn68YxdHD/saM85IPz8l70oKEfxCdVUbyDcCdW6TWRdG9V/+bFBkY1TDxGF4N
nOMxo/SHCR0UL1eU9IJSat68yQ0+a9ohh/8Lb/cvWzlWhIjt/s94A200dLkvWQNe
gvaWkxrcT0HTkcN9miSPqRalB96VfHi3xZTCJJbv0QfeBi8TZoEGlVcVlDJqbWMD
M0ZSru3r25Lh5kLrI2ws3bqeh5rCMX7tsjArZhaNBKmT0SPWhjcJcL0TjAAvTWM5
i/23G1WjBHjWMmo5eT2qLjtZ8kQWgHrI8eNYSjaPu/OAFleR10asjNM89FyIB9sI
E0s4/cq74dgvrlzBX1rfEFIODa5QEfEw5umZeyvvUuTpTQvxbTyXAJY/OjL8QQWu
aXFRCVNf0TFti+a5E9zRFUo65KsJvVvDzyIKK0WR4IST/oRqXhdTztt+22AClZ2d
X6VsFf7ncjy6D6wMZdI5Gxr3HIV2W/q4n87QDHhEEcawWVtOASsEbO3FgKABvz2s
VPwgEVzqgqfwrhusmjgNgkeH1lf3nssyERtaD+A/EhaxBk5Fezhf36oig3FlKtQv
dYShIzSxh7+BMEHfyDoErQtOqjbExIVmk+S4dWnFz9wgP5kSKQ9Lbv0BYcUDi15c
uo5p7y5f+b8WTrN7m7l1zNdp7NKbWdRQQb67FgCTmx1aOhp6C19UabZ5sjOgn22I
FedmLBj+bR3HKRu5qYnNdDh1zNCpp+qGBdx847stZJ51z785ZteTZDXU27pJpuQG
wd6vLGnZq+GLc82eIsrQuNCDg3cQl99DVWj3LCqisrBN1sxmX6/HR2mUH2xDrtOr
sqh8zOj0R8LC3JEIQNM1KKnQW2cvfh6EtJHZPar46bHpdiOMwnLt6cD8vI+CoQLt
AsPs+tE63OAuaiJth33Pzni0Zz9eUxikAaJx5yKPYlzUok4LkBsvtf9PnbhT+2Me
B2YO3RkryJ345t2SCDP3mS8dEWBzxhQNkWWdBt40sL4NChNh8ymoUpI0pbErZEYr
WxDajDKiOlvAUDQmodNDpGbcVxu1MMjKQ0YfLHybIJ/I4wHW3vCuHndsg201jdrf
RJ5EOnn396dUGHVz5ZAc2nRHqJ+JqGagpm7xbmsu6aY0UCOKxoxUnT7S8Fqr/ABt
x+aPOp6MGBPBf0CGWUnf1191hBwxmJb8I7kjjZEHgThczmyfYLtKjwXkXk+sgGrD
fPH0TPGLlJofBsUa7sfU7sfhRnTMWqv9Lf8SagMYZ5oFmfwBYDZPe9zyiDWOTT0t
55RJZDFYrTXFBCxd8tuc6ol/1QEwVmqXEpt13MaxNu2DzE6AAy9u53pypDsRhgjR
4f/zxOWrHNVKhMxLSWHQHtLfl4/RUIt7WDkLptqGPX5IUMJjxzhBCgf/zmZpJKAQ
6Eu95UfzSpTMhdkm3eTSKoNEktEzsVPpXbjJVEaIk5O7DlbQRFSqSmGXA0rP7RDQ
djklLfSMwKciFxCXuUfLReqemEOfelpfKcaWhD3AACyJj0sOBIW7w6h+mqwc0jnO
ZjNisz5czSx89Qz/xfF8gdF5RG83B5kR7YGlxEdJMCFCdbJMmGvqb50FbElIT5rF
e+jg09+vQyazT6sV9nUbk2S9x3qNYrx7svOazmjkuJO6TAUiYao449oCV6mltw1u
TNY2YpLQ+PQkxQMC65HfES9psedkpCsVm8kQPL5YlzXJq0UMG34Mhw07PPCAIQO4
VCfao51WQ4b7Og+kcbjty0OR6DxOUlI/M32tuTCrb/Kv6jS6gRtmI8vkrIwpiCW2
j2XXzXPBTXNPRQHnjBlbow5KQnFzKX/bH2JVYJSjW+jvZyNR/0Ii5ikGOb6OxorL
N4pTZCbVuyWvzZhxUnQZhpd5f5Mhp3lYo+I2de7hjTtg0nAWALieoDDu05LxCRE6
yBMleAExJG575ivqtEZFby4dIKV5oHT67OjyXnt2hdRzXGcAcMPt6bHKqRIrIxx6
Epk8nA/X/RRse+kVhtKL7pzSDYKvWGuaW5FnbujRHhXisY1ilv4q4fpxBTqG/cb9
KC5Rkf0el36lPQO6gdSu+rT3cPFo4noG3J3QtSoh+tMxw56Xyuz8Oe5gpVA5HMJd
sbvaOAM81El24kjlA9dPDr7cli8Q7gVw/1g1EDQGW+rKGuuEoMP4UotXAAhGCRQe
REi5S30ltVZSFJuZnAAPeYF7bmchvi6rxoGzV14kwZJoYTxWRrzvZB6za2PDgFQn
Kbn0zQZ+WlkBB72Lo7kRfA90MjYsIqzl6NfeOESvum4wjlAU4XbdUEtyCS+DaGIX
SL9u/vFfnIEta5BcOFscBLt9ZLSO06KPY2jWQ5v0S1YGOKe+NFMDR3XaElhFZC1D
Ba2pZWvyGZzjJ4LgGYS74aQxo2jUuZrypvSx5D9zTCYfVg+xcBnfp8uMujkIfTGF
SVRmDrYoXzzwU6tvP6Kkvl+LkP2gDeSXaOgEEZ4ARpdrVBaVcAwFA9NI1PpJ2rsa
LC4AiemlqGDWTTfxxHnb7HyF3uK6VoemcEK3hm1OXo8m1fT7dVPIsY3XXKBgMuIr
aStPMf/X8NhTA7Xr2Ubo49sIwVpZUMTR5T0Q0w4Ynixd/OiSdDo/ITUrWeBYmwLh
d9qdW4FE9mBWxg/w/77ymzdaJ8lc8Yp7jWZZZcwmVg15yID59Pt4+Nn6sImjrI5E
uhc94W47GcC9jWOre95eyxDr+XfQL4hJANkLBl0eYF3Jx1NZ83FVMc4WVdmajr9H
Rg98mih6TrTYrWLur2xQlyjNuQmNNFxrHQpuoKnbMYfDhrenBkFA6AAgxtxqnYoL
WmeUHSRIK+UFlPLvMuWEm1Elhq9nkBBUE0vjO4z0YBrdRggKOTLm5cZVOp9YaG9i
E+vuJ4RHqXoexovloXBsOKK1ravKHy58fDwi/dQoi2mInYBm8ORXQlvwg0GFgnP1
6GKD/yUGQQt8vMJrS8bQ6kKNszBjisUd0rHiuvDF7+to5SrQa/27MgzYLQn70c1b
6BFY57JTYpWkidXMlyHcWz+H1/WzYTymOD4NEO8nXlSuv3+CAdPOw0OAxuXdqVKc
GRK2rf2zfRXNmRhxLYRg6xJldBcG2twImOluObRgQlsUmTnRLty16PnYOwjwn9by
BY+Li/VSK3mkE90grInY0a1zmP/AL3QXBqkthBWkxNQFu6i2lGW5omXySdbmVQQY
tGk2XX0ca+K1UdW05M7wGXv2grdy7KxGmB6UgBVHtu0Hgh0bVA7xKzQfTnzsXJpr
okzQuSnXJwuGvr1NLg5AmBauFvflBMkOFi0C7ZWxc0DfP4yKcUnGdVt+VJ1Pmee4
NyLHlW1trOo2HWoNsRaHLZ3VA+Zayx1LwNPM8D6WLi41+otuwtn/nuI6uZ+9OjS8
3TbsL58WKHE1vjt1EQgvrQw0Rt2NbgS2h2++i8spVVisb4ikgZ30I5vkAuNnUzgb
v87iH2BxgZUufqjBh63a/LNJ1Bw+OeJvKpzpk9a8QLDacrd1h+HJz7PgoWveZDy8
xSfwiNEET9N41aipHWIShP/Vv7sRy71bXuAcwZYQ4YoCUFrKFCT8vrRMcf+O/ENE
xzHXsQ6ECK/+kJtRM0HU0gsin0E2nxYN5E2wh3sHFndE9e+QTyRSNn01/w5QHSXn
ovhkNYcQHxwTDjiptaGyYHHemMFnKT2wd4ibgCZ3FE3V61955RlwL22WTqnlAWaM
0FF7W0+U2smEKxW1SCshkJt0/fv5RWSqDjCnvpH2TteOItzIQeoFkfiscjBSByd7
VQ9/3Sm7mRUMsEcNrVVS6Ki77PBDLkyIfhf44qioP18332M95w6gYv9mLlphbTEd
yhU2VOtwwcdAqFaVKmetYsKAaw6bVYp4nbmZG+75950QhU479T8ZkCFVbTCbN6Tu
BQidc1t1zfkgf+tBeqA24ng5GW/Te5MOQTXYoDnS9wWFqZ8MhIxxpxC7K08tzJqB
aApspGJt867JUpCW81YV0rvHjxVzBDO+z1VKF+Twaif9NTy/104qRkJKmCR5iqsQ
mNzPyKRvIADnbVZK0XlxvX6zyxKb5sY9+vGcubDcvQyxae84PBGedIhbdfIQf4Re
ctp/PDIa/WaMaseD5Vcq+51Gd3X1a0AVd5vbIgq/4RBdaSZvPma+ijb+OGupD9vM
GIm2q3REBOcto5OyKhYcsw4auW1e0S6/Vmngi+jbXuNo3A5K967bEvm6tcCxldIq
Ht/5R08DrpnqOv8Uo+x1Ii09mXAq65UYsfPM/0PaBbxCUtz/1iCH7FCdl0C5hqwQ
EyHpu0HkuXBA9WOIgncsEV9Rpa/bzyZD6AnjO6HSp5eV5LDM0ZiP5+TNxr9PbvhL
6Pa5rSaI0DPAm412gWFJw0GE3Mz4qVNSHvDiE+WjmyJ0PZRvu/km+yEaHmRrV02f
dK9wGYFM1CMm1az+X3J+9Nb+/RLfa73LTeMPHZNxXQWHO9ovtGBUp08901O0MVs1
z+Tj/p3M2EwF3DfYE+8kRRAEH87XLPQi8uZm8ElUwjAXoRbirrxT2211jHXO0Pwg
irCGShXBDXU2ZE0o+OxRRCl4uH+kZZ695TQFmRJy6mYGtGv7HkKp1lkmAfsXjy1g
8e+nOg6zYgg//3NTSNrLcBkT/SPbJDt5AHSMTS9Y5GB9tyKN4g/c9bE4sSvKVCRX
o00r5N75tPXCFOcNUc3laplVxOl7ESPQCzYTmR6WYy+hp/lDbwDJazs+z3p9bXyb
5IOldIm0a01BdDjlFgS/Z6Bred18I7ssExMZJuTh6nwOnPMv4ot0TDo5YraLo2MU
wIOwWSPI6ZAIfnVbFDTZhRCX8ah35J32+mmwZZn1U/MAdoimaP3jPMGJKJZgwXdL
N6EYjhaVnrR2lEb90QQWFdIudkxeOYFnVesWbQF6wvtFkyDWMuvjvEd9/L/Fgxfj
di3NLHJ1BRPi/wmy/uSezSdUpqTzR46SPOTLPnqrwuTjXfMtwSAA+tLYfI/xtKQb
koAlz68n9p7KJBk9JZASESuw+CZLQt17V9pLGGqnFlrXmRlQ7mgNkOKzc2nOdpbP
uk3891pDZI4T3Oi0wrILYheXuc0+f6jeahcYE83S8hAdOZIWaF6wwU4WeIb4DDvX
T2qfKQPXji7ty5qqFzbynIP4oZruzYDMEXRqjDNVB5h/gJM/gy9hgcZIRpPVVjKq
mhJBYbXLAwXqjJOZlGC3u50toQW83vQGnbTVDZkyxRsSXCRf5rG8LGQ8n6c5yts1
LVQGetkR1gcYpJautITur6N1CQnQKvl/pdajgHoP0MoEkaGYFnckTrWqH8RxhOnV
09eLobRs4YEmCyb6DIb6JEm5KrWHNlSAO+A2+MsYvpSKqFUoMYhfcl9e9VWowwu/
UFTj7kYuOEoGSdc8pdEQcpQ3QpUv8nqYRFMEM4xCxPIn1gVaSXtL795j8U8xVTn4
YFn3SZD7VHzoRq0Mn11cuDMWCGiIKFm6siHq/UBerHy0HVBiIvd62gOlFg3ksGuZ
X1w7H+cXYmBa3O1ufFvywEYeQdm58A7kyRYDvbzqboZk9oy8GHR994I7RQBzxbb/
zPyLAMsbR3p/A0Ufmj01oiZKxKsfFSzRLRCp2msrgkDf1tjnorvtzSSkG27JU0ZX
L0aYylhN6hRRFYQ+G3PT22sB9FP0Qj3R/EOmUeYpjvFyX37Yld4zXyaAm5PFuLcS
LXEJ8Oej0FkwnP9zIKpKMXu9Q16TYNU9jhWPtCY+47r+jtORESBicjAJZjBZVhSb
A2fuyvQ/UVlWuLxkZdGLWRhjq7x6snt9Q/1Yrs+rD6fhxbhAtxIsNeBGtCZ6tTCM
YC4aZ5hbWz6f1PGSikQvXOIJjx2xl9z2nEVC6/obxvoqSTQ2Bt+Jd907vT4Qo4Lt
yKSYbIGUfQT4R6/EqDswZKE7bOqU/A0dT7Kmst2mvnklAh7CAk4ivs+KiOtf8cxi
BctQgfMUioOaCGyH+Ia8c7/b+UFxJlwymxsCI93I9Xxx6qED+ZSLJbD3jLNw1bcN
Fl4DRZqmb+tz/VJ9eBfuKD3moJ4rR8ehj6rSr4MLXltG1xEp2M2/zG5tt2Eba8HE
p3fk53u9NmjXdMmtmqoBJLOEbP4DQzwhJV7ns8seJ5WuDtU6OOLd8tM90bPngJLJ
kiiD+TtYkH1p3MaH6P1Wr9lYRUmal1eASbKvIwE8CITrLe9WthL1eZ8bYf87EhKC
ODWUR85xWprHDaUjKDO7XoCHSv9KTT8myiPwDiw3h+oYb9ycgxB1utf3MjArH0rT
V0xE2QfNNrECHSi5Tymji4TysPs/Qb6eo4yZEj11OSg2cAM/6uGAKIGSvr9VT8XG
XE0qLJX5vk+IEP8TI+/mOp0YFAyDQzBZMRuZ1gIpsZ4c/bv4VI3D9tCypidA9AzQ
P7sHJ4s3+vzZEqRbCSXNYZ59KhUo7KrXESCY9cbCc2rQsbFGJt6Ik0zBYAgYOCWc
6HdQAK7r+LC+Ht6Qy8+cVNsp84a3hX6rqZH4xLf8J06EaMe1EF//quleQ0R9r+zh
Ayel126Q4j0f7h/c6xTEFUYoITnxf1c62BMSj/qW++KjS6ZR2K+iviRGPB+AwpmG
i22Rrdl0f272KIWt9EzarvrmglkVOPrM0a/NfNxrdzowItJ33MSK0ggOVu5vkLe+
du+5Wxq2nHxmuFHwTcq5GiLmr3uqAzhfvcqz3KfxLwNKS6WxRgN+gJQ+joxxrOMX
OverdDzAgVGGvNJ825azpjZuJQzfbBhiMOcGEo5NX4lAR9qHYa5d0EbHe9y+ct88
TerZEWzp8ngwMwA7LMZH+LNFgC3A4P99eDLhg6zN+IBYK9ghfwioqMjlAIvIyzSQ
Dii8X/EipGoZzTasTxPwl91k2/XpuGqzFIuJzY9LydLlnDDizxYH7EvxxvXWTef1
KmpPxSL4W1kPfTTdAVY4Sky9LQKdPf+SFnNEYqBa5kdQnyrV0LGCQSdm8s5G8J3L
nCc+0Vfa3RUB66PwO177p+CIsXUp4Ib/qPsuXIR+ZyRDihSUJPMG9f56WcfRR03P
IYJjmoGIX3UIG8QIiNqQn/r/TnCtj0yNe8ae3/PBPlxTcFwiy8qjZZjAv0NPUABV
J9dn/Akd6cztfwzihts2kRDV2wAokmsBPcZwrRzSHiwrf7Rfe/OXoNWaTzpHt/kq
mcxL/FI+c/pyuFEc6i3UvO1QkCfxl8X/ru2I4l3cZ9OcUK8qQweqMqmonjAOofwZ
Jb+KaPVuYQsiE+eDjznw9zkZSxetIywoF0xJvfRjz4p9lgI7ng/qqdIA+69fp7IQ
aeu02gHsQMLH7QdVyWV7fCeKj4cCywvJB6h8brQZ5YEU6CYgnWDrTWIGw+ewZdeq
dpFu0l7Uf8noilfHE12hyN51QAVgYdVq1u9Yu9UDZxhQTkgLioYnEk3s1Lr13Qvl
8qSKwxhZxjYqQKD4+kU50i2A7wJktErr2LDfT832GUk/GIvrP7TZ7pQagmp4nuej
OMhjRnYc6W65R3//+nna9O5/JKDXMnkciLG5D0JItrFZzEHzwEm7O6m9W15rraI2
eqpnvC9IP/d0XBfnkxflLemzwLYZ/0nIThmW1jl+MYGAfRi1kVW/FYfRXG6UhGXn
EsbnGF/7UxbOEjQOaUBeDks9RTigk1N1qA97bCiiXK8HwXITaIFKuiFNcRCZyNPN
h5KxwI0XKMvzkPN47IKDDM2UErfev0eFbr14ebBS+tAstXON5080T6olO4N9ddgD
eGjTLjm3EPnpP75TCvoKmtWO531+Xr6FgXHTmv2SHlfhakocHncecMRu/aDFgjKy
7WYdtJUygZKKZPicm9XWWgmclWHpur3TSoF2KtsgTPHNMUWkrt1xwEACLbTQpb9S
kt46UCThliYifLdqFRFhWK6j8qIGcF/RJZTv5DDNAwea6S2FUvChNSFZPkxfdFPO
4LHRrfVY9i8Vq1m7hbmwnzLOokA9ObLNwiyXZO2PMn2wO+6Q4aqJOBJCmbglZhp1
fHgCs43KXm421JF+BD5gZn+gaV0+w7vUVzT03TwFFdhovo2hKfV0jvfo1Q+aIw91
Yw74HRGS4IkSfqpybxAlRxjYuUhIv8EDMI5RS3bkztfmEAw21f5EFdbeJ3yhIxZw
TIn6Pynydk7+DRzydvxU4Nswn1MMSWF1LwQERilk1xtS1VPJY0oa0CUirI0Hq/RT
Oe1HrdvgBrEn6ZTuPIQtT8pMpyYF/+3bVnQkzTZKoBWAw1sPPjJNGZqUOh5MtnMb
J3Zu9dT1b6UjXK4VhTBPwqYjGsXwAGI5n7NTTtKTyVZqHpgtwR+/0Y8iCGrSF7Xv
lrIz5O4e0b9UFXaH3qM3jibkGbMEeWtrln2WAI6WgAf2uxy1N7DEBUc/xqXsWE0E
C5c0Nq5w9lPyMQ+sn4oRDRt/IEMdgD7oFLwd34rnn6DCkGNAjkRd7ecyfM1cGlS7
jcASA6HEdbu2brCHy+3dOd85LbCa3dZJ1hOvXE551j+cB76OfndlUGfrZdO3Clyr
IMVjFDKBcD+fokl3iLqeOlfUulFG2y07/Za+U0SObnio5MkJFY5KU3P2ngMm3pmR
4P9NyNI8Iz4lPTNo/4dCDlDXnFT0T8tJeSfocSVwJTvKVjElI5U6br65HMPg5O7P
nfqvN8PuXJ/lRM2ziXxT74U2Z+15Vbf2GoObJzSURy1gNXHtZ5YIQGoMbtvbJNHa
L3ybGWcdJtmL3gVkyzMDeqgz9caoGCGTmCMC1roPp2EKuI/CjbYGajIEI294sgfn
WdTNqv9PkESJQIIgmPLK7qwllLSb7M21IzNdOhJ6U8UBtDrBlcsqR8Swz337FiBC
V1AXaD8BerWzZ9UzAcFQmte0KqjGDfe0B5R5/54k/4J5Bp9/HgIAk5sKrzR0XvoR
yqj2AMhIDXzOQm4INN9HHLs8iD/6ugRxfubKtw1L96o4lH1ZfB9UK7UqLsD7pGMp
EmzvNKvEjic3mZZOcaBPkHXEQ0KNq7r2ORuhPECyscGUSkKVqRCweaYH6s046nVy
M5o9sXrKzW8Y71kTGF0QZSsnAANZk52aoVsdU5H0CPkA9FTspyw+T9K7/708HhK6
wbXBMCcCOkzZ3K2TYwx7I0HelCWUUh2OBvsmn7eRWtbfHrZBf0rLSkFknVAEA6s6
1uL98MvfqJmGCyuDzyJai0qzvcAolYLd/9zIG8aClEZsxcG8tyuA3GMzILbbwOnE
PkSU2Z02mVDcTyjIW6M5l3b/Kq3sDInujO7s8o4JwRD0SPRKvwwajWfLcGetLV1f
TD9QVzRUPGZ5ivyKTbr31oxRWxwDV5vi4br4IludJVL2Dd8HitKbGsYkipr7AaSq
hlx/jSFFALHLRzHPb+Z+a+M2dxtyXO9gSETZDYf0ZYSnZnhU/WXTl88XwwI3Vw1Y
8Sl5cLcwXPuts4xoBcGnBRcCfQH1JUefm2/PgTWq/Vs45wXwb0gauPq4+u6mzZQs
Tb9Tso1aoGah9HCG3eeDvsuXuwq8shflgYmMPlulEtt+65Nbv0sv0aeIcDROgORQ
f/FnVCODGbMO4QA2+JM3eWDeh8iooF+cY0q6pQg5Fjx656tYP1b0VUD9axkL4bVv
eeXMBiPEaIYOtnWqirUBCP6XhAOWQ6ytwOzQcz/QWUX3+/pWnevc0kdw1EzLy8zW
03gh08rKR0ipcO5WFFeuOsrvkFDRCUj2T+ctVsqKAfgiWxGgDvDEVX+ugN1jcZps
Gjxpp9nhGSVYVjdyp3CLy44qE17uImzqCV8ZB1pjWkfqT0RpJQID2vs0/y8MT8WH
ee4Hkc7y+EYWJ4o88G+lRrvawnkx4qANNiQXyY51WQ7v1I1O4PnHngvAm2Mcg/pe
x8sbCqloR/rzGAc8yF1WNWDDxtKASm3pJRM+kmOVfOQnGoFMX+sqQ9g0ows0OdTU
+yI+otkmGCfGy+al0cd57e46ftmKwMdYGb/51YtryXL4/IUHQzEJKGuP/7jR54Sp
uW3YoXGFJtjC/Og0d6Eho+avElxmHoZZEocuYbnXc6uIFUcDTnjYq2gZfNv7wx+8
dPDwuuGIip8y9zm5/Rz6xQ9sWh+4owCXujMLf64wsi5dpjqv9iF1gidIOZcntWCt
iaFH1MmH5TQUrDndQpJ3pusXJFx6Bq14+zYAMItrDqP7b/4uyGg0gC8BqqZM6CIN
uICOsML2+9DfuQzYGNB1B/KV0gAuflRv9O5eGqa2NMPQKVcqtjKHmJ1WBH6XGU5S
8sQ9p0u5SYQobQG1eqX3oTd6tw1mzhr4I6e7BzyCHA1KZ3zOGzlzrvU2lT+Xgzl5
AYs8d+CF+91HOCwfUTHWDwF6aT8M7mYaMzbs+QfBTaF2FH6SxQd5Q9sJvFnFWMwo
zbM34IpZh3aHNxM329LhisxFL27jyLZxN/jE/jPNi/tt2shjIXu+0LLEnZZWKrEo
ul2EAIlsnenKUEZieMFQ1mVXO5XoWYwNzpp9dTiUaWCjOsY0vR/pTEpbYuuW1/g4
wOYh7jFpTvrvsD6O+r1jrN4xBIi04ksS4sWyZCncIY6WUGCdZy+FTueUNS74JJID
YmD6LaadeQEMXwzJ/2XTn4/SxRH6sG1FsF11A6esUmdNitN3Rl5UMRpG0m3/yZ3d
dyED33l8CuevOEbTbsk1dkUZrR583XCUzqqhjbA8YGl5+5nLldPNcYYJKMkxDdID
AlIOjjf981bhM7YB0rVNGx3urMAuHPKA4wJqFVXFeYEE/jgOI/zyEY+nC8MEq7jt
f5DMp6hYZsgmLdlGWMGkfSx3TN2mIhrYirDzzSvpgXzzrL48OilqEu+CGWEmMqVw
3jetq8INsnX1PlgYNjNuqFRVjSvjM3kxfTUoVdjizUaV8L/pMDTNrRPfO6ICiSyJ
P7vyJBLyKPtSYoLSnyG2xjtdDW0owA+Lc1OnRrVztehO08vMKREejRI6H0+1T0qC
EKTOAL0Qn2k/ghfBu2DgkbZiCLXRn6Iv+l2K8JDeKAMgW91Ff1IxKkorcOo6XjRq
ZnWEkpEy08wJT5cV+bFVkEY6DexBVZYHFOTtiL3MjP6LR4GlmsNC9EAxFn8r1mWC
pK9WhLfIZHxrwrjlVxuJk9JC0tbyrWHvab6EWHIy+NjykndRvK9rlQXM/wgnadpn
GoqQ6HDlx/ukhZngO8S5cXJnTkY3IDnmFuupJCvafrNO5nPykdEdTfkogOx8gXpu
BjyuIjYLWCz6zvrTkpkCIWYtncTo5uIaj8zZGdj06bm+eU0nW3SBY5Ws2aOdB4af
U1tYGAobK+B+T+LWHj8J68R5c8AT8Yf5/J7P5lrgtduvOvaLPgM7lS3vmb5o/31Y
yvNR2yhsNfMeCLJ+EcKFflTdyr1ZUd/tBUEBJOYRcRtvLdSvkoP7E+B5vGV7h7zu
lTk43iJarUcZecEGp0UpzZD1A0b3YbOoIysT/L4suRFfbkELWITIsMCdwqYhc2kE
8OsadhQB8niH+8cuBJNV0YjCWOg1G/3Yj86FNB2m/jJQKytON4iygFs0ovKXc0mO
RC7hsV/OOiyniIPxibOGE7MGXbReARrx0frHY8ZXX5gQIrKvafAFRfP9W9LAoPX4
pbSFTjhqhd2/Z7yA26VCdHRFHFa8NylUUenOe2NUDr8kPb/aADd2i22B/G8ZCauU
glFy/Lw5WcNyUYxyo2Xv2MpZWMoy2Y+Caiu08W2/fS/A2OK2EDiN72cinLkKwpPx
rxWnl5mkxUcNfo4q1TK0zviJ/RlWLD6yO5oF+LXJF1dKIu8CX8kMB3nUKpsWkilu
voVXXa/F92lzYe08ZPBJqYMi7kr/DNP8KC/dVHXKbZ4XsUIMUhZOCflYLUydgCOf
iAUy0Zgoy1Ouq/3UTvToT/pkIpxR2bBKNd6F6ZWXeKcBib/c5eQM17+IDjK2m236
Mvr7ecx8lB+RvTubotOfqpRZHyHMvv0p3khuSS09lUS48mlWqFpuyK2UU/6H1Q+6
f/3m4ByVEJQKkhhcx3Mh1onIMJMOT1MhZIGm1BTjlgL1DG8kepqBT0KyaUsWecOO
YQfNxYtgG9XXFQe37vE4Z1/pWndACggxuhf+JGkLSTq8Bl0VNAwiNnyrfqJL0x/i
jvqXygf2GLDaMyXgyjIjF4qMokjq9fOZsj96EamwUEAUF3Zy1Auks2kUpkku+fTZ
D0dOVl0oKLQ/vKXcJHmRmE0fP6dc+cGpUuwgZxsCEIthavEOE9N3N4AT5PNEnfxI
FO9z4yIqaJqXFb27fqAVZThZe7Ih26SStUcvlBTVmpQhTHToL2mHi8C9evHoFfCJ
aIN5kRhbZ+j1kPa1YTcxtyd5I3GjK+cOd61rOnZrgi03GILJvrAkGUX2nppOcK9q
LZ1+KWLhrttkS94hP2amZcO9821WMke1O97pOJP7c7KcNCMeRYyozOgUYoKiD6nK
XoYHo+s0LFfUVMgunlrNKQfzCVP1CEUWsH+nZyeMcdmfCNUKECt4wUUeB4Eo7IEG
bwAuCxmG/mQmE5wJdaQEBZc887nHLDP+RIFjmsARaBKxMwmu5708d0ompibt+yq+
AFkTO6QfaybeLOFmaAYElpcJvnLf+clNsyqbgEaOnKcGm5euVZToxydQgdfB/Im3
eJvIVTkFEPta8qJNak7Y4memjXuLR6265url1E3W654nOs1fl+dlCxMMTSB+FGyK
8g+eXHmVs/uemmfAfEe/R5st21204rUMxsCMiY21Q1WnFs0WrJPogkhkAd/oo8lG
MoSixXGWi52cyfnax05FAF6qOPxqesngf8jrT7sQWCeWkcTO90PxbZKDPLoKxnaD
CafMccHoLGgNSytLm3oVaQxT3V3HhpUU3UWJxpZ8Xw4WSiA4QFZu5Px7I+qPfYP5
VUh6/ocJqqEr0G/MeEuDzvrp3riKZ0bVD5Zqn3OcmsRDsgSFHFQOAFCd5OQrwT7O
5vvvcygimbkuX0Ok3xkKKyjY/h8L4SQJbrwfAs7HRuHskodyJGcKD6gZYtTDEQOw
BHO2dgKF8xO/wGnWhnL4l3ij68ovhkoMIVsQUUddtiy8TexbgqikKx39/jjUFq//
Irw7MjZqFt313RaLvsjMKqiOTcLOq6C2pd0f5J/rOZeN+3dzZpwCXKAngoMdlBCp
vKrFUTlXVJj7SS85YpnPbbKy1i2NV7zwm4nw+/INaQQZgOEfbEQihMtz35A9kfas
GQQX3Uaf+SbHtaVsISJpd93p61aYJVmaGX07aK4zhCoaR96T5mNS3sIlr5Hti/Bt
8prR5e0ExLSarkohGcIzOs1ArrBcMu8c9XvK/jjabbaYMJExne/8g0guOXWZbzoe
HLT7NmA1ccdj5BfJdFgvxy+QfYtz41ctireETdSd0anF8qZTL5jA50mtHD/UGP4T
fCTkDS7nRCXP12inoAFfPhqCZJhASAyfTP+6YApegwMrHPxn2hCBfGUjGaERnGnW
cFMePawch5s22E1tAHtjG8cwcc885gtbqeyrydEEWaAT4HTGUYJDRNwaPsYb4kV+
/bIKC7P7Ros94ZMFh6XOXtNBoCXe5w2yiDov/+MlWQw/lwaTE1+1Rl/JgmrH0Dxy
EH76K0Ucoz9bF0V2+cq7KSUxCPfqYEVMjHk1ZV8hNgSnOzBggwNEvkbIOtTW9eUj
hSJuwqRqEdNmsz0mCRubkzXuOPpvGV07VsypRIgUsSGg0g5UyT9VXlVAfFPFqrAY
qb19I82VjLFFKFlVTBnldYuW6orycOJnkwKPkANW4/0ZqlRfwgNTe6TNls10Jzl6
raMKicfj0dwhHsgEWabATb3y5cdbw5Przjl+PMqq5ncfAHEPIMikRg5EwDCTd1N6
eBrXK/KtlMPNErYi4IE4tCRyP3Me/2QYSqE2++4eNvyfsxHPyoNHaDPRvefM7eAJ
LdBn2Y/TnjH1sTDcjm/VKEqpHJlDGgWMK3seIkK3jQpYzqB9rH4L7YDHMyUqHQWk
aecRszONecGYXS4z9Nnqtza2q+va7isjYAPNKWMcQP+PD8QXZn4SwcHFU83bX2EL
mMpOLNsHNgRNehbLVdQe/1nDvbC2AED3XxvZ71lTfMsg6vPApthj1ghVJrXI5Niv
ytMkZgvVHB0b0jCqFYtkehhYizzESK0hyUXUruKMeM4wM6rDa5TOWQ/CY4zTMwwc
LN+DtY9qtDSXqVPh4tWTocFP1KJlur18O2G+Zjj9zKaSeNr2W2EKPwi3JrZmKVy5
WI0uDvhjzBvN0igS7ofuytg0s2NCTVoin1ksOq/OCfa5ZYY3e8Lz1b5kU8ZRWWdf
I4JW6NsILsvuDmVKWQk0Vshg+xIduEpFsytSd4GJgYO83N4h6a9981jAxuHaR8B2
91OzRcc4Ha+aDgmSLSxX+xTMPHM9cYsh0pRQSoCmao0sQ1IJcNkmwK435bF/ovOd
JkV6L26xVVDn41hI02r1pbwld7Tb/DQV7h7seTjbwITWdJ9Ti//LwEjR7+T6DE4C
W60ipXUDqUo1nBGyl6fvONWARznkFyUI0ikbrO8ZczxFxk5YjOP640gU6Fp1TFuh
5bZxn4vRaUv9PVSMymRJ26Ov/LiyRQSFgUXh3al/CvV/VwZyghTs/ucpE62sQlaK
hEZz0Cr+gQqloIjJRWp+iKjswOgclPNDydyEDGAvwJ0fzrlqODY5TB1Wn27j9AVR
QifPkwwdkjcc0IngxZJPY/qFeylWbbHE0kgsxg+37xQW8un9VL4Qi21zPyS3Nr+E
nzTMFCZMN5ZLRCMvrWmTMHb28meSElqDXQR//YLGBOIf4ffp1vDVdXNFJcVCeaai
+DAq1mgn/tmWNv3Lxt7cZws9EWKpj5YSCFV49ge0RdlZdd2hbm4fUsEBUR8G1eMA
BWvj1TB1bAjp5vx6NQuHtKb0+RYuD0QQRK5cxvvx9hdZjtCFV4g5OVNpLzfcF2Rl
9Ct0zcD9gx3oCX44YCUw3lU6pIQrHlYP0sCPM25Eacb2ApFeBmh2XLBfRCvdTBWC
bJt6T+vlvwdhJ/Eu694ngYevBlgWAalIQ+bU9R4hzo6XrvEfPNTtZMqP1JiwGaqO
5ggDLZ/JeLpYoOGzZ3eggG4CLqJH1ew77axnbJK4GWniXzUfJUdFYLw/a0PVa+2Z
RMxHRcThg1SboPs6+LvvAYZe2+RU9y19QTNjSj6N4wEv07woO1sHNzGvMif8GRjI
yHhm543L5Ja7HE2qmGobPri5z7KnNuMrV15kkPqOkY5sD9qenaGSgkWqGuBrNkSa
TXWG13Ayy7GQzs6dKm+DuW9Hck6wC23caDsAsNgOHn1OXW//3xMgxE2FybVdzAdo
ViqCCimKewBjc4IVHjjAId8+rYWws70fJzhfDuGT6uvSSD89GkVrTWeKnUHQwzJi
6JICkBcpTeQWWefwbIb2RIWfvTE+Ru2BsD2upVlBiwUb/Tyx7R6ogQ/o3drxKIg9
RevhRHwLyBO71quBF9dOLN9qLXgMoc9DI4xjxnkJ8jvDNEvgLiL5M51DTDKrh2FZ
tAfA6jQVFXUU4iKFmVmE/6N/eBChn8kGgmjKrSqOWpAU3zppIHdaxU5ok4KxEmmv
/b9DDQUh9TmvhIlTINkvjKF9JhcdGJCRfnTghuHTfdduSo6CCosriWWq2QuX+bnF
arvfNBSb96UP/hQhTvNfma7aCijcZOEFKGyLvv0jPHUji7Q2mLmAIewO9Ay+p7h8
I/7B11DnyXUTOua+IHGCvsjr5WdNUCqCPZc0K8Y5OiX3B01MtglyHk7fozmfR3no
xoP/G0qd8lZiwe1teUK45EhNY76jTVBMiraDRb7g4eclOY7YuD8ZImTfMy8DRQrK
e6qNjECrmPWVSmuIMVhYwunWb94QYu4zkN91GW7bBYabfaLtj8vzqjFv+dWbufei
Sy4egPU0hVHmW51hgzDxG/9XF+e+1CCTiaCJ5WIZrTnU82Kn4xndkg4cwVQOEEtb
rZK/cvmF2AEnvJVGR3/NHOFDFiUwOd0udMu8aUEiqbOMeBqKJEVOdWeyfH6xCjN/
/EXw6GdosGFo5ULiJ6Lh6QzOkCowsIoOytXpjcQhPMQtIU80sdrXIHxZCDTyRY2g
ZCzBRjuBpA8W+I+zxTp+VymEdIPzdrnTG6D05KtfStRpqTDyNdiEG7hGyuEkTnOL
gA+UwJquQ1cGoRss112X215XCacVkYfgTTZ0jpwgvlNNsBVAHOZdOR4mvGRWY4UF
Uk+Iw5p+3LFl1uppEQjdYoHTA69iC7WT3sEMrZt4tIadaLIVLKJLDqd67XKcH92d
xEKEAzstE6RKDai0Erlg+5NeC4KTun983+uT2KRrseTR6uTL4nLfttn1AK/EBonx
qG/J6IYbYs0saca0HS2gyU26/Z4bYuwNy+RohHHYtmiZKoAfINT7nlb4FvG9MuEu
ESdjWz4SZWRvwEPBkHJplHnEU/hsDcBfeWyWt/ftQQOzCV/y7odjVkyPun2KgWqb
p3Jo2rLE8+/JDvlw3FmvHyVtd2LmIIA7Tz0K/z0EV81wWOZlpEGnYTzjwLOCdAu4
a2XZwcL2BaCZ2lEIvJ+FBbBOgM8fgpIywBWQnNAwN9gOqdJ3oNcl0bAKBFL7bO8k
aXa2Sz1eDT0PbVMXVW6BhP31gXxw90HsLJsiL4ZtlpVjpbjVeMCX+OtVjo8P7ltA
dQv7ps4uJk7MGYajP8fIucMMuzIpzAMPlB3V/eKe7VWcLx5k+xFcXFz6XK5E83ys
d70vARvl0wGvWZWoF0NDdUxWkqJTGg9pduKAyq3ZrUZrsctvxNYul8TSqZuzh/Nf
D/yRozD2EZHcg9PuOCXpRD41g/cyApYM0fbdrq+m9vEzX1ylNGfWOi+WJvyfMcAF
JGjQTW+eWEdI8KqnJHOgNCkCiOAsLyb7w0/Mhk9bpFxaLtrpNxIK4tT379CFe82r
XOV5eHbe0Zyd6dOw/aMkuzblhaUNyjWntFrBKNX56qI8exfjPBM9XZ1gnqiK+WNM
TSbOcqpj7Qpnj9dxTOlyHZMevOHFlWIhJKZzC84xRRaxIellHTmJlKmAS4BmoPrY
Szu4K4FMDL1A9xOYNBpaJHSMOVt9I1oIOACHuOkDGYDIaVhIMue5InnxOnxVYgEW
eQL30bdMuw0hVzjdP3BYK8LR8bvMtQHQsnkA5cOiHlYr48nC8nh+zpchYkwUrS9n
KipvrfBIa8t0JFcv3NvlxhVEcBd0dC9CV8i7qGB4e79gw3sTFAddtrytvBFO9GGa
7zzM/kkifeEYLPtf39E70uukvBi9gmD/s5cWbIV2QDAv7P3Tltez9YcqRXX6njA7
O7FbwqXbt7zHGnJO867xZrgZ5DzHpYhQA/Vy7xTaoHEZL/oUbNi4jS3ZYfygZQJ8
FqWjxUn2V78uL8P75cIGiLmzOdDzLU4Nthi7V/pjsKc3VqXpLQ/Up8qugpxLYpdI
4Z6c7ES1JBuymZIzkssEcu/lssi9WoR/mUh/UvKsdWllXVy+THk4YAUQq8vO35ip
cI4lP0BuLW5MgenW7/2O90MKlvf7z0TFelg6Ey4E4fblxwEKo/Y3u3DastUINnH8
R8zFoKr6AOD1op8z1jV9dAk1ukN0YN0BF6vCQl2fyOkzqKKEtMcaansTuf5KCNqZ
LqCi5/uiWpAceXV+cKPmRVmZIdkA0eK6r+83cUfG2C9GePum9PC+Rk8RZV8PJGkF
SJYsTyFjdpLo1DpSw/liQe2nWA6fzU47mHyd9XoMHOJ0y0DQmAO59izOT+zIZLW4
tVfLG1hTghB0uMoTf0LEJoo8q1ZSrkYqqUuQd3d/ATuU7gxbhn52GgTDpol8PIAC
bEl94ZUT8rn/S47Q7OfIbSr0QxmQY4qn2mf0WowORXcceoks7HQjl5eBIRJARj0Y
qVMGm/Ph6UzFHBcgVqscpPZkgkY6cDhClaYMJMp5enSvLlnRGuMqP3aPMqCIXJrg
Z0/ZwcMvtdM1D4fvxOyGkgYda0SgDOSqbS+KCmjb9qjSoBRMkXsNh5APkYWb3rVI
7pTOByvEsghUbS44LqrFrvgtLCueFgZH5py7KVRJSfV7v62MlqGSW5i1TsXHmjVy
QfgmZfwlPR3CLAFyu0UFqsCMsvAYU6WvF45J+WpzmH8AMuyIUA5Fn5rlH3/yk0FM
YjugYJ503lVHNFQQkLkLozTQl9GvVdvKZc2Wb7cqns4Dz1tyqnBSogxn4/8cYLIa
g3Nkv0ZQrVpaDAzHsoR/AOTqTvMZRLkNG/uuPllVfnyamkDDOoDucMLG243NNpEp
YoYmGPZeDa23xQ9Vq7F0DcSUWeZAxh2Vnv39uMJTFQ0vZ61mp52j0XW9ZR/wwfIx
/qaiV+naSSgl88QMnqG9PFDF55mZ9IL98H42gP4RvBbMbss2+QojZfQjnN6djDKT
BehZtBzaENkhqvD85JZICaZjhyVFTqbsqSUusTWepnY5TNPjVM0Cqpe3FEGnDO6o
NCOlsvpW47slzJvTGVlOXtosVpE0msA+OymFBGASqyg30T7jNY1/X4bXaZSMo6RC
5XqJDFDKUUGFSh6wzmdixoB5EUpiJDURHjNmYgy+Q11zH7IKIIlOYNsVvy9Qpith
dVI7PzHX5aLNCdqC2ghGApo+UrAk8xfN0t+vcob0SMrDv1AG89H3Xekw2BhZ8hO2
pizfhrzidStsdLObuQHDVTBoK7LyPn0Gvneu24a6ZisxUllwZlWoJsKw46fDNlHZ
EPdQ9lQZobjYAC6FIA/TTzakfqYv99ALvibYcFz5gZ8f3TQA0N1muTTtmhk10rAr
vQSkQ47qxmZ0EpOrk6tgXXG7N1k2TSZdKkvmtqKWgz9s/NQciWDMKSXW+Ps7r0So
ijy5qd22Sa5R8vYPVFygFg4DLE775UXp0k+B8N/6JoMOtcqKr7Dfk7SxZ6EKOS3R
Y3cpF1MSdMfSSjDQPKBlQhmxDmJSKXryOVJp3qhNDujMYeHirlhveGUV2DFRmr05
qgJY31MJmQS/9pn9KReZVFKvJE9NKOfNDHa3unSsoQOjeWMrBO5wOt3+W70Ti+ag
zq/vKXEcXwW97u90M9lNdjqTvST9QUcwQgW03XWylc1L0dSu6rDaFNRghTCAx9Fw
gJ0z5X8+1uo2eEKccXiNE32bQLkz7TQKT3P4fBRuMI8KY4DXlaQpLEVPU5w2b4zo
p/QSHpVPqt4coPMpLJnEymAyh5AwZJ/vQ8BczifulUgoDBTxAt0NQPa0XUUOc7JD
F/nsu2R1bV1Ad3V9KlM5083RTuTizVAHP3OyFwxUZ99yjUwJwlzJD2vDEv4D+4EX
vL8nNe87r21kqixAEO20Y6+k3aUDcN782EAGYM5bek6izb2TciGAqS/qnSMscChE
gV9RoFmDbXCvaY98ZflFYx+JiWpyiJU538lDV3QMzMQwhTkLCqjIdcAomZCapAv+
9mbM6gCrtbZSV6AtrZ67PMVIAu+hLIHQfGdVMmt5hUPHAcnsjGZsctL2wGUUW63p
VRfab0gsyN2ikRuLC7F0ZAxDTkN2eSy6Suz0Am+AvH225BJJ/d7g1zHWCR66ab0P
w3pezDJfZQ0i/eptRJEn9iMCLfXqkl2Woybup5xA/ejRX3tw11AN1IR0VojHFSw5
fH+aLhVxlcit3qUEldIES0eO20V7Qhk0641qJ+UB5+u2SmvK2C5o/Nq85wsZLEQH
fTPm32Qi4Zbvgaxwz03FRUUyBpkko+msFD6Ly3y9+OQm/W3K8Z0dudIWcxIpN4TY
imctrlOllXw473n0dnsRdek4DwQBEBW0hRCuzqDnyOinuzM3PDklAl29hT0peMw/
Pf3qeE7rofcw06edOeWbrtH3lgQv47iwuLUjtip5opxdU6qeIXERUktAonr6Mgwc
Sx4mTczZf+emMerMKl9AR5GzZKHHfUmCtjnPYc/eAkgmAi7o/XtukIzbvD7h2zjv
wuxi4UVbnXJvQcDsDb5ffBbotiRili8BhXNQLUOXkzgtH0hvUJu23ROgUn1mhYEF
2zxXkYi/1QGJK+hlvfkPL4uzls2FXbmb3VU1hv1/JWxuZwSJfj0utl/wxdmVYfkS
RcTuxYoQuoqZbvjCLn1LgL3TFQbb+x1AoLIYj/xHJWPWLuWYgidTZRD8ZJ0j21b2
d0QVZEjB8Z620fZdF4VIjucpOmZSe9LebshqwHgm4jKkSWth4UFmTY5aCMLwtWoG
wZFs6OibTpWXymEZHTjTffeLtV80MqC1mS+mwOywVv5XF44VMsM+A6eGMkGYnk2r
CvulRVC4mF2xjfPl+AdarAqkJEwNiYROfCNfVn/iwmAI+kbk1xuqxZR1DA1Jn+7W
iCSdIkaaT1NTdQQk03wuKKNEyYYUJlHwQfwFYmtwY9ws4M2YFQTfpwdb8fiHzx6b
H3EeY9Iac2OepiuPVgTlF79lZM0Ug7fqgXCBFoxZqnjJM36vRKsB/x/ZBt9wdbzM
jcGE5PBkcPZhbtK3R3/7dRGHsxLucMgGSMsJHaBkjQez1eTuL1u4XpcUqZTuzKIg
qqtnoUf3FhvEcrJjjmdf7DKWIStHh6OkakeuxpaI0B2G5JmVAvE8cnm02o5Kz23h
NL4b7fXT6ZMnsEFic1wCno/u/UE6h9InJDAga3rtZh8h+tMkL58jm84C8pjtbip0
TYQ6ijvZq0+YLzcmwm7ZDuUSHUkwLMIaZVTFrUhxZDXClAVKcNKO5gUorM96iBA2
+zcTTdQrkREyEKDZUxIi9ANisr7bcnjg8q2qy1lgprQGy6Owz5h3qWalKmT8XFME
+xPc9lqDNhLtEEjQn8vkBgY2NwtLnTZjX/+YSk5lwauJ6hJbsoHVII1WLFE3qGBe
dKL/rblnHvEVcc1v/6ScPUYeUNsAIC/Kg64qEbVFGomujEHDdRS9ZJHGqrUXnAdG
aeMGbQo2piMiL0Sc3MEiLaAH9/g6ZcsVGcI/YzAg8HpprEiLowLlGbOyb0nDA7Pg
K4zp94FMJS6ugNt3KUnhNKpFEpJpRwkbOnGHl07iWSLfMQVpN6lm4dTARsLyEPAt
J10qRmQ5/jZAbh4/t7XJwAZCa5Fnu2vwc25mdRPGVQa98dzonShy5+wCEfvYo6xV
zT3kc2zlp+Y4lWfgLSg0spG2jjNduRr1ku4fWpjpwxjjpdaBDhPdAhQsPBs+B1Ly
QbDJ13HUISYOc9Ef2lZyj2ZPxPV/fNOph2lcQQ9UMWfTLCtSlTuYQ/UO3ejXrGc2
HKy4UKUPjhspNnR6NtwOKy4PcIKPxn+v7+b6zGFl1G7kO64YXQP++NqcUhPmDje1
pg6gmj24t55onBWggw5mFgswPIHTW++1abeR8q6o7cmi69/XfBwavPtwp9y0eBJ6
VclBU4IkG2LTgiuB3p5Qj0bDbE+0qlyJHvwav+U6IOpzVNfHFuZmeNPxMVYmWPIT
l4uVs3RAPqTBsPxBzsyuUWe8NMaYZ9tfiM7nRUd40VQNvvEIOpSTG4aWB4CUI0PH
7KUQyaBspgrPW2wPUYdagG0N568gpNx1dVDQfof4O0uOG1bH3XzAb7aPY0gGnSPf
O4OTBHJkmNeoNxRqwINZUz/O3MBdS3Lbja1gWQfosgske5bAYu6KV1bTSFlKp+Ac
DomYOGv47Sbm016FR13x+Nl5AUd0I47EG/HU2JZ2Uk9Aucy1vswEiNfW4kwl/OvN
LX3Wa4yN4v6IzHLkc2GW9jxWhHKc8YYB6oOPE9u5uYap4GAjEo5qLbGN96cUDVFp
G71nA5xmg+Csoi2SCLGY8PpH8BnqkGd0J1XxeNmiBnLQt99HHOYz14s/AJpKqVfJ
51laPPaKVNUUgtehFm44H4cLi49BT3iF+d4i4PzLm/08KKVzsTwHGIeY8diOV4ka
/CIaBbWfMj3WectnYoxs07ZTKPjLOAICB5qakz132IUruA4meEMimvfTFz/JcRtf
lAk4zgucynv0ovRHz+5uOT3zh653mxauFqHFAZBFWr0B6YEucuCnLcZ4glnXuH9x
vFLfa0z0UMMtuJmkMEKGjlNjQNKf3IlrzFM624R7bGLCOozRpT6jQI30Tvb7SO8m
Qeb75puJtzvXNn5JThKMtbZtWKUXFyN6lwe2FCRyxTCahDDvYy8nf79xxsd3sN3d
+kJbDAcdtY+K26RPMPRprLBZYsRXgl8g8yrOkDcT9Cg4qsg+N/Uatk0dapBz9op+
wr74KYq3dN/uuTWug2sceDvXXaOEHxJ8dtICbnGA2OYfMKBQLHMOADTm++Gsv8FN
pyF/Tj9QLLQiNYjqkYrTcp5jb99Frn5lrf9BjfWEsAVB8ZND4d7piOSrBPXhOwNd
amhYkf80I1rwxXb4EWR3951nJGKptdclVuqHFldsKDPRDJFN5ahxjThar3kK+Ym2
DOmbL8EcOliLUgciYSKK3K+hq8Dvu02KWTf8CwgDXZdIbBpnHEtbHeoA1HVPPN7p
11GIkd8/Molf6McRp98BmBdgg4DxV65rm7CORhOmBFgOWqUbugXya4wlJVVq8V4A
gA2EMM06ItXfdYXPyQv54i2fjbvxBDECMnVOz4hhUSa2+3+M4M2e/ayVAfxujEpy
pBZiiYS3MT21odiHN0mmSyfoB/xC9vEECzMqGn339Dfyu/lASdt+jhiIljNbdjuT
SkfRTPXih2lUZGFncoc/1EUJpdIo6qMa2iLEnvHXIx+4rRjvdxOzfSsfANwTiegp
a+ZYcL9v51QiYl8ix3/Csl5PvRn4HKttqUjuS4a6wv36iv2X0MwJXhNUzxT56TbP
E99adyuRs0uhy3ipC0sntWXkVnos70RoLpMl+O+gzbeULGPyUDcnlqKElMIhAJTJ
kbRnP5DYuxv3LiwcGhIQVRxPx+M3v/NhJJ8kxD2w41ww3wi9dOziKI25WdExvl3F
P7mFm3giueBN92WrA1si9S/lGvQj8C1FbBFZok6X0Wi9oA/+DGIxCA+hvpMAC4if
1iURMyrVWlxvijCFrSIB2OHNcqWd8kMNFfXxObJTqdf6LrM+7EZXTb+xhmkrFMKb
jfYo6Anvn7cRpx3zr9E9fostUh7I5crUKSYz9afmMVvDRIBxYuoIsDaAfbFkspfi
yvCdwhdHMsqUV9pzTILJDQmEmfT9cjNiGZBPqvPPFDVbFFqXSSNQX4xdiLA1+awX
PADHCheusdq/ips0L03L+YzfRdEiRtCHCO93QkqbzYZLVb9QG1QdOEr9L4JZ2BKt
Tna/y0B/VuFu8LK/g8S6Q669Qc8w73rTg3uSyhbWTzBWizmUJqsIRZMnZJcM/87V
xb9Yg7DWw8C0J+Of356eORKl9Jy9uudjR/vOQ61j1meGMP/dkhsloSJh0Fh7EsUr
CrepicM7B6N1RdQdSgA0Zx+LV7OPVlJ8uYa4ndEfIVKuietqrqwwujz2hgHryazR
Cq48eLCOrecx1RlVmaTgZATmY6wuPGtBY1MCStkkWRwemOFs7c2d/8wr3Aa142K1
XNJjbqEdulAbjUyb03TZAPzGowJC2bh5rFVgX979RiwjGg12Vq4KN2c+2KXF144c
kAfOjn1GpBXDhjd4brNsjcb40Yq3ytt7k1uRLNcG0zBDrhk7iRadVmhOynOzFntL
pg8bUBhd1Z/hO2qiX1pp4pu0L0fN7nc7J3+of+AmMluM7Id+OC2ULxh4AGfSMqPa
phVmX9PN2PS0Ca98WU8+mP3J3NTQ7LVnPXLD3y1+gA2N8eG7Pdz5XnmDldB08Jpm
CMGkyozPH10hozMsuXxA6jp3GxqQ+mlH1qyq6rpZe6I29SzJY4PdfGi2a8jTVohf
cphLx1B8HLX5j0zWDnqHKIVBF3QmFKntpXyupjwFaULVUc5dO1o0dAxVrmPeWnDT
hmNKDlWIThcs1TKcdS3hgdu3k15WyWO+GOnEfMrgmInKx0ZxxizA4YvOAXCsTNOR
5tW5ZlBba0mF76RC1na17ixHujVa4euvrGl7y35RdVxF/7eVqaZTlWOe1XW6/xcF
CY9xuwcPA9HGycqtgipHZyn8i4zly4BSuTifNUxd1BLmpZqL/I9oYIoKP30CgvLW
KHmLkfitZcpmNXXi+7PH+6GoE1e/hIc9jNHRlMB/RNDfB60hPcTgN+fwj32KSVjI
XOjUtxselNsPFS3mvwpMsE7qnhPO/dxJOb886q0mDRdfx6BUWj7ygNJGWS2kM6Pv
uMMlSU/iZOZbOuVKka33U5d9RyaX3+UFbX9gCDzjR6lB4i3bsgS4TJi+2CuNsXOk
GAS6S2ImTIJTqGUh8/wmtUSc5XY8/xjXh6wvX4IiH6mGjR0+GrkvkLYeMepR4RCt
VFPpMHq5ZTmBTeJ24rxAP/sfrg5Cl+ZsFYhtcnCwwalPv+ACk7kfHM/gHZkInz3u
4fFrnVLvm9Zo5f93TfbLj9F43sFBuSra+QW9aU2ifxLtyZGOKGOZwRfuhWKon4me
ezLCQNPFkzE/c6LNcycNWkuAWOBl48rOYMAlJzd77EG1F46/810iIQWE2IpSdbTR
TmjunV0ApPqJ4QJRPN1zPKA8mnXnsmJ8bXqJrfFgFzyFNtA+3cWK9uoYRQGOYjJ0
N+kL5nmhZ67pahQYvN1t42z3oUDNcghdLpy1KGsKu/XpoNcJi/+o5vL+yLxuzTQC
SOrofaBK8rP1wyLLu/SLHbn7ogYu+sBqShyf787r2ER8sZSBS8zSD+rDadHCwmG9
nT+YlD1R1Z63RsLaZH94GCihZpqV2FRDb5pZ/jmCn1KYAlF+cqixSeZbc2t4OWPn
bHs/Sb39ZY4In5JUQmUqWcEXmRUxwON0c4mHZTHOWb3y2XIjE9PTem7OfbDU/bZC
JQqMr8Ldskr867bzyKpZQXZG5GJOoKcwpSHYK2h2l+jaNAuCOSflcTQPioFs/Mh/
JCfk9sBMbQ9STIc1Y/tNBk22023FUcKz++925MSfOKIU0Q2V89THs7KKadVERnhN
VHKxcbK5BfV1MqqwyiYtXBSCTe2C3TcuK553jEtYqFh0lCs6RxGLaWeF4cTcVblF
lzuhv4FbOvN46JkGL9mAFZ4eBF2tFM/d00rRN08GHftSh/IKJXJ9qMZgewLvNL/P
3unt+X+V0nvyTKr50R2YoaIOAki3DhZ0GPOv16HpfZwrQKe3islph9VWqsG6fXzl
moEK9LwCBTIi6DF2KQViCQ9VDnezNqSR8s4eLZWbLhddSS0gVwo8ddCLXC3ic9Gg
A9Bvbv8wdrZHnFXFUpU6PpHLpebW8cZoq4pulRMfwSm2aB9D3I3zg3ALKEbQVng6
mdq7kPF3MNaQH0X9ZTLBumLe7vZZgTsTsDP0uhw2qj5t/wOxz7ujOkkIvCXWHYNJ
IelmKX+gEutBEEzy0rPNnDwCQKw6Vtcw5CYZwgLPESVqwCKTt7c8CUziQkWI+KIY
18OzhVKs2oLB2W34+bh+GnmvogMSUikjmS42Y1KqGSCcuA+n/INhyPI7E2l9IfTq
fV1FA8AZ2cltMECT2OmORsgOCOEHhfHo69fm7vuyVfOlX3Tm6IsKY6aTPqI10GpR
PVpJh96SfnF6RFXTVl9q2IL99b5igmfiwYzOVALHfR20Dek8yVF3l00VmBoN3qHV
peB0VyLLHveRDRzif2VnpeDuy8xEBJQJ+JZKH+Ew3FU9hi9baeXVCMfIpROmrUUU
eijayTmfSn6cpHFIZmQbgrnuh0RN/AS1Pm63cw+GrSUiXSR7HMTpe0QI9JRbn788
XANloKN8hbhFbzzZBhurCYQpK9z2SZ7Ifh51+rHhxNEYu6RNWQsdBbkqq9HrYNdp
1KY872e1IUNnGYenA94nwV7s7C4C8YjhGJAGpy89Za+94fMm4lwHfgGdbV/VW3Ez
dOvUIDyc1/+sC5xSKifsuT1DYLVqALQAIukBRepaEJHPasxohTFHaZXAN4I+94t8
EzESk1NFWhoklTonVB0edSndL94Su7UI7j3SBlVRvaAtGSkK1ePNRaOGkkZ5GSaI
nvKrECOFN9TxPucEwi4IUlbM5jInvcbSaCb9uCxqP6gNDsZxHMgVisF2JGE46y7o
XyhX646eGCQC0WbFuadXS9sa3EJwigchw/+T2KgIBwiWfYzNq9CpBWVhviXCCBHQ
h/p07N+16FrmYzbLBXoccuLjNKpfTJQaJ+DDDqfPgekkJ0b7vuj8xmveAJigg9ca
pkj27Am8dtM7AiofMES9V3fRCs3oWs9P0PrIgWvCA3V2Pskdf2czh5E2X5WCw0zN
JDCATDSsXxlPiekv1g9EDft92T0JC1WJmOE4VqYTcq2aBNkoLv5ijiw2O03HBxr0
ob+3eIFFgVupU0AkP+P+jfOWQDtVIKhNLXbCuhX0q5HtAlCTOQM1FD6Dej1dsg02
0IU1PzeVBD+tfVD9U/m1N4WaRi+s2j30+pJRomO5/uD1ukXB+IWBYWo83jqPlLHn
mAKkQ0FDaPSYzaJqrowgohKR8lX6xM8RF3e1/rz9xIYbicNf3LQ9HKIljdljMBbs
8EWp0HNlvGE78yTNYoeSb2kdWcQ1z6UwBnIe9RBYLnyt4FH8I4yskun7igUkkIgp
8sU3VtDeZe7BWmpNqYUD8nlQwjBaFo/ADNP542BmuObdUjBmpJmyDXAS4GB5RyEo
tzhDkvmhY/xG9TtFh9LQD7plyt5juRCnz8BstRXm0syq/tNQBMpyvBO6Lp0477eG
LJ6lU5qj1Mb+pOuXVYXzun++9CE6R4rOV9BHlgswvEfK2rLvCSvVwX5gKf7WllPo
bTQOCpyzLnIpSgvEKqbrC0JxnCdhQWCkG49H9+qAl/kYYlsJxEMxsXpGnf67n212
EDwXi+embLE4YsmukbqWsGSgVNe+Hq+2S1qMshZD00bt+Ws3NSFdGjqrQ9jfDjXb
nzGYOSz0LUwxYik7eDifTWxmIYWNHwHImtCv/8aQ+Msg2GyII1j/7RTxJh1+vgsh
wQ+eTsyBeIxr+d2N8xUUHxKVj4IaDf531vcsXGA377L+AClyi0mDQifhNYNooxnQ
kPkQnz15n/R/3FgfARzP7GpWcfvl2BdM/abNjqICUyu0p04Nn7kroyfhF0HecB9A
rPIBsj8S2qyz6XVgI83qG40q0o+zbTYhlWCQX21sWa1OKQQb86thX3E7lbUl0xlw
Oo5MV6gboZsAM6i1H0Cw/ThDW2SiwNN29+HnHJO1fZHiRw0uPyscjYIHHbVm2l3s
Z432wqVGN4kqfLpTSwqsmC333+9lExl0FI21762uUgAFTgsnSxbLi6JK5Andke5Z
HbE0JArX7zjgI/OWP7Jb8B8hRwUa6cULMyJh4zMZr5WbeCjIBjLwhE3hOHjfxZ0s
4ocVW/YGyXVlAZmrOcaKiETEy3oGDwSJI349N4PH6iwq5RgQvASGVPqketa9TrGU
2GRf1d6mAcCTpANINI48W37LuqCwgjbhrgvaJH9uFNPpnxKwV4zgjbXS7Qs39D3h
u0p3mlDygIlbr2K/CebvZtxN/kLFW2MkCF59OwyHbQKfE4Y8XqdeheTAJWTq5fwM
t3xNZBAn1+LxEaaN0snwO1jH3P5vM2P1QBtEYst5kdbLzMY5jr3+izY5xmNvRcyu
cErOj6xZuWP9R0ucHaOYBO3rhFOzqxRyjYKkKtp212N/wkLnFhqr4rmADNVd59dq
avqtowU7Bgm3bCsFiBe+SUINb29QRhZ44Eq6LcXdO6JljIrME6OWfEvDrvRQOI8R
PzxCCp96/WBmpOgjhzEYjX1CumvU48zpzl4gsw1RBxr+CpODSvoVMEqd80pxmesq
zm0C9syiaaMjr64F7tX/+M2pFHXTBe+MJM7/t7+Qti7rqY9sE2KXlOXXdHvQoClz
E4ekXRiQkpQU21BP1swIBlUhOkIhqDUYzbckPbeIPFMu51YAf2MoBqGjj4yCdSXD
Tkw+Bxj110vwSUxxYwe5shf3dRenkwyetzCD9EgiI5l64BMl6J50XJj4ReFmYxsx
sYavO2/TWT/uweyqoFn6YiQlA7dz785IrXdGy7gJYQM+gD59lxrwUYqE7apdV02/
BAx5l+wZHrLtLZwXaN14IqAOpsGvfPMBNnQYb7351Nul1nknWG38bqEs7KGZlzH4
kCwYRIyEtWbNmA8Ukp2pi54frPLvlj8vbdY5NdUoOKVLAP7bIhh+ZPm9dHdCnsXV
/DYe1/EwnVO+kW2Si3R4yzq60jAD5cselJEIJQoOIWXld9kyP3rKJjG9/c/FZcPO
5FztZZQS1Kujozp6m673WFxwSVeWcyDCVW20u70hLrSbayTbkwQ3VCDekkXHbZZ+
n0s1N3Nn13Jsyq6lk/gZVqXtsSQ9bVoGJW6fT7ehufF/b7lMCI7rnfeTeAG0HT/Q
wFaXzZqUkbShPBVI82bTXPV0IBeyI6F2AWdLRS7eUvDeV5N21Y+h7mudnJGzna7Y
82tA5CmO/D7Ep0Q0l+X3oVD9Drdv3KwixZCT6FaIoaynmcHOdTzT5UnpxXJpAGo7
zuQyGAXmfXCcFnf+s7VcjtA03StjcyuI+pwS5E8VSkDEuexKP+ugrYwVuk131H3D
9bBVsijbsW7/HOBT+3eTyKRD051XQe2R8yFZ8hInlhQWTOmTb6h+ZwYRRXWtZi1m
9xlYHTMu7rsPGy0nZLJAkGHPyOVlThz/zHkFTwcMgiTxXJX67e8WG/CDq0mnmFkf
XBZj9RODiTwPYHCyy20XLtMW+FU9Djxjz0Kb8urKda/F1E03ZKDDkr5K0w5ravKf
VGjcADMHubtrtBEukRB1ROuMrj4utF6/VvgQybbjGpv3lN/oUqnKlF/9jffK03l4
dwI+iQEwuPRO0JVQCMGm4di8tGy3TNbPX7fbRysRlQdHZKTyKMLSHwk4zo8eDacK
cjVTYR5qBiCfUJTa4s4KV7IeyI2Jb/uibhjGIHpEbw80PrERSqbulDQyvIfLX5Mi
YUPySsgLh8wgpISELQDBJd2g4QFoV9SazHrF2Exzs+XuC3DrDzDUtjhfP89Ds4R1
NxxRGS4VnaJAnzvaLMn51H3XN70nszLF+gGD+IRe0ZpBzCFsgUtoIFjtC3XpAZz+
RfMnAguGrS+fIjIJu90J3Tc2lZdTz1G5w/q38HgdVj/EZeYAdlBZ+UUxEOljSDvH
jQsG1oTwjT115R9g8GF2um4fqQl3FIA7mZWM5GBUVMNhJj4JJ0hn89CJDpqEq4bM
IK3kEtZ+xXJlxasMd+N0+rHKgigP+3MAn4agumMEFMJVvv57o3rZS1Hk7KfVD32A
U97UkTL2uBQYWD/D7G6rQBS8PLm27KGtY37ZGHvaPeQrKdWWfmfSyF9WTj5N23cT
9oh6Scur+HpdNdr7aHtTjoch0PojgAA3V/Jp1MkRt84AiW8i4S3QjdSkbDjj1Viz
YmhG7IXoo6NHZ7FPdsvUMOnq4PmpnsXSx2Gliu1YcQPHthqahprcHZ9yQiBIt/YJ
mzC4W5yX0vj5d6KgGIGK/O/CiH0bpSaCqKHxqAuiJR6FAAHHROZKIYVKAvd9hWlT
xLOL81EJnoaCkPPyzLDAR4F3QFgcLeuvVZe6ezSkTdciLtXHC8Hbe3DsJ6J9EElY
LKsuETSksryU/BYIrN2IWwqhKcxE1yt2wA7gyrar96dZH8w0+ieEOU2EJtOdhkq8
5lEZmM/6ScrG7GYhHOXnkyzH+yf+mru6FgBWOMCRBiUACTwEQj5QsplPw7E7jnPj
oRtyVe3LqVlA5n/fdFLe3a2EbjuU97KHrreTby3HmnHkjDZ8R6f4Nos/oXvIAqZD
oY6Foky6tVwg7NNcwaP+gorobVAdXX4dox3gwva+fRh9wCpbC2BJwfZoa/uWPnto
bud9460UUiqYfQPepDkyv1DW2XgUKiYOTYV4RkFVMgX9AyRZJsBRvkTsGAEZOPeW
LSdOcn7xj3yfQ23Xf1wB6oKhSoEe/y//KOq2R0fGqbhKB+gVevkukDCg6ftTd6zZ
Hzqk8b4yus6z+Mk80k8eBsJgQFkhAzBPZDnNZ9V1UizQyoPSx41K97TT1L0mFhTM
Lh+syoVHFRn6j/NKldmbBZ4NOLxwonWOZrhD319j3neEfLbhqmgXbSupmKwUX+yz
/Frk+5GENaKEb26mPOZk7xh0GLctzW9b7KlOfvyKBlF1zprYIR1WRtImoCrWPCz5
VEjpuHSqJkriGXTK5XjgcePnOflveL7O9roZNMbuA2Bd/O63xaPtSuJs0xmBWhnY
KwqDi1OlXuDq2YHpZZbJ2TM1eXylWK9jbN0AOPXlkNrVzBrfgpvBdT7j9eOFNXcd
H3N5L6ekRjGfvVOxZzE9SuQUy6FZa3u8NjlKogdhhOLYxNck2XCrQwQHm1x3HRx0
GHOIxpgrKlTWHPd/DrhDu3Xqv5kc6EgSN6RoDXV+ELQXV11lsH9UjLJSklX76Rhk
vuZI8BcHjYCqy9UDytzblv2ChEX1M+XqEjKKA2F7LOM4MBr8IqGgmgVQPHC77SJV
geLP2RTrJzzYmsfLg6MR/VvYe/cS77EjWVDhCMwTh4kSXcb/fuV6goFZwK9IApnq
vdcd76nZw5kmf/Pm4hlGvKoHIpYWaxU6fpovvKlO1fdHdm6gRx268hSZBPsYkgjB
9LFlCYpSRvkpG1AwVGoZKCKuBsNo1jXrMgFRkr46jg6/rYQVcRV5BnXH4me/i9bv
9UR8bikfkhFSJQWTbyC/VAMr6SFlohztjM2fq4mCSh6TNwEqHDRZjd6HXP6+Ma03
da6S+tTCVi4rkKRpJcUTNT5g+R+RaRCutYCdQYiCWwZCqD9YdXFzqgcV3INv6MeH
hXZ3C8PmH834WSxgOPOaIzDfHeooRry1INKt51Io1vJh0GLrWOuUnExyGMX4/YDO
J0+H9r7BrhT/mZHPisTlTRA1dsAR70ehVHlPkfWxMs0+IgQ9NYV2Eu/aZfsCbfpo
Uw273apu0nBXVtddvavzfqSZvxaa+vFHw7U3t+Thpds4252eBqzj18Cqqi2MMEm9
WkuvxusKNswkPmE0Cu4xN8zaVy1nH2tRaSyQj1c4p6CpxTqhVy4uSJ2XbOEp3Mat
4ESi1OBOxCo1TaxZCzQ0m/9K/gAsB/m2vLKZnTAgiPth4dDrHVht2Cwida5qNFY5
UoS4m+qdpTPrGp6JQ2AkE8RXFk86gorIoCLmdht4Ja4ZV6a7y6dglSfwCL1yn27p
NB3R7KsjGQePZTeudyuuDBf9iDzsSBIP/vsMGqGj8cAmmZLGFT3SbqrWBGvD0i5X
YX63EwFe3Ak1a2hnJK3eHVXn8VMo/WpiUGsfnDA3flA7PKYS9ss6jHcttZCU9irb
qos2Ss05bAovID2Zo7GvjIc9wwilYYHESzVwb0t0MO5OhiYLvyWfF0xAxgXfcvvw
+TYPoGEYrv/TGQyRQGqvZ7jI2fSNKjo44NheynmyRQeSJCkQyebAXuIjAQOGMXdm
TFak+kDKtB1MwU/SjtPjOexi1Ic3l+oCEgNYbeBqYZHn7bxBGEj1NMkHK7mOXsaL
aKpkkehTFnk0jH9rAJATqt+XsG4ggHEwfQMG4ED6lHuapJd7StMqUZ9k1T9JF2cT
rKfcQmuzsZINYmxVW9nUOo4X+FAJa3H7wufO2O+VOlHm7K9hfJzwzEFbnve/kKP4
7QG250yuPPlz9GK3qejgWrotNzwU9CPd01M5fgghgpJlS7+JbADn4vBAV1+BOpyl
helDT/KPuDR5zpOdzBP2WcAp4uS7NRLD+34hgw77UHqwINhyZhTK85wXhcMo435L
SFtbD13DhYsWc9PGp37ePnlfY8YOUsCG1TAoHBYUT3wWjvBL8SdGMa5DrDKKWEcz
Wm4DB/KtUwrgc0wDzOrAGPwad4QHORJsYHkG4zs/xjYAe3I6tWyALKgsPUN2Lv1k
efohksTTSQ0FFDNWdzwCG+9KZpxXnP1GtQIYeh/hr2vci29VHzButyC+U0KqmJH/
gxgzw0nGLsGVk0hFDHCwuWdz8+zFlaM8pl9a/N8o3kj86x/e2tMoBsIFc6jepbAX
nxLG5bFzLk/ONQj3QbRDtsCqfc15QWlm4jdFtBdIfP1N1punKzUT4dMJTpXsXMm1
UYcSFpRry/mfAa1sytdbWInDy4FXtB8uSsW43zPvfZYCWuBjZF6SICUlhBeKZ4nX
t7f+c86rpHBB3Nm7fKmgr6WGwmCBAYqryOCL837AmHaXS02XRLiKIJ/I/KdqTKGF
FWBKCCFDKTodYERwWJ5FArkkcqysMwIJxlY5NMy79wB3dS3cb63dlrVwJ7U3rMsE
7BL6WP1ivRU6iK8ePiOLgqUohCcsiqKmniYEczkU4+AhK+L+CZmvTj0KVhnHt/2X
EpFTGt2FNstgwDatB5/JYLo3PtfdGsZDv4UbiGGO3uqkH5QbtmmZIcVJRXbG3YIy
db0e4DeosDMkYqHe07fE1/h/yzowaW+sru3iMPPybkMkA9IX4J/JVgDbTmxuadIp
oBhnwpVYmZk7CIVKkggu+WdAUGVBc+Dtv0ChSQaykP0C0z+Qk45k5D5WlrOF4S9q
hnv5TfwqKDadNNj5o28XccXjV9fVKoJSSPYaAdsawvd7ganR2kd7i0G2NfNZ3EWr
QY7Ke1zUJXbyDjmLEQYgIzLHqfCn/key+8lGe3265WHlSjZbB2foLPpbdoNxj9sa
4e3OnnX5Gyl1KrUI6+pr5JejkQqV6yLGtlBUx5L4wEQ1cCi63vZ7qtJ3f4HUGkm3
97NM0R/of8YTDQaceNOKnr07w4ohq55BOuzidU9Sg7qUsUBt8I62RhVSgCfg4VXc
MaFJLnhI9IPAp9i65oNXgQPgol2GkIkLNAfQzX5LGKr8PErLvTVH5BzdPLZEGaN0
bgFaV/nsAm8FS6daPyYc7fklombGJN4APT8ROZQr/aBFLt/MrZLV+6s9gD1HgQ1P
zfOTJTTeo03wUhfTSV2Ah1jmxpR7LZkItb8RVMJrgbFt64zGRSnOIvgm6Etkh+k/
uqRISwJ2d3T0UVtpUAii64ZBJ9M3eBcT3acPlzT6KPknCFSqYTPUuTig4iTlQNz2
n9ieCkm4ZYIOqklrNqHtJpBBtJxGgev2MmAMaDURRThdQHm19fLgu8WxF5a9egFq
m97st+4mX2USuvxJQHt4lrDnjQsBtm8arLup3hiqTl3pTM29BvNMH3V5g/Wr/Q6q
s0XvBWBsA1yoyF/2+NNMHLY1U1lebbLHNIUcHhqLvJz+D7DabMSdLgp4id20v3Ph
n/xfajX2ADQ1Kj+05d7wfWSEixc6tB0/o0IJTiviXSs2osNID+UNVWPZ2FpkJmfl
bXaUHdVj6Po6bsN/zE4MlfiJLOueoPig9lKQb1iqiW83vjGCO8Vtv99vkddA7BDp
hLxcEq7s0LiVDHZ05jecqu2QMNjIcpSy2fXhdmwCbKaFi+Z65WRGOl4JbORckVCl
PwV6dr0CYmFaATR4v4x6JeHynGi3kDGDtlJvIv2EpOoXiV6A649l7kbrRWSwDjzN
ybHjbhFo+padwLlObe68U/qQiqftSNZcG04t66SVBEKOIYFOvfsQm8pkl2R0WX78
6hLh+O+RJGSZwmPoKLOW1oIsLD8atA8pxe/f4mTP8VV7qF0hsme057tHMKNStp7e
gW4ZpDwccQeLlrPFrpQ0tDqYXyZs/2fUEO2uaA7NjqGQ1DjQ414WHvS34DLo5NK1
8sD5nDLoYRteVLORWsgzCBJe9dFemUhpU5aCRjQrzkhCLwlrdnX+CxHecQCR97pm
gl6GrxCxePGiTNLB+uE16mHCa1ewdoId60q988/9jw+Dr1gnn/QLQEk2nCc6PAbc
Qu9UZeWWeSOCTxa72ydH601Ns8LnIeUGO4uR8OB8YBe1S8joCevFKsLPUM0gQM+x
y9jnD0P+QpoiqsTYnEkU+mVCkiABCIS25I9/MQmv/GWRgA327eDvzqyd84sMolR0
p6yOXZnzVT9f3ffh9FIiJddVkhd9oa467klDlKxcp+J0/TRnoDgCplI/B7/zF+I6
LfA7jFsyAXUkvBS6038lc19E3/hRQ9AmWwevjPdqmwx2R2aIUs4ueDMy3+DLwpzh
aefdlb1xA1ku6J2+Xeo8GqBB68rz0thAPgups0UDr4XoqSri6/tN44zwajDuFeDX
6fYQvvoXqS0+IGvL6DN8u53JPGqlXfRZLfwiIEYMCL2z+OSxFVP/OjkxQuKbki32
2gB6MldACGYsRCVvppG8v4t4PQGQWTnVyXA7NqXduhseJNBu5mTSJL8qC50YoWkY
f6tLjM6+jveUobgDVhGrFYGdnlgRoqp0jeuryPZm9ZJjsSloWJCFXQPjBIJDcOG9
tQ3AMbG/b1eNJ8dVyH7SJJAXrWnTQegAjUQTxLMtaP0KFKb6oxHEZ+QvuiF04fDW
FO7HIwHnq/1wzw3eo3gTNH+G8FMkVotAbR7EnOPQB61bQFffj6O0QsGldCcCOnti
1ICwP7G4PtWgujARYZhh7r+t1JtNAsjFh/Lw9dsWytSjGy0Gz2iNVUNKmcIx8go1
x+I6sJiSTJ4OiHdTDTvChbMxsB+KSyJQmeUsNxY4nfLQhADVLdLegOV8+DtwGB4F
jYI7i0rHmuxf0TTsOrpf3pCRaABLr7aMZK2vm4ht//H9gv2vZZ4p9gQhmMNX/3Uk
vKv+5ji9d5nXkkHdXG6bN+o8HCcvZssPotFRa5eC+RXllhif7bFH2na2RFb+uNjR
3+GTSS90ThxK2u3wQaCpL0W06iKCF2dQMWmC/Qg03R7f9oBw7dH6jCyVcYCTiuHj
nSCFR5vSFtsqm/jWOcV2FxsYoTQHuLgEKS8LbMm78nTNwM6WCx8EKcyLbDxgD7uu
01yV47IihCu1uM4fFkKefyLE6zr+VCFlBv7fBXdwr1C1CyaTdeIpr+joODO1DyUY
X6xXXBWAVzups2Wqu+w/CjHoGnDkvvv7jHqYqx0pGrtUMLaIFFXlLy2dQJtZEJyU
RqyOGMw/Kdrd3DtOvq3KBnQc7dluZ/NEMV6dDdzlsZOt7GwOcC40K3RDI1rfXtfY
dmzV8UKjdFaefZebsnOspWVdE+gOVRHVyv6PafJBz3mQRmtmSarfKsuPzX80mVNm
set//Wu+s8EMSbZZ1glk7PajIH03AJcLX3hFVCV1ieXrCqfZy0SEz2yiGV2r4Jxy
UdvfcC2Resj7ib3ewq6GGWXXGwOFVclNwCq7sFSOL9Lnm5XZ21VaLdv7fUM5AGIs
PSB+k/Bal7GZVtT6RUbBv5k0e0r2xVuEtwFlC0oy5Qe1tIPb671GzVnj71laywj0
CLVGUXeH9G1W5V8w4rXFTMDnVv6GBayAS613cYQegZ7N8CNuxlvoSkRoXAt/wyiL
tcy2ViT6OqqbvB8KaVCn4Y5BSYx3fpoF1AW1sFqWZ2YTeUDlAmEOnaF3blWmiMGO
8zeOVhCw7rC/8jQegejfCIIzKcd7UtXL+/Xuy2LXqVPF+IUkevEVXRgT3BZOs7j5
isaJs7sF9sMq+/FgUo0EeYK0MCWUl7QMKtxl8uu/DBAiCI0oDt60GydsC1h2zOuN
VmPSsGxC7JlVYnkHwgr+3mqfXPT000QPo4myn74YWZ7GeXGPxF/utYL3nFEBg08g
n+XIv2H9Zk2EoP+fAPRgJzFMY/pCthLTqWnxVSJv6dA/eKKwm9ZlUzIqwY8IEx2m
PIiMyBRcVWLMMSv1vn0Wm/LYfIODPFFcCM3YDXJ8pNBZORbTsbMQ73KplZcgzX62
SCRvLHXRvhDNMMHC44T4b1oEwv8bDPh2RiXjKDJZkiQXiGmHA3jefkVugPgV4fYE
P+/xLJjPN64sj8bdUNbHRfEjyq1d3fvvFKHr9uiG/cQ1xJjmFjys2J70VHFhYlvc
4psjL95rHLA1/InCjm/C/D6hqrlk2iL4/Sa09YcoGIt8oel/7AIwToFJy7h7qTzz
TD/hbT7o3y8KHeGCJ9WjPQIryt32QjyAspKJM3IbSYabZRNJjoLRdSTI4yJ+T0EP
8ZiloaSkH9noi1QJh2PBAmHlbdHUUur3JlX/ryYHhTFCfo3t1CXSWPmbK6CAGfF9
48odIup90YNdkq/quT7klpI6eDFi7Wp7FDxxuYyw1E7hNEucqpqU0mtP7VZWl5iQ
tXMDt1LeBLhNYW5OwCXA0/oB2IWnWgLoeGheRNkadIlyHftPdxSLwqWwCslFt63f
9dC8Di0Bzg2ZWE463YnOnZIkHghBJCeC7c1uZ0ehGv1M/e3JUCRzdRW9tYjzxf6k
BJQeZHk+y6WleiOjgFwFqZ3a9TW9/dK0hzxGOf6LTDNd/xG8bsuVa0LjQHvt5Dc+
9JfaIPqLYX+G8v4uinx7IjmmUWkV+xuDYvqv3hjFy9Uzh8y6S+ZSAGXglGvEBol1
WqY9DRYUO7ZdQaQqdnD0GpcE57TNSMQPOLMamD8ltjwPCOCxlP+TjTtd8MJi4s8W
3ZIXParsInZml8lSDFpX8Ix1wyYZMsnq8/xBBpCrcWoiHjdGPhHoWzSvm/gf1RrJ
xVJ6nwdIVgFtk0C/y/FlN/PWl1iFbHJzfkIV711NM5A0dtmokk7YNdZkOPHDv66t
HbLOLt+OboKB1hGblD4Xhg5BwRjJoJzU3GN0vZjrxxG5JL95yVQKbIqhm1V5HvVs
LXADH7nP4WmwGVEgOb/C+bbh7SH1P/0fwOIK5RbKBWIAPiyTJ16bRYQfqddVmsoa
SojIVlKT3Y4OFnDKR/AvyUmnIzgGiK9y4vV9LJ9MW26JECHwnZhJ5uOQLLmP1Hs3
qjE+kTUJUT7api7Mc/gZ+26xec5A21WZjH5DT7n68Q/d6iV3D5CmGVCMeZ4kdk7b
kwoubPpxnN1lS9xZmIR2h67YZqhtwwYwFWsFZwwPlGo53tmIRsghzDijW9Ng/qyo
vCpYzolmXUEUoS1NQhF2Ybk52dXKe/DRSLRxJx/UFx3cyZzVFo4uetHW0bbuK4Vr
Wfj8yiyXrzD46TabAE/C9/QJ4BUH1nbdM5mEJNXYxvLLf+oFW3jPydp+7rTZXSvU
id8Ncgp8VVscIhxypOkltN0+IgWn3cFcIBnHhJgqYTufhBJuo1x+n5k2iswsjrYV
E/sVYu2mIiesP9tr9nCs2wW8rfEL/xxCahxlVY+AGXhUrjhJyhwhfakeQiie3VWA
5YeTvqZ81+kvHzc5ul4XxQh5o+AXhGnpwoKSbMkI+0iPzvcl1F0qA05+pHfk8UmG
KSxH1Ms/AVbHX42/4m52q13w7Ixfyp2xdqhfyMpomDYmZtC2ZTJZgqDMjKwdeMvb
y9GTdTnUdtzu3lg/GKpIy7PpsOVUyrnC82wept8Jn9sZ9QuBDCLW5nTZibE9hLrj
ijhldVoP7kROY5Mb14V13DHRt3iUoUl3wozpxffM1gal0N12PU3c0SAthHV9w9EW
tO7DOMQELg0FBUNOJMFYP+Q7X0/1fKpCwaeMmyPfyMkF1IMzv+DyYc2mWeuln4sv
h2EfLgoZSSTCaFufhQbmV2P4z5V7MijP9LuJyyBH1bGqzYJsj+ZJns8HPJOPzpa8
JBFidek4it2Lp/k3nNzq/tKV3CCUaGCBtWDSbXPAD+w+4X95e6+7oqAsjjpA4sYD
USiLchiX9JiJMOq6nev85AlLpwDchTC43dZHrJECRgBTe64E/eX6J1MAKUnPyZwA
y2UWJ17ywtSFRdlsB2K8E3OWn+V9hh2NkrQpMVa/L5JDCha74PDRJCTKSOqngTkS
CL54K5go1nWtCulZgAOYZjZPvdbyNOmZjtDCutywiF2niVmOp3vVtpT9zblE5Bx6
/+CCPnV8HqrO/NB2ZAUWMwD/DGFSzYJd+N39i49BHAEPD7sGoHJVQarTziXdJFJN
LoITYor63J+XYQEwTck7ULdVIEPOVrzeR/cOWyZVAIrFyOzi/uh9gqNe3uO8YsHk
R/rcTcjBQULWxxC9wimuoVijguISJRb4bgF84QtS36rW47PMjnTn2VmBpQRwhvU5
WbVgfwkhXP5PbGb+E98k8/ilmZKr8RL6KoXVRYzoYMpWYy19RNG6/Cv4s4bJOPYu
lILK0DfBqeQZ7umxB+N1DHFcZVkbvOgF6DqVSG9ZIu7u6yD37nbOfum3i+X2kwrH
h6hrVlJaNPE3CygPL/eDdsjphlkD2YjjlSQSJ1LJtxemeKjxQjspXMtjlZNn3Ql+
SiFCTN0A+Ier3b8yRtpRqaTyhZLTkrOvq89My9UXRT/WqovLk+ecUyKTRCaSVJmX
4SJC3esgiyHaivW5aOJtIUMj6kz9XeLhHxiwm9XVzLn9X9vjPZL/gyp+DX/rZRlq
zibuqqzG2ssUvcYfgbYKsnJMyY/77UIJPXoq8GOhKKCQo9y2st7a3mDLCEFZk/1a
CvT0h7zKKLRIwpHoIsUh2yqo8uW8mPCZNhmow9oJVNaavrUhJpRS0wfPgklkCwb4
RCFORRQM5E1QS3J5wi7LhlYWKw39YJArw/5JBvAaTilkQwSgq2rXfVA9e6R9l64B
t7LnJS6+rY8npy+NH+u819OzeMwuGwYg7cDZB95f4v2KEXe8ZZTV0b+KXtrvZ6M7
bM2mkAldqXrGLyVeoc2mqctbTFWZhdOWd/HJhCg8m3LwdhpJr6SIhFYWRVXP9wfK
RUGElRHSrd9v1pZ3pEKLhm/mtt7hxmMd5QXvlidmTVAbKv+eUqt7cMxhw/lZn/VS
JFASY96s9Kl9WnoPgbrXJZ3SAsdhr8vpXEoo2MmWDTKqX4RtqzPYMnEWB6luZtEC
cih1Uy6vC7T9OIfDLiFo8bX8a72JqnfYQkE+oGCeNAeFTQHVmL0HeuPKdZoaCH/u
hYai4qwrPPBIeJeaGHuf7tPo3x8w/KXa/NDrTixtCFLklWSmhGic2COLG1p/OBo+
nQ1YPEMiCPvg3en9h1fK0T1yT0WCbjxH8gSFACCMhlQrYA8ifF33yiafdxD838e1
KXibUKp+xu7IKRLI/DLoq8KPgUXBWx1HV0mX28+y4aGOkoi848aJiLSaifHbIRM3
koqNSTi1SX8U/M9J37FxolDvZ5U04tQ0SRu4bjNJOwgfyBeg6RMmmiTyDI7oMAKZ
jS1Ef6cR8Xcx6rzgX7Yn+FfuSUVH04QDg9K9cHpd2BiQGjvy47YwSRR2ZmG17+YI
HYqArsZHWfNdCxmLbsCcrGMKT93YSZ33Cs2OlCVUIMm/ENQ0uATC9CVTA8CoHLfV
4P1LZtcDEZnYOwbtoI/upXp4LpJbnQ2LakN6Hu60tpEAIMq8CLAl+W9hkdPIiHkJ
OjKPY8B5vFe5/FeNJJ3fFNSkcbl+ahDTzY+VqM3JEVcYfkLzJ/lYFzByv91KJl8K
McsFI55SlNAZsfhFRPqY53bPm/OkG3YgzD7ZwunkFjCWPQ44e1CXsIZUazxw1r4C
tUyOe/ErHbUGUeO9hA+5Gx2FsBRbasJ78jnv2ZYDXDcMwDerLQUnmslkiOrvudar
gTnMO0KjnnQ+bRjQeMLBK9LWbmVCAvQBQo+xO50hjxY+z3r/p9fL392SWk13PKDO
e2TJcQS0GbTKSlQ4juRLq/7mQl54s0HkOpEwA+aqYce0VbOMgEsdrvqdii3f3JY8
2vm7U7sUeaHrHi0on98j4HJe05Us1KH5/dbEiDKW2QYpI7dnUbm2CsbAdh0F98Kl
p11SdlbO+eotENNbZorpL701fo/VNTvcDFBDCmXAScHqNzP/FKAyveXy9gHakVTT
DlrSBVhn6Rv8zMG4YcaEWZTd13PI11M/cphwo1cwanbHhtJTud6IDBqtuBVk57Tn
lgsX22eBypg4WAGpin54CybRfCeoxbQ3RKu5doGB8qlY3duiGIhqzMwYwFSUeGDO
wGiHYh8AjH2er+6ZnKS6jwdwBJThhR8GL6gNHmMHxi6VV7T/3vw4xLUHaRFY7sNw
3VNglmQmzOL0twQagqNwecer6/AIo0NAFbyDcx011axP1ZmecKrYt3Z+OsjGR9iX
OFeFKJniKwrnvr8mIza3xB+McMojTubTK+gUO0IPqPYWLrrRUITZuGPU0RRAeF/h
2Uds76G262nr+1xGpiavyVShd3CnPf+Uocmi0EhFwG5ZhmvnY09fis7dT4QWuZ4B
+P9rGZJiDqXbXLD+V0E7W1VU9i6kEyP/7N/BwyiFgC2ScNV1nxNRxBf65ROUKNlC
Ywmyf9iT5/6pULGMugVBdLuVR03OEbPmGBHjiElXqXwIBm7RLx4zQKs1rGzRNcJ7
vMld0U4qLYDUCxjPPZkblva3g4A8+eUoFLopJrEWNWeSBtIdYJO7sRl9WwvPkSVA
D1JBQEQJ/t11aaTuoRVY19HRXBb8E+wpaAAVVlXYjnbKoZ2SGSJ4aczsNyCHRtFV
UERIGkxYq0ZliYD5K7TzotGwNUqPR7xUuj0aY0Ly14AMeeYwGKTtcxmT7F7S3/Rk
oQQfYOQgWfmnf01myPB1uE8XVStFHj41AUPg95V9bzrTdidlKekJDCFidVsgyJDq
4t83ZtTDGlwrbhox+fToiK6NNlXUExKAXZVDTzcdOQA5bGX4G0WXDJecprKFzANI
7NBtIQ+PNH2EFsjFpS4Cn7XiLiq8JlH/R7xaxXm+JSxkucNCXk0JGUfpJeubQ2Kk
8HAaVJAx5fmOBU8J5Ie0UNtXai1RDbSGSeTXYf2Tdzzp+UsXjpGrOIPMN3Uwba3g
TPKHVFUkcdl2UIq4LSdiG3PIZRaGTpx9EKGsSLeD+rigbl5BsDScfoBPfdnKCiCM
+xVaZIqDZvmPOvdRZA1R8RHO+bnZSbA0O3z+0izfyjhyMrqL8aXE2P19zg+/xKca
KUXkd+x212IUE3wBrNLU+9cgdDeB2a7MKj33DaGeyJKQCbjF6RpVBrYvwZN6Rhks
GYN++7y9a/eVV5EZ+dtsllM6VRbxfaJebxIsoANJ3abln01KrF55ruOUA/tCwGXA
94ExAlERUv1a3rgYNqjIXO/ntp3MCAS2UrNZAFCu9jh9j+heSSi+rLNWd3G5wPHk
USBHWNzX/tRBYlCa0gTUlyUETokLj/sQ60F5Sa3XISouv5L6pPzzMzWe3h4HnOhw
8n/H1zInmrAEAtJoFr8n72XS/UI2A1MvgSvblMpqTULFkYb0zXH/LkDU/fG2/JZH
zemVV9z14tcAYE4ySt4YgIPXrTG56bKldqtLX0kuVl26sYnFXRFXbLyB43paaWiF
qg+Go8DCGhR6k+V8s5iH4Y9pLLPoDQwexxkPWt9yzBYV5QBcFF3Wn+/SPFeghgvt
bV9Z5nw7hi3imIwd+Q53uoCrBlOR2W0cEmXAn92DHzc64MNjNYeQ9n71cHHoBP3w
/rYh+XMZnp7JSZe6Jf0V7OjsCG9vrgjOIAEXPH2P9oQSoLSpnT0IbkgGsnIx3shL
7BF99SrepOI5Q5JWCRK8LwBvOOaVQQ+sUjv91x3/hYo1ijAsyY4X1ab8GVo3uhHB
jNJC3AwJPelE+zu2Wx1GpEGIWhNcxqXFys/4giEXnKqrhPvouIqtQtaylDX/pKzd
T4+ohduzXA1/E3yh0tsY/EQx+pG+J3FSEVsB85MzKycZgwt12hEx6P/2H6EviTTU
w+WKjJF0f1Iib0Vo5Ugynn4D0qlTERdkOQmq74b9jlEE/ziN5LYae4Jn5cbrGofq
vTatddgJxDI6qXjhR4mmpOwAq16Fp2iFcZ0SFxy6lGmFKGZ0GuFulU3+3FEdE0R/
Ws7MUWWNBNWfntAYucpinLtp8XHDhLpl2ErFeb1dW32Yc7pgMM99H9gh/xuo2osL
IA2QHe0tTid43UqXKh2XEzTJ77ReNdhpYSJPzTl2MaLXds4Yq8jJLn5/Z3X2Bi0Z
lR4zXZ88AwEJyANpHEBO7bhWxN4PIJYQWCMjxdtgFrOMvCEDxGIX8goBn22aIWRv
wAZtjgT8i6ZAZ8wTmGaixEYCA9a6uYl6l3rmzzSdNj223sb6JjCtrH0fPp56dBqB
sJS8xrSDF2GwUmf3cQ6yfKIzOtFZaPktRp/YXJhjyfLbD1ciwTZOlqgXLSjimcMr
8wMIIKFqqDnXe+OdBr8LD0TW5v6khKzqlaubFd7D+qP4yh30Eiha5rScnVDJQRVS
g621d3SpXjOJYhpvjXH8Wqa4gz4LQgzFoinMniSlnU4rV8/PmnDCbqEIsnZI2ywV
w5EQhMuG1E8l6/rb+nTC1GyzPvmjftA9qLBOfHCPQGqvxE0kzdTpJKNc0OoYJbdy
iTDiS2N/HUW70arKdK04p2t4nu3lZcSDgQVo1TNt4KXOyChCKtQypww85qKyTDxo
1lDpA3bhE+rTKRY7ej9Q8/0p5AGct25juy7jixdkOQrHcTH0yLnN6PJntAsxk619
29Hudd+vsjLvWP7UGsPbNhTQOoYeRNHYWFLLJDyNaCKXSlupHo4NJosoEC/Zcoy7
NdDqdVwyPnmMA+6Dirn7ZccuIbGFHCcHxKKnuuDLuQdV5ndyl4egVFtdpHjm+KjQ
vblZMhJ6yLwqZRnJP/yX2NwpyT/0FBEWtizso+A6qFNW8SJQXuAbX4IiJOzpPavD
N2ePYNEO2G/mVJo2LF4LlzFZKtiKJ77AiKwO6e7ALLv5kSkjyab5ePg6siZXyL08
WLWWYLea4P2S1Y5y/Wafe9MD29YHYhl1Vc5qgidzH+5EadNoO2M1Sg3aWjgL8cBl
XEydi9oqJ0auH9HORBljUHQDO43IOK+2DHjzDTfZ4BNl06aUjl/ZAwA1yTFvJLq/
E28qsU55XojcVnHNMo2yeXBK/ELCVxg74is2XJDUyEivs2rYGe+C/EamjoLId7c1
+KX4B4/NdDWkklnVF0zIRmUSo1IQ9FIxV9HuZnvLtg3bA4WgfgBYCbqov1yjgLrH
ufZK85oPJ1D0dJsYqYYY07L+S0+WPmrNSmfbNwo0yDvpCWQS6IxqCGfiJ38/8UWx
gt5l/hnYkUJs+jHAHRGdpZyN0waunOh51sLam+kLpVzakQ1/Be8eS67JBxSWUF2r
0/OPAfk95Cah5c+PL3KTteB/Y52OcFO8Rp3sC4O8HmYSJOzNgF5OGE0/h9yO/QmY
d4t17GToMh0KfjqnfAqnd1tvT3ye+OrYh71kpNaWxHm1gPuejICvn3xH8Jn0KE2V
pMCDwzkIuzn+DA/OHBNENTJ54yO+PqUFoW6XNeid8iEktPjM2e3nFr3B/d5mwx/8
yJ0ngttbFtkmFLCuWz6XyFpoUYpNcrFjuNhK6Ap32FA/f9bTMBCOCtWSDi46/1iD
hVwOZdi7xwiPuzsIeTSs+gTKTDAA9aCZCjKv62BchxGPnWqJRv/0eYHnHUwiVXtx
DdZVxH2OYjQTosY2Ag7MqPfx2GywFuyqM9yTRmZTjjCOGsGOvKZvcl9S9vm5Q63/
mBXI3SzI+ZFzjn4+jnU8MbTTskBRSD+/8dwELJFLJGSUSOtuN6evOScXd3P2CJ92
3dYM6ksaTS9MTkXLcYeqtZ4hDLxMjfD0ksJDj8d30oEZU1rWdc5AabCLKPlh4D2f
NbQolNnc8yrwyY2Fe5VKqkRJ33nKE5stxox/dKo5gA7SqvOyRGuYuCtitjOjIJnL
UbXrSKK/tWD2NyrQ/w9NrvGSgGsIQFxRU5/H1xOrE70j+6mHc1Wh1oZFrHssUM8w
Bd4GWWvSpsZa1ZfUzxkZUxPHlMAkoWcwggJW7PMV+1MQWjbITXG933CRl2nNxY14
zwgclH/XgBBcrSP/qnoElEjOeMs9xWomK+6V6RE53pU/clyHSJEvslqppdLAaADD
mkCzZokvYMoO/L/gb35urWC3o32+gzU8/84vxeea/dY380tH1TYzwFk8RxbHwBaY
PVbFPybZsvVHsJnPu9UKktY86GC0cMDmLT06AfkW49vPYrRhOGJTn4KhRdz57hq+
0Yrk667dBmR3zM4/yQ++TuNk/45u71FvI6fV6SJxhpBUu4H6YZ8wnmwKTwhDG/IH
lviNddXR25dBoSEtxjBOlEV+/X27YrrnN4FXbyZTykrPx+uBZ8TeHr3OcuS8yUBH
LdJw++GqDzPaLOzCg2200p2VrPjmieBqwMgTQNm01BEMH5HZUXyOF7BZyIW9XBnD
rwxSUto8xe8/kS5HUaeWSURBiBXTV22TOPaKxsPxgFtsClmsL39SseraDvtpFmxS
rPGo9asSXLFYG46MA8BwynGa1UYEKIe1VI8oLZYRUAzLT12YYHMSeJr27vwSXcyh
gd7SvEheB2gYhNN45UnML3JoAtSn9cax5QK23QjJWaOBtLCBFnoqdpAmwJucLejk
C9L3hyDMRWup1w8g8wLmr8wQsvL3aLUiwhzOLmeUmJ2pAcucZHRpoWPk/jT9DYml
zdvOZeDWRdMaWp75/5rncOtGW6yYcllv2K3nuG+5YggD+HWvoWNPO0j04hiNaUbZ
FHUVrthG+98nu4tgZHZfymBX0NYFxkuIUHIa/7MCsq6JPxepf1saEfswQ9rnOC2i
aXXADbrPktScZFZC0v3u4+ZvS4+rNmoYchh6LL+9qjOutLkQumv7qCCvvz32Y156
tMDIKwWhmNkCcy4CiM75sRxdMKYa5OROeTHpmDGLNYmMgDvhYgj9drFj+PRfXz52
ujPOqP8GZpR7H6ycVL2RQ3s12nGcNi0OYXiMSeJj1YKG6UXyAzjIS5u8OtoY6M/9
TQAZLJhnfnUZ54A2ZO0T3T/FcJYsTuw3mFmWDSjEtToKOvw5kg+VfRVtMCgDv4VU
cTu31TeZk6xz10t9Pfk0tVp8fnhWpGbXbvvYrI2kJBPq8xqH3ZH6Kdc6dos+fuKI
ktLk3OBUqw40Y0ll4faIYnpKAnumLtsPNPbnojxBavMxsd+VLFB6BHJyAwim+XVg
ebzA4DNobvIKZXiDiNXKguuHRiMzBrLIaEI5s/xWCp7CWat52m9SyFD69FvK5Mke
jiAG6waOGAzS+1m242VFzVwpR8ZW+eWxejAVItDtS2FGgQgjcuLvmlpLRayE156P
ePhUT3XNq5sqVf4GgLwxwtqhHDA10fizj5Q3scUMcErHxpIcFqjdu7uPjkq1J9G8
Kyhn35iffmedGK5EL/VJsqttJnNoR2gvNSb+Vz9l+u4QS1r1Q6AelQoc750jG0dB
SS/q2N4cDENrU+ffKwWmProO1TrZU2fh8C100iFKiHdjLZHDXIhOqWeY5gKx8Y7G
sXvR5wyyly++gJhLnDEXtWnsAdjNaBO9QInBd2JDI8zLNP2SEDIjeD+BvV9ALgdc
WJGclRUMmxGkrCH+S1X7JnNHjCJdrrv3MwnuQsChzXz3YBdy/DUwkbwA0FGT4cfU
hOunpAU7jtpGk98l+0TyAFY6T6m0V/K9w2C+RxUdNYAIEFt6fOgbD2AFLLmpSafb
2TW/5szpn4O94h2Uh3deQoSp05ktdkzFY+b4AzwlsaI35hi5cCxo4kYS7/VVpUMF
PKx5umkCNLcJHNHc8kBy3Mv6bFIgyXV2jJ1YcqeXqvC6zdkoi+Jx5fJUfJFovQfd
0UaKUNGs7SmjVivFDKFPRUqqUT1KN7VAXou57q8A6JKahzNqhWbmgB8ZTVoQmaBf
TeEbSAux57XcO+g+e5LF9wWqOhzzj7Uz4nfJwsTGZDkC+AGPU7UJ39v9iWtEglK2
vIoREwj1q2KagMnsT/3Kx5n+0WAFpvc86yZZRSRBHFtGsaXQgQc0VGVdr034pugr
Y6QhrK7PLo2acIfOmV95FSFs70VR1mMZr0bainCMRYjKsJMzQ8E1aFyobKtYz0ob
JqgrfJZL1wr8MQFpebX0kOzjT1WjxlJZ2/t+jQQjR/BO+DWGWpSE2DRDCsVe80bw
rUkaq+GujC1GQkOcvmJ/5Sx/Is89IBxsusdrfNtVJQdVrlgLrDdwi8SCk0zqG1Ok
q6+FSaINJNnIKArmIeerw6lrjg+0KGtRvR7HK8Z57mCsddQGzQ/h9lofpKgT/Mmh
Sjh3IjOghVkDLR/HplZ1ELZiXoA+mVx6Ca1G6GMFfMAsRNuLmMGY1i3Xgmnb2NDZ
jhM2rk8ccPHTsdeY3E0fR6XOplhGycKPLN2juvZSWbxQMtvABHWRNXedqqpxct66
rpxC8F4VM6SEllo38GWePCnX88BZbhILghOlLU4I/kLGHUfnDPqJ6CmKoYRhfUdT
HKDHqNqh0tyy4noPZc1OQym4br4icun4bx4TnopFiOolhd+ylvFx4H+5TJcbSHMs
e2cnuV2tMRsyO1WeUPyqrlTcHD8kFcbgtJcL859ac1FXMl+HPZuMd6zI2hSzBTxT
/cCf3chd+1ZAD8rY6ETcB0UAWMuXVOG9NRPlI13Xoi89VDW7X8RYLpyQ4cXxopHl
RJRNfEetNgrGb+rUINFr1eikpnVCDftOEewr51O6PVdMarDYTthRm0qVx/xK/1Qo
RlRAH6+3MBELfZ57Gib8GO2PhBQQgqo/f614PG5RnnwJdeCB+v1DW4GQ1vdB8E9t
55LHNrjV1zI3kmvILLk7QGPeP0j87ui0lwnbZ3Cn+RTBy9MSBbvmffpaDyg6kGA7
zdeBRwBb8mtYDGoV1KHtszmCR5AohCH8HtLQdWMW12p8Y2U4O9NiJ3ZCv2C7nKzJ
tUWRGLlOqw9sgmxXAyeXD/qyKWJLJEranM1n+ePlMYjYftRbe95hdtShqJiEIdDB
14JtS7QYqb/OMrbILanLsWWRKDbD8sdmfeleueyW6qSUPETvsXZDi1Jjjd9iVFtH
DLZxv7UURwtjlnxefDCA90zpOmdm/NgDcwXOTOWnOWj1H3sQMDZwQwC9wC2o0WIY
K8wON2U1fARgjJZfdctcqX+o3eznO7fckHIpk57PsRWvg1L+LAR/BCSkgvVzUHZ+
+I+VoFaNgykGtNqNm7b7YtePBTvCukyL+JqHxc1d2Jw//I7m0vMRvNRtB/a9D/5Z
9tTQBXH1QeunPX7kHiyhjfZstqjebaBnUFdWYlL0LEuAlaCsS29xij4UvCIZC/GY
cbuXyEME3bSe/R+DpIpJ6/IPx4ypTNw8sQeDm+Tjq12/HU79Kc6ksATnNt3xLaVm
q+dz0eoE4nrki0E+CmyWZc+5ebH5rJVh57Qw5HuSmU8QUQb2SZXZXmnI6ztm/psp
+WCM3AygrelZteubIcvskh6+4kfJI9f7XljJOR4GPM5iRp2ods/y/c8XbCtd8sTn
OD7nxuIBYp0H/QKGjX5P4wOjhs/cXnWeHa5yH6XJmrZny1AX7wJLqyZwyL3Pc1fV
6gJnJIFho8NFhZB+HusWSLXOXjBelPaunHyfaFBLyt3oQB2AikOx7ZrNsFxL7mdM
9XhBMYsLZnmTHdfhfbwB6U70GaeSuBA+dWMfxuJdmTpy7iOIoNwJHG54YbjgXdHz
H/zwd0Y1kbGVVJDhDmIWhvce0wC7Wo6Z96kF5toYoi+sZzpYxIvqKoJca8LwDhi7
+WDYN/yw5IGciHK7rz1vB+BN4JZ9JFC5qG+Ipa9DNywG/WsakDdunPNpjE3hCJl9
lshpoC1JqIH3UQAaJNSYGGiyT0gApmlQGtpGF+nc+UGtgK7GCdOW8r2KOHgB/CYv
3ho06OHaNObtrOjpMq2hdCS8csS/w2hyQDUGjJ5w0lLRl7d2jeEKaaqrcoBKGPGs
SMg0TH0tLlfo7h/7Uf+zvjAfVh8jgxwUsKwd4/LzHHheRBoZI7AvHbAPJuDBwX/5
Fq4phskLJG/fDJ7EVGNn0Ff6MZ811SeGSolgkbUuQfRITAEMfUCpDI+noLhQl7Zp
eCUBwLIA1FdTZ+LOcjQbLF3MlAAfJS1VpwMZVj3pPIncuBeRtm2j0ImCwtUzzOEG
Dbmm69KEoe+qaqvY2wV56ZaWmAPfLDgifvQJ8PKTECqp1X4FFsQ0MNM2znvQ+Bul
b1pRlrUHPJqLe8SorIaW2ddetchTyUbVGSXhG8LUwCtXZnTS9V+R7Pvk3rOUTW8W
E9exj/CoyeITD6r9QDRjls88kwHCeLKNyEKZEB59w5pECWZ4OFrmZfISsnwPGI8b
spqMUwW2xMXMJpDDwBmTX2DJyxcq3653Ec/Nk/UZMZHyiUgJy760LVEsMCwsp9Vw
JBlZPXBAk6Ou5nEWsog1LdLY7RO0GjwGUeWGGW+QpVaoLPBYlPzU6frigBVW+0tP
yjPR/LKkJlKBkAK+EKur6t5iv48O8QiADkOuRCYP+TvJXIe43uosk5XvC5EeGmg7
zG2gMcT9SCuz/1+7i86rv8ujWidVt5A+dIroa0U9jqP5U0Ib/Msz4NO7eMbNlNoF
F2m8p1hwVjqmgwpstGACQbXiZXCBevt7F7vlR0tAiKGCfrVGSgySpHS39dmU5nbw
We0DOPdCQDJ4n740k9WHoJoJ5gd5XLxBsSQ4XBd1nl6a0w06x47ykShqItnXUSWu
1zafnrf/0ETPONPlWmjOfSQSAopQn7VBwym7UtYZ8OIDiQzxoGumsv+nj/ykJ2ox
FQC4ByDe4UwKKLBWHj6hfv14Bvan4lCqMr8ouNCKuFTEvlKEysCwQObEcFORKu8y
AmChwZaXgYVvMQQZ7ovGO9qSdjVdSLRtJAWUHVCshNpjF78a2W2qhk1X3h6ROKaY
e1QP7SN9WKR7ZyqKa7E1Jnk2He+/FMK5zlz9lB5IIWGHneFAG+pCnYHe9WWGQO6R
OwbEF/CtS+Jrm/1V7BFe5/SF4ZGgc6j+lYWDc1svGth6KsWDa/b3rUmH9F7xLyAR
zlLoOxP9UG6H8emg10wRRHucspeJ/kgtpFkDO0ogx+2jGGZmvLMprA9lMETEFbbe
ExAcqRW1bPmBkbZaDsGWjZmv/J61H5NFYNHmMOnsT+lPSXzGE4wRYs2UzXz5UsTb
DJeL2vyplpcsFhxg5U974tDlgeX25poNNqp1eecLTAIQAt+iJhvWthN5aU4wrhL7
djn5G5L6nLz5pwr9pt3xRpXJLqH7VGxiEwK3ovkCNhWEu1uuHwSUEITZJi/Mf9fj
1OMukT7OZxOBrIMrwzssgl+O8GCB4HqNSmMtgcnrRfTj0kRMEMha8LNEqlE7SzHW
+eAfAPjU1p9dCuhvEszYUXxbj/+ER46f9b5YXHkmRUHMZGBdVwwqLtqmi1Z0Vi61
nxKyTWeekFAUXA7YDLeMAzzQf325z3Q/+SKksNkfOWPeerRvnQiwPeu+51TNglfB
YHBHrPbFuOJH4CkbzeDEKcwYLYfWYwJxvxUp7WyPHlpaKbzirK9UlmGIIDlvYxOn
SpNSEb9Mp1STVioBY07Ebh9/YHaJfCrWIAk0nj90c8Im8AV4MbivKH5UHoOo31ku
/s+Mz5rGOBiVBO/KbdAL4PF59qTz3EnK4R+wrpnYxZuaDZiqQfoz4uDT/qvUiEdw
qDaBQwPmvJIx4+wuevEiSSHIeNqcNm/5CECjeYvt45StXL01S9H9Jc8AcE7WtJVy
fgqwHx17fQGI0TMUAjFBWjOyjtlsg6/WCi4l+QNdvRMsxFcylniuS9vESZ0E0IcH
ULlw6yCxRlxh52TIROLNngbuNjgQEQADxeY1yit9zHdg3HgjzLMP0Kt7fLVpPuFz
4LA6umN22AYyQaIMprimfKq8Pw210qtX4xup4LJKrbSubs9KhH6fZdZ16p2z0wkl
cm5CLK8kf4arcGFTZwkTFKPZylYRdy85AT4PFvHNZZbn5ZAiAJmPZ3HLpInS/4cr
veZCY0zDgwFJ//kFXiny+IDKIKFmTU4v3+Isn77WevY8pBdoH0EGUek3hVuHjugy
QkW4Qs2wYOA3PZEj0C01FpFwqxV2zxwGNdWflDbgu8M+mqcrk1Wh9AhSGBBX+zjJ
BwSFwL/gOz+/4WNH/Ff1bWq3brie0bkLO7lMfvbU5eFYqTl0kHg7bRUAc+xtyPaN
VVK24xy9D9UphgAgXx7y4O9Y5+AgmH3Rly+b1qva3AT4dfevNO03oxc9AkkQEILZ
iLN3F1qf+0gEWKa5ipH5mC9k1I5iPkzFr4gZ1Lt3nVW6aOklcjPLPpkqxiIwo84L
PxTjdjLKJx39ODQg/B8gZKrVAYPLg+IdPcfxNxciYONm6YrC1uiHyL+6Y15+drPB
IQHXZiKGMuzRuIpQcYQF24DAc9zAahloAJ42MiR3g8WzMsDy12NIu9PFK2T8+Aon
VlMCRuV08EsJkXxWhjxPbtRXwVYZMgTb0V5VQncKByJlOHIUCkd07RsFZFlKzQIM
eYZ9mBEN9mTBgGuSZm2r0SUFiBoRO50U1tLp83xU6XRenK7oj3LNspfO08coNnzf
U3I98O5Okr9bis2HW6LDAZDo/DcyQgnjpUrF39IS9atR48P8t2mApIp8ISbuHBd1
S5tSsAjWMOfZhDFc4QBdtx+xiL80aEtTMNlj1qy9IJTjrD7ZPs5J9pzSW58Eu4xl
+QaF5c4h7zEUMcOjeoUiJl1cyZx0w5DJqFrfHiuU1naHzKWpDs0inYSbZNyF0DfH
3Zgvarii710OhqoUIDxDk0S0qzJK+oR+JT5oXwZdAyhQAGhMU3K/SZt+JJvVwkXc
pxGFhFWnDNch2/elytYi5HMNDL4WVZXCU2r6Qulvw7GmBxApBABbNAahQiq0way2
0hiaZ9sFL1H34ZBrsdCMzVPx4996tIS/dq0WW0lpI6p6LQIIGW2+8QSYV1fayPd3
m4W+aHokwtaJDIcqZdtpXzaj7D+cENXF0IpTAtnaD2v6jmn5EZ47o6hgKEe+Tenf
rpo7lmwaPFptadJW2qLi9y3k06HyGNVAckZAJrQG29uGjJ5v4AmcCM7RLZ22+FC7
LuWxaC+SGdAdqoIqEU/oc8EdwBix5MQn2dwoFDgEpcqfPFQptIGs00HaJUt3kIvT
/oRSzIB7uEG2/9tpTOIKOfGKfH9jNrrLwdcgprHQjHtad0/cfjqzM1R3I2G1WA3r
drq8FLWid7b+/wE9yD32XzaOGrkcXMP/Mqotur7plyGGSvUxAJbWpy4mihyaDPHP
P2RW0mPdiNO5z0/4+b5rJdoRsCNkY4e9moBQD/c7cyZtFvDTfcQcl6IOpoZqTCwx
N0ALIQJVSvsieZXAIJbwFHmoJV/oB+1VjcMSkOuC3dZEN5av2lEpHwuN3bjuiG6V
CuGTXcm3q0bIkEg9/WzTugQFVqNbdKWLzisvYYmvM6o4ohkolkJEwMuCdqBy3hlS
KTa8LU2vcv+wx1B3RmLIvBrtNa+79U+mOIHp45dzbm4yHwomukkvsZVsH6YOVdiz
3T3uFKoZjk2nLyO+5qIzYjyMRHR48y62bIhsygTJ0hdFjhKCGSz6OUniLwTwd0XP
Dbg8xYJtxiDbSP7oBnlWkgS4nD6hxf1p+POo1P2qq/I3GZMRG2p5ttJi+r2Zb8SB
C50lzVflU9R5M+gSauMkRLwCraee6E/HsF7Et3Tt9SHYu9Niu5iQvkIHy3IZhoZR
tEQxLJzOjlenFyEfWSIgY4jlnUCTzEVnqWFofEVx3ZB4uS/dcp/WuaAZQVLOcPzI
pL6HwyIjVHLS0tUjxTkiNJL9YMcqUKUzWVyjYQy4nxmv+pj/DCZ0U8nlzxMdx7Vl
kZ/u3y9njXwaHRxLC0nYAh1nN66Ag29rIvRs6FN6GO8spYpYLfzuWv1v7wR3mIik
3jfgh1Bg7ZC2pJK/S3C2wCgB5soGwrqNQDR9EhtnLdvPRN43RE8Z17VNBErZgoT8
7H/pr9zJqUpIir7oFZ66T/ommXZ2rajORdclR+Ne4bKcnJmqeISKvWNDuAZwWfGn
w8qcXzCCd/8oDpLl/vnjaLYoX2oIG/HRPDFuUng7bdg/slTbqNeyMeaNGx1dgaDl
wbtnsmdZhFct3quZRJudTp1r1sl4tdy/pZiSJ50zsfjGpnyCK8l/r8Nn6u0HEC5X
kjLzr+6mpCI80laPMAMPD74r58tJoIMtC/RH9b1qZNA24WMDDGHfnLKV/th9cPGh
Vn7mWOz7VPTavXAQyGY4hvlxDRxDksWz9UcO3YTTEUOn4ANI8Sz4nz3txph0VHKd
WS9H/6HcO8oZ0DJUktEffn6Of6a5JbLH8mVP9lMzwbMXGVzp9mNkig/z+B9v3DuL
+A7ZodQcXuxd+76w2HYGM91Tpl2Jnizav4jJgCC8djSZsYkc+0iXcqw0AM3nqpel
mcEOtlPU+UppelW2A45TIXcoaGT0/hOLXsj1pa4qQW9/cymfjSfyijoL/bxa/zVx
GnqqtGbh61YEM89wx3bJyYgGnd1Z1ckkGd+kaGtSgznFzdIdVugVmmcRDljwiWkg
Ti/0c5tsagYPNWFVueg2T6mxBk07ytaxKRjg4/XDlpc/pNF+U0uVeNM+5YK8jpRs
IkZliouPSsbeElaiXLpMXJ3zE6tZVlplBmc4LAEfkIt4OXlQpwEec0J05app7mA/
5wARCKzrSz38ulKQ4tEix11aqbtDxdW7iesvHHJgvkU2H79jlYjqX55q77L4Ijb2
xTorUauLGKtd+fbWTCVIrlYt/ftl1pfhEfxgBIdJ7cdBqRnP6lsEEYqnbLLaHg2d
kMrmvusDq4vNTC+3IuZ0kV6W2dMdMTh4nchHwJYFoAjTUqV5XcNqJoPzW5ZapUq9
lT4OBnn7yFFT90XA8zZ7HnDPIbF7vv3uie+PPFumKBvPGbe2koKXdn5uOvvMcvTW
94uZvePyVxMizj1W0ae1REzdOS5XBtH42rMJVYu6qBXJHXjjI+BCXH13QsP7Bi/v
JYfiArI9tslBPG+5tmSnK+h+ASMEuOzEM6nVoSkpTISz0tWo/+OHiIouvG7f828B
6MJPtgQFkESXpuEqKEMz2I6Vt3eyGOqJ9ithv72LQuyxtPWmA3W5fuUI/kh91hKG
1rKRNVExjOGCtpEN3cLc6fX011aogEgCz3HtaS3zoJW1+l0VWWdUVv/cqrG/GHAP
Ne1sWtr2dkcYgVB8APIgIYpVA6yqnip3Z8cvwCvsfp/OEhrPirM7srQ0xlhsuVdd
ue/HpXwDIFQwKbZlKjs/zTbnYtmM1W+bBqIJuvhWKAR1iO9qb/thJzn3RpB4G1ir
xIeoNZAjFYQ/BGtOTCliudDu0b6mnLtpdpCjU+IsgDIAd7kKuq5ACBphWG08npFb
SsogFfmFShGvlaxuyEJiHCQZXABqRrhjmwsNnQ7tELTZKoC2JSoWHxIVgdrDVy2w
cBoaj2yrScnIOrvPACt7NmBMFPvHlEkMmE1wUck8jn/FO8oieTSH0NjPEDTtiKvu
qkRb2ZwqBdrtwhbrn+96h5JZHb5l0xQCFI/9a9oiHxCdBlSdWBtxn8cl5mcTXVyD
BRIG2thgIuMQz2FwZ8uxe2n/u/o0E5z+N5kotDVf+VPsMUgwsD0lcQgr5Qwa7EM4
94WWCQImM9GVJpnTvjnyBHMEbbpNvJYMtmbkYx6a/l2FT2esFKbG0q72gg069Q2q
XRNAdm0DKIbZqO703teFNyHpQeWEh4pL7s1afp+Aq0FaWSyxYuDbVeMM0xd+g9OR
DvIrcGcUEQXZQIPb7nsTvJNqCT49ZnCi9L+Sd3+bMwuXLeDDM2Qx/tLePb1e7I/P
5yG73hgHtbFfAv+Qda728lcGJf2Yteu/iePBxkE4Z1P8Y6lglF6r42CgTsUz8GmV
qbZONJPyJwxWOthTN7KN3DowjRbis4eIoYfSU1mRMIJTJRNwPiJsVpmfgWu+t9sZ
3e2M0M2cGpfZr1B5BIlGhe7M+WImZZnTMK1JBQlIaTGgcjY5xE4/B+kc/UB99lKJ
nm4X5yi8foAqr6b9Edv+tWnwU2AASlP2OeYR966pFKcvOv6ow2Tq/g659OLAfQUw
P7VO+Ty70zcWV33dt5mBNNH7/vZUiYmWykeiH318/IDYz2uI8+n/stR7R0p+Ey8Y
K/nSVvndDsMqXm2eZcS7djOaaV9PGteSiSLX0Ff0KiRmfHyq/SyFgO4iaW2DZl5z
VNJ9W90RJhM3z2KlTrzBoaFbqoGpMs8u7OyItZxgV/qEB6DuONfqH7y3o41zsBH1
lbJGs/7cW7IcAeEawnjEF2/KWjqCb1dydXfIcZ6UESv/TLy1x7x+tp84KTngR2Oz
+wRflvlvb5sNKejEGDNhPD/HSojKK9COi+77TATyLATpPgFcKBfE3qL5gFOMV7Q3
0rZ+GZocIcMyxApvmcLRprL50S10Yq/k+1SdSOyNZgpRHDi4hw/e6tw73WbLhFNW
YZAtJzIbmKGdNUk4yGQUASC9Az35gUyeDlhDsXC0js5YKbGCE2GJgARDckooXOHB
bDfkhBMnVZtSANYKslQ2MR8SZsJEkXcEMa30fSafnVBcdQzPBHV0vPMeVHrmUH/3
nvkwcEtUL3UJADTrWd1fHtSA0nLbxpisw3079Gz0EHRldeX+uKrlo5R8OspSLRH0
7pknngpZCxx5rVDLS7YG2gJqBfom3+mS8GTmtllcTDgu8bBZQu77QdEln1FUfP+q
HtDI00xtP6DvxwXeY3U79I50PV5lo3EbzeLjU4dhdJW6moiQORI/wtD9mhOvWEx4
UhnJ6oW8K/qxUk8IjEuFobiNX1GF+AU44j6DL8QoaIEeGz03UQtNVw8cyrgjnacM
YQMbnjlh3VoYC+QpmQ1TwFGp5TZeRmwl+X6epxSopqPm+TTlIv3GQOIUZrqvYtyv
Njow5lVzrSIEf1diO/j4InC7BV9f9LqqCZ/PGcDD31gDjsiP/xs+KmkSPy8zKyoD
YE6F2l2hAuUu/9XhaqmepC3dgJc2zS1T/OozOHPGkgV/rrmdfweyY+jNoKi20ZYC
JLGWhcnwMQvo+yzMA1y6Rp438OceaI5jwR7l+Ey8Gk7gjKCy3mF9QFX19K3nT0lZ
acuXxqxvBwNx6rWKYU7k2K7Lb19i2dANjCeYGrR6JkGJUzwoRKGRsKQsWKNrAtO8
+c9UEXhdxtLo1SOs09X3SsdtUF8mj9Ax4pcdKx0nfyzqq/g0FeaCRARovuQCuFGN
C03RO4dhRLqIu5fPF3HqGG6+xfXc7r5aUv5SolEkijb7tnmB0OBTfavp5yIZF3TO
PsrZHgqt3s+AIQ+qAVm+ph55MJruYlcNm3nmdJdvjxahqagbE7T3566LwV6GC316
+HI9ZkQiCO0Bg5ruQ325bJaTxmcmG/rTwREzgODuXkrmYoi8MrTEnKL+iNuxlMTN
8NqpS00tlhyjTEEqSRlX9CVsf5xxkCRKs5izbTYtMtH8lTRB5cXKOGhP/66jb4uy
c7IQGYCA1btVWrKLPjYhsML5+1q3w6nNeaZmouXY316O7MyOS0GpwsriBaJrbK48
OJ34I9LOQ2PeTjs717Ai1rUXKInKsQL81cGOb71qEFMLe60ZhjqVYBaHtf6rt524
q8qSK9DoiINftLwaSbNoxf1fhlFl0i3CMak9VrPirMEMHxFj7Nto049E0GGHJ3hb
OXQD/LpGG3jjXKCarIsJIT90AsFJMwfMx2OdXBsGO9EHPxEKTMGUDqntofYrk6Tm
V9w/YTNO/j8tPoYs9H61kFEDtIY9ls4XNS4o2ZSg1pItKfIsu8yt5/OCNvAduitU
EPdMx98vqcZxk+bXWs+ei78Dv7UBXcRFMUqjj1nBjsIRjVpwjRgyBcmw1ZlxfYPZ
JfOej7bcc6a2AEvBPbeam3qa+AGsBQEPDWcDgASWQ7d1p3IfGffv8D+fA/fnCY4U
261d1hww8zIMGiGJtAVHehNVfbylsB4/QHhZJmjDv4cnHkaQF4WFrKB6c9xkHVPf
DUIYms03O21mssiExPr9SHM3GuAb7xM/Kk2Z7tVIYeuG5UxxEYa9KjBGckF+7WmO
gvjvWJnUclyWabmketJPFJvBQB1R68b04fHNMbop9/9GH93VQ1HoN8QD1SfQnzj7
GY4mvpAKeJ7J41D6vxUWtlFzFgq6cREfQytSWHV9fhb5/01+b4QlG0slwD2zTNYF
GSnStMItiPI26GAhFEDxiRwmXOxJ+XCVtwpbryynblMs3EAFbJv2PW1H373IwmXH
R5EDaqIpYSp022Tm+ussr/WOZ0mA319gGfDuLQB/F1C30nEecSeM7C26bzrF5Fhc
yK+69CQ8xgJUf9yCInDeSPTRPdTPnxU2FQJT4g3YNm0nWqSYwv/yr4O8fHEoklfW
9si8mywPAINfVdUSaua79OVC1gDoA4OHhrrxcXYU8AsTszzNZ6c0rAcyidO+y9ZX
0QfvF4Sy+jD5pXu0hXffCvM0NFkr6EJdXKJ07wHr1NOQ8SmY9K7JjWkUkNqJ7wjb
aekL2TUOmftmIvF4YAICZW05C+VrbWvQc5pA5Qtn+0Rr0tBZ6siOz+uUp/vu+Q6J
cKP+MO63BQWOwFoRfHwbCym7OHNyKU6n/7nmeQ2E1POafoQpC2uWY7o2NJy9a0rX
DGQKPpMCqSXIexgIvexJQgZBDx9NQsTZwUEQlJrdob4GidGt58fRAI2TsVJsJyDM
Z1yQ1P6QPoWS0n8oUFS21SgfctyioFMvptpLYauWliG7t3qneDPZZzNSLVdc+sWJ
E71KtiD3LZLWrFcHAi9nizYjBoHU/0ZvXZPkVxFIxUHNnD3xalDcg2SwBN/ErnOQ
mMk1eS6JqjfRrPTQqbdPQFmkpRC7S46Vz7c1gBzmqzY/3GY7RArd3+JvQWzbgRXr
AGe0oy86fThkUDb4kOjQmkGX61DDZ1Z1QyUllDIYAcAwRyYiVVcsrA+1QLTFV9xz
seE5S01BLdvhqZNYdmciPnzWz4FPA3yHouq8TXBlcqADhE6aXaOgqzS1fx6lYvuE
Udc6O+zxD7sOjKCdCZ3jDV0k8/JfRcT6w/479WO0t3qD63okSWfG0/bVXd/NPrrG
0P8YSunpGjfnm/WguKVLTMPxC8DneyL2b6A+XqBUaoKcHVaT7lyAxol+g3FsIDBi
RvRzWn8jrCrnNKw+B3rIo4MV7q/BMJwotCUZ+lZ+GKHAWw0+CoYuTH2T9g+39XNJ
s0Ya7HDzLua6VekeeAd4yEEjEoRDGXRT6giXtB3N/hRkeE2LDLM1hERt9YaJ8ysQ
nAXerrJH6qXgLqz1vkppcHMlq481odbzKi0G2NBqRsk8VfkAV3dQ7gWHdeJKCcRB
6n8VIB+E10tIbzTnDxMHXrxpjW17CrxN9ONqISO7q36efXRDnRInUpgE6ilPz3E9
MzM4tp0ATQNZxyxbYxe38OGZ+v8u2IYUWsnYRMW2d/7t8GtI57OLG9lDkoxNoS7p
gV751Hh0TGzO7w46CbdrpX1VQiv1gZ7F1vpD3hBxCvRrydtbRit69mpjetixShzo
GFaTnPn+reGIm2aJHImFqQM2CBHc1kjU9qhTLa7ldRObaV371IDHEQjsRlK5iIHw
qo5LtraYJGLZHqUZiUbeyFmafWl5b0h2NgZ3E3eGVsp9QcIaJ43OVuO/U05/97b0
xi35jSVPUUO3mkH6BKEfzCVmi8cCvFkY0b3WAlkFouO2zP846kygPyuDxAWB0dQn
fm5VX/djTsIoXrvj7/ik9kTpK4A3sfHAbypYlgT5rAeXvZFHFOzCKBYCR4vEnfMe
T1FrtQqQ/8d2d0LQNAiS/93LQI7vTenM32u37kPuKtTt7JZKObKnOOsLqIZgsmye
gNOoXAe7FpSrUD64tcjCeXkbzqZjZayb/mSyZMGAlSyq5XV+0jpkT5xGfnLhJVOb
43OI8l9xU7EaIM5tkdKIxu+0uB482SMydKrkqBd/00JVPckfCHkhdwAnoelXRsVk
VKRRwAaCf1/W2x3zlgjRKk6ktClTJLBtaA9bCWaXLJ7HEHB4T42N7Lsk0gaL7Mqt
hH3QqaqQ6v8/047sHKvM1Nqu6REyN3QDiqokBOyTbwtsPfoHKt7IByPpaf7jOrX0
BUOAYvJczo5NKKhep41Llb2yIk60pjRtE3zRSl5HBQo1Xfj8xnBT7y/P5n1w0A2A
g0FCXOO8eiWUkXqqX0fEiaUIZZWQ+1z7UjbV1spC0ED6m+w4uj9dOiUgm1BM1adz
dQasENQ9mGLmU4Djkk8hKXDuA/lHRplTF6I4eq/kR1SA17Wo01rUvNVYd21ePp3S
9I/mWRp+2qhDzMPDVA0cPfBKvhgEw4BuVmyyMAhxsPi063gtu3ljux0ZmssuCkfo
oKjXjYrtwtKE+q1UqOfbF05JSa24I3G4pv/XU7/Al/SufUfvFfkls72bMr5ulyrg
yW/fzLnkmRJ1yl/HAiRFf+bf0Pomap65d+6cR+zgaIkaWVVFE1S85YtHW/XvZKgE
Yx39XMsufYNnATXdxW3oRL6lONLOA6gfVcZYrysmzKizBs7m1J5alz+llYoFaPiF
riNCKCi3/nhgVAhqKPBlyISdnzCuOy3F64Ny1kUOrKXQ+XMD4mWozzFSHG882zoV
TJDB5yi57PmkWrmV+Us0SkhUsX6OwizjmCH2ng1h5aVAtV8T6K2/eqB8BxJ8v45w
hVjin0tL63sj7bOdRJExpJvXIbyaeZWV7RX2+rFIZ9sVw+0eWn+SkpIo/wIw0Hx1
CL2HySjLpVf1q+h3V/hAl5l4cq63P/iTh4Mx7IWJE4hSf3Z+17agfOLD69vFLDdf
37KAXX0UHzqWYz/+iLNMYtem4VdlpGbKy2fzZ68TYMYmCA2mEKiLVS2U9HT86TnI
2MQEWJbGtZ032YdMY1xAVmD+Qz5l8wJuRTGCOxVhcfmuZsKRpjhhPe2V/u0wCsFZ
tqeJcdnDihBkRO6cZrp9/pRd3sBgm53I5rpkCB2BadTFYHn1bPzC4IDwh8fpkY9j
o6KkMjRXmEbjxLLiUo0EY7Fi+T3e6veOuYFLdeAFT2Sbi/bKrYcT67TBP3nlstIE
73En4WYTJ0V+izdV42kbOMADLy6nbad8ONRq6pN73saeqm2SgGjlMy6V1I5qkCCm
WxTdlw/nnIj9VUsWjNDUO8F6WlLe93YQsJxCoIL2B2iPIGu3V2MNUwpaxFwTUvj3
ZaKhLP5N4rayYOP2wCyWu3B2Vw8v2eIQdNU0sWS/tGHthDHpobOJFmIQtNZhctSw
P67X10ZUKHuUKggE2syQd8CgIMITvQsrQdk+Aeh/tBfgnAea0hNdfDchQoaRp+C8
dAKp8uygPDN+LnuSEAoxCmxSH8dtPe7r1Xbchm7r4hQpQN7uQAmaD81oeQEOh5wi
FuyxXr6IN6Fou+Qno5gqBnOdOoAtjEHm7Vj4/QMvKuNZYTG112BjiIlM7nf6Jkge
mU3tqwyWIdWReEIRwuYGk6qa2syEjUuei07shXZML6J4UXtya7t/KYUdWkceB75m
62Mos8FczWJYQD1Peisv7Y7SUGnmz69l0pjbJReSfoPNKPFAoAOSNcjGnyoPPrkD
hHVtM1dTv1W7K1py+yQ4HRhqiNFNX4z8r0/4TbPixtTeOdun0U0ROie6aohAt3nS
jNJXSvr8k4QG5r093cNrU8XcoF5TBvFvK9pQBdgtGfNXRGwGHiqHwOWVyoC9Mega
ypEaQCS1P6R62roMoV+n44eQWDUKPdkWaXKsuLZl47aMSzL8kq2yIZjkrbELq0Ll
qnnRLUFcET2LksERUm8Ds2JWElOXr171oUo4iD9ZEWTnSP9wFWa8IpOgRs47cCWQ
LMENxQkYYjsb6he4NweyjQg7O8IHSzeYhFGwzuJrvOGbXKsyFlFRHOzIIMsoiRcv
TlVjKsuylWRttJ+J5Y5re8RcRvtytdJdFnnBCel6ocuzcmyxGaRzlYv82GhavJK+
dA14RghFZEIQ7rPJ1d/fUgqOQpk43dYSBQ+gnwre5t55k6OGku2EO9LPTTI7gaW9
DnWzu9heexJclSkZdi1T+b15M41QDDhvDpwknpxsV4zMFYkmOAtek8JGkBJIL3kd
xqjncWYYXC2lTLrFTv/N4WbiyHJH+iytvxvo1p3w6jLRN+0miMw2IgWQFWle4AyS
vfTp93AisaREKmFrXQ/3YiVEzW1Dod7U7a8Ya//AmHelWvonHW4mz8aetGnf7SN7
PORl3ZobJS4sA887gff2BWWmsPqjPSC+dtDaDljPl58T9+elRK0Ycuoikch4ICR3
QuP/kHhqQlMPG5Ngfs/OaQJsG1Q/GuLfCWidoTVf9y5vFY0kwRRmc8vt5tbU4J7M
7CsPtHTd9ikuhWkGSTO09pNU1Q8ILR+PfrWx2/OdWPyyoXyENhK5a+f30a8Zyhhs
VtNMJ75vowg78lKV2fmdUJTZ78mUSAK9SpsftXV1IfwN4u2JKnJbcKYngy/4hgHU
259x/f4pZkCl4pOhswuNZqfP7hFgVektC7XDm7vToiUDZHXGsOfM0C0eTiN2FGMY
pO0k+Eq77vuhJZ7A9n6pNHuk89jhPYSAnRrqEYglihuDdZmSH8EeRmrZdES0gT+K
xzmttc5JEaqILZJDwIs9o6NHg0RfobZ/vBr/vFJ4q3l5Rl6Fcs4+PnB8Y2NU65oE
GlNMJkMd4H1lkPN4lvv5urFQ9JPTMPlG8HMRjgSRfjKdLU9saPGisPKw5t6azwLQ
v17OxT1dr0cSNVgAzGp7gER9UO/8fCArEQb6FBMOB/5mFC1m+U2JmGZh71Hme60/
pF4dSqutrWBce7CZMA3kFcYhsbLJWlEdBtchoRcgiOOIG8VwRFW7V+dwzVkBsVQ4
qF4u4fb+9795941NCakak6joEsQZPXBtxD/mtldDucMdBBIz7QNNCOtxnt5Cf44t
Yibwv3oOIxfWBTpTiqUMfiNDT3FjW/jtgze4RGnhQnhixkEgpLHhT6DKnTvUnTUX
WdjWWzdfklpHvBMa0KkPHaxmK2QAm5elzM9ls82mACn/wZr1SuLivwNVKRoclahK
J4Y7/XJhjVevzG+Dv5ZgM0ku9r1gkegAk9hG17cF8SwvB5z9tDx/jm2e/PAqCv4V
TScnHwU59oVd/Fa/0czdvybF1mtw6s6Iacgg9feiZGc6Z8KMjD6mEqdnAByb/HAh
tnGZHJHJoJoM190AxC98JXjFY6tuhprkWQI6cr81lkBXD9O1ZDndahL4p8UvK6d8
czeQ5qD+jxJ5+Oo4eRMGJZPkfIUnOsieEze0iBkBTBhqPAYMyBNh1b9lma3KmArP
366OvcFjwS5CGXphoQAbxveLjl8YpZOsYf/fP3RQ2p+rJLTRpncI5+Cg+dk6FyFN
QwJtWP8qenylrvwb2CR2qaz6KgLk7ma4ghOWddce3EpwsPE4FjRuPm4wDjnaEdQT
CBnIce4U9K4fy7/JqBvcwVD7JtviNw/fPytYbw9Z2mXQomN8OQrGQFV019gSRmWV
cK4dWjVLpRYhGo2r0qoBVxf24cq/2kVlRzOvh8X7AXTUoAR1e2DrZydV3Vw3m1q8
C1Ov4cr6mXF/ktiO1hf7F1Q3U1Ohx9k51x5r3hHEKPW3cSqsE54y0iAjSJEZiaXr
Zd48WCo0DIEr/lVYj+lw8oLdk4FyeY6LlWzusUenvesjxZ9dqbcOxe6myKo+KwCV
ExqYoClwuDzZ+8Rn0918OzEQ1Z2VWAjc/1gYx0bKO9SPtD3XEKzrtv0UI0wWmpmb
MgTEMSSkc5Eu8nWCAxLcSVuNE4WLwh7oNFLcn8Tpc4k8IT0FN1oDDrj/VwTwwmqE
2L9CPx+QO5rW2D6FdUW2atxquwRwL/XN2UaX4I2sHBiFtNBz7CDiehejL56cesGm
Ls4lTuGC4QNgV9OVCC8rLn6wQLTk+qKHE7hVinJhIubbkZZ4KCNMa/XENYw0lIjq
RFbobPcXWnVkHpc7L0GIbqoxBh4+rR7HpcTjmKLXKCPCBtA2YgVFEXoTgo1HH1uS
MKbnM/9yR7dXyPdmta+qVcgOUe9T616OUUldCwqyg8Wkdj1xxwe+at5tSr9aoV64
CNTEwpE+i8boJIntZ1Uo9pSnooXSg7QY60TKg96TDU5DUly1ZnTzp2LZ0Edek5hA
/uarHeO00vbqp1Om6mAQJOOsxBno9yeo736C+PrgjTaSnbB25lMiGz3CSnxNhTyc
/GPl9SDuvbDUjkmNUr5PDC2j4gQI6nEyoU3Hy3+sPYD1i4QhUZClR644O9vD89mX
GwcWtbDdcB+o80pyNqzQfzz+gCzz7eXnT/3AE4jRuE4K1Z5GvwMwYjBEOwi56q2k
QvB6DHhkrqRfghj1qY16AjHoLuVE3r/xRwbgBg7WQBIRTySVnKG+mBS0EINrOpc2
OaCVtyL8c4ZfMZy87AiOmMPIPYHQ/dU0E8Ip+2m/RDxwU4ByeVzZkkc+Ci1qSZ1S
aXeLhrwSeEnKEgeKXocv7ZZy68ZbHOspoSWlvJyz7RKI8k4OcaGkuLnq7zIG19Yf
jgogPavUB3oi65rpLGO+vZOh+WEc26Qs0HkITLWJ1lf79KWPRvnh7qVoio4rm4Sm
9zXSa16jsiFKprbBl84oHpwVLFBU9XiqFcQOLgNxXYUYX30/BAiHNwPauLj3/j1w
kHInzu/yNKUuzzHWFF4ue0mgTCi41thTpm4FHpZGJ1PmNBQuiwQMp2WabOlfTf0n
Oj00LnkuCF3x2WMijMvY1hEQtELWg0TDtj9r5rKQWpL4cWE9XX0cFtOi3cK+3Tcc
KVporRY4txfbtAyxhf5iJv2R+FKMfdEMolJi77SkvNJiXuHx/e206wlcaLU2TjU8
E6HwDz4H3j5FL1RFSuSaODwPfYFDrTHi3kZm9ByaUIujDLU7NDV6bdYUtW6aGd5c
OTp8cAIW1LW+JlYNqh9eorXatquQWyqwEqE8B17FZBC83DlN/bU8rFVGH6Obrwez
xG5IRiQe7QBZBfTc/zDQSzqDM1p/4Q2qDSvdhEwzT0Ss2bdOkwKzjXhb5bIXcD11
zd6hUzEez3Exy3mt5B43gIAPXtCNDTiKVpUddUmrncQGSCP7IxkePbT5yTLrAnWm
eP5eFuA1NsKAcTfzbGlVSH6RbodtMtg6et1yxVrPAFPLL2v2FvKrncndmMs0qyjW
f30dxN1BEw+tXfr3nljvPlUGbKXb68Ny0e2N3COAyQd4j1B/lTrK7vILpi/4HhER
Phct5Ss4YDTCqZfRH14Scu24PNSK8eSrm4/+LBMn1AkIcyKlhWrhs1lkc/31GUJn
oClidtpGfSdQvG6ljsirZZoQ9vxo7kTo/fzlXgWqqqHAQJHLOi4Bs/9H/CUCKTUr
Up0xjRyuU7AyELNSMkRStQLLIZ5FMDcZjMyJGpyjinJBqjpvJSVz+Pn7BgUGkgcY
iinlzsKIqWhcX4zDMugZrbCVS5q/f0RI3F3psUMm7izqObb/qWy4OAxK5eYYFENJ
ROPSVQcyLFg8h6kD5svjs01iaocjehi6HlbDlY58BRTRz5aL3bUgpsK6+jLj4m/8
9Uisod3Gn2Lgns1oog050u6cXBzkx9Biv0CGJLUynQhshVu78l4H3PC/DU53TtTA
u0//TnM3QGMFx/3JB6CbJCZNYzYhNlahQD08otD7TD71c/WY8ALheXjqW2IWp1Kt
sX0VoYjtJl5Blr/q6r9UgytliClNci+WPstynA2nn1dppSAmN09wRUPqfRqMCUfL
pybLbLEYw+hDJ7JMjfL3WfT7uq54UACZWTVAhRn+82ZHl9I3YdNd1+FMOSnH2Cos
eTruu0z8sEdpDzezj5m8bD8QaOjPpDUMGoEEWFbPNMb1F/JhPQS9JYCOQReVPmZy
eGMact0btYSxUjoiVUnRxVqgYwDblBIQB7rV9jcsWxymlQNoXqAEcHS/WrFxcQR6
Q72phh1xJ4vgNckueILQFMyap/+jGEs+UIFymXF0gwWBa4RpdgMMJKWWB8OQJ5Py
SiF1HI43X8L4vRLNZPSPJcRW+KWKp3+HeXZnvmSGBzoXwmWsBpMkG72WTXj9UP4Q
UN/Hq1AQhrs6PDoKZD5yRcD9Fz6UsW4DZOOemxWSsoPFf79ikoYEkgB56A0ixyY1
gcCXmDp3ed7SsVRzLx+1NSQTNMQvlAKYadq0qaJju4r92BSBFCe34hWyyckNyhQx
xEbW0S28tPCvtrOYuRZG4tTVUpG9N5xfxZofSQvU8Qy1suKNvm5vpsYuJrHOGlTk
Yjt6KkRP1WKFcVYH6xPEq0BWdQqgdX27H3qzutECB3DgVO49Jc+uh56lJ2tqFPjj
wxamVxdS0h5us1ec01O68i/naXzO6DZr6evAJ/4LTg0TmEtMuzTv4lZNrPCyASUG
F0nn2OqqL7fvWP0WOpLVp6HFq8ZB5+ir6XwYRiLCOx91fin89yMtOFTTVPyEIP15
ssFH1o91+AwAdRgc2HPblRq4nZa7MPqG0QkB/C1njGxQu/q2bPHNtEKB4Ju4xfNB
8p29RISHhifX2VvqsbQaeeE+uHXtOk8onkV+apkacm6A+7g+z4LGCH4QiKfkjezo
gRkWoJO3U9Nl3saOXPOMQpwNANV9uMT/I/PvcmG3RjupyKqHlZNynWtlNB+Del5C
SaLlRu2MnAilUCHEouKoVohwXv0j9t/qxPXezrPRTcd0vqjnBE0T/do8RBR6S6cu
O2x68C+tWw/Fcw01b/UEu0PXzi2eFmA8ozpkZTW6uU5kIyh78anbvdG3P3YWAy2r
xl81x6RHZe7kYFl+YP+kNb4T35U8Aj1SYlp92JyPMqebDAH+vLxGpcBBwb1b7kD2
d+KMjcXkC3pZTFB1bHKBSPQmBkVJW5C0/w1lWZ2d0fNat8FN9RQFkD6ivz9vDc5A
yox8VEToWg77wCbbenGc9Baodq2jDGkEqonUJsrKDZgCgjlGU+a7bCI+tiJ5DfSK
VuK0tqlps/IJitFTfpQbknic369uhK1CeM1yiMDP0vk74+syUAyEewHSdLkjqykt
ANyfvA1If31BkgQu7OCyGz6Ct99+P+OcIIwboy6UH8f6tGueH/Sb5HPiUVSAsZfN
rdIKXU7+H10Fio+hMi8pvEDcO5MzCV7gakHgyqOlovCc8u2XQH2OTTnKWA3+U/UL
TGBiYbczdFE7rjDUUp2pTqyrXqk9k6iPHHgK/iI28KBc8UtfrhXU3HzSqr0zJMl8
yDDAw2N9LoIoAWYlKPRqjoW/zucL6Hg1Iy8cvxvVcO5R5oLuaDqBLX9QV2pqOBBK
HFJ//kvpH3WcxiNf31rXvCV/6m4ksVxMr0/WDlZd/YE7j5aOTuIwUfYnVVfCenLX
lABFJSB4poBPGOrA4hoddCXORlorj0SKf0C6yyp40304Zgx73Qm+eR3vFRYvoDOW
TH5FlrP8JNW23LTWzG9DfE08f1ztka+TF+hSrK8pwV8Ben+F+UbUHu2r2pdNZ/xc
lJvNwH5Z2NknAdwO03Udt2MNJFIAZU959KjGNALEjB6u/HjCjx6D5jvfs32gM2Ma
6UEK5SYdKgEoouaiN3vXWCI7fSwfg7FRfNg4x2bHECTKaimfLGJ4NzM399vCagV1
EgOvpClmZa+ARaUhQt6ckl2YSrTUFV5084WBJj4cy1Jw0HEKreF1u2WONg0WZteL
jp9XeCc3NtUhmbZpCNNNevKy/R5o49AVM0EvgLPa0EYpkqW83YPb/lys2lDRdwDV
64Gea960bzxzp8tOu6AiSqrs49mTyZddkzCDHE2dw48826OVEWMs4++3MQWERWow
wCaSD3SzVnMSk1w7QdCU77iXdaX0vacWhX3Wga8DpsxpqFzNoozWZ2YZaTNmnZ2O
CV/DwCMYGFrnJ9SEhRkx1YIkFUPT2GtqQzBoOwqRga6JZ2ESYShkyFMcAk0nh+Rk
jlrg3Dpt9RxJ+c/YkSxgn1W7mwSmaB4/JgRQaCCJTYEZVzR1+Iji7axW63u5Y695
EfrVPWuuFsdQvQ4Vciz7HDVCMAZFvTNAomzC+24vVsxx0R/SRodKbZEEVLjQEhAy
1awCCjnTRn+EL+tiQfExKqFfPQhsJk56pMM60/+mR8VHCQQXF38WbbmrWTVxwgvy
ucBQLIW+wQ4uYvlqUvH1n7rTv48efUPhSOM74Up2vDX4qxfGpL93FUoG1+5Zu2rS
VgipKiHyeZbXox363IjsF+TXVKYkTNFYRxEt5At2ZGKwROU/L2dMILLzZLtcBRhe
b6Y8Op/tNdc4M0P+Usv5o39KcOAWjodifJbdMEIDVC0jmR0ata4hjLKHdPa0Xps5
+t48b/NmbJ0YSTBbYQKwVQr5zoXiIG1LOP2sdsaMzlI7vhw0LXZOEuMUbRB+fJap
ceX7NNyW3ztysyY4d5uPpFdx2DnVtjGGoJUSYeDetuoV82u0V6XXe88ek9V506/v
gPqPLGeEsIYXKynKgF2mfRGtSxUfaUvlHj7ysTsXwcQknbJ5RFXqlB5YqGybr5E0
qGaJiQtbVMKbVPDsa/yvAXZw5701rb4IK55IyYldzsBwJs3jCMYMjyw99SukXOU4
MkOkMyu+jZxDLi1jHWXJnkAbh6+kho42UZLPXzVkeDJ0qlt/FyxYSq6QQ6V0OeyD
vUi3l7omaJ4+ctRfKWcXKSrUYjYKXNRwc36/U23aYR+1yVyW6ITzTC++NxrCuS+g
s5+dYYsSTm8Cz5dVesepiJWiIdgib82M0HmohcQdpWJnTMP06g7Ne5pyjAXBbrxH
obTZmpMDMRhp7yRQ78U96C8aHFTQDVihu82+/1Ko8xgCawLKp1t/o4t/+BGSgbS9
dFeddwZ2VPMxSXRATLdQ7CobFpT3Yqqqx9V+lyw6pktarzyNvBCkC0JB9YHywSP7
h8Int1mK+SII6ZEPjGfmhkskZ3YpMFqGQyds6m27mOXJrdchFpxEh6dhpgEtQZTL
2Tk7KpcVTQTdeZRbDv14vedF6knDhDZHjT5OkdPW9bhz90wsZ76HktVCP7uQgpU4
gbLL7LdRYTkaXzPi1rQSCjS1POmBTLleJXkVug4nq7Wt7AqP7AUuXonPEgp0W6Jy
Ul9lz9fCt2Upo53eaE4fhy48M+YRiVINtJEsV9l0CbuUmRTmnRxMbE3ptvK6I7IP
zt28fhMiAeMY4SgxJFk8tJMhJRYcfygt80KRgeELs1yYv7gOy3yBEGElpAHqN4NC
8WR9y4RW5fY/4vCA/M7O/8hHs4ppHgG1/hkhSe+GRC2lRv4XEn8H3yuMqPAY2oPZ
EoMKis81cIm2EnE4pudaL1zttc+Bq8YT+TMKMy8/INOckQNRIiO3KWl4zGBk9Gd3
v09zpcLIwD5joUdm/j4kbOHvWA0TUd2XDz99U+FXxvgHXGtH75zTZJ4B0PBZVRQ/
oQfS+jBKrFcqaS/Nwc3Xkhi3dQ06tqVtYLTss1vZhlKQ+aG1XS0muIu0P4RaqSVJ
VvH+z6+4uZdi54rr+gj0eb2AxAupGYRtEkXUfh1DwMT/YGP0wwg28xuHPlAZ0tEn
rgyig7zx9IJXAD6n3Idd9JPwQxbvUl/rXKvOP6RSSEO0tSl6JeZmYiPBkMTPm1Gf
Ql+ViLuF7VmY8+OjD4/TPfcGx02/G+xVehSUWC/bI7kcsqgPj8kiT4hhqj+aQixI
/I+2N1eS3CSziz9fjwJQyGth5wICKUi7YqnGWNDgBVYQeEkqmGa29IwzTIpJwcrn
WHcys1l7Sm7TB3dhDUQAUBBA6fyhB8+RZWZqVPJXwKdhkAnC6qYyaIn9zavYc2Te
95u/1TY6BB1PmiHO4kcNK2ydCkqjCc1Sg3EcXctg/gfO7uZR52O50WilZgOKt5MA
bo0hvSwTfy66VM07tHbLBwN8tJxOe8kIv4v2iWFndDuDFvej+pVcmvOmpdksrnTi
LrUu1nPMKj0dx0/bg/zt4aYgZivScghUizcPIF36jy54ysRGKpgAzfx/FNioswZG
mr97CVrLvUfbwBdpgfK02TuW7v57k6VGRgcfqWqwStIL5OcRCrAw5lCNEGNQkxCC
uNt9wDOaJRo6OJu/SZOZ5vJoS1B5LXQUJ4nAa58Mb8Fu9HjfhSEaToqKPfEKdgz5
qqvzc2OLwAUnRNC43HJd8USxC16NTaM0iihA2dwkAGk7R58dCjAf4rLurBL9ZfSV
AVlT9MAg/pK9NvyWmF7v7oJ5VVXixjrbw2SfawOoiZt0kjoD2KCLVVEeeWagr6nb
O50FjuPUeUksrOK7RfwCa/Cs0SG41JomsuNT5QSutSrYlOopBFTVOE8/5JuZ9TkE
aRWQeaPSV/hz5XL1JeQmRV+Ojo4JOz+XjXYVGTSHzOAJh+j6XTF209Q2ePwaQBgy
CQ03EejgoO/2sCxFxr4U9r+YLbunzx/lzsXolnQzV4Z0GjNzR8dH41zgoz0arvG5
ifE9+pTF8qpS5OLRWJLna5cH6SlpAxiGCwCROueOANLDhMqqhZ1J4KuVvBYUF5B0
hSW56PQ79+VDCrRv2XvEuc1gJWIOqPwu9VSmWHPg+a4dP+cq5nKlprrjYuprmuO5
qcuWf29/LJoCBcu8L8MyaF1wj+DtWZWHRx0mwI50GWMigEUEztZ/4BZyzb9mmIU0
BBKyH+bsuVvVAEdEJOx1OrIlsmsoqXcGQjnyQWc0VH3gKJ95tgnBcm0j+V4IRLSJ
sGXgJ1TNoqBzKSnllVO8UDL2XNotgWJkMDxbmv1jrCyIwoutfJr7WwxMMseoAOaD
UzqHSd5HyzwbUHtXqoIR4GqEWd3zi+FmeKfbzddMmGjF/y34T06j6xEsEurDYfOC
EfgMVB2Qmxujt4nKKl8RtrFCToDhY+gb487FcSkJvQAqLGqNOJfvvWIkQlpV7lkW
8bv5I9PkzqSzCsXQ0FsBnXn/qCENzc85nbpVhoezO9IJNETJZJMtENqJd3lV/Gp9
GIq5u+bFK0qbERUAC+KLGGZi437+RCdB5/kdDM4PaqxqrGDrZrAYSgwEW1F3qsgp
g+30VyEuXsi0+DfA1oVUXQWw+arIGaRyPrac+qeBHjAipnsggA7XHsIriZnH5EIe
TJeJPrunp0HfTwLQb0OrN3uM2BALavBKYAEGa08epHGZyHMwX/uSYE4dmUM0srF9
5QbzxqIonxSgBMY4D2z6GT2fRsL35R9psDcOxI4KsTgx1StpFs6TmYyC7fEOxx+O
dyYAuV9r8+n08Ye2uVTkwKx5eAbsFYRu0QvCb1hL5jLPbxdfCwYZJrR1OaKKPde4
6nq3wv+081DTgznfwuNFOYDeioSDZaFR7jIQ6T4eysKjE3EX6x2ZHZ1Q4b9nEQy0
Szxd2bI3wn5BuhSB/Q+Wj/zg8qu8f0zXPaU8b+zDUkEn6qCYo0Zovwws7DEc8zUb
hb2unQkJMfW1sou2WbcgfPYcl2t8ISlBFqNGH0WXXmpeP8GzB2/kkZvg5+VgLOe/
Y604TohbxoRR35FBXK+XgubDb0A9bmcu2f9Irz0H3PLdXVu4+/Yt8VffcZ4o4rWU
3tbZrPFJ83zvSAgUtVMLlCq0rhI/9zUmGZZWitC28big9AFDgqR7jWHV0cw2xn1T
XPBN5SCvxQ1k86nGWDz4j+ujTXAC501kPgEFsw2vhd5HQVAuqwnUn6kCl42rbXy/
QkIEZ0BAzPGdmW0u8f8Mujp31Qyf3RWuVUPXVnlAC7OvyWu7XjlhxT8rqEgukRRy
SgFh6jE6jAsduwtODf+FRn3TLoqHlklqpB6EtrjAd5WtuUyij73HwZiAb8Giue18
aWl2gqYdC8IYWmoe0KJiKSz9NYj84j6OAf9/928jVHs7viz1MgrTkWpaNC3h03Ba
F4ub7a1YSoJDRcVeDBR2ZEoFcTXVhg0xNs5FJGonaChFF1eqKTggfui87b0GRqhK
auwIOnUgEu/hsrZZ7WLVahRwTm7FuMv7kJGRfMQjTqRvSWQOW/qkSpU9RfwWR0NG
yfELz9Jplu5e++7XHl4uzeeqE3eqfVQDZHKF8P+H5D3eWSKkZkZAMQkS0GXnGp1L
C+cxQvDODwGo3OiYvkVZuQl41c/HzSNhuUR4Tz1zzeNuBh/KcU/d4sC99DKoPzoA
SXp1854muIEdDe7tGrrwBCEySrI3P3ME/osW3RE764A2GHfgapcZZkWNUnHh4TtZ
RS/4lE0e1kZpQPqU1j7QaZ2nOR6y2BwHEJeW4AAB4Mrw2QeH5fVDf5s7/jdHd7lh
ySJLQ8MmS8ib//GzP8feue5hBEJzO03U5u//rRGDxSWr9moNz6G4L7WqWdq9NHsU
kHckJB8gjI3tMQeTXuRGTj6EGWOzbTzx6wyumTP6VHglGoYxl5Ktfvsp44QbGIKl
gPRGeepNz8nMOVQcw+AB69da4NlusLXgElfvSU6770nsJvX73jnnKqsK9T4mfZcm
rXctVD7FG1nSvXUlPbngc1bEwCR197xLEAAQtejtwoKZmBMFm4PWTHGZEoQLjveW
wa91Gn4BQVNyCooRlkk0MHc09+c8PiKxTBViDfeNaUK75DpD9Al+Rti/W4a6ENPY
FSZYGKDapvxUH/t1BUcxS0LvM6L6PtzAfDYNF0+gxl47UQHmHOPSayexTFUScp/7
BuTDbJMK1RknCFCZ+cl91a9vjRLPjrEkOmobzWsPBSYwBzEPgalGmJQWsBzulMkO
OtB6hP/2Q7Id9iaGNkqhdnkhcASV8AYcjKHZqPaI2rEbzJ1SLm8fg3SwVR+C2o9b
AYqnuJo4ZD19aL69F1gx3a7F6B8d+7JYnevAU0M6lkVuJAPpIvH+60vp8tZA5ybD
L2StEdCZThDnFlIXGWM/vX3FK1sj6GZfZmZU6iZavKQ8/mRHhJ0r5KLluPls67Zp
5UwMQY4CnBLjffDO296Jkv3U8h2DIeFtsa0+NLQ3nVqxECcQQiGvzNx9uP0qLsKa
PSvokVlkb/1nZ4Y40VsZqmAk0qp5rLdTSF6LbFAMoahElMIFQJZmjgVxVi6Xx213
P1ZzpVzif/30KUEtpqEuf3RnmAcXI/kJ54ZVxzTcMN75oQNHv9S2Rn4vvMWm+K/n
Fg0mMWPdnlKdZ34sUw2nv7E0LLYEV44UUdwodlUR+MIavxAB9oSgh/5cvOivriDE
ye61gtC+mhBkYnPFHrZ/nTbf1lbpWDhMpJdtgI82/SgwxluMKmHbN0vP5UGgSpaM
2bHpCpN4KshNYthjCWTS/i/1S1bxqh/OIBP7kkBFtSCGSj7a/vTa7Ds8czJdcD1O
cDCk1rtYXmP7Ajm1bM/dHfVKAlsI4dlAz/cejG8SIu3a6wyZAlQUc90UZs1Llmpy
xJQJPihVJ663NEUo7Xbj5YRCheiRu58KFTyVyWBfRZOFk9tzI4zn5H0sJf6kDrvo
l0VICo+6YW+MGydqufsZahCi1cI9lnmWqKYwreGdN2oj9ZmhmLGsGSJJbNvE0q+i
xCwzyj02Vx5OEwTm7fCNuJm1AHQT28wzXIQEMPqEFrq68Zq7kTGep0bSjZP/1+k4
yPboDGZw+8EK+jetTE2+wc6bM8sVWmYKQaUuxjGcyEvboSxMBZyt8wcb2KKwZ/jY
j4tW6a404yRjPhiwE00zxnyOgAeT4N9lgFdItW4RS26YpF3PAQ/kulbTKyNbx+Ua
A4/5eKB/dY+Svu6Rgv4OqbGZbgLp8LpEeVoa3nATHH7uvnUb/h+gjvIvd+3HyVBa
+sq+HfaSD7IdgDYeCXDtihos4hY3WN5kcaRI+MwvHPfwoPYLuRMRUGLVFNC0tw84
1wFdGkKCyPE+9/iV5SnPOWt6esxDyxF/Ta9jdDmMamm9HxPGIPH+pT2KC1ht6G5s
aVp/+xhnix9jRpKxIylxwufiDXiAvdI9jG7EZSp6q/bgkkaonSEzrdz7/lz3hbgY
52U3Szko9CovATS7uq2M/NMoOwQKzegCrSRLsU34uJSaWWrSF1JjQIffB1y041rn
D30MZCzjeMLlO2V/+7OZ9nYtAYLcNPnAo5vRXNkvgUmrawcXR4UkTg+ObB1JdYM3
annPw3eb8vbfTLD4fvInyBUqoofLc9FVieYFjUnUkmsG6rXW4xFcMrVwrhbLIXqZ
9lxB2Ao/UhSBsz/lF5i3V/UtW7Ve4r7FUh5G1qGuoZMhXfg29dqyeIEVnNYfrNKl
PGrDclFOX6nLAG42QANFVZEj06338RBXjAiF4b4r2NhCfKAMG9F4HoxL3orOb9Yd
A+eXL9W/yfVQgM+dHlS5t2aUA3Uayso/NBf8roADDjb7hx48dPJJzBDSQqmyEPlc
GrAcIV0TUO+xdpEkS4y3/rMch+Zj+Ma8cRyTEQw2kfvR++Weu/3VJPOQFkwoeAll
SVFJg3QSp7SYMaS8X+eHEEhgo0P/wiOIYPGsIpfbGUPcwUs3nzqNjk27apMxwR+W
wK4WW04sga4jfAmXSF7lAEWgHow3MnI0jKCEcPTDsTt9ISIuKOkTWQ6790I7EFKY
fVfs/zfqfbUOdc46B1dkndhdjU3Zr7cGGO/0LT0GXSDTBtmWqmr08hNTw+j3Trzd
HTWSnSdpK3CVYyqEZh83zk6Rt86cg420d2Aoi2ZRj9knxTDNaUWGVXoOtOjZDNPN
+zUjZSGzp13+8/LHNY3AaPGUOo/WZ8YckQagKGNbWrY+MdcqL4nDDYbVRrEw5DRw
rFcKwqmyCXZbw/51QCenBfz8KqQ80NSw0fV8Z8iPN514EX1ZP4pNcpDygQBHAMt1
Rdm5PpEz6xa/w4DZCuwG64OC04v0oLGNTEY5K6lvkfdPiQXmyz3aFXtB6Zcub4uM
KxjY+4llOMRJA1irA8WGTTz0XgnqTq0z0m0VSoYRcqArLU0/k8v33OCQFBtx9zD0
W7dVpV9FWZll5XtVXYkeiB/PWd234gg902w5cSpRGX6+zq31kkcgVJMPSmdGPzX7
nf5LUdyGogIPo2r4LQLYip/ypgSFULkbzFRx/fje7WtmU4EWd60dISoQmHp14v7m
DpeYdq1simS2SIUcAq2f2bxbrnfwRX1TOWC7kGpiLB4YsmKlG1di+wR2LxG16lCP
pEVHCgDqTL//gEYCnd2SihnVdHZ1NiruGxY6PNirXPZmwShXr+vjsQlVHID888lJ
GxH+q+cIkp0ArMwfXtzsptLv0Iu3ww0T2BMmLqU8wJ3yLcnqDdZo07SJfkoVY4FB
xsNH/l6DzXWn6dwNgcOdkOW1AnYJlbKkqgxyKorsNyT5c+cmYbdLPg09B4PJRD9B
CzYkK6FUzw3k9P/ZD3WCweav2gk0QSCMzt0ZwSKYlWREoHCvkFVCkUANb3D9tbAC
cle6QEyDH4HvGo79SMI+fgRSalWH4Z5NZI5qt3OSB1HogrZ83igLUnyUGxOb8++Q
pu8XE5OCUA2GrtYNypGEfG8qgueoSWQ8Cpy0F9kyDUwzQ/qBQz2ZOgkJf1RyypVA
jQVTzcMgbFJc4/smXzwHpfTPJDEKkLSqqBQj0j81qU9MZntVZhtOJi3h/kbokRwM
2++y23L5EpRuJ0FLiYKgT08SRZfLhU2JsD2MoGFmR2D+jAQxeLx3+03+UnoqFTo4
cvG/SNzzG+o9oJ1UpUQLONe1GDZ8EwDjcD9EV1mB1EaukjI9Fa2wMxc+o2enQsDO
9dlsaM528lOJzO8j6tkdzDdTleOPMM9UF0L5fm/P8OCIuZM7C/B6rhq68hzEjhNl
e1H6dlEhqtfLSO9pXfbMxlVIZmxxZ9jet55NZFYzNB+M4LEzr/U0Rq8zoR2BKUbf
NpLQRTo2aFm0mXAYo1DJb0xSgqYTb0ZgSFISXp2z8HFj1UK5YVCxXXiS0no+uWuh
mXrLo5VKnqDEHE9B8Jg8obxkYjArpAaliNnMQ64tckjzdtUWIO9sn16Lyyn24hMz
8a/FLBpNV1RFfPAcHE7QShl0KgTST+iMllocfWrC1D5UkW4uFh1KxyYkE+HFCSzC
aQQBmBP35dgSDYY0Ev9obT/RplGxpjeILdnpsDekjEdklg/XJHASVsl31A5yZpE4
vagh3b6JVhF+6hfjEPIkAt6RZRiWfwffXZ+ZljSR213eLos+eGx8nXYVOK1k8BCN
z8++M4faS5wlWqtnR26A3+PTafmyp/4mKvTynfPhFnbFMBa5ygcojZqhnxhpq9C4
s5YkFalF5w17WEf+s1b9qFGbSzleb/qqywOxxfFWZvlGPpl3VBLG3Zd+TP5Lz3sx
fV8/xzoYRBhyNEeJZFjeOjPfayjswWlTAQVQ7kQfDFOQdyLM0Ew8iTyHHcrmlQvL
VYjb1bZHOYflkUVyEMB9vJOL3U6VLAYApw+Djg9D01smIHZuOJ839VYMGBC5+O4Z
xgpkrtUO4t0XF1glLZuy9VVfa20sQljtcey2OfXVJW6ZLwML320uNXhxsjH2LQPW
DcmsfkWbHQ3XXvr8CJ7RWnkITqrga6CcUFr9lx7f29s0Y4kRlioHN2lIBB2TGQid
ofH8hjZXl0dBPOv3KBgsc/ma5jsa1YRfIbyOqhasxNuz/KslriD6Hr9AyYOhSIfq
2xD8wMxqovxA0anD3btQgYkaCuM2iqXUqjArCSxbNxJiEw1Dw9TYstShVnT77lbN
xdb/P4Lmn1IHeKadRlwAeu704RgNLT6p83R0bq7hKAITZm62/1Y06Lfk3qkFi2H0
Fc+FPXx9AOIxQ2SXz4AYkbDgZY//JcSu2n4FmXArizchBTvnfNYNBBN5OGgtB+Bm
0wpwYtjcgQOmQ9cBboLJChQ5MnFqM/soN/U1NeV9vGcbRrp8Xvy1NsP1bXsei2di
66+nbi8+j8i5+8sMoXdmnMCqDWE1KkV7fOD9ny1EazkHw9oGT94lSO/1fn0P0CZv
PW1bCTb7GoS8cOnqe58JIhRp2ZZfi0yZkITQwsuIc/7Tu3OO8fsOEESWSq0+XpYv
FtaqLrZgWbONDHDDgFSk8fqHasYU9d2hlVGxio7M/qbv5TJPvn1w7tqVfoG/ORbn
1h8ddEP3E/gacYCMpMkF3RzAiL3Y5CWzH9HZ6KGOXFbpZlb1vRtoX1mTXkiBL91O
IpQupGbpHTMt+PtTJazTbNs7AO2/AnFLI+25ndxzL6ukSyHSbEK5wWihP743eEpu
cvPMVomZKJvsql7qLx3lA+GVii4GLL2dk3pZsvxB380qrS4vggXMpdQVeFixs7CS
e/uAy2a9xMMqVJCs0ZudAX8p7RRuVy/6UehbErJ+2P+8HfDQInI3SIV5A0XvDHu7
4yCt0hHxVjtmyl/Cktr3cdgUR/riAiDrN/x+UTTgvxpE7dDnMfoiqQ/K7Myig7P7
DVhRKouFLTni9qVVdGMRwwSg1blGDXFUs8MmdqIeApifbJKGJ4xItAsr8PDunUwf
1Cp/4sOJo/mKB/2a7Oz8d8eDSDRxDdC6um4Ugo5w3PH/6lNXHct46DhYqVW75u5J
mgurxFzzgKuu80HJrKEbHKQ/QfOXF2G/iVeZZpOn18WyOcN6C8DVnN1oUMte2E5W
Hy5rnoptOg7+juPqygBBe0uUSwLYg4b+OCjO0HUvIvlhwIxtyQvhakog9E7ULyup
TkTWedZvNCfho768/I2C8tgh+Oapa5pVH7cWQVcLhXviKDXCUzp/52JwTLBGYF1u
DN0zdIQNGCcn+WateVrKOalrArXUQEuq9fXGkll0UISj+TmN3dMgyhstTBmNgyB+
59/on4pxASxk+4VFgx/I9KxOH9qRfbjAP8LcaDhbsxH+E150r0Lp/nCmDRgoqVaL
Yt3dv+rf418pj41l5qog3EUsXfMeRwS9gWuVlO9GsBW2t3H9lh1/Gz2pgSD0KjiA
JDJBxxP4xS00SjOCrVaYLy4hercJbmzvo4tSS6CqIhTN3boCworKv2HbDubomQdv
Iwbxu30oqfC/w0HPGQ0V98GGwoKwGzw5I1wNXdTFxtDuYzUnBpECtqOFlVUbqVYJ
EcRTWDnhfguoMyxfRCqJBXSxulhLELsa4wOXk+NBfSGmDguh6itSpFXN0HPBjTBW
ElsqvA++6md6C2dnfPyG6OoLwc2wZ9g7nKpqvHX6yaGzYJRhGixl9y5OBH2a++jQ
6pa4pbrOXhc8AN5ns9zRDbitnc/+yJQxFFxi39MD7pQQE5XFNkIha4ZrYBtdgzxn
qyNQ1nkGhPPgRNk0AauAlgB9GYkyL3dQYbrCNGXbUpVMLDnzvIkI+/D++W5I6J/k
AfxlzNxs2xc8CUNYTbne4Xkmi02A26jagUyhMUXbNCm1MMHLaH+23PFMfhB3EFrE
6JGddBjkgvmmB4/VwesW9SQdSBwGgemfXuxZ1QnPQRP++MrsVUbPMBTKo7R+7hmH
s7KTuxotIubomnOGA5VPUxZmOCjDGN/xebVuGdBBjPO6WmGnkS9lIaqXfzuJRkE/
aBC+y6U0T6jwKAvCTGwJGIo/6edbS+o+xPh9yU6nqA9rzUaDBnFnoSszh+Y3qj28
vdEyHJg1U0av96/dEkiMN0bheU/iHbLODKE+54c4fAThCEPLgUdLdfe5f/0FdriN
oQi0NH3qhu+rYckk1jFu51fxpdesrfga0w8C9tre3HH709piYA/qjkq5hYq0MWuC
Xq963EqnJFzGvOolvL2FNUgU8uNiDxlJZxaDy6HGRUrke7Y/SuG5VPMj/pNW60XT
l9+A6AQYoHfU5hWiyFv3wv8Noqbfz1TAVmn7/YB87wZsfvHqcyXqt81HYaMLZioc
Dw/Su/D3iA0xADk2B4RDjsxhdrF4R658NtWPDoCA7HeN2/Ak6TE/jnyBqiY5I7LI
QoxN1P8MxbZI8jA+qQjO6Ck3oB3cEst264mFcDxB3bXgjxh8amaWnj/tC5/1TgCC
DVAdgEOZYeF4feCFAFpPAI9OQF6bFYWR/cEjQu0Z3zdEAX6Ozdm1JXzk4/JVsNhd
oegaO3Dwov6hgolFYSpat/eoRCoUFHiJ4bn+uKU/tkUebtQZ/bkW0S9KrmpOUY2U
c6qACXKmZNjWCWX/6FKG9R+2O3PZ5J/pNFiMqrj4mLhzw2yLPc6o78CkV1FY7jjL
GGVrmfPHcQvRdgKs55vvBUNG/7xm0mUKqPpIG+pOSB2IJiEZA+3b0+uSsBxodoc3
608bLYTi7cnsTq48lZsBwRMubygiJ4+4XWogr0BW55e26XbEZTMaOPXeQog4jgDA
vHUV1dMVOPJniCrg5W7C1r1RPDCNVtiBxA/s9OEhWKyH4phSzN/4mLq/xuhYE0UA
Z9GCjML37YKcUMzrig8bEbxfsnpHQy69dcIvsRbDQJfsQ64OyBiWs5FIOoRY0DSE
tdmHN5dqv/jTQGagBYZhPGwtJwMOxEt1im6buFDvM1opRZej9kqVix+pXOyR5C3M
1iHXmqAI1ewe2ibG7T9qebaekyg/jfLgzqSd9OIeMEA0BTULiC8bL2zxCOJDg5Vp
x6xcpE4m/rzY1zhFpdDZRD95FXwUjQeo4bCAytBdI+TJ+p0dJI1CY1geDYtcxCPi
uNNQ0uPf51wGkCn1RSREv1ukHXm+vc4DGekdTSu76/ln1kKRTzq2aynqh5E1OYZn
l6EOLeqivMZZCP8sjFRB0aKb537D4N3nRvl/uOm1Y8xiOf9iwS2KINqobGFsPFJm
cZMZybgQaH4Q7vdaRp69hdwYk2xGVc/YesWbTCqpqttIkVuS7rjJ0sxOFDE1iQ3B
OaLkOgTuFrvh2lulhokaYs6meqrpMaAvERRsarpCurWybLR+4bfROWGo3apuRNvt
aE7Kcx4vc0h3xzn0ch1dpuwf49TaRIw+O1wxytShAZ3QlyfB+rYdxeGh/gDBx8eN
h9rYeQCQqs9NZbpHfR4G6zSIl4mMdEo0WSzpsbDruyoqspZUHDB3HywHIJu2lGLF
vuPGkeqgeTqsemhRXllVnXEJ82Cp0LYkhgF0DqoabwgcL3Oe7/6Jc44irSY8DxWF
xDo0Lft4sZHOyS+G2G75ViCqSFe7SgWZwpNOxHVHwax/wUqBsNcmsTc3PGPIiCsy
RZe+9OZWDFK38cTuAwVIdF3E5F46QH5dg0ZWetZ6kDVoyUPf7SBKjIjHnRrTrq/7
6UtncgfnXjWqT1gkE3H1/6j6B62HTlb54iWDYts/k+GufbIQlk9NYSaJR8YIP/vN
jf0uWuFP1SzMkeZXgird/q2dOPJ+fsanpuvW8IYueQsiCAcSjBSxcazoaQ2ICE+l
V+GLYzTR2YulISQaaYex27ToxbpwVXN71+P7fLTzKsmZ/ZxyYrsjK34ADfqGEJ9n
QDzL9IkiQjYaVh3/NxbJrs0sY4M9MwUU7zMbt0TVPZDBgp/PDfExLeuC1xXD6+7F
EcXX04kCdtiBTpNcy/wcDss6m45EjkFPatBq0CR5uOtQAYq2ss8V7XUYuHbFwe5G
Fy7B8GsghR7/M/LSB16G6CPvYRsxOTW6c6OYRTFNoSAKSLgw1GzgNy3tq8mg3O9k
z1e78Rjv6k0KROCAHbxFlGRyarO7/w/TFvD/3ivDjvLMbchXHg1+AKpUpPekCJVq
I/lKIaBxqUgBhrR5uUjkF2Pn+mx5b5vvJaafE3+7gMVL/JVEEPP5RUAzLfrSQqKt
ze1zktwlieCAoba5h4ONXeFvpuobqCaWnwUqtgpsPUaMVHZo4pku1JRjz2iP4mES
6MrVDocHm2r/0OzKmD0UjmdXVKbAEpGORXkKfHYuppg11MnINPaocEBeB3zwp+iR
xL6IrzB4f61fIS+7VlouVWDVsD/txnYf2+qzku2Y/CKU/EB5ldIgUpH8jTEVzJf9
mIPHDqJVjR5h2wi5+pUezNl5IAbEW406HxgTpLfykB9tMEZIUbur4koNE4+2CTbg
6h5wbWX1SR7T01zB8BoIVldCFFs2/gshtK58YStH/l8NTDh2DQYckfyGrX4550c7
PvpvkinRHllrKK/J9sYb6wWwR06JhBvmejTavP0js/2biNzkycZbFP3jCuC4ZGMs
JXrNRa7IZc6uPJ4dkjxXkX79TuVnIoH5eUuKuWdtO0gFuDvDiG+6oVvFaifUtjK2
uXZThQ5zQMTn+4R2cDZlRzB86pOMYmzn0kvRd0nHnWc1Rznoupe6IEof3TEQheXX
rJTiBdqIQGm4lhgsJ0HkH7UUwO86rjl/TD2ReHCPt81V6Gl5iu7LlEzvI3UrJo1l
iV03pbF1HLODypcQweBXEFQcsRAfuwk1LAmEsg/EMT4EKVcXOBOjOBykQpMe9dLH
m4AgeW6piwdE7DrHXjtRGiHoixwtoMTGgcPJ9D69Ck0Jjh5AN3pWMggh0qCO8LDY
YDcyxbbTnzey8I99PYU5fr70YZC7eYCeOAlJzp0PGgD99Pm7K8jg1uCYHnblqIVA
/I3p6KNGUpYsvfRdJvBukV9eIFA3KW5WbZ5gZNp8WAeb3cZIEpqmorFt3Z2uNmpw
NuclQK5sNEEbl1vel6NoImLtTJ86+Vb28hjdu7GI60iuluf6yDMdHyfYkk70GLbU
7zJXL9VZXQgx1yvIJZlrR4C5OkL6hk+/wJL3F+sV61NBcyVTrp5/awYZOPHHAHOP
QgwtJ/mOiyg1fWDBSm6EnJqo5Y9VPx7VC9FxGlRx46whMzfjhymwxP1W2+ACDdH8
VN2DfyDkchKNQlvFiGGVGN4R3gEjvbzbSiv7b3AmhVlqEoYCJEfsEEMNFXTYPLYn
eq0Jv7sqtVVTV7Z06HQRsodzP6U2h5kiTjsOUiAwR2MTll2Zv/C8su/nyiGy0A4l
i6sRHukaS5MfaJiKljpZPe3rB7RVCHtKRR3VgWzoT6McMAUsUZmrygyvvIoM3fjy
J85dRPqnrh2tswhntvtgBxSKr1GRaDfaeUAlodVMZe7gfhLvsfYCt96Fd0Bpf75z
2tfJaj/oY9Su7PYp0LqPhxcPsnI1REMvkM38wn53RLkiwr4djouyOzjpNo3NVdoa
HBwr/Rf4KlM8MlGAfHyTfDfZgiqysPVlJ0IMXJJI6hL8h62/wcchVZRjI7fvKdgl
K5KE8M+wXcLI1JRW0OfU53NF8uwv0we5/zYZoD9Nv3axbLvziinqocev8pvkFF1m
LPlfB9+r4Df3YyfFlsW71asEfALL1AZuPnedDl6Riz91FhikOUMl9dC1fii/IiWb
zOESIgQbZd4TrKb49hq6FsE8tx3DKVgJBLyLOJcReDoSPaqUPAhlVKSvUMVQycbO
6PlPEysdcbCLa+J3eyq15Dlj3pqKaORljJlKCxbJUbmiQsp0pi6jBxqpTDsfwGY8
gBD5oNtxQLdvW69zYfLRB3YCwpCHrsZ31+56P6VNZlg5iV78dxFZz/M3NaspG2ib
EOwf0n4tYPaxKF5ZdKTwNDUgfmcLXLhVQIpX1RRuRAkYxL0Ek+L31w/L1U3o0fMG
P6Nkz+3Pm900uc3DEDXFZ5cnWegyCt8XqVpU8i7Mr7k26xUCtzYaBcSxxQGwgDjT
YfRMd1m5/dGGg80SkOJ9mfNIe7othUlWs2JcmptIfhUYdWS4SQ48FVpOrHStuScw
6AWctfRCk1BK2garJbQC+RR6C2qLgAxmyZs0uAkDFBlOR8YSK6Y35qtqWoM0Gn1o
4zZXBkKTfHhTFV0j3a7ADqb5epu1j7hitCCu0Pytac44SZ+wP9Tf143ia538Az4K
kq88S5vpOjQmbIhfde3F1VooCGVozEniXGyTe9ap0e/+4rz6yf5gHj11OzIFQIr4
Uc1SkkeqWaWTpVPA9AyqA5oMmSvRtubDfEdjwciWJ9mNeS1cuvdxuWH6yhaPYdVw
V3+hwrBudLN4VIiLDyLzNSNhDPbaQ1YZy8duHN4gw+55HfYUCAEYkXTgk1T5ZtZE
0rj2wC1RXD1F9O3Mcu5sZwGko8yjzcLQ37exqXjAs9aKnDv189xGYwOAbc3ASXgg
/t05l8O4dy/M3d7OBm8XG3WkekOBy30rw8ZILRmco6nmOrXKxyf5gW/AEpKN4h+6
tAhcMGm6cB/1OaYX8rH2nUiKUr1QTTxeEs8JPe0uQPQk51EJ1tHYCSSZiAmSNNEQ
7O3BSjtu/zmC/sgdbnj2xtLMVfEe17TUPUebZnU0SSzKi8C895ajci/MF5Qpt3vJ
tkWpPetSYlsM1cIh42OkVTpZS12iuBg1WmvqaV0dkUNLsJ088O5j0StqmgqvDflM
olPgtnHvzd3O8y57ln4cpi8EKipnvMq0iIqsJrEBtLp46gIZgEvQHv11c4WRjjbs
xx/okwg2IsGTjF/b45DgNov9mbZHaE/2U8oI/REwEHLLm0s7kaijtV9WWwRt3GJm
7qbeXHJeHa3A1hXWFlyRtzOU9GHh/2hPEZqGpkxmowJnvkyDNY618HsI8Izf7TNV
sa1bpcOk367paoMQEdYCgTZEGZIvoKDXZ5rhHNoWFt5tPP3Z8x83TWU4hlPnxJGg
a4TiJaz5S6GudJda6neq1+fe76nlGFHNhVvtsgs3bdYG7AAqTtRWWXjkQ3I+gAbS
jnGhc9vk//uHGz73cMy1SnoCTVmrbHPRA5mt8cL8r9ODTGpxShguQgsncSTb6kl2
jfzR1AFVSYgaTJT4/zxKnvByBTG45CJ0aUdkv0Z1qwFdnXWzsfXMmiN5ZvTsSqSi
XrKbMoukvc4MhL/boyXzZzigPHy10kDEr3o99WSIF1bgj2ipIV6nO5EdKm3DwE61
94gAc+0dxhzk4YEemh7Yp61x8F0wbLxQXditIkeAC4NX/zIZrU3SXtghmJ3qk9gm
HWxVNm39ezi/FuDpin2kQYcha9x4nwKqBTOorrjgb8d9Ws4mnzGujKkiw6G4RW4h
5QFLhk5f9+Yzl7OyLH5RCBaeSr7s8MV3/sJBhm0YLNcHxSs98lOGYi+8BO9jmE/4
/hMDXD6SrXKuZRFdb0RlvIv4bb41ZUmcxuQgjDl7NTenkPiAbu28lqlYfKwN4wwT
2ryZQMe+B/qZyLvI0HID13qwBn3ItDl7mc1MUVdtrxNtiuhOaOkEaIT7jBzA0qwg
OLbzo4ksiIESEKR7zw8bpRKtl6QtNy5NMkR2TDBI24NMhi01hlj5UCz9f8TdAp7d
ODqq9clf0Q5P7yVDrEidIuJgLSPLMAuA1xTjMdmWO20lfX0qqLew9lUGuuonAsMK
eax9WceJKv0/O6dVOViGJlcKodnN5PG7ImBtZ9dE3zTLtyisJ7Wsg8b9Ka6e9yPe
mtGiA/ToAbeEnYF0O1BABQ4DTvZ3rqMln2PZpMEj1ohHzDGawLVaFoZp5ZrsXyJi
XYVdXNxdxvN0axAq/a/DiOV1EanWBLCB5YjS4WPpa/HqpsaJkFlEV3baBtZcEww9
8cxdh12i4QeIwHsQXIIqN6DVVmRH0VRIupa6WCiKn1wM/OErSDSL4tApFiPMkMAD
xfUBxKbmwFTd6kivnmeHv7eqZmsnmbREk6nKleTfwN6Nc6orf2wdMoyvCAcj04YS
lVaUCMOx6vITg2lYEaBB588y5BJWXRWDfDV9bH4fpM4moZbL+v2d8EvfVOmAwub9
iS+mOQJiqZJAPjydIKxYRxZsalHvE3P9ywWj5wBH/T9wP6ydqjnubesDgUjtMTpt
oCwrhm4jbVadMR0AKz3ONvmjstk3TjsnxasQ1j6gyMque2zYRngU3QrqtQE3BWsg
g5eZkx8dAKiQnax9qgyYzfEkmsyUKGbPlqe03mJcPRhFryH//DUg6tEkm8Kw/86X
dq3UnMy/WS5Q63TSyZRN2ym3DOXIulJJJWF6ZIXmoN+xCi+daPHsTbHSEdzQtXJM
JUT+v3th6vI0FxTMy1Wnw4O4Ja9vY0+/WYPfFGtRZ5/poMCJAJrZxYjJA+5BevK3
DWsKiIZv9DHEJK54UM3s1L8AYsrJqKuKmEdnmXHF37Y9PeVf8uwo0PqcrK+1rtjK
EzbjNjcwjY6pWFW3fyFUUeGE6U8SVK/6+WxLavFyeiXA5H5NYR4sX5wh2OXg6O1x
l+L9UTUnLggesRoYSaCAnqdnwnkOTPaGufSxqve9tHDKfoFrWYNsH4ZAaxBG193k
hO9tQAOlRi4hM4EHrOtWC899EfLRyQScI92PQdIk+xOqSalEixRRLxLrPTlIvSA1
mpnHdKuAnnq7KUc+n/CSHCnWaQbR5A7sN0ImIZwCkHgwlzwyypSIjz1pXkF1ax+W
zQd33QrLKW91LW0zHC7J5enFftJuY6kZSLmJJM6cZ7OraYyGtarnmsM4zmJo6F+Q
vNcLxQUtVTQEQPwfY4avMnf19WtcoxdkVkqi3DBBcS/72uiCt6QwYlLUKleLdofK
CjfnX9bHsb6jNbX/pTxKcd/mgIgQ1eKBi5TmLCVMC6nQL6JjM5zmpcH4tWZn2e0u
7Mi0CotAzjyhDAP6KRt8UWiSDPzGwDwWB8pzfVdkLLjQmCg+AtAqdJCsOoriTiMk
jj5fI+V6D3SgPt+gUI+vJWu4sNQ9EZjHrZdaUqvtSvVjokaNl9HSEgr2QhZVIX1A
TA3EtMvZW9z8Y3/FgYR8ozJT+nlCtJaHfplIh+p61nQla0qjwYDxBEz0nq3oJnpv
oLRlzLIYaohgd4rM3kpZ81Oa6OCtPRrimlzEuA/HqbUEXj8MV2jfHhSy/6R4F3Lo
57TIGDN7T09/WQ6AaoVD6mXSygWTEJqcsElmrCTx0rKD2eC7V9ybZ++/E4nPEgP2
12GJ62OvJ1RzJlOQcoMzbY+Z3RdVSWbqLLOgLLnNPKQnD3eGrXnc6hO1Dl11ZBOn
i44GxJw3Uir4re7e1QO6pK0Mjop2ZuaA7t2a/a7lDbkP+Wx4NMdqVKGVi7NrLM/S
SzPFQxOcpJzMsB+1L7ws6TsEkEKIThFv6ACMYBPZOKwLZFDW/IlCK3hAkQ13aCLk
jULGl24m2CQfz4+4OhpQkr93jp1eqZm0BrkU+FMZcZpB7dpHTmTnxaF+9e5nxGby
rAljbp0qd6IV/v8fPWVCph/fyjeEllb3zBKXNWG1bYL1AJAw4VW3ajYSl4F6J9w4
H0W3+LbEzavqfjkjhlDWMU44nOmmJ8m+MvDKurTOBfiaF+Rew5wg/spbVbKKAZty
/yQjvCfMNS1FupZTY0z5/imTW4+0GV7oMheUVYRKxDjKdKzC2preWSVXdw2q0Lnb
afz1C+/KU7H87ScBWgwDv0w3IKuRDAqqoOSAFNd7z8hQn2ra6O7qlDy12yrQWwVv
6z77KXh9fnG/iJKXqZqJHdhsv32K2xn7pM2xSyfrM2WqBmNo5mwWmVNt9XIAS3E8
t+hB7ca609GercKs2zaaQmd9QpjIcm/bjZAPvLnvs4Fh2dOAzJrOk6VEoy6t8TOR
sqyTrusWvSctBwppXPU/9vVrP+NbSQ8cBpJIbI5EWFAc4FRyEhO7wWqv85W7kGGW
OzMhoBEqxerrRuQwnO0RcTirDdFkzo1l8+BFpFsI2DGvKqagL43x3pIRPba0dzJu
upiIAR6RLGOGJ5HCSGE3hkREaPSCN9w2mj4IscDlXRgWdsN2eK1um9jlj9jR9P9l
WIT6OaYUqI7UfUUnmVO2cN6yt52rxz/FtdbC2ado0mNlD7RE/GhvMPeML/kHrHvP
21wMRLKuxyA0C39jEGVI5wJIupdD8AJfEXJEUp1RL39hP/24yiQn5cdbbyFwqOrM
wnHmuDAFEWXjSIAYw9goLkQlTqnyids+JTZ2jRp0w5yJqiZBVF8X3gPIq0tiHzW5
/R+4VrEmk0ASLXuLwRerrF1VQvTuZdXKGmMayYbezsG774xpsefxiOvjpsBxcoMQ
cdY92FfC1w4GPcRevLEiwLk5O2jAth/2EPNUG73ryTSs30oZvmEBNN9uLZome7kY
w5abTx5u6RZeP72hwIlwldk8c4meVvFmj4tO79VTOfR0kHYAYgSyNw9zI7AbOhvw
fAn/1lLX3MUie+hPsHNIrPCRN+jGft8ssYEOMRW7Br/mimMaFq4Q6RTfrMzkx/ME
Ij0LFMQJGi6pqh29cZh/EWyd7Cp3VBycIYHAIKU7ooCzl1ajd6mD697besfha3Mc
6bla683RUuoCJGhiXiyZiIYffARZMPLXdvAlNFLhfTs0H8aFpRK/04iq8ciM1Gwk
lNwxkgFXPk85IV2rpyr/Djh2bvXnMinlk0ch1bCl/0KowG2IzXYfhfaSKm7iUxnL
c28MbCTIcppZU6LXmBrWLixWvlrhDi1UkxRGVc2VljZaofGQAE8BggdiFlA3ILiJ
f76RiQm2IzWu6H+H01KynlknJOgvDd/fkY5nVMpMO2xWyX/7gWBe6jnSaPNTIk/A
1Xh9gZpXLCJvZrU3lnznnIthN9yQ+UE7x4u2xlq+CzAwtxSsl36Y7jgalw+YHY1+
noqkd/WlZ17OkslX+0n2CclhlauXm4Au9FCt6oOZ6Vgz/G8wcD6D4uOhb7Xw5woy
XDTOMIEADM7S6lEFMAUqEZM7m8V/FIYPzP5ISN1EekMj16fpIX5lanCVsCzmxDGJ
NgnjQgUeN76xWazEMIGS8hc9x83waK13QRawA4JEnp3Anmb4sUSqcE0c+LBWLchh
W6CvDvjPVlwTe+wOFnXFCP3E5clKTq5i0KRChttWyv4g0gGOr5Ct0jjiD9QdvB/x
hlp4gVKlxqmg1YF/Ah8NwzFAXj0Ck0smxW6L4fg6ayC8kxcCkDbAc3c/EiD3THPY
vUtRDZ1PmIH0hBpICjBXRgQvb/8wDX0duju6rwYInrrxlDtMWlbo+hrPFtGI+sf8
NSizTuL0vs/l00MkcT9MbFSjAJ3PNUmL6OJEF/7ur8iUf00xkiQRmNzSk4Q9WBwH
ZDD5YOibOfMO1p8u+xAISyCf6UTkHWh6bL6ic/GbxAa1LYlRP32crbYKHoUPkzte
aRJIw2ciDrvgF/9g0YaxEaXo8UDU4RWwoy/dceRpcGCU0ZvTKIJeXviQIITbVUbI
Ly7PtJvguEqT6y9iNiMF5nCrvcVSsaUs3EJUUe3429PcNRUFxw4cS5cnOiwZ7oKr
cA/xDBYBPJVIJBYyoKY8wm/7IJnI1wOpWG8BCxS9q5G7m21Ei86YUXL0HRV62NF5
lzvezerGSOw6Mdu+W5SZUwTlLZqnVBhFncO7E+6IvQoQeZ7t1qLpRvoRwnrXtRY5
BtC9kjbCF3Rfp+1zfqRJlh8FDGISJoLXrDaigI48O+YpamfQ9auGtXfumqtMn7QD
p5UMtKE842mTEzipsiFQS6eEqT/UaG1mBL9IgAxYaVf9pF/MzkbY45f4yzIlIml6
vulSYesLdJPtylyyZyAIVpHMew4M7BpzJXJ+sPiCoUWlxflGYqizAiYRVamDFQLO
P235x8T7nIptKbDsDa2PtDg1k2lRsk7VgfzLlh2i5XwvQXTMSKsKEzL1XiC938HI
1gc5edADqieQNFfveoAGCxPDu3ZYEJSgc4EXrSSOWkSSUmpKKa64wPCoh0/C2QnE
42BxAOiEduBErn6dkVt9CImub2zcBgl1E08/SWiwZKjdSOdL2WEZ3jCUeTetvSAx
jzZNDBiSz3JmRPtbfi1eB3dPAwBZAkYVvc+9HIpJxK4/eCv6TeRkRbU8PAgVo7fw
XAPFH5JMw7nAkxTCx5rz2oZdzR6xuJJRUf+pDNbSdxrADMxckHrnfa+678dsWrP8
3lgTjYxn3ncUI/26cn79cU9gMpqATG9gzT3+vPkgDapzX6449c2sYOw8wpvSEF+u
cZjbtOu3AyNvOBObWc6bba4Y3RNS3ZGk6F+4QRYz41Smqg6KvaD9F93gQUKuTX8r
RyDORbUByMyRJ7hlRTGEMFMT/tb+snzUbRdAQqE01Iiw/1pou7r9UWTDUntMpgh8
q5fdcL5zNQgqV7VARlFeduTuCM6DbDeA3HBa6e6vugbNeVQWt3qPDmdPiXXOL4LX
z7bFwEZo9grRqflD3G+xM/XhrW7/ir9oNXObWAgEpMVPDU2qosx8jAEybnFN1J2v
aHfFcmjOePoIIIIEUZjNxT5RN9YlDBgVFP3rgjp4tab9d5vzzgI6Pi0+xkigjS66
QmlnyTcrs+446FXna4wOiCSove/dNGUWF9Ij6caU8Dzt4VuouiU2Azt122aGOUGQ
MKEjzl0v57dHrl0mx1S+lVRbVZAYT0F68+sY7QxA05fawpNpVxR6yP7SvZ+MT7ZK
TVX7dscqO6+LyfhJDdZrm13JqU03sNwi+bpTQhwu31n0Mb3QhscKg9qbaXn+Ij81
D752crxuyguw6BREwZEwvIt+rxVMj0QSfhLdSROFAJzYz83083Ou0eNQXdruquAu
cfBMDLh14YFuvbctTjq1zSMXjsmcx3MZEPPLcwHjGdsHZwRVa1dVFTHqPyZpUFDF
Gf8vzQUAZvDV8FvQaKr5OETORF06c60zE31uyrj0jFDcHkyOjD+lXuniFuysBWBN
f2BcA/1931gR4b2mif1UVYsIdlYRBoEv8mTN4FCqQQhF22I+2EZu6U06C6SV7qin
zlseB0r2286p5qBv1/xucitV5kSXq+4D00UR529TeOr/upSA/vijJM1biJZjxzom
GEtNxWDBIE7ZUpPRc8vsLCqkcdc+mBIp4oKJzJb30q11mwEqn9fl43LFMlMMPIwQ
+WjdHD61sbrjEe/WidrMcYfjONNy6xRWYKRMOAWfpIRIP7iTSk5dim54mv4Daxza
ZnJbYHoXlrBdekz/jDlanZeZSEI4G80aNikIS4gHH8dINWJNk2oYu0+a39rqV5C0
KLA5NVeYXc/ZLI75yD8C4IgAe3EUgatJvGG+z1DejhM3fQ6eoipL0pKhmYquMQUX
PIsVlAZEuC2ZH22cEJjRma1MfYOf5rrNmcLucMJrV70p0pyX66MWLYhG94x+Xqv2
ZgnDLCW7kY8pEii24QpQHv06LjZo9reiX3PXt+ivcDP/4AQs2viNvGcUAtSmo4TE
zVMp1KbTQzDQ/nA1KL9fei4CLcLsL66dOAHtufKpTC99oL1xiYyBn/UE5JZYk7jO
kBk+B9cO36Oc1VGRc8ddxzlyBZz1UjPZoUFbArCKi7bvfD53bN9FOJk0KGql+RvM
MTnv6vOaTMM6OkTfu8j2lORaYQCkqPvySOi1Bnq4BFMvY3vm/rBiQpyFDHEnd2+L
FMgCYS6sFMvrriSvzuwOIw3kBEnB+PanFQurAtInbUFyDKoY1VY9qEnFOfwWl4XU
NoX/3a28B2GrWijCYwJN1piz502wmc/LPjv+o5v7xAcYKjlAAVbxyvLDbP7mH6fe
WzkFp8nmp6IGG09UeghqVHPkQiW4KMoc7iF6qzIQ1mKrLooMXIGliS7qTgpsX17U
PwGso9+tGwpnbEVgnooA7SzUiFwq3f54wxXMkjLRyF1NuWI8u7Wm9qNygwpj4v4O
bgNVEAEy7qJO3ZHRwy1r5EDpGZIwbbijjWMERQp1Aatvw8rsDTlewEBsLycqdfg0
NNoM1AMH+rBUjM5B+gacA5rSnMtEr26P0WBbtKhP/yXUQnP2NYqD1CtNk+WaHHPF
rkwjXBVe4ITC8tmRR7ECzINQbJXDuLvnQeU4kU2roX65jsFaj10ZjyG/CNdSNWkE
pOb0hg5eDVnMFsm24GH+7T/6o5nSPSCiWakQCajnIfZ+qqKmEFf0JgZ2KpzcQw8e
gHutN/++KFrqs0A+5G5B8tVwvG7j5rdgqkhcyBkjy9HUBSyDQ77HYyd6JjSGqOd2
Y1KzKseXYVKJfMxtSx1w9oRO+StVAMquUiaZZ6CcPl+TK4nidkxJohjQJSirNiwl
ey9jcs4rJ54uDFpESxJyJO7dyBtj6gYITiBlapDsebsNBSXAxj47fI2gGaRfCOpW
64xCwFo7UIw1IP4O6TV515RGBMh8UTKzWm8s8P5RPn9k83bC01FtknuAeCJz3y5e
/sSyYIKBKcoGhD9szvZjQ7NisW0LDhguBjbw1EuK5qVpy4Mptgt40rJPuPSdqvab
Uzgk742aUUKe/+m2C3JtNDCs5oLAU2moPHdypSfu1p8ylYPd65kTojRRt0ZyTUCL
LaETF+tWYyIVBygPqtBV+e2RUTeAWmNee+dMD9z5XyIqNZwIYvS/KwWaJwEP0bw8
HSPp/AtTEg9e2/3gUP3BBi2CEIBHbQucR4kyLIoTupLJ3JitVVqXuvD98Yb7X0+7
k17s3XgIwYrQuXQVxj9cdbDiyknBTNj3VMUiganI1/aA8w13DzBYvFmYqjZ1PkIw
74D0w4OF84Qi1OnkYgqvOYnvHchRrXwKBgYGZEYd8H6n552LPe84mpTGSDGN2CKM
RmWPS8eXBAIls8Wap7Eb5yU+VNhiYhIZc5nkcqNemIT1BUPlFNvzyfj0ohygGlOD
F3QOC4klezOWmX5Sg20bjCc875PpWsRn1/EukDr2uHm8kt/Cuv7bG7Ei4tIyuQzO
+FH+DwvXtrNf329t7Lo/KiQn8ZDlRjsaQ+5LkTRfZ5Jn3OW7Ez2HCcdREolhX+nr
2My1FtEUdgMtkkFj38zZpHRkW/f+KxbKjEpCdzqKftVEqF7XUnMEFoMmLpbS9gqM
9uKihzwD+Kekwq1L8rmvNjfiOfbYnhq05xiFkAV1Q4JlQsqLIxKxTeBqacZSA64h
ECxR9fdxHg9agxRt5MYE1aMVDLgC4NSBuusTk7lMf1FlEPMxGlJGZYY2yRSVYE5t
wFMKyj5fVwLHNfxG1K7GG/zPt3vlVYyYutFc9pLAtsLrRlOrv5z+UutRQDzfYBpT
YQQR/U/6hNugtntrJf8EfHclmynkn6Db7ardh1C6WogBilyp7zt9aaodUMxduYuT
LbMCrZ0Ze4gNoHcpW3XH9wZTjYtr1StqCXjFY6Xj9Synma+3l1MWe0dMU/fEnuYc
JcWQrPVVS/TDjFkAwil2NvIcid5V1RA19RX4VesYFmwRTTh8JivfBunTl8Jg7YtV
IKU2KERTuSs18KbyrCytFhypG9K4P1u7pb1R0do4okGw/5g+zUeav/yo2GP4L1S5
XTtbjudBNEsGL4jtDa1jyj/0bttVXXdiBoR4bP5L2x+nvscEpm1iJpPhNd0QEfzb
2HuOGc1wHIC1ElwuNZBafFoD3o9srueWYF0KgHVzHyIgY8w1fD3yhJaJGK4C4+Rp
18bPVPUeFO+PYvS4sA8Oen7Ji6AWMNkko+2VsRwGhpqbmgW8xwX9zxnO5kd6/plT
GBBFqfCOwCfqC7mwyU/wqziSWp/cFnmw+P3KEDsRvlpuJBQM0jfMEucW3GX9XUkY
+uhoOOliIE3TK+fazzNHOi0iFr1wgU0XmbpWLClfH7IJJHPVfXLJ+25IZHPGLuE+
p1KF2o5c82O5fiBcQ7mv2ArGgLLppA5KwIzoX/TR01TihfEq9vRQMrSdaCKY7IUn
/pq54Z3QCEii8QQM/wMvXpyGKTKhwZeB94c2cHbWvJX6zI7Vg7E3fgTXpVoSu/OY
iX5cLYQto8yA57cbRxFxgmhg7K5Fdr5GrfEWbPJr7yazJtERpZersJggcst5HcqO
V1rlB9ffiKgH8G3rFcJ63DNVPYpUyvVuJk2WVcaGn8yF08mTDHhauhaA5BBcOt5b
h3pikVNuagtbBh2dXzAbsdxekoE5AlF+YB2lGYChDiycw+RKwgyctbfsLm9DQPik
8rEcip5V1C1DuqktsNc5bjgYJxB4ZRPckZWfW8yx6V+xdmQnE6IEd96jks5S3oEV
88sv1qrK/i+ht1AoBUM6viK8JzJXw6GwSakwxQCyGLY+uP4mJy6R3RaQ82vWozlU
MpPu0716Vs9SxqS300DpYDm4bsq+uGefjOWlCW42BHq6qd6k94oa8V8BPoRImljF
SKkvCvY+uzTj8GANsDFZ+CFXxbcKFouWRhGM9+0h5cqeaxlsMdy3slQCH0R0FC8G
YHV4d+pIBg2jEc2+g4WinSq4NNr93mBY2kcai8QXGpZqlzZF8z5WdIvEMbUv/OuM
Xh8UbdQhG+YPQxy159M+5ITJm242odlUdK7nbG+oQDg9ourNnpenbANUNAg9QElh
/W5sKMDTavkh9zuIt8yw0OE4jvsg2I/EUZpdAiJnwlmxVFMeivqTp7F8mYIXnKg9
+njwf6+pqWOI/xNGSYsz65t7bceBRQ34Fp2Mvy0E9kHc8y+IgqgqKtiVeoAZWK7d
MCU+K9CyC5uPwaj6sbEcgLlkPuFg+UCAr867IAScijerI8/z0Vz0QG6udEOL0V8H
qKg9PxrO59YYvtHQpmRwkpn0sZMMe/ACYZbUTYZIPrDa0pgfEai/75ekFjCAVpjq
8Yk9aiBtybOmkJYJ99FXU4tUPUv4Zi9QmSZW2kQrW/wpQL/gP369jzfTM5QDUbdP
Q7AjaKmB8oFQJJp6rGn6qonuvbY8uuMd9pGSKVsXTYvLT8n8D23JP6PQhuQkrC8Y
1IJ6Mn0UleiafPwSWzu5uvAif1e7yWRR4DOOlmuMLL1FESrfkyg44F77KrjWDVoC
sM2HdG/CcIP+3TOj63byNTD+PmHbw/6s1nOjqRX+7hmQYEloODILn4tDZOZSBGVi
0nXLE+BSjeg7mBCHcRQOtuL+0FIpPn1NyTmJheUchBre8oiY3Et1cwgqZb5y/paF
W/Ls4qlNK8zPgJ/puv4QsXKlsQA0nZlsA+kFjf9JKUCodeZR16Lb7twMfHz3/WZe
YvBNOPC3LY1fIOzeD9u6AkeAJqc0lRDvr5rZ9/EvpNc8sddjwIvD9uGGOpMSZMve
MmbtMBnJYuEcSJNDaTFQeBxslDWRdaA1ILKssNXjazWbTbyR8tmM4I7G5yT3H1Eu
uPhlJV24TiqcQVMnOQgNzCEBVdpo8tlDdoZstZvNULB9vx5j4SRokUAbFZH7NWsn
j5NHNnEdWnjHfgvZwSTwUcY3jbKBBHVIu5nQ8BB4jfgbOwP66vcVtc1JtyUWnRR0
zKsQF9rgpQdcCDW3ZMLx8RKD1Icro+dReJwIh8LoVibeHlZsTcm4ea0iXaokHATk
YB7DJFTUR4XkPCLkOIr8uXZOWzEFzD0x6hgipjJmP63zqi94CbPfOoIZM2vlXGVR
2cJ8OQ7ZSodmgUJAsoiOBCA2GhblqkI7j3pvHXFim3NX9p7CRqdg3Z9DFEu4AxmA
FDzTdhS5E3ARgs1gkE356G05ZQHhp97i6MjLOuw2C9Nt+fFGxGZEL2vKv7fZuFh1
Fy0aQE6M+Pd6WvsSmu2S6ND5hBCVnqjoL/1UpYPVBx3T+gGk7MmNRQS/bPXRxOTR
ukOG6Gepj66TsTDRBAld7Qeul0ZdW5+B9khkoQRyaieLF8o2DfohjMCMavdTAnbg
89VHwCFaEO4O+Zv5TqhC27QKAoSKzM51b2lrEGnPTBAXhm35y7DILDvJiK8uWN2s
fgubXtlvW2cM9WMk8EdPtmMnUYrIFyDzjzJd+JPPRVBMZCRPS4MCas9tAEQHf4zk
irolZspTUnG+h7DzHZlWZ9RCpnmgLrE5NpmJcm93HVIp0bT5eL7LEMT5h7thKlZC
vFPu1zOeHk6WlntHJI1ViobMglzhClNmm51wXlaFx2YK7ir5cK0SE9R8BXTVpJJM
ey0iu2hLf1H1DA+SftzEdv6BNUMkh8bZDwLHJIGDjj/xyWzb4oFWqnOgvWPOX/F4
Na2CJtx5/nPmmXTRNCWqK2SjWEdg4WLUZBW4uH+frcaG4/gjxRd645ee+VhtZ8ba
KpYEE4duZatFj081GaOnDZs8oVypDtFnrRtN+GSJsb8WfbYwGSOV7erxHpeh/ih4
IOYxmXzLchIKQ6UecK8ub71eNA0zTUhu9olglJPQ1ngEZsdRUThn51T7qJx9/jwK
K1hv8HrlC5Mz+YLL5wWrRItGL7OLhzjjG8/pbXOIOosIHITUFlEkdDy3IA6As9IK
D5KO7iFOXdZP1ls+o/wJ9lOZIGjDrZ1XK18jOJFBwesAhIBpcQIjXdO6Y2OYO/ma
j6MoAnuBMS7BRz1IjLhZcoB772BecC4igpUcK4OuLFlWLVDwophLkr8bwaimuFjc
DZZvw8I9uHYw8D73OnIWXUe801Al9FXtaEDVXTWRsv2D8VS2OpB8pZpdvErbbG3M
/0GCztDXtiWnd+6hCOC6SaGuF3/19cb2Pl8vWFxpQ72kjrVN8CpRwEbVDcTqC+Ij
qz7ZE6RfQl7CGPqpaS5lHcFgtwic8rv6KtutxX9y9ZzDQbNduvmBkdaP0d0WjtT8
MdlHSuL3mCHftKZ2C34yvxHVpbnxukaPgQwLtO9xPuOz+B5gKJZRHWAlmGW0jhCT
rdr5ZGBS36MKwgWQNgG+xfMHaMuVfqKqjizDAuPfYGoKL19QK04dnH9r+RyoWbFL
f7Fb2e8OhIckqm+jLL6WqQIvQ+DwG6GlbdMGLQghxssPQonTbVJzjaXH5/8BzXTT
020EKr7Kv9HCM+DN+atSgJnc1paap82+3HtoXThaq91gu6Nu2GaMIedxbORnas+4
9v+dScOuBuEqiidh35lb380ZZGgiqsYlDt4Ncw59S8LpXXVb3ptUCjfIYSXQh9Uz
OFJqNt/zDW/wPt43M4I83LGDGa+T8/CUFIG8kTeq/b7jSJhtW1g6tq0wDXkTPBZM
V+8H9rBUPAnMtuMCsExLXWhtwE0jHfBVCg9usGx1wOc6WZSsL/oMiTl+Q9Nu7q9E
6wVi8fODnwNak/gm+duexWvY+LUh+6RXPhrtw6CISy0bMBdrnAQhYOodLVI7aYEn
A0a7fCpOF2zk5yXU0mJLsiXSBm9MpUzV/rj7A6DOUMlBQKSBJp6K8ESe+Ya5D4IA
BsqBuXcaeNuTtvCz+w2wAjCC7Hmd+5OhOsCdWVnoV+9N3QqPo9VLsDgmp7hWK/95
gSxNq6xmvmKyNkrTyZ/TyG1GgXI52DVtIMIw8djswqUFo86HJC+/vPar41KXVTCO
138uv9lRwn2DXt3PKB5Gd7ern6pzKEeF7mQj43I7gLVfUAIreFnmuq+zqLXv7xqN
OG6hYvA0P5pasdTmeCDO0g7yhhCeg4EC1bwckuV6kMJUx0aWWaXuYXatN/PJpfuK
qGTsi8nNqcK2o/m0bfMUmGmP8soD+X8/IemxrA6NTfUt11RtYGOxS9vjPs6ULpEO
ccH69KppC8V7GT3KjKhAcdcRQ3kjIEnFIUNB9Dt0AqW82XQ1X+F38eQcpjd4eW5l
D8Fks/PIbtKMAZIXrJY963VJ3CNkJ4t8Gxq/YLJebn3dMMbmpqSJo9tClde8DXo/
eMS8wcKqbESSmP5jtCK4PFUchognjiMvHkI6PwFokXwAx2fifwz8vWeYG2jQwd2x
kvEArZb2vkaF+8zuNtSmbtLL5UbawsisGiWqGDAAFfYX6vmOUJ9Ml6Y8Ou2aa1EB
2VZPgB7IvGtYXmc2q8e1DozK8zf1KyO7n0oEoT5nQ+rOqwVhteWAGBl3PUeyEz8U
2C6408ShVG5kh62tXn94EbpElxY6t6ghSwS4zxvV1igEW+ZxwhrHLLV6nx7+lbIw
uVa7jJA+F+v2OMVS/PCv/FiNzEIFPekgg1HXcMMFGoP5PqnNGEQN8kaSMZ7ZDDzX
koBzaP4vMe4J9VdRVGmKm2578tWkWRuhrZdNFUffSCQC3Y9ymREu4UYmk70isZrz
8so+9AX9P3fo8qsKP/BKNVNub/jJO6eh0nkExpbuiqPQsPB39pGTV9JNtnpbAMXS
DtIRYUM4ZSL2HdRJe4RxVKp98UCr1NKFxw5Z7nRQ6Tgypif+1tkCyMlmp2tw0iY0
/13Lfc1GYjriHZjr+YGtybOh+wyruIZzDakaz/ssaebT9hochwvC8C2an9+DoIU3
yAYEQSBt+Qgb2HbORdCm9KrTHQv+t7Gu7WimNugcy3j4GDv/CRsPMQCxhHyRI7EC
/fYPgcxmAx5PRhY5flXRK15twnLaaF9pX6HtRN//DllCM+a29PC9b/ANqkNjXOXE
7u8FkKkVa2A4sB7ULsDTdlsZULXPHKtShyINPN93HDUn7GSsau5bkexovHxT52Wz
d4bPYoAQwEdya/WdLfRuAzNumaaI0jgxbIg9yAm3wx58pTdup87AA4r297zpqQT8
JBVU4rEBJCajkgvypKuo1ZTXGz/2XgI3M1p/jO1xICe4gckH+O+WtLaMgaltOiNi
1laBISYL75fy+NTtvtccBWFJZ5FQoBeyUdpD5yOb+WwfGL7+MIreDQpo0T+Tpbb3
1n0OSRygJwvhy0zyjs1UesAWG9PegBXCVbz720dK602oUBbvS5zCplRm9RhEPMxK
Lsq+5QpnFx2S6m7vim+vKgVdRhOe5P7UMErhPonrAwsBMCZH2r0hcwlqclpvFSEx
KrbTPY80wL53VH9S4WrCvLs51GseAo9igZxI2wVt8M3TvgHbPY0Vqf4ppnibs/bq
4AuNkWYVUsAeybgKaqbr/CbrazRBzGykYvYXWbqQwZfiqET0nZ9L3Ld94Dk+ssrk
kYNYxjOr4aLZQywX43k4ipt1yd0YlaWoBjFI5nvbu7L8Ylkk6Go5S9TonXINCBv3
47FYZ9Jf55pLtCKsbG0GMeWuLok9rUZ6zMEUWaBiN5Sv/hCf8Pbo+SCTNNBqP1Yy
ni0Vh7w9GnHj7kUg8Old7TS6QHj2BXzSeYkHuJn5OKMuZ7kGViJ/pxsCZSs++wby
7p86xJaGdP/ph8w2W3uHmIHYRacBY+Ei9saXqHCtTKQz+wRk2kSI01q3ZSetmd7S
ZRq7Kf37zUrYX7e2G3XCShigHGRZcvuLZhDrHDtOWCKm2caJ6WU0ui/SeatOeusY
Xoe9ClK0qOvnJgJTCtY700Jxbvw76Mb5m8JrHcUryUYVWOOCm3rpHShtosvP1qim
pxIq5vIDTgoeCviGP0CwdVcC9nH/NNpzg95FqOEQNnUJuHCmZ3bXOQ2LYKpgDOKC
uhmmUIan9mGlv8BNx0Gd4F37ZnJ2vdQ10bpAq04wFcJ3iulGThceFrX/igETHpLf
buuDsyZWSkImopz0eJ0fkkwYb4Ob/cxyQ4zxyLZMLW6EPD6CBoaEOl/XLxIP2RT6
/NWUyoQ4HFRlL/pP+nLG6bD0TeFZImK+wP2m8U4MZH8vuVNnVHkLc/92YnpjtlCg
mJEdi4PxdsNxs2cBzPq5pLAcuwi1c+WkQCIVg6gqyoP6LTTK6eU8XA6enuPk/qSr
yPHEVtRWR0vKeXanFJ9/EvUSPm7MhU38FcQOCfF5S2fVfsbb+wiChTpgh6w9ooeV
dqiFfRycIFkIUh/DmB92Q0FctjH6TDrgF2AjWISWwafEDp+2ohTaNUiFLYzdnReF
JPlxS/jORGMbZpAyBOVYeyRiIul3USO+ozMHs2ntLD/AXvkKnX9WmyzXa+u7K8/b
77NkiKNWsXmCkkdg3ol1WpOYRpzbNl4/k8BedFSTYXwneC2JV3Aw4hqZaLuGVrSa
eVuY+jnpVebzqxl+b0VW7mQGr/u1dJo7nCMnhQAAIiYuUxWBXf31O0myTN0UHnkA
6+KvqGZj4oulILdAJ1BdByQ0G3aUVuNm933uMjLdklNJfMhCIsaYMmSboONzwwT5
aA8DSZvSi215a+ZIB075yF/zR2a1bQ5hmW4wFk2l6KrXdGyYokLvNAT9lwTww6ep
XS6rNYzLlghOcy4pTjgg3oIWIidtgkKt/0saQMqV00cJNaHnxlPKEkEOEqmoql5S
cJQPsp11K2lJBpUNHPtQ+uIqyhGhZu0BrEq5pQG/Rn8Uj/no0lYWVbBNRHhUdxck
S6NWcI0aNW81z3c7fEzdBX1EfRXnq6IuwL11+I5BA61Hz//1hZCSvo3mWliyvbmz
IISnIthueRAlM7b1p2sZ0CWw5QmIOyLFMZgrecKWRyF8LXnXBsoTo6io7T4RXHbl
y+9K/19xws8OAVSh+ZNSsTbqkIXYDFYKKTk8Zgt2cVGKM8rT85pSCpZtBrinPpyB
MFDaSqEI6YK/ouaqRggjLlewkz/GtV+nPHiBmcFgDUQ+c3InbE+sLYijR7d0ae71
sfjs+flgZk5ae6nxvZ00dw/r6xJeXBa29oZ05qNHFjWpHocVaoK937xceFmYTNpl
tPlon0syr/RCANngKsxDx5UGSPakxff2a1YK1yIpIeBtfgfAm+qKOCfc3BHhp4e+
k7FTWprNi73r7Eb+8/AQ7874qqZKvxfxbDPlQdBCcUZFA/ySX72STKJQ5Bu2MaBN
SfE9hy52bR5ji4meIFFt8jB9xwcghLcej0FX3NmcmPvcQUKZSY7VZfbbfua0Ys+Y
QWf1QCpK57Ij431iAZB1q56IwRBM3IqtLVpLe26TMwzDTdTM/VqVsMPJnz7L6+CD
yIQniRm/rsi8nzrLzb0s0paEBu39AL0rWsq1a2N5aU+5DAuh0EvBBblp16RLcV8m
Z23YItZ40FqARRttb42undd4OlmY0B/t1rTpkMfah9eMlJaykX1MQow1XM2XSGMJ
Atja8gBl9J+IcC9YjjgPg039xfO/3JIL5kSAT63KEv63B9W5QN24449+w9NDibe+
SJvRTbVs/YfilDD3HinNL/0zj6aXE0q6ucpNx2rudsJFbAWXvLQ9mVF/YzMdWaax
VGle1Aqger7uyh2R1JJOVCWv46Q26ncta/fBQKbJhe5nGY1wsKm+u/4bjF65duvL
2TrIOoreHR0kCTZT4XNj28N6JftSPi5FbwJdiySNI5hSzRYUBDkS9FirG9Z1/4gT
HfaNdSsGEC9GzP/rpO4VQjNEduh9VFeo8mxkBXfTLucWfvr0Ye21MV6eRhm2hYEV
6DXSSNKlU08nsybfXcyXs7P7VqQSFZIVcRgtrNoqJwMSsYhy6y48i/8BTQ3noyNH
qP3cJm0qUgxS9dPLSNNYf3M33IjeUNhunsAkQSOh/tfPUKev8bE3pqoVWxWWRixB
qDv+gZ/+Co5rq04QqY46OwqzFelgPBrsxcmGZCc9BS3poBF0IJrW9GwlGVuRHwp1
T6YOPamvCRjIRkime8q5BD9cjWFDHHMWuh4qj+uBCL9D6kIRbCMAmFsn12aGjHH9
2wICxmwBB6OxHbO0LQJz+EslMoQGGAAwzArexbZUEX5091jDmGlN3UeyTcDouYL9
sMf7Sip2elWdHe6LHw6ABFDO9gk4q/aNFEcmUO1vfKs+rxkhoS/zPaQ93aX9/60O
9DVn0v0oL9CSzM2afm7zc/4NbH2hfo5o2mZAvmg5cRtfgszn6PfLTnspwgUVZ83Z
iHFus0AxjjGdWi6dtfpRDCBLrv8OJsgEpIWVLHmr193+BhIe4+7/cprr4V7/FKzI
4+ZUSlVWLPK+h0HDVRQwTn1kvQR4nSfxd+9FzHx6V/aQlYtekSzlLNzkVhLaoUZ5
6Pj0czGuvmeIrXdipZ3rsPBMwynKRnP3COFB4IlWdQFBTyrx/UaFW3MGEUX7YdlN
XiATxZcxJzbkwXT3nZ+/VMbo8B2RP7YqrD+sTgbz3k7C/REyoqhNFNqPmh7uoLU3
uWoTkih5CsUwAXHzvKpoYn2cqK9fawfQDC9Wz09ALSN4UejFmgcp1yTth1AzidL8
v7a0b7Vb91zcHK3D27Z1VHHCfrMvL0eilmrCRE0eJE0SZwmvWtnxDcjkqCPHTdOm
XXlEiBLsTMMcgUYUGMBssn0Q9j+uhnGXGouhPofLnvMVO5gh1LrSX/WL1uTZPiDR
YYWvu5PsJUYXZjhNZhwybLcmME8orwFOVcm9xlqdWKyrGyRQ6NivIHBwGDEEIScO
jHHkE38hcYhJ9ikFIzOnNLr70IXKejJmBlH+D6KcLkFo7UNnLfaxPtKU9CXJV7pO
Va2+kx4QhEqPKqJqA6LIbB+2YmDf4nEkv9cVZTpnqgLCBYT5ubDZ20puGoUYmW7e
JYSxo5lh7cI1zcD3lyQMHxvNoPdBIn7tXmZYaxAsK8OfLwcREYQGS5xLY8OE2Ilb
tdMUZEv4+dqOOKqnpzl2+x9/JTBcbOXn7ElChuxJ+NOGDbotileb4B97rL4h36zk
UlY7gIe6fOp1NvSle/cbqV/w4i/3yUUsGlAgxWd0XfXZrRGGOwhyOOLFDCzW+6Ec
9Zwqg3OcDn5vgFGz/w3iB2V9w80Q0xvJ6HB76wunIlVhFW7R/uyAoS8X+OG0ZTn7
e64yliG6GaLUVZkWJfSanIVGk9Lj/JFS9ILtn8vWVFDYykvxo2NoSMxyb9qiH45c
iNbNeWp4BLiCx89SMWhB6aonbvCVB1e2Z5PyNgyzfbATyI65QmgRLwdOa3OfsUIK
DwbYtLkv6SDZ4iWTDi6IK3vJy2Arx0z0ECoyzF6Kxb3oICPb291i90geRvCLYK4I
mWXmlqcOS8WHO1Zjbb+HrWw3wKRzzOQlcN4e67P5wR+6GmbyCf+K95qEEpLfdXJa
0O0BCkGx+BdW/hXchixKKBFsa2dfB8ehyVSvb1ZRQDbQ4lO4dBU6PongNkdUK1w4
VHv4cGAREFZZ7/q1uPmx0NlIoQmKAddbwr5DmHTQWWjmz7T7kMsMTQhAKM/FoCvb
NzYWGdU4ogHn3XkqV7dN9qxezGmvfqfvWMQXkmkhWDmWq988nnMw0ULAXe1l37+1
OPpxK4VW8dRY08wxwwwrIMALKxrCOMuNcmFHi/vLok6uCNipaqFouf6NmZ17dty6
vMv8uuWSjRE5fIYvdYIOrDYKuulfjK06PvNKLUH3WdhxPW07Qxf+rYJc3zIpaLv7
M7X8AXZMCTspDqajjKZW4INJxNHUFMSW3+eu25DX+al7GatG0gyDrueKHa7wYgTx
BTSPF+9h3cY/M0aX0sdZS/JVART518fBKi9z7G6jTJiaMfRSRz1VJpskaRKIOJjn
ss38z+X8IN3bcE66bwLZ/FgEI0ynYT7ccIr28B/KvV56c5V7zsMsEpCgakznZXWD
yl2gNGgnXeGlDWLE10GQZvpHNLzlSFKnc5c2xcekdc6stwsMLE5opv5iWqKvtNdf
FHSAgkLpkOdRcSL8MANHjt44pkzQd0WD8l/+tx4m0KXluLN8MtKqRo8rlS8alM/1
qFojSpwb9WHbvntSBxmKTLC5YonJifFOxSog2uiB7cCWBFaweGLOiL326pXUTof/
2D57EmQUnNp+TYd8ytrvCDR9Eg0vSBZ72wFMzNh7h7D4l3hI4tNwXB0vyHUIa+xe
Uqx5AHeyw2ZOuR/BXInUjfypB3aPf6Su0W9Nb7vRq27ENxj5ldHQv6f4GfRzhTBd
BlyHlxSjTLXnfHtCqu+TyIwXMD+QM5lw6aNuCtfgyuPf1sKldhVUajT2hxV30d5q
CIO7NqoGnGbyNTbmy740dl5UxTDpbMExlxpXNePffGRHdeNTwcZFKEFaJMRYNfmZ
DgCEEssR4RkvaBRjolhfudYpo96cDN3DIXTHl1B3d/YkTPb+2aGJlv0RXYAj7lKu
NHUmPcgyarHi1+/6Cmd0wOTQrS574BQnLwh3ggpMrLzIwQtjUB5x5rA3Qdj6EaYJ
CZiGRtCbpamaai5zCgKQ4ugz3rmv6bJfg5GBoBe9fDJkb9iSS+ITO2OcOEcbv/V2
0JA77cGEL1XcI6PgAX5eQBG5GzLV8E5tt7235xMEjylsAwXOFyv1zEY09wLsrq9O
IXlgg8fYGNqwDyQryMjW7ZZpRpHMHUNNW8C9TmdYa3wB9vHEfqXycgdSQ8ANTAtY
pxJ6/ZXrTUANjs3ktycK06v4ofhYsWfymcZd+H5EUiOnUDpPGamCpydFwzeLir5t
zW+tFTfmns9hadjPIbzYlUrx5MCIQ6T6yQn1MR+HDOAsmMgt/A4xui/J8Akakrxc
s7xykRTFubUARgYsn0eszl8GaqGhM3/IgjBty3QPKdvKd9MAvsIsEdL1do0+AFn3
8YjfMF3mXSQpXTopUeND9i4oQ/sMlsbx3MIdkM7ULDdsG1J9e+NUOwMUh0jLPpps
1buThFFKD45OznGy1BMDdYLSgXOtcYrJpGsfSsWh8XtISI9BOC7tKptk078LznrK
c2Ey4RmRJaRndwk6S/K4sVFRQZCW/dmGx5gVUPm/4iKQNsqlbMrXmgL25rU3eXD4
TQGVgYA05CrH0vIZsEGsrRShZk8iGhmNYRwMydXwRq1Br2ChvUSRjs5syrrsONhU
qparId8vJSm89zpiMM/O+qy51Ma9gbrIWzES6FLSYMF2t2jP4z4Vt99poUnkm3iN
BS1Ha8M3CZjJzpdSvWiGigdcrqeVp2ql3eXYHlW+VhgK3kvdokr1/3Ncr4D4vCTA
7YvskdXqpzXJTFcPJpK8a19TbbaMgo9Dxb2kFmCgEnohFKGuib2KqaAulafrIYT9
RrsC8oa6/XmfS7jtHZAY9vVcEfrpV8JkMI6P76f8uNN12ddahHQRlBJCBOr8Wj0W
+Wl+mWgXyTkl1IE51AbtGqdhDfelUMSXQAG1y/aRsuwYNGPnEykSNwWoiO1znYUb
GLasOinFdjvN8TNe/IL6//4GwSFGwuw8O1b49wd9wyepfO6iM/8YVcx3acK8R+wX
jC0kBmUMkXnNfNzDTJCjxWqR1Mf2LavA3yHmMeBzbj0O5s4ivISI+nNq2GGxBAXO
HlkVIcVbnc7R7x5EUfxQv9d0IYj+r+1pt9tx7vy3pw5CC9eRUce5fAUpNsnHk8nr
CgXQigPQMy9s5lScQof3DV5m5CW8MIazKtmxaH3Cn9yZ1tmrnIpcDVOcnea/L9hT
hAXQoY57gpThhXuXiQsC1QqE+54v0L1t3wPQ8JkcgFpwnJ+uiq9gjCfBelI9GsDM
4RhF7x50IVOQYq6x+fx/Ume92PL1iUNCEi7GE3dUsOx4vDXwqLVWKzKtKOVLwL7e
f3SCjLrv9ro7YXv5m4zKTnRS4FyeqfeqV7XM1ZZtwkXpsX+HeVKT2ZR1ne7uCFk1
h5JVNeLqsqOhTIPH8AFNRF3THQl8mHenNDQMnPFPCrZV/utNwOCUMC4mFxQUlRmU
2KhbjxDbDLrSetAiQa7dTw7X/AwAh9wIXT4XYcn+S3CzjvciivK1fRKqf0PVdPDT
SYx+aBTiK5FROqyvVPaMLpuDCh42pny0AJ5wnyJlO0q+rJlNXgf6ScfVBYEr7H4O
gFb/Gv0hNfhpeE8ggPk7iQMMxYnALIY6uI6sthCFBg51amZCQUoJgrWP102tcPK8
uKcSJwwKhbd2sr6oFa8d3ftTosCkS7exOiDJ1LeZkBvlfJ7IaH4ErAobWCA2uLp/
bgCSOIE2iZICS4V6IxR/+jzB9FUo8yrFufCG4am4Jjwt01/KMpg4jeEwp7E9uL/x
kq71o3ueGMZTH9JBd8Rd5/glbk/NJrZiGUh5mxJkouLmBxXpOZNMemJ2Ath79D86
QU2YqeZOCdItR+mcCF3Bx1zGsSGKIPjDJE4BtSmMlcJuittqhdETNM26swKgE80G
HR4l3HUva/5BUFFy+SN0QRfTAIBQL8NvSe61FpwHXKsMx6K3wL15cMJizfzMI4Ee
3KPB4TUpBzl0i3igCMLM3vquwiNNQS+xYBFDMMlZMuos27Q7xndWUKpnXCd06bgk
TFGe47gHBcUyHFa7lSE3CgdRtXZEtparzveisQTnkCaAHKivKsldMJoeqrHn6YTz
gE9OiMn2f9sXycjU97PHpgfJulECmR4bFiseUOgUsGL633y9WAcMsJgtdF0A6Yfo
pHEXHRMUMqOzUbo7vkCkTI0w+IPNBvCUhbxINeMt3qTfYSv5gxHrKiYmQPDNjczI
DaIumVhpx1e5jmjpZLFhJtf0K2yb02Pb4MqpQEzhULszywymTgXcG7p+HCy72AZw
13mDqsmuSoY//Fn8Wq4KdpD5OTXV5o2rET1BNH+BBHG+OkvvUskyyvHh673z1x1b
XIwUX2fDBgjAGZ73pRh8jiVrTKHEBpBdiR+GMlY6F+Iy9s96pT3Pp5V1BA44RpV2
wPzdr3LervPV/aJWa8jp5Pq/iBr3Y9SZEKFY8yz/5l58r/4o7Gc57ZPyY603R778
j9YMTA6asOkGhhE5IdfRI834FAiFXh3ObI2wfIquRbFtkZiLzD9ow8P4akoTIlL5
LAd8YSOIZE4Y5N8fCJquCcIqkvagqP6RrtDsODPwSag6JxwuUPW6Yd1y8BgfhrHl
76u9pc3xBCYG+cwmMCqH73nXXZOY8cdo73ZDft51COLtLLKnoALhSoOwWy/O4thh
JMXcescffJT9feOvpev6DJBC2Um/HI1f9t6WfAuZEMn+UMtxXHLs4RZO2FczitZY
MfjhGv4ctRbFwO6pYSZlLti01LDyr0hj1lZOCra3ttSyDFPyuvQ+8bmg/QUpiDks
Pbj8PJvBOpfvDB98wa94vGqH/+Hw56lNW1bGZgL0W3lvvnVv+mkHEm0lqiiCD0Rv
sFqSkvv6Io6smVznfjMGXSWtLJKjOzI36aJgSFadnJ6gCRzk1o25VFVIiMiXbgTr
HwPa0rQEkiI5HetH51D9QtVWdI46GtFH5AnkcZSgXRWN+h3+rzK8hFbaa2K+gtEn
V/4SHSYE0wSt7bf1ozv3whvwJpj6dF2ckwibNBKfVT2vRKyDVUDrlVCmxxFFCu74
oQjQwdo4Fp8Z62JJ/rucFOilh5ld1VvPOPLwmyRKmKrcGMI1q5UHyrRVO9RnjS2z
UshoTX/8WOCuOnUzA9O8x+YNBI8QLv+/ieNmDTo3C+EkXYFhvvV3WqiIwieqKVzk
2ZA2KEAKASMsvqsHyL9O8l6XgMtzfHM42N+b7xXzhE2pilM9Qj0izMD8y9PFYw5h
6du6LlCRmQZSL3KXGGIlRFyFskIvy6BJc4OK36Z+iszcXrFUUmyk8rmy/UA0FNGE
7Q7eEIRig/abUxVD/Zt7B+KBagLdS9+/os+ZjaLYUSH1BL9TbkfXNbd9B3eggCng
MwGveppg56+Bmr2J6T0TkS1UDTag6PhET/+ljSW1uQ+KJ/Lxt5J1vHmPn5gRsEuh
OBvujgdg6Rpo5RqpQurHkgBRbU/Yz35/WDhBTtSuABu/O1hVdzeQ7TaSxC4gsh2G
9EsmGBejji0xeBVdnb5JwVPfKI1vDgGhRY/OCM/2vP+4S0yjrqTasBWyE52wfP/W
ATbcaX+pLoKObtmL3uXx5GVG3H+IV6rJNvR8FhqS16HkmGB7noMqMDvOEbIlhSQi
EYTos9+LwD14f9CWp6wCRqA5uWxcsiVGamkTldgSWLyokjU78f1MIL6wp3w+3YGc
7e9ffffpz39qCP6C9DLQAlrawdv/FS6RQoElWcnFvIzJVW6x8NRhmCtaVTBHQqcu
q76qlb7DAu1ah3RYwBWvqlGvteKR4Mq/jkNyQqGFzI0VceN/SXOajsPAlthq23BU
nl7jzNJkTlsl2VQSyoL+LGtdCwkOxxPTf+/hhHCxmFMGLh2MKxBCOxroEyhLlSTt
mdtPIMAOANXpcLo5qwEitRDEm2mKM9sBhxzWNfWkUNT5hFcnnxcJiGe6FpF0SqV5
kW2yLcIIcQYd0qvQVbuNLldEDR3/6ttDsKppqYAhUV3TMj0/m26df7jlwnw6XXKx
Th4v6zOi6zs9CUYnI1NDBbxqKevS76LHMH8mxZ7tJkmrw4btATqNx7L/75URg/1r
L4E+us7349M76542OBI5la0g9s+DMAZsZ6jhRkpSGQqMtJSSGkZzDCxssw/hTz5u
jcBIKJNOXGMcdTG8N5rN+9IDMudlmZIa88uDDNP+HRmnd+zmonyfsVXUilUyMvH0
W2YiqXYG6wI+HCK1RAj2VmTKnzkM5ae1bjDJPbtyrHejXKzghXCfNp8+NlMPrWEM
DY+c4KwxSBkSfk1pKM7XJae1R4pvk1160FGl6UUgyz+JCasTYsOnAr3fCN5CN1zE
0VsiemeSO3kxt6+mAkmIvtqmQsTN3YHAwOa3RLEy6Sx/E0FW29mHjAE5LgBTIWoD
aMYXluHcYPQeN9kMQzSJmjgmYqJVjM2e0FR9UcHhwEwUkVQjsWb0SNRYej+zfNPg
k7ZRrNNJ8I8ZG0xljYYS0CZa/9Fx1jegXdcgs7oNl/gbO0ClCqywlocf0g+094lx
qQUhK8J/IClP+0KWbwF9BvALyr8wYabk2iKLY/MdzSKgZ9Jr3H+/smwSOQOnCZJz
psngZriNU9bVaULjBDphIWPfyn/2PdI6L7HTLJk4OuN9Zd5IIeG0y5YsTod03LCB
KTYw+GgWtsQfjjQS0Q3tSJ/DuwQAX1+TzByXajsDsWFpIARmSvQvKQNbzIJzhK8F
6phoev5Dc0+6kwe3Ud0N6fyGiIzz7yZqIedu5sVPW5y5gvrCGZk04uWbba4EnmUE
QtmCTb0p97V5fDA3Xm2HjHeo8nISXraCce+F9E9URZ4BmV9woBWmcLBedHGTSqEJ
i/apZ+dSs3TNjXsAPUu8wW7gZuHn6F6Te5jS7Av51txDsb0GOHfJ8xtrImFbDRbW
zG752abt4cWbp5efuBKOAvni/piy3NKA7WGybOxULPondccuo+GefPh8FP7H4Uci
pn6wA8P+U7inN2LDArBMrHT8VYsqa8Mw+J50aiZOQG8Wv3rBN/H1YbS/izSVNrf3
MgorthxGHdnf7OA5m15i2Pw61ff+TfLhkFDLwsA4aiUm4ZywFX+2g8ZEDM4p0zu9
tn0R6C+RgB+Pi9tO74vxituCg9SX4uSo0YUIKvKsFFWE2Y2OhqT2hDHPoxW3om+X
a+lipfUcxi6eRR5NOfs3Wa6BcSDm3UNqkX9VBX/6bQ2sYe4tKDd6UzEJpdudHVv7
fHPv9lxN0Ihc/FDxRUu4A7shZoRmmdRard5Dw+dWND2HjSUQxF5o0WfjzAOdkZSN
vjQvpFplSCnXRJNi0qtvYMNDE74/Kbcb2Blb2rnQ29tttTOqdZtWxr1K/+zq/PnG
1cA9OSNw44wm8kLWX8VpJhZeMiJztbi+K+7pD5kRAt1Fa0nZbQ2qELcOY7eYqzky
VB6JVmj+rwY6yV6zWAStgzO3iSUpmWBfK8pQPriLwiI1tLhIzQESKxF5HTcxc+bm
hQXtS8QlMLjUeDokPlVUH3ZswXoqrnFpuqam8jRyoS52Ehrhl0uE4lv86lcn+DDE
BRlAKPzdkKlieUaW+a3zuZDl9XozitEgqBeirO3qRIMc5LFpjXCwcL9IwItPuXK2
7eqkEbqsI69IyOC8FnFTnwIAKOj32nEyHg1s7L8KtT9VVIlQIhcCGYRRURU5D9ZY
mPrDZLBEH1EYVg2bDYa5TR6Hosvcm2S2cuQCONPQUZu46Sb038nfty205VlFiOnJ
NNyvijB/J4r9aTYcbIZioXKUYGh3hLPUaUUJN21cddiFgkGRDoGz65Cau43R9ceJ
ZRoQDPWc8ZyEvh1PmBeZve21BcqxW4yFOIXzlD4kqa04Fz8gAAOVptxTy1jvYs4g
ui2BgBY1ltUAb78mZYf0mMN6NbAoFFWuBqDv07T5Jcy7eYR8jGv0h6zOf/EODkqR
r7avJD5qIlDffmb0aN+SxbG/5uTAhJmlvNN0N3p2hfezCGtGQTvP4FrDTiLDO1Jf
y69B/bgdErBZjtwd0vVW/nIPtyHFj6FvXtxaXy+FAH1YhTBc1Kyu+HIv320cpvFk
iB5pTQ3WIAohzSQvrndtQ2y8MxGo7yKCQ6keE1vWUS/sLHR3mp8sT/g0J0kXoEC4
ywQHx57022YnFPeGWULxGedGEWfIe/y3uSsTU+aDNabbVHVYqW0TKF2Y+hx/doSV
VTMhixAMHBsKzxg7d4W2v1j9FLnwKIYC9a3e715j9kOnrE2FAZnz3QanK1PERLoR
dXKpTGoO/FeBUmtOU0bHuTw3gA3Wkv5Gr6+AliCW7q9z+ByhRF1spvjJxzltBd2H
4uUM6Jfl1HzwatfZLQ0wh9rZezYtgqQxMJ1PDVgYKLb5S9SZFq9RYObgeAdQZlEc
Eq+GExY7B8tTzQQYcEy2CDoDnvv0lh5JOZFiQdm/wLAXj5WSsizgdR7vBuLNW/hl
75/5zSC4/yXiuB66n1fSr1mkInXbeOwVxhdQtKx+mdzUcTtxSdus2oMq3yuho8Ma
ZtQQguenlKEq4zInz8sPhzfnP7dY2rZpnprz5ELdiqg8NXBihtKW61sa6DIzflQh
0/eS2atlPxSnGLtk0xHhPOeIXSvcAFg3MZu7Ef3Eguf0gtyZMAWj9ug6yirTwlq7
sdYHMQf0HoZM8aGO9jLDTh7zvPVRmbpQIjiUd4IIiRLv/wWR7dqTNNZT4era0K5Q
VPXxmgo/qkoy4AvbKREnQPa0jg/KtB519aKutuvTZGIZ9ko4X1AN7qvbey9zl07B
HwmZkoqb7v8meZw+2rnwHMFjAT6bJW/t3Rd4DOha3Mc08XY+btJ9u01WhAdRm4wt
nREAU/Gh4pLqYYOePrzr6skLPBUs+zHhabrjIhZNK1rgadXhhFbmoTkTGLkaRraX
dCSD+opL3fWiCY2zP5IXmNsIQF48Y8/Fh9bDXdzteaRtH80HqhzRvdD7SBBcJaJs
+oNAH3QVVpqsFWvnKp8E8cnOkm1XTCdEP675457yPzJo3Av2BlSkvfVHOcjPbrDB
paHFU8sv+c7CpRyyVNpQNuPN9nOLEIRX2wpU07WdAtqR5F4CYmXu41wSwmF9SqBN
3NjHpo/tLp57UEnl71rEux+BjQURUzXD5wvm1hfRJMlklKuCXKk66xTAV20L4K7K
G6akuc0AOgLPHESpJscxq89g6YyUsdN2SI+r6pcRCfSeuWizbOg7YL5mUnrk4UsW
nBmgAG0kzwKz44Ju5Qe2YVKpOZdEKUkbEo5Y0YmZ7um79a3Rqm9LPbVJMiS7DsfH
fUgdmC+VFDT40nJIlM7nYsZHCsx6PLz/EpQEG312YA22RbCG+S6btv1gJgTYWwWy
XeuVMVaBEJLCGBzdYeYRcGrTdh/0m1I9AL2z2kao77jhLutCTFHmAXPN4hh4eu5D
dE4+cn+nkTSh7UnssKXXyvy7NWt5nc0rHLO8vDWdYk9d4yekeYFCJ//1Ax/IDRGt
k4BvdnKmLJ0IRLMWzPtfIarYXnsDanJOKxPXTJYZksuuO3kKf963gevGArhjr3zM
AOoeest0u6Xbkdm+0JsyBBI6FG4/sM/yvbAwzfdeA7fscXdgI9QywDoOtcu4g4wP
zGPrx8sCiErXd/Bwe4m+OCOu7xTn1/i1dq0B5VZP7lqeRwAy8WlR0vPQosMmcwNs
v4nAw247YERf1a4s0v8S81voF/GymcsMDHndsodYHV7k6lD30RenGArOhLVN/ejz
Oo2MsYj1zzkjVaxHjF+FQ5akcMWT3e9hagbry+esvmeUVDikxOSdrdsf/tPuKWaw
DMWffbgzdFY54MgS1g7EYpALqMyOD0Gk9jp2v8xzROtQ0GdwA+F/w2Sfcw/4EK+b
lhBHKaj/Kc6pw96B8Tlc9i9ZXI+RWf4mONujH4QruQvsfl1UznVjuPfiPykiYpnB
ie2YJiohp2AQLcWT3aVweigIIGyluXTQFQUxweV0w3rhbA5XpzPT8MuKHExp4t/z
KPfQy/SZWQ9yYVYT2Pxb2xHmLWljNcxgHtFtMWU0ShwiFOLX6mfctOTlM+pD+9/O
twdbTbXs/6YfMJkDxTkErJspC6Vx2uqiosz9abR0tVtjQ4/4fgR6czcR4ex4tGbb
TVixF2q9ANevwQMvPAwCWKovLh+fAxfHWLJbs/H702PDidPNB5ZO3dxmpxZIWsJr
nmNRhJjN2mUOBNZO2VJmR/vbvSU4l8+N3k9a94/Ay911U9FXMdPZcgnHCtfs9LAx
Sk97HtZ8u2cRduex0kOV/Me1r3Js7q6AtDTZv+nYcfFaNH5ppf3+LC1TWtGEaEZ6
wPp1TLcGAbUoEe9uVvCqAv7WnijS6bvlXuQwJSBjMwWvwbChsfVJ2ekwr03UJWdv
eMitT1IjiAokWlVnxbsgDo+EtE0KQKmUZXNdGYIiz7DvZoy37de4y0fMyMlDh3LJ
+tTqa0ubeUTflZ0uothEvbxEA/xusYBrlBVltqH8XRSjtb+UwghqI5UbXRfkgh62
9nPV027dnrUG4KWuqcqY1JF2MVRx652ekrIQ11vxu8Cxa4SDTBrznjMo9h+X5rmk
STryqx3MwHELW0rlvjrr2l07R6g8rXyRf1LvxOYM4P8Z6Z1yv2++3BzWw50orC3i
f8paNZjRVlvDrUxdDihY4hcju4MAlSfZ3TV+UmwYLwhznLAYhujel/4amIO/0W+c
v/05Gn3/MdinduIoZremSTxGWsM0GaYEZaYFb3JaO14sr4v3vHrL32L+8B8Qb9R4
2qMizaChnC1TH9GcwBRy0P+bIWkC4Welx0XU8s8/LQoW1x92hUX2AM7kw5IAFNMQ
bZZYU9yB9kKqWUs/ZLGQ+LgiWbgo1RjifNRK8IAMb27XLtcNcBG2YBoDFf8BYjqz
iNiVML+nV9A0zHiTU34MZQHj+apsyHtEbryNc3jUDvsscRAFLMWpGWBj2rA7+dGQ
LWBtTKAbyuRQc+KMEHimSOxqEA6PxiPqYPoCyV8mj+SCEy5ny2Y38GUPXPMGO0DV
t5jhpwDXT2Xxkev3ewxZbWu+h1NmBcVyAq/KnI5pb8RQDZ+aQYAsamsmZKPp7jhO
Uz9sTyDzJZrC76HINNzMmj6BuUnHDdef8RnRfSM7Xhj21Ba2NDuMHMH8quvNI8Nv
V75ifEdTeVoIwhTfH3M/wGiv7addmzGa5LwoxMyWuat8sRQMemIKwQBnVwHViyne
Use7OKSXrbZfFoUEaApz8ykeqY2oF91I6BhwEAkE/CZyOMWlo6E49cNu+vJYyc0s
9fpO/FvVvmQ/UsP2UYbsCNnJgY36VThNMd7Qnpdlbjlx5zn1DUnmfGCWTnlNPpcT
T+ZPNbfEPvkRBf8ruJcMjBpwgwlMLdPLsD83+YksSRj05NQ7t2I1brcXwWX6YU6d
YooiYXK/SmeNCAVO5j9loPEz803SVtFshSFzG+QULTtVb58abJ+bcsDUhMDWz2od
mJstIpUfpy8S78PA5oh/hD9nvXPgv9AYVv+biARcjz6YQ2ZoeWDPQg0G56xsjczs
muHUpJrwiPty9gGzQ9ZDbwwNpb9aGjxGVF4qgsMPldKbF5yK0HdYswJnk4N5pBYl
QnUj1wPZHzAyUQgSeYZIv5T8hxoD7XDU7/UyFH35YwYi5fP1JlFa91Fl9heIvx1c
G5rHZctb8M45/N8aI+wcx7Q3wReIE+Y9BW8rfa/LfqegQ47XxjbtD+qwPRgiZ98Y
liuILqHpYZxwQxhLRFQjqqdEhcjgBuLil9Gsdz2Wun1/I66/+PWoS8Kof4cEaY1T
cwZbaZ2lRGmVSAL5fesHKavctuvW+MS6rGq8Pz8Am9t569+oxx1J2PmBsezaRIte
901tb3zs92mm00tGZ5WhDweCvlQchRXh91fr6sEnLdlgATJ6rEz260iktFxYVq8a
StN2M4TDfziTmubTpVgN41XGGN4lU+2oB9zZLrKWW+gFlbzErAsQ3tRddjRKe14+
eCoirbvdqz38Zyx2OcObyDoGBE1vqhSvhseWf1Fg1QU4l2TvcOfBvF0O153KJBYN
FSNz1nW2zTzjGuZAH1afhB87UF1mSAR1gEbIuKZWX8saFy+jl2pFEkBglN9YTqpW
PiJ4kpukC8sldr1iuJ0k7bf8GR04Kvqmy0UnWmjQfcHbc2HKZLL63ZS2ppELLbnj
QMnKHL2IYSfKVFgGM67+kDV0NljZ5Jijj4WNR7WbpfRxVLDaXkyCUV36avcaxAF5
P000QKNPJGJAlBddXPfEEzuxaFyZw5TqGtVSD63gNMRR5TPuNI1Y/kfa/ZerXy54
SSHpSsvK8y6uQ+UXN575eC0ouTGEPxgeBHNGRgR3v6xGbIqMIpkXeARYwVh/SfmU
YzvSMpR3ix/GOJPxl2VgD0lxd/JWnMnxBw7mUNrkoZQi+E7zj9LM4jb2YF39QKb5
k9UwqYcS3dnCtDXFfwVtN2aiJU8CZcjTdc8/mtYHYdFmizmZukLOdTAQ9hO4jvro
dYMWrlBLyFkCKUixOYsCZVZbxsvjN44Yw10RKux+n8eZBwyWWYHygBv7Lglranil
3MGcCAoCe//odQ1oPhjYhZcspnpx5D4joI/3UCKqeutE48cL5iS6IHBGINhcwkqv
Osa6ey9fgCu+HSKfHrgFt0vKKA852R0OB7A9CRRNuPvpCgqdy46iGnx7XN6udA4s
gAeO/Mc/EJW6ae9FDh0W6ajCG12cUdtz1YIgFWl83pqIdOxMXWqzOt2fU5L9cshM
IEDoZFLNJJpazVGNduWBMYH9mdgj9o2aCgdwahwcACFq0M45XCGlB3dc4WEj1QMt
OCYKyFagDGjFD3nhY8U+scJghDJMz4uMROSSA822EHp0JB9lq9Wl/8tSxVRlhywc
fmJcM/UxjmVI229gPi2sW2MMA8rxYnjBXO87wchnLNsYxx39uDN8wE5+bL6tVh9J
VtX3u3Vr6MdMfDjpTVf52Pqaum9U8mkokOYqhdWgIa1ZqVReq6YcM2pUVh7AKwLg
TOueRFTykn8Vu/mDzIXnzjkmXtfJ6lSigZP6QJxxRdpNn4HXw37n6dzXJn+IyKr1
5+msm5gDbK9dY5jT8EON/5kwTD2PSkIyJKbq8jHxg8wJIv59I59CGHx7sWGT3Jo8
APVw0FKPIl++0mNydSMDEILEeMtBJbLIMJzFv+n0WyizTixkkXiZ6owAzAhvzm8C
QPqRPSkmflH4VjJTyZ3zxk9pOrKzhttXeqQ91GejSGuMYrNRMK3hXzXV5ceKRrKS
n3N2/2+2knc2YGfgEehEPuCV8VeRvo9ZR5PQQxRhBJhAl0aHSHxos8Vp35W9J1cg
1NsE26U8gyUjCEDoqRc8NBUQqiLAvfGkiGgJvLkamFpfHo3xgGnpNfa1kYE5ABZ7
piUmzT1lxnW49AVP7/U5Z7RNn/GP3d049B3VC1w8eBdgL6V/Ki4QeAAIGbpN8yHD
nSNA71uqZ8dYak6f6ngVp963+jUM4ELzH+yRT2TqisRYC/xG/NWmclGpd2XyshAL
Wuny9ni3xHOQK1P5lenBAzNHzfzcoTwuBp2m6pRJra/6sc5E0k7zTRGm3oYgO4FB
MKADmGzgSdsnd8XihO4d3QjY27vt2PmYaMN+mnrrrh6zyyoKhV0gj4fl3YHhe7ki
H5IpbQkJhTtObQ3EcuA3nUpbQLuKOu1ivrZzOuQtl6wOnsKRc6jhfoLdiLCpbo49
LZaal3TC/YoHY3gRg3hrD3alYsAe6izPPyY0qWiypYBY4+ncNOJZBmcGHPgBTG3Y
WBcwq+MGAng+oGjRkBPjz53YQO/V2W6Zo0VacpCtkKkuH1yyP4OWa1r83yFE8phT
H6LiaUUzHJKGEE7W0w1pdGA5hg+nIIwV7qf2JyAcTGyLJTcfY/IGs9lTRMfov8/H
2ZXvfRnq4xorenB2PMkRUTdPY/KTZYuj5IHaRgq6cJoj7zu5yAWk68Q772h03QRi
g3keasFKk/2Dx8ir92JQ0nrj3cZlhIe47r2hrKx6KrLznzoOsj5ykW3NDMWzHP12
+I4fiF5UEr7Ku9TJ/CJnhxyW7W5Z3aUmsR4tEjC/uNGRPBlErt5+pg8so4ynlfYZ
sZU1/EkHMTodp1krOdKTphn1zWd1VFRX8Wn45cEKYn9CKiy7wxB6cnZwNEBPS0Hm
MX6ZhtuWVbmcNzNYA4c5+uvRDx+yWh0fA7GjZZuQqHIGTTePJUie9q1bh52VRnC9
4WfgCXHSvVJIKZpeY12GX9qs3CBHYbc0fC2a8JNf6c55F+CiTIvWA86k5BKzg0zA
xp5JVmcF/0rB5tgdFHAc2lm+i3RHnCqQIptaixXmw0wbWYAhPChnxTzzMl1vwqnF
XaO5LQhshPq2caBUa+I7qtPOkw4l40HWIUzU4+6hr74CsbY9sKjdzigUVrYTK0g2
WViihqgSHcJO+FIX9o4cqcgh8tOMVuXXWo9L0rSJPkSnI8W28EffoaVLYZVWbR0d
6XvtfDNWnbJMnqygEsQunzn8r0IKenw1S49C6M1+qlT+SKVfWydFdBu7qkeguO7e
xMGAsOz6lCML92+QWT9x/hKMBEQF3MP7Onr2v1syER7HSGXJmxkmhMrAm9vDRnaW
qca9l2rLsUisJaRqZr/ISKavsmeVtuxoy1zvD0RG6cx5zX5zf5BlGk17p7AhmbvS
1Hyr4QYw8Nefjmv3CBPghFqPP8gm4aqX140SVyfwfinsab4998y+LF/bCtsbQMNp
PNIxnje7K6ZB9x+AFbwX24Xm6xIAseRbhbnMbhST0EbzGE+ZBNwcTEy2gH7c7Uag
sxBcMuk9f27QOclslZVU/5oTVT6Dg2XmWKX0N4rEAP1CAbpFsEuEKdUaeBTiqkEy
vfHruqacw0Dpd7TmqN4ONCCF2QJ3KZeeeDWr8sq/rmp3crqCEAf+EjYVoaVSVhGi
v0exiCVqokIPFDdUPKjmG9cBj1adBVU//Ks5Xliaqc0ML5+Oii0I0A69yoXEZTw4
FnuDSalupVKHJ4/I74TGZWQesEw/S1wCbhvaYJvh/BMnf0u0gt9VnJFExPZKk5pz
sqhdwzwxiuL1h71rn/VkXzHVsOEwNltWgnx8bCOm6KxCX0NEFRLpd5TpuYrv/Rjk
4gky4s85a4UHb9AqIdPA4mCkgMC8i8/UhK7D4jBXBNLmnlHEltIqP44PsjJEX8Ei
4YeJu9fKC8EAlbDMvrRAWu4XBuehN0L2K0pFNz/Q0Iu6hV5p73y28TTt1YgYA4BD
CFRwWSFVdKTvlGYBusXHfgO5q+R+yWb1WdwsnWHcQUQu8i3qx3KLfjUQQJKE6aqT
kKuXRmkhVDvR7jYWw4jXGIi5srBR0gXot9eaH1+TI5yVbJRj0oiEY7/p2lYunYNk
qM2KITxNRQ2P9rWpZGAX3fmOt9kDtnMRjy7y4YL6pMPAztE4g4BGXocW5ElXdKL3
nzI0sTFBIUruPGV/xujqCMpvUHI6EoReIbXyPIZHur/bNGeeYGUOgP9TlrECuAxV
YBtLu/zZrrFf6to/vFTvvfI5P8ZUMW+1JXiuXqDCqU/SOOCRt+d+mb2rww+YTFXy
iINOvBX8rDU2nAF/w4IcIHbsc0piBbGrR5RwOPiFuJCSALhjaWkVyj08vat0wDDP
/ZUIyXZ31DKmmcNC7VyZ8aym2xmaS2rBkolotEpBCxp4syOt1UwQ2fs5rFD+eXhW
7YtVkkr5zeNc1HZKm4I63af8Bb8hVxpcC2h69q4dOKOd+jfW3SM0DG4GMlyikUN3
S1g5ldEYIxXwJR+nKBChFqv0izlKVN+Tcv2drlSUtiUvzJWOC8sKVz44f1DuGxDJ
cKEzh8fmUF5Zo+ZxPzdx0/Y8VABv8fEpwCJqIfoAk1w5kqgdkNEFCSLUC2cy7gTk
6tkgUZmDrdSzkZMqozmXaHTB2m1mMfKpya3qjib6YaselBEeS138i32s5mHfa9Ma
oMbeQqcnTGvLhK5ZU3RP1FTGZizjVMpY3wxLtO+0CRbxe7VkalC4owAwXFPlYn7O
q88LhrVAw39slSVZn6oOBJOMUYuI/mkS8f63oTGzdnbEb+6Yqa5Lek05abSKDUNm
AqNW7FKeY92yw3iCKR+nJYNAkzibyQav0coGlyuTS/SLlqegU2lwjO78SbelDuRf
3DPMdMweXrQhMGFA5rm2ERSLiWKFKzaoG/6jIC7DmpTdwl/dH1wWP7ASkYpjDRXZ
UrZ1LCbHkc/UuHZZ3n8QogxNfaCCVrV/XaU3Yz2ByE+uIqV6A6bbY/ZeqGXHG5M4
C8U1yJ2KPHggJ/5dOWp6X2CKpbH9UENx+2WnRrekPcvuJgDQ/0JHZNzfbLY0nszJ
xAxj5X1zGZaC01eWHRt4pdQMEi0yWAEGHZCs1HCOv4razszIaIXBSWZiP4dum7ap
iPL6HLob0O2b7i21umM4HExfXMnSuBgMRgniuT4R6MuR+IqR/DP0T56b5E+P/GZ2
TVbQxwC/cUWMzGGrlnT2ibVz6OMMpdcp5ScpPx5/p/0gRtpst5LYPTE2we/9+BBJ
2G6OSqMQanSCVh0P1TdkPMHtp4dxn7Uc9S63Bw+xb9pNXWkBhxzfMlr8uG20C4pk
Gw4o/Rc7PJ8Wfuxg0im9iqpB/cs3rTm0CACAI8PbJsc4p/rs67O48/vZkzjtOy4l
nbp0AjPooKhIl7zpIy1A8eml1hKbLWTMU/dCrp0TiLvoBfQlOQT829fa7ls1fNZd
tM9qrmz+Jxo7dhLf3mbpXAKyEpUjhT9TaWq7nqD/mlgln+Utt8dr07z9NpljCdHZ
VPO1QmPe/ExrjVx4zZF7UtzlF5XK5xcb2U/GAFmL3Itg/Sm+ej2dZLkV+APvf3UZ
x4DdXvmVsDYLJFknVvHSBgmHniF4ICcj93myZXoEsuyEuikIhFLWCPx/ZesCCY4H
Wjt/KGWD2dGndSskzU/kZkLT+37rrvhiWbmCX+g7yGbdyIkmCN7UtKeuwGM/RA03
CeB7fQ7Bx/dDMJSNo2Vkl+6IdULhbTyiurEga/is5p/BQv2/ZCmfImnKPR8T0Q0+
yIMPGTc6Fi9IZCvq3eaTKk0I8OsjmLVRa5nfT2ukkRYrAeSWD4wwdhOMroaE84A7
h97+VAUvLyt31LhQHk3WI8LSH/GlAejdF6v5gxQC5tSMOU8p/NfCj2g6S+9n3OJv
mC4a6M5TZ2IDMNGKl9uEExU97Z0o/jOJH7WnSoal/ZDgHAzyV9GUPu3bmbj/Xsgw
dlrJQKE2ENCm0IfcnFwNLksL2tLmBEN/zuIxx4KicyMqR8uoWjnqBPoQrdPoP3Ms
jY2byLqamp1zrHTCwYPmGL42SjrTlCsVe3x0r6ys4zYNS3+TfMN1xyFYgI9lVROC
xC+wyNxuSeFF0C0OcDRsrw1mkSD2ifZcaYsS1omwzKm5U/RFP/2SMdLFXKj4/Gyr
2KN/hdkgJ6RySIhBNk3uTDPjF1xNzIbNfeYozjfcuv4r0EiezIafs1KuOU8ttggm
PbkwCbKuZm7+JPzMlRcV+sbC+KFgiNAiAlhiqYeHciypvby8JYlCGM4pbQdln8pY
z/I1RF08Xgoo3oT9XrQzQPSFEnE7+MOKF70FoATr1tE1SYIr46OsX+WVmOsrszwX
Yoc8RdRGQjfPoKfoV8dQPB4CdP4CIXOBVDJ1/KXKyNzTShDTDpMVaygLnRndZgPJ
tbbbdBcDx81sm3K+dNZ0JWEM9kPopIYiuUis4z7uJpYHzXgsbS9YfkLQOStePzWh
tJK/FYuFyo4+XuKCFJCqowcvpJa81QlQth3eXy7k+ow7K3hzNqYL1B4Xrs70UY44
lMwAo9brKO6Dj03HTywsOHMoGsflMGB+5WWu/+9C87QbnxMymC+1asWf79tHE2fr
zzScBQhf1KaDDfaxmpcxNpXcMxUoqeuMGDrEvyp3sCDPMEAKcBQ3vO4fnDpxiB8W
R5duhV3Lq7vXqcI2abPmL/9RPyf5SVJjdF6S3JIaj84qhjQDaQtgLopL6gOMNQOx
DMBNlDAXveZdK/WnJEm8Mc/wECEBqN3tT+jgKJhqIQ/16JukXo/3L5zVfciFrpHt
d695iHuip17YEYgea7Z3DA7cNujOXxghuv5RITETLPk66CGls9agYFGe0l3emYpJ
1qpdUEXwVGAYdj6zpplboVGWPOmACtb86o1qwRg74vJMJMNXk+l0ptoI+v2ILz5W
bGe/7mthlnxHtBA+TAybxT+K6COEG8rXr66XNYPjJSzrP7Sd2GVkNFf/oz8pLp9W
kpSbEr41WYIJX8H3XGuZ4uRqZ1mrlF4iB/u3KW1lMy59dDqWQag3mKQ9jWzLAnJy
CzyaZbBCutF7KWtUV62QvyNfHsUlphJj7ecmIh076wD11XRS2JqMByCMPGFPrOuw
XEgC0kjdTKXQFqd+1ZE1k/9CUwrL3aDDHKtg6501CkQQTYLTscFEzl4qovue+wg/
cBeCTgCM3j/Y+zCz0cIYenurMkRK9+kF6aJYhxmK6KCtL8ujIXcq3kMxCIFvRmfF
f5nvUkH3T5eLMKLTV/+gVENMM0Ql2R9Vtn5UmwXUjN/EKjYbHoUhDJoeVNc4geU8
uz2hDt5V2JdqHYl+a5R0OlxuJqKULY5kyKqoQc+RSlxffmAg4t8A40uS3tOC7Gur
mCvu8IhOH5KOy/LMUQERxB8xW2xcg17T9cufpOKKMQDi4XcQvmZBCyNOU8QoeO+9
AncAH5V9xF6wiEGk33U06ESEvhuU0/6MRDnAIIXpcxdbySF8wSLdEoi49DvtirGr
mRP3scafBqnftY1KBY0mK8mOeYxvhMc9JUoyLExFSwSlAfN0VVcIU8kHixr4aWt4
ESDfLtoE2bqj2z09ufjcsTAj6J9bp36uk0UEu0BBwg6brORN5K8YlKLl4vBLYIr9
+SngUFNc7qkkgNsEfzQM/GRwYS/h+7+zkpnNfsWbIOxY8WGJm6qGaCq5lQHigXzl
TP4ywgIqq9wjUEwcmrOe9J4nURl+GgsrSwP88G5RAmbxU9ogFFYEEd5C8JfTsJ07
wDOlO/qIgto9u4x+DdPr512u/adsVEAXInr4TzT9QokWSXi4G6fJURuU66bUrOOu
u3zvf92s4ZOhjGftjAKgAm2UTPrqu6P2uQKwXDQgw2orWSoSrO0rwafv0/NCUaYa
nZsNAVYH00CnP0z8PWwkmn4O93uw0FiXrxo0uTqwZLSEPi7yIrkihy4d7N7INh1G
Eo6KymhmqizaBgRUBs2YhFqQCa+/zXE9Z3f4gJIhjyd/7/l+enEQXhK53KocukRA
95VS+EKJvuzfneB/OlKH5GvyCiscF+M2y+wJhbPGWG4321j6Cb3p5PAT9h3fM/G8
vzeEI25KOs5/20RRhG7vBbi8nf7AWoh8X2DMdubZnlwfEXbQwsaECjOUROUtiITL
M4a6KcY8525DZL6WtMdyc8qOKOLmr7gUs4BR48iWGh/YzWWug+noISFa3/hz/qkV
pI7XFif0AGNgQTcn2GXYtt071wBMaJwNrXGCdsQQV3BEN50qBcMfG5RUq5ygzOkW
Hn52ZAKFILogqmj+Tr0lZ2UGwCVCqWizNaIj/QNgRLrBOI4dqrPoBxRG5sawitqV
UXoVjLueF+idSLvYwO2nVV/4pi5SyBM7iq5O72+joEX8wBkpSFN+uhN/Hk/FhzE1
a+9ZbSijRs9tVaAHoAqtS3JBQIuEtXls8MWRROHNtIdqq6/7kxzHbimqaJghh3Fg
7cgkXp21lDQp4ZDxOLUO9uoSgG9Jj8hQD72MTgPlTPD7ABuBs9nCgu/azD3topGf
4egifPxTqfQOAjZAvo4LFryxAhpQbB117ZdblaGQStUNFMUoFTf5QvWkduGW9ma9
9UUXzR/qBiowDTZcQ7v/P5MkdsTVZRWkOn3iIbppSFnntGUXSRVUvS/C/Qyn+2+H
Gqotj1QWue5gIM+hiRmYd5xD6I2fBZPVGLqVTrVO/Rv3TZNYoM25yLaX7YaouAoh
SGJckDj1v1oW5qJnW7ycnbBL5ULAaMp5TqIPuhAaVJHArAtM6B26siOh1vG1CFyr
O530PGQvRqX7uMqKlraHc0gY2r2Kgz7Y0TSVbCSGpPHttJg1muZ43nJ/95Xz90Yg
GCOQ5BsNa6VGGPL7Vkw4QM/S+bdVvauY3m1nFdCWuteGnVOsHipi+2WidKSixFqv
CKqdknDYCGRSAps72qwKdeAHwE60P5hWAjTpGhlvkTPy1D11ZHNWCrGCsiLYXwyE
hRlBX1wxNU0mYpvp0i5ED3H9gIa0h5MxSAk0C26mASULxesPh5UEtz9mxwl27pDi
tY8j8pr/I9zde81QeSUGoS5A5OHhROvI9jkC7X9+LgZpmxZ0R+mfmPoBIaF/+1VJ
PEZD3rRVPDmvrgNF5KuJCCtA8JIaOdWPh8iLO3H9B8JvnfqI8K/AFRyYIJCLnHVG
9KuEEC7DeaxfLvuGcPujxrTJcp0P24IzHVRJPTAC4sr1+obDszLfEzcWzaL4NrxN
2WMqRBlpJDgyj6DUnU/bVqCV28sdgrdk1o7h2X70BiZKrKzfNWR+egR9185nPCJ8
EdDHtFISHUe/rilO1GW/98lnC1Cyhqjo14yhGZYJ09BgA1AZ4QcUI5y49bPHIvWG
jApB4jbVsic4stqVZWiWftESQXEo8iPBJ01hGf26NbPaGhQjmAD06gysKo0QYKmq
zh+fM85CNMxALq9FjuPDC7LFD3uR3pAOvfpWNv2BDlFflktoySORiYe0wDl/THtw
k5VoDMASkvYT+gWfSXxwglSzlvvCz7uFBShvs+3wa5chdursxZF8Aoo4qnVtk4nU
izZ7NLmFU0A64eK1yKVgJLnrRsbr8rrEYBnpiUQ5YOjpG9U/KnEU9x/cap5nOMxy
7BwugHVj/rT6pizLXGidCHN0zLuxuTjszjXBzrC8Fw53Q3VijrxHXXIAyMADXlzP
+MnxQifBxTV7401IXLeY/tIw8alJCMZ/82xS5ROpsTYBcVz/AUW8EHJ7ii6l5LyQ
oBt2JSLyTdDtkjsy0qTba1Ek/xeRzrPpd0W3Ymop3N2Uk5HowHShaTOmiQgrgo8u
oCWK32szgznDWIC8hCY3cPAFanNhcqf5odZnC05BPqejtJbgImMbj+9YCH6AqCo7
uB6m1BwE8U5dTquuazKu7NwD6dtfBsiYd+oRdfpdsVSmdJBLIXFHMFSrzv+X6gju
HSc+oO9RmmF8z14/huJiBF/s5oUZeymnQG2LL0g8MrFUbQd/2cGcPwO28b2gRxCi
iJFd+WFfrhv4xsKGBma9MxchXM1ExeSIMCSPmdqyuhg2LbAAvi+7YOFV/JcM0uBH
Rgt9g9g0vexNgPuSKl5vp0AWYGMwvlyhbnP6Q+AzhHJP73Y7Y7BFeb8cR2mcu2ay
jRFLg8rCUCS1NrBenVj67x+lfHlPzdTBLS9fpyDSbxhsfNz0Yxeb2iB72X88hxob
6/edI+jqK7TUr4OR0Z9vIN6kKJ9J2h6qwVZkZVkZ5Pwow0vhuSrA+/tTfyWNawAN
45cu19J64AOl56dBw3KFLBWvyPZKGtPzRfF7stCCMHNGG8eFHyPsLeU6pBFodJYe
ed583aVpsDraGz61hRsD6laNjGIWkXpQ6VIXMJ9ddj2oYE/Ry4aCnmCgkjtdoSBE
NAMQhs8S8fRKjt/aA6Fys7sXR71jQGalfwfExc3IbFxrIkSboL4hhbZJHjD/139b
avtkMn7PJmrQJorkJxkQfznuFS2qJTQtJ+3cw9BR4FN8a4f2TumVOBvgR7wpZO7w
XbjJcLGLjvpfmDMjR5SVtGW5Zj1f+5wLGyaZDTI1K4nzJjs56TBn9G9H9G6xTbHl
Z7VHBgZhQJEgzPJ5EXcSPuaHskhOiHEvcJyJUb1Vdyt7P/WM12l7hvWdzEixzWVK
uc8oFvOJbWmBeOSFLPmkeaN71zndTOFuGnoYtb+7boL57ZLt4nNEicke2A36arKZ
cktkAquEWm3Fu7D6AU3FqZ3cBMkzBl3JSa3Ndt3e3ahw0wKWATqQmcAfAP5NkuJ4
Q46NO/Oihzf6nKptAD3g27yUy7pObSyuBwJdAaI9f51AuHu11iJwU5cjL4bMlGTZ
gRMjqQLdN2VR1tktwppE0/WFccoSC9uR53rMYhizOCHg0Lf6bWcjTIbov+4DKcl9
xxiPzAk53KcwoJnwhSEBZwsf3pYnW5Fji3c/dHa3xE+RD3os6UZYmA+yEuXYtmhq
qcc5fpeEtTdeXhkYFtn1WSzm4BlR1gg1sNW8OWOpthr0+whGNxfQm3uuk7HZo32r
oAbu2k4m4Bl1Q8sOXAUf+iXbLt7BIxrP4v6GXwBz2E37KF7Aaq/55DFQWFvbTPTw
M2+1Q3+kFMp8ic/mgdvDE4QtO84G4hnFQaWuzzFLq2SxQEZLL0mpx+Q7frbwFXBK
BfIpHdazCj5aigpOT7zzzYNN3DE+nQW54xiRlHzZnlj/4Az6s3eGNkpFz9ivYrRe
9r41okiGxEbDJRxjwh0+qgCr6/KD4IMKYx2TW0SfL8p0/vYCAjwBsfYUAJHbdYjn
fdIMD2nppNXoKQ3HJdR6gqPIieAzej5vpp0jHipgTTel7xEgw20EuGEag5aSX81w
5UiyDljJkLOJ0WQuz2v4tfKDkZm9sO1aUm4coEkYDi2GfS4dL7+Cpt0WFIyEej0v
S28Vu23izGsSJM71gbM5U8ljVwj3s2Cx9jl58LAxulhqC4NQJhQZ77L12iVmu3l2
SUpZwbahVKaYapbiMUQNu5/JShQkZchxymKr+dcNHWlTHRUzu967/DABjs/E7xfh
LCa6EbTbQtOU6EiBwBt4QpJWX+caxsl41JabmRHvQt8rTPBQe6Kg7eqn5mYZ720U
A12youStzDND67cXnW1tIeK4r8hMKuL1G3mQPMBm2AKgdyX9h96rISghox3/Y2eY
akKIcLpmBim1LEMrbOWJUC3XROdpngMRJTnaqufuWm6d0TP1Gw9mHS6nPpOExdPf
z+jGR4dde6d+cnqdtSfl8oc67ucsmSQixlOER6CN5880iozZpDf2ozHo7neznNwA
UcbK+XLng4n/ErRBNVbtKsokgHc7vAsnNgAe7yq8O87mDFC88E6uEncC4SW2101Z
Z3PCi1c60jA6zFGV4fnKabSDQf1G92xh1ahKKJLER+x4DA5st6WCa1BNls6UZbat
vW1gcGA14o3eWZKINWQt9qq/xdss0wWW19Y/YWy3E1/F5W1GcYRHS49HlhAO296+
pZp2JnYII8jzo/l3TW2rvwUENEVWnG3bRLm/BHXUkmm2Mfc/h39CMVfpa/q5emyA
I1esK+wcYHFTVhHUHtEXL42P2s79f5fB9+LwylKZZnIh/XrufxNLCkO1YwdCc/UH
v2P9bFKVZWlOe44Jr4UTyLcWyFu34GTg5VtwxQ8z7hSZbnFwYB6NNCxFRQEbe2E8
FNoyu5D19/oEcor9O8seCEmTq64ilEf0q/ehbvRio+GB0/JimWSgCVOcq//74y3q
Io04TZI2PeS7TGSGK5QCMZ/PZ5a/3we+KpRsG+rgfwmB/yVDxo/hrOyLFna8FxFM
GIB1JdlGZOJhLVxFRGYUcP6wH79R3E3tltg2jb+GzwKNFQDNmdcqCIrdYO9+Y5JZ
bLaL8CZTi2ni0LsdskMlxOF/TVHGZqArrTqb6fO6DLgaSSOdsjj+Cekfp7JI17FI
+ac7+E4SNcU471qc7jgIlJk82gzm4ShKzXUP9XxlcExrbIndq1qhU7WIWVB1LOa3
JhdNKP4mH1XvzHtRWBWpLAQ0xPEjeZ/G+8H4W4+AVV0yijzUrriQc6+3hf6YDOLa
1ciG/QZhyQqJBckjeeg9Cu3my/niLHeyGQlnVc82WjxfpWddedgsYm8Ou6r3GMhB
MzFcuvaPLWdMowJyh4zTG9UuUNPaFUmCZsa5boGa4n8tD9qVxeDeck0yRtqod2Og
CWRpDz+e5wXYEffzYyZFSrrSuvtPO3KfLOtzq1bjm5Fo57/UYPNyyAQnQ/ZktlXn
BAUoRukyV/HdDeTZ11drTFtuBUzXyNwAdv16NQD1pnMHjiEWL9I17O1kQH5uXpFS
O/aisR2heO5g7wVX1haxo/8T2Lvc2wZXsMT/DuzE1UZgXcLd2hgaysPnFp6YUSiG
mGmj8zSZhjqmO9/euV4MzOyvpMTeULMyGjszk/QgBepc4SceV2LaSeryIvtwDnOe
HEP2k+g9e+CWSit0M62zV5B+1JzjCA7yftdLOfanKJCJP5ny09oqW6Y4nZdLhT27
l9lzGCEXUVOyG6ITncVGFl13LwXL0U391xY0mP2ogwyS4Og8pjx/PX3Rrww0sqse
tbueIUIbPPgfSt9HDDV64bHn+s6lohmbXJUnzYT7lczFNR9VKdoKvYqMcnXM96FJ
LCFNxrSQ8N2fSDv75jjAPrpOKb9mmsEl48//tBcb6nTMxm4vI8wXL6ph82pd021b
EL/JeA4D8WWUz6Snpq8wIsskJ1ifoorNDsjeU7QLezWpBzQ+hin05sEA0iAOYXZe
eO99lZo4nNULivkLUoMVzcxXpBYzkD/WGKJiZ9UMuu9S4zUZb/GwyL2T+Lxh0dEC
IUkwqZiCC0WIZKqhpi1e4oiVWoBkn712pBI6zt1f+okIbqO4Pj//12mMgq7ZFhIy
cVLRIzT7aG6suFkP8pCCiucKWTCPSJYwzGpZa5Cdyk1ekTzjVqwLPUQJYZvukPBd
p0suDqj8y9VlOXCwUqcZIY7d+6cwNwx7vh84Xc1tHwT1js3juk2g0Rwmt0DKdFTK
5fI2f69I4Om8hWCN2GZKphCgICCCvb6oxUz0u+WOWNx9PbXRLkDCxa63YD9fi8K+
5HJbdY723BKhs5C52WsTuKVelhuF/OjbntCbbV0H3II+OlqMdRWkr6uQi4Fi+yTQ
Fi0UhYUZ2i1JM3Q5Tt8u9tl/tR+124Cx4SmnfSKT8R8u/fENSncepAIHxrg/p+tR
W/UGxc0Fw5ct9WOeYoZXQQZemwzOMBezOBxLrZyhbDN0D5EpIyMZiHjf0FKAt8rS
mJ3VMoKDrwhq1EEJ6PRs88qN778Xc1uFzNUKCcx7X2vcVesyac6g1E3A05SXhMV/
Ygqpg8uyvDXGHcg0Izl5dcyLAueEWTLEwEeuEPzUkK7sq1vmCwKtLwJcCwMy6ed/
lqGxxzWtVqc8JP0mAxeClTmfc4CQeVwyhogOzq4XItvLvAvs7LauwgxEilqGuNvd
65sR2uQ49HYoakoDUIl6MwXNzeGE6fhgDsihkXDuen6ldp0ONwY8xRku/kUJYTzN
Dhgyod2fZO7QdfCXRsyRVo/LN1ZnTVcefnS8iSbkfsM9G9VkL/23TUWlYMdgZabA
oUXK+ozbCx9QhlrzuXUOwacXLZL4vkvc6K8ai+56X9iByhcjP1WW6VwpVRk7rkF0
3wSUhnu17dbAEO/ir64iLNnkPBybaq/5BpnkWjDXVKTPagTs4zYsdjHhYrqgX21G
AT1ewEPDd857bYWY+QI1X0xDJf6QJvTICL1Yj/gb9bqhYSVgbbhyyWX40th9HFTZ
YloAr60K65XwH6FYbmPC7f3YSKnP8OnSedvrQ0O8DkZsiaXASoooPt8tT+k3hMAw
TJDfhL4MnbHnH1BIpwbZo1uxe6oYqHAEb6uDqyoreAZT8FiEP0avxqqP3sYcmnxs
g41+wZ26r/K+slq0oys2J5MMALNZ6dKsfIEJ3XPPCfSDkcduqOqPuRdnnBWVfNqI
Qll0JqQmmNid1LczoRxGgXMIbpF+gYrXe/9OO1ts2Rsr5TI6UR9h9Uu2bXmS3zFL
hPP5JwGieRhDSzM1s83jFu00xbpCyhWDa2QAPCRecRKZ5vrUxN+Zw/amz4GWGFIK
blyii4oLM1fwBHUR2XnCe02+ZwxNk1d5EkL0yvsC/PglCweh0OJkSzhV7KpwBW7r
PnFAk4G8EgaOF0/wesknHDJyskcYuvi4gN6w3+KWGRG/nAwEYRhZMMCEAkNwt9oQ
fH1hWJ4PplCDQyspZ/TTleSWfL47i5rh+ZuJgILAqccxkQMvXuil/hFBNnwMExRP
fm7BRorho3lcVMq8VxR06b2P0RrJEv6NQTDB/p7ioTx1WP1o97zptIaddbDeXD2Q
G1YR9+jm9W5gfZ1RKNTp/5nzztbwW7psLhVx/RaNaJzMLQadEbEXwqvg7MjaX8wa
y9zf6sKDLlX30axbEEnuvK8vuSAamWcMLpy1mkwo342vYXSrQsODjRPTXI4PvSwD
u2tBVdveR8YV1sq9ldRcWhHFZhVlXzC49Kb5MuMLw1gFZgPSi+xOsOEMp/PEsaz9
h04uTf4fEXnV4D5HYxDbykalH9RhUPNCMYSIHBF3HzVuZeBckqWgFx2hull+hJwr
3AOc+MlF7ySoDSG7J6gCt4S4OXojbGcuAwgvtzZBB4W+qV3pgALDMydKtK+y0ggk
ACQjOTQffg5k/USRo8rS1bRC0mN07MwXBl7AsSI2wxlp4DsgdcK7MhLahN11HEUS
jmaLKSsnG7qAOBjkcGPSI/b2onnlgieoJsgr/SZH1xF7HgQ4NEvtVQ0MfAxrH2h+
PRKKEmUP0Pwh26D61es9SvztLk3M7jYxFyp06CUR3r0RNbAov3MNXec88CglCrho
Er5/tQdc61pgwZjxLZzHBoUucMOR5JGxb6YmHL0As+pP/5KtloZOKmVEzvs/4wob
ul9AjEmrDhEpmLzsAGilk6LCd8zqnuRL10DpoRDr3OypHuZpX8Gy1ICfJGGAO/x9
76gJS0FWr2VkxkkXhkvluvvP3qfLkIxfq6lXk3ypB3bC9uGNESWb/MFUJlAXf3ip
V1dy/AQIvMtGvxkgEzXomtqCosVF1OrEXLNmfvhblAr/cF3EQpXKlyuqWzrGZ8Ay
trbdLp0y+4jComubvW08qHIWAM7PhmCQWwoSnKhxujvXXYj6eI9+hvo/EvA3xAoI
72CiuVFc9TNCrBpw4AnfFpu07cI1wU6FrjOjywctJ9kXE3f+HSWKQncxLzPd5+OF
Bv9fJK7QSt+ZOCGpH+QzMMgLt1ZnyzPdTgLWHCZxqyZEmp9HhRWF60FgszyDby5w
xOB/OX5qZwHH2bEPaJ/Qdz9GGeMIZkre3MLZznjkcXX7UuOAP1tvm79aXkACrqQS
T+5KvN2rdM2lABkKwCxAzDdUyPlQgFNSe8prDanzThyrWIbkJquYrGkqdTbo8KSk
c0PsPkvURQ3BydOiNjqrMKeoI6qcrYLczxje6E1BCmwO9U5IfmywveVnWzMakJte
TpfHwfTy39zbU0q5If32Ej18T+SR4jI+QMeilqLE03u+1jpHReOoEskbxEA3LFVr
B/yaYdCI6goVEMgwjkh8BIP+Fx426+3uNpwwQZZKDtRgWrHhYV4Dr/IpeNd/v8Ql
eRlr3a/gk0jYb5NKJUdGoyIaPH4NPneQQdjJ7VrL97PKjC/gBsENjPWb4XUuCWs0
S9d15zkdfSoNYSD1rNGFk0GasVyY2RqYdDOZf059+5HETKcD7K4IabfuibpEJdu6
POQNqJKADWYHOCAhd060DrHFNdFO3QpycNYLxUn67khiMGGfQz05dzCP05IkPQU7
XNYriIc8XRMjF0Y7baxysUvFDWG6X+2hRrwjBLuEaxCmZah1aEsAPtDvrh9z+HtF
hNiNubWLNw4OsW8lI4fEYwxA14wL1hPFqzWHeW41mYg8FHOTT2sZ5UQAP9Z2CoHZ
a5ACSX8PiNYcT0IhjWz470NMSiZrPoTRQVUBxULSrTaT6tyRXOqwy7eZIosw5efz
3vgWF669VaItfeE1vinNSYfcj4cjZzq7soD9+OTrPY9DO2tTVnID+eKSweDxM/IJ
GQ+sclDLlmSQBCJAM1efDFG8BZ44Aw7T0FUt2IKj4GgrNcOdtz2r8NccTqhWodZa
RP5qGnKmTMAwbVHalqtzPhylSm3jCS8aUmnC3imJKh1h8DEwp20wHcE7vmaDV8Ol
hXaKoRNyqsWbz6NmjwWJNbPUzthqPcY3soZ+ta5P5tLBzJxvLphPKrG5nlec3Bks
ZT4gjYRWrKT6ZdwzdMIyXFmCZy4V7xa0uE179LkZpQ3akalKJHUE5mehf+w9SQOi
ZfHJKsqV3chvkWlmgeJcM2Jov4kj6u9rRsRAvTKrY1LGQ5+5ZCBTSL4bOkwQpY1r
4Xe9jCpKvdr0qqpzo/IQq7fX1wXMbaf5vldOEyquVcYrCqYPXYK2+4hGO53nv7ti
C+6sx+LA8llWgIO8yOY8gC8bRGtguir5t0byaBA7DdBJvz3XcowGefNViE/4EWKk
633cJ41Yfiln8yubCO+3H3q0HXfyN9LKZYksF3qytqnXJAGvDtj4ZW9FJu4qVZFS
2TMVM021kEBEzAcyxBGqwn/XFp2RHBbhBdlWXmWD+lv514paiht9bxYpkimA96N2
CMpyZA7WExzJG3E82qVKQZEi7nl/5iaRhti+kR7SUzVF/djQYjseo+tNCUwDP1xa
l2Dr0peSRxgt/AHBZFjU4O1lFGvd1iR3Crmr7012JEcHHIpe1WCZnQJzOpjAXnf0
gNO2EUCbsewgaR0mPvG+FNLPlv5czFvN9enJ5V4fIvQ7TS/MRElf69Az5UnSEwes
T/60sJAhrF+d8zu8djv1f66hwIGa9ImmAebafwkaY5JrTkc8QmJ0EXKvQzH8Z6a2
cW7Hu9cUQP3yDrNVnPbVNNrrWLyWeN8KGxbj/8jgIZLwAvZcAJIyTeh4asg0qDRR
QeiOnXz0E6ZI/jfrPAPeyq5Emw3T+m506cWwF5lRBtSJEjNHqN+FTYcHicEernM/
Ye0GuysU5adAnVHw+1ZoZzuQYqMfhY9vwsuot/rza+FYfTJAHjN58sxvBD5ZoxbO
w8fIezv9jLMZ5fvbm8KcEibwqTFYJqpVJKbW4iEthiNjqxzwdh/cW/juXTy037Zh
8/kXPRuevuWkmD/6AzgW4CAfm2g85pq3FEHdjczqgLqZTSP4zU58wGRF3IbCNMem
qoWkcpaWv3KN+Mw3OG5vQUWwElbiHfnb4UBL9kg7UpGmifC4sNcClIMHinrpwCTE
JwwsLCsLF0PuzoaqhWTejYt7bPkZvwNVjc6k+4dyWjEiUdqZxAoKoUCXTwq0PI3l
yy3Wp6utOsQtNC5c4K45dnfpwDUaykKDsp0O1f1CFPh8+sjeWd6wW752ToHOzMb2
odjlUsYKdGPiFDS87iqwzEkHJqummWAfDyRyyR4QWKpBWksS03gyUf1VIJ+TUBLk
y0GQnDa/tvFJdRrEMClJ84X8mK/498GFojNbfYP/I76j44x4jVqecF2vi3SnQFHU
9HFSZPeR8nA175CzTGp8M+QfebgRIIrsbqd/fZK8Q+OPvMxysrD7ptmfd2BtTzWv
n1XQ9TUE6I8iq9SJMfYXONccGWo4kIk/3Ok1e54/yP0VHfHSqwggNyqFhQrfLZgA
/zDFYg6k7H7GogR5lU9HawQgrFD+uy7n1EfyC3OSyj4T+dYh4/THJpbJejPZu2mo
U+NnGK2FUzCdXAfICUZ61nQ/6m+ORr3DM61RYynLioo+V4CYB7JgO5dRozANywUj
ovtwi6qLHOkWVWMEH0UbJP/O3xL4denZzDKVak6wgqX4LJxGabJRkc4Ws2EFGIwr
LybRBDugOKjf+d2OH2I1a9vc9zinMAGoibmWBGGrIWMDzn3i1v2lyb7rW7VMCYcb
9auqeTsI4Afmpxhq1eKZC4ynYZe/hJNdTnM7aMXvVbrqxzL8KDSgozOLSVh5rHBr
nHka8pD4fj2PDRFDOCPC9txoqeCxsBJAUOJb8mbxpt9+ulzTSjKSrHXPwCCApQAF
ymAd3aSapyo9bUcm8bVeTjrf62KG9pk+Fu8+kzdNDDZTJoq8ZwRDeIngSoe7lNtO
UlpzwUKCI6/q1O2hqRvDforzmrskYx85F9eIPMeffn9aiy4/aEX8RPGwAAWCoNtn
IhoLxcxEUpcpkrg1QMPbPwyNUBb+4EvniQ/ytJkYC0CtzAVjzM4SMQ7aHRSj5qsn
BlmfC2EQhKC8bmTB0SKDMiq9BBZNwDoItl6M3niq25wDwpxLHDd0/AmHoWYz2Yua
u/EwBHvNM+b2jARKY1pj1fSHXsj/Sq2nHx9VPMiB9ZlLMI/w9ZwCzVB8tbo5V9tS
/UUdGb5lOJlLGuymKNzxIMz3IpDZRsVoQcWb8JwaXPy719pt8uSKZOLKC88cPo/H
o94Bmck8RdSTHCf2Xz2ouRhOw8jGuhgMWpr5tQvMeSZe6qO8iim8Qv4mZHRm2Zns
31eJro++CY5ZqNEyadrHttG1S+7bRki16a1wWjJ9hp9BbruXl0a65/AhI1n+PAe7
UNgcnm0KB8Kc5l1uNYfrumdanc9uM/rWdWOx7mmEV+2kqzsTPeIFchxRz85KkYwn
6t10ihsUKyvuibm/CBTB7qpngCu1DAhsSgZiqsyjzwln+RYfZbrDDg6eArboeGlT
UASEUiS0KD8d1p2llPHFN/2dYSlwwxaPrgvo8Qy0ELnAzJ7xGBX3Pc7xJQqOXElQ
SH25bz3OBgqRHI0MYqBmCcWMdVOBxovVcOyV8Ku954pB2f3FZ5XDpNUeaiLW7Yhv
0BYuYt853cCjg7DbVpa1fLRC/dqAeuhlAsWWUkH0Z/hVXXW3SmrUacaLfMz10wzK
NK09fUIZuFUoixjCjNJ6gcsY9WQsjeIArX9K9pxWqIUQx2MnE+FI2CKZSocIDewE
Mk1e1O06tsOILJ32LnRLbNVtzqQhvofwrsT4zvJ8DH2Zqgycm/jzLWGXSVmmqmdH
FUjxeaD2xLb5UOhV0veUD3dC1HatNdXss4bHAoBFA+J1/iba490bKDyU/JjVFz4d
mD3e1u7JIljQSDVyIykTPyLCldQZwh7gKKNdK8VCcs4aUot1s7UZ5MP9pxr3AN5E
EHhwDZw3ZDcrJT4NzGXU9O0mUk2y0eUPIhVUEzwKOBhAefFdjMgaPWaceSfh5tVp
XyiBZWikzPzsQJ3ZerNIWFNIqQRf80DsCeIjgJFCqHC1u0xVCpwxQrJeDpduXyiF
ju48PM4V6oXGUJeSHd5IlayOaVhtCiI92RTQVwecgvnUV75KJL55BJekSgyCcQCQ
V/0/M555D1UYuQxfhIlAnzYE7V0N81X9GkQHT4hg+SFlmO6bsK/dsZB76P0FKNXq
/Dq913wD53PjuI/9N/C62IYj8sCK3RQDTDBCBFpr2y5HDanDVBRO0Kiav4rsNutX
giQqYNRoU0+9ObQFpEgmFwUWg6fpDC7syCzLf/PJyHBTpo3e58LJn2z26gBR/y1R
iZEYCT+4clSUlQJEHaZkUTCCRZbi4wO7HvGbSj33yk7wMQiNpAi7XAhnKEdPJN3m
RpO/nnYxIxg0pvZwKGyxPn1T5HyVh9Wqen5dX2VtWZId9IT9KY/v9IlUWZuUXn1y
fTdvwWQRa1b3nitU6uCQ5Vmu5a/M8ByVrrugTLcQxl8MgnBD02YAEOyom83gn6EA
yfJOULmfHgVVu5vK7sQkEaV36xHWu2f5bC2geUOA9RU5k4dlq5XCg3Fm97IYhSvN
DirRDlwwVT6KPqBp9hRFV666Xdc41QwUiHXzCFxo95JtdMvaxnuUvJ8dhPTIWvxU
m8ApdtuCzMmDJqKfTkT7CUPmiFK+79N5YjhWz+jVdHS/k3v3c0wMsrqNaRDomf4J
C+sxVAeAfFHj2kfLIie++zw4RFVzmbGPUkHU6YpDRaNgtrzctnMd+wRCanPbxxFH
nscOk/1lv0DTDt4ITOYUXdeqeZLvzzYVBeh4EWrSQHai5UZpKQyFemcOxI1M8U4p
JjonHIxzYd/Hk/Hq8eOrmTjoPCyVc3LDd7NmbXV99GkCEPLWPAyXpste6s9/QgG2
/t1wcr1AXfseuVZRcyg43yX4I5NDLbD/OEW5Gk96c2ggoIibkrE0PTMdnFD7igNO
PbYKpcqV6uLqA4mK37+zBlofYYPiRspYuUtXfJE8f3hDd8q9NU4kJU/0oEtQFFmM
kFgfZ+RkV+Y1yYtSdUPwihANS9mK2FexYw4MyBMWoYmJjdA3L8TdqdYhwGzGB6WV
ObEKH6kZ1oe5Q5EkLg4f2dncRtiYnhzOoAa5QsPXJc8BkyR1EmTlGufdXBiTxz0r
qNHj/mgty8qUrO/Z4wJ+1cI98/W5OvnV/dqRZ1+yG76zm6Wcvd59co7lMg4v9sNz
DJ0ltbhLRNK7WDJArPDJyFjmdILaF6en7I03gcv/O1CXtz2/kI9DVUFhjJZE6c/z
rPCpZlDhLr60EKGeHSRqG1rtWv1xvyjeVBKoudJLKJKHxTMG15NqtojUrX+HlalM
krEKNSW6IUlqvIn0CzPRs0SOPZObXTFu9+NkVS+EDLr56bGQiYubwsPichOIiPE5
PIoPYVFnyatls0NcdL5jcTOwi1RKhIJIyR7TNpmE0Qqt3Eq5ej85h8etHUCnl1BK
6fc81evIbA0NThKofrxQVZmIVS0HuLytG0H95tDfaVILwejWyQca+LOFyBXquXrE
C3Clt66xMK9o+NnEv5oriD40LJplQbHREYB2weHrkqyj/7JI7prLTbmkq+dfKt4f
pxhe1/exr0zEZcdzjl5sfl3EOMoFGb+rYEHnzJvInNV/sktRTIxFuErSNHLWN/xj
kkAtOtIc3Vr4KfKjH1XGpm6mHff3yahSxJjBcL4IkdP3XKjtB7UcjB9dzVov/kPS
ccEx0QQGblHc6Uc2qSWTboXWfdBueIAYzggnZuuCpf/Bs2jivVfNWjVI3RzLBXsf
ygwCesX3xmwy6/aRLe/xd9qFSZgWZ7/YfxOFLUCrmvLvJLIXVH5tA8jBDwp2BKBM
5H1+S8Y8w56FPWEQWCXjW5bJ6G/abhj/byueT0CS72CtuaGcjQPyogj3RXcrNkvf
K37fI0Sfz5FeT5aWjGh6AUuIbZwfooexo30ohu8MLTNBdiVVAGf0UzUBbTiW/u5W
0Kyb5wNiLAcIn5q7sGlvVprDII087KFv2SDy4LPOpf0QE44Uyd07HSD1CLSTzPZT
ubxjYf7MX123pMbbswJYS2DgCzLuKj7gx1GzR2VwNtmU5gv5sttsjFCTAF0KDt0V
s07b6tbKORec6yJy1MSbEVKwjmHPdew2+5UzeVrItS6PnQ6n+QYZ/kpGb8Ghu8+G
iHyei8RFtYehPahjQ2A7pHEafioOc9t/TAecamesO/uEWrLIAlK7lppOcqmqzO1z
s5j8LRO3schDW3aNsur2MOeZx7qUXCxfKcacLc5VTq2ccIi8oRceh2TyevfxzDVV
KY6dxvhWwyYR7cfOMhdZS8bWqy/fAXftZLlWHeut5ShBzIjZ6RLEZ7+zIXIXyaaU
epuiSzdZzgfJBCq2waThX/KWIvwv8fnzovwwJ2DAjOzh2mGpnoEvm3l+HndjfhpG
dPnTLgvSf0S9pE1VgkAFnLzBRuaSxG67GxFVs+QZSRvUT7qt2bRM3A5TXJrZlA9F
X6avAaaDc/A+sNx3gXXhFDlcqiaBjHT4vm3Mlj6Vyhb9/FX3TjYfqYJBwpLgIrG8
I0QbDjRDd1awNiW7nvhwhqmFLBEzpl8oKASxSKDMQXmVmxY6DnBxeFSzIqI+d20x
dvbNbN6EBz8/TWhrkptvVkImg1fj9rWQCDO7f9BtVOyq61ibWHvwv3cKvdizUbRG
MI74LSgtfQ5kNEtEm1+Yz/gHXmIuaxSXmf+guSOuAJqx3k3aMQcr9SRLChPOUIGa
XQmuB2PPz58t6VKx+3U0LL/HtFrNavqEpJkRyPzCEeVO7E2AhNiNco1tMBXAfMw2
MzdHygXxw3xeyUowB9Ie4c77oiZ84E7tFWLNQ/L2GtQ0Lze+wrGkkcnEGmqVOdm1
WxYvAtGAQx/t5i7MIgY5NZ2AZ/EQkBOPj/JsJx156BPtlddLkFsPzeMdVqUdnECY
Bk7sxRfFF1NpnQubz6XXEYqFz4dFW4gysfCn4HfxnsscOj2xM6MGiTdgPpPcvJo+
LuD0xlYeNHJTfDDLNw30CJuB4tnvmt470I8ZrGtakHqXQMbss09aG77GjVTHa0XY
dMzvtSmZZvkBUVIMYHudi4HUGrC37Wq5BxwXiXf6RuRttqSTZWJODEuxSCtFDcbl
SQJHm4iPGFCT5i0aMsmBHySces14EhpjFKbBKK9IIYS966yvyCsrRWiRTpkafYF+
sS3gqA/YE3+ZMzDbZbTkTezgyf5cxlXNJ9YY22wwomkH54hTwKqnpy+qfXfnp/CZ
tL+z/0alUTK1ZKABUdNXqUEdXy7+3L2ZRXvJFNN5+cdebRh7FH1kyxKpuBf1oT/l
EY06nl3tSiPf+IjEiTSQhye0E+m3xa1Gi7WYk29Fl+KwSKEHH49bUSvSuC3bBsWd
VmjZS0jmN2+059kYY+aMg5Iqw5zHrmcszKacnx0ROqyMU6/K6iDsVk3M9q+ZR4AR
nfHH0aEkepB09Eh4zgybYBWfj5VHzlP/ongOH9efP1mPwiPFJt/ifwdYmSVPLm6g
W4Ty5mb8HO+fTXQdZ6PpQk2kItrw7ODwV54272D0llVNOnf4GBNEGhbp+M8P0h9W
WypsACK6gBARnfLMEki6bAfz9ZzKz7QwdDyIgmpbT5IRwjhzxv9DsFQ0gHuzvmbs
henWFpcC1p4TQmEYHXKe3VHBF9IXhyVn8897K7njcPiDCy1rf8te7S0fjxJYG/rD
pHpkHvvkRSYK+OYR98pl220rZjYi/oM3BxAFBnQ2/0Q9c7IewTXJDn/yjy45VByW
+m4Job9BU2aSVmDKjEm+uDGGFLv+gcCV1CmED0g5vCoVh1HC/JIWhCU9TJkTjQEl
YyPnfE0StVOv+Q7mqctcJRyQQNTL6GSbiATdkoWpT81jMJKx6hgvchC3qfiKM/p7
/SAgH7K4jLYDkP+MtHnvqtUz6OEoipPepMqbWyQ6UfYTmUKqjW+tj8FsF/Ao60sx
Si5uTnru5eQutd0Dm8TIu7VXkFbKKBxQ8fOO4Ycv6zj6O6zmKd5W/YMazwGKuYdc
oa1Wu/PSqpoxyrs2Rw9XATanvCmTw7blJDIymsXemh/B7vbehy0kcP8Iyg1kg6eK
uZK3dnTLRmFiiQmUKN2ucYF0yEhSjkrQDn2mvPld0ilaW4fsp8A3PCdoO09p++FH
wL44SgTazhwdceuxVZrFJUI63K2kx96MeOzKIPyKiRnNVBSfXPk9txewBAgxN0iJ
dncMM5XlKWkY5QN+O/rr6NbjJ9v2gdTr6yTu7ZW7XA2etoXaIP0EC5xT4L/kaKKa
2e7lzeE+pc4skjre8znlNI36rPKePbVSdlHC8aCYWDHQJ82/p/yT9ttzwz6T2FxG
km/PBRSHXHqjiRJ7KHu+a5Mv5KJVVOgGnLlGe2bPRUCyLo4VQHwy+/mrR0VNxJqb
kl+e2YijGKbmtT9VUyqQHLbbVrDaokBeTByyXBOhAtaXir0LZliV4eQ9iQwK1gP3
tUl0mzoBNRF1+F9NtvfKRqQ2SJiOL24WBqqW/qkUGlEEz3HttSu8h5ZYJifWUZDE
HxJ5aYSAITv0stHgE5zuci+5WtCZCmlKXirhJKCDqTBWJ2g0c+B8GZa1RCOhCNWN
UnfE+4dMzBIkU5Gjc1pzkNj56VR4xBaUKgDyqNCGfkyHVsVJZCGCdKUWFPO3Pqi9
NM6D0RVlVB6ZqC3i+mZ5Lk+T6ViReBqISD3mHVn8C6KeIWvZDiPP8FhFhV/hQFdD
oGJTaClh/XVfjoslcTjuqMDaDhN+1GawzA6ZmEraqka/YvYgC14LsTUbapIGHraX
VodNV9fJCgJWp8deZtdjUdSttw80JEHlP94ybzjxnish4OFeLXzeD0zf0T6qTq6l
fbRw7fe7twMcqQWGqKglU3BBDeiwRSzAjk65BIwCL0lBrXawrKGKzKJ9BLktFg2n
BSyDeBYN81c67275M+6iFcPfcGYvlWeZXpWygqBfgXjirTR1DwGzYvotOixhv2h3
K9Yb8Ecmzd87XwbrUE+e9DBV8c2mUamB8AbonLCAzH201aC7xRZFyrDr/ZThcyIp
vzmdLrqJQcyn1oqNYyQYMnrWUcIel3kpqiQOY+n1Tgc5iJUgK2GfBeNfDgEpsrxi
L4nhvHHwEj56eX0gqwWM9sL1uoskZKqEgcGmaXrqDBB+QfqaqsjkDISbua15jreQ
4gbHRFXggQa1JoVOEe+6H1JQ2viy6eGynlg5J+4XhcLbh7OH1QNx/fn7//5kJd+9
eshmhmV0xg4UFzjTpXwKZ45FXJhyV47V87VQMo7DUQ4ykSMi6Hg4b7Rik6jRdAzy
aGP4BXb/ng+09MPZh3fsAhYywp4PIFzXqg6VVtnFiZ76vNdjdwMihIAWqYsLt/aG
gYQTkLJo8bvNCpZDwaUo8g115xUFgWJFuMzZIZuZe1HfY6CLF0fWK2NHK/NR7BNl
OV7F2Goz6u/GLwwbVW1ExsRx2wePhJ9SFFiaU2oBW6OquZ5VllaaYMAEnU6EJ5hc
25jFztG8nH1aXuX0J4OLM2aJhfs7uZDZ58Q27D09hIHEx6LcrsN5uLk6Og73b0Am
y3NJnHGkH1NRaUMGb8WKwJINXS1R3+04BlDHBJiq4i/7IHSkD5/2kdoMcLXj+/BF
kDUQ24sXr3GVo+4OBShexg7kejPcfUiKtqljJ0tfCVjYrnEQWVhHZjKfPSUHYwdv
aECM8HawPyw+sjp/JVt80GvV9N8wtC5Mbh9E/0/5HgQagJwskT7k6l/FVjN09mRW
hfUP5G3DQAI/jLQXMEAsmOtBEymU4dMuzjdCK9STzkVPrdlYNGPbLw5h9CXzdq01
IqW4ns9zoCokam+OCyzgCrQk345SbIGd6ceOqF+vjMWJuO+e69xyPV0Vg7haSRQQ
qujT5RCUb6VTT+eV3K6EZhsNi0G75r9qr05gfQZUaX86p27iWm+YewKXGWQTCneq
pLmlh1OBTfyQSgHnh6XhReW/zt+SrVugxwbYubbhlflf57v1hlQa3qvD4Jmf05sN
GNK1obnmXPscA18XiHUnN8F4eunFtx/9BBFZFJAZxoQjNYIXwsTyse0JDaCtdtkb
wUIruT//cXunM9mknsRepyR2Zs8Ad/RbNIr4ldm8WX115VtZNPjXadoUlD/0HQAU
Len2Aob7ZK+FOOGvWqbqP5TYwxEokXtdA5/xTV1r7qPbnZo61zpJVeKgjg35pM4x
4c1/IU8U28jk1qqQmj2dQ0mjqs0VU76SJ8hXxxC2u/L6Ri0zHp/Btq+jlqUiwFOw
Te1ZMfGbTwya0T5S5kkX7L2ZhsBRJqgCUu535Pf7Zj+Nb7INuiViiDON8gVP19Eb
FB6sbLyM3VS9W6Rz6Cixw2HmAMjPnR4Q5YzeqSdInLYY4Mwd2rtrkvujyAF1+igD
cb6hKiwwSHciNvcxv6T6uvTIUtfcNWz0ANkDta7ZXj11GGiWVQeZAUhWGcAy1XvK
myzXfydy5f+MFHe04/1xU6n5GJwei9yY8PprR/jTzapiuhEpVFSrSkTJ1ItFApJ+
uiJ1I+xXvwbJjWO97jyBxn1Otm/VqpeeFhpaWkB8zF0wJGkFZixSo7etsn/5SQPz
tCFpulw39I9ma3Adh7eFtVcn/9VpxbxSEAcpNe7yFH1G/oieCaw1JsBM9P0L5Vhf
DYd3jF22q41Lbd52l9CMAD5HSJyV7I1S1SRCn+rrxBnjVaYQDTNvBUmY1Re2I/l3
UH6cxzQGLGyL/b7um24+9++P86WbjJwYECWGJIJZloTgZYbHJIFASFnf3NA4uwKt
rfsvUcQNfMXnL19p2o6VPkx9kCSdNGrMN5qaZ10Ybhknj35szWVTEhmSr/Qt1+N1
JGsBJj0mSP8gPWlYjigFmO1OqZVOQoHbpzbZZ3vKRduVGwZkjeMzfy8i0Xs0/SwY
XfmV1u2GgY66QDrBfIfNZqt+oqHD5K1YzF3AlF6Y9O5TTYdVPYE1AvvhV+QGQ6O4
JbFyfM4arBB4rNyONP0YjHHQTncKcx2x31lkb9lSngWQKdmzkPhKDITaVQWN/glY
b1a3rSCxJHb7N/N73v0KODEx4HQh3QKVEL46r8yXGwqc0hZcxQIn9AcnK1Lmgxn3
So5kIOqzwJrim1FhMKpDwtXgBHBco3RJhCpfGcbABufYLIBc1kIRUDy3tZA5aKqD
wjutaUbPewgHFfeGZnWXGw94LuLIgCAJvuK/Ef2iXVGNlOmkSheHN8nyXUyW2EtL
bpJKv4r+FUzqjEKjgWK/gJjHQHrqT9YH6woL4rdezrGZ6Na2GDoEsLR1rQOeQDzf
ROe1yuQn5h05Fjfjqa+Pw2a4/KCpokftsQDihq+kjvTQETZxQ6tzQlQ3MP1Ey7Xl
zC7XLu21v877cHto5Lft5UniAOG03Y158FlqNhXIU7n11Yvz45d4mkLWVEfokOCP
GOJV2f6QbB+icg5NKxNvhXcOf/QfIIlVSaMlVIebP2HoJonTmQ1oiGvQeQQV4B4E
JT+zcPYKetT2R0P9FSwsWmMpquKhmSl1/qd0wAokgpzZPOJL8mp2p03uHACTO9Bo
eYUM57XoUh3m+06EmTmxekwyQm08QnFokJ78at77Hw3G4PoEFcI1hkxO6s9NP6zb
MQStHTQjVNZiel3F63NkGaD1yX3gYTf+padsmxZuyWz4LXSOMIdxab4qCH9kiQGS
UJaUe2cd4Ubu5KMgkTnlJI9b2Afku98Ilc1CAfUB6j9OiOjrhRq02C2eKeH4IRfp
qQiv4AEtoT0ma/ZbZ3wZmGndvtowMhOLqqoq8sTMVeo9QqJfC8HhHGeT9ve/Fh8k
JME4+EeH32Jwwm9F2joNQnt5RJeFCSNLJH71xiPz4ruWepyCzGTKlHNVXwHSRnCm
WBw/FVkEJL+j9OtgT8+F9GVkwpj7RK3wEQzXlQr6MkBioLbnTYpPHbi3iYqXDj0v
hvnnlmMsRBOAQFjBvbNKn8zigeAzsaFHaWdB0YmKQn8+tNCJ+L9n8U66JQSLThRj
Q1YE9FqNBjJ8+FxXy7/BAE6n/Pt2S8HHXlr4tSzJ8Tciqo9kF7kQMOuD7wX0SGuE
ea4NaTKagSg/S1Nz5Yaym5R9LkTkeEMNObRswzrrpAXg/UyO/uo52Q3u1x4rqvkX
LaZZ4Vtg/c/FPlZDb3RJXhWxILNiyvADXITCZVTASLgL2YPadYk5pE5B33IvznDl
NiiI37RhZ3FVY/yej2HV5nJWeMze7wdQZdbYecDs+b7qzOOkPUPXprzBhBxQ4yWA
LhC6BMyE+kndKNcMpkVXWW7pyA1+4t1jH3jpaDZ37C6vLXUKTpbTGEm2QYVR3OKq
I135+qkTJZJWxg/p1BaIzzOu96OuDw6JbutqpwLC2xYEVdkzZ5tSkHe1ovzCHmDU
ytlXLPByGSvQaQ2YnYNTnhSaHxfyB+b5QhjtY72hDLX6UVXXBiFD5sslXbxwX9B7
YCHM+HCrG9vhgAQfZJ0uSdx5obNN4xGEXEbLZidVtfmvoeR6JukCRl9RIMpsS5A1
/li9bIleDHE5MEVLrOTY4pqyw8pmFyawnca7dZnVdU3CHkzFO7Cwd9QzAUB5RuKD
7caJPlVOeSzkgKqjN3wdGpUvzq0ZfrDwyrXMKoQgjKtQMG96TuNjVHxtVV25ECvy
yLPr/KfVAf0sj7MYBTWFi177c8zh1EypF0EOAgwWi6dZLHRqF5Z70oMwBmHoUygZ
XFhec4UVy/4kaMcI8ZhSSPw0B9Xzvpflt6F+oV5wCFW/AJ2E3HtLof+n2SYRpb7B
nHqDj3tLHMgkRCbwQi/mHj1Kvoi7xVHv3dYKMPcP364nLU7SSs91YCLejD+zw1CE
eDWSg1i45I1HpmMjgsVezrDBk7r41k+754/LHU2r3OCHJ02h/dBM4/dgnPBOo1KC
bB6ZqaL5qv0RFBqLMFpYcwG5zkCCY8qINYj8n4caHbr2N36Xb8k0HRB0ITz15PKv
qygcpt+TtQ/bzMUAFbARO9TxyASNjN2U/cCtlueGuUju2oeXYjAZ9C1hocBu22tj
Ub4aV0Mvs6F+p8862fwGbBBcnAkxPa+6CABEJLhFNoF7Q1n3WsKi4MY5VuFQ3MJ4
fjd0yfT2YuXMlnxh9eMJKkMiUUcNh+XNZl3j0eLdRVXRrwvAWdzScVomCefQLFtO
AOv5uchP7iuT0UaIbHEMI8MQUPPA260WkH1Q5ZVX/CutBqWWh2iZ+Gn/1z1VDmCu
dr/N774taZkh9BRFoqiJC23LPyxugoCseZfUTP1DJOb9ANkPaon+F2pqw9VgHDAt
La1bLP3GarsA/A6Koly3iWxig9sEjGDEyxrwqUGpjjwWT7v3HpIhGGRew9Q4jemt
HV/1zaqLfZ592k1o4E/rHAYafkqtP+o7PltM9SX2NkGkwCmvmgmJt2+dZaN6bi+S
8QSeVLsmhNhcsfXDtP2GvUfcY9U7KWhBwDOOgI/yEL/mSrfJdqY++ZAydLSvqNVq
ZJawl9P5gnCdXKOelV1dfIuBID1wqPbq7ehQVYpO9KEx3glEC0TmlehpbuigHp3X
6w6OlLZnvy+CiSm6+SBTzIkv4AjgDQh0Mp2Cyw5RWtQQOJwOGd6WF7TXAoajtsYq
SkrhgLuwbHFuvvIEgaaIs4lpFQIA3FfrxRiP/xFMCkbHMRKJgHMwzgNGQyyiNK8m
mD5BY94Oq6nqrD8YsTRl8wxBiD8J1ENWLynApzgNVPVIOxbjdaiqfCYwRKJPSNWH
LJ3CkgW9NVao7acux9BFQ5NfQfSCRtffr7sJRa5z+TV8w5Fe3z9oOFfcmpJFVJ0i
75gQSrHiL692+OE2A4np3dwPlkeo4zXat/mGjqbHDJKjSlzK/Rq7JeKRp6Z6TJhZ
7Nwk4PGi3FI12kniLnmgAJdW25TUd7iuh4NmYDJzhOcFOzrH9E8m+rBgcAbDyFKn
Q+EZliaTkLBFfc0sk3pwp/XNmExMFT44Sx0FeECJJopuPxO1x9UZvaUQf7oEValO
4Ib9BLfmF2ZTGmbOLlIXtLeOjXBbvUWV3xLR43e5D20idPuVc0sr82VzR7MqA9uw
0YXF5/teTVavqc/nJ6t7wLdD8kAMqTEkavGWYQslsXTklKKQTqAmMoPXfJ/fbN9W
JyWtcsPLkEYtSQK7agACXZ53gRvkpWPVvqgLfl5k+F2qJGXk1+0A5A0QsBQfE3DJ
+m+zS5imcoeFVsDaSkvMkc4N5Gp/ywhWisQhn/uLr/+VfHWZJDGeGdMba4AzQsl9
vnuEGuq15nHYYY2bIoJyanpMn0ajN9FBBnBmp46stZ0hsYkvhfoVkjQHydZrvvIL
WL18O0nQCgZW4c3rSYq6VzcBw9g4S71VbQri3m4Mn7wgbmyMhzU+FLV9dCwfUiyk
V3JWUqGR25PyG+e8DOoo/lmuxxEkGAgkce+GLlc4f6YzCuTt9UxwVJ/NyxTK6rRO
ATWTPysVfUdxYwGbrj+ultN+2cK0A3FSOJ7sCKNsfE8bsX9kQy9P35gDkg7a1gvz
0nuJ37LFUkfcr+0t9uXwvxahPQV//O5dqEPbNmhqm54dfBfNqZq4P8feoCzEBotB
exfSMMdDMnDqvlTUDzYag9F5KVIwF4DAUQmNPFWjuBKlSVU0VdRK8GOPyF3q4bZf
g2zs1goxxZ8CslJNgoYhsZfRl1Qwyv1ICXSvAdFN/UBDb1zuAwo6fINVi1FPiXP2
oCKxusfV2ru7ekvtMhgMsJwOTMvR/o67rj5rMWVIseTdFFQVbgnFfkabXHEQn3rl
RCESt4M4Z8zXK1xJgNLAZAvn7phg/2X7Tpx8fdlq8g66k1VYFfEeAfQInkpNtXel
fD2Lim18UdQKwOn8cJmEEyiTCF9lpBoFOanAKMfSHEbXXavBrehgW5S1TLiL5TC6
3mUK67bzlJm89XYJnAUPCjQFnxlwlWl9ozBAR89IoeUsrXJsbSBnG3rwXss69ZPE
9Dc2lcsa/eE9s+ele+aTZ1VgRsLAgRu2r2LAQUKir3V1wK4YZRW7jrS9ma0pSOLx
H7PdKbzEomsmWzcj9oKtfSsLydFua852Rmyae5EuuoF24Qb4yycYrVAJgrbTuqtw
8AVDtVLFVWDIYqc8+mXWR3Q1WqGpkr0H3PTQJ/B61bI/3w+hTiKLvWwCTx/k7hmf
bep30yAEHcEgNavbgYSAmYc6pFw5lzy36ZVlteQZDENZsEalF3iMrRJ38yHub3cD
3CfjJvbg9hg5MWrsI0T2OBEeJhXWL2aMTewZxBpq63JoFmp9rq72K40Rwe7QWFbb
Q97z5WIYoK14HxS4VgLu9O8d5qGACvuBFRgEBU/XO3E2KQg0pZnbO+obhs1tcsrh
AF4/NekL43Y2yOQbzKMfD9y0nq/YOcydKsUTLAsd3/ayJdQ07Oa0OwmPH3GNrKcl
TRPQQw16u6fth2K5uLili6wP6rzHaiuiZn30GaDQRIl9hDml75HkbK9A8rSxlu0y
zGMnkDZYm0G7Muc+C0W68UMCLsih/u6feppcdFO2D0sVTJci6+kW35u5+xF+vFd7
cyalgIxNN59H8DEYt+Dw5sait6Duom+Z0atZwTjZ0e3f+MN/OspG0tz5/OQe1VT1
fpCIRxgH6K74WjXzYkmOLXyeaXwI2d4TQ8FiOt7Lj2aQIKx2UKf6AViQL/VrBNce
sl/yEghdvWUA5QDZpugUVxPC/DF5f9n3qUNAABbKMA3k/Syd5GucFsgpk0yWFjfJ
+aenMoHOknDlFXUHg5yVYkLAup82DQwZjp7Kqp5PKah6ui4pc1ZikScE9w5Bmkfq
g5RlkcOYtM0YN4wKrGZ4d5r1G3eQJfx6c4GKLpWFDqjuUHiOXkM/r9rEJ7gBTn01
T2yl8H/TLULm5F1/c/w3+Swr8kQq2Wp9WuSJVAJFAHn9iTwOYCcBr0CT0OEUj/fB
R7X56Rpp6/QQPHqTv3rGsBB/W9nyZ9S+11EhnSn4/vwAyNB/gwl6hYL0+/vuo3CU
PY+/tpqyCwyxSYb1ebwYkhnaP5k7yJKjFA3vIUaTUohUnwrIVo/C/Bdpr8HtjsUJ
d2RsmR7/vFDRgM+fUyQwRtNBhH5wJF7388AYRJ93Kwr+Ar/H90i6pg9Qs0GGzw5q
GxXi+OWGe2WCvq8dWJzWrIEGZwgUF7lTLFNYkyyetS+/cCfDIkiJOWQCrAdc5B9J
1PWA45MH9CE7jWTUoMIlF9X2irP/1dsFxTpBLhJYtJ4HbjapA76A55e8nXqY8UZJ
dzx16dGnrZpRJk8HhNHDP6IjDFPrzxhLCOm6PVcEoDBdcMo9VUSvqVCROXTqhzUe
8mbUsR2QFXscuBI1vXqPSmT9miJdPCvlh/Sq/VctFIDoBhwSH8O6SbPFk7L2Mh0p
N+nclgJGnn93WHH3fv2QxLxPFFevS9Xtm6qa3huGhGpVdeIAeebIlPi6aK2ompef
aq1mpFkF1rpIUQKt9qxotyMLX8VAdVAK0B9kyZkd2Ta5MTVEDIH0QE0BPYuFd+uK
fmCGbSTOJ6HtFrilFlj4C74W4Sub/KGXboMHV6de23tcfGyzZMYK8HiOWGn3Bgpx
vjbSmOo8O6ewl3ZNHsw8cAvtm6vmmrSnaREo39U5x62q0+mN+yr5VVPO4y4L9iyU
cGpTBYPNU200jlsFwsUCOMfvQZk4/5q4r8hXTqt1v5FXF0mb14Mdpbm6Mbgoo6Rb
9RBA/By5rTZkSfiCZTyPCpB/u9jXOj/l4wR/jm2UmQdV1bcguAopUB8gJtnXP4lt
ciWfR4fxuzhdN5syqhJ5orKLTOeengRkHFcmFz05qo3JzFLEbkjlj4eZfuIQ/mTd
N4s+IEKpIW/cSkbCO0t8bmNQOe38yPXO7DmG/Y/jdbv4SnG2T4O4Ht9bgDhggZgE
mfeDEKQiQtdiOE5nyK7L7tizitUH8xnzqWQxe1GnxKw11ulvtIZ1QLx7TRo1eo8o
THL6W9/oulUHsDLnlExkRbAy78XGVz2AS/yANFhAe+ZpGxLlfL/rXSsby/4uJ/Hv
SiSNoFpR3abTkcNEQi8IScbyrfmgDipS4QGNQhc/64LU7DiHwZg9wzmqO6EC8JK5
4iQ/wCWTO/P8HL11J9icpdwd5HPApBmAoUK7/FUW8TwqeETRFKRXDk/LGLAKnPVz
3GbWnx7Pm+K/AdOUrLI/a1hMNoL+KFPu9FzQjT7ZUs427vhc/oFlImGXm+6TfqEQ
VvYEYNsGogLmZMlMTwdF4bsqzU38kLtqAybFlUiUFPl+okmEOxNrbYkPPEbvcbTq
PYwCcRaJ2N2izkaPgLmRTRxj+lHoUK6+JyoQ2QbiqiUgAvRyStpDXVLuKx4gV7v/
BhYgMXbHtCmeFahTqJ2QRI+oU6FG3JpTBip35+lXgtvn372tNhvV0djX4D80WiaS
z0XhPrXbrT3lK8qJElVE4iKFz3fSz6oB/8x4LpArQ9dYOj+3usRu0+0k6cAWCOwD
hDG2j+bUIiaURQzvB/L6ZwE8YY/z7SAfW6p6pnc1ECudM2UJRtFz6NlWj3B4O+hL
XTqfnvnvf23zKUqgqY7XYHLYhhj/k1drZAcOYRARsgVb9sULXm5aV2xPpx0QG6JQ
AJl73Lj5Wn4xCAY1K2J79wfAQJ0iXrqyu7Qe2k8bLzubYbXcTydAvB5tnsk6GnJV
tKOKfanaLO3NfLKFaJTknx1T0ojQwMh7uApXnPtO+OnVqoKYxaS3b/QGH4YcUiFZ
ENjY19cVSp5JBkB6835gdAUO4oCl5Mvv1/JisrY7XFlbIgnj7c0JkgefxsJrJJGQ
MnM+w+EVi9hZw78YAlAn4sJ0fV0gA/74YYA5S5bWh3gPDwN3Rk/QaCsLnApReVpo
Rx/nPJNse26D6WcoadKgnutNapEYWHuyXkCB15//m04obOXvDeB3u8bRqMnvJBbB
rw/wLjZN8aA6fD4FeJIBvpN4BqjMcoX+0X1qJRRVlt5QuHM7ogr/x6r4rNFil0Yl
YZ2xNgC45/Y+AcUOFtxVuXApPcGS1eNNJ8RIezZ+YcVAO8EBPndSgIg9v9cWv7/r
ce1/AHnkc733WLReIpfNDUL+rPNw1c2EC8GU3kLqqDEdzFUgCZ2l0CXWQVFC5K6F
V5S28HsWmTQsjLr1hF4u0FkRtczboAT+K1yXZ9cuuCsNtGoTFzocumQywoQUegW+
NioKPTPpeWuHV+iHRLCISkKroKNeL+ZcqH5kbLGdNUi9Ja8lsFBU+gxoUCBsoxNG
QCED4NxrNCZyngGugTw/Z69vefK+oXffzjniGXoxy/ZUp/u+5ovKaa0nvEc0Lsqg
w6wAj75KdDn1Dr7Dc1sl7ik808PZGAcvEyK2b759oIgih3sIaTBfMf+86Jodwv1D
Eyp2Ex6HsWzPkOI5iawdqLStvMQaeTBCbqqjbQn1wxyIqXz6PJswLkHQ5aQvQhrT
lqDDbc5buurvZfzeC6btWHVlAvbVr5k9y8fdHVmDf7UG+pS1l7ihtgy3rnT2qnkc
Lvj+LnkpKrNOF7cUxD1SWCrYIfw1vjiMt3ewceIIyTjl1Uv2OBtwtTe3PneyTwpe
O72Vgh+YeCZ3jNv/RZMoEn4maCFyTZbdcinc8IdZjxKNWZvnG/uEOUH80Y4DA9tg
gAWub/qaowcaqtVIn8LoJRjG2+uwzbqG0D4w+0MDFzo2bIGj4Fi2PSFcmJR3ANk5
clTBEJz+RZoJ7Dbdxo/Ys5dPnsYpSe9QbHtcwM4oYQuxBxbmUUvnZT1+Qo+v6cVf
pOXIPLjK5M4e5rapO3SOJTCK1KAFq0NfL0uLfBwTbedr4QhyLYBoRvXg1f6cZu1m
J86FkD5BB63XUUpm0+0AnQY8AcTEJhHFXNUBl8srESVMoaoe29AAlSOYcdrWo+3x
SsoAadGtlLqwtBbb5lLMGk+ZGUBVaBUxCI64uq1QspRwevraaOXQFqQhTEUxOdis
yvs1DCBrILSi1JD1JeY/II/2vbg34iPf34LazV5qjnM6Do97BxIS1oklSu812K9y
fY07HJmSF65iy3BgYsXmKB9y+m0duBTQ3llGCV37rUdv/QUs4gr/OtRxMimOzzXK
3awPfyVWaMDDMY1s27Yd4Co4voNQwzzH75lLWrv4xKvBa9IDwcxvqkaAiouebAOk
TePD9yv9YV0qJusEWwrZyUWGhcNvZMYmaSYRQii7w94xCSUJEM6KDvuHqR2n2bv+
kbuCgnv4BT6VtSH+s+nnVHn+VYfV35VU2PShIiQ2Jh4I5glD3A7cAn0a+X3ks/PK
8sRCgCLjIRzW2RlW63hvdr0NxBdsqzpu8bKWiXh67o5LBEWxx/tqmtXacfA2GMtc
NhrQxVq4yJVNK0w7oXKvORlg/wjJG3uSWgPGEmDQiLI5ei0J/zV0Lu7jlwNxVhxh
41DtdpXxjvsvPkaIs3qKjykaJT1m913pWp7g6JZaKH6gPvmn4K+4CtuYzIzWg1Qg
qRhO24wJ8J3K4FeTIJSrRIrBVqbCxFRixrY6rZ3atLd6NSqV9zGS43zoVZYTBIs8
uEb2/S0+PgPX9/6O6MC5+IerJ3GiRQly5sGjtpjs+Prokg+H4XWHjd9VgJKBACE6
1maKgY+WUvxyWd10g1K4ylZ6nirlxZMIhFpL7Ib5kp6dsVRENcu5HbCbylTjgOzy
KEhFrQBZbiRaHJqJmMrx9upRxpEOeVux9lzzmjgvhgr1MbmutWgN4sunpfDx286f
96W/idY7M146PGZOWzx9n9WFbUgCxWupH9NiANy5NAG8QZ9InYMfqGX/lGFwdSYD
17ezAcjvjlpb5ogvNdtAbWjk6Yp1QUcrJN7FveARYNWPFKWPdP0fE4XYLTvooHj4
RwyLlyB5ti4pdIglyw2ICGY+JsbnFmAschZV5JzniWe+bBsUOCTKnDdNOJ3j6flE
pp1GijNUmdEc4D5G5gGuRv+mI1YR4gnnzUJQf5eXB6ZWwjU9SZUzGvIKrxNHTErz
BZak7ANihI9Y7Dubaqw+g8SVHdgwdoUHUCiwBz7OJcjXEMayxXoPLnr7ygiM5/34
ndE9u8SFv+/bNin1AmoM8K51gfDpa5stDKeq6WcTUp2C6KuWzwowQwujmdDnEHcz
CTxQp5ijcxgm4fAmNcGqvSO6sjaEGd5h9OldiOk5+3JpaSwjorecV8GYRfNGFqhv
KBdMNhA6OQBhSxB5TbA5wUkZacjPrVUxqDt3jJJbSt4zxSgxLNFeiGuR6vowR2xV
hDTZbfqXYU9b/aBC/wD+1DbYTRyVFQjOuBhcm1ME5zA4PqugjDhCFfC7OkFqh/T9
v/z/Qokt2qJuHqwuy4WiOBVmJD4xLWh7tYLzxaxT4evUQCufPOZi73ntbgvA5LWM
FPX4jOs2ZPVRiV4DPoxi4Ysuw3Gb6xRmRO23heps8wxAefdMFw/WOBM5YeBD5VPn
qVXzlKy1c0iLYumEQpaDgyp+wdYm6QTWYxLNktYSIC/6TvS4WxfPSdsf1ge7FRAV
033uvA2w/oOdw43D7EB7dm+aedCYI4JsEZ3xSd/jDSPV46cewnDglj6DnuZ0jvZu
FykDRGpx8a5isxWs4AD7xyVm9WGymIo6rKiRMspaTACuXAEh8cnrhAeDVJbD0Xqi
6Ze5yPDRO30Do0M3hzTPycBpPj8BA8MffXveVCj2Z5n9Tz0qPpB//p3ekMq/x/VI
o7PbonnB8fmEqxP8Lepiy6ZhEKNvk8UM5U9Us9PJCJN582z43M7sT4+aJPfiwBvZ
gUgdiyzCmHL4jatFOhwMxBbGRCIuVnQICaa4+a4Pf/2rZTWok6to5kpY8VqPqoqY
zloLrZDknHV9+B3gJJPNHL+QpAM3jtldsQ1QcSDIfO69zI9Yxsg3UWAktKz+HnWw
sibqfIrRAkRPd+eYmW8zf0yIfjwzlQ0N0ErCTQ5XCjfwDLiSwM90jrtwzmsq0o34
vobPnVg8jcIIbCsc6XVAuk827p/W5XT9YvKRDJ3sBu+XeCxSywnPUwxZNUd3zSOQ
sviTvZIumPxw2bwV8lFN6s+IeMs67Wbz/qkgQk5umVPn3uUoESoiwJVP083ngGCJ
CVEYfEhHRF+c7JINRgX8hVqx2rcF9V8aWlBCnzPro81ZaWM30AyqPOkMgFdYr5+f
JlAnZQZcXQHTobRPlhgLHTAxVBmfGtqzazibUV9kp04zGdaUbDzIBgQNbqsENs/q
Tq8S+zX8FTh+rzPDyr2RFxdxG4VrqSdeHCCQHBHYoiqK1n3KE3GEmUs4flzKKIBL
fdG+GzPIYJdVBFgN/cxJOEYJ2jlr5h/ZuoBz5SHlVfPIfKQAxcaqYFC4APc3wuo0
OduQpZnKS3UF/61IkKQ7ulPEeaH94XE+eUtzJziy/sSniPSzg7yTqYKRG5UFMSV6
xuZE7vi9dhVIZjgI69WqOAJfNC49WQpnFLfEd2mLnqGrMC3ysv04Ya/ox4zpWvYJ
2jAUmolEEPgXWj4Of4kc/KobdKsUfA9oX0yta71CE2QgynJ3NKfQtIw++kL4CZ/U
/TCrXEeMexMpC894+ugNnp6cL/afa7f8aWrO3H6KNmujwxSGoYIMtUEXfuL/lXUq
nND1Us7YGGZj+nek5KrSRIh7vam6GBPK9g1LlAoUnZdlwDeZ8jUxPvM3VfDquv8o
KFBuQcUpo4/hpNa446p3c76tlB5iu5W1hewo8Mw/wrYVleA3TO0mpn5erBiwwKvQ
g/xiPupxpLymmPgrAUcCl6BCaergEtCLyzZybTtzIpTmWzTHcNlSRkOa6YfYdDmI
c0wrUEltVSORoIMnr4EkaHzA5QDY1ZIe4ttRYl/Ry/6BwwB4MDNoXm/Dyh2x3I5c
RwV59eYnGc9QBxsibtB7nDhmLxwX0ZXaFpmTaZxMdGTHF3Bn4CRMsq/PYpVtCWHK
MvkcFhf/Jf7Fy3EzFhew1l23yHwtFQBzvaWB293gbjmPWZsSKJXsuwNxeWOt4gO5
NhfXsQcV+6IwTmkkvqseVIV0FaP6ftfrAhiJ7CVHUd3Ytk/9+UYU6hgKOdIDCwNQ
lhHg6GEgrKclodmaVdlBlI7pQH4WLAqG7Ya0shS4PNrbqtEd/avPkW1UfesN/xBj
L1HfFKlRomCi5edwljNpimUn7B59A+5pd9It/LPPEt/y2VpXBhG8J+Wyx+bR2ha8
lyM3pGd9MZcWBAil2rM5/5P58s3CgbYvmKpK4hkoREYivFOVo0+dn6HoSfZtJa/a
5EhhHhGyfVDzh9C25j6/d2DkoM0low8nGzF6v76M8A0xzTMIQQuk3Uoc3i137GeZ
iZLUKbwdMYGoPHyy2kdsQZQRpvbihguefzmzLb2jITeqivOMH/U7kFqWgmBS1NwM
fYaJOCVlGv6zXFS3zslErrG+nNWOlN3d+h8uUg6CeY4by/7/SBJ7gnLPJ3sh5ydA
TjVU+Sys+RxcXr+H2bluod1ugvFU45UwQBQCGbAVAYFvjd+Uaz1YFR9+dpUT2na/
3GPgjko5SHrj9WwmkoNI/1jdd+da9Ok1hObH5ORn/RW/SwRv5fchI90VyO38KMlq
kcKCky37ihxq6GihhG8bV065q/lwYzDDFw2tRJnfEP3v7uo8k6YygXyLbHGF/Eak
rPVzSGkYKoy7D6f29jbrAwN8TGkApo28u7taYCpbic6cgZlPp9Wgg7NnjIFZhOUU
52Zb5JzxP0FC3asufNFgsnmM95AtPGBgLFCbVRPDwVycI5py8B4RNW0vo7TL6HI4
wLA8d8V3cr7PFS5CzjlwwkmZWbPcVfQNPXaEM7hpQX3MmbaffhSyrGll6ujHo09G
rED6O1kjEp+Gndms5VrIpsgxhz/gF1dHlsEYIrJAdPsblMiuli2Om4P9k0/inFFm
BPmJLnmgudSP27N+bk7qoPMsJkgxGfW010N6jeCKJAqKX0RSP/L4c62tyS6PEF+F
HTvf8Z81Hgd8NjxhsbyjkZ660gBmAEo8pXAL1/wDfZft9NCL4OYlm8/g9Li1EJXa
GCyfPzXr+tx+qeHAfYuVZnt+GKPG4zL3nutF1UgPXHWAsilj96LF0JNok9H/cVjH
fk1WtU3lSAa2DXOq79SvLo+fJy6UoO4WNFISrqCBauDSGK1rKbEj5ce3qaBSh0Aa
daIbvbK70BWj6PBUGe1c2pKs6YWrw0aht99YE/v3w2bc+CXoxcyHEsdN3A7NTr7X
UeiwJQbbgdNo/OERDneiv2jpZ5QEFuhapLjtAYKfcKEOXy/CXsJbmIKhUw/LdDOD
V4HXBd6uJ4F0aLKQRwMMQUAoK5b88YaRXU7LD5bUpdcCr1oJ7kb1nIlKb0PAmOv0
am0IrgUIxAW7jDLh2tPa9PnvIodtJOwl6ZEEhu1jrZ5dG4+g4MW4mRo1trUq6oUd
OZiOfS9/2MZNWKYSBEnBbbywliiHA41keEim01xExxRlg44phFFUF8L4NMBOIvyX
ycJsOJbDYT3R6h/8/YJoZ/KAEnxvVlKQKMWxuG3wt3+4m002o1dPgNybuPOfjvWQ
ka7VaIs29+P3on5c1cNTHAWrskIjzciKjcV8RWpSDkPnv9oE4kAMng633ykbdirH
X2ee74HUrKO1r5fY9A9ue6q4YaDuc1Bmtur+lhXkBHQaWHNWmvfMnnUsfFoneqRy
PeEoLWEX28GY8NKlZjUPVil265gE1FzrL580skt1Th3ZEc11LKb4Bhm9R8Bell4d
edvQPAipDD4eMn0NwAXI+p0hdbYSElsYo6mPnaLXiAQeWKGAo8k5ta9TwGKFPYt2
eDnMMyQu86bggkno3m7s6eqHDummEOCm7IkUcpfmJAKxMfl1kmigAHff6MYbzngs
I2Ib0KFdmJFLRhJfWl4dMHqOVpixSXX7H+liBnN8FXmRPeG/sddGI0PMKtFzShfv
ssmXV4eamFPyLAawibB22U1Y4ZD6HFPM09bj5swG9KexP3DMVgfC8M/JsqNAIC5a
plIYAsZfa7QREkysk5llbMOAdhBBM52OP4P76kopAL7btUv/X6Be+AcShv2xcRoT
PNmaHSW+wC3QvVcsgabM0NFzvkfHl6TPYNf9rHM9j4WzwKS5JTQ9A8jKbT1o4O1a
hYpMl5CX4NFpMvBkDX7PiHY9CooTjcTM3jDBflWCuc3UvYFSfVjH3+/+jaPaIV/G
O73KmlgqPmr5oY1aOdbE7q8GaNbRur574Y+eGwSJIUIrw1oSou8JSWzTWWImX4Nb
ZA2e8H9Fkqk0y8C2RBxNP4J+xJF0qAhwEh6XfqRB3xfkowByVa4qu5GNcA5tluIt
34JmTxNtMCRZtJL9iry9hzZy661Yv8udxVgHD/M5p/GwsUshR7sJxCesxq8RveuP
3z26jWYn6sklVztgjs26pXO/DaupTgj5bETZuXaHNQXkAJjk7wlgGumKC07UY7QD
vhdCTEhIlAawzfWOTEbmZhso7K4PHKMHLOiYm/i+NBOMP9jZpyEIafyg11XGAijv
vov4bDZ3jlJ0UG1eyl6OfoDdTRpeX3CiW9gj/pAdvR08es/KsyK+uGQFt/t8wuAx
YXGo2WterPSdsWsSQLIs5KjGfvZPvQbNicHCSPA/mAEhOSvDH5s0+pVp+05QIOqw
zph0przrry99mbaP7W2BCDbxg1GSDw9zw0i6OerlPM6rLWTe+xMqYTGjWiPX5G5c
hMtQogx/XNt0K84XthfBnI31r1BHCR9xvUw7GSxow+5AnUZ1vxvRQbfvA9OSQJCU
Z+yn8fOFHP/m+hjAnng3LY0kXbwCqS5Z/IYOADkRzTv/bdK/+oLRKPvUXladrIjJ
mcRlWOPPc3agFtzD67R1gtu+I8UW9TD1PbSRiZ0wx8L+lDfAhpqrjpKyo+mD4YaA
lroQMtvIzxMe7oIZjp3uFDqo0Ac8VuDIILD5KsGrUiaBD5uGr3tsbVV8AdjJHiSP
XMJ8OCnie51n2CIbmov1Okm/g2+QBgWWIK0zFUSAUSRAS6hGZ6F90/PBFqZ0aW17
PImyfqwRlp4QZO4MtfeYc4qlUV77dh0kxFkH8C+GgC/LmvHFjQw4Ut5AvUVHhik/
WEVGZuatn5jHic3WOzfTJ3gFtjI4z8ajTMzlAvasHIhO5VfcBDyhe1sKzgyJt+m1
77BAxEzLU/ITOJjbbFWADZotUy1OdPjO7zWkoK5FqYK3pBr1tG95I4MtRRoMKvWN
kE9EaepAFYiuyPV9OG8c/LbwOpJCu780YreBaIaJrEdgROdlV6E5lH/0OFWPQY8E
o8dh9VnwIv7rgQpSzXcTFfbv3pJJmJxMTN1/ggGJ2ZLmT++giG+Fb/v9A2pedm/X
rz6bKJM+xEpgsWa5R09OJb/RYSjnlC/e00rHeajnhULIDGTQHlFzBXhgLHnUXcMF
xX6fy4VZzev6yZ5jVoIFWg2SLohZzHtFtNDmFbncnpdh92nCVsAADdPxzYzPS+5P
9S8iKt/oJH03qwzdarURNMwcvZU00qXImR7I1nplCUoBL/gKjVc3A8udpNR2F1CI
WxGAafnsGykugBXNKeJa2/RM9mUdy7O2Dt2cgyDRC4ZVBzgGMWz8VDBE72xNjF+t
su07EVYR5Z6dH+UrZAvBYAplnZRjM3leMkCmEduvIRvtXVBxNIb5rjI0h7RpD4O4
49m/IkaZ55MD6f/COF7B3eD0/54ta7CLnoT7DuotGSAbAnSQe55yUxVz1uBHe+Gj
m/2wFuQmywN9LtjEUUTjHzXoV7q5TfxEpVoApf/2pmkJZQoXjLrzTSpOlvUigAFw
6Er+q9T8Zy4wgo7Y8YGR1humUK59wW+GEjdC1DwYBSO+t1egbufPMm5VY1TNxyMJ
wvVIHdEjDY0Opu4Vq2QI+xEpLFH2VvcHUag5dynX63Nak2px6JZj1KHXfrx0BQsV
RkIRq49NTyXnsWv/SRb2CUD8e+2/s08hP8Z2Dk87PSaTP/dBgvF6/5NGKBAk6iG+
IwTFmfq9vDaiOzPel8ro/gAN3/1CWDNNCYAotPeAGpMDUp5nuDaalR6rRJ2+zAGX
Fr3CwI/yervxuTfFL+5+v7rKc2XWAq28b/KCPrqZS53Ky4t3wlqMRIV2cs3fY3jB
L1xKW8P503Qq4Gy71D4LWisRcwsOkelniVdTWr+g+ihsvXQXXu/dtu8gWgVUDMkD
avwOfGTWUZQmnEtEbXND9Ai5YXHZKSxn/wo6RkHe9Th2HlXKS/VC+83eTt5IPL4j
JxfP6qlLIUdnHopQ0mXXWTTAC2mtkDPO9HKeEQw8lN7A9MglZq/bQ+VYEC96dbSH
yDKuvC+2FcfOH8w7DBNYaT8rXty7v8xOgAggSMmzvExfTVan561vPzzQPrL5i8bb
9VlIvQCylhz/cGxYOQC6EaEc71DjdW2qIpJQhRn51GmP+4G3vw+S84xk930cUYEb
ti9fsC0tQ+0LgyJPmsMFe0oO+3AexXI/UmMDPJpFyXlfpINc5Boe7MlA+fLFFfGW
NINWfwSazqNJU30N5NVCwR1qPpLe/iCrsq27VwGqpisKK/fMhOeRrOtFgc+xPJbn
J4WAMK6qnozwk5sIFG9ISqqiIm57ZLE9UvFYtPSVgpXjmLbZZ3lNJBmKKiZnu4mk
hj90T9xWgIbf5RMwQDj4cDwqFsxw42W78EkJJoJaw+TMul4zLWzEUgodzvCRrmmi
IAIbyQKJeV7GqM3W9H7zsti7oQqnkl3ow2U7aqk+0th/aXo5L89FBFdMpalMbGuZ
ByyLUj5ydAswu/7Ex3k4JolKHxEiynG7tzYWj/pkJSt/mIi5FZHapM0ddZLSktlY
E5APDosXiyJQ5Q1pGb+WIObIw9nN3QmP+ADjTHzaJUXlCur07xefYg40u2ssnuKC
5wbrRyKP7paUVKoOtZu/62CMBdJQB3fAJvSw6sQlFMjuZTwwU5RiG47xB4BHHy56
PXX7t/krOjmhrXoek67C28XfYphHT1aWRzdslZCKre0NfjUq8mUzY2G32oVzTamT
84+dGc08Z9JmlSIzimXC0WX56+H+rd/7m1l0IKciP7/9qrCJm28jTpFIRUwVw6rC
S/klx1GSmeuFJbefPYajIxomi1annnCC876SjqSjEsDufmARLpGtwxNQJPP9xv34
JSGttyvmlK89LBLjnTaoV3x7iBiLecKux+l93j9ZqVu4ZXM86iYxEzsAXsXcD9dv
0Pg7TpmDz5jwyzg7H16NNUH483pEXlTLGgJOmd6va9Dq2VfvwTzyn/zqx0Zh9/D+
CsrLCSNkM7F2k3Vmhe4GNqSrEuwmiS5JZ6vPutKdPrO+DbI8eZbZoKYZkVY1af0I
rC5gI6rX3rLri5NRR2T3Jmvq3gyLIC6+qMl2lohz+kwaTCJgm8DhsFcKwcGGAZe0
bO4LQjM2NFPgUVonJPa362HCt5naj3toVBkxWkGDbZnD7pWdBGiMSUGmMO6md92L
ZK5SPkBmqycYusckKWfmCefnxiCKU0fCb/ur4oMi2gd53yPcblHzZXK6rIsdNQmj
SkiNwvh8nt7RBYG/z8BSjmw30PjyVWuQQKtA58t5ho7mq9CqwfV8Hvi0KA4hOwNJ
Tiis6zGmtaRyOruenSi0r6NhevwI2Dpc9LKSR3eVQtzPLYzI6xXEfOCfP1SJdipz
lPmwIIv69cMgjfOKjLkCgPoapMbCCinzeXFjtBNtG8E0vIyr9feejPR76rC3SLgC
hjW7Lozj9Rz8XXg+MJf2xdA26Y8DqXE8b3CvTbX5h4kVbgGD/IMFk1lN5s8Q/I3F
MxW0mM2E+i/giLlB+UPP1OA+se5JGZtm46YjcjkTk2KjW4eNrs6svT+UH4zcKdmO
wbQRvoFFlAnhdBmyhwKlr3m7mfbzwwfrh45LcirhRs1sbcdxPj7TD3eK4i012tPO
AQr09I0cAGDyhlu94ldlP0yWirS8I7YrAO6VU4v/YOPnx47VjYfKxjeXw9/O/ve3
5ASItH+c2g9rJ0qjpPYEOBHx/PhtCRbkWwsUAULdSzjsvNoqlM2I2Yh8ao9LFa/U
NWXDVrDT6EZRMVPZfv3Td7K1nr027wKfPEYspjLv5ZCOu8n8hRtZLAjL61yF0QBR
6CYncwQ0TrUeU0TUeupQpGOM3q8P45DlZqjIbAGuILd241AQbZ9+4DsuMs+vmOhc
+4Uy2MeL5MREjjfYMtGo7T51ZOY1Q4NV/d9J7z5gbxOwoHrHnS50w3TrUzS67rfm
c6ci4cs20zl99DiOuNKQsPhACP4t2n92BV3fzFRIBYoAiu3uyunZcZeuCHveo6A7
JvsAKLS0hW9tX7/wCg2gBTcSmJs9r5n/asDX74JMpshryN6ty/Xzarx0nnFSFpAG
8iQBOseM8DHFfr+sGZzsrlbUhq/4cOiUwGmmTklfo7yhynrZXj6Jtmp/xNpAbDdA
gLWOFkRgViUALqR19AifsnIrqpqKwrT/edFz4LPfkbC2tlV7ceqBgOJ9teGaoNmB
dBF3Mg7sn/gAFjnsANoW2tmD6Bcev3v2gF8ihNjAUskrOvpvsAPLl2xQIxBQMT5n
gwArvHH4qz3dc8/lzh6G/rqdVrRecrp6duPmbFVp9KY1U7Jkdg3NBG+OGS4cy0vZ
z6/ec+ih1KZ4sPbaj+BkC89fKN8VE1TCac9R6B0HmeoNl8ZIUBzWeX1F1zfROL4t
y0JnmIHH8YECFFf380oy86rtIWBBbgphjlOupeUozFa97Yyt4XwCIUNX5o9fm7jR
8dBj33+bIk6KRq8YmKnbk38kUBrR1x7WPGgNujnMvZIJWzpjy/PnD3PDE35KkNmx
a5UIZjG7T86lLyKKORtIMKwbBojvjC+kvz0LSKEtlMFlwlpSpdyw8L+/h2gmzlh6
p9MwwvcFyH9utnTNP8HM/vC7VHahISAthpW0oOVBrgUYCHMqbhCpEbZuXUVEuGNF
KnZuIMXivR388cFm2dECL0Wz6nloJ9fcziuShBcswFhzZs4pX41Em1w+nVlmGUYw
A0FWg8++1z4Bowv9Dj1iwwN1KTI1eamjm2jYLG6p+1ipaFM2K+MgvBJo3eS91nA4
uoncRpWYk7GVcb07xQjJpNgvuwKq9TRZGFuqUEHzgc7MS70rOc8RU/GxBbmTwgsU
ESFQV+aa84nOrvmAle+tTsmq8BMr0jUgDzMm9c+e3QAVlD5hhDGUlRiosBXOAjjD
t7IzUDY5jXXHQYHLZ/c8a8ilTaQkJoKsgWVkqmKhFhueDfHfbYNFvxIHZed223+V
wn6kB1kXnm3YI7QnfxK8oj+BMSG0axHD5jXmDHSHv97ab8GJN0CzH5EmLH1X8yhU
qokiO0fItellca9looqR6F+c7T8rENr3yd97/SfMPTdFlIIKTuc1py+9UyL0fiIb
IzevrbkbduNbH1hdxXLn1Bb6PZH9+9Y1EQkfZOrwP/Rusj91tgoaW5tVXIIwHo8O
+oXlVNisQTOiczhNKsGNVDeCywRO86FJgYzJ2GWMdkp0Fy7d2DBcLNg7OIOC79Zg
JTJ3gI7HfbYvX8JLGfoSA59a//vfPcFqPKfoSbUkP1FLyYlMOZgMD54nBhg88sMZ
fVRoK7VllAxpEmsbSB454lhHMB0gYpRObtoyGe4mY8rp0pi6NAAvoEo4VF4BkZtD
0enH35LSDuKR7dVV3UQk2s7fUl5/3xLEwPj/eQ6Nda0MOrN5i6KQHogCj4HUHTcq
2WkV1c+9Dy0Ow+pxMleV5CzC0p0+q1N5/5apP6u+43R1BdB1VPr8aKEB9kw3KlcE
oIu273oiXXBKbI5V20JNHHgTNrkU+in+9WBKPVPgGXECkSM1jJdccxeD/LRNtMJt
0vmL6DAIKrSF4LKZYyxSAf4mtpe+4Fog/J/27DMVrAUOmsQYl0+jS5TsZr+RXsRV
9eIAQRDI3fX4h52hxylN5fu/1dbeJZ7IlQytH3zeN0yTgAMfdJzmgdVVQZm5usVT
/s29dCo6TPoysG6FvDyoY6Zyw2PeTt1RKzhAURbsR5TxbcLzrRQZAj5v7De1pCgm
O3TcqVhIOGteltlNtWjvM7+kfFDLdJt8AmyVMx9kEAuqnIuGL+QY8fPlgk0oPVkh
RaACIfFJhVMVtdVk/06wauIwnEuHvHFY7oNOnjwmaW/qlQitoPV+biGNLHdovShC
nzE5dXN8Gl89SwvjkmblomXjBbrUql0XnP8x9+kRiTWt0gjSUlfk/gr/oCqJpchx
Z/mwsjzAIqu9mvCAALHFFlNqNNYGGQGPmr3t2KP7K4a99OtFFddNlD8/wmSOz879
rkcoWvBpS2oXzzBUrcNm4nyeSlwStFNsmYglo5VMUWjHxEdQulO85RbRCQZtYVd6
MgRMAgmd0p53B0HvZaEFZDNmNYcJnbV1GHvIkpiTraDZPerbNxzNA/xqQJzyb1nP
NVpJnFRZBou7FMcqyjT1BlxtgqrBUEhGV+ycSvbu33LfhEmeevm3qjNoCuC8fnis
/z/bcCUO9wvD+Olo4AQmMT6PZMFhsEdB69apzSfSVVL5irlCuXME4KZA7MN/g85T
xTp2UzyqJEX0UmW+m1UgraSCSvqYiKaO9/2HfNF7dAXjv3Rk2IsDu5KnCi23ksyp
hqsC6CxE5R7Zq/vSeGvkGdi0UH93b5+SN6ApcrOEDM6IJ6hqY4EleqOTtv9vlEkF
dkSGGeIirIzD8RUtb37J1LlsBAN8e5b2eCAhTaV0iiRX1vOeCIoolAP+H5hN+nib
ZG+7+IRZ0hHuLgSfLL4BJ8IX/OTHFoFSKqU50treSrL/chIQ6CO6pJzGVIqfgUmd
VfDvkB7fu5GnpCaYeP2kFMe5+jWc2D2Yp/Itj2FReW8u9B9gGt1RXP8nnLNgKrPD
z0CVfFi503k+xqKPR1pgGGbSHif4tgzP2iZAdP2drCAGJs3rFw29R+tKHVtvrvDZ
kIW6qsu+Bf8bRmc7dnSvCXD9+sP0G4m+4GM/ha0bwYZIkK72nsCd///FzAULlpQu
TiOJnRYuUQDpUrUfn6xIx8lv5s7WCdHrlWjGRSC0pzZBUughTwq4lQFuBB6y7M5S
GSkcdjbP6+puMALWYF7TaSjWNhz6vFrAJVMpNDYvyMIANyWc9JJ+VwuBiMpe0T5J
l8iBjeoftBNeVsUUOUerKFEhnsNDkgnGO1/WXZxwefYho9zjYccA8nmUPphlBdaF
nFFJnC6N32yWwAvn+7IvBcHgygb53ot2m69E60P9b7dYZA/ND0oO80gK+56RDiGf
RA9e60umNFsSgw/2+D1WC0UYPihThJycRc9w1QxEzACnTHbqXcHLnzOvwpsW3wh9
xHOUPT6c0rXyI7pO1YGdkJsn5dFJS4XZcO3YU1O6PJGKtLiyf5yy7eW9bPLWUP+2
LkgKaFyS5EP/NCHgQrZvDDsKqnQyw4RGa0Rnbg39wMJGRtUSxR1lFtqeEoImRhOu
qrjfEvk7FNWEBaqq3FlKo/H0KN1ErEcesZhGOkOY1zRmg7bWgH/joq2mNgZMzacV
wMaJLPD2F9owqpq3tGK7dX0m4O6fTUqbdKB7WUnQq0eW6oBhYZYOhRZOvbQx5/dD
C6zZ/Bv6x9R4MkHpqbE/UD95FQ+/lXBDe+7BKVBxoyYBc8QcWH/f5F2ic917VfpZ
DMq3VXkSxQVksaV1lGbypVIgOpcozqVqBRKnAyQ1mkBNfwiJU4HxWC1hKwv3Dckf
cNfMT8A9iKqonKRLw3xcheKZ/9MdKc+KK5KzuqlbT9c3cQGOQQh+4lA/dSFTEh/t
jq18p/h2NcepCJdlkIfFowZQOPT08jUOJW+rV30OaG6exp3ihJu1s4TkyEkDY0jK
HURr1cdpksvNm/JgS0y/Bhcpo0l4/DDoaqE1DrdxKj7S0JnbCeJiBLOjDb2y/2Vy
h+lzdY0CfW7k6R6cEhA75UNQe2V8rxGauZGFOdkIXLRl37fsJIt3nKAHdvxpZ+CF
OBdM+eIA2oQGpK2RSAA0BKwapAKsd1ychUcGkBCjptp4wbnEVegKDeiN1m/D26J/
EuFyGwqkIoIDtpsQGD6Mhi4IupQZCQ2bhdanMOJtv9NRSWneGQ7Hd56xz0FDTAfo
T+6aTw+id0Daz4iB7qt20vZZ/d4X/NZy7RqFUzJ6QYQVNCtg7uafu8WQ+6M6OaBS
xP5PNja1uOTUb7gXsgd/5N+vx+IAXqL3XekMppA/vGIgGtJrsgZ48vxNzsUAJ5G6
wcxHOLxH7b8knBI51b8h8VFHi/FVnodvS/Lg6YR7m1W9tv5QCSjsFWYamJbSFeTf
huwTYCky6NHPz80XKPlV6fyzdA8NiRMTRZnHe9Btm9UqjmjlndyrJWsNBsLk+pZg
Mam18gF3ZFyeqTLMkip9B6g4w3KpUkkroWTPyqvjFu6/uiydt+F9BhbHFs1nexcy
pqwlafayRK0BpwbUXduJ/do4TDWChoKx89JU+mlvO8sR5n9Mx3GMR4IRzdhjFd9T
u3s92vMpKKU6r+y/mOCIAwnZRggfuhTj4e6JCnKaaerR7hzS20QEPHY2+G/n4WiN
LY0JhrQlcEoEMFVu7MFhW04t7tRyUdBKva5XdMof72ygIGPebUUkHMumJBGveUPf
rw+NYHjFPdVVLSj+YtJDK1epYYKrk1x/v2PLbK0TOdbMn0/y51G7cd+q/2ywVm9k
wQQ2uB9sBIWWb5kYWIylleh4267rkzfngQQ1fBMYFRKjrrm04qf3lLqO7r3e1GrR
pyij2AwW9CzVg9ScZvIEPgn9o7YLGkwF0tnkP50lK2Ta9IGicvzviQMT5BESfdCk
tNwnG5JbmdwKBtMLfWwdsXH5H5FxNCPW+u1wECGRP3CFBD2o7yJSaoLQZYiLqgC/
AoR18UlMGuovrIEN9QZFnDFk3/0nWyX81xxpN1hEt27Ht1lZ7amT4i4rdP1LEJIF
j0tGEprfQs/BFPRXktvAO2WuA6cdkON9vYRk30zcA2sGMR4VBZSxQNSvmEbsDdoB
BmuPDcSPFB5u6XdFS7D9L6TpTDxGeP+dyB+5VCV+WyGueR7ogvrzTSFgvXbvDPxE
3t/bFGeaiIASi+fZ8Fv1Z7peF8LXU/c53L01qYE0LQktDZ8tHcYY1dhO4/3pILW3
RWubZ2TTwK2X8CIFm6eAIhGv37sqnN5T0UwTH3KJJZv4Ni8RxzdvJe8INh+BjMEc
xZB/Npc6U8JaKRbzOq7uOHbtfe6ENUme6K9DJj8MSkDh5BVkhCNhPYwN31RAQ63q
YALLkRps8HZFtcfWtdXTxtu9BIdvTHOO4cd1E2M1W8tcA15BjPb4J5ASvZvVub2l
6E7bQGhM/xh6OVGg44KInfSrEAR3b9DT6MNMrmQh+NZD5ZV02sDBe7OVvsxld/Wx
QOq8RFpidRs8lapOhgQMPfeviByHRNhzqKEnELe7LaWAj27gE7zmnt6EW6I4oy0u
NF2eiljt/YlymfiMPOya/Oxmt2i33NXMnmQuB2+QQFWa/AaafAhTWOzgUYEikr2D
R8e/auzrNNAb4BK9IRkWB2OKwLi+jLOXNJWoDpE2BTbLo18LvgMtVpoA5awEchEL
yzSP0EN6jB8zMTklFi5uq3K8J76ajGnezK4+OS6Sq91DRUNHt0gOfRqZrQVZERzp
n2t/3Ls8zE6nmKbsYRhar5UAir2LIbST77apQ+kWwqQkbno5c2OPOXZOe/PnIHvK
KB567C5cOVJwr9g53BjfOrhKghRNFiWCvXIrDXQ0e3LnJ3WWhu1KiwcV1O8D5ssz
FEFDX33iP0bsGl8sOyA4hYoqzC+Zi17OnAzfuawjIODPhGAmegvxCro+Ikv8D+QN
ZtqDhWZxSeofcrwuBnHudjH10C/Vi1CrVC1SKrClDWu0kQ1zViOGHlfGAM4OdiIn
yV6ZRbaDdgTgeq7FrTNZ9fvINYFgelsAEnfx+fPgSjkiGOzdBwiZAaA4RzBQNBLW
hEux9K13S93FMrHvM2MZDfLqnl+ZW1DUj/mwnuPtG9IR/scZrCo8nwnR3Td13Tn9
KLg7stmMraaK+i/Q/V9oE6I44LUB8uJhTApa7MKhpgvl397i+eXIY9h2WJu8dPkb
9W6NYH4z6iKSkaUf1ALk8HzLVZsKo/ZtnPIE7WkzhswDPYZQ9ILWBiDvN4p+M6B9
z4XBytgF+gsCcACFynuNV/0hkaqEfKfTOiy4pyda/YjlLbWOXrH08bCGDB5c7h0X
+ZnsqtceM62UBvzk9sZ9IKBJ5Z9pwmZDCXys2zzX7h3pChnX/mRcGdOVOAvQjC39
GGGW5hk8PWG5SO34rNzHS29yK/f/EjX2zAxOfOLyCUZPzqa/cO1jEKyHkoz2z/Hd
lbDFdVH+ynBcrGqcXaAF1xTK0yxEvpFJTmRahVoQ2VYxa6ZgK3qVKdyUib+N4sjW
QR0KN8V/OPiUN/iu0Z9xpE2J/Pw4KOYMlwaRa5Xp9n5SUFpV78dUsepLreLvhhHz
UQ0lly9N9+TWQmiTAY4ZyoX/1nCQ/huOS9YkCM2ellNYZqjw7iLxA+dvDVRoNrRR
6MmmZ5zldDTkj1/zoPFJcPSlt9hpqQGWEH9/zeq8RgWwUClQrvE8kHAoYrghLIWU
hF+wRoJRJ5DHMjW98ZrYU1hObCwsEBAcaEIHQ7SIld/PFLlSByrHqGO9l9tMW/ft
NmBdymBLWTTA2d0cpr6szukIL+LU6wrRebBqiigYycGl/l0wegX3WTzyy1hcH5he
T1bTYQ+Zcqk8TcEYFDBTU5MOIS5FDiXRHSLbzdUBcfLaAeX3r/xg2wldphZUh5Sl
rlgLZSi7OlswN+gIDq6oFso8g9DMVc2OQC4NI9Vzi3fc6f6h7SibhzilpKqI+g7U
Yp/Ma78XngskrE0khBczEluS8OFbfPNiJC2C9WmaBsEjU3hsI7LaeJ0o5LBf6Upo
B4tj+q9RFo1Y9fqe2JlpbMkug8/7M8RBHbfletrogMAguIvnareSJl4eagkb9Rdg
KrZbxFdA/tsRkJrutdDhhB8qwKR2Q6mKyxQcTRlxWkWiz5zTTXVbEU73U+dKQBRU
oXzRCGt7d8KyzlRqbI2e5cvc+SxuXcIFdWaoqQvAundNxQwMOKFxpv2nEvjKqWbs
6BBHBUPSZBgXqJE8bDub5CG8VkzQxXDKPYImcaTJOJ+OzESvftDu0TmxvOpTtLrh
zQScL/DUvkacqvIlEJ/tozwp+RrF5nNZT9D0FMeYromPjZ4w4GrwiUuqrUbdSfDL
kH0Cn6FhgHsYjyLJFkUyr93M9+5eT4zW1WotwmNkDv6qy72pzf19z/hrBxni7EfQ
zUDdzBL3fAnQQ2IkTw+NC/i/KsocIy7anJKQG3rqE9lqOOKYfTgho5krm6P6GFba
S7H15jIwbgECowkLctlKWnCvJcjY5Ckvr8kSk0QMLjklt24f5Jgtr9o90uJWGoe+
l3ZqZyoIb8jP0W+Duh0ZPGZOv8F+ikGYxzAO4c4m/nyA4dvm3ijVau7tswoJ6wa2
r8LgIJQteY9j5SbObSvgOWKdljJW/uOb/Z/q3oY/KrhB9mI1+ZGUhJ8m4oFALyAk
bVis/YAgjW2S40fXcuVKDpl2dd8EIbSzooZu4ZxP8IhCdO1Xhqh8Pm5pukR0vRnB
p1hLFDLDiEvBOov00wrmfxntMNqBFGuYy6TC7x6Fkjmaahj0uFg9k/vjr36Ahp/A
fy+wU6fqmimGdYXZUi5OyNeY0Q8ecbeIO5AnpkqKPATKzDLLTzNzjGs3iS7p3y28
mdSa1g0wykPfkeApd9HyvQPY2JIWkLXKrOi9uZHmAKapwi5pkJSpHP1qw+bf0tMI
YsPD9LY5EzKmCQ/nKJP+l331kR4fsZt4tn+u32RQK31kDd1OLJ3mQcoqntuOOM9M
8bGcVZ8DsjcTqz0maUn7njAvGFrByNaIcJ6GfhFyMJ9PSg/ugipyBQBTIut9iAqc
DBWYr399L48wsgsUfWXFR6ouNhN91T7qWzgpQd0LesOOz0mlWHSqcG8tgE36cN8S
Oii3YwEDcXbrC8orRTsyR5AFj78VNP9Ppk+gI2DKQF6VDdfBr36AMN3E6+ABnJnN
Bue80FpqDvcCfirlFiyw7IgRpF2axrf58UDsQNDvsv0oPiDAsQ4gqh+O4qVVPZOS
/1yzn+uh7kCJV8ZL/mGYlhlyn/KNzaPtbVXYt2OK1STRj+nXHdIXg89GvTy1j7uN
g9dSyij9fo05yyGwCfhA32drHsWBffbgsHohBvQ1AfNruwQqewSaTswcL9Cg3h/k
3M9Bi6tUH6e+xRuaSfj1BGIaB1Lru4R+fFRGzBlsAoqPB/jeLlMz3AzcREXAVeBZ
8VvQe0ADqeI0CcgsWhvCTezQWK1X/OGnqX1m3vJSFQL6c7vh1kshIjdk1rV+oGZd
+o7bVX13Nes5MJTHm6l+U4v+RQ6X5zLkB67wyBtACWM9CHZUxuzSzh4H5v0tCoMh
FJH0SQg390ywKztnaghX3XQj1AtzAqWtwoKN42/u5IGveO1bue3ItzYlyQ38N/Hg
MRoUYB3crsZVrcQ6DuiMA2lTAo+daDjt/ZvIaMj6ZuNUseHi4qPK2r3aOPb769GB
fx8zkOGqsqVCUUqa3OTjd2N/nc9Ml0cjlwibKjNUzsuAnXTHVaUwCjGBP1djF8/d
Fee/UR9rOVAoTy9Pz2jR3VjtxAKeOMr/AahIIBZHodxPGEnkFOCUR7X5J6rcsvFR
8RzVK5c2V6e5HgHAJzEbJVY/NmzKXzW7mosg8Rx1SOqifH6YgPN4FYlvruh2wF5V
ttS9ZnDlWLe6sMKOSxTEWGs/TM600v21Fo2woBM6rJxTUHtA3C/W+IY17O+7Yd8i
BZ62jTUkNGhuUkLp7iUuIcz0F3r5Zpe5jiJXXeTkUb6cJax55zzdgrTATJRYLOKh
SzcgPMBn9PjnrTjtB0Xv9dQpNjL/72Wl2uJgcKbehuFAycaY+UcegrZAkw6NPE/t
YXu1tuvxp+1qZ2lI0/a8opM5K9vYeM8+0V7N2AhtWbxPLoEvERtwh+Ti0YyP/7Qn
8BCJUabf1gwAIRVqaEFCFj8gGfSFO+x06SgiCpNMJ2nkTttCahimg12GKGyH7T7g
/pubHx4HVhhW1N60GzpbK0U++0gFwGhI5/4aMyW/q3PxKWK4WTVegqEG7LKaQP/4
RqZLGtJvamTFDvX8sjYRUeuCCA8pzudqZDJ+CBvtWCR78Uv2tXpHOlnXz6P7bRgm
xONwLc5XHzuJvhLTYG2VJzqe2+x7dsf3sSlQ6JOKgy2cr8pLK2bZDPSb1UzLkSf7
jCX5cucMGemm+yydRKnD5idSYqrn7qgOZ4vOkxECAoKtUYQBkc5GiGxR//5s5fB8
e7TMjSYHs1kvQZMA6qO1R8qZ5N0CjhhWiP63b7KYmwiox6gXcDwGr98joUxanb2v
weExMKBo9DVCccUVHYWIe0XSYdqdkK+LGxUPFbmlylZEHnDs2H+5P+6Lnu/0io7N
knFgELaChVRDtyH03Oo1Id9BLrXhL8NKM+01ib7fKjFDteZoyIfXGhqoLHoAJoXa
ahd1xfxJ8sXcGRktyethVFSqIUsmHFsnC2TXoLOr9P7iSwrHmZYjTKGuyH1C19f3
xEFYPgiZO9nJTSGqt5Gg7vjZ2IQyykJXLBFdop9R2WMag4F5IaEYemRw5Sxqix7i
GBa2d68n7ySzI++FIFsAoZtPFvdt0gtOtm87wxsXLmJkbncsHdnoYeWTSDainN2y
378CzUvxlAQQRE+XeAnL6/F+Cy8uHdl4SzXiSJqRNVZYOZLovp6qKU97uaQ8Jed4
956QUiPjGVMqO83VAXU0J+GzSN4q9bCMJ51OaHVHBJU2xjJ8zW2u0/l6w8Bv2Y7u
o6pvMcLF9/VKPr9m+UihCSL+xlJmG6k3OYohvbV7twog+r4tzN3A0CXsiZssVhPe
+oau6WGeb5+hwodOIb2Ii+3Dp3bZSYAgqmIO1ZjYFx3dY9chr0YV6r4mkODq8eF8
pGFkp+fpOvZFZt9uoRNSFK8892p5n0wmT5iAyc22LXnLR9veAe4frRfMWtxFGPly
dNh9WC3maLAYT81XYY9OsKYAuWLGyEzdgNeImZFpN8+vOmsrL7oGx7047GfkHneP
gzkYcVZBY2NfpeDNtnL5hayFZg+qRL5mwM/81gQ1mAysBAxWF1x4KwnRkZGNY/nc
wPYb2xsjuED0YLkWTysbX8RQtT5oCoiNAxELjPFXBtXtvkbDZkQoclwM0nGDrqYj
G3vkEn9pGyAAwPLMefGWXbFdKKjm3tAARczmLqsNYCHkpfKuPB9N1EPZY5bSAtXJ
bD5wBgtzvA9iY8+V6Wl01VPAgnC9dKBhULVJtiOv6lCvHIiPUMhMPPKlLEM1gjah
Yr196TBWKAdLDa/rfGeZTEMuxTjHq/MQ22y6kx1jsE67s2EBwAi6XtRTspMqTBCJ
V7UXKjNv6VthScHqzCNPuX093WoZeiWFYKHyUek+hHAJACpeLmS6r2/S8LYjrnvU
mdSamy1KRtDW4Vy0iOhb8U4KDS1kTNZTPGNPH9cSd9bdy5oiwtTtlOLLg5tqEs19
wSKTZnWxNdQZD1K8rzcT41iJgrTDT0IPn3uL7+upaH98FYoXRpEZ4n8A2EIrSkaM
xovP1AVYWjU85C08LkZMAoklSGMRKtmJnxl6eS0LWi2DZt0OncV0KsE26lDBSyDu
XYvRHGAudLoKJEqo2PWgLSk9VUdQV8B/WEoasYnAiRTFVpWIRf9zvj0ST/wCeN6c
VYxqjuW+hgNaSB+Y8bEpNPBqcl6HRNuynugLPpFoYgnLIiqB8zBpfYCoa7I3wCJ4
S+ne+dk4u4I/xMo73JK9Z50oAxxLSKB3XiNtNnjJbbHwu6aGwm69NYh7zqWtbZ2n
pe47xTeLjxOpzjXWCQ2V10rSZ4gRDELf+fWTt8MTVErP2QmUi5j4MnbPw/LRHSot
EY2DpumCd6FWHedQDUF4hx0Le7VK2i3lV040k+WW0BYM80qelyNktRM/psirhduq
0wkeiyHUVYZzCUSGxE1U5rWvHS2IgobgZp6GU+IzHj7QdtlJqj6WIWzvHfBJJJIj
Cs82Znab+J6lguxSEN270dPNLo+1qfrMFzCcZZ9V4Bsoh6tIAeULBQ8AL5F7gEH3
byarVnazIJy5pf2Y7G7k2R9iGHyZ8QsmR3lXEKQh8OoAPXF+iKFV0ADHRJ+r0gUj
keAsdmBg37isd/ztPlDNnWRw1sxfTr2IwaHRl4ZIcpo1VnNcXENUlAA5LWmROAey
qMF42xyZM+DiygEP2ziHPgXs7NEnbLVOtgmweJ0x/2RBfPl1lBvmmkAvpHNKDhUK
VOVkdGKYd4v8D67nVeN1g/6doF7K8R5GZP84ON3IiIoaSmLci0A/LCWvRYGrK0oT
3/VF80DxGBACLYq0LaBS4VptPssjt2Aa8MhnryjFvgp06G7WTaDvm41XuWte8U0e
4NHoAVXETpPy774qzWfcTaNhDgkcFTG6kCsY+ahF7pGg6v+HwUT07f/YyuF4vKFU
5gv6RkPSNjQYP/S4d0J4dpyuN3y+0xlCAWch9ngWAI9znxqtMMgwvWYY13K2c3RB
qbnvgbKYI8C0mzcRuM/8JxsNHFkq2Ay+7GzBB+4xGiXIGTnOeLUChtBZGgxC8t5B
aefw9JzN2ist0bA1by+QgrVc/l7IkY70MQ/W3oxV0Yp1tR1eRJ6nR6KvjAsKkiJm
t5r9kmG6eBtevBKx6jBOul5f22c28j7HWzRL2qe6K+NYu2FAYv989rKXmYNggjHe
8zrn5muTG+PK1GXON/tUVOifADEq9lo8PRpZI6KhFWAb2dm/RtUTQj8OgOkiSdar
LueV1kFavSWnPqjdZFoxAL8GkXPqw2a1oW0QTiIzIgcTtOI93TjAOTiu/81OVwcD
8EQn73ky+8IJq3D1T/ifaw+nN3ATOQhwunRPNWh5tx4CwoZ+Et1m0EUd6n1mRqLa
tIelUeVj3EeMwrlO8tvMGAOMzvBmeszU+606J/LZmPBItvrvEospNfabsmnne1w6
6Z4FClePbbKZvmrtT+fEg3uCdG1uOEyIYZbWM5I/aLhdNsr/3JldbsitwObuVYeL
XZ3fUcR9I/C8p/+1Y2OQYx1eQXSD/YFCAKbLaYaK4hxk68rOIGsJyandGKL0EIKC
XUbUzRAB0ke0YtVGYQkVMlb5eGM8fmlzIZuwZCHmJVftsWUPvq9AUKQyIh/Yey7b
vU4kKNE7f6el8z8oHxa0yOOs8mv1Uno1R7r/H+3rTrixzUiBW9CXQSZgbcjyEZE3
lzJ4/ze1lWDDa0JfBBWb5z2Xe3MREObG5iMjGoJKw7kLNkkp2HHJQoC5cfZV7xSZ
izjbYEBq4dni6Y2ahEoWIkhlsI087WxkoNRIcEOXfNVpfolKoxUqLlpQECzLcrcK
CpwfeanLo0a2Xl5iLQuoBeeqK4qArkcpvuZ+j8qwqrgAJFxjezUT2/duAzyETi73
hnHTftSaDAgQ3vGB3/MPicYx44JzdnKA3yl8uuUiYHp1xNpcY2i3wMlPYeBOy30R
beIa2jnz9xgAdDxE/ujQvMLR2Yl1uU8L6wgDDHdzGave4mGO3+H9/LVAKtdOdCRY
R2wvSqXFxKFTVLkwjgOEkDIQP5rzBEoGd5wIRkGL4+ehEySrstmMe69l4yorjUjS
3REBt1PJAIuF32nsEnG7mWF2O3ooiW92qiAAYneYK2QT8dKqMuHLzH4qqVMmBF49
GK5Zum1QjFUbLLyQdyVdJvjnurVa3R+bv2rIeLvzm8nIZE2WL8B7tixvDiwi/ULr
bm4wZNvWgcBdCShiaVdh1VFLjfjXj7f4MeFEfPHOFTL0KLcmUMrtA4vAXN7WPDPd
AnWiWVEi/y7IjC4j/uyWAguSkixSThHZqnRXn3RpTm+E5RZOwWMK8vkloBN4jz+O
HoDcVFtQb6IEOusOhopYM5BsdgRkINrUwTLX661FBqGUNT6lPUNci7qYu+V7o2A8
6l/UFEzNJdNtBixUkKa7rnBB0pECI6jxCSmT2Vg6YMK7AQ9196oVM500/ml+auwR
nVg0wTmvSzBdjB4yGueY18B4EBYfO9A+x1/UbCYxuB03YijNCi89TCR27EMMyms3
rFGmNV+Kv29GHYqk44DiCnfpOU1q3oBfy0Tm52kuZ6PGjXKj1tlDz1Fij+Pkuyyy
SmDDa8xPzZldw0K/DOlhYE3iwXuYpyWJhFLOkHG1z9gnfqrRElCkm2ks/wI0AcIy
sYMZLcPzqgR1/WqwD6xSVfBU4K7eJi+Q1kd5EVZeKoXKFxJIwxyMCYcHSQXpcK14
LBKqiR94WdmaJRC47Chr93zOmpCK62bzyrGb9fK9vfLUGRpCZtbByUZIoEuwPT+E
a/OiO4/XUomvEhcixDlBiECtXr3GjlqImsYCamMNB/XFVi+uVMSnZV7kgAb3g9oT
xB1pnsUURhDHNZknY75KTwEKddDbfEIH8vX8Otat3uVU3xxeMb3Wq2Whwt1spgxm
wVWa9FLH0f7qf86vtzFp8Ha6oIyh69nYWwFio9MgwRRXTOTADEcKI/yD4PwFtren
WJBdBv/513RUGivDFOC61FjMXUrg/zcDhK2efd1I8XAzWsRJVp9a5c6ZgCR4pX/d
AN1szBhQSiwnaGGRxBBoG0rDI1gbQ8xj34X5hdfZ3loxA1HVQxOBuaRCwQqM8hNo
aPl/55BabN3y7xigEkyFCRNIn89sZc2G7Uur6LMriizUwVibesgljVOswTpJriJe
xY+8IROWk9rLkSttqC8/+ZAdsPkU5a8B54iDN3fQdVnPSYrP+kVWW9NsrQVJ6yBf
XxygmHBQmqTAPEwUlGGab07tHAj5V0sIPLdBR+PoxcX5inxgICCuyib5riPp1Xb2
FLo3CQWNv1cZMyFPYUydhM9ca5AeabsZlfhrwHL+z/5nHZ3PzTePjqWWPqDoJdmo
12YUy7vVY97/eUe04pqmFdEDu3MWIM4PnH/PbXGdUyIt6SnvjmK1QVWbFIKnzrwH
ZwJ9b+tqXpDSj4kZ6D1GNiANdYbpYKww4ZGrf+jYjtWF0I8RLOYZ03XTltP7m9es
uHYhzMK9ptsippmYCb8uFNK0ufPixJX59hYEBJAbwV1JKzkI13zcMblDZklwFeWX
Ot7lGHZ62nZrbvhMUfoiN03Lq2ST4YOgBL0Jobk8vvGO044ahQp9Leh/9Q5tCcdj
tvWuvh8thebGPJ6Hr9r7wb5gqsCVhdcsUKtZB9CNGCQDGQu3Tv0nKscoOvXzd9Hz
5p5MZKxz7krTSSKzbXt+iIvoGxbdPJIDbTxWN1TnwvPrEIOit8rV8XwK6L3eGOnd
HDJTVeoEZmi+m4IRJogFZTOTkWKq3u4STip9xf41pSQk+Ra6lyLgRd5/cavoyrrL
aL+me2t70OCrOrrDIPyT8K6EbeIYUvQvZcSdICMIlNVABGbr6HZ/3E1XBLW90Eu6
7HDOqXJ2y24c5E9A07/azp764almF1ahMQ0kPBzjdu9tWJ3EwJ0crZuPWmfzb0GJ
sB7sXWa17/LV+2mgSzcN9tKuan6jg4y++rcF9n08EjzF1y/i2JX5ijpxJIh6JSVq
b5XZ5+ADxm/SW7Xg+cGWVrT922wajQbvS0TVxglgdhpMK9R+SPr4xocNQo/1Wna3
tzKrp3fA6TS0p0f+1niiZ66ejhJFGnllkm599RlnLPKOeHowCE/dj3N6Ar2YrFC/
vvdey13SXqfEad18cAxX74G5XD2ayZzlbmqMeRsZBPARCJ3lUzIKfxtjzRm31L9r
KjV7bGuLyY6AmATKg4cuTErwf4zpmn5CMQWSG5les7lRM7kt6gMmRiR/BHXVzxFo
EZJ0SdVbdkMr1JcnXAnWixRH0OUREG7BnESjpa0/4hj7bR9pANTyOyuyouEQd2Q/
8EzWjK05Q3qN2VeFtfbptXX8Dsj2ggVvQ6lMViqmh+kNYZd2kBSR3VSjpMe591Dv
nEyMj4JL76hW7Habx3xQRnWId/PnEfAe0tv+hN+7Hwql1/MUJMX+anvQ3f8EBgI4
fRRfcL1Raj28Qx0gU9nxYZN47/tt6/ZWBp2IA9g9pYI+mgygHMyyGNcfANPRjndT
z/GWm/rte1vSMyG8i/jRpBAdlWYHZiMemsTk5HsyXKrrRYcCT/sKZHLmaZIpdV6c
Fe+1p0+nxa7e+FL0i/Fu2MSH1kn3Bn/YT3cHauziFjQj+vowgnW4dME66+GH2Dur
HRIIxtMwH1vNyAEm67WQnZssOpI8ukvlHOXQBv2LPj3els965Uj0KUp2zH1rQRqD
pE1R/16wfxYV4tg18t2nA+dUBciLLzPoXFbBYs5dGVn8sBEIwC4lWeLycBuAFlHB
Gj7uFhzoUh6cUaPl/HJa2fEebR8u66B+Y64b1m8pb3o4w37DyisheTOKWPxH4xOG
X2mOT0i7S9Euap9ZhMH+oWcNu/rQNtWWYoZIZMD1HvkEjbGtI0s3Sc+dceFM6QK5
CdB2UdA/hYTv4KvwwiBQC8jtsXkZ08n8yEZxWmkZ75NbdFX//M73x/ZGLgJIjGb6
CTHlK/RZBXwZjshL/ZmTJYUcJ+K+vGlu9zAvDYrHcQfp2LQ6H3FbN77rzNeK6+Mi
y+rrLInbL1aypItdhW0N8lHF6sFKTwN2X2r9fCUigijk2UAt3Uat0v0cQhCbiUay
YnvtXTJlIkNfJdLAfXXrK0ckezO9Lfgw3bXKY2HJaPSVsMizLy0RKmAIXfvYo0SG
Geryt0ajqvfDCsIGUL9LuDeXBt6aXKWJ3at0SLcKY2zZags5De0rAiaGNf6XXYYU
m/N0kFAYT7G1k2VqgDhLYvEbcUabn1oVTB5xI62vsMI+2dJC8iZ/vUp9pLg+udQd
ZlMowPuQUy4sMMNI3+FP5lNGZaREgwDOMVztCGAveG90xg2spgIbX7HUrWBoFvE1
DMmF/8/bcBUyaq0V+AeEIzM8vxjnl7Cl2QEEojUu2O57LffUEJv1L95yhhoZFbag
Rr3iyRiHTCx88yT0kfzdS2p0VNzDK1WhD0mutAsuox3Y2a0+dfzWtWSzIAsZ+91T
xc6pzTuaSRkjayrLLkFZQaVV9Gaaj46zSQa5CjpRzlly+oXEEPyZRu7LLefZKF66
dMsIdCyvZYN/vduv4uD2Az2t23iumiWxzfiIWE0hI0AfJzSrpoMXvIT4kM6Xw+Jo
PcZose8zp/0FkuiAIMBtgvRT7jYjPOzhXQaln+OYLYR4k3ZzRxjOH+mKmdhljZJd
JzbXkLxuW8kkdBChpZojZ7zEQ3lbbEGWoqakr+v8BHvzEJEEiKsaQIdCZKS5bJRp
vW+18pNVcbANK0hnIw65U/dsXrNKmjqcv2jJi/0m1r5baAEqTI83faRfpkMIjuqI
IIrSgdHTXBz2b4mI9AZzMKGX1DE8GsXvTFiCuIOVW1fhH+vghJvqXfcJQf/xEdw5
Evycbt8sujtBkvVz5crUFsQ8EF4hRhBQrNIYkVTh5WEsXfsuzrTmq44qLAL8nzWz
RxVio0pU2XZh2182pmv7OZjAORzM3RjwSTQx2crze+bO+ZAnTWDGC5jS5Z3lVI0M
yJOlYgSEw9mKtFNYv6EXD1uzJArexrsbBj8OXah5bOmw+1aJNHRwUOAJgPjeG3WS
lkSDD27ROSWUNG8dRiEIKlKGph4rLUIMgXl9lng1EyS2BdtPvk4A/ximDC0pDGQ1
8DA5AJhVGaefrousYjbFQ207lD0221YyDHl/qSgHuhNee2xljiRNI5dyPXEqNNmi
YUgePvRol0aZ6BX67MoAl/Oz51OOh4XgTTQokY48fYp2yP0ceuv0CO5cotJEHbI3
utSrLAJRg6VBeeHmgQQFjg/muK/CAkg3/N8Fs9CiJGJrj9DO2VpK5aBLsYTKq6+x
OZZ5hoJnj8RAVJPuvZRTzrbnoQ3yMCGbXhJ7ZAL1lJZz0bjzkYjeb6bMtxRJWzz3
zd0RrUkWND5uhPNbcm+RxYeAHir/ZkC5ZfMMnrYojhF2UZLIsbua4OXG5uoayJdM
a02hOaFXbTJRm51cmh6JcjisOO4lYzPnApU3XV9KSKRCRuuMyAKPIFK4qLUXzPUu
ad9uV3Frt/ypCcB5+a+Fll7yHDrkhkuGROLvT7h++huwgto1er3yy+oMNR1d0iYL
EbcWHj77FCIjetXbIq5FdHq/9hioRurnZ9PQWh4YGjvOgZQ8fOMZwqKKAkojc6jJ
tInIKadu+pFVJ+tAp02/GDzGGbZl8LFGbAWUSfg8mr9ZMqNAfPZJnUK49xa/skR+
8rKPKZghx5G0XxtZI78awA3rE2lP5v6dR+pBbdhy9tUswmhU7UwBijgDBIbjNUd4
RTFXdatMTHT6BbbxjAgeqTNveIZ7gK/SoRv1QiMnMjVl37tqUPcbDZEXbmd1tCC5
RpPQH4HJDtqDdkP/JtTgoj8AxGU3OqpHGvkojNT5AFElBvuHUPIuXvSbquKD/GCg
15aV9Q4EFjBuPIVktRuCjLxZDZMQ5DDy2JY76uFvMi+ApvRlDDr1upjL2HwkAbAn
5cZCmOpazsYGVtg6DitTe3YxtTKIm3pIgQQhESmT4QL5Bp8s4JsY4PK+jZWlJWiN
/cffhjjwSJRibfReATgGvOMusasJBq3mKKHiGLmydscpEp3vFjVkaTe+R1IpkfY/
4i4MBzM+BVwH/YgHgA4N58qWXmxpU6WSKOfSFqJvFYSp/26V+cA/IoBdFa4P7nRq
0os3wNIjcbvTW+8eaybm8HiKljejJgQ8Oe2ZNEyZ4VFHeNzqJH5fJb9BqMqI6W8w
0+EbI4EStRIYS1FZ4LWvJqkjLDxTrKZxtZej7wuwomg/TGXcANOhIrs9GSIhZcYi
vSk10Fo4gaWfz8ztD+w6fwwxqonTu+G+88rSCACrzjnxsmxfEiAL/VfIZ+t9cyUN
otCHgcYWd/O+trV+46v3/yPoEDOfnCQtSNnZ63ai/xRkAZBhYvTJ32VUX6iIkvOc
oNMwQlXNrxwOIpr61DebLnLdkzmMsrbvEGW6rsy3TnS0qKlmhTi5bNcCPR6KJDx7
TXq46tNuWqTDkAXiv1iwzVIZ5H4QJuKgd85i+AwQVUBGZ+67HvX5jX6VsGmpiPdo
XAUYUdN0hBO+YF1PJSVotByvPF2GMQYFy/RRYsICVHoI3jGryg9IxxaX59U+kmIh
H7gSuU2i6xPVb///WHhbX3ULf1IWHhniO5e4AerGFNAbc1l9cG8t6PwSsNH2UGz4
LNJnGN27DkSJf3XzJUK7eD4aZU7dtEJGRxeq5ryeorZ14bnaLxCW9i009jy3/fwW
ANEeFKVAQwBDJgAet/m6Wex8z5zIiRYuWeUAIZgd4CXP9NY+HVKeSfcqMP7clz9B
vOp2v/lDvhLC7XvaBOyS7sLmkFZPX4hcBzSVvj4Qmy88WsnF4B7rqdSQwimCn1xp
KzN4TNfWM4w7cYN35iFicfE48pUFIjNnDrr0SSoT34/9JGaZ8xH6Sqbi40WQaLqF
gIKlBMKolHeuOBvL5SiP663EQvP8S5ZSzAFMYjqVuz272MhinJQ2D3+GdSCzOTWV
Sdpzjnl3MUdyAULnaWQQ36bu3UHKlHZ2gFnfw1DGS7HiHmV44xR170/GrrjcLk4C
C8YA2+DYDQC9AIc+UgDM8fFqHRgoYMWOXtX/A+jY9dtRvGvWZijwpMnmnCzp5Uso
TAf/UlADsISpVKqjAE60+86dzYXb0hlNKnbatrW+i7idDVNuQ8wvrxMCJ42pdtYv
Gk5NBez6w1sdM/+9Q8GtJHqf7fFvs7Q4IpM/cjoz0987XMcPs59nHxMIjYMCyu6B
QntnL6IBy9W1a61rG8xEibvT9eeJQRZwYc7ZqWQxtO1VkAwR+HwLDDW4ByF6cGNn
qW7W03XAmZ1n7OIVgfTqcyGBVHJtgOwN44WQV/iSGijlIc1rzonR5I6IzFDL2rMr
R+vrKC7nwMI7mP08/ZJLrg2vPPTvVdEd1P40iDqmQd/R/KNrG9WByNfem3Ieq96v
I6eEQGFfCWKOpspxmM8jpTMjRNcw3mOidpkVCIG1utqi8auVZIfIl6Rrm1laCDfd
fTkKTsw9TkewO4KRXu2VeAzDLG2E+3HCso41yFqYFW3E/tHbnXPxsjiBHrUeu+sU
O+49AImi3Wpp30CFlWIdydVYlJl/WI4fvhG/ZdW3Tg41K0Q8wO1QtzDlk9l08jkW
qGXgS6K1XxnT7WtF3ZdLUJUIQa8tPIg2cCZ9QUjy4Ak3zG2YvbxxT+DRrdAEXMZy
mg8BAi0lKc6IyfABYtTmCS2sisTnPapPjfwOzmXhLfHX+m4L2pTOW9XrF7MsGrrE
FzEavPd/XWA4Cc3ZzWhIveci6nUlxvMbPQGP2eNIREA6E95mNxJokWAnyL754JJG
v5tvwL7QVSv4x69OL/U7wKYgzaZFh6XqvKM/q3gmm5psbBI9zizn2G1nNbWTexQt
gPkqTM5G9vNBGPtBMCXqiGIGpLaS2MZO9n21Lls5xKpVIjKIJmSn0Axesa9Cb8Xz
Xrm/+YZhqo7gvJiZNRtYhnvIum0FUR8EDHAy1Ousy1Uyrg8BF5TM0wvKsizA/c7K
lvwS8JvUBQ1WCmQs1dr/BnfiKoo4WgK6mPEQ/mFJS0x90B3HhUOccA3rAUMxdt4x
WWiiy0wwqIUrLXDsJMg4CkczSyj5NhreaoGUZmih0HBFl3EP4TZ9JvSWuMbs/q3Y
76IgkoKLY1OO5ZRMq2Ijsw4KcgyJzk5fxSwLCJ0KZZrcn+dTFL/rpCB6niuUv6Q/
zx6XBE9PFPBiBfoKm1ejvBf5AF+Ngbsmn/bpPoenW9slXqED3KQmSKN46rw+Ws0i
fnOscgewCRZG48N3qVzvrabVWqy7lQqqCGpmR0Z0iuenOFIoNE4feTLkhB5wX4FV
g/lQ8QPdRAqkR1VEBacMFNfs4WP3qIYE+EUJCgQGAZ5S31JGGvfSzWdqEF1DwSON
s5pk0VecnCcg6FUPhTXFKPtwJ5FSUe09eCHhzN+2TDA8VrHnXTJivcUpD4csmzma
4C3+M7n5f1mLv+7tEVjy/PI8nDWhpXRuuxBNajaFHibDLcW7sSyfGiN05kvADBh/
IdsNgkeWdtv2++9J8qQYSfLE3spsJwA9xUXU78GxGt5uKXZQ3QbQAtn2fJMwzu/N
rdfFWkyYPOGIWXkblWThSzvG1luuZtEDxu2d+phWsbfg+Hq805qR5KOpqoYzIaFg
hLn/txFCWRXLdh3hqtneyoQdI8LUP0gh9NgX1JKeVOiDHXCS/5PSFjrAn+SDkNia
iEEdnlBUmFCL8wPTM+UKw0dQjEMeaUXr6ZzMHEOfNAx1RvhuXqBivgePaoJtJMgF
VJATsLptDKSg2IPphQAB1AwyieEsJx2Yer6r11He6Mh1pLCXVkJtVYlqVU59PXdk
tVZAVg/C43gQRrnIwUSotJqkc2qMVTzhcruZu/nx6Pu0e69COzap0wMPL6v8Qdbe
N3MMCgAxh8250WXmCrqaZqFrvJv8J9+MM0DAvc1meFHYCQbMadp+CbO1UOAx7KQT
t3pJVcat5VgjvNFagiUOydxWBzQY5BgEo5wm5NXlpBUJYviuTNWHdnf/4BQ4KKZC
ObiQOlsXh235h+a4uyw77LK3LO4Hq4j3DpdBHGo9HLcrTdlzlkaFNRJJ7g2Bl+lm
Yt4DTRXrN5VDy/GvI6raLzWmd7T0CvFU2yUCoI1Ate4zukExCzOdq8JrJtozAHeN
l0P4+Ygixtr4KsY2poaePnkL8wHcOmsW8p/BnnLB8NP2TOFCtTg5aRqcIRg0EqUO
bppKzcw6Grw1k+2/pye2k6qSpB2Dpe0TYHwggnVjCnmmA31ZQ5pmJQtCu6O6Tvoo
kBSNRTJMhAd0397YOUQJFKp4fI5OmjjA4yWLazbUNrwMD5kovWM1CcpoUC2Q1Axt
FVIAybl3DpM1MquR5O2EmIYTlSDGyLKHCrR4nIQJgpTa+JRNEoFWRp3k6gjqsbvd
38F7zhTQyMKgJOHkRXYCvjSeOFhMC9SXq93SK1d52Ri9weLReuUdcdshPyWRf4Az
EREkltV/3fhSd9sY23IhurtBb9yCO3JkzMsh3/5OMR/UJhZNP/zX7L0sg/bqWpJu
HOwmKRa10KRuwlMb102M70b/icG+mgQRc3GT78YmL3e83EH8zAqGxUDHGM59LmIM
wAmJgB+Q9WW68xo1RQWMJivrJpD4PyV77PcNapm4h6aOkNBPFC6h+SQQV5jERMVU
yeh9C1JbHgWH4/+QxdGo3l1rv4YbPrQIh4JGEcda0VmDkeJfLeRfmXHc+TK+qaWj
Yv1fzFbg0K11u+oGY0h1lbb1YM9fADmJJJlYpM7BS3PWY/Zjs1RCPxPcoWHZUGCz
UpUH2JdsRSicJ8d51DzR6ASm99RQGAEq8V7dy9lm3MDIekivsHJUpsyky1GDNjlV
7TAp2G3wiq/BdPmv0SBD1JGr0Gm/Q3Sc1CRBjo/AFsio6XaAl+U/Dh6B9gdTIAj2
Lf/5VYTVFcHcsNf8UAZHU+KHoAgZq5lz9tOI6s+Sm/+KnLLVb6tV1qmspOibWGcY
NTAUbfJi7MNac+D6Ebls1d3AA4/BgaV3ctEb+FYNJeJpHh1/BLQiIo2BW5jZSurj
rZ2tNqvru8zI0Mgufg74boHsvQD+ere+gZF7cLQO54nJ4FKqBEPaB3LVYRHmuxN3
v/xw2I6wcBNoeBSdIwsyuYIrun9cUe6VTKVWM4B9WJdtA69nw1I+SLaS+pRB2kvp
S+bb+dsFvHj2+TGE7MlSi5AnE50sBl7N4I11enjliAoCGet7zh+QLazgn/7+50gO
FjbdLz9X8xjn1DhSfyLCmsk536b9boPUiKp8hQP74+n5Zp00X5HTmYhcnhmz5cfD
bCD9M+8lXNwC7Vq7lxQ/IX6lKwIy5KhGh8xDldjtJoh2sssp+hGKV+u8weWv9Gtm
SodTHBP544J3IliRtXXhsASGnaLEFG5yoyhbZdoLwRivh2qn3HN3XntzKxWir3/q
JYnt0kwZqkY8bJ9b9owBBMrgYtQlHkA5Tz4yJLHDOFbgOt/BfFFZsy68yXglgkZF
R0biZSXS9nqNArIT7bGhcA40b0gWgEG1y8V3bxYdcL1GmoSl5OwdkEL97viBl5Dc
id07qYTM3zv0X6ghWoechcplqiCsWYHOahtWsV3o1e0d4idU2dPfEgtRXXlcHbTD
tRRQxjKPzntcRgvrFgnfOHJw0iniFk7cSh/mHsV5HBX7llcVL0uXBiVbzcf0zKhL
/ZsMudjvLnnq6S6eywaJtC0e5R407Fi8rCDQLhZeKDX4DshCRNdjo4lB26sdZVe9
x44GpnsyNicUrbXQXmMfm+xcizD4rNmm2mvxAKN/9O5+lN8+bF2GRjJZrzvL4ulg
sjDPFiaWL27qDPqOe7EAe09olS2RWDGGVUcqrAPrCR1n8CiA42TnYRUBMkE9slMT
rrr/+wen/zwVEr5Uz+EjgEjBKlucPQgmVweNHQVlzbzNAMbW7wcoFx5BxVWZ9dy1
SwGkUVdiAqd/GSJFOKUH5+/YEdiAUaGIBQL+g2yTt0pBSzMonUhbcB6vgPMWs9Dl
5Ut0c5bx6UcwlnlaS+MkE+FLpxHR2hKGTwhH/5DLhnUGj4hHaayRhOIDysjpxFLA
bUJaNHbI9GPRdeh8B/YhzWcSCDCZyNjng7dN1k5dZWmOFaMIKJcU3/62KyK2hUet
RtfcazuGy59R2Y/imEoTfSucGnuwdchqrqcclvDeM9vl4mVLMd2DvYhP3wo1gfIt
ZYP0FZv5rNULlHW0POcw73xBHLl3HR3jt8kIaOHqJ2Z/n5H0J3F2B0dfhxYNV8nx
CDTobBx+93Z1h/HWNCksFkzAEhaj3Kj8exTWAUqEbBb23vKUHdArO38Eh90Eau8q
QGz6heTVHGhSMQct5B0+8s//N1yN08oWeRjN8bjtkv8gYwxn7dL0LzAZdjUzAHRn
hkCmAUvPF5YZG7vlwpXxPU4TM4tEx1wxVHy/HwWDXR4gECSatdJN4odh/hUgnrqk
lB62kqFeVgcu/yUa1s6WaOY/Knt5y7gNqFfxRdvut2c+MzyDGrZcPu+1+OMRr6X2
ifp0ZTdcUYTYCUSss9i6xkutXiqZdNif14MEy7lBqTDcLBcept+BOvU5udznZ69c
hNoew5l3gcSLpmkaE2KZ4mmS/1BgAvaQqQl4DpRLAFrbK0PZjGodbffXu5Z8+nQE
eAkd4nhSxGVkTHf2tdECgJ1bb3h33rdBqS1hYm4QLpD6QsunT6/lywjaUMXE1Dzk
RUIc3QHM7512tdCujWlbZXI6S972+mtQPGQdOgEtXTOALPga35bAXt3T55XvfPNU
ARqpqN+CoJSkIXGyfOL8t6D51nG37ZPmORBrcKls/QZlN62md1nzxOm2wB3Y7Wi6
2ll0FdXnmpPQmym5lx7zk0mtkiddxuu2cicU5yUcEGqVH5Z5ik9CJGWlh+WzOB09
TB0kSLnPlV4PA4MV2vRxnOKxVJaYuUJbkCbQW7ShV4+E81QnEP3Upd44OHt88KxX
QNjtpy6KiAKgxTM9Kea4C7sevBRPAC0RHYJcQS4szNLHBB8AxP5L1mhiGgnNh/ct
H5YCGTMQ2VBN/cmIvwtJLVJWVjti/InVGKrLDtRss0+4lSZg2/fRDzVcCWqTqIOG
HJW+tbCvrSLbJshvLjel0Pedrbij7Y7FuVpZW0xPOZj23o0H4FKy1YxCBV/m1Kpl
KS+tdCvAbnu1QVdWPF2RtPpv5oNopPpWABQ2l1ccThG2vxS0BVoIOdWL2GiIv3r3
cNrSYU7Juf1+TOHi2XBp6RW+cutabSx7PNySSeXTrGxNFwhgfTpKEgwohmNTnKiZ
VL/tlV0cIYDX2EhYs6whrjHrnLMHSR8doQ9FjePjbwjN1XfsDJ/PGE4dIyBf+rrv
+XbSZK/rN1tP51utXnSqhLh9IdSinc3jRw+1QfBvpkZu+DrC4RnhwNSiJlqxRiNL
y11xVj8H8mbhIAT4x1RHYXpWh21VkcCpyc4X1zKZns6p2rQLG3efOM8VR5+zpD+S
g/FXw+mJtbg+gcxEQLwxgqDa3XHr+4ga2hnba6jbxWIqQFZ23Cv+4Gacj/8a73T9
wb48zzkpC1KDIBog4arjCpuxnCDQec2du+Ad4qq1Q+uxjpYk4+CeZQt42pR7NZ8i
4eFkFyrZKnhciNad58znrcxgJtdUc/KVlPVysCxmBmoCts8mmggOKpKlJsM87hgd
BKp4se4Ft94swbrHbxj42iCvXswCmGDGK7EkVyYHZAclSCATInhCUvkn5+w9tdv1
T+e+cs43Y8JpHEqFNCtUaQtRbvvMnXMej4jweizVRBbi01f53yn4jGm03dbS+DrW
bkskR46kJfuOmpaEbmFLiYcnganRLD67UV9xZNl101Cjjrmt6NSdAxCH4F1WDtLq
XRwG3nux+Q96BtMfxIH7CE/Moz2XBrpyC4WPlBWLSBVAfkPEl2cK8pW275jig84u
wjOpV6Jc2EBQbi3110ES/4bRi6hSSwiJKENMtWa0bMNLwgrF7TBm72EPXefXhcD/
NN4U+dYt+iNuqaPUDLUjAZfZBhvewVibKHfnMCOvDFHxCcORWvLFwOeN9aD7SA8/
R789mOl1Ng3zqNeLARuS2gA0GyyZT5KS+4r5JAPPVkIWdU2GWSt4UiclYR4u/RNJ
ZeWZTG3gautS6nKzdlv29/nNk5uHeOqUfDzNgmFZfsaoX6BBD7P84BvG+9DiLMGe
RFDPQrsnd002HXIIV25qk69HtlSN/t/v/BmyXY1zMtaMnVtpQkinHZ/r07sgo0zV
4AwCmsGtyDxDsni4D1gX+mrccDs9lN3TiwEdEzBCAunCyVFANCX6YgeQ6jfXmDx9
/pBHKKYJmsM9VyMBcCcrpgcLQxB6GpwmvprxDCwD3+lSkJNWu8cvbziWQ2CnFtZ1
wLYFGGK0sxyMotbq6vh5FcatxjMMAtmm7ftaZ1H27nytOPMzs4MlSgNKmBysdTH2
AsFcT1nOknl42OOI+BMMxALYcv4P3XfAZ2Aio2lAsIM9MmSK5QSyUmVXNen30Q7U
qESZG1DghG1rTJicotJsyG2l39WVS5ojn3vZyHK2UQmSR7N8vbQAWkaws7VOSSgp
XxXqrXTN3bV2trqeY2iI1116Zn2UlPiAfSoruu4SpkUwCSMud8uXRE35zC1Xm3Ua
aGy+GDuUPrsh9Fmy35tZ/plS5eypoi8UU0S0Rx9Df7xH2rJwF56VeQEjZzyvffMr
Ma6XH9qlTxMluEgTU+oMWrwV47MNvun3Dz/hBJ7d878tRfxvcYdxwSBwcwVZ9QCR
cZ1GaZVxXaGA9Pl0kaxXumeMEanhiaQIP6Eikab78569kNLANiz/011MQHX8ju/m
skW41gCHgwVu6X7Nz693YmpyIXD13pfGQfkGkKFRN5fr4BOXvz+mo9zBgA2VI4Ne
+LzMQoFLjvfD2OiSYcX86oNCX/FGp7vylRZnTieipQI2z0EHaSqLNzP8uF/LnES4
yxsOCUni5eG89hWzHLUWNdoRoPE+ieU1aPB0aR5501zeqMfKVM/cOg9nlwvrz5ja
f7qNe7j78X8jLLPA3zzks+NOuWBggnz9PG/DDO1ryF8hbk/ud60/ZCU8DtF24hoE
pwNG1q7jOB35jCIYCtsuHO8VPLxOnb7A/J42KOM9Lg4XJnleL6Y1RILdOxQ1rsYS
tb87xrF4+Hb0OhlusmGVgW/hkOfm/qTshaglKLoW7wzgt/8gw0WFlASIUxhVv/pa
V3kgu8IE0LXEtHKYexl2Bxlk9sBi2K8a3VBV1xYFnqlviHE8mknuHgJoKToWhhst
4vOkrbyU9Imv7ec+XUmMa7oZp681fuFpMlDkogd9gnJ0BPpxKnFWl6c0fY07o/8P
sGAgegm9zdAw2hHmCBSG/+RNBE1zAJefcxBZ6Qllsb3Qd+maMfxuhpsbKwxzxxlq
CMRw4UyGN39/W/muIa2IxWWRsfg4cwYraMxZTClZvFqM0BQchHLsSmt7lPV2bMKz
VtFwUXiEaitSE6/P0NbMfzZusyf/syF4TajYXmFK8CC4/TZghQLR/ZETKY46pdWM
1am6Q+yQcT5fdn/Li9IL2L4GNVKdvfD4ur75cJiYbJAckN29HdpdNqK+Uddv46Qn
sUM0f4IWqzTZaYY645yXTmz/zWHVpbUXpPzeVfS/82qk7Dz7ofx+eKwHz6DcNNcy
gOLL+Jjm7LooRJUzLq/BapOSxTP0VFdNVpKUJ29QKUcfd4TlrlAmxTQkisTBCk0D
eChjIoDE0419G56IKB0nxNUYDoXb+Q6li+HPT3KpAdZyzXT0nKVApLMoT7zIwHbI
pOWlbFQzubvNPuJ2rzUOIpgfw6F3QIwBAOPUPqpQkBhRAbh/TmyRVcPoTJiw7Z/B
WHNSJJRIFtJCef0mdDjFlg14Uu5iyWAgN7CL98NvFaz1AMPFKWR9dNFCgiJ0mTcj
SJhxzebBGZa8Bmu+sn5AwcRUIFAUI7Qhm0CXAN3D0xleumKOReG2Xttf1Bu8nN3e
g7Uy7/MmJ+jIk5sv+0+Ts0Sf6XuSCEOl9XDFtyt/+1K+RX5b0Z3Z7L4QkTZkm3n6
KK9pQjibtuzHR/eabXm7uxoRgfywaymadgENI2cT68PtYRjTccCSO5tEXMrjaR+u
gYDiDeTCJKgFyDhww+MnkRsAQVFWgCTw/TcYuEifrYcqWIdgPOZLBOR+jAlhvxK7
breMFtOYDGr74H6t8FY/6AwKxvAKQJDIJT2uaYW340Eer47yDaDXOWUE9T7HZtEa
wJx0C6bvP3r8it7fHkwxEfnt3kW2JZ+zJoPoSHi49KEEWu+1Uhz+Xhk729xEx5Kx
eLw5P+/8HLutvqhvxw1gVIrdKM8jH2lxDy4DsRSkWH/vwwXoMe1FiMZtnGR3yKXx
fxlPznr6TTc8j91ySkvHvQYXZ+7J3cbKRfpCLUO3gCi8Tz9oA69t0n3L5xiVb98T
Lb/TqCogBL1fQzgLCkiyr/VS6Pb0GcR1l493mJS74/2rRIh4W78KmQSXYhGCCA5J
FjxHhAfu3T9C9mGgEU/1Xla7/AiJDMjEFyp0smEcU6WsZFLg1AwcM+QAX96FGM1V
dLfa5zbwyn8s5utbpexkQG/cPA4rhLhsejRTN3EfFmfRhmUmB4pZNbWquh+bKA7i
Qq4fRgaazgZ28gJU1ToOKqxm/1NuLvmG51gU50Rip0DXF702uX5bJR9ap1nEWW/4
R/bYQb2iRmXUpjxjMb/y6yJ0Q8M/TpkL9bwMLNN5xi/dAm1aPZQolYst1TW1n16R
LMeR5ACvVrQDLskQSiRdHvGCi0xaArD+FGLjlHjopfZWE+x+YkJq7YGZU3xXdZRq
YjJey8VfiNjUmv0zxpKOE2KXk3dBTao0lJEp9OUrqFzehP3bcIvI7u7THFKOst7K
7MtCdL86qJBVuy84MHI+poV73Y0bo6kDtQNJEtm+RGTkiX3Tru9y48Jb8ljm40f4
nAcoEh1ldSfA/kAcpdyGvgSEy48B3xv+ydRplLt9dYNjzsaoXsDQagXWH3UQl8bu
ycla4ezqSgEGvDBtKJ2UJtLOEFCSrZahpr1yiQJTNNwSDJI4e5dOXPt4erlHg5N1
ny/iQxwvO9GGB+r8HGOAfE5tLhGZWponZe96DH3nF3060zyRgcs6t8OKB0+7l4Hr
fs94MvG+N2fieYURv8mxqZfVGhbbzQ007yobGZADJiXzgCu5M3ZcyfW1mTZdwLgT
dDsXoPjdWkY7/vTVIh4K8SFtNn+bbvUg1uYTTfQnC91ZGLA9vnkwx0KrLnNTc2/O
8G9hNlYT54wO/+8HUJ1cfnsWv7CVfOUHCo70scYt4wpgeFlKhk4IWzyf7hdS3wPU
kIZsigFjOhu/c1Eq/oHhm9fB7H7VfUkSQ3j+mu1Ej+7YXwjJ1Geyt2P3e1c6dQno
e0h5hoGK3y6k9/nHA7/aCqoGEGysp6E7iiCj8JYP7iuD0c+ZHpuSzBk4hNvj91Nr
TiR1MsHTHTBO4awD4jwKcOn5h0ImdaIPiBZ4mbnvW3PAAD/50H+78UKaIU9jWhJ7
QFoB1P0hQ7B0SvXR6h6HCLiOIC1+7Imh4Sv7uqULmL007fnDXe62Xq8LEt7RJjn8
P59cldMcYWMAXZ+SFy2kstvzyTP7hf9EX4QLFQ6VVYXhsGDvfzdX5iUv3ty/33V6
sn1T/BLE9qgPvTfjZlrxjLITxw5Bbn7GZmdtk0/H+EEl6RdUdgjWN/76iPCzr9gp
bTSm/azm0a+Dd19YCMs4qYEjPYUvcGufW6mBj3byPxhcHmgnleocNjn1TGWyltAe
44h8Poji4AaracFu4J+gHTijuAN2skz/6hmlVTh19qCv3aYlExJ6iB6vLaJK3i6W
TSa7dniBcgtZWwdFPGMDiw4s+IIN9Ff4trHey7bWgvYdkpeJO3U7jkLaJ2hBu/zy
8AcFNuzIjTvJ3vEgKDlUUM4kFOj7g9AGINvnaZ/Suv4VRlazfadeJjlGiCuUOXGA
6q9TLA2FlLLwH/wzD1z6o4cipumNFjyZOHbCoCm9XVvUyp0MZ6gtUPwz5ufqOLVV
0VpGB+qeT5qHJ/jmhzIm/KTk0MxdEQh8H6r+N0dh+y6RC5VSJz2Lq6K5G56sWxIh
1+g7ollx6d2saAoeXCTgUNArxnK7vlro8LG3VzqG0QOKqZEBw0M/POvavtwKjp2D
nWCA/5ZyN+FYTcKx+UXermIVeyxZnGsPbGqh89W/4BWJkP+7tKe37WUokIji0djb
ttKDhSgFtnCrBNRxJZIDkWxxeKo4urh6N8d+7ODnbne3l1QxnvCbc2868wogOcje
roGyBbdD3opENsdZuF5t+hNnFyw2N0wtGk+TxBimeE7Yp24vnKtddbZT+SUpsTJQ
1MPG1U0v6g8KOrjWpWbZSlvo4ZtF8F1ON3yMIh2jvO19p12Tc2QgBsgGrBUYJl/q
mGIrt68VSayWmtGn56arTZJxnLw3voLKM4GHx4bA1b6Q9m/bymbrIOQ6Y9QWHDQY
Zg6tPY3Z5jQKaxCIH0obv9gyoxJmvp6oHNWH6xFf6TLrbJKpoCSqMJe9xJWkJQt0
mIDOLl+J8jE/RR89uok+jIUp2L9ZhUL8oEQ015VzNfN7W9lZuz3/7GrOl9jQRrC6
ABYw2sqRqz8NdfV6MieeKpkb8g+rJUrQlifjsp8IZJZ5MJKr9jzCwbCSrC7VopGE
igvYXYFKuUlJgkK3NPvqshop/KpiXTayPxhPYfhXf5B2AegCNqwf5QEfasjsc837
KbMsc+XHM4pT5EFnD4AOfOhhWj80YjPXeV0V9QLH9S/q9wzoKVuzUj8//qaVOcpy
fJQmzWlwy0cxPXdbGE9JFo+uxIvvgpERinZqAffqBSq9mCsDbBwNvlDZxcGEKbzW
agx+5/LmaSv30b/jWrfxUKZajEsj/WXRHQMbzHI1MdB4kcr86JjIOVp4Kmf1cHOJ
P9gLiE/r+5WK+NxTWgRK/5HtSzKc8YuERuQZku7L3A5DECiq6fMVfTjDAKBxNGNZ
xidla8tXCp850eiFYP4NTijN51ndACC4h6GuGHwlFbvNa9JsOInm9UBmMNlFIq31
BT0Cwg541iPmYgtlgDno7CAM2Nk12G5FAOi8Et1USsQXpUT3TB+rEvPfsQIShATo
17y8YwiQAASWABdUlifrzuU+nezIUiyurehNWvGotANQBrnshAtqebey3rfUTuOL
CoYTD3aBUcVts7+V6XTKhirpWVe9BqqifFXLrB/5yS5osBUUGSwh7dwubyjDgVDD
xBg6ci5pWkNgfu5cab1E6DJBYFnNxUwDS97U8+ZTux/0GtDkc6ct7qss6meL948C
xdCzODjPq3CA52xTAp+N5qdkzjCu9R+JX3gtE2gJhguOXjVwKX71+LwtbcQ/WJBa
prUdx0t93/idB1W+0V6PNQyvic92vTcdVM78cwPcwbnFuKamY/ZGHwPjXL3MJ82X
oITVOZqg6Lwnop+oj4CvdnQMWM+UQqj9cq1kqEEi9X+ehOmk5fucejvL8gu3WWO4
tJcHt5TNTetzNnh5PNHirKbXUIeSKbzqPLLDtDnYp6Ib6rVQ9IC85aCSo/xuaRWy
APPXxLKzw1IzdsOC4ibkyBfvg1ZVdtzOtldqN0d3GUzl8CLEqyHBpS2tZjnDl72N
rom1fEdMi6rU08RfqXF+xNKm508lCnw/mejfTWTw/OgPOF1GY+QPiTN6UaYlXfCo
zNDMZw/iQMu0wmDjCLMpOAt3TplxGFmlvbky37UVulVz/JwYIrmGekuVoqanLW4J
HjSHq2K/SmfdbIXZHzX4Ie6Wtwxl7uCm5W+CzERPhsB4sWH51dcEIZz58xZxaNlc
erZ9HENb3FvKDh50vrKPgAqsN69V0137cxYcoc5hNitxYRC+Zvz5JrjveX1wma0a
Cjmd8vZ9y40JH5AeGkTHuL9ZFCPunLXvhLYsR9Q0nspVDj5qupcqRWFCbUZ9npgR
yBfgXhUxWxiSQVCLEqfGDcK+pH49e4ezan6tqpetAU2GVsVNZ9cKVrSHQzyDCr8p
dQNF1ttZCbeOaKIrir4AL0UFN+6we/PXBYEWZwY5rHlBljGvynKFDzYQVMcRxaqV
UdSJ097r53RjCTzefNe3c/QVseAuWQwOr6V9kROHWNmJsukPbyVa/zH/0T8crMFL
ZxyD+dg8BS89LUnqKLvrZeu9iTkHRPhpka2N++So95oXiqZUfRUa26teHNFvp+S7
9Ak88pSP2vuGCxfuPYQD6pTGGON2hahLGYFAhRioy8alT86087vP/ZRnWEC8yMms
9t072HSLeYnxkv1YZMSixqDlTuhjMl7RuyKWr5/RIzshIWR0s8KHxsHa3VZVBq9i
iX+DqHUWyluIVyZVelrLjwa5xvFxQkrcUMsvX/LJQAjw6q2vX0RTZOIhF2josZ9+
dVFJFJlw35hV9zPYuz+od8Xxg3GE2q2zFoc1UzUbPqoaLTw1zD3V5tMoNAgIkyaC
+HdAWZvTkMPMKvvTKG6dCPRRfO9RhhgMv8vO06P9gqJ48ydNCKj5D5J+Pw64ygG6
16+/oGnizhGvvDVA488PkVEUklpj4JIp+TeQs3H7gBzIQ89yjEXNmQVz1l8q0KCf
mc3z2VkruG8UtiQok/1ccuRlZKggGLXAfUbSbNi6amXFPWO5pZCbINx1+s3AxF9X
pRWnmNd1A9D3kLA1Te4c78qZEr9wSaUD18hPuO6RGU/0SeA+t4a7+GQeXA9/FpLB
bqeNr2vKvb0cYLXWdCC//oiW/S9RuAkCBuvHUPcraQf5pGTWjWryBXELrzgWpIQv
vFH4QlWb6tPdmKzdPoNyMCEqI5+apaMnxu16kiA8tciMplC9g16oIYntnRgvXEov
sJnni6K0bFBqn2g+3RelMJ0DGLNVFdMujvXkGM0J+zTR9Ud1TaDnkW+vM3kZsIKu
iuHixeb47SuTLQ02kYQ0kjU1ntn0Ya5Pz6A9JCNWEB2dnGc3cplyOflr08y3JIKS
2kGHwPdjdNyn/FCqlfapxn8Qla9ldFeQrcxr7L44YhCh5iFileUN1URm0lX3JD1M
Kp4sK0ML+/ws+6IsZz1+jizNYbVAUJz8WwBvFWMYU2HnGw2iexyex+oA4tfpBePJ
zgJ+Ea44iVIkq8D75FJTh8ms/qzLQGXRRW8TQYpUh7UamqPfFlusWO5XTV6MTw3A
iG37zHmE8cwyO80sdLmedni3XIdC5oHekjgMYJTDJEj5L6lFeEyFhO2UKcJ9QCGc
7lSADIu4U9VIsym0hFftGRDkbD9QveVVkmaNTGxT1ajWRL67jePQ9dqSv4hcjQGz
PUrOJdO0Au5LU9lBJFhzCBq+irRBsSp+wSOrfNSnf8bJTXIXtQyqaqEhi0JPtCPT
lS/eOFDlwkhRnqJn7Rm2lrEv1u0iDHziF/X128vm6mw1Byn3Vq/yvDK7OhX3SeF9
EYVvcTbzxqYYzftFqGHaJkqV6TfLb3ACpZNF7JqR84UFPGsTpU4CcLHIu8LnRTpr
GCVOa/xObeBJXYae/tbyzDPKZ1d8fxnOo702IGkPI3BYBgEs8tLnmaehBKSgt9Kx
cf9xfsgIhYh6yDhW13bFBP2UvQcAZmauzMG+Tuskb6i8lNaQq/EU08KlfcPXDBzk
bHIhKanFUx63qScG1l28CpW/gXWUWX5u9kr2o/P7sGLA2tdXcZNJ9wlczlI/Gi9g
R4YdBHo6LJjxJiVCx4WLCwbCWm49sKX9NuBUOCwnkD2RkCu4EufWLnQ3MICFV307
WA/uvnCJRJIGKGAv6XbkYe2H3IdOta/GFCTB+Vawet8WBPV0GvdkN2fTAjzRaE90
XDqrA82HJf3V8tMuKueA6XzfYsSUdosmowjDxILRL1y0c/9AR3HOw/2YYoWHNoa0
ZFVMeUuUv4hY699Zj1TwMCT0NPmpo7JBEJx6K8bSFzl5Y0tEAw9qcwXEwUcRzF7u
IYbvC4gdDWbwCA+py6D7XwNF+aU1hfnJGMnxSVLKr9P6oacgvrDjUYJDAPqgDhvz
TzFI6IfQpEndSIllpIQS2W7kCZ8UsuMIC//XotzXU+qwhZ/jrwwpgZxIMHQWVMOm
5dTQtr6kMhVF8NNQsEMiUDbbWX3+Kz/zBXxh578tu1wUp6l3Uo8CI+iZ5Dz9ehNM
h4+uaOxd27GeUUPF5muwXymmWBJ5faIfkkpK3CELofYAkVozPTS2FHH26O1PZJ12
K9cH+RcXJZEsVAN6SbvXO+haXWAe+GTDFt/Dm/lj2oPmJK6tOMClGXoKIQhk2Qk/
M/WYLXrhpXofC4LDCcZqhniWul2yAe7F2fh5hFJvPYCzsWxwWO5ngBlNZO+FTWxL
iYnxgRHM8d3h+7kHmqJ74lQqfIn8kUWeW5t9+61jgrlIbC2ymSZGkr6VEC8p0Hee
x9JNkuabOfOkQjaucId/J+KzVKMMqVs0Umpf6xN8WNfZKV4d0jICcFD/lqHnLMbO
zB6lc1UwENMmukd7iC1stNFKaMHJl0ZrFK5LSiaxwZD35TtvB9uxY+LwqPj/jqkB
xMoV7m9HjHpgO+eUfAoB5th3FIV1qoWMfQZV+bvfjZ2BeRa5VbHt3mBCJMA9DcsY
cGBSGAm/G4YrWWJdLNo33TVDmvr9njtR7pLauF02sSWWEeOIVd0q1V+j5O8ceJOq
BQOxU07+1pjyksBVF7sXuYDtraq/40T/KGg9g9taDfmMkL1585ATG596nEFim5mE
2Qq/gFNWtDPP5PFyqxWi8D7EyhYAIOGWkKWvH+khtLUEFpmMOTf8Ku8QUT60mpKL
VAKHlGYTQE3NSzJIYMxqcus3URaYOTqfgRaiVEYIayAJPzvnE84uctWMaTddE0JR
kgYkEYdIaxrQOF1rI9JUmR9SBIXAcXCJ8m8iqR5NxYZ++iWP/YSvhc8a4RtXwkYz
L6KmoqY0kVT2U8o82dUJBaZ75ANoqGoS8D2i3GNArLQA6qGxD/jz5dYYXGuSey4j
d/XflfoZ/cc3BuVRzEi/NxfmQpufCnifhJOZWb/j+hE3CfjyPiPo6xFwNhsX4lfI
Cy/ivFL5HnGCMYljB+XfY+8c5LI1sj5i10j1mY+l8uOI88dnB3Gv9h6POLoaIIkd
CelNeB77Dv4pA+DDQ/qGeCFhB8QIo4bsUMC/NNP5xk2HlQ2nTkG1U1bZqNG8SiPx
kLTAwd/XLUnUox3Tyk4Bl9opR2ZU74HT29UAhWx9r0dpD3q/Tq+bmq9ILOM1PLLR
fZo4Ylvg6c6hFApYbvNdgaVjmCegMz4QbdHGO/qCOSl92j3zVqe5z05goCAXhXkV
iZtMkRXMz7pYtQjAJIuoEyVhvWnBgm3qbBJE+kyz9wZk7uVms4K3HZnPO1EzxKgM
o3aqGiT19uYmrsuu/oimLFYutsXANItokCSBAPRmiN3aL2HqVCinBqCy/MJK4xMJ
SHQ2qSCkn1TZ+/JFwyeKrGxlyz5u8jKZensKMei7cNy7wFuSQK8Gho0FpvqG3eJW
PVlYWjsljUkTQ2msGUeC1wGN9ntj9S6K+ksJotVwFpEUMucPbO722CtNf37cSh42
wD09l0+Q38mv7iItobeKQ8vWqXpd5SAlNEYG2cVd4MT9cEm6hJ8C6Q4AkGoIRJQC
9oVDRGWxAPoJNpKw6L8TiAoCYi26t71Vgr0PGhrOJBQtQk0Z6lEBGmcJ+7nC9gNa
pchgZFsL9feDIBjORDfy5tO+OwRvAfpeOsR8tuGSM0A8IA0FWb0Sp/bOOjip9DxY
4UsicN6qbjSreKUUCSWY/gIk2+diBtY8ZL32epQ8DI5HyabndbRKHgpPeShcwh1b
5oMISgNSwA/fpJFf+VOptCguCm75HTPJD44ur2KzhxnPs0RXgzQD5b+ToEretsQG
1pNIv0YGaTJljYtme2aCJpj1dL8kz6zJ6s7bAFIdPRY4/mnVBDrzl/yPnBwVzNPI
iSOGlP5c8B+KInJT3lfIYWGpyKXPK6ImT9UKv1SDCmNrJ2MlDMATZwayx6xI8xJC
J6riuzmmoM5PSMQWJuV/MXnSXSy2OpDHTDmXRURjhBjCnEM9pHP0M3LWcxcitFwU
0OK30MHGf6hDJGMlBPqMpShFy7AFCjJcT2OtLR7FKvVi7lq8ABkPTlVmAl46DNn6
4tqgZ4K2DP57QqONcg1DAVInDtHNr+1275bfusUnYOcnsIVHFonLllGz4SIWdqhJ
8G2r5wwDwyvcbzEsaSLaaIeDD2AkQVARnKRB1sLnQlyEczVzSNPH4Vtk1khxcTGe
nm4OGFapOUzIumLAoCCKs4xlYtWHaFg2CNdmxeM3SxuKNMJg+7ov3vJT9+uatqSS
890gaxzqGDWu5QaMDpGsTcCv8xbk8hlzVE3P/PbFgfLHvD9qfD1jArcGZvuiZJoj
EwfL4dZlLgEogqaZnEY61clMW2GbYOerYLnGtjYWSGmMHoHX4FRUH71MdV3xclkM
LqTHYqPQTAYUO9u/2MuQ8JmFV5CoFoM57ZiSlc610yeEYJuS744m6s4bbE8cxe6h
+vYqF1ayb0DwYIz61OKFrcEs0euLMLvpZUFj6UVUpYmGXYmfI9+AlfG3njs88NpM
7dDKTLp4lceS+Tvqnk5sMbwE9gZYqSeqBEjcwJ449XrF543gx5iU8H2Bdej7Tb1z
zbQUwdax5J0UYfjUrLAKCsIILxZdpOnGAF8PQoJS61+na+r20WbBeX708YcSXg0X
ToVNAqgMnbtDWyrYe+cCRrd3cTVDBRCCeXN20CM2NJSJpvxM2NwYppnRC3AbeyVN
s2hbjW0KZ/JyD3l3Oj9FLvv0gXPtp74dI7v4hS9LR1uuQYVFGmx/TJ81BHKow56q
snWAht1tpRtK2+1iOkeRE98IWUgu0Sv7L9SQfOmMyryCJs9+WcjUVM99MUqOPm9K
7VMM7aoqpk/EZn/boNJm9oyv28WcqDrQgoWKspkEfY6tVGl6phHGBtFqvOJwgWGc
c0ZVsfIuQkIwQhJ5909y3X1/nUSXdRZFIM6K1pywt2BBLyONiBTi8IKdx19DEDH5
t1VmHpgcpWpBAA2J97CSQvyomCcdLXTr2dOUm/dfeVnlYEnonmMJtkzW4fWw/Wxh
8Z51Ak/1TEf3eGi2ud+wAUgmkdKlbiR2pu/mEZ3qGPugqe5ChoaI5LsCSSqdgf/5
W3qf2+OwGqnn+GFwFbXFhpb8cpg4ilKHSCUrYVAoTYNT43UObnYs5+hgM7RgKUpN
yZoLek+Ji9m0Ao5/KbQUQU+C9CKXngKsVq8LqiQwTzKckecNZHCNlKttm3c9n9bD
NPyaKB5RB3IITIdd9/Lq7C7/pc+5o/MU+rMqG3i3tg2c/I2CLoCWtw57e4d2uKei
pJyznkG/SgMlUI+f2ln+NvU9KbW7mIkp9RH2/TrHhRL+8jJM+BkuYdlCRM6uq9GE
plzfTv8OKWff1x1mp2oE5SPOJCN3Fp0PZCcrS+6q2opc6P/yJt1lyYx6Py+gYIRP
t2gDqusA3Y5hYEWcuHO2aMKvMtweu3i4QPOGLGvJsKu7yn2HacGHeaRnFBuxLpfE
AsxMJpNvg+tk9siB2y7TcDNtroNcGVL3YOyEeiE8a0CvRHhSwNPGFd0e2m9At5c6
aGd0GBY/FZwKaZbLAKGLXePqCFEYZ9GHzE3lSzaLPHMkwB4b6H/ETnlNC3VtUqiT
R5wDudV8ufQnLuDRFkNNuGJpHxk4C2zJZORNly66cEJjZF0qn4+q46ieZNHZBxgX
sPgNx5NoAHElk+k7o024ZYJWh/G5K2Q16r8C1kbcJHdKl7iG84oTLEaSdyExW1i2
uoublRrFxgOaIT2ndR7ZQE+c2kqaS6ELzbWGrUqHJoz2MEVCYUvf2PLJqZVdEVBs
PVqrtvvfVYxnVezMVY9tGa81h4Ujy2tykmTEXaLfwWeI7aDF43/RoZ1NG45Piido
QWUP4Z4t51vnjE0flbhF/b37iOsHsyTzt0wFOVFlbcBN7nk2aFhL11mrPKJaPPei
25N2CfOphNhF4txWRRTT1lA8UN40RhTYrYMAxLWaO/4KJFGxn3o8nsS9sJvAk15C
t3vm0rDoemePV8iadyGZLoe/MgemFfLIPBi/xQ0tKLk1jVO1GBUiLp4KAQQQTXIv
WLeWxupOQzIzQIG7Jg1eAKP5T7WI3DfhnR5HDPwjbn+gk5G2uAIfJ5v2YiCzqzQT
HGDXZqz6nLBtJU86X95WYYkXh4dDGm/lWbxlY4qxIQOUD5oHp7em3Z2PhXWZ9QG0
nBPnMQws7BwiVMZ4dXUSEcWRi/XnbYzigH1OHStL+9QWQ9JYlPznsqhNfhj3rODl
V/4+jxk3+b70rprMnxa1qtZ6c5fEDRMDEjQzVwW/5ZhtbUCcI70dCk7FozxgQ4dj
rdYll5jFBs234ebnuUhI7TVj5Hj+uq9I9BKGZqfPzV34tDj5FJtFdcyts60WSun1
JRujp0V1I0x9yW7E2AEPfLnmZoAP/oORpzV1Cz7sJvknlbc2PAFhqMy4mrbwyaBI
ImVQJ/wDtXZNBptlT3ZwYpEZiRPQOoDV+UoZs5nXOwrKz016HQn4SV74ECGSFdJv
pANAU/q2zt6TSB7d/jAU6pVKCh40ufb5lDTytxOmEvosaabgNiUDWEpjgJIQLQM2
Lf7QrKbKZhPK6zXA5PwQ3VoGEewFOSB9iGExmNiYq+WDrA0ksT17rmrqhbDNMIuL
jIE9JDo6Y4PtO6jOm50nmaf8ky/+hq6RbaJtH6vqbbj3TgBWrgVn9uG6gQLyIcf2
ki43Y72jkrFPkZpb//wYEfdKZnY5J5DjyyfrEA3nbJ4N081eevGcAWcLepwXI2ek
OcsUQeVWfguVJkWnGHrwWR+Av4Oja0d3Iu0C1Kfewyrn+xgWMJ/BfQecMyxm7AKo
S79OSCsfEaEmPkYGtaGb21JfNlYoAM0CR4lsge1lVk18atf+wcRbo4DZONuCON+D
ZHGwj685Z7dO2wXZZC22zcf1j68T8oUHoC8tfEazFYKlSYgEXlQX9TNQHu02a2Id
dMh/FUAXZu049BZEgX4qkWylON1llcnsY2+1dEtLrDjhGZgFOiJ4oaYCmK/uswKQ
U0rf1Wo962uCZve5gusLA2W1v/k+D0Hb4rEfNWB0QPEJ9SBSYGWpKlc5EWYuptsl
kBufdhZx7xFza6Il4UxRbWejTGPy6UjtPcMM7zxYUCZcAW+pFlygWDKUv5JFNFkm
7ZPyx9d5c9ESJPlXF8x6zXpERj7by8U9IeIZImaHZowfbfrZsHoLoFoIk8bwqCGv
ojCmPuxmYhr3k1n1yqldfnD59RtDc3qMjB4aSXBKd4jy0QNiIbN4Ili6toG8myxW
OA+zHhyhyfhEi/CrX3ZN+AqSI+D49DmERcwPgF9dCYIEGtrjDaBa38kCFbimD595
619x1lmNdghPJNsOqMPAF6aEnEReUDRWYdK6zHR/9IoSIYeXeyhhObg3CWVmMU27
jDHhST+u4RDWddatgSQOcZ/NYhX3/P0jZSsdbdzUVS2Dw+rw9VjuUl2w9mO3pUIO
0KjHu1g16bn2Qx93/VU8YGEe3scc3MBqzbOG3QHRoKt591gXwHpaSRsdOE7VhD+w
Nc82lYCHOIZPi0MArijzQqxNWiPZ9VdMkrcAWZykN5VDmSRmXVYyasRVG1Jc6VgV
bAPyQYCsuOZeXo5gW1bXokPIMB29c6oxBXEAWZXWfayZOre6jqto1ZOc9SY5RUyM
0nfIc2ip1pOHEiOcVsVhA4BJRocHDc0F8h3nP/nKo4pOkMwwAfdzaOcHFWA739hZ
eXcxx4U8prdB8/onAswcMwdATYoH8736f6KZQc/Ybpc+wk7wMJJJOMOBsm9Z7wnB
XbDyqjBjrUyu6lE8Q0CkU4ncwuwSXhNyovjV9C8t8tnCDnl59avDsTLV1pAtkNWC
WeklTq8wm+u4+GGkQ8gFcZ+0kPWiUyYscAqvq3mDMgpV9rhfwALevwichETH7CvX
OD4oMxlWefQWMGRkEosUSWTpuTEG/6nl++ZQ6vznD7YBSRAq931muyRPzV+qCh9O
4RhqADX81eZqhlU3UwKOlpyjV5yU/9wMDbpK3gg40XVbdZo8QLiEzHu/Y4ngemf1
JfSlClFIJfX9ZJdXiHaE2U5GwugXZqQTJ8cOhWBv4wsZ5iwoIorgJnJ/4ikmdSYn
tnf6R/cidPsBSZqh7CV9OgFI+5/L+VH+IxdOll84nOPAc/eFi4qgvAmnpm26HXZk
zmklYCbakAvFpGkyDAhhIkmkr2PQ+Bmi3jUbrHQxi2iN/IguMVZzxd+kouH2V0GR
QclAVEKKrMnelM/8GmFTMhfo+SLga9xC8cZXmctbZXc3+1irgXlfK0cdL8cWlxLV
IGtJeLehw9q2nVPRXLFhg0m15tXTtn3MG5jHs/B3D9cAjV91+atzglNy1ricQVR8
wvPByvYvOi1FiW5wXjLBbg2MQMfQOo/rY2oIsCF006H0iRFEvM3Kx6zgLRRmT2AW
61h6wVVm413Mtgeudwa26ujzwrAG8UyXJQK/8EIsf4L77nChP8Q8UEaRtcM8A3Ku
vD5E7xYOyEZcAbKITVIhEpdrvhmWO3hOYXPb1swStyVnYLIM/WJ02lLsd/Q58w2F
lnBxHuT7H/SE7zLKlt4WnLr+Anm0tWcTNxDPYY9GyWE4jOzTSkOLYbiOYilQFXF5
eULi1Di+TDS18JemUx2K8+QQQ9H7p2l8a4tKHfjbKo3Tk+T30PF+Kq90PUIywlmZ
vcqCZmQxtb52Ns2nnHNfaNhY+5qknZ5ZOjdjDXBmBOVwvo9PbteavBVFiaBZGgYv
x+8nk4F0k40GglXZwCRU7tVHjbOAMMXUVEBpat5/kKwKpUyF8Xo+il4X4YCuE8WO
p4VkfeidzSs09HwKFuDv3Ja5B5Jrhiq75tfzYbQoIdZmXw1Foin8wC9weUfp9FGm
fWEUB+uaaEWbXwOZ6MzRdVFmGfItcs540goo/0M21Osocl5XQCbZIghjQOqFUtez
I5iXoEIQUlnOJClzGWYlJXI89d2uqz8oHbZVZk8pJv8HnBw4EPXp7OK+Gt8izDB1
PLfAycSS6iwllkm+p4MnxJHmGWEzSneFp4yCjXrNQiYIdTxSOBgFrZa6RjQWZojC
Vwp/nC/nppeBcPWoU3pbX0ppxkpzDs6NLo3eOyck7WUzS+l8zLCNBiwi9kBQTeJv
gjHJxMu/t0YxbL36f5AzaEG9WRin3SmznUmB5Hyne7mkTLw/cLebjnH0QZ3N/qUm
4AmwDF3a4n9m4cMabhs7Nj77TIUxtuCNgYhf1V+BF0d2JIXSiE5bjgAgsJ7CfTpP
MaFiDwRCM4Suz+RGBTY9xAOjcwzPtkY2KIPiYMiPnlVy6j+8V1fEWdg1TLFifsfU
WQV73BWf8uZlkmXuC/LPRsQRwIc92J1asV7QNgFpGDt4zu83k/cjJ724dV3VM0kD
VeZNJKKOWG0hZVAFD0aKuMkUCQruASHHen4SX2Ue1ffvmG9hNfBmmDsMj1Kw9B8T
KrH01eG6H0FtUd4FZyTYnKCUabnfdIAs4LcXIm5ALlD319Kn4PcCnZVR6okzGUUW
4jhXEg3FJSvahoggikkfAVqBHqBqgo+gG43YT3MLZV8s+GFToKi1MBUFUkiKwanX
LkAC+ztOA/sg6OFPeyjFhJuYvUb5UPuuSgMcTkY5qc3+YXHXQ3USUd4TUZ80E/WS
/9RJIs++9XRCX2fAyULGSoJupKnREHzHvsoxgAak0OWUWI2KQmvdRt6nSyd91iDZ
wYqlCfP8nlLSyxaEZDuBvUGHVv/NCUNGcM2zcVQWKuF+xTnMGNG0DYs4JrhAmQZ4
hJZDtR3Z3Li0wCAOmvUBDYAYJlAMskhkHc6of7iinbc7MxDcXAftFB2AIiKkKNAF
97fPt+k/v8cnU3Wxaz/4w3mj/CCuEZin9EotsT1v+hZQu3Z/uG7N6g47mr0NfaZF
uEoktVJMZA1mQQ3u1ikiyFMbTCciZ1HCNbsA2a+awiusR/am4z0LOpn5+kj0otov
tkVQECpHtLgDCuUah0GP5J/vnxNyPy9ttmcmOpOPzowBRi2F/feHUzeq9CfR9G7i
Y1hndEXJrS3D5qyhzGoSdWE/YgWvdaBPygFwGBhv5usKYyteHWdlcFySnVFYprT/
AXnTO8Ge+/nVdcfNzgJh/q2sFQpS/6EBBk6ULq1hiVvVwSxm8TBKq6beHoNFIBxv
B2PSFl+uT/wEJZfq33X2oeUteDyJEVTfIO4vVwwtvpDFU/5E18eGVSuNv55+ZZGd
mHMmShktFo131WUBdrcIqjvYgjZwNEZ42neeyMrNFwPW07FWj8lvzT+9RoxpB2mx
LEcfgFLkEX28b0W2giXd/APp7GtBLFnWNhUFou19hfWDLdo04ICqFJMARpfe5tbu
zt0hUsuR9X+++GdjVBXqzqQDGEgLDTpakPUrtEYaLRxvqtj1VcUmIb1XSnkzjSEE
JjUyus5JPnUkMVENS6e19BMzOrxdKSteAFv0Fj094oPcJ5D58/IQEqXGqXJLU599
WJz4Z9NW1My39vU9PeKcNTWZWB+z4aVqSVpbkwIIohvxH9mf3jDAqJMD2YPTbxTg
UZWMjYUsB20G7ibnoOawKBPdkMb55+HhJl8qq1GSiXw553dN2eBknxLF/4BX+UOn
Xxi0bNYvOHPrBswXK/CVEoEv9qF67lFshjZhVyCoM9nPWgBjA3vrqk6U/nBFoZKs
KV4uPgbHVAncBjA4+IBLGPecPbDG658Jb4GXUkLJhSJu4scC31EnAjdxqptPrF6a
CDe1Gwla7G33zSimzcwe93v+g+lMxU5WerCoTBr2ZOsCpp6af0megM2grBnJ1JQ9
gfkxtp4gRxT7+zU62Z6D8IR/5HNMQo6/UURXKLNryU9T6zHdxhAdbL7cbZLTq5/q
4xeAcz1znZe5XCHVzDhiU6RCMc7kj1cQIBZvGYSMrdalSFswY5Um5eGqy9ShrPc0
5RUyAsoZeSb6gV2VztuBDyc6ciKlJ8ItXDMBlRvf+Zxrq+DpfUvb5xVxSokXBKlU
YO6+7xePLx541havepAMbEtN12RlIzRoL1ykwEuA1MllNsVLR/gsQcjzFQI1txDs
dvt5Nz4qZ41/fKpkxH/cH/UDhMgRFXZloCx0y0DJZCX+QVi87CcFmIuuDhcSMsAr
bd5ugmnsH7r9vsnomNxOpDaA9/UNsxJDJhCOjKmGWt0loe6kczEcWzd5IhdvR2j8
zblNpepkCqZ4GfLASpmTwoTwRG8GM0Fxus2+GGHbVKtiPGHSQUeuscYt+UN3wQpV
BTd5ti0+0rpXO2dtW6+Mpy1ft8ezNdW/ZtzxNwVtuE8406oide93uFUKUjM6W//m
hx4A0uypya69aHH807iK3zQVuTRUIC69D/jG+iLyMXelqvlRPAZuJC7st6bJfGb8
mJ+2W2MwwoixBPinc02vzdbCVFD2OdqRDWSNZ0MNvU3eSvmCgpRY9xODpLzKuyCI
Mp/VL+H9NUKC60Nzm16DM1FfnU41Lea62DbUosM9en2Cv6zmKIdL+vHylvP6PQzc
PZZBq1HyVfeDYrSLqFXUv1Xu453gvcC/dOuQ4WBCm/prRxSLVye4N286aAzEeOgJ
ACXaNBDW2FwlyjoYac0hFxOBUASg36omTFTxegppmfcTmqMHcNrskMEYsieQ0RUB
o0Qdsc8yiO0qRGFRBLyZBtMGe++gQitCCktBBqdr8gZQtC4jyA71aQNMaNRRB6B4
u8LOXpc77hUZ4SgkLAqZLRFIdID0bZimF/ll/4e6PowEKeeNJplzjGPwoTUHIliY
z5VKgYlZ+DnbFjBSmEzTaSU/kFxf+Wz+mjAM3vkZYWZXGUhyV4RRxMcO8PKCC9zD
+tv4pGv15R6hTHX4Ekj3KDARSZb7Pg5jJMVJP3HF2TFYAlS+Hbdf+JyA+mm3koX1
IWG49ngOU2FNMnNJ7qomJrixae6ehjM4Rwd8L4aLqZ5HvFoeU9fDKEBoqlrdfRGB
zPJMX4dsh/9BXccbWsCs1JXj5Asbj8P5pUWFG7dOrtH7dkbP6rbFwuF3eWPsS3xY
Y5rFta7qojnye0cZawjy6poJL+dtt8G4fkGuPrlrA3X8v61s0dkyxkptfKqVVQlM
Yf8yoRkK65CMM1+hgXW9BRJVS+OiGWtRVaWbGWXnOYqV2MignI6UHSzHDJktdEI9
ihQRrPIcj9Y38mXU2FBi/GVnKgdE/kTKisebX8quKGwSI/ZDZgml3tAeha4wOGj+
En165dAvHYwr/Nn2AnlFm5IznwsrnXjtXAHF4X++2CcXdYEjg/12fPovld3rw3I4
nLbCAKwK+k+/SKJC8oqVizSPR2asoR8uZnqps7l1jZfSpjFYFZl5vuRA3MExemb0
C10GLxf9xXJ6f9WvZvYbKcAkiAb+EIoVBpueozYZyu2LJBQX2qaclxiUZaHizEpe
HsYdWRhIM3djbmWwig/GXrODCm9WbMNaQ3+Fb20Qy+dxPHkh71AtHD4rhuLCD/AG
guoMwuGYnwiB3di2ma3EMFHash5sP2tzcA7T6Q9+hYLj3k00w0y/HLn9Oz+TUald
kFPjd2zinEFFvYhc10YmMwShzCmmddpLH+x9UGn8k76wlqqPvPdnrHXeIsuBCiDu
owzS9FANFRIuVnGmk+ozchuRhZzE1cDvwp2jAFXSQFqENPoSWv/RnkZSuSjIZA86
pYkBkvt6bhxJl/pQ72Umr5HUSY8rw/UD+cpA+h6cnI9EmW+l/Tsf0SibVwpzFAu7
k1TxrL9AVrixGy9BZ08OPMtyCtE2tkJO4rlBt2m4aV/skzoIu3SZ5j+9XNM6zbr0
K6lnfSQJMyHguMe8SYotQLrETB5NkC4vpg8YVnmrRpvM+llJwQfndtYXKaCTkICS
/d2j0EwUmYwpjMc5I7Co0bNNPZg5WBxAis5i242fcGqvW81QnkNmqnZlrw/dk4+A
1AFB0Z7YA01WDFJhVSjIap+aTKj/Xy+LusDPu1w7jn3zeGqWmorm3THlJeEj+1c3
rzkfthqaE6uJsKCHjK9hWNh5s/bbW0WDRANs0iMSUN7jnxlZOxquB07z9appcYo/
yLc+oD19ulbTgQE3KBIiY0hTHATkii9LC6qPqVWrTtYu0xpyz55d31Ekrh9My6Ph
SF7lzyEfWTg8t/aTqn0Ed+GZin2jebUYvf5crokLW1WyH5QgN7eWVhr/QetqneDf
GTXXD5qjTx/yOW17RsVyifxLbB+dsDONCePLfcAOh6mvGjREtlQq21saoTeF+iWS
VpMkC6WnpWR0Rj6BwAxJi+Uia48Iobsh9/ETyffwfVFlrQJ6HuCQeprKee+OCcDc
wNujdzbNkYGN4ias8hnIEN2dTdasxOkLSwZuW5WGbSWYkOxHfGi627HppoYcxZMU
bM7Hwoqu379xvo0uGK6Fvlk5GteWgxwh+nTo/sWJYboKXVY6IdJMjvt1OEN7tiUa
xLbO1kTdTVkEIXxMQ2f4Cgatq0Aw+lCRciP5n5T3n5vFcPChb4g/capnMx425wCi
Qaf9kTt5DSfGfol3Q+m5HBWnXfMAxPJS79wv8Ggt6jAjgdXnWzmAskI92whgUneU
9D7W54s6fyRz/XTgy4RayezxhGySqMUPkEv8QxcVWW9nvczAKFPatRJZf9J50huD
h+Ov31auPXQ0go7r0lCXvzJpQgRtabn/G8+t4j41fwvFAkeJmNiYaUTRAEOEb7Xb
LXZjT3Z10ksS86SaWUEDze/1wOGf5WmlaYWh1qJ2aATHmlqj5+Vv9N7corHB4LDe
/iVbWtnwRUvzFKL9I3W89uK4XrJhwnOGXfzJUgYHvkR3Df1SzrEDWmjSJ5+oeLSD
XPjl1+3Ifk5FDhYH+ZiXDTTHfTGD5pzfLgxGalOaSrG22XIFWstolykX+KEQbkhS
xEDxb7jC5PamV3TEnGwLifMQFMRqWAu+MKWMGchebVmajTCDM7TVC/NYmxB/Z85q
RAN/tyNv771CFJfiF9OPQUxeAM9WcPKfHsqpbKHUaciq2sGaZlMfqIv+rSHGNpYh
aA5TvLtpfPTe1pA5kWGmx949+oepZl1zdYz9nWrh7+CHmOrJluC7y7E/2s2xYlcq
034X6gr6KLhW36Il4LC2ooVD7731PN0lUqL2IpW4LqK5fJ7yu4anR1N9lE69EEPs
6Nr4Abm81zyS7RJF5KaCSIT9BahVV8Zz+QDJ2KgpdYjmUu3Rq1TKNI52TiOXSqIw
ACMEj6xGp2Dq4M/vF9+EMzktc/gtpvY3mZu0PYvhYVO2/dhJHR7/HriscYaAqwq8
Ky+auMFcKFET9T55flaWfIbIfD1GbXSVaSQlG9F0cZ4OqXoa35Elxb15BTiOGwzL
LP+m5mkucL6McHrgRGqBhQ2BwoBPhW2w7AX2vW6svCRbdMHdsjUfSQTSmUQeE0Zp
+o6kWhYrC43ryMXHSKGVrHsJaD8SQ/0GGPp8XYn1D9bt80KrTiiT3A/tn20Hy0SX
3K50TIVm6jWuvxUurD1SQXI8jtQ3d4TOq5bIWwToA/+sXljO2yt+LC7q3vbpDpwi
nwbVERUsUSzDBtHkkYXaQ00wRfnBqHvaPsPxfyp9avL7U3QGsnKujJThoBeeeHyY
R0bMc3KsKbwSQyZalI74RexVsMvGyoF92dYGY53ATpR6aFRAyGlZY4+DMpD8KEv2
cGeu3BSL/W7/D+1SuYZGGy3KzF2dWqVs8cz4CoLAIXqCD6KHBxsUM5J4k67IW7fc
ES+g16V3rAEF/gdduehh8ZJTQRGysy603UCGxn1bSi3cEaajYNsUO5LO0q4PNYub
Cq8K5LAwAxJjrnA/kSlmGynBnUaYf7EBJTD3tX5Mtl04XEaduez9KWYwa6dnzDyO
nGmvFCLR69cV9SIm7UtpYSTlinqhB/4oOSAPszsp0tfJY16fKEqm2m+2xpW+EwKK
TaFaPMyRM6UT6xaPznLfnQjCBBGBdBaBJuXqQC7EoUuSeNI7CQZTED+QeXQdj+ad
Mn4pKYFsuTrAqNO/3OmDt01AgbytcwdY+ahuBeJVB+V/gsAD26KlBgzp3ElP7mn4
8CHEBUglUbm+kDzO3q+vOI02B4BZvEpPR8NU/3NG/oPzwc8Dryu3+gtvFLG10yzK
L2mLepksaA8ImmdaCHHlIozpAx5IrP9irobGiZDQeYR8eg/hdF04xdC68Q5dW0Ol
7XYIO1mzw5L1n9TN13sd+jWhVV/hvDLYAb0KZuKvEQ7bQkzvUtaHHY1NZfk1g+F4
UnVR7HN8/99RxGWmQyd3rP1CgGC1kbso54vCVkYjwbGbDD47vG7wm6dzW6yRxLG2
KlrQsUwGPYlMkJYbFYJ5whacQwlRFHQzkvRGZ1xnenQxZn3WHAI0BpV3DfIAh2mb
t5v+VIM4PcHTbBgKog7Pf3SZFMfIF4qiSRKPwfCs/frfWv9L3QSUtaorxUPKmkgH
ZskRCaE+XExb3hLnhaouXOFy95/NJ79Cw34tyuLlUj+b6skJGN+JvTrLbwDUjry2
1dG0GmMG/ucQJuhtm2N5r204tga1s+2Sbwo8zlByrEGmNhAZt/Q9/S3+btKVsK+I
drJl/IbG7+4KOoYSIPNu1U+PWBeesO98WnyGSSVYWE1cvLjSWt7nelXwiqJXL1fN
eEJrhEvivGO4Kgfe8iFTmu8cCgYQPJ0IRy/N0U0uHv1c6gCQFkQQoSG6wH1lfXTD
GKiBIMLVL7Eh2IZIK7QLLcHhqDoyLLaQMydvfG8oJNCxZkLS+/Cb57kQgBBk/Aap
Gvu0qh/6wPZ5mz7IoyZiZZDvfEF2jb88R4s9nK96uSld3FsX6WadDtSxn4n1U7l1
IMlqCkBO9E/ns8tc1fHXKEZPw9zA12VZ1Jsdbu3dyXgQpWb+vSeT6bjr70layA+8
wYIGenkLzJUIVi4B1WuLHOTH7kZfJtBASa2bT2GW6tVjl1zZ5qn8OB0EWYRVw1XL
SRHZIAQ/gSbpOQcHX1ukIXjbFwfFQHtMPjnSTk7G3TVJkwh57fW2dq+cNmo4Bjk6
F1sRb4n2v0DBUDvrqOLV3Q2UqFnDewwbDVi2qbDT+FkZg069E0hWVw8ENwhtCaUt
CGDrKomxlgA6VlnU/vBdi9lmTf6seJkVxl/eqTBZXmeDky0klBz9VYdSijbfkkGq
tXQlHE7eno0B2aCC8ZV+TSyVXtertf5ajlTGrQBiBfE2T5O/aCf7ybSKxR3njO08
9a+RRU6KYTW18S89HsFMVrNJDgYaPlYGr+UHTrxgEWfbdtcGpWod213oQbiVZL7M
pcEbntB9lB2T5zLxzsDviRgVTC53hMylZxRqyuyexvGpDmR0woV1+BQq8zLz4+i0
6J9KHxOEByQ0aCreSqB+IKKvaIGEw5eggk8ipdNxnoPA5Ob3rME46wxHfT/O+Pky
rDutuwAzTu4uK5lliigMppSSYsANS/JzpY9uPui4ajmGoM5ZpOivMr5wQu1nzUsO
x1qa6okvBYKHGeNhFqAerRq5P7h+/jyWIjwSIBo9Yu/OcVpeA/NlXKC5JFpzAVAr
yq3WJ/pIaNwL1waytcqEdz/97S/UKxxXKspf8rKa6em4RVcZzDqTSRL8O55nyMIr
lesel7vKZ75G5kcj9eB+ttNf0sxaXPdCM21Hc89gKQSxz+X84idJFKDpVN1cpbIJ
HqztHsGUJKT77WCk8N11TL6MJcpyRY178DzUejgJENx1hKcyT83tawsai6FTP6eK
BAx6lm2Wpv3+A1g1KoundOIAtGvl4mXT5pLtQq4//y8Y5G1g4VPxyhRb6zxCXF8K
HmWuMSWe6lms0kU7wDP4moB9Sm5wMBr33DEeoCHHWc1xmNX7N/fPQTX12kM6fovu
iz4KwyUxC7RARBwYhZINqqFIfjQ0vmYyYrjTan/CnxUHoT4lL/IAKyG9Uk0Rtkqn
sg2A3amHoZRkr+7v5kwm2z38VdZVqtXHyFY7R5hl7iTMj6ivjDW8xaL24Uxj+RJG
u6jpKCBQ9UCIftOvvfNktIoHj8Gye/skC6RU3La+p9Gvz8dHAlkjaFF6py9YyGsL
2EtjBJpH3mjGBnCWDTQGtWN2EtPQyXnTnfynaZn9yZ9pmMdAVOdYw7b08eN1B67M
IAyOub3g6B81GZzx+pbsJUFhaKvcKGZskZvfB+H60YQxfBQBADX6ZYkBhzlav8si
ao3LOUuf04Li6uaxVsg9Lr+HQ8nmLHXB0dW6OcKxxiq4nxMCuoHiiclJHgxXg5q6
VQaueJDRHAJLxxkTsV9twEiqaPZ2siCnWlQP+7mT5upy3PYvt+6ORO3ttOX83mDS
erAdyB5lPyIgfD50X2QaW6Ffl5MPbTMPD9Tkx0mmRdLihL38IjRxw43DzAk0xPR3
RXGy+rFbCKHQ2NEZ0kUueO//g0qaR9sXXcttFxaAFBa6AfOkVuJL4nSlwJdh7vra
DPb6+9AdHCbueiBEa/Jxhibq8RUkjV8FtkIqs0IUVwiqS0E/X4yUIyDWmUUFv3Fv
8mZ6PlSJX0BcoZbLcvNXv2pR4aAqOdKujnYqWh3QF2T+anfbpmr5gNOhPc+n2rl/
6B+Sz5VuLZ3AylseEVaIgXB+FICl4J66QPF7+2FGVdYtESd2q0A+dAPvDCowcw04
L6C2rlz3q0oax2aUKmCu3nkmDJonKL/aCnaleS4bQ81Aeuip+dsfoLysaRSBOWNA
sLHOUX0qOV9zqE3W4hsCwDdAi5UeMpfC9PCMTSnctcDnuy41oXD98zF6w2yf0g0C
kJaC2XExhYb5hgt/PVklgPR9jvXG6qR8U82vAaWb0t7KtQwU0yf/+ZXaAIakpCOM
/BE8ay8lnF9HA+p+8WjuBJu18XKi9PW8lBEHMVr1arI/Bz6BXzdceG/bRweRlOCV
PdyhWznGHIGFMVJdm7O07Y9iOweBv4RCSuu1sadz9Nhze41Sld7NQJUFoNyX3CbT
PhV8zAkANadPNrvFk7Y+lTEuVasCtTfDipNTpvfUOS/mZFEy6JyCvJiRUQCSfSVz
uJKpEwavbrjIyxUgXCE6WsTuK4h0h2+xWIv+Z24MUxu61EzAJGfK123A+HoY/aoD
V773aRoNppVkH8pRI335GxgOUmnt+Ruly0E2T1HZFAzdek4AKXSIPsQryejs/wuM
eQ84iE0dg+M9bz/Dkdeiegf3WVLTRaqdUNwaJxwkJ5vAqhc+SfhTUjsrleHNhch8
CuiP2rRKAJlLDYPD4zsjCVfdE19jomJq/BM46wTbJFQPSaRtNLrhae1Rqjr0Dn0b
svhJeSGTsRqBbcSdrAIENoLayUT/RnUYN1sMpkfCoc9J3FFvByRsbPz1kDr8cA6r
C3fLVAFx1IsaIRAjtyLWF3eIASnFq0vsSOWyTli2oUIL63aHDh9DsptlJwlEx4/9
ivIsXSiHGrXJm9X/M7gGr1Yr/GGfHkt8lXHkLwpFMuwKuRTy31Mor321fHbJezOt
BfkSCwCRO/I9EskdTDdiibcE3njeRGyxvjCv/YCKYXEbPCzKk/v8K5m6fDbhsAl0
9WyKjWq29OeTRHoIdZ7Lmwoi15eMeU11SoKjRGrwXLn9Unj/whSxXC3DshRa7XVQ
RCOxSJE4F9BtFn4NctFrtHkbSePivGWkpWuL5EHjLqKj/HfDRgnYlVVDxJVdi7Qk
KZu/ek2zFz2na+2e03lWr8HV0MJtWfDbPRLkdtQ0b32tsUOi4876f8qH8HFYPlsW
dYeOkU8Xc53qDjdpoXBBj98FIlWk8rlV16OP4p7lMaAFCyldUKFuP1OeEytbIErA
wHRKaH/ESu91QS4lxjy5X03APY+9J4YqYLlm/WTL33TYhmQIeqSBgPIaTxn2iKfh
gJzMw9f4F0laWr/mth1wwiIy3brF/PIjs3vBWQR90UvU7D7ITwVB8+0aFvjuhkyq
XdiF5BeLctIdp/FAvdlKYf/lrGglpgUYzdFujOQzCqBXrNW+l5wo3cGiSNfTd31K
k8qge7rfJZ2d0rd8rfkHa+hBzBNvt1T4D32Gw0xTmn1IvHvIxCvvowQcGj636NPB
CVAcPxOBout1Gq3QtURfslSXe3LUrvnwa3Y6gTMwVB2MgwJscizUJVcA0PJuzxKc
7ls4aT/hqgS/odtrqmFUmKV+on/OD2aoSuey/daurWmuIRIh611Uw5z+Npa8tb5E
/WrKdC1K+bipdTZ8L1vpug63m3WgMax9c6O2wVvJCtjjW5FYTlqhL84ipnBQr/5I
iPEa+vlo79sQ6CFR0B+Rn9iGGOPdGS9OaARhVeAnTEwOxy6fVLBpksP//PAXTa//
nfbSW70CKyuoON4553BCQLkqnPVDaFSRbfMnPcBnTv6OLQ1s+1/GyJy1xXZgExdi
mTXaDb5zl22cUDcdrk3KBXQZJAUxsHTtk+rbO3tm/Gv31D1eioDgVIwdGqrhg+NJ
VoaKp5LzBNUS5LUkjO9VGhiEPdXubcTLCLVPe9OGMPvLsDJds+GLO9ZWz4b+WiVH
XN1/Vyt8/o6ltxdJSPRkNRRZk+oLUFfQkOgAc1EpgieFYfd1yTMa1kznPZzoNUmy
+zC1XBYYI58NUhLcGqbcPfPbS9wkxsgIfvnwfHcWWAAho/fqJChdmiXZ59vvyB9/
2logjyPMSYAPdcLWCGy0QaUAP5LwqXvIoV2kOiJfVjlhbROG/EdWKalkWN/62eBd
LJExH3KkdgIIc0ASbqCNPs0FNuvlCJXmH7b7K/NA7jiTC/VOXxM6woxuDQQxy66l
AYkgq+Cb2z42xkuniWPaxTpRcnyzjc8pGw9Wfau/W0ff4ctlBBzd4/9HK3CfT45g
L8LKOQx81F9lbvISDJsk5dlafgAsvujFE/kZxOQmocp+hKj3+bI1s7Tgf3wz/dMY
XwIsoby/abPJbdL51wIJGFOu2aJMgJGSSdd+uIU/bahB4vnt4H4Y+e7xCiFPT5AL
MA1/ntDnJ1f76Rvp+ZMgGey9QbGbluQ+/yiLkzeeDRyN7emUV6zQVfoPlmlfQWI1
Rn1kqDNjVVHB/Okjpf/QXGRb9dRE44vMoBZ41IsliyNVa8CFzMmqPeWUkumzt+E+
AK4PaPXfItS3mqKlUGsSZ1hpNuuV6f0+vKMT/hyNUGerB+Ogc755U7VDs4KT4ax2
9D/cmZzph5G76RkJPwOW3VM7InlAHTKIfbnaGLi3E96DH9aoVyF9hTsbPL5lKL5q
xncz8Jcv9GS8afR39RKObmwG4aHt97klfkOn9//oAGlW7KocAlbeEE/g1HlSl0tH
8SgD9HLjb0f7kZ3Cz17qGcV1nPAFF+xOUQVdhF4njETzntPQRJOxVKjuob6MJp5H
sx7vQ2RQ5t5RuAaw6bA4kKYvaTD2K63Y58LLvLztWB3xIBVyshsgBnKNj7/2kJtk
FvAD0k1X77ZTb9FtNEJ/InHGlw6dRA4PzC3uA5bTlhj1jC0o5bqzbwLOqljMutVO
DyCBg+bvNohuX0joFSLrAzd3MhI3r9/yViXDTJ4akyDpYanAvNRLMOJ07/0puyxC
z8ey5QIap81fCR+KI20q2I8tppLuRzL8OxwvHBMMS8FKLSzyeVyCLBMIPpiYD6zT
bEQ5kAuFhTuXaOpnvIg/j98k4ukDXJv1+IkG5x7XgCl6fFlbj9HWPXU+h5tG9Lqj
xopYn016oJXM+0/ASD7waGRIzGr3w78/KdzKGWJZ8hZgugpImz/4ILCYFB/of7mY
yt5orykoLJCBqajS9hmZCX4H75fQHS1pUBalYq9SCJELqxz7Gm2vHrJ2++SvsG6c
4BXurxnB9gsITKmTnqpqhhORwDYYA08MeUTp5CGh+V4SMLD5UaDtOBoxeSRQIKIV
zqMHfgYG947cSffCjKW29LIyyxW2FiZMrMX5JKaKVxl9vYo5C3T2T/Cwkl4Oan1O
m6ag4OuaTIakEAVtLdiCLG42JQ5vBqqJAVGNcG/dlACTXW7zybiKunanoI7B0z4d
IkfJ2oCChbykWXqPcWD+60MXEeu1fhmTlpM3r6cMWsh8xlNHRj+5zUXd5UMZSH3i
yD37LMnq+t1dUEtdBG8rkKiJz2+7tjbEsjD2J3I0hgqZ1gR7uw6x429nmDCLY11T
B/Od1yV9cOGK02mFHo3t9lbQ5outw/sATnA29LgC4GPQZkdgc6vKBdSPOB7FPS3g
6OZ1R5ksnWl1WW55vmx/wJpGnrvCPZ0TpSI2kINSXt9jmqPPTSgeKD+VVR7fJ3vk
unLO6l/om7rBioYvUt96U82Aa8dEndF0gZpEejy5wRDjJFTzVDQyypkSdwI7Gz5K
KHEDbthZrZjnPAj7m5qcgc0CAnJLQi4Qpv323SRvRmoTzQDdklYyOrGM2QS6G8zb
VpzI+bUVoLuf0CqjVnGHLSOmfLPicFZHVbLw92bviRaGn/gWE+OW4/26gho0+43p
aZQ5tDWVCv1fLVVD+hT1QPvLoxyaGeqkV5hvX5lORVbr8exL8SLejvTFmrgHuhH/
z7Lv63raBDNfLev/JjJFFzliOcgcZVVx7RvXdOR8RsXOiWWRtoYuOMrThhyc425m
uMu6fpjmJi7E+P0Ah+ENK9weLaF0767y22UFMImhUnZZ7b7FUGlNSIVJ88EEeUT8
CbERZLbXVBXkXTjrTke55gdiMB0a92gP4Tn5PWizJc1vqwoRwfSvORAt6LvhJF8r
vgXK9SZZcdjGvy3Wb1LMzVRY3nb6yJr6Kc+2hLOkOnNa1KLXCkNFbIZC8ctEyruU
0/x/dJqWMctB+gk7B2y17xDQXG+QaeHSTNxl2Ox7G4Ksu5iZdEPnBKmamPIf4IT6
baf23ZGQfPFN0MpWSI4J+1kdcT1eKwSKnnPq7rzHJ/U66OjEl4lYHDrRx6T2wAzH
luFMRKuTRxa/fs2ziAp+JXaB93fYDMn6TbRfN9ziSlSx0VkfXXko3cGY51M97E3Q
pYVrDrHer8rZfBYGV16ohPONab7vGq6ivSIQcGc2m8DZ8EAyUZAK7WCe4a9vzF5U
AJO01BHDAXLwqNTVIxjhlWPOEqZNFLne3xWU1uoR7sSclCP2/ajFyocK67Y0IKKC
MTPTgYctRUf5Sq26E0q+KPJfz0+OacsfZD7PPTEWbYuiNE03jbuxd1MBIVhAB/+0
sXdq+Ehz4JAguvBvCUluUbciWexNaqiU/UoIXp0ruN2QruzT0t6o8fMU3/ca10P2
r0E0lpA7e2eVhRAJT8dLCAkUDGSithX7ULB40IRTsS8oHKcl2RWcbe1KVLRelKT1
f3SxkZd/cvfwqlMb2r/oArgNOCuBhw/4OONXuiLkq+rvkp0e/ZDhJcZYzHUROxxP
EmrSbRhQpTZootPuVfSjbAg3WO+CpWdfn4EICihheZJWQ+icZiLFoLsI5S3i5uci
YsxBi4MI24oQklyP39MxgcgbnLTOD2UaZUbR3PEgmJFnIZ+PHFg3EKXLhjCvOMNj
vvLW0QCnEFJ0d/rRb6iUZmkx63sS1A5ylg5CUsRfHCqf5nMcNnMQm32SuKy03yLu
fwU9rgy5C5ZnehLjw/Mzi0shWD66OEr9JPMbm1FWm2AOw/H++2nOO8aCb/L532F7
0qKPdgaJgrAeKEJh0HAm3R7lp9uWRpb6n7IcEF2d6M0Btc62cV+R54C5VWg/fu23
uGNe7Cnq209CuNMiE3KSdiUAXMEYjuUSbtwAh11451hBMr12hvnZupm/1oXj4ztn
K8/WqIdl+8FCyCnIfEswNFMed12vmZemZ97d6PU5QB5FOlsyXxBgYf8XERY8IMO+
9LpsHEYPGpMJcwaMXWuDW4B6EcVZ4tTtKdEc7J997Mh/PFE+0DcVxZQiE0ZJoXw3
Kn2qfjX4QYL2SCy8AxRqt2720upoRh9Sw/3iJEgGOzyJlM9ajFgtHBKIg7p+SzmH
RJ2Awof2SV1vBNfoK5B0LaISZOqJpwdI6UdfjbWBb7J65LXWnNXTicrT+jS75OCT
Zb98XnHaokTpw0qdaCZ97rZvSfTJEssbSE9ziM++kzrkCVtboW9JTPc8G2jKLe88
RPtO+ELBc69f8yrnvW/83a+As2hCaSjSfjLmLlogtXfDKbaB/hZA1pxBmgT/RF6O
LAxK0EbnjXjqRCC1aEj77YuPoRf7IyrPmS9YX/95JuZJkPJWokarKrQtwltTyqzo
X6Vz4F/F/cci8u5vGGa4+O7zoLg/9A6vpiY30KHvcKm2plJRy2biaHe+yjl489Qk
2oC+78nAWruPeppUodU5GtW6WQ8IDTHMyvK41GxuQ0zkIsXmJ4fo6HSCfL4oUTp9
eBJEpUWkDhs32hwaWK7SVnC3Ux9/vsDZPX1qF2qFNKiq+8lOVKO8UMJojbAp//4S
4mMWcydvhAdAFUbCqiBXk8y3Cu3OVbdekAVdy7W4/uMhYSPED70F1aBpzeVaVOtt
Yr8IUIkjFLmKhEIN/axTrsXpe6ABjmxPOvyzBf74pu9fANIewk/n14pxLkP3MF4G
ywGey5m7oA5r/ypUBbkil5PXWnGyhxcKfinA4DpTpI36a0njhLSTuU7D12ka/yHP
J6FhuZ9OnUkxTghLEKe3dCvo+OwBghza1f8pen1baXGk7LIhi/eV2QuDEmFq+FaX
L5oKJripKPJdkntdA/BRPb7W2COI3U1h3tVtGortDkMCoqJdoNo/E2h9ea1PoYtF
TvWaUbJuMNQxu+Nk9t/BZe2ETw/hqPCiiiv/3WBtDQOKTP3sk6Uqx5PNf1wM6pSZ
fprFxNGI0Uv62Ntb6Z5l6kmrMIZCGtMe4DJPj5MKBJ3279S23jaMKgn1iZEu99SD
RvDLj30yr3NR2LHQnQDs0YT/lswpWW8bNSr/+woKpXyeyaZv7adLp6CIsyUBWvpa
0kxY9mF5Jxm4770ea7AflDbPAlwCia1f1Ds/XuEc2QBh1fszTZmpZlZq4xKWHoH4
mtQR9nbZCMDWee+n5FjADyrztOzJUXNnrfEAKqV/l2cUHBSFpMk9BeAqSe/32lGz
hnwHP9NjvQM41XihXWOM3Edg0dXF55f7OjSorVx3SbUm1xSblDKIvEV9N2YcyrOA
bdJiuWy9/5gYJ/TQfOQPM/2Xe/yKA3QBRYn97zXITJ22wrLgVro/HDumzKzYrqMv
/+GLzhOM4uUOtejb0hAdbdaAkPA3OTTnkEaoq7CYLJxKV0an5YtQrqhk4rSz58kn
QPYgRvO4dR4SLJcKxfOYAaDGsWLWkKQa6LunTOqnbIOw6yVvUNs41m20IbaesFCL
fBDPtv5gF4wtpwUtxTUun9q2Y4jnDQpVGoOHxvJsjYhO5swqFU/nnKo8cB0tCbhL
faMDB7+WjE9no8Cw2Si/I8W6wOIZvECF8mVZMr/hexd1LxfedS9X6SJj63AkDt1C
D3MCbHLbvwAL2b4/ebzhxmr5KXG4OLGwgDr+ryLIZ/FeOSxXdkzBMejzAyqmhXFC
Nci5tpwbI5NfTAEMQPCnLf7Shu/i61c19bd9YlI0HfLJpSLkhwIqDopfYcrHUebU
sRC0S3ibAMcfd330/CusVib4FtrvhbCsUR52p2f7gUuJFxy+5y6IxgQtMJjIeDj4
PoX4YGMqQM8jGfltSG/Blg0jybsfG/WDCOFuy9kokqV6irPOIu+rdaOxADKdBHCj
gv7Qs1ENdexCAvnM4oGwJEWkeSfV1XRlMP828bXt3bLqugserXbHKjH4RjbZv7QG
qq9DQI/cQMnI00sRiLjIIV1Ajtv0ijROe49iEcOz6eZoiMBlDgIYaKMl62jwgVU3
sqi/gPICM6EUQZeYqUM6+q00fj/nM+FKaUzLMY0bL2edNzoydpYi/FYVHisDfQh7
EWqjSnkCvogJXZcCPfxvEc9ZVBUm2FndqV7gTNXVDXENzmoSB3VzowmPZqbPwNns
gzYT8Girt6FOptYigektsIkDaq5cpGO5h7IsUeMd8zq0DfqQ1UB4ayl1ZYBu5JUT
giK6Wc6gegBp+sUj8IaSQhxpIdert95nwbDXuTztUS6DbqO6vEHvE3/Bobn8dPH7
qBK8Dj4VaCLwcyLvJgLtJudxmBbgxNffwIGVMqzZWj/88jrkgT5g+AtNV6aKg0ez
//GwYZJQOIAZrDiGxcwuudoV6HdKtdUpGGuvhtBdVapMvpjs6z/p4i+tJhyhlVJ3
Ta8Wsu+84Su9rTyog77SyHNhcZGYChrxpJr0MB3LwSIfr5mopBMrMV7GKX8MVK8K
xWasmNaYp8SygMcgT5BiXI2DmymG7An22EhtLV62GZtKR46F3nJcPYbjsoV0fVhq
Yyui0bP8mfXFlye3Qt1eMzjky4ZqliOsf5ravYsRQjreqxB2BqyC0iaK1jaG87FC
UKjNvoiPm9uAvk9yVxNA3gVYyKZjxqE7YUBLh/a5a2CFufeQNL1sLRG3kbyFEnGb
RkYlmIc+7vVUNrsKHZiEoU/fn4wlSO7jVtv2nGYU4bQzgKIl8seSoZ0oIPrmh5E1
jXWwbxmK13vnHJhdmG16fyYAC4u6xtS+p+FyuMS/25wHvgw9vNTkwsfP0ioHI8B9
xyEh39ATThJmvJrFhEuCFuwY0ayQPGPfasqIPrGa3aHqLJqAe1sEfp8bUe/bfvbS
TNPuUYmDcqfKKVzKiaV99tBNFgy0dkKAeQD7NQjQMu5gqWzizzsUikmAXRtbeAnd
yZmmfeNcQ7YFHv55l210NXxxYET6//kgbVM9BWQT0tK/h9BRSuNbU1yE9Xe9uUM4
P0C/X9fozrsUNc3pgVsxCX9BF9u0O7n3OsZhmDECTQ9uN62xgug53l6PCnTiPqY/
ywwfJXn+dG5jHya5KIscwfj4xSC1MreFffrfCfz553FniQtkL3kzycR1E6eAt7h8
vAlAvN9i306ehQRmIvViJnRcHFvNUcMWXmOiKGnCpkphM/BmZIlj7GfNrIQvKTy/
wiz9s/ZZJVcF/qWt/cEMI7fFNjNMlKlB3P994pMOJQDpCdgjuiq31S49yoZYWCsV
e1Pk06sdSo0N88jYuKNJP8LN75YEcKPwOeUSuJiklStepYqXkJRPsg/l9z0VnPx+
WZK4bOMFB4iCIVOsWG2eSIIg0sEbFiAclDwJ5bZu/dlLI3zepy4M96/2xXNKNIl9
nQOjLD7qLdzei0en7EfpmPw97OmNxo3fZMD5TELGnZ5FZr/QZv2BYCeXzmDqhy47
f7oIrNCuuw+TwNP36+7w+Hw7uEVRZ2AuQ+egc7CKcxuah70jtRFOzwNUIF1Zgvoq
8DYtRtmAqdgZ040hr5YrH9RqnG0Ro+rQW2jLNNVg1crsGSh6bIM6py6VnuwZsHyu
l9mt43yqPIrJh8hMR3E7Z06cf5AoDJy4gSg/yctC+znHBq6HmME8hBahzIdD/Qc/
2lNKZ5Uj0ZRxpmanga9KpNwtIvu+PVCOK24sqFlQdpg7aEbVzzwLX9B56tzLqFQH
tN6PTu21GqRA1vU+zxWt84l62o3c1cTP12v/zFRtT33C9wRCtK+6FJ8zp0gXUpy6
w9FgifFw5pI8giplb/LpDJFO0DzZgI3Dc/rbrPBXpbcwqwwx7Srg94wGpr1nZGF8
1rWuR2B2kQjB1JP8T2Q5Sbh3kdTg6DDZZoJbplZpODvTh3WTse/V6iM9Utl2Ko70
4sJKM4sdD5e8PIXz8fT/RM2NjIAn4Je54dJ9QP8lySfyzs0jED8y7YwUU5LovdTJ
mzk9v+dH75phFLRnULrfXrJerE+1C1cKen60DIWkkVwguEQvaN8KcYIwddzBF9Bv
WrYglNT1CssRFzHZANrXpBgnLOMV0M6OUymEY4eQS9zgmanSkeuyiSSYogdyaDUs
9caXDa9BVNo+E+6vunnzjWZYnpS9EuMyk2sjTvTssx6/Y8K2yy1pn1nlHPhIQAl+
nNKNucXUo1UfRYRmR7pwN8kI6nSgRBXz/WKpkrM+h0Ext8FBNEWXRYahhWj9HKZO
pbt6BlkhK2lBcrn6Is2xMyxPCb13dEwZNjlnX9MBNF7pYys9jOOQx+/BFaI6EKMy
JEByAld+rUPH4GyqAFog2W1yazdqy5iTa3Ydj64NF8wG+qJOdMQNF3WA/+psw8IR
+D9W2pP0LM4fc7xxl2z4T+nDzyFVdxP0bgfdQFqsvwZHcVXJjVqWhR6ch5+Qup4V
f+LhacOPVEVqWFWPIv4yPeFW/W+20n/CFrxWiekmMpQqsBPH42FItNR/vognX+e4
7i62KydYTFY3nra8mhJYAKvCTBGWh/SGQAXX2AIOvJQVrUdRiiKQS0ZOQ5GPvQLk
AiueY01mgEgLWKI2fQ/aqF7q6fBQW3Qr9rYabVP/2rW7OcEKHAK64elLF2rzhKIz
X4jDpXnBq3hbdv3UfmWYRVX/l09K7e6Rt0yxBDJ7EbwYldvHlZgAaPKG7KfYtU38
L9xWT7t/2k9qJYSDmqhc2sgcy61uR3g7qpaqTCF2GMjR5jTtTElgKBGSOEnMPSXL
p5Mu3ToStfvsQSAIaslRgdOtxlLbopg2+ur1fIat9flRZLQTz8I7nHtiZwIxA+yD
sUTZgxJ1ZRxekNV/cYoqyfOEM2vH5NfEQiJKnjLUkalqasIKuP9GO2IfsEdly2ds
WQX0dpFxG61ZzR0Ec8bbGaUVNkpbGSXZwskV70HX2O85IQLxPSQUks8lSFYumZGF
OEtGAluwWSwLHFYWCATRMQB+LrXmczFSKm3boWjZLlfQktpAATWlhitQZRmwgoEZ
FCHdB9KocNWMo2uKZNRkEEwa+HkBl+Moy7SfMq62Y2miXcjUVW238Wf4+LpqiBFM
6ZBrnH2K/fwhuA2uvxyMuxolA+Rvr1Lv3WIeY9yRgOyxKNukM6qJt29x133u+WVL
ssK0Lh15GuJmH4S552mHUYH03JcCdcT/xIJoEdO0V9j3a5avPC0L4bpcewtBV1y8
h0nmGZhi5CLz5TxfxaoPU75RcskBe7myBnLElooruX1DjzDSyQwWw5CQfOnM4TMv
yIIV5VDPTB3TVobSsQUojCtqje+qSdBHI3YIjKktpgDBSWg5rs1n/w3H8daKKPV7
WGJu3MnTTnE3+HlEJcl4IiZm6Ya92MFrmluq5NB8unesnT6ATxZLwpsjEbXD8jlX
mL7gzJyiyo7MD3Jgnc9liCHcSwt4amtDgYPxKTE5+QmEEclrNzpnFRh+2VSfgy6o
o+VyhI3lu6dldWqXQjY5AdGCCKcA8pdHpiAey4VyxGHuxEGrIt3yijde5TXMFfMx
Hy4TPSGPV+dNGo258DXpA01Tcpwbq4mzF+vlfL4G9lyktd6pHCqEBVPumQjq7V7g
6NeKNX+i0p7ikhXmY8yv2P9eCHIK0Wlk+k7J4Xoin+V2MZ7UkHzpMVYK+3kU8E/H
rz4+RGCXY+nKjmQ+0lNcxnuC0dnMgfKDEIJI0YFQCKNQdwasBNDlso+0Bxq86i6M
xAkbs3Dm1GnEvGXlJiH/E8+K8u3XUXaVP48/aoQO3PdnBTBq0EjlyDdcFbxJgfwz
bbzf7XfuqRyDXda/3HsIoV+lhGkrjlKDDb8XL+ZHOFQsHzSjEyPLFltsV/VZc2/o
NAoD/YqAyzsEA5wFuL4EgWzNYg7X655E2WZ1z/cAVd74eGSJT0VLyEFV/OWz++FA
WXxyJsKhLacPDvsN7zFPpPK2JPYTa/L4R0RS0Sl3hD78ivfh3a5b2ypnwB2MkHms
7riAabG0c0n22lhY4Mc1kIMu2WzhGmTEyEx9zTBLDLsDg6alAzDjoklvr/NQueF1
2HcALFKtP/Sz1OlUbq8qhgCZ2OcNIUL/yMfaDrFRKRn3K9nPoVaJnt+wDyqRLMm+
AsIHRxY9tnkTpyZrUN9oceABk5jAZVrmPOIu1goTpukR3+Mx8ZJG5BsC4gBkz2N8
Pj0s+w3JfQ5otSf2B2Wro1ECqVo+vymRj4bIkIXWEXQqj80ULFCnAlGgPdhK9O62
wWYaFoQUaE/kfTbW2uPayfWGb65kx4VxJOmwu73UtlCf/l8NVcM7qLJ9UDZcSIsc
JRZdCo7cuHZcI186DtINKXuNleRhn/bdo2ZmwUXOgPdRs+1dcN76jcsa8uEWpcWf
flk7ieefoiGOw84DTTixBaw9tu1rm31IFI26ZrUIXaevZLN9vTAZwutHRiGF3r5t
eS8vy3k0JTWuUhgh7EKtQadN+JfS9nIhh8KJm7PmuExYMisf7QE15G0AATJjv72y
nTXVF5jb1LFsnEylgGyBA5+fGKU9H9TBVhNuWVhN7CKvqFbZHsdZsXEhK32H12L2
mZZnVTyTLFd7QW2gXW3d75jOL3jxR15ng2Sj28rdHVeeiJw4G34yXsow+MT3iji1
9eDoapOHrzef9pSC5H9mg7js6QEUxLJzXbEQO+QU+rQAgXWJIZ6SQKM4VJFxM1zJ
5HNOfHPvB/mPd6vseU+zpFPnuQ3sTHRPTta8THrHJ8Myi9jzL9GCcpABNfVTJG0Q
TkHTkbGTQyTBD/53BWQmSy6coix/qK+j3GDF0ShQx5sAsILsQ9qTE1W5uRQ2Wrsp
q+ssNmapWx/AruZiHbBp+KsEny9dORm/JgjXCPsOwQlhfu1SqVf5v1znBLhxmSMo
JBMRoE0K6HMPdoMbaM86Ryj+gODfpygbjzd/MSKd5U3+jgeKqd4hZh+aFuqTQ3jp
NUUn+S3ZA1Ytru2gJwravARo6PvFu26kF13JucqK/rBzmbkC4z1yKKQgx39iZdXx
CUP0ZKWnsNCrix6k8XmrH/OmEC4fTH3MOC5bvRkrWT4TyXA7EtjEzzaYcDI7dLfT
PytZ6BDS6cgRqdT8f8+PYxnOe1C4h6BGmoeT5+wVE9dSmsTCeN48XEW+17l00TS3
aHKeZXLWPyeEe7yqVaWEixCIG78sT9m6fTOSFhwdIUdm2SPTrmJTFv60UAMgX2SP
uVtOWfjYQqqmaKEFaDA62jsGJQ2PB+LQxfm2aUzzjuIxR2dVxD+hpU/mXmLcFyHE
FHUF4kX13vMyj9x5V4G/E4wzJZKSdznE0VfSv8EDcFPqbZU76ERom78mwC34aR/L
fzqGAAyxbf95c1r4BAn8Fj4Z/98OQvE9I5oxmnaT0nkXDgyCzWkhwyrgX4SlCnY+
ISJ86tGPesQZ6/wZnAu6qP3k1XwSTh9l+uFhPQUEeJXzrug6tgMaLmfoeaCNXVTm
t2kONIdtZOU56W1Ok69HFfqFubWpCHvv2D1AYBt94QSsPh1sNsXzxO0NxDSsZur/
cmh60pqHuRfuAovwaSe1VlS5lK69LmpcmvF1px19BZIRzJqg7XLMU9yaWoCI7DKa
1F05PxrQHSEvZ+u6RDh/Y3F4maLk6g1MtI3GIyS96OCI5qlYTRiInPA7P1gNfTn6
+2eb6SZi5nkk5z0X5a2Z2Ys+hOeY5cAgiW6be9rFqaVnMtD0K7Yr3MPUiyjl4+Ll
25gUrPdxIwjE1sWW/JQvONG8mdoFceMyUS/30eEdkZVZoiobzCmskIPsoIYCIbcz
5b6ql3EpuyRbdo9OwVClPs/FyyfHBI6pBWGLe3otjIHQJxM/CSDapJjX7IAC6Kgo
1FvGBBflsmVD4ZKVYdP3ivzrDKYCmYfn3cjw6PC6IDFYTqVshK1rcPz0Jo8esOsa
pLCH9ejdzSa67/Ak8tLj3nMbdsxTq9ZU7BL4lposwHpmnnzSq64ofMQyXnQf+1Vo
n2lipDr6X8SrTJSibeB4Pm6pOJ1e/vfxTh9IBYW1sOV358ssizWPe4YTUzNvbcpj
up12aQcdsJPETQ1wMpWJ/kEuP2bBP8Ko0s8bU3+fbm3gEJlxvP0+iaPMFeKUjKGZ
uSPm2XmMQ/zdiEtvXEbVRMu+k/MBh3bXJsdplIKwaOo7+iEiUyeA1VYhuVBihJqc
fKa5LqdK8Lzheipvu905crfBQLjf6xnMHI3xkO98FTLJjjI8cL4GMTQTA7JwmO1P
lfkLYdXnqBYmvAAmkx5pFYdaHo98pobb2W3gFiL48/GDaLknAkGptzHmFV3+BS9X
zagFLG1vzuPKWcSKDDKxKEYiGiyKgx8U/b8kmRydYzODJPmYcE9/9YiK4KGotvGO
MnoUHVSmHe6UtY72BTgeD+/pUssT5Y2Dchb6dTlCcqnX+Wlk77dQbvu1G8F/rP5M
tsEQL85Nx2OzZpwJvTuynPIrRBxzY0lLUB904DVuzsO7u7C7H0Bz3waGx+p4RIOO
+uvq9edtVWJ6Fb5wz2DJhqBiFzde0ERrA1WoYM9zWf0Je4ub+wuSzeNt1w33MNRs
PW6OoayyzBArI/I9KKQID7ZCgGfHGsrD2kObhobBv9WGfu5+40YjODPXv7g87du8
wy5gA+dUmB4hd6qv5iu4oK3V7G+g+nk0PL3X+UkORHaorjsm8Sfmgb1fIaMvIeuy
FzbuTYnYBY+yTxeblR9S3wSdE5HzUk3FifSTnpg/D0wXVRck6x4QQ6TmVLa4M/8/
hcsM+DI6VX4k65AaxSSETUViJ8BhiJOjclFM2skW/6snLY3Exv0Zp4L2D7Ue5wcW
9VWz7hJotUU1Xll2lLewelchwl2k9C+lkWh53f4oiGfRja9iC7n3dy1Px9MD2fl0
oTMWZsBHX26isYM5XHZKbxbl78KQe/T3uiA8NvRGt0ViA7lYSj+pYlwpetWZzPRP
yBf5+uFkU+FApezf++eCx1E0Y2fHKZnT+872PtCEZIbUfWnL03V9Bm22sOO+6tDG
LG42cFVpwTn2v2yee1WjaVe6eqmTaXrC+iUQX7xaovzpL40JCGuLcO7nJbPMmo87
p/jjBaeYUnQs2s0YU2nBVYhtO91JdZa3QgGiETFx5LtlHM8RaculwKLZX81fuYHB
nzcde9FKUrsXDVrZKAL+jU9UzVHJhWGtUTqCf0bGgSY3m7bHIhM8RblSU8CzNok5
XqHPLJORfpAoIY0s+tKn92hTvrX40ptz9od6QX9qwoSWJiHkzaepseQKAns1Q34N
c+5I+V7xRiZ+WpNZmeSIGfMeyIvae6n7gweU95GzMSoWiz5kI+bedJaS2GdlVWPO
eudnfpYTvw8YWauY/qoWBnXdEPd0Ag5dOwhAFpWPcy/LFKBKfI021hdquJqt7zIQ
d3EBk55JyLauuNqUNmrUOFGqyS1vmVEx1WSD1jQDY7dMimDh48Y8+rnh6hrLz2fH
NU+lKg03BYxWQTUVLmhiHbjpvTOK+qNL6nltArxEk1EZoh6D1P7nYJtsIN2e1VOe
PX8GcQassHPoP34co6aSw/Ctny7dEmO/rlte8NZWcb+kGGpkKJLGkdFvmlrzsRcI
GeNHZHMaGF2572PEw1aCtNRZ9TsFbjJ83ROsOhnSVlU97Y8iNLrsRDl66oyIJ0vW
TQrkcXOoByDSYN13KvJKMF/qX19+5Q2vX/qZwOl5eidhOudQ1Gs9RXgOJsk16ZXY
XDH3nvH6LMZ+8uC9vadO4FkHpyQWNSin9N3nEMBORxm2DkeRQUGnVwuUgLjwp3l/
NRLBIvFphUw4L0sRgX1J33HQw449O6rqH1vtJjggnwbtCUEMLpxHRyvSO9n8nT/P
uUUwh5fXYZr7t2HmSNsxWC3hsY2256y9JlDDmvdUsvfFnytzN1eeh4sj/a/1Opvw
YsKqHubBN0+6jjy0frHPpY/ssFuJ+9lWzQFIa9CE6D7P7bmrgMVEUhIDgjCyRc8t
EwFSQ9ttOIywWKceFbmFM0X3vKR/VMHjh3LdkcH56zvBxNRxEs9Djs59oyxKhtRm
0vezXa5/FhnuaVGnoms52CP6DvxCSSjSRznwf9Mr6E3nzdQFC93I5akIWQP/q0J2
Z9KAErXSJnVYpC97PdgNyvfhli6NuBK1D0GiKd3MHhdH3DVQFeCFHLKSv9eLL6wq
wItFpjXLGeqO/uW3nUbznR6WUH1jJGm/Z5q3Tapl2lu1D6tR6vPC7E0ZFn1v3115
+kMwG/nEkX6Dnw+Ht6T8EdrJRvbgpf32S5drFik6Q52RzcWFPstKh8ZBk6tfwIh1
BqkpkFV80bHbGHbDqTX9I7qCYK7a/ghQ/qvjhRZ68I1lA+uj0V0dnEl1CUQ3yJ4I
T6uCCP07HmLiDaE/yJMz66KlCiOal18NAiS7KVhIfwaZF/JAG4tc1SAiadvTZMt1
dhOh1FcTN0oDth4GQ4Y/jslK+DXS8JBVc4KCiwu6FU0woP3MmLfozgeqG/YaEx4K
mj3Yl+1An2WLRk3Jw9xUxDoXffQDCD0wBnqS4dbzQJvkUcc0cQYBmAz+0vdyrDdr
DM1OtEsB8d9CDl0H4UpcDrUP+nvkrEOJaG09XsUCVHUP0vrBeuQLixkCqwhrKiJ/
jjTnk5RK/aXUU0ufE6tt/NhuyFyWdLPj0GAs5nv/3/oKNLlymnWQngm3bmtj6c1V
P640BVWPiNwNOjJMegidaR4CCUc2T0u/2mh+ysMSSHHkqbrgZCVVFGCrA6O7bSQr
L9msis4VYMF/2thmJT9rXpRQ3X/r9YVsRoPtR6cECouGSCpWMviANiNK/W+HKZqP
NZcX05SBDxApCzhBan1e9MQq4xW8yUvdD3M0OtXNN4MYIpIBXMeC+mpOMOmmuAp0
tFYlwgNZh5feIH2g7IXnpRmlvTcrP/QftiH8ZnwGvaMsOXPE4Irt8FD8nn4pG5Bd
u78r0M17+db9NMHmSibUpIOAOpqqNk3a8KyOKxprGyfhd101FdXq0DY+x9VxHFTl
WOgnGO5w86Y6eUUTDDy5HkkZ/d/C6k/nxOIJ55AlhGr2lMOpCHyGlTp32DKiY8TX
8M3IpQemKGGNeHyBflC+//I+gE94G61dHbBt4n8zxRiOPaNyO80FYLT/DvLly+1B
3L7Y8XSOdpLraNUBv10jnwBO7yWlNAeWObyLQ9SRij8IqRwmd78M01mU1BRwcGzi
AK4z7LE7vFC7oTSSf8vy/r6xteO95PyPa+DqJY/pZFGpH7k1ykH5aeX7PBVZ5UrI
WNUWT4Hlhun4oinQ5xwixQUiAc4gc4NUnc0lY7Iqg/jIJAyIkJyY/sbHXEfRHViP
s6o8CRIjXe7TRQx5QjUGPAhJ5bnAOIlwhPh71ovWdE3DGP3AaPqZYXYQCVBz6So0
DiCdzUi9/DKa69vC4Glc5hL2O6ZcZZlJU8tqofoB9tSZ/dLkgwnp+8EuQppIL1gN
QeT716VhNxgFdnjoAVLEAHOnHCSwY4M38NyL7aP38/JQ0zhowdrkaJo+zecSa9vz
Nf9hMQkEtAcUx+K16ifxFwGGhLicCVDBz7ubnGDRvQDgS7t8oGhTzf4QVGnYJiwf
fNMJTz1lnSefCYPA/4ZGVj3XgiBPb38tO5WwLf1ptHd3Bqepnm/w152ScYecp3ev
fbovjKvQ3xJeN7r4GrIzeo5QQfiSz3cmLnEnr49e3B+hCpYvf6mPSh5Qgx8/rQqI
9YDawx0qdtyHWHHEduiMUFoOe7HsuRdpBUDTzQOxuHYEZj5mDA4p4+zuwuc5AMpV
9ytKDLZIUlpwu01YLSB/TUEAjdXewPeN0HlkKO7MCV91aMKlIVrZiH9tgntsc0Kj
u80Yk+huv1EnikKHPUdeVIEy7wxvDYAeoBmxjf2EN3qHHDsS16dLlGvxE3LhVYRc
71yIK4cqLfaiq4pssSYLBnzgzqk7GA1UeDWd5g8gN7/lQxs/jMVJ+PyMyepQh/+5
Jc8H0SAAEQyPVCWhWqzOo4tZx+CBV6yYCMWSOixfpCotNWystjRxNoP0G1wY5YFD
wE6B7O0OWCoMbyTNnvetj2zVOh9qAF/6Uqc8hkX/GuwnfF8jTCJA+EOal2n92OpU
3H1n35ojBA2erf/Kdrbvv0kZ4iIWaZp7r20Lcy6OiOwivuYL4XsfYy92z6XApET1
xb8x2GYVxGf4whXVSqKH7h/ThgUT+KEqsULvhmlfikRg8WBTmBBrC4h6n5fdHPPm
ApkLii68P+bGeygyI8/ui3u8qJvOCV191g8QdeRKn09LG90hy6yUaI2OLYTCTkTx
DKpQsxeHjSIj5LsF111jaQhfx+ikQldjPkf5dWJRewmg8x0cofWLObKLKELwUG9E
cNcGdf8IYDCHzuDp3KFI6qyBTiHNuGv3f1h9dJpmr0f23g7C/bT957xV1/BilcPb
L3nfexKkd3vX6OIIuZBUY7Mh6B1TltRoYhlL8LSov97xrDKNrmDpdFR/sJmi3V7+
UJE8Uuy6kjRLjB67Lg8Gv520kBCO7oIhcT2KVYBOIP97EGDGcJ0k5LtFPMghW2Xp
k9iOyDOSqgxGXbiom2J+0J0gB2Funte6N5J7u1yufEUjOpEe4paKZBq1g1ylyrGX
1NfOyPDWLrYO/WwvWDimbZFXoqL4sy/PxJ47Z0tbEZP7bDmJoUGepesRQ83nnew2
uTxpm5E+AeMvSTjDBWa3UUftembNQQqm+Ue1xu6DQETL71u7fll5IP9c7n40NYYT
DLpshYxg8MzhvI83xByTt+XhTW0tJU1AcL6zgethFaU11fJtVYnU9g47Mg712ZKA
a3Ai7GD5WAjhZKdMvk7LGIv1e2nHTuU5K2sD1A8Nc0GL/GPUsugaFycpi41v9B1Q
m9a8juknhfcU2vspIJiZpncTusadt4UC00pPUDPo+kjoK8qfP4mDOgoZwZMAJJwB
8E5aaM7aN4ci2d8atVKDu6vHfsaC0qeIvW2zAWfxHWeTHFdh5VWPQCNGcD4ZAdqc
vinjNpGFKO7AmLvt0QoPHNgd1h54n468C29FbeKjBxJN2m779SjPoc/w5UlFjE5D
ZVDNS3I9bop0VcVx9hDXbImB9rfEyYd4qfCF64dU8tyUVWsmr+P1+M77urUnqgpm
UcE6RZof7vW5YSMgbu1BYcmk2qp8qjkPhe4AlLFgC1hCb3w6zkTbWZX68qixg0U0
Qr1arRbO2SzBqQfLIerz8/cfbJ550+iAjPkXbSK5izwTBQ27tlZKS+MRdo3wyh7C
/Eyb13oIKzR/qrQLIjG/HrUuq8Z++A9glQfsi5j6HDJPTdQWgELqnVvT6CYeiVaW
fYZxRh8QK0l7dh+ciFjv46qSaU/atK6fIf3IZzM/Na0z/vUi5VQm7fxx5Mn/yNl6
YX7jDBvic+nlPv5n3mvA6L6sMfc0dp8wafrAuzgQHSMInJMQz3tvG8xznn2WwqUI
tF6cKmH+IYmBQJcaJypqjF9IyC4sQVhyGMHF6xEQQZTY17Mb9JKXaDvtj3dZb8Je
WB/jTSPFgOh+aOPOOhEnIaQd3fVBxzOH3ZyEAty2Id4yi2/rXcHqOo+3ANft0SDt
PC13Tz/cCeF8vkZoYEcdPO1vFPAimOmCyqhioBFxw6N+ED/Al4xI2u3edFDlfzPH
ChKcYm8PMag9e98EP+h08TZ0mIaHNmy7ywa0Py/B+9igr3D7R6Rgqe3xBKb3v8xs
zr3JvymItKTkKzAbFARoJVSCGQxvfEvx0G6rHVhVZh52Cvd1FdY+ENR1FhCo72KC
ipak2YCG9jl/6SauRkyhOOS1YUtDNP3k0h8UiOl0ur5JNBaqPmrEZmk0qshkdwXd
mXwkB2+kHxenq136PaoXjM3p6BwfbLrCNra4fBpg1GCq9qARUnophZV7d03eIJIA
OaT6oTGV5sy71BtSOLeFKPpV9F5A6ToNS3EH9ugf+VX/Ew4lOzT/b/Y0yegv6+YV
aIaxie677Gn9snT12BIihpzd14uZG1ipSpJFE99h3grHu2oh9k2qllhcLCU5T2FJ
mYuJfuw74ckS0y26QhKf0Al6tGjG6COK02TBMhi8pHV3ZauW5sKs/e3j3By0P/Ge
xQ3xg+Y8D+R/aAgLkGYjzvCyhx6Zoxv0x4956BFKx6TScGCc8JpEyT2xgPQ4AFZG
TtTiJBIPt5ksOdxFYJuHPe5dneb8Y1s94BDrXec0xX4663Nkp/efE19HDNnx+4Bw
Ocg/rts9qSR02u5fQkgea59xqEHDJSHg+uB6XI1hk7BO9sFl3iy9iFE30BqCcZeo
CBW8rBmpgHC7jsylR3QpM5LEkArpmXDIEH9nL9IS8ANjCBDrW2WuInvdzGq70we0
wopGpFY7BjJDwC/4avbMscqjLKPvOTdmPqgjtxQXaHV6j1TKtcNkHFPaDErfK2dQ
mjmao8Grr96bl7oLza01wnntq8WlpM5R5/w4WJ9c8ThX04gp1d0JMQDznvUs/Or4
OJDDCvvLkLo1Vg4U+TPurfPQ12eXbhsnokw2uVtwwvPzONJuliJv9o3KpIAlM3Xz
p5z+dFdCnQBktUNVT+RIojO9fSQ7ItQtP1pYzyR6/G4lR3D9U5qLXEULMeFJVqeR
NE7s3SIk649XT/5/3PI6PLanW/zvzdtc1HMgF3gGmbgH3S2ER11VBJf8kRcqTgrZ
VmtNoQWdJQYUMK+ldxRyqtxu5ZeY60xIExihEe0ZpiE3VICucRmRWZYYgAGoVMcm
l7YXenT4PNTXUsNJcT9YQ/p4IYqjDhddnqkavZXq4mqP2Zyvfj3N8APwBQkUrxbv
AB0FIRKHmvoHSgiLPWAe3A4Oo4YpnfgoktpWWDdZ5n3TYfwNjWBkKv85RordfbsY
g9Eu6IvdNlhT1C8OgE1RbtcjkoqtNF9QbySJfjWnAv61OqQX9pQjzrW4ro+7qc4h
M1qAPmQaxCsIKw6f6/bopAHsAfeFbTTYXcKRxj41IFSjtVhHTzO4YQwHptdVhVlB
sp7ceeinwQpO9KMgsqcZZryTsZPkLv1rFvO90KxJ5B9mhgBq8muI8FPZ1qhPGLSQ
7XjNoKuDAbXqIZQ4sJf/eYlRU6ikEbWKoj0HjoQCxBEU8m4D5QWMSt7Qxu5oy1xL
oh2FKWjH5Trykf6Sb5PGjhAhhhyzDtwSo+0oHljgPjTFacsDkEg2CwatLxrk4tmR
Hfb6SZzVk4j1+Y9YELy7g52h4WbaAQDbgW+d3z48urXKeaYv5bpSBgaB33a40yAO
p7WqMkYER7bCETw7P6QtVYWuLslPxsqkQ2hp7FKdq3js3R5xLZ0k8az6FaTeMvFb
qx++0MmT05jZX19SlFcmFRO3+q+eurvN8J4ernaIhQKjaizFFufB3M7FV0AGeHPN
sCxklEElUbp4GZP6fyewQxteoAa9TEjoEvEyC+SnvI7qTTnZBaO0aTNmuQKtvhFp
DEBFvMbbGtWxxYgCOuvf1CxxAUbaJQlR6nVyHOed/CDuYXOOoS7suUE9E2fOExgl
lKX2m/2Y2xtB4QLE9Ja04bXZahLq5q7O1JALjwgp5WbctyhreGtd951HB4BZ9oST
EiQDvnZqSbv5rbtn2vtmEeUSof0B5ukznXp/2gQ5ajk3J5zmYHTwOm+fIAdZXdTO
TiLDpOquV6JkivyhvDw0toCzG2AN0e857Q47IMDDc/UYij+zZV+ppfTTJNAWweyl
HzPKdzQoxkk7WJYJcKYTe3ayT2txk4YEUQYneDnfDIh/bmM5DJEU5cVFW47RIEp+
thqyLs17o6kVNJ3GHcgr6WGR2THiIfB1dNagC1TsKxs9BXgv10VULxuWyW5I5EWD
Sb+xQBaHNvt4jIe69f//+RrA47RI3lBrMU5mm+Y5J3vj3Ah9t9gPLSSq6M0W5okx
Dbcd6NaYr9s9apG2Gl1tErIeDyx+n82NyRG0rpvBzj6RfDx/a8e21vN26+QpUecp
axtc4bHtJXEm0kZvun3El8/Yl9jiNkpvr9PFMQsBChuGqtrYBtPGJQOexumDEAhP
dlUseOEMa83oPSNNArlaWOVkPMiFd8/+MuMT4nW/cB5hcecMYr1CI6ytbEupeiBW
82nnsVHAnhb1Kg/10bAYIrJRnVoO8xmSwaL+Pdy4qx00H4c+jAtE7OBUpdCjJuRm
c8opXr6jCa9myuePFX0QwYqiUz0HzELZPYrOKAIuRhS31E8p32L5DM/7GW6yR7rv
/2eKyr0k913Lxt8qOENUt2RH27lNm4JNLLb1NdPxjkM+Jj+qc8UmzxGmrQtipqqq
6t8eD3cUOOiqe+uGMmGqrpicrPlZpu3lZAj1mCsj3mSK1jRILGmMw9Uc1xU0uLPY
ae0HErnFDVEzdbUELppQhRyHsAaPiqjUB91hYUWeoYqR/U2X0WrBRzWqvOrqPnZk
3484GdKRfdv2gAetmXeBkb8L1dhUG4fjChwO9Psn3QduoSlLOrFQG+F9FXMerobL
5+VgyMapVret8LnCJmQxC657KCZcw1RxtkM9xlJMHBiqra9TUvhZzWlrkDVMcc2s
hOy9PZg+4JkEbKmOCcF5sNdaxsLtV5594CDsqmxM1Ro1Q+x92/tZDOg+VZ2ZLlgn
KA1wyuOa3ID0GcgYfjFFA2iC3PVnz4nx6dzMyGBc7B1ycijhVzTCFwE5rEC5iq6H
Lpdqjanv0LNrCgc0B0mZCqFnGHjDvtjk4phSZUnQcrBpiScRC7e110VAVj3yCGDg
gEXl0qNTBHoaNsbqeeHRcde/r2tXoNBB7nNJHKsyVvCMWDQavRHKqsmWj/tOcmOZ
7oK9grjMhZNqCWJhAfnjtbS+KeDMqHTOMGeDl4lvdlB/PiFEk7370E8550ivCz/t
U+3hxbmDmUsB95ZqDSsLz1DsxiCNQ0WT32xWJs+g6cMY3W1CsgpYnzO8c6hLFxYT
OklT+09wFyxb9gZHJe9G5DM6BQia8toAffckJcEc1tMJyS45k2xqMmdx2p4bb5y7
VS0+rTbEWrpbAwCxgV1ebNHqOFIBzb+bl7k2WaEU3DbPb6yjOQRkyl9ZCxa/lpQB
kWzKTycjUajmZS6e8l/Mgp/hjsDIAGgjCuKYkZe4V/8t2ZELUTPUk8rAeZAM6IgI
X7i6a7sBawn78pKU7jefHIIjxjllv9er2YWT1Xfp0OuW5/l8uTonF/Mvc43WE7i/
tD0mo/48oJf3+8wthZ29dDc1WXEJakEk31PnkLMj6jKwROXlKpjdDGe+zuD0MTKm
YoA+/qxFU3XqQS0fYWTDpR45NpNX9lOaf2OeHwWCJQzx3D7fspTLjeofswfkERua
9EWPhuKc8vdabdJJczCx2w+WmaKep9WtP5Jq1cqRAmHP8h3Cq9Uoz7LBeWkO5z4G
YLFVoX/XeN7EzWAtizGyg5tFhWf+w+hFCWdnAsysytc1VdOPbBFZjvybu94+RBCj
WQoepgcxvqLO/AM9Z8X+r3OjGkIWyMwlI2V+Rp96P5T70GQmGsYKkpqpx73D5CvT
bfrTUlSYLYeZRcGSQBpqB0GEjSxneSwWB0+d+DlYJWq1IjnMKDIlCikWetXPZ2zy
NazO8a5OGkNHmillXOKo8l6oM4HQYFpIQu4/x4fHQ4MV39OLnGFHTFH485s7y3m+
ZXHH76CBoXvlP7DcO3HMTqziXnFYJgG+5Hm69RwvZ7qewTeOrAT/Aw9ujyVfGPyG
gKAakr14+NyTl5ulfibYjuWLOzifzHHPzcYjCMCVAu+jbi0RfSxFg8ndySqQylPY
iA2eSnUEgCqHzSwIQ6aULNSntImUzf5yqlseUMHVYoJF0AjzJ1UkDoo48ktD85fT
6BON8poMkmBMyHQL0XK99QWOIiZuZm5Jn9omIdxWtUSZhrUyFBVjixaMC7mQgdjE
Bnzb2EJXb7sqtj6AGyCeG/1KEdwmuT899MTuARJwKlfAPN7QSco/IbZ1Y1UBJLV7
r7zvbAy/8irDuu7CdawAhIJPl/UEZd5Sz6jhMbJEgjtNPrQygTAKe2Xjf1SlX+IM
s7phPHhlZTeE7ipI/bLJXhn5DGmPeGDHlY9gUnepGod2sfJ4NcYd/ziIvjtl8Sf8
99i4vEy8D+FxmlsXs1hQlFG7FoXPcmTgzdTVio1foevy2vU4MpS9f1jkmOKVujUG
RX438g0iIzDuLh99EV/elwqp/mriCe86kHn3FRxnAFlo+JgsSdZEHZIzJQYZzVtF
0PM3RLy5R93V0ekV1OnbB73gy9oKy5KXPMDI9fOMk0DUoFrkD84qrOJWeMLdpKhR
lcAJZ2f6mUWKeoaT6pXfb9fxe+JzghfZFp+P/czx/nB/CtJEXvE6LBXZKEpr6kTb
nY6Y0aeXhIeybXK8Ca7xfJfvUuT93kv3/syQeE00kNST4o0/47xIMBm5azNp/Psh
H8s8IIEfc+6Kipzh7MyhYuaanYkSHOI+ovnWFcla28epRU426i8hMm6Jv7bzJc1H
gyxncjHMIea1hcuaWHM105GYxMeAVEooa07efmKN9+C+OlMhKxKWvlG0Y3aLNLyW
dT4UsvV5I3npWfRapJ4XhG7dN/rHAZ6A2sXstGxorrrmUe3QlDurteCmMSOs69tF
dqBNlZffoWBRQD6tZCTU569nEHI4ML1jFUo3pvC6ZJZYqsIgTAWfMysnC0hTU3q/
ZUHKIvdL2HR5cn/Ddr/H/4Q84CQNSc7lkcVzdwmyA41BzFAsHZhEec0+LbPFJrnw
XzGZ2YWwLoe3ZdNdAc/mI03Jx/ZOnO9wvnN67d2mVW7fnPs+Ivl6Q1SMCf6TyhW8
I+Prs52YLF2TJQETkX7l/LIuyoIBdSTb8k5Json3zErX1nVT+eaJ7KiKnmvw+xto
pGr36uDIv6TOg0AJywg9FPb67tyCkYfLFM3PVLChgPiLrg5D9QYyzfNiyk+ja1d4
oI2zrZnB8nvljOD/5yBiz4CZ0CZl8o0DjWMWBLPSjv6q8b9gDTfOdyAG4D/Oe5Mp
brjE4Jmj0T++qROxw0l+8+/4ZsrNazsrWHCKRRo8VupvomDm3yafkK5nNPd0geep
/hBV2Gy3WZlIQ62ZW0xwBXzEfS86E1oBcmVnnfRiAc12xkdB6RHYTtc4h/xpu1kK
vMpclYrllQpGxtzg6r2E/JBR+ZVOJnAd/1+7UsYcVh5d3qZMoODQt7BrRk+yo7KJ
PHzkBadSYboqhA4EDceh37A/ndg9YUop/P2KI7JeNSHmIsbh2I9xLNS2sjtIuz9Z
CL9FwT2OzB2zcGiUgRENWqDJOKSxHdneJ94/rPdAI+isqxgxb8wpaHNc3N15gxIK
IWnp+O/dEgDT9ZP38Hz+BE54ZvcWt4qOcrHGO7hr32h7T/ZUHTf+xTbh1dAUFEnv
iglvHhB95biipvjHbWJ095tsQN0/TMkD9TYzyvAr9TZ5s+meKByVq4Z1Wrwkxbtc
ce/RqDNd2JYO8SbU9ICjA3lGUsFzs5UlXHETefEOsAtdMjpGm9xREKTkO0XcmfhT
MRUHSatyfYocslNQF8U9HW9TsZppkF+fD5zH1SOkiL8ckl7RIyb/wr006Xwn2ZD6
zeqSjl7WHOKHcc/Eq4pkqDyjce3vasbRODB6+6TZs22Ec/gwiYvYIuu9wZt6O6JU
tR3qwjFLB9/SxU7dggKjMW7A/tSOzCnqzAJDMCH7NmmxxNFh27QRoF+2VjNKvVuY
JD0VO+mS6MWIkbXwLEofVobTgPPueWd92Vxiz7S3S33AJi1oz+zCzT2iTpod0LO8
h4NDhP0i55tMhZi0VNCiEm9ShjlB7wdWMUwGSLsrgW3+RVsaoSKsvGdgZL9XAJsf
Yjw2K25vdKmZe798rTNJgptKt3apH9M63xAkmmtwVGio4fePuUDNg3FDiiuxuPJ9
sLBCDzXKH+DayyAPpXtfA9VBppfyc3h63az8F4CgdKsfK2thkJkjAwC184Nl0FLt
+YUcQroC642tEoP9be2qYgzIluEeZlhKSDBkuXTTLc8B0Ibdm7xBZ+2OVuc4bega
VJF6lygkKJsh4RmId18r5/dhL8w8CBtZ6FvKnyaymA5Lt/MpLdc5wY54ckfXC2MT
unsIz9J/q60cJv83CC295VDYFhby8MZC4m7rpGmfKjyDzuoKjCXyD2/5gHQBZ1Ao
IlvN89RWf1427DugA845Z0VwN7KH+vNteK8MnlTTjuQ6cKwtjNbl/F+a6Co+IXu7
F+RHFiCd3NZ8XA9QUsjIWJLAttufCsh0w6QoqqpHFuWlkEENFCryVPd1uai/jTVC
JTfROCL6d7QrqIj0dQgzNjU6LLvAdjY3mJNFcVXOhUVKXBMTwhSF5GeLrVRyfVZ5
QuXFShrr/WPyBlHAVpgPaQkg3XpxbA06aJpFAWGGfekUM/X6ai7FcnQzxUl7s6Bf
T/y7Ejw59Je3ppWDlg+RTKlLZeff5THoO4XkEWNtbCiPNYUls6toLTR6h/dr4UYe
HeSi5rt8CrKt1jSkddbzsSLkECeE7ThzdZ44Erzi3dFYy5hNTXSAbjiD/fruk+OS
8lt/470u5qQA+N2XFbZOsFOPX6kxCO553LSckrfyscAleq5CpiYZkmsYRx2saCYR
unQL/m3+IYyp9jjwc6kEqUkGH9wK92ioID97ZqyhMeGwdCxEINeRbcJiIX9h/hbH
QVtagOw7LDzMQVpVJeirIqXPLOTHaE6h2SG3YKVzPRNTsaI8Jl2I3uVKKEDwaaJR
bQqDfeKUXKRLOO5LLh++SnhJ+mkVnG72wMI4Nn5uRzcSMMPi8kTunpUMIW4HikzN
/cpjUigMFCxVgXVBfADB4KfS67xuZ9dYaki1TCI5K3XxYtiZR93m0Sd9+9iBnA0J
6vFLuZEo+TQvwBCl/okbVpWrQ+N2v4fksXBiuq1FSoj1RzWPKzFqbNYlgEGZK9zd
pHYgg5c9XDYoVzA404BkaXpKaeOuFDzfTPwHZUX5U2Bvd59qARZ5nhPRdApRcaw1
LmTMoo3n3JufytJoMCGxAAnsNBv5LUaaxFDMHF1IARHz7NDePaP1jlYWzqFdXSIF
czIEOP1FN8uyA/PADmrBraUJ4kCTuRVfq1nJZ0M0QiZrAbUPdOHxhBfjLjy7FN2N
vQowTsdJaAWBYDQK4S/WWvRa3vTjXtFyHuVUVj0stUbFyPV0w53V49hn35wg3hEC
L+iSYK33K/HgGZQIxfPpPI5HAsBotU7rKdz1oEaQnJox/cE3ExhwDeDjRKVd3jLY
Fb71x1tYekxMMlkq4W9x3yD2if2TAKISeVhla9Q/+XEYLElQ1509d2Fl2vIF7mAH
wvJBM6k0ccqgq/JS6Urp3k7NSkgEtpRogF/pq7WCpy0TL9NR1ND5VmUMb/fitPQZ
6OayAEPsJTscG67iOI8IGgacsL9fmZgialHAULCmR/X58r6Yo5cB1X90K25fxfhx
NF8r5A1YR/QcxFTbbOfBEvrr87SFgw5jwE6CPlxASlnvA+HHvC20+vI/HKlTz4Jn
C4qOZS+f9fbpRvOYlHVewjRniVJM4ZuYneysKOkVIvSg+Sy9UwYeBMBJMNrXK8qU
iqdoDfmBQDKZCfqAKBo36XJ0cRSGFmhMzAEGi+CVMhAeIj+imSxdtvR6qLEfFw5K
o6ZB88n1zPZ3syhckmjc5o5GJB3dEHD3gghWoRXmp6t/PdiUXgH/TqhDv3jv8ocg
TagcSaUmf6kp3G54bn83KjQUkdk39WN3MbuZJOMbDTScWLfcGBPkcDnJ26EOv8Kd
7gNMhAmSRZmb2q8TiEN0WQ/D2lRk9zg/ohnkl4eKnbuI3S6mGiHGOdnSxgwqMqOp
DtNLjN4EKSBA5KO8cgEtzrGGzDzuJxpSM6oSgtdFes8P+E9qLOntU+4SbmTetJsT
cyFJoahoEX6AvlNFm01upCsVsZNe4zgmND1QtgsjrCxfKavvvqqwFtOPQYD1Fdou
pnVf4CuxeRfbjfUfMnNLK4/Cn2RnjebOIEjBYBOdtBNJVm42oVebOKbbfZh5Z64U
ExKYFdtENOeAb34q7cxbP+so/nhJ4kxCLbvYxmE+qTlrfqmQo93+f4yqkvtpJ5Zp
7Umjeq0C5f/4MzKpelSdqq3WYRset0I8HuUCDSdAZHyzlclgy3Yx6M9p4p1EUUnE
HkcZYbvOW7AK7fVv6WuJcZU5F81IkZWyqPa2n1T22FrqhUhdb/8rFVYgWxQxQ8CA
NQNBVE6/WmPkk9uM/wVZKw0qFXG2w02M1ah/Fd+Ay30Qs6KV3t4uvr3FEYk2HQr/
jbZXulowwn+NUaxx7x6ev4F1uI4PYDguEpg2xg9zIFErcKcJoN6O7rvXzwQTWFRx
yBjukw46AKXzvSBjGsk0DWpfeM5GZ6S4Pb3o9or6WFwPiDfz8mvjcGZI1/3ONeyo
agpI5whThQxXOHiItRJbkgAO1wnhApZyvo0k17RfOohqnRROxDkoW5L3Rw/UZfrs
PpBLC0wXnWbBatq18fB33M65AmIdOPbYkkyeL5oXyinUwOHNlKR0UM6mrCUW2G4m
FlAH/X4NRB2+q/V+fGsdmllO5gQ0aanOQvFu4rBi3mv9xe7gqeQIQ2kvifSB6LFA
CLOjwRJJm5NzexFtxhBtpGsjm40RFH0vp5Rg10IRzV/A9o0cejhETwQRtnULr0Z2
RUpFEyx16BgKP00A4sQUAaCKN4JsM8weNOJiFGugsy1oAGIiMxZtpAIHr2zp7oZk
F6S7HMAz4FFaGZh6gXn9ujhSxqSNIDwe5zS0IbbdG1xdEf5VyYDL14jS3/YTlXkl
hjBm1UePrwSPGt4Qqx3qcLtjDQjvT5xvPUjBFOg7cHR6qPM8f2VqeEDm3I7CmAea
swL80cAAdw7cnKu+7oF7Rlh1Sl3fy+RZaf32Panf2ptWq9zS7Ix8zU6XyCWAZ82R
G+x/lnYnJq7KczW3qLEKb+hPWmMYdvLboncDYR+BxgfEnvVzlMm42bSnzM6ALyN9
qAD7GOdbTSHzs2CQfkeNaXSOM0ryK96hAe8a1/H5hg87GIJgwLcZ5vIQlXW9OUiy
WbR+GROWIXtO9kxU8un1KGn4mBWsVYn8BCLHUF3eIlhS+KdTN89VUQMe9i1AWQ63
fXCivj9H9NFaag1aEEeAiYN4OVeG6s6UTaRyt95tTtrOrCPQ72JJlVZfa99uG+FP
Ee1gef0iKW8+An9YYxlMUjG2hgY+yUakFvBf6XYfR6B/W6HsChXdzbfGaX0gU1TH
zOjWE/29sEltU3Cia8Rzplqu3rPMvNutkk+SPGhDDtMrB8RZQsTVI/5vlbLKU8er
gD6S8CyfRcnib/E6xG1F4S8xJOQxWkiuHwPv/WBiE9212Cyk0BmRoNWGVw9BTKGt
SNM3JMdNzBkWMl6I0838CQByM7yNZ2r/R3wXlBQpx7bch1dqMG8zjwFeFWu78syL
J1KreIZtAd1rFpx4ssz2jE1viJAEO/u//0i15nBZVPPwCbElHu1n+u5aCWiH+N21
raRXzJ2TXN4Q+lZD3BHRDZimKhqxvXkc9O3iES1CqpweMhcIyInOFIo6txUFZRJ/
lcF2gTEEZtt3hWDbf8iq46bfeIMqddr6UeAAVdubwekyqR1bvB8c0cLzbtz1eaLh
R8zyIVrJD51iie2oFGI/q7yX8o7b4Oa5jsdIOyORqwuI9G+MZnbWf9KXcEWtdOc7
wsoZNssTbfvtVpQpAmLasBoHLxdSHedIBE8lD4r/xaMRdaJyavg2ySDnc18wRKtg
mE9tW6jdTvBB2ER8c3eiX2Oidt32H9pfR8T5nRsFdW6fq+xXFDrEtZepNRRE9zMs
PpzxaoLGjLHJceH/hjmv2kGA/P53fKt0hjxPgUKKj8mwS3n3315Bn2GzOpQ18XNV
VwMEgRb+bbQSY4ZAktWfYyxZTQPYtjZpO1TuDFEJzwulfiYx4Nup4kABoyVa1c9B
vEnhZGhml7Yaemx22BE6DAdkvZNkuQkZLDlZrhUqsxZ+P7SI9b9L1JOqEbAqCez1
Y3/KjZokoYmO5xwQcExrdm2GmgpjXEp/FIflI9rbTqvu8ieJ5wszkAzGiYDLL6TZ
n8vCP4xPdBeq/+Q0utzBt/JOvGI5ltPkk6/py36cWYdaDZFlLcvae98qJYS3e1O9
WRDPXZZ4eUlZm9at3bp2cmXovHhOPMXSmV9q5EAqsAqwFhblhrmfBspPfP9ZWoRs
Mu9UqtFRC02/iczd9kWCnSGbarLS+bbTqa2ar/fGzgnflIU8nbTZmvKyF37m18vf
kpJo4G/QRZOL0kdESZrBWhG7pHtrRHiJcPC/VlQgrvJfU0H1TzHGuY1NuL5h+F6v
P+jTU/pptX7YPAOs6NuAXwZUeIXtu+O/IA+CekiXZKFBS69hATRHZGWD0uCQe3Se
pYl0wDGWg3E4S50ikAZrZ0jV00iL4/5bQCWAQXsaqwB6VfnYIFrgJ0/Mw7Ohbfxg
LDSch1sI5Wnhvz05Z1bBr2HrQ0oOjCA7HeQ890Qhs5FPLhYV1RSqtECS4/rT8ioZ
Cxd+q0yvKmZlHKXju05JEH98WjGO33SROGL0CpnPXQs8eOfmul1LZvc+HVQQhS7k
LdKpKDZ+REmcD2VpJ/hndjMGnwbr3+8cjvfgf56OSYHxx09AxH9rkUPNvitlZoaG
VepQ47feSuB8xLOo9XXgga2tq8v5FptjFhhrXVEx8JjemQUNOSsUI/gvePzWE+jD
WaLDd3yYVUny5J2L67ivcv7sIoXSQWkWPWFSwgZ5ReGtQ1T3tRZNTonmNKGw4NZw
EzvpZC9uCTCAQbUG6rCV7DgBTytJrFJDeNUx2An47cUdLT+Gpbp0sCtWsKj899yM
v+7cMlqJ2UYYI9RFcJRc3Usx0ZMFKZPtRvTHy0Not4WVGVO3ETu2lSDfA9ZzTdnX
gUUmACa7gIUSmEZ0fd/s8ohIxRromtqrFNUBIEogcAQnrUuFhVfd6ryD9Y/C/fKs
PCqVvkwn1FrFYc8PlbYPEdCWCSh2UedsmXoIJGn5pz6K7luQJv6OulEawsQq3CC3
JEfHYeTBBeroZu6L9BdZnWkU+nNZDoxmVoE5UveVJScBgVkOi/Wv7uwhpgS+5LqG
1um7wvUa+engAo9aUJaWHjMU85NO6Bj5cKfr0EkXJdFww4NH9PwIiX/ZlqfdZMG7
ePOzzhxvIEriljYrycwzU0prwQ77FecSrTqlpsbzYo8tOY0ItdIA+63FBqSybu/u
Bc8XfD5Fi4z5yGGXte//dlp/or6mcul9nAnSq142bAz//XBRrwc40+vhmakxRz5e
1EPFgpDHs4Xy4CkicBjaIFVRolIcGUNCrwGe0IXRdNWWi0AN9/EB5zIDwSoeHag2
0c2hwkiNoFzYFW2pfKHQ6iLsF1bAmHrQamFTVruMmoOhVqw6H31exFipSyhsa1IC
9TxxGQ5D+mVDWwOMmHkIfz5/AZPCuT6T4UO1SaW3JX3+dEDVhzJTFMrVG8gojlu5
ETzuIDT56sxz42YI5KIyIi1HT/wbZ4QnmQBv+fUyMkWOYTPbJ+QMnDxBrLyruLif
aYFwBgz7DX3Vs94t7y5poDO1LGhE3r36um2wnPbgMdRJc7vFY2ieTi0sJAJwudSA
1gBk9vQsF3o/NAkhn8UrphrI09zh/CEx5lz5nATLImK2uBwE6ib6hR+DdFraBE9s
luWEsD4s51VBu1LqVj1gTlTGOfTqNZtadSM/pYflP13P574oKtA15Z7nvPb94AkG
G3h7JTdHB5jdJbqQbTKFVLukmC5ECUVXSjiGAtR1htckn17rfIlahnx03XQrIIdY
vkVuj0ycbPOQHeHnL2ceQSynvncC2U+yVuQfOKYMHz5R0linbfTZnWdsyboeks+c
GRrVO1xlBrCGnqfUX6ChOblG1c5HLOTcWlBq+Ed2nv8DQuTMP3frrdDepIcF4XW9
n8UaDuHS9NvUxThPV9VkBROc99lzTyqsVuXQN/4xQ602QYrJmmLM5zDs0bil4gPk
5HOgQdEsCxs+W/whaHbNmiRyO5MpK3EWYzSmW5TAZfCRnJNjdNpbUSHCCc6E0bWe
IPC0m44iVyX2J+N4VE2R2ALB5FLZebRqVftzNoypxsLbFBxnEpOCh2sP/loYYU7e
DKbeJ23IVvf7SLzGKZkZ44k1YWaw83hCs1VSey+2KpnsYxUO3Vf7WryEJ0x5pZNo
S6SDVSQDMQUT+0/fhbL2jLF+gJW3Iu4RMGqsbQ6AcX2MesL8ZgvmsdeVbKcysSmr
XRtp2RZS2FSlWQGFr4MfAe4c6TWQUyYe3TJolU0j7ZPcZ9A7YsMxn7jx1+7/q8e4
aXmSrOipzr94L9aVri0Z5cyEh1dXEd6nghGHEH2cc4yUYyiOp+eiMiYfxH/60IcP
WFQvUNXa5cGUxMtEYrHwtBHDnaPMZMfDpvoS34TNQQnVWhU8gqoo2E/06Qv+RUWT
C+B8EL48kLFkyhYwJAi3FoX9DA7lsEkYbZAHSiccG3B7v5581b7K5bIwN3J15ZY2
coryYcBXPRMsdIkkB4YFlWmdpzolYxlL4KLNLcMNRUUsdmD3ANF5sJealDIJha0O
BD3sJstXnZf8dMc5zUh0MnHn1+VUXOsII+uEAcpQ+zKfz5JiStDEJqA9K5nm21sZ
sFJraHA0Ap9pYPlROXCzrFWL8UlwnVf88qfAZym340ptcgW+0//2K1gNH4TzGK77
qFy8/aQr24alSSn08sjWCOo3mtQi65Tz5X3MQERS+uuCbL9HOI2SfSqUk/mnYIou
8tqFkpor3sO2GuPN9mx4g220wZnThhhJoFYKUxbDdhZVzszI/CrEJjDfEL324hfO
kkIZd4p2weQHHy9ZTK3AU1TZPxgd3WTjDOxepU644h4Dum5lW/4xBUN9bOIK55Op
YGl6BPmfeqHmO+wUDohtyVeftJ/Hj9AapoYhc3oj0OD5nqgKTBIvhtrH8tHRygca
Kp7dTM2UciYDUVmOMSeUOn8kNPM2MuOvF4PcFyThI1xKNnjvBx0mp0Dbpz2OdFwi
Q4BT5OFymFhi78uoi2p/Ug8rQpuftnaYv6lRKThuki/6MssWxvYHhTLpvltEF9Uf
F+7ZPcC1BxtgNwGsA6cMQNR4+wUNB0zSS5ErEYSfn4pKnEL/hgOIM1QdvN5UXAUK
ptPLYRSKGrRkHyfwi5Q+Kq4AxkAnlQbjQZAmP36LdbakfzFTxM7fJ305BBFNAqTB
dOcAs/OVUbW3RXV2z2H73CHs5tLu/zgvVwTnrzl1HN7bHmmdTGmzG8aZ5NchNKC6
g8aTV0dEVF5VN+AGwFa4U/2W65eDA8g+tD85P422XouDbaqT7HDYA5hnmkWRvQtM
fQKhaZ3KkTiDk6jxKXl1wFGPWtUJAfsgZyi+NambLaGKbiB6E6WTwiou5uBcLvl3
cKow9VXyziBNc6/E/QWph2FrfPExa1G/muqly+z4c6jzWDVxwb9cVULLfj3a2u1M
G2kHSPSl9pa0qJRDyPXIan3Y7oruMfjrbMojAFLcQie98QvceyhAiuEJpojaagOJ
U0RzQvrdFLTzfekEJjX0E42MqSOq7HSwe198wM1r6UDTcL483e1lOCiSyb/s7Ww2
qogj81vdr77HnUJySRoTsIssrBLjcRoCb8RJLyuLutCxJ8QutUbfrmf+Jj4sO7Uv
v0qi3Hfi5xO3Zub+oIIsgdK2gpSZYVMVefydFD/FmfHUQLuui5N8HpNN01DUAYNx
IhoOwrxz2P2RuD+qZ6pRbNrC2m4QgOE4rkaTNl5nsJyOqsmdTiVyS1nZdUiLyAsA
x+RRxgHTdkjULCDFOQ3cFi0utCqb6H4S+mhfWWhs6M5frF8czwboppCJXvpiopLP
tWYyzP9BFAGo9SfNC2bYroqXlqJ0f1C5n8UWQGk3+iepeWnQqv38UZYdz2MNljJf
Lgqkhp6nyyTR8aEQg122cdIEsfJBFkQ8DlW3nc77X6Rw9EezoCeR6YrmrDPgfZ1N
pd7rk5OA/2vtzNedTm55IhERBQ3hU+AHnU1vK/qrqFn8Noek985dpN82GoPyCXUL
MjNu4VxK1a7DmzmI++bkeeR+HegbZyWcJYYnjHCePANKuoEAUYISd6I2jP1LyA82
fVkZIuFDqztwOKXdg28nuqD5qiiFVTmCCPQbgMKY2TKNIPu8FjLMEnIAEbe3cNBm
LJLQqTj8qimy8thnTSh55jXbyFC+44ZrPBv62oFYk6I70wEEiKqk23mFN8EtoUa3
vdC5rMo60vDfUXOg+l5c1MDFN2/Zrnx82qCBZIsDeaBGmVqx5pn35IQeW6KmToiy
OqlBO/Xz74OiXxfiJH2EsLXdmhnDHkxlNbgHVrflMRUN+DnoVaChdvnq6zhw0bjV
2pkuGzoDCM93TR+ZTgATzgD+qvQjRiLRuj45Qr4b7p2pTGzx7e2s8nu5kbukE2EM
BivxlPzzjkZCkSVquKJFDxblg964uFqsZNXsBKDTaHnD2Aq3dlI9GlfmgTBc7xVg
2l43ffWBAAR6Z3qb6n33QKLoQ0dZDISg77lMMDF0qxPTYZddOrzFJU5ynmgF/mcC
jAsXU2nrpi/WdBhy1flpREroR7Fl1QxUXVU4ng5OK+MIkVx0AUHHVsyQ2Vjjo5c3
YUjw2lf0DfS0x/sgAv9Wg25g0mgscwtqDIcIeLKkN1a1F4yLGQe1RgIdXOc8S+cY
Sif+rhsP/zvmRDlC8rVG4UK4T7AxG2VhNAs5F5F6tTXEzPvkc0tEhJxqVbrBGa59
9G525DN4bBn1qOOHQhOD/5xMa5unks0U9uCgTbEPlXR02qDfwyTgcoqf1nKRH+ul
3HmKoqppAxj0XzAHORUmDmhfbi+ctrTyqskjo3l2y8Uv6kpJGkNQA2oX/3WOdA2d
TVF7pteiH+ZHO41XS7RJrJx56aV5cPi3qgIcUhdhZF+n7VMPRpdj5Hj5njMUUBp7
wD1x7tyouHjoDsqHkKf5scawLRqVTPrigzrscoHHhfWlokNA677nosGPhw2kXcJm
hfZxs0W0xhHKkQoGZtgnrwkit/ExdGAfuVREyc6yRuyBE8f4CMvimBM09ykfMiWF
skZn0y4qxbyJzRpLSYRiXhSwQCvc/u1tN2B9PmIx46Tf7dU/nTHMHOaGM7wEryPZ
rzlqC+axUQhh5b2ns0trXDaDzFxRTobst5QBpGKrLNYy9WXj1ajhvUhokAU3ncYr
qwDpa9S+7vCA3q19yV6VlXsWoL30Yc+IKXrRThFi+z/HHNeWiBPDIks0l2YbieUv
/F4viV3EY7rBzKOp5JpwSFkO+IG5x2r3WFc6Mg5eejpl8by3oO3UV4Hxj5bBqig6
u1bu8YaGcfHRnd98ZgZcd8kGXOqw+QOPiTQw+aXCRgpQUoMASTUSVRv7t0h9O82G
BV3JIP9tMI0x6tc99dtG4bZ1jaROJ4pNloSxVoPni+8ILCfZ1hZ/nshJoVa9Q8KU
e62brp11DNKfKV1DmLFEkwrMfhk9OkCONnx2v60fQiVAfc4dLIAtBWTvlNN0ypPB
3H2o+KdtDjmXmibkAj/ty3GLCZv3/q8vKx+8gy4gK1K5Xg6WRb19H5bRchpFMZUZ
8tYVdNfZc1cg4/kS2TgT7sD3GBnAjMiWXB7WX9MaWx7IG2imO0FM9T3xYNQt2Vbw
V0/jABK/+Hn7PGewLQu3yb6avBSDvbBFa+TH6PxYcSI5KVZacL85lC2PMySJKibI
7ebUByyoN0haWN5J0Szl95bC7dhFtkIKXgYFld6oTCgbgYwhkcQuFWNp25nx8wP0
0q2kSbXvSgT8p4XiyvFR1bBssMKJCjGKWVF2jU1tKXk8SHaspw2orhDHJ/Wa+OQc
tw88oTstbNG1peq9CD50oGTuBQVmwnaY5qC6UVA2lrHc0jHCQkoloIjGWXZHMMVl
Sl+RoQejnPiWR7C/EA9WwHe4I/bwtFUQxwWK3uC+KogeMA2bBc9PF2fxBVyE8Czb
+WZO1kAjUKgUm/U+OEFnn33uan5YnZEYxWPadNzHpXhzKekVXxk0n0eiHm7anWlB
y2JpUYpKXNXoEQzk/uhMyKoQWXYRM4tmZCOiULSiDWOr9i18iw+nZflN2lUfQAyZ
GPAcdYspMtzVborzsL6wpQ8dRSpXsDiqe6ixKmiIosApve7kz0JC69fNx8JmWKcR
1k0evV7gq2dv6GcHMwiZsolwOUQ8CnkIMb3ZYklLMJhEQZfRHiPFwx0b9gQmZYhl
T9f6EPbZ+zzyyQk3j1WOr6+/Y0X5qDeOKjGU1UIKYobINo3QW7lCnJunZr9Hq6Ne
XWUSpvDEqyD8RjbhQoDIBLX6hP8Or0QDjNlB47H7odWvQa38A5E/hF0XruQOldDO
5F2+Xy8uynTt00wrJg7QF/mamIV2nTHGYtrha9mud0ZMpYStN8AenuvUAJHNCU0q
TTClyExTILpWzUF3YfY/GtUh22HodxlHGsYiKCRWQY0XRewCALeEv067xML8rp//
V2U8tL1nZilDwGwLy/+XHAe9ZLU7OB73LQf/3XeSHjhlCytbijOJQSml5O3juCMh
3qdRKjOC+v3KUfW59t7Qw+kisZrnGl+Nk/M+Q9zleskM3elnd1Va2bXSV9rItnBL
6Gh5ibe4JPWMramVZzTUrZ3rJKsgtIlkeNXJ4EOb4Nm9vA1/ancmtyQcPeZE1cnu
dyKyA7qBTOz+h+NrnDweY4GD9gJtgcrJo86MrS+YSId4mc+xpXyDOI5oE6Ng0Ccj
AQTMYiqMhmQWg1VbTkhUlu+qArw5oQ0py906MBDj5C0TU81BXlFPIRyCg4JahJRK
0iiRKwGIt5iE8di7SaZzqH6zVGvvOJfUVlX6lIC8Lco7WvBOSydAeOczhB2qqZPw
yPHreVWaMxzIxTeDON1ZZVwaAqS2uBCyqheDhbl5K5nw7wpVaW+itlSgm4CMX+C6
NGpLHWRsKGY1BNrlUsMr3/lB9Vx/lZX9zm7GWvU9sRZshg4+6YLHFqe363U2WBKM
RO+0PqfyG59BFYQhNlCZG+lPoI80uufkBarf/mQJWVJbydd3Ov6m9/3d+SwFI6DK
zq5GXlqyLi5fsvtN1puY14dB8OQ5ACmS/F9PEufIWZGJqBIVvtU/HmSXJ4s9YIaL
AbR/Qrte+BF1JcqtURWci1CFlhBuMhjFBslHtes/FzZ9i/PwBOqvARRp0B+IVKmI
BoaSdGNs6r7nYSWOyWVBAgaeAncEEok4NvSsc0pNlYlKKmkxlzXuXRLdg2jK+lqM
awI0MK0ZIHeqTlwq58c9d8V6+ESWB2N3lcfLKWc1G/kvtsziK4NS5ZGX0RP161MR
G7dTyu3dTFzahCwtsT6IRHt78X75afdxKutWP9tFAi2RjgXlcYuhR63c69zSYan+
lm9CrxjPyLltxXwYUCOqXLeDdBliFlQv8KwisgTTza47QuA6D8thcYT4x0tX0MQR
6LKegJ1opuE0lLxDnPmC8Bgyuf+B9NP+x3x+F7ZRnzSWCjMJwGxgFKE+ft4Fkrev
8Q6qn3XrfMVtrtmX2L4Hr8rh/u43nT4J/EOyaPmU53eNvi4PV3tzM0H3BQ8TkMHu
LJ303dlI2lF6xOgoEK/Pi4xDm3PkRu2P5ru6/e86a5SqC3Uz1XKX9cj4G9Idfsxu
bqUqRY4t3gDz35Rko7n+DGxdTvUz4sLV2Pcfmtbdpp9MNjrS7BC27cZvh82mLEr2
rcx4vA4m0xRADCO86jH+8folnk2OeWo6ubb65dZlWs24LX22LkI2U+AgNxAiTWGM
Zt9x7uRFJ3B2HsH5jma8if8pqN5OUBbShaWtTDPNSJrrmfXIqdsyhht0BxMu4n5I
cpbIbkyGx9O5osFlyasekvLiPaHaeQjYybgFhNNTtW433FAyhR3TwYTZukDQlN2L
r+2nQ1DOFQNTFNUxV1IVw2FtowI5mwxIqykcS2zixAcby5MQ8cd++OlZBP7WDA1q
XcmppeaqKlzPW+g0C1MhyERM6prH+vIrwtOrdO77BNtwBtg6VQxUOij01JHJylIz
oHLYaQrKLCTlRS4TjILZIPb1MT36fraiE2b4yceA16e4GND/5bx8fF9tC3BiLbbX
J8kvYtIQiLE7cyA74Z4gN32URnTlfy16WPgWhDRg7RvSj56lAP9CEYvzyBeFSjd2
JTeIRLG3Rk0wMMFJULKqoUx3pVa/mq2j5Hvg5aDVAkTmPkE//SYhFm0NutMQOzPm
b7hOwM7YfJ+PtInrEDnCKBYdTAJdqu1sBM9lJKyyENgtvSdJ53fXouqtRgoZPQnv
6C9ixO6cn3TUEbEq3m20+EzCmZmD8gJm9+bMiw2hi35/c8aigDavwg/1g8ewR9gd
zEKzWY4WD9Xpf4oM8Z4ohVjlfkE2pqnvVF+5iFp/zJu/+UlyC2V1sEzZ6BuXgP+E
YGY0cGlY8vrS0R2D33p46eq8xo65KBORR8ARXlJC75e0eqfUXuDCmAc3Rff3Jgiq
zNuvrGlaHrL9NuywgV3VrF/B15JXClpK25cq76Qez82p3zgCZ5an4GmDLBIo7mlD
AQhaeqTAsuz1/VKJJSC5gkxpeXNG94oMphqXgr5fZHbtwSSBa8F7XRus5+8EBvkh
MaystKy5ExZbmLLzoT3+gIGbI80I9Tv7xxE9O94qtLuS8aZQ6Rqrjjh68GMFIpKr
PvcMNHcp63Bf6nyg8w3ZjZdc4MQFLv0gBgyY45UOVVgVtDLuMEjppUjO/CkIoJ4J
Iz2wnEIvQVGZPd6r/5EeA2genBaO3lPByyxItCCnuY9hJOSb0BuRazHkgnAnd0rL
jVP1v6t6YKBjKEOGL/jf4cr62QJ0vgNRlsp7sTJMMLR7ox2vX9BYGpn5T3mGWTBD
A1VtvgSmZ9gpZoLKPkeQIoSU+W3DqLYF5PLunYxI3RR6Y6OD9NrZ1r2plgi785bz
He+dVB/Urdf+m1JQcj2JuyhJJJgD16EANQLhGsqwp7yYeBiBRsB5BpDYqXu84k/C
yMBt2CvVDJU5EaxEhp0i8bpbCrHfKU6/oIttUYSZrmijl7cWTOeQpV79IFUDEnYt
BuPPoby8/3dyx9Q/KTYPAmLYcQL4SCW4TtFyI8JGTmbZda0UQ5+IOIBapa1zZacE
oob2+V+BkTjl79Qme7BZBD0L1xubBLCLTDimbaww/Af4tnQRRbtOda0rHlYWj+IE
DxsAqIHauKCRODEUcaqKd48PdWJSZ9oABC64oDKkvJP/+/hSz4Geb4kWVpHIR+Ok
/RU0Vc604t3o7qa8KlstB5T4Ax25wCcG4Ew2A0be2qZ4Dapu6n3xk1E5B6+Tii9p
we149qBEdcS7lWTDQAkHws9LKgXv6M8dKZb7vkJOgV8APzvyLW/Zi8ZPaIgoNE8p
Y3+JZxgg9Qne7PF/jRaOeBv+66Aar6Tsc4HNGccfkZQTHHB80vmRfGWoTj9l70Cb
5PWCCjrRO//HZkwBdHXqY+FRgKPvB35s400foHoDtP0/3kFPMH743T2PPbRvjpvG
oAQsm/peoq9cyPU81Gp4oFbHX/0GhRiDJJ20uTYGNWG970UrxrtHEky6LRz8YNUs
zOVWBn7aYi9KJMzgwpF+5x7ycQIE857VZ/cB/nTLmsOkG2AWG18nj2YYQWSUGZVY
oVWyjEZUb91CroQztP95YBwevMiBoEHsYdkLj1DGxIheaC26tVecRkQmswIPFcY2
IU0H9k87XL+Zyj7zFY1wjbAmfRhcweh35fJeSgvUfBhf4qcrstU0p50OersUtd0/
FFoI1uo23XTRNA58TrZ0AxTr8Uyjz84+sQdqvE0jYz/yq4Bj9rj1hxlZPtper/uD
csHGvU+RHNxeH62YRtzWuzSCN6ID/NAH+4qNMZJj8c9+5fQTG6RYxiLbKK2X/rLi
awSXMgzPW845YpX2otpEQIIJ8O9ZCjXkEyszWW+Jh8GGqmpk3ObikB+WDaOAVLfi
ndj5xhWRxgmONrJpecFzZJQZ67LWYdGmFgEDb9L9fq4VNxAGUqwhGUhnt6/2eedY
K5ElqYgI8BT7DdbHcDlwGw/VWaAmLPTLETa86e4x/l26kfIQrOA33oocP3Avy4fZ
NlW1i/arnJsdcKU1RhAmPN08uY446KCA2j+R6ATWaVmsROYPo1q7BngsjTeJ1My4
t7CjTxxNzQTdoPlAce1nPrQaR5FI6+iutP1m8iOenIBzqVBXhNGynXUiW9BOSF1a
q0i5S2yjdD/umW5+dQouNTWdKBaWEmbOz3qURNlJE+dL7MUO9TUcygmQXf7CLtpX
dRQ1FwKo8I+XTr7t3dXxkbasUkeip06uFsmoyLgfanzvrmZ7ranuYPeSY3AouxB9
h5jO3J4HF9PreLs+QlFK8TG4DZODgBz2V0XQx3ekvWQwE65gQNZQiMHcg2K2chRk
OnBqYvl+BowtZSZrl/OPrmV2FJT92B232Yygjm9w9EXKpby0Dip9gOtWrCsqfzAG
F2cBGYn4uxW1LXXDIMbliF17IHMgys7nS7mrgChwlQaIuCJch29j174FlY36bedT
taCNzpjNKjTyLWvHJzpOBoCh/FqtDqHEyTFnKR9kOn49wGozQJT+wS2vphJFHMwa
5ool1nqLUCuhE7dcNkq5n5MpPM0F/ypz4Ja4gLjmAu9BnvKq6qmtc8yXhnSQaeiV
8Nugx78oFL0t1zt9iQS688c569TUUfBzeREXO6sSzgRjkM3SBZga8CdxUmY6Wx8L
OKUQaHunEXrBb3/T2odGO7Ew1VeDoJAFmssp5SGeD7uDJjm196zjPogOO7c1t4Ro
YP2+e5AnIHb/BI9oTBFT5BFhQx4Xiza0Q03Afg+mdfPJra+HxxBY0rxh2Mq6dvb5
ktbgWHKBrmedFhTpCq0VFVr04j8rjl1FxPFb3DUW039VGCBv1KXbYCh0bffOO7hB
PUS1q+6UCWxQ0tOfV07I/qGPdHQiOAqud2tOhHIS0pM8NQwFGAlNqojw3xyKZET4
2hzxxG3cie7l7Q4TJs2AjhPxdFRzv1zbUE+0K0FK6XmSsilgSa2DtrxVSFT1nFZq
NdJ54R5uohj4317LZ92ykL0UFSNwATyi9Hby7HX6QuMFu9XAq0dSXWOk9yFjpcOp
c9522IAyXkt//GQoDCZak41dqBhW1IIL8Zd0Z1tcvdGl2hG/Hyx7FEtzD+lMmzdQ
FuOloVSzdkIaNmwPyTw2ikOh7FFULrDNLLBXM64zzhjdF5O3GSpzpKlnNUy61ZLz
z0Cx+JIJ6qlooRwIIiDXzUI7gN6keq0yZpxuEQpXzskzs7h90ZsJSIElO1/k9ICA
gPke8Mz4mhf1UVtMpnRxeIv5Z2UA36Egj2Ac+TITSYjkmgG2mT+Myq2O019tUN58
iWnl2jsCzvLKNYLuwsXrnS1Fvo0P1/gv7LiOdb8s4davSORJBjkjRmXJ8PR3FUNK
cEpqSjxW9MImVYKtz5rLKIBPlKdz4t0vtpACTWJYdOwHlQ/+xp2K+2G1QKAWPrN5
uLRd/Juk1kaWZCxIdjFXR2YUVYesm5Ust4Ge7YT4WQ78InAnMr+UFGdqiGXEdq21
cjnlEYJ25jajYekRziwSHj4alqzgN3Y1+UejdGbtcV7Pf6BMQ+P50sI5l/nXBER/
wo6qzPX++Rgg18tmXbiUaNyFhC5Xt8rjbL9MObvZ6eMqSwJGV5uaz+fsjFUX3Fp2
89AQD4Po88B6u9mIENowG4I6XarTC+Xrdgr4WviPKqUwUqUNFh+ibMqEJoxDmmIT
lECrJ11Vk4eqUAnAstfKjWbfXVBkHveUnuI6L2WM8ELPbBtFEVTzTDxb5KKqKmYE
OeT4WP0asmEPYehC8SWTfMDZQ9o53IJJP84KCAfvSUfZUpbgP4kPaNE4TL8pspUx
mY4xoikCP3qIMXSN1VFzKYIQmj+xGsSI6CwxrQ6Ci8lo5ibUOQ637cv4wL//k/R7
8Z+TqsXGkVjkC80BbNc7rsMG8fH+y/sBUMUkrAhCXZY0NEvB8hblJC24p8wO7lr+
Aw/ty8NjxZJyY1cHuxVxDwMyJtr3WeJvsyq7qLGZ8hwPSM2LFOhPFSwNfLS9S5Y/
997kKuMg96J90zAJMLlOYAlN3YMEggyTh9blfep4S3VoYo6gu4gLvmkYy5EawC6A
ceGiUW/2hfdKtdIBaM0+ZE/GOmXeNHdAWdiVQioWMVebxWKUwHMtv3KTNe/Dixkr
Nn5Z4/rN6DsDXv8HHkxVkliGUigDAyTmPvgY38x9pNBaGDz7+4Pta7/JjHcMdyhB
nO36EH+O9tnOElT/obDmHlQ76pRiTBob+9YwbU4o3g7rs+2HGTEWfletzCGOkwGs
v29tuoL7hwaGRMxWS5HTQCUEROx0rCray113fzrkBBFtt/i5uX7nj9H6AAKblaf0
49OXYbzJJZxSf3TFfuhlhKP1w43JGELSxwSNZnoASH5dBWktZqjTGGNDi1Ibo3iH
gOgCmHkQfkpWgJy8EyFsTrluC5Is9lhT8++jJuzN/4vgx2YvMFgDDZWhkSoLFDeC
dvO1QdTUxuj9cUbZJWUqqMmnnM67Y77lvrsS4A+NvR3KdM+5GxUXqFTVkxNgdST/
HfyvZKFlDXjRsexH6iJRV/JLAWQbx1Ug5MxYfO8MCvKchWNetFbfEGy7ZMiwOMIE
PR/j2xvt6tef7ZrqtKiV+rVroAyldkWkmI/bfpKlQfi0NXnQEgjolfBfvf1S4H95
MLJSn4HxQvRkVklIpBoJPtnhmSyrYh6KxiqBtthdqQrpkzai4TwSTVtqN4LkQ02t
zoBvapfAyHegSKTZK2G5/0svKtQMlO+wnjMKP4+7hDMwNbXXg3Llg2YDMsHUal59
XKiLOP8i862zBepIUuIsljx7WuhaSzEDDAObAHtUyTcDzl0IbBkNC6BKeb4/nwvi
vTSXCeMn8ZD8xXctnzdMReQBNCGhB/vxonhUe6BMx97PtnCrROlSuVc8wUCLKJQL
9BhHom4n9Fhpu2Nkr2DjO4h4kVUJyMhE83LOfOJ1+rGSGwekqenQqw8Gjd69g7sY
LMkzT/NvSM2HRuRfBEtu3+VNrIGmoHt0QM2kVmZeG6aKJvdTtUeQOaigtkXqb6R3
sOTwVyiW7+DlqxNJ7J6/n4vNAXeKoBAGDGz26A27YqQQjUPodm52JSrd6Xh0EHku
KMlfT/tqRlRvOtQB7aMaXw68IMVtx0kQxF4XC1k4W9jw3bzqKwcd7OD9YbDbTsLm
pDz8/BD0ib+Ul4e+d9vV8YgDlnEPX1+QqymUW9y3tmsdnrx7vOWbrGRoubnKElku
ehmgr68heWE1N0hYo4BiVBClwdiw2nJb/GYGEGLjSFYZ7qdeOAwrqYiS+O/xs+Uo
xhNu+Fa3peOKDjHSravASELwnvzuDtjfQKXBvu0NBTf0xUtCrbRPnlCYOCGQWjgb
dD5qsjJKQ+5VtO6889GKv9cMSD47g9+qSruXgjuAcR5+QyTFWQh99f8su0Pqck7M
qSZHLJ/9EVKZGDtGn5Piw8HrmoGJkp8OzDZTdskQM02DASxnDtNQtTHvpuh5Vwpe
ewpR0QPV2ErSJL/A+4KLyt33nzBMlnNvklEr2GlnTSQu30rEVCrC7g1C40Q9z7sY
hSM8cWeHnXuI+JvG20EdYotfLWN7f0U5z2PgZwwvZnt0yEazzIbAiy+3sZqMSSMV
Uw29OSXGwwTyB4SiS8mmnLxxjZp+EPeMC4nM4BEzUrw47smU5OiVyKN5pD1Vd6yZ
QRCe3e8pRx36WjvjvuP3zMYBDQSmuNyb/CPphjYXzmpkoVEjFbcJnwaBUAVHObOk
04B2K1D/y3w/AoLus7WLhzI6xSUc1YlDxdCfB6L4dDqm5YDNHGjEpJYLb0LdoENa
xmsXY4A21Mj9PwjDmv3eq8kn4vWKACqLth5+ALZtBZMSlhNa6zzflbFAALVuwTzf
mIkSq4VjXN5t5Yk/GbBpdoMOZrTJ9ansPPHEJuBtOnr41ah9P2ZTCTVrMhCUjpNx
NS72QsGRtY6Gh/o41aspTEpHGiQfMIjK0DCtBowH0ZKOIB9ZjGVd26rxZZnIZbVA
JBRg8vTNqGC6Bvu9qSQrqiZwdlSBifmYUHxu1Jbg6guDJ3BUXONKU0j1ad6ioZe2
cyEQ6Z3ny6VDsd9RDcCyoXsBUpg4QqvbJax+eapf3Bh3+KjTopijDjnL6NwYGsmR
C7CAGKd55N+BY/MWjkr08mda2aYZeZQkcxYWMXLFQyaLFneOpB2MpRJk+i6V+BKx
HBKmJmoiCiu0CX2LxsRqRAuLXzbH7Na64b2GtFuyOisjZPY1mLCIKSxxG8kV7R0f
zayIxS7BNawbfeDqT2fL/5ERlOBx0ysVjNWkkh/dg/tKwTfg12xcNN3nW2HsQAu9
eLjEtk4/US1dmhVrs4OXsgSZ8ljEqOeLvH32Z9fytA1ojYU/1r+pL7a9cB/e4RRJ
h7xusBJ56o7hmf/4H9p3LYnr8SfT70eFrsRGkTEoRJEs/dVsFuXCXHraaLdmRutY
Wyf/nBXO+42xNDGz71OY72zQuTrestWHD7pTKXcUwGPLz+OjIVHmoz0y7BEcsAoK
W4/ku3pMwLvr4WPxzKYT3UPD07hbz4bMeDVoF3hvf5DlD2Gj5aBuZVRS6ziWDi3Y
vCU/TzZxFGvFvusoXmKS2zSLJ+ZlqpMuqfwYBWnqN8LGjSJJtLed4RRHMoKEtNMj
aAfUhZITz1a1Qwu+AqJL32SxHZnUBUkkLL685lsT362pWp7DfAbLw5lmKFtl7PuD
0odQoJ5euLxLlvND4kfN/8N1FqjWepeAPxq7Ji2jcme0p3cxdLrT2HZEMZu3E0hV
hHXBcbxUGw8Vv71j0pwK9BSPUE9csOwUdkaqRBgbFyIatBceNK/8PVgliJnzxq6i
ZG9nDjod17bT08LU7j45CTb1KYv2IVUcLj6TwPrxHpZgmRn7B8FoH5UxYWmHEbjV
r+VOfAn9v8ZiHvtqQvKRyxItNvvh7duKaWblH/iJBbyp/QDLqGb8CejpBPGLNplf
hpf0307XR2JHSRRYCigBmsLOVwdA5PLNI5po+rCFSM9LEwVH2LfFW/+ek1Vk661p
ViFK8b6RVrFh6NjARrMMG5jL9KSPfjF5iCHeP56mNUSbOIl1ivkOZLzw4vkUtL+/
CbEBvLsdxxql59OqqXod+eVXNUuZUhlq08hutDbLTg2BE/hZ+o7SS0tFs7t7mBmY
962TPnSXBuQQVBBA6A4C1rFSGU8iXaPPNCZgDXpKFP6TVs63SfJ2C5TqDtrwAKyp
X1gmKBgLuYZki+NPp4y1YpZKY2ATWCD0yUDItj7YC/mByqTT0u+sWLffLzxllTFa
8uyGBQL5WzQMlsSOMPYI8zUtXL4OvukTGgESHJ0zvJt2kkuJXXGytGGxbZp9FIeD
1Ci9alGnmjtqsslFRzsDW23tPo5L7n+WLAqMXjvTcChLIvXYVFZBPHCLnXcVSUfe
r7g+LgtPPZ08wdTNSXAwl0uwY7VFPOugfk/mKOt/j1pwXf3e87YrSXsvAWn9KLlE
pHmoUlVd3E3XOgq2IshQ+1SPaa6mlLk2gF867Pia4x1AJlH8LHeBS7mMF8l3Mwee
O0qVnAI1Vs27MrB0wv1Ngrf2dN5f6Cyav9db9J9F43DetPsgLG/V5+30cnXd8pqS
KqRol9bG3ZHsHKPprGMD5gYzeJ5/2yxzwgW7TcyqZgUDuJ2AQkGxG4Aihbd4mpvQ
/iHQMJ9nlMS1GfV0JaVqZtFsMk4BzBJaDXf0LEZ/K1VPCEBYs5a8y83yJr3tseC6
mqGADTlEIIcYl7P5rXqluDO9Wf/nFAG2N+iHyNsv/Ziq1HWHY/zghBDuuur+aT1B
8h+px/zWjGSvIL8R2e5CP/R3G/XrNd6jeMKF9NZ3Z6MB82fPoEv1+7nu7Dur6dHM
9/Q/tdL/TwYEFo1Lu131FJ4Vchgfur1+t3NX3OwLZKo0gO1ynBkhZRe2Pn+sMQeM
M5gawv8FHQ2oiW8wc6YGfiHdmXQB0b1AmEfuQzJl2Q/5XP42RnIrZr/m61gjlX3Z
dlzobUzVH0VuYRsV3aLbrHxWYvedqgHeXOyy6kfBwQ/02D81x8jZBgrIYMOeoIaZ
UHzqtP7CIqFYYhaeCt1vGkbdISORjwWBR5Va1H/yWmUW7GG7dMvX65W0di1/ksgx
1TrIkCtk9mV3iatFbHonfeg+j6zvUG3ik85TZh++Epd8CXo5ISfiuMjwmyACYned
Bv4W+tMA8TzOvEc8I2nZEOQXvW7xkmA/MS49Sl6qCSvRS68JNlGQ2u45E574C0cB
mvhOLPgt31Md/BfYX1kHo4RJP1tPymFeYz1bbiK01RgQSIZIP0gav43U4d4igW8w
vp90ueigyTUyhj/RSBeJvSP3K4bEOUpJ9rUcvA78IswSfFbMCyZN/kgMWMImy5hx
QblqziIQIeK6YMKNUGZYbTYFMlbmBaG67kc8GLaIkr9HluVKHuzwoNOENdXO/mc6
/NHUU5xw3VZYOw6ZzufsP4GTiXYjxsn3lkx9WQfMWS1f8V+L1xizGF2wReEen2YU
iDgBlhehJ5a8bnxY9Ecw+YmhBYmPnuPzFagAd5wxb8kSxizla/RfDIlcW+ukl1wU
VbwNVSjUCu7Mk0yxXI8j384dO68sHQBq/RFyEkXQgQPTwj7cDZT8tMvomQLLNGQN
zlrKt3EfsSO95L6TmelusNz67vHA29nMYXrUX+gWoLhK13QC9+fkOjVyNHCfcfeS
SowQ5Rs9UdHwwW/qlhUroUMT2k/vieTJR++KVD1lYzISPBpxGsCP8UooneWTc9cv
QT2Pw66FwDy1jpADSDlKGORisjFteoDzm/1CkftauQOxqptKsKpL136vZtxeX4EH
J1rO5tJtjP8oSx9o95kFTloQlrDsDRm4ubUwXUhrNPesi5wLqPbQwfIDNTwD0kpS
zHc5Ntt8bH90tiBAoxAQiYB9P4wOc7vkrceAgkN81i/duHAtdX1p9zEe+1AGLjNs
vxL9EI2fAwPYl1x2LCDA/rDTOK4djP2EqE9aEyKBMmlBbZbPhL2/V/xGrq891NBF
gUMLz0qvdeMvZV4x6ukbBnIth31j+fUUDYDa82/8LA9W30WAGmFK4f1bT+G0yZAk
W+rRLIXuumWAsWywi/TLjtr1fhVTlj5xY1JCpiGHGO+RT428qqf4AxqKIo6Z00lh
51dLU1/Rf1Rhv3kPyTSKHn+8Sg1RDixPmMLWN4R/mHfbUeomG8Zc5jpPUTBnI2Ht
ouxJWWkpSR0lQg7p9IyaPSVZg39ndcjKme77hnwpAy5XrklzgjJ9lKSvrQDflHrM
CWS8in69ymjKCnBdOTOfaeGodHp7Jtzn7p76A9uYXqdrhY5ALhOkfMD++w4r6re6
d3hrr3ymRdFwb48YsU7KTATmilGHw/Vhz5dSuK3YQH99Pp35+63S6qkyFW9wBRIm
0pZqMVHVRzotBCi7UGAB4dQM3hfl2/ABt6VSyFhDI/r+uycpPCupcfJPMqMULT81
Bw9NbrBPIA53w1Au4BmU6NAHnz4glVSYNpJO/Aur4wgD/jIcNhjCeffHz9cFxwkp
QMdZ7BdEPoD3HORNANHOXCxBs0VrwcBvTGIB5CKLUrb97kBGThVlicH6LQzQiOuI
2TH0hiWbhf2whHtH8rJVAzT6E5jCtSQlF9zRUV5dTx16bqd5CxEXnimqXbzdhn6C
IrbjLBqFkIv03VWl55E0M9KdmIL/SKu3p+Rcu8Mezl5vr5vUYv/leAHBZ83yf0z2
+QLnLIj9ZwpNgFP8eRq5WnJ8xfwsQGlAy5Yo2riJXCzxZQncDzxqrpoSblKyr4Uc
j7D7U9V81TkunoF61JIU7MY1SGcV0mWT5fxSienPJ281MdtYiZlTthq4miqgZWKT
YWb/MnjTcWo/kxlzvPmOr3ynqIwnVTFak3Nq+q94e+cGj4hfLZHakXEXD7YvWd/A
SI/FS6wFT6M14KmCkXqNTxoQgrYMiALKhRJccyyxn8FHEmzUj+UHVfFiQ87umexN
v4z1ezI1kiOUxwpVA0WEe6eexJu1zxqq9VfKHKprIu7YG9wfUgTc13YNB41CfVtU
5W6bdvjlTg9rEubYye0cjcijZ42KUdgtqkCKLHDD0lx3NbEbM0eoNMsJ/7iUj7kX
AS04W7NKAjpbomCyGs4b1HwCmo+qG6dV9nDCSyF7ZtGtLSWV5WA7YJmvtRw6MoT8
2oU1yAdZzhyB84pbj0EBFY8gGfFLlEHUv+qNvnJyD6ztbwwKFKLQxibw3BFAQhG7
tmWMo3PeGCH7f4FuooExfAvDVZST8U7SurMkbPK4LHoGQjSJVpU9k+T+kzQeopuX
iEXjwK8GpowwcstmqO+iGyEP+qgk6AkUHhylUholxG/7HSZL4Y/sgjua6wLycyki
hsrB2wWrS7b3f9gCS2zcmh+TEyIZ6GtgdWGYso6oHxXzKPgT19NB4P7ct/Vez7WG
V8gyf4DxQUvSwREb51WVnw0o+fLvAacWT0hPeqMQ/VOooHdyfquAHzz+yXNV5185
ntsm0QoAcGELztxEs3GCyHiS3kR2OMogmNsQRtwubtCh5AGnMnI4Lh3/eG0odMZL
+BGOEbI/Nkibj12S95l3O4AqZ06HbcbHqpItzSVQH05+zioOTbItvLK0y+xvYpaM
uoolQG/Z1qcE5kaM56ybdGiIaziq910Ht+4RcV6BhhTy9hnN/nGKXE9b9CIacd68
4fY7AIkcZdA5AbaCI7odhoPaB1ZDlMwA+sUjN5RvvTeQaEY6GjJeb9i5ztvhqP+2
aOgmhQYwfqgEB3XBBPwwuxRxgq+KthFbGvtDM0BMpt0s2nTFst8sMnMs1qdKmTLx
eQJ611oahvEOdzMizOUfmUaMBMals2wV3v1tJDKhwfldIWUL5e0HT73DegOKJhdj
CyEFoTonIveZEHpx3UykDoU62890onEH3t5dKKAZDM2H482ljIynHar2dyRXAf1I
eBrRY60b4t0NFEcseYfMZqCncI3g2+nVR2wWJyXa+bNudpodZ/9XfTUvLLPEkbjo
coBh5bSC5wOXFTgaSGCUud0JifdPOxNbz5ixH01Ze9nZSYWuD0Jq6J2iwSAcqJeA
V7ksBgRSpCpCoThAFyJ8tG610dym9j+sQoUkPvvfP6yl/wX416al3ZnQdG6QwE0f
AWzjkJWqJocewnfLM6yTnrKZomIUq7lgeI8q7272/im3JMl4tII6sDRVqvmBEmx2
12aB6oS0QxBe5mFy7Yz4LB2m/ArL4Yih1fnoImsLO3M8DJovo8YXGxhI1VUL63L/
YpJpx5MYD0969IGNucr8wKna/ozcHAozuxsvhf1+brbeRAiQLEpPcBHbvo6aYT+6
pnFOHL0gui8u6ejp1akawcAVaDUJND3cUWQS5pi4jPaRforZoVBHKW9qzCsZ0/dO
9cLOaxsjHdf81SXs/1JQrZC5EKtY2VLlq7WcWwolobOxwL8/Zl/Q87FsK7GhLXm3
PuH+wdwOlURFGLrNhWi9IQDpsPoUalNmjHcCcLum4T/Ax1GNVRa7FNVbqgY56WPx
wFJ7nbnd2fPVx6KGTOZk1h77uyx66K1DdaSsAWK6/3e4PGcDE+qP14ujIxXCcvqe
2bhESs+os7uDOAy3jYDYvzPP6TTH9rhZjUPzXiy9cGTNfzCy3y5r9SWSf6l+WvIv
P6LajRn9lNVey/rhrgN/I3qJf17Rn05XZDVHnIEMyq7d/Qtkfpzt8XthDTi/4KrL
8bPuuyphM14xvNNYVdzSbWP3TOcR6oLCxzJ20QWD5q46srey1fOy3TadmdtLYcaI
go9+j5QX4XVzFKKaFGJxfz4R1yCsUsjNNy5IaPhJxQ8aDP1No9a/zhHp6QayGwYJ
CTAV0NjieVZhvVtPpJn3yLN5K//1wNB+vRhsvIa168tdEGDWFoVO75LZPi2Neokb
XrE6bzhLqCueg/1OS2axIpfb3R21mQnXLnOQwwZnAzbIiFTlZae1ncq+6o/78e9h
WhlGQF6Wmu3cz6jKS/P1yzDh593a4+ZvX0ZlmVa5CzHKXBJtZh9iGtWdI7WNW2w0
zGBKoL118zJlUSfCZaVxAMV7HYEGcmgHa6hIL1YjYUKjWH1CTJgUTs4j3RaFgoW9
pi0XdQRBQe4Dkc9qRsNy3ZZmWToUg9HU8CQXYf1fOW8qOwdRio+pShYmvO3uwGBV
WXdz9xhSR4LMJT+5QoyxoNGSDivS7TXjcXoq5vuDVQShEFf8rStetz480W930VWy
nSJCvn6O5Gv5T8RJMCVgngIB14DOSZiVYjlFXPMVnpTopoEtzr+8J6kcqexLelse
lgVMS0cmDFQoaPDa0Y02dolOosZ6QK/DC4AnSWO6QWlOAxfFkd4ULgLXgEzYTauy
kTG1+NeHAEEjBB0km6aEIgUifxRnsBhSgDIHl6NRoVIACd/RYpwwIxXZVmKOXyqK
Y5DL1PD6SLekLqQyrmVo/RfX5qKiWm0MIAAK83PPMLHEGvglnt996jW5KMiC5w0X
Lrh+tLH3jmkpdIyMy4EdAFvk/7URInn/kSc6WrPYfS/l8NO/MPZMzBs2LOdKbGjO
bXl7eE7ip2WhMA26Q0sVRutvgsIZV1ZEho+3tPuaVqbWEiuZZjd/bTl8Uw2ZBsKE
VKLN31m9DdIXmngVp3jemqBjBL+tuwfDA10mbKJeqmJdgEEZ+KovVhtEf5GeM4CG
Vj5bzItwQ+O2l0ZfOEbi7TUg4pG5CyhkDJc6EiPJKHuXyS2CpoI1bT2ShAzUnkWa
0p5x4HuSbh9jWnMgEfhoPyGcSEJwYuIdql+VYlhP0WC2nu19riCQJKP+M5qXCuQe
n/hGYxKj8k8UNlcYGEaPPLkuq2G+HaoiLYVqEVHokSbGRlXmgCDjd/vigpSsKDsM
YxIG3sxXOTQdATxr+xK3LzlRi17UoiBi4T6oKZctzEKZvLTwLX7FsD1CxW2ZJP7J
VWkpRNoz6P1jQxHZWB4D/FcG/BTi5ypTjWEbEcLt07SHV0ipGIo4uyfCxUVwcX5H
V9wRuMXfFfKaFy7TnRh21h8oS4yjKvjX9XXX3yAvmBPnHIqrRrBvQHADbXfQ3L9u
U/1W4kSkeAwle09IafFIrmcRFvOgQmkJ71s09DqplMwj5BNe8lIt0JLQisjn14mG
eUhTWbkew+2KK3yZWmttk/vZkpfZoQs0lOevhbTvQwv8dEQJD8eBsHa9TMuVJ+dJ
CvCeMbyAKTwcJrsZRR+9oUFhzNTJP0e3D3cxj8vFTVaNsj0CtOmIGBc4IMaaTyr5
+SVq0yhKwstWEW8hrvtDD0UvxL01Fz+JcYhvC77sJ8FzbJcc4Wri76oXqApuTGd4
engYWChijRjI8UlHMp8aQbgUIoUonueUnh+EU/5DhUFx2oGS+WucP8n8dOB/LQsB
gX+/39ztz74oNtiofvBhLJ/9O3GZJCFRkckVWjWcRghwmaoScNC67gWBL4g3ZTXK
aM58UwJfjKYE3l5PJSel4M/ZzKhKi+pLRZv1Lahr4qJ/IDPQYtv7z1AYWy3FLbGB
YPshO/UiuaC6rNoToeQ9ZarKhXbZ+FVzrjZ06fhTMR9NmE6l83sLUKAwD6M2ZTy+
8nVS1oLCSt3g88IevB1y4FtgW3hxyhek27Uqa7QQMKmGJNze4rZKfcGseeVzjDLn
86UN0DJlOOJYE12ybJPNvsDExblANdvKYGhTSpl0biOrZmhZGRmLOoFVh0N9nCzL
xSxgJzqBiJlzpNksDcbLR377bGmNC64dp54X/vsoF9Et3dXgpd1MuxrCRgi1HtTL
Z8F3WO/SjwxlXP+Z7+/aB8v8WnHYNQIitCX38Yc9humQzTClNByY6hNJpAm5CVnr
M+q7OjeaC+M2q6BBASTCXCP62O8qyS5T1VSl8TlC+LXvZUNYWhPIFCi941nmupor
3u/YGUey/mjQzou78TI7wHcRvirZrUAjkaIbmdKPyZpR10IPODtlQJ803kkjiVfP
doCYpdvdIi5BFn21ZhxKN23G55uZYbZ0oV6ZmwDG3cz9swwdY9CTVVkBiZ7Gyflr
DAzhFplNzmZd85Jqp/NZtDsi20PLIyoVLFn0vc5W1fQz1DPJ63b5NktcECEcFW6z
Eo3CY0XS94jQq9FwjSZSlu6YeHV/Xk3LrciNNdKh1fZWD0O/n+rkIlXuzd6zDRcH
v+8ObfrxeelLTle9zTu3iaY/QzPLJnCE2FV8A29pGkPgVat4kfCmIZr0wsrH076n
G5CuBGZTIuhr0RBSTJbid57CO4cV/DbjMpTHAxswHIOMaBCOdozEsoVmX5sLcDyo
PVkt87MvM5UQ32CQqiy5fePBxa71Ok9+PVxklqIXMFkJYCyDflhBFMeZRERbYAQv
dBil+36vkMJdhEPmbPcw7ONVrGhY87FexZ1y54iLQLeDYmH9FtWEdVvApamt0s8G
BLlhCUWcNndUfic5mCsCs3/8OCoxPjxCEIavekoT1YJPQr60bljBU5Cpj46bgbwQ
6Cz5LO2/dTNkFfma1o2ggo7xk1Rw0Ur63HCo6zs75HwkDfsEBNIdjT9hrzGmA0i4
EmFdYDABsNMnvrL04iACIVM3T+hz0XouWGGFpp8ckTR1km/NwogkG52Ke78GIz8g
Cq4X1cexq1YCbjUgRM1zr63lfwtX2mBILVm0SwrAWzW7EVcHAZsWOGOmT/aqaM9B
FMhNOMe0FSA6JML9rcToBtHd6/YH5R5ey3gHaQ9naAIC2Ub9BPM5Z60g4IscLRgh
ZzCN/GXx98eH6nHGXowx8TC4vMmYE1GU0vvh4Yci7DAEt1QkDRaDT2mNnLlX/1fR
16w2lydj8zpOHIFN/uwezwydqOfye60SaiY4hwZNrgZG1F7QGsc+Prz69meZ2KAN
t2iWkMFRZOysB4GwGQvV6jiGbvoH0NzYjnSZYcj/+oWYhfoSre+MTaZKxkySKLg7
YC9IvlDrRq3igdOjCJKF2AeRjv/keo0+8qUc2RHKDvxmRpOMwwWnuzqPj4jx/mVU
Nt43glh5uR0dYiNQhpkra+tKYJ7wvcN1+zsDv0htz4PhfN8H12+RcLNM6UsAqKKl
kIbyMiBneLL2qCtQJLhgZNzSSXqAMNFtjjc/pOA29GOpQy/SEiBTOieliMftNhXY
K2CaklUT9gubA5/1ebRSTJU1aBpl4qOZWOrPCjSm0fdFZUdrgr7cXDDJ93ZYj47V
NfimZDmMI58/Z1Tl7cDLGFxMJOJ5SINoPG9LKTZxSDcu725qbJbhrsyXVRdtLAGx
Dh7G/6GDt+UPdvSOrC6l8GZwRSYEPvI77JAecxbkro0G4v+1XfJWPtwuEGQfvPIv
qMN0qGSTRqaK5t+jbmbhXlMw46G2m82IpE6uC0u9DnZaQYRyhIX1GfVGqfmZ4g91
30YCNJtkKsi4Y43ulP5lG92gCgQFUkpsWDZj1UdjAArxgsS7P2c96B1wdhgM+aas
TS0MCupCfj/MvzhPqWNL6Fato8qIXwXFQVJidJEJuKuUubKv+YkTaTUZcEMPg2/m
yqvQ+6tb2mZv6gKtWZYDvJ8puLIiUTdfTxAgdOeOoSF5mXL/gEG0nMcTfyp/HQbS
R7ZKWSfHNoyz5/nRvxo2N4xBg5M71yEzgtbVZVPFokK0pLQWI9vQotIU06Q25IHd
PrJ0f9j7Wd7r5nrwpOlmlSiUfTbvDYiFJgGX2WcrfH/YlQY8HRk2q72eKjzaid8X
5kX4vrAxlWiqQfDuRCHBcPiKLGq3lQUYs0BOsADPIQjvUxtnVcYcpev1Dsbo1lIj
CxwYCCgPfpsvfXVR19sOYbl4WOmtDOCsxs25RwF49uVoRkuyol4D91e8TNJD4H20
zS5mdxvaZNwAJM8SNTwk42upuIjH/ykKcwlxNJUx4tikbt3VeULp+Fw/FK+XMMU8
Ug/TTJNWrlAjKT9pTl+NcZTPh3cZo3UykdCic2P7GgbQqXMp23RBLn5UBKh+lceU
WWq6xnl8GY4P3oRbIJwvEZB04i/JX7wx5Fn9wgS6qHNYOtz4MAE0VMJjqB/hJF4c
/bMs9Dh7lMqvtFdS6LpN9EjG6yU8brTHoyAN7Wbz6nQeBEZMvJBY7rcj1M5s+xYl
Q7XsFsaAuN+R/pDqhE9larKvs2KMeyZjxM3rhgejD3GD29W6dwUhF4oLGflFuTZW
Gjj8ysKwe2tEWHrev9dXL0c1BftjDtIPF7PfmGhJshF4+obtdrMZhaCPontE2qXi
PPYTiAjYYnDvSgh0w1IsvzkKg60n4EjHlEW1kM5nmBuXDOlL+4oaqHhwwhCJoqcR
4Rn3mKjYjdgS183BnvpTGZQ2Sz1SdIdEXi0d09nYF0zLOBSCQKX9yCmF/3OqPYb/
t6vK9Ya9uN9n9sD8Qi4gzJ1tMi3qFeeubwv5YycxRfeenfreuJY8QPWJFS24M7b0
avtoCEABhxQRt7ILgFAdzFniqNOLO4d4FAdyCTFPjLLpWi2jnjHZg9LZl20kLt+P
kaBO7NXaWdVzi1z0mf436mJhF/G7fwy8Jh+c4+2PnhVuQk4RlwJX+XAH/xeEQRqY
oj71BPnMQixCvPmN/bPN8dBhYR4qHie+gzeVb41Bad0CxuEj4V0zSdqt4ds1mMw/
ZyKhiilmryBkqHp44pTUztMzAFC9c5gs2tGO6omsYZNKytZ5A/URPCm/J29a5oMv
Uh+kI9GfzPQXz1/RWtX7xiufMPVzNN2s3KQ6MOfpSv41mr0Qmw8tpS3RtLQiayfN
sNQ33gfZlM8D4GpYLX9evvPiPGV8wZtjS931B5ulzygFzDFB5SOS6ewH8EPeMlkO
r2CXy6IlOetrGm9JksrbXqkt/VW7vsKXwUqT4BQbg15oBPykrLnyP7cflLams7l2
FJTDfv5OvP/+M6abIqznJbE9KI6OKmcWwz0tnJsFyi3f8nRxX7rwmmN0WwNsJA0B
chf0cA0WNdV9Mg3EDzDJO8+POt7DfHL2B7u1oA6GmXpDdgzpzTqYt9JdqVrUul3y
9vvldDY0XoJGMrJ1rHR2j6RTHbA+ppdNQGmkgimpac4Nmqb/ruryFKFXseBjs929
rE22aYyr278RBh6e47WEmeCMcBDgt4dNj4jJByfuhruG+AVlGa8sFud1KxzIjXeR
qxoDZK3aOzGXHuRU1cykX+thtXcrZ7GHPPIXHBvIuzjHEO/j4xYPVPc2RNBUD8XV
JqUDwL/DRLAnAkt34i6pgGkDDHJtJn452FJHwGmqIPi8GH+aUQikAwl2XaayTAka
nfhUCsVK2a6tzndrJYjJMzjwUp4rM4ht9WzwHM+QAhHn/ouJ6u3+kZT/hs6BkueD
Q+Z23FDqVcPQyhpn120jTP/Q4T9IjbhUwpXJ0e66jebFwxwKApBJ9BJRlrNDpOXo
LhRak5HPbgRGVrTBY4WZmw7YSw2zgqdd13a8Gp+ZxzrOuwj++ZTwRHFqvrRhQdUN
cbqaIcKyDflLByrjm1fXHDKCtbqSLf6KdEwOnxUqnPzaB7oqFDlqOVxR3GVwP/pl
K7NJN8jymW6vH9GJS3dR6LBcOe9a7PMFoyK+ElpNhNcRnsEDUHY9Nh8/wfXM5L8E
pNOwV5oRUVmGlcRzK2yWytUXWOJMA5oCddxGRyeKF8xgG+zBUP4N4mwMq9ob4FzO
Cox6HWAy48/FuPIl7BrV7MjDtgzhX5D66AKGVoqvXeZI7Jwb6ElNVZ1y8EuzuU56
U+dnbH/12bWIcvkLO57hQvuOmjXC5oDkVLgaqEmX8aJgIwXSLwx6dEXc64PPjmRN
hxw9hCYT3H6ldZU1q5nHAbexWDund0veTFzAWKFw5IiKRyh90DyDWl9SkNHTam80
PcHJbWgI6Z/uWxsf3AgVp3quO9vUWjIgsYYxzzs38th2CX5PiIfOkpWfnJWiEkpE
0Wfq/K6wV9vmW7YMtXseC7qoLK5YGNzbR71PU3qBfUREJADFbARz9kZb1c2DGT46
JVGrBdvO+2iMsRov7FriCvxXfrnI3GhXNCgAwrTSo5K8046yvuS8qTy/FWCBSmnp
h7o1pnKYXjf2AZVgadgmFYsXwOypZpMa+z8wXKSdqvObxjMcs/iuw83KK86Ozq69
GnOnksAS6AygkhUIXzwSU+AvYOlMU1kE5Ko852SnxQ7LFZ5zfrVFOby8BNRnYiVf
cmdNxDOAREb//tExQRyofQzDT+aIUUqo9QV3bLilDkNktCCQinm5VbfE3/G1yfHO
zQy+ks4KSAr7vqi1xCZgcjD/5L6X9SH6byKwGhYJ/cJik0uWyCNAdH6VheMscqyu
f71WBFiCol2KPzFNsxEbnxfpK0XjASdo/SPOZOEXHeBIqo8grY2oKvPOUWxPCyzU
4ooc9OB3OZUY0Wluat9scQOEprXAH6edlzyF0LRTuqYhwCSK7b4LNz5c1QTOIDJm
I0AU+tcwUPQSworHRLElaSCuhtOZrFfP/+U+VCOD2w7uldAaib7+vUsp4Li0YxsK
2wqMNM9qNEKOMdOuRNv19ycPED6yXAuaRklKG5b4Teox+5Osnm5OUq7vP0Mes3+p
LoDTAPipcpKl4K2LbC6znS67UNFFX7fNlezC13ijCGOK//CpWQsiAQXrOkarBLun
vpHq264AibxGyf1f1CzQ9k/dXnw6ElSA/UOGil7mpVt+bdqOUAVHZSOi1wC8bFaU
rzhjptgrgdQq8A0tPge4NHjHXX4OtgWajivaMp2k/rJxQEKUpVP6ghruTFabG5GX
OOGDpMwgBwbUKjSmF2qD4loOwayUMt18BsJyMCZMBoG3Yqbk2suoU4xOF3EuxOZc
eK3+oJH9uRPxRowUKrVpkxxm7hYUtCpWPd1T/GMKEPNKSgGu4ykHm0yZpvzsOmBE
z7uIWsYgZDGWXN5uBD+r0dk+CA4GSQ/uLjCfufPSF3kbZEvOVX21L9EZLnAHDauO
4uOr/yO3gBLYV/e4MVBdPsYXGsBypp9FdKf8AH3ejdhlgBeGv3Znjlrm2bl46cd+
q3iCUSAl0/j4ZtIlg0MfMubcDtsvwY0x09bJJeX4XqTJ5bH7zAWs0n7v3zpab3KV
b71ZDWN289gbuL+2Ngx/t9TQ6LYtf7G6HycQX1nH0UtASFgTiqFPxnfJ9INLmOR+
4if2LaTmdT8ItpyG3yxvs9/9D19yOl6fE+Cz8tNnSQ8FMlPxv64ZCPFeo04usOg7
tZR6Gii3gU9gmCXWBgAJJnmvaNk8gCRD68vosT4lOrfqUhC9lMxL7ZW+W7X6vJHQ
RJT1pm2BOCR6qMkWtEXPVGQ489Ksz2pNeeYtUuZMGSixZ3yvwqYLgEpxFYxnrfbc
fm9jMhEv7JUJKyHBR2AO9pf+gQWvhG0jmB/HRST/JshDSHDzeXCDwX9nVl0XPYHX
KScB5WzTxcHJdnI+GTnlpsDV1cFJ/KZ61YNwymwTAuk5qT4mnJvhUnQqkslqJNoz
UMdQ4mpdLGHaZPbg7fNUwzcgjOOXoBhE+qPqCr65KRQPwyg5QGW7f4G3imsCd2fo
czlRNvIFc0mY28bMjvyx0Y8nyDI13mr+RXcLQICXdxN6j72sf/CPyrRJMZR3fWPR
v5mlQBsjQGvaj/440SJ9xHTB41JHFQu49m6aasyWGozK+QPU2lsQMywe3ICU/R78
ecbNKkUGMSw/A2hBR1FOJYBNqhn9Rudl5nmwM4doAIrRZ6TEjqv9OQ1jQfzJ50X8
X/eB2hGnTgGhyG3oZbcW2q9tvK7Js2Kn3XSlOgACsXezQxdj3muWrcRHgH8Vb5DN
tWpFLGSdlLy0M1tFW1DiHwUpIBvtyONSxFFpEKYums+UHdbi5AgKyJfp0qkDJzJV
VJbY8gVuMY8U4psmrMq23bKq527ss3/k9Wdbq+JY3Q4qlfJtPXNm0CC5zYOtj5s7
6dEDG7eRkldQFLFx7BJjmvQlKKIMbysc+mZYT5bg/WJnGXKQGV4v7WAzL5G/d6a5
qDD5BrQTlhO9dVBnqw38xTTrUjTOeC0A4v4VUn8m+0kpNcowr3NhizWbElBhJ6vp
OdVs5M33E8OsvzieSwuJ0gBemK+JF/PNos6tnzZfsTsqm7A6IHB10L3ozr5BzzZo
VhrI7phfOKzGl4GyzWM1yzWrP0AYyPKjsD/RIxP5GwO6JIkFpybvtmd2bA2+CEQC
xRSkWvBTqUCa2DawFLhg6E6XHTnQIwJn2KoqnreOX5bTix4sEOey+sU56M4EP4C1
abQYoRmO7QPKelypoU7IURACCd/s9nx7vTJVaiMwdnKd/n9S8rlSrYP0r+O8ucas
3Zctv5+SnQfNqbO3nYlf947AYsD3BdxV/TJg0W0/R12YA9BJWue98P3PDfaBl+Be
/J7rN8WP94oQzNpwOexHDcx9zPb4Mr6HlloQnBXhxsBJbTY9r68l4hguwfnOILKQ
VdJyhyMHvVMnq3gIXawjv5uc/HzaDM6/iSgBv+5FSPasb5+wYEdhx6ck11QieHdL
S16raGvNXanZrq1tYHY4KSgm/ZSVG4u4TEt1oW/RbZdzjnfMrCqtsealSu49d0HT
VNKVQ3IX2Wr9r2i5QwEXdY8PIPGXUUO4rItiVyUGTFU0sNEDr2HvcF9mCbaFbb3g
Z1fV6ge5rBH8AvmP/XfPu7cVT2abRRqvMlbnC9tXY3ZydZewgQvwBQSphQEDVuPm
jlGvn7OTT6k8VVbWCzlmkcdRN6YLQL8qp43lo/VMks9e3KOfTzMwth5z0qFw9+dQ
MIqdrkapgGz5e6HS3Tn15JHlc5KPw6jZfk+fMzR5XWdrtY8+2UBfBK6nDi78UOLb
QvwCs7MJhjUQWwNgL4s8ZpkIKTLTU+GNkf1qp0oAYnhTRWVOmkuJ8f77nPiIZ8RK
GCu8BWR77BA5Co0PTQPe5Eo3puSY961/7vn7FLZwsrOOCA1z00PTwZ0cE+bKCgWS
aYis/Ek35QO4hrvPN76M157Lelf1bl7K8GnVRxt1jlOrg1bGx3rIHhLu8BRlwgS5
2IJbzddxnoXLRFVxWbZ/rwbtzKMPQDiVrDdaaMQyEz6ukZKD/EGmkpf+O+nYJQsR
wTdGbhguaTV+be91JRdPRcG+Oi0x3SOWlB1C6UppW7CRux24ajYWygCEIwrL6I5r
gAa+SpLt9Zj8CDcW+WlLZzgLf6vPAmw3kpVJwZs3lHtz6ugbYUuQHG04GrRCaIpu
PFW5mz57cXvpD2EWwP/9vkAuBsvegQiaL7bzEyP0qfErKNlQWAGnEl8WypeBF1y5
eM+xubYhJQMQFXVB53W5+xY/B2dCVqlM3JnZRZqzYZfQbIZKWn+OgoZu3zOZYwmg
tOxKnm20feJfxMqQ5wQzy8QhtlQBn+CUoB6PbM4iv2WgFwXZmFukFYMBA4zkRnVX
2M5HZ4LUZ3QLXPkOP5DaTFT8x+WlsBnk7JioTB7RbUHQPF3MyZJjy4aSC9ZzjmJF
ip9s34GlUu1oTmekbC74dcsl4S4lFoqNmmMfeDbnUBGEw4zOrJirr3S1m7ak47TT
x9vhbs+CC/0Mx70MruLLEnUt/905WvddxCAjf808114LF+67w/HwjQsE4UQTTXUE
71wLDvs/jHuH1WF0/c3yviFcT3tVR6KmtzShFrx0LoQpYnwj/M/nJL6iR+o3EXkJ
VUo5YJ/CHchRE9EpGXFUpWwfYb+wptga59blYiZOnhulyQuAKExBv9WL70CsSTkw
0YpQj3Oi2NmkvoBf0HdklObyqcs8F34XeZwpx2a8+6cnnby7dfUSN2u+z5F5haMW
g7u6JKnJE4NdaBai6a0Ia7RCKMcXOmsDfH3oyAJmQxAiaxqNbw89OmPn9cTwCySH
CVI8waiFeVeM3B7yTB93++ydsZPdZbzDBmQP209Gbor0cAdTb1uPM6rvTm/0qjdr
qjUSOfhNqrb8dd4NlZvjcs3q6g1oKTQmG9M7PK1TpalrXReCj942WoGjQ75Mds0S
vO6z39a1MaSMPtay9G6kozn69nWm1isecIl83Kr4Xim5PHvbQBDQ9iCu70dfBRqP
OanV9ed6tuE6XHSkU//VEoUWEt7iAEGXxHfSQnvZ6zxj2Y+IXsfmcLtLnFp5I2r+
2v99tbXh8oxZ0QW8+FbL6R6/1cSPoKQstL0/Bapovge4NXec3/7YfexW7w4t2O1T
iQF6kQwE1ytezofL7tbbQI5yn3uMRcRLwRYhtJtB83wlwmoU6RNbswaq5IdYQw2m
o0hgqnmjnIMO1u/SgQ0RosLImNxil+n5smncn+Jc7Ehad93FGYitordph/cxeJsv
cAxJjuQrKrTaFT0a6e1vkZFfxLBbvGXwtC6T14KCKi1I6IzVlk3qxCm+qhazZrQA
6nG11ARaZhp1NZ177vXyZ6DwsgDRMJpWrDKzU4qb1XZU++wVXJktUtNs6rf4JrYv
LtSZriieF91Neb/Un5K0H4IcFBXJ3J6zELwHhPZFpE+H7rEVjx6REKBPyx2XGiae
9yuPaoH6JG8XvSSMQp8TqQjiX0mSq/yKVsUxgcUwTPJlvS+rydW6CiJl+76XZnf9
SQdYG8tmKdVVP503cZBBeEnK47a+lzDS5y2119mza4YEYb4O/T/mG6SysrBvRas3
ydiDS7IDI2hWArztyJrSaFxbHwfQnwf0HyBMWJXbGW00cvnh3XluVzFBCmgylDJ2
MjIh0pTU9aJDhowM05chsGjYoH8betIZrhLRkuWWsgNAqdOMRX0MfWuYS7d84geA
3WhNUrpXprGpgNkZElPhuh4X26Uip3Lq2dzQ2794CcX/ofYVczG8CfDOm7OTFuCk
BhPvBvGGThuByUrZzIDXmNoKdWMe5k/G9HUfCYX6GpoK0k6IjLnRbwffzhRd3k6v
LDzjUSGUbZ1kqVo11udFmRrB3uDRDOyao+fJgK6z1tpnFxEqacDjGeK6NDEmZA4C
ZTbZd06umR38Ya+yaSA2dsCW9XxBQNSijzZiAHS/k4sVd/CwleYq9WWpCbiPwn5n
zD9chbFyXoIdXlrRajRZAdRfrhNf5ZQgPVvWW+vPvuB3ZpjUPp9KYRZlsgUyG0Tw
TVHoMrRtt87FqREzgk+Bn1I8MrU6YZQlI+ZncQwbZyIfTNnCuvXGQrT8ljB0MIY+
DOBgtYoBtAjsK7DGQQdojlQnY0egrukHILwLZ/gGtN6MaRb3NCdEuke6OUG7g9Cd
cqIQZ96AGxkVXvHLm5GllSJKk1XlpKIrWTDa4j38HU93yttyMo0L03XieoiJSVdW
/DV8a/K5Yrp4dOSw7uN3vFWDvLzPXn0GxSt6A/DtKCP4U2ZmyFeL0Bg3kI0SoPTH
qIq78gdOVZ1PNBOFu+SUsEcKTQ41gUa6SoacIEjJPMV/GDHvciGJFgUVaLnfJz55
U4Ut+wan6AJB8A72HCBGzZ9ta3hv4/z6hKnu7CRpHmkMwFN01m5MkaJSJmPJvWU5
nbiUsoiZf76h4a0erfNQpbgVn7riMwxaSgTVyVHo5q9UauJ4cHsmompiVeOWFNhH
vJqyWXlQVCVRHlgliotna7BiWf+XuRl573NencSvBmWAA3s9hl2qqaj0iP4wnrNk
QHbvLlGw9BHiuqWKYNY/ZBCFhkA9eCeCFP0U8JIJN1T7PW+StLT8TF4ieP27199g
eut5Ikn/eB5vIH1wm+i1CMfJABpO0vv0wbQ1rg7bu3pydP69L/8pHXoTzkXOnAtY
uNhnxWOXLDBq+i+k0Vvh4RQpklCaVGCqZvMZMrmDdgnD0TYLsaWul1j1F9vk6CBL
fY6sybMY0nbldwca/iOosX2PJph44eubg/PKqBxzjPSutx4ajZQHoG4rzxHhUONq
q4+OJLcJrxXC1eymQvJyasThXN1PH3FVYb3BS+h+n4Z3UGf2Q41fouR1alPpM7xN
ZFsBipJxbkqKtH4rHJfmlyoCO97YapJZg/6TppjbPu2sucJY3R9hKojr77TKcbxC
kC4WORS270dU7/OE1KNHqYsoGZECEaSdiwX6/N0oGQYn7xHdfBMZXkaxEvojoucE
+wuLZedXV/5kseAlXh9niJhyddVC+jIle5WiMBxtvH+TUSnwA5slQXo0xdyYx5pA
frCaZ8d2dDTeb0rXbl3Q91S3KdMKgUdlKvV5W1ekNbnDmrK4A9XiKyk5DGDf66WO
xJYO/BLUrD6zz2u1bzKKUxo+Oi1uSl+v08kgivDxvimNGbAS2XienkYrjS02Ijg9
V/t4KBfCmXR28KquknRbQCk5aK5awrhX4gfpmzXasekNfHayH4pQKCZwARbfqCKT
l4Lv42EHJ0caNRXRH9HiEMCrQyLuJcMDdr8Q8o3QvcGbuwy8zYmf/XRrdXSPRCrW
FXjPg0wIkOd+gpaG46wu1yZbHei2hKfAklL/zUAroPnyZ2Y7E+DQX2kKcL55IvPI
hFlUM5zofgtjpxLJWLIxM9x3wudb5ORKJ0FS0xTpUd05rfFBcwHX1fskeDmihjI6
mVXuAB70jcpgttEXBwIfYJv47ZTE++V54DfnSZmqUeZsSArdnFrxxENQRRX2gXnb
nJm3l0678nwJ+f6RFsCw47/lqOAeFiD5u9iTdgqF14DHBFz7WWEeeqJHkJTNrx9D
vixDl1Vfmn1B0y6Ojc3qOqiLO1X1DAb90rqGRyfB2Lg3CWBardC0r7ojw1b60tK/
uo2W8GebhBVqdGtTuwORrlN1aaFi8Bdy/8RvoxKrDN+ZxBaZdfeQJYnW8HH2Z5HV
dIGSmbMv4CTdvhpTXr2lV8g1AgAhPtReVnQLRq6NBlH6XVBV3CoBhwY8eSbW4Vpo
W1xhuTUmAWeGCHszBv+LchdVLV1CQNN70cT2h+HcGQjO0v7hZnAISkXoM3GKxI8+
/PhFXNB85lbndbq28AyI01iZLcy7kt9cfoaZUqElD4aHlSwP20OkYUjP6miM86zN
tusOchhbU2QgU85vCetgtdN8cuFI/vZMzPhJm7D8J774Gxzis8D2P+hf1K93KiY9
8IBO12icF0/NM6m4h2vv3fX2PRoCQUhT8oxypuXgI77L8EBY0TjNB9B4KRu118wC
x02iYXEi1KD84xwK9IFhPv+59ABRMcnHFitFlh2v8SiI9F7kgRy3uAjgFg9arQr1
6ux1smk4UStibBE6+YrYpLkoeVZ+VDJ2txyVpAlTdODDz55uAdvsLt69wp09PqPe
liJTC3mca19skz5sTCeLzEcM8bIC9svQZj7z9P/YJAekJq6scJTrVI3kuyhAqwvq
X7KEZDLuu41VfDKuMgaBOZjQ0UH7NIEm1yV4u+kkvnPihPw0CTg/E3xqLLAg/kL5
Op5rL06znJHUfu3h/IhGTdOD5QhNC0pSjZB+LIBc+VQEJSVRYFaMRQAGmijQ9Szc
70s4tE3orkX8c5+jWSTgp+nhvFcvxmTpB0Qfbnn9qYjMVFLEmf16nP92GNmJdFyT
CRibbLptt2qRDgtoNUbrzizVdBd9MqwWbANJ20YgyYoT91Sc0eI5VXNVk8Bw0xoE
EMKSIUkcthPpgic3ZdYJWQ0MWafGFTlijOZAtL/BmRjTPFtA+FsbhLLGBySSaJMX
8r1ZiBkVKKa+MJpGoYSGz0BayltFQ9QnEhb9TiHxvHy+qXVirdwyolzb28lIKJBV
No6DIb1S4L5W1mbaf71/BXVvsbfGiyslDuUB0Guvo1rAlAEzEltJ3ojjoYnL2Eai
9/xH1+jcCJruzsmR7ik5qJWOoBZbs/o2Q4DrV18RuUEPMFAGOAy1JjbKlmnh6Gyz
PIQ1r5A99WpAv97tHo6x8Xebto/ZrBOG39X60/VwCAXUqEEWFTquA6WS4/GgNKq0
eQxqUYvTn6aM/TDv9v3qRaumK7uDv5C1LxxjbjOkHyGb1qeMOEvJL+fCsZRrnHsf
t4DbtARyhUCfYsVV5pimOaShXdzyshzeTeSeoNTWrLFJ/tHizR5gvA3Vo14etJ0L
caEQ3N0OLZBVRsxayJGTOnrIso8ANNKGd5omliL8KFYZFWj45WGSiHderj2AoW3K
qi3at2mqdPrQGg1uD/OyapBX5hqvU+sl38jbgoEf1csVC6ii/MQY4D3GwwNGSbOH
sy1hSwdr3EHqW1dAboTN8i5d4mFCk51U+eG/CPsH/cImNLRH6XfDwwvdLn+l3730
fy1286AQxw/nDnxFMIlw5iihezrrfTQnjXUrlJMagUdVAyNkmkt1I7MUzLJfXORI
nJQSi7wDyb8mf2lraYQLDVHGMTMl/WEa5wqL3Cxw9JXUxziji9cMWM07HRxqvD/I
ixn/2q6lNsRXMoc3A1TGfhHfCNzoU91al1+MYfluzNMNyCY0JNcGX6OKxHiDiPci
Nqd7/jTvIHcPA/fY+lCbwnYFuguOTeYchCkGlL+TfSswQtYYfTLYBL65unbLZnvt
/OPWBH5idSyGVNjM18Dbo/uNIevAcfWCQWeSXZJ9O/c8Q0l4UhQHbHwsSFcIy3mn
6/tzKhcstg7ChGPh6bU/J4BcJ969d7R7jyw9g6pLzWt9yIbyjeDW9EkpsUv1+UF2
H2osAXGCl/0WWgcg0Ewnrs/tbcfTZNRruCYo/QNEpfUCsCVWRRjPDI2l1Z8Hxjx1
Z3EhEhKvVv2p11mhvG9CWT826hGD6vhq1rDALD5M9jF2HBoEQGzdIo1HKdmjhnRm
EyT1ztG/5cO9zaa+yFNpC6rN8eTPLVIQRNr9sjfvU1mJHMhLn+x6UgzdqgeMzOTr
hOg/BCK67X4hpng6m3AYBCjNZEmIWUKaREzanBEAydn21Ue/tAxDl+IqrbEPLTuG
4wZ+ROUDNOGvL2UxBv2Bi7cJh2I2BtfK8Ir/qc/OzayrGOrtjjof/VWOqiOzUw9D
zNYONzhNBLsrs/rw4D87WWqS8Uc2znmrfh8+AJJm4zVWrQTjKmafKG+v4hLgRRJm
XtAXsYXND//aFgrzuEMbEyemW/9atJuEK1PBtuMMRxW7BY4wgxCxcC7s2kTKzLvR
UHXDpMBE3Ol1euOyuprMQ7k7+Op8pApldP7bZ3WR7+vYd8bvTVx840w4PyxlD7Mc
ytCLUXZhSEd1ZRY2pilyCKzwjteWp7tZnVR1yYhhweQ4/RlXuOfD6KhJb6/VVnsd
St6YWgB88PgPlFom/cOFwSIqMq48xqyycnPvE3fTtKa8rl/CFsewBQV1v2aaGqo9
7YwhLzjxqqobVvJ0aUzq0OWaDYYVk7DtPMyJukoZ8+1W3XuCb85/YcnR+zxXAdbm
DV74N8TCO/6arTqak26glBQm1f/gPzOAjNITWE/5uC83Vn8R+mQLvfrNio4PFvrM
S1oS+xC/kPROeBiJQXKTnF7R/KcqnHJpUSCDc1VyRH++JRLpJhsuyYmDSXNzLc+x
hEbhhn+vHWXneOeXYkXJbHbj4OgqB819DBspFT41isrCmFwYXERIKrr37IPnZMhv
KfkDmicYUG9WFEoE0XbU/XEUuQW4yfaW+59w/yLgoUfzxdtp9KO0AIwSV64e8ZC+
KqXndh8jll9X8Kf+ytStg3JuaSglwQPzh1VqIwpmfqcwr3mXjepubapNK7NYkYPW
Y+C6h7DJSqExvXlOYlDuIDEMz64Sq6bhA0QqHcqQ3SwjB/6jjV4rxxkSoEN2VKtH
WK3I/bn/SYpWyHHoWUoneWI9S2U5xJXEGICBEe1Mrzs2jueFz6HknZfNbcJjD/2i
xVRj0SkzlE4tB10Xnp71+6YsFxefYE/Mkm2Z8Z6JWDZBhDHq0+rxYaBQobQf3NWm
Ah4LRbdpXDnnXTX0Quk+X17atwDrjUpO5EeAK+juSp6iJ6lnxl/WrpZYpNP8tgnl
YNONG6HM1dCxRH/mdCLIZioovjfq0A1VPZeCRuy7vWKLtKO0aBhDj5vV3Oa4SczW
gXxvCfm9iUumRl3T894RmOxWVdwzOW4hYlfBi4MCLmyXapfSr0gJmGqOvPe8FpCX
nKLtx7cVCbaBD2YNc0p5msTATmWOR/m76D0RgTouJvYS1ozXk7QtmCJ/iCFj+Tjd
xVBkoLa5E3z+rsa29ilKNt4dbYTBm1mijLbSCn7+1eYSD1snAXdL2f/nhPN8h0yV
D0R/oDjk3G5eaD8dFMGB/8S9nxf82iY8klEUR42Bq4dOnMtfo2Ti4k+Il9l0ciPC
beVsjgmnpk101RIB048CKGE+AiX+ev3Ki4qs+gnKzxHmpwrgUtpSnT7AMLRfPJO7
QaY+bKyyig9uIFoyM04hneIuxqx4+V4AeLkvDS7ZZrEnwZvRPtLeQuxm8AwGoMFY
sxey0y6eLtPehab1JQ6RchkkeQT1eBSRQrf2/4JM25rparejbmTM6drdzuIhF9jF
2yqG8noNm8pVYgyPX4o5acmbmYusJl9eOUnYydjkfEmahNbVHtwRZchVv0HhznZR
YZrLl4DUf7dAqp7YVA/GOSu2zXSLs1VxwnOp2fAymsisnJO9mIld2WW+596Osapv
TpGQ21Baj/cLD0Tnwkg2a4zsLvNyw895wyxueKk4UPCygxzQHp5llXeWcae5anRr
I9UcF8auaRmz1X0xehxCvIpZFFergUUYYDTKWbhvGr4fQNTx2ecIFyBjOYchG76w
8msGKI39x3qGbrcmOdjvgYu4Xo6eHpG+qwrD+FSxSkqmBLy5fmC1wTutqhnA2EP8
mW3m7iUf4XN8sP4bp2WNxCiteNoORoY0LTtma4iUPtpy2UpbMTClYywd8vXHIFjy
ZvUa+jwn7WBf70gl1UEKlBAWZ//bdGv3iSwH5NCXCm5aAQ1PrE3adRJgO2z1v/Vf
L7tQL1QJ2SJw3h29e76HZZ1QMzOjVfuLnhikUipmbztn7dnTB5gBgWjPFywMmxTN
RVJNi893eIO8WE7SzTz1aVopciTYE3wGKI1rxcb9mTmKo6KKVHIt9YZTwtyD3wH8
DoEejW1BjqlwWHe7b//E2IaM8pjC1K8KYM8YA0A3vKyRRk0SXex83bg3Ywd1OsID
7atpJ+oVwTPrXgSnnLC72Y1QMyLCRDmtimuCnCiULTef6V0e9qadCFv3nZZaV6sF
Dn0SielqSIE/EvDBQLF+6a2WKXH/YWISvWrl8cMpLvGgcc/RLAHlkwcByAZ9RV/Y
kvYG9aawV2wVh9/oKCsCHtfNqLeHWxprxIFoimo1HrLXSQiZ0myk8wufN17ysKhc
UMum2Ox/x9jEoRvuFhXMJ3iSkDIGvby4J09O4FA2i5JuA8D/Uw239OWiMWM+fcsz
xI5JsH2PJkPfbgbddf6kqiKRIpZ5c/RhyLenKJqyFXUbp5/546PbDdfec9gs3XlB
T8Cds+kxp4Y58PusHR/+5IVOJhDJgKuMa4jJKIoRKQxYXrQXobBlZGFqLmVckVTS
zpqJTb3MkWCvQARVFDU1Up+Z+acaowFO8sFZDpaNDVgP0DFYn0ttx6waT8AQ9ebK
ec1yqY9W6U0JingKkePVOzjDGXASPTFkIMFTjxyBJEhAWwqD1grfX8aXWqPzf3Eq
ZR0cljX1SaSeq696tGpxRvVo1tiveMcsS7nHOjXNsFs1nXOj3OcWBegHgZkwOv0B
ow8AGA28sGilWD44Bu9x6EHqCPxcwnWFbfcps9CgE4m20Y99RwbW4gr2FFeHU0pA
ztlbeXq3rVbQk0vqx5ED2UdMiN5lPMnEoCx0A3V4MtKlkumgw5fHLw9S/2lpCyeD
PmNvx+TCuDM+GaOrgl4uMvNVT4spOe9wJMsyD+6QyuBHvtQESmDadnGxrH8fmDol
01AMetjE4fzDPYAFrxDqE1zvvnSH3kpEiNtF6K5kFE6zd/ST5LozbwOFtuR1pbMF
+aduwzi8BlIAxDVqGWKS0VRUr+M1RiKP9kQ/SMPKlvTDA3WF8FmpjmUmsCqmtrEF
8LEocexrAJln2JG5RWNhkpewbLGkUaCxLOtdReAMuA59oXCi+09Sr49IXq2Q3WRq
H6DAr5XCPdzewkjP114TT5/zz+BkZZ8KGo+f9P4qOZcEtJZugBrwmuqN43Twk9I9
cgZguMVHo9TwTGMN3snDji0c9OjnHNwe6JXJwxcPjCTxNvOPi34kopgVq5vscTbL
gyN9hFfFQFgSa0uOU2hy88a5y69Qo3Qo4hYupn4OWPwjiRXGcjkc5VGi9/Po4w5C
gmzEwLfEPSSpBnSxmkodOx84lHcweh0aCoLEqfnXu66GmlRXT8NJIVCvNl4cvyIv
aNZPWKnNhLqu5yi+vCKyPQ/MA/mOnpSkzl2Xs+4nPLdJpFrdwHj9KJsuOTNwpLED
NBXVSEzI3XI4m5y8KRwXKsi1FJJ6KE8FNSkgVClr103Nm6Sl5cTGvCsmNZFz2jW9
DNZGT9TrD/6k/ptt02DHECYURCwb8L6eVrQ+l8ua96u6BRFUNngtYfqM7yEHFqkm
+B81zMq2BxDEhlWjVVciFQNz3ao6sg9WKlNb+i7qKXXHmFZwqDecU5k/C4H9rCiW
aqx2uADh6THCrVN8idWg3OCiIxz3dI8udmXPiUGE0LaTlK0AxO00usqa99E2h5Q0
IrVPNohCPUKAmdryvu5qDeeleT+NbfKKN3CgdLRJpNNRRs5P5oK461PoQ6Ux66d1
lXOhZCLE3pqYSVCOhyk8Hun8NOcX3OQ0hSVcIXuVwRNVdAXCnhI6fGrL5WB0SI9S
NyG7H+eQaejpdfeOlioB22z21v9Lk2Xx7joXr6AXrQ+z/ISbJNlmZ61a9+A6hiA0
QsTCtYYzUTrQKshhHeb9Znz6VfKVEjryicbnwrAQtiGmLAJKlXHqEXqafhD/pcSz
y70iVGFqaYBXU5PUxDkHqptydIJU3EKDU016s0wkQoxVJOvVB/3mby5161DR/EKe
J1rA5dPiPqT4ZPgj8t+X+a5OoDnUzyMJ0NHzcbVHthwZ4Sb5yt1w7uog+VL1jR1l
2eXJVRKOhCKDP+EF4rBbfttaE63SSQI/2TzuANh9kBAJR0o8OPIexAAIahPQV64b
/d0t73ow2Xc7Gtwp8GMXUeNjkWY/Wqonp5PoTPZtr1HVDfN8tjaEHIsNsKe64+G8
4ECLLdMXUUGSEzIaAplxUPGueL2NsBxXxO1csdwDNally7+bErUfzdYEzEqCt6n+
zHmvX2TrLXJ9uDumxS9Fn0ATrw92/upEam70eCgBlXQzRUr5KaAC4Wx4kPsQe82P
o4y/Pka1Jh81Gin5J6X/Ty0w+uywh2VqU/655QorTq3+fi9wHNDRgdDpuDF2ZzcQ
sEvgoZQKS8Xo0WdGnJTdEOlnMqQ57kcOy7UM7VVUi0ETJ5xKGAo/rDP8mLAKxTON
SwOuPLq9TsHfLJ+C73cDslk110jM6vCcB+mq5mcoZ+doGuSxJa0eVe7ePwkg1VfY
68k1UgvrGq+GL/1wf07if9DgqsaUjcYbVtkUEoACTyn+aTOEQP1MUdZYqbFi1d2n
ovb8+l7bi+CeVALk4znGEaSixUELMgnZjXIInKEYhx57yoLfXSm64zf+CtL/KkbH
s0pxyy8KxAnzbRZCVOyLKu005UiEvW+SPg/ZRwO0u/6T9SDR+inFLTE7RVYwE1WE
zCRk9Gr9hv+gTyp+umeKuTQPOdNhieulGOawuVR8C7L6lfRufTQIwVBVHj6v9c4c
lMnAySS6FB5i6y2VoQIFt/aYT50ELNHQ1oGZcMIieEBYw09dIoXJO9C4rfNYojo2
fvKo9dcxBh/9xJliElebWH+yVSmAY/vZJ2ss/5UcJIyu9FujMKAxIW+AonOrk1BV
FhAaAo1mbPt1OMctv+Q14PzLfIRm+ZW0R6GwDLgCxthZ8l2zE+gmYzIiIrqHQNsl
/iFNzvwOJWsgyduZU6pkFlM7qmTz2THvSRnN7fBfjJo3+PI2L1EazX5KCWpg+daF
zPbNKsIueCWbH3ZSQRV9AlzS7nAtEOK84K0Jcu8dPDmCqptpIYXCAYxpaDzSUDvQ
Etj/EkoHuX9PfYW1+byrBkjZYnU12mdA4BrzGZZil6iWZGNyB1ZQIdZ5i/WG04Sg
Uhd2lMLsIgWM6746QqdLtEaSBo3PR73SeTZO+S3cVzemY/mf0YPP3DYkNc9H7sam
YTur1agXs2qH2isAF41kKz6n73VYZ/9aRri62G4Pt0Z8TBqmYteMw++UMBLsNlOF
X7Y+TCFMdqp+jOaR3TRrtNXjEtx+GMAOjv3bM3FTqHLZoyKYgVtkWBtmsjfWHRqh
leUkYnYK3WrWxg6H7wOClJ9A/oXKxIyDPr2KXYYN4Y9kJ04zc/udRR5zzNO0iCGB
zsMJIUrRCo+qgYKnR8PxAHk2VtZgoTFg6ZuUIP0yPRTLy2YwitJevc24kYRdCLtG
VtDW64sddujcfl0l41d6i4cjckAnsu1s6ryZvkU+krFb7IacPldk9xKuhNzBzJ+f
twV0GyDezzfm+isd9d8Y1v9QBPXEdpga/DEz4pJc1ThqL68qFfZnyslrrzXMuo+k
NbLzErRoEhfyHyGzSTdMaELLWfXDAz17/mVi8/W/7ccKnG45wooOyzZEyRomk4V1
u7iCjRAHxW64uSyeI6zCSPXgRcdZlXG7RjTEjDsqUIU1OX7mtvdMpb+CGDtvUjjl
sSmJYshYkkavp01v0QsdunjF7bQHChImTbCPil4WA06MaIAbB2gVrmwbaBiC1FxF
amQqViYUZV81xG6K9JZR9eKoXcNYY4rpKS0KzyRpl3pg8jImEiQDqfQPODWwC+U6
rXW8DsxicPB+gP7czpMQghoVGMp7gzqRE2zMjsYQGaVsJEvFLWOEoPVekPB3N0HO
Q3oAbDJ+r5O+NzwavAOJgP10VMFub9P5axOuMkdBdPYegTRfM3iXdDFgU33uIjWg
6r4KmyHWHdx4FkrHPXuzR5aPEs+zlDNymykUJQCeXb3U36V+p5jtN3YbJoRh3aXU
DsG0yjdJe+jl7KLyRrsFyN9cJZ4GbUCyKEAeR8AgYW+g239j51FElUsdxUp6XFNL
ZtRGkKpKLFc7HzWT8ntpsvV78C69O9jqLV7+wd3rseMIgVlrIOn46KLAgLekpPVS
o2dQuIXdukj/BLKAwEDFcmtqIhm+6AUIgrZr89dCeBQ5UaKyznf9gOTswTteFRXi
6kiWzRkx6o13wE7BCUCVEh01yHPHqr2w337OU9VuAxEFA/R+iwNLBfBVPPtVjZoh
ukxSl9hAEuu8d0n/ruQr6LDQMIO1lm5RfO/B1f6OSRPqgWPJ74+De9ykkMKLRCuQ
5e4l2J7kOZkGbK+IbVrRRkNZzEwwnq6naM2TrEhXOGZDwUWDEYnb+8Y4Q75HZGQi
s+f89Dk6G4UUVy2LTaiHKA36BGMKFWjVBLRj8Bsv7LcvD7oRF0TeQkjSmneSHV11
wIFz6sCJhrqiFqbUodKT5IVY3vAST8iE26vaMpdrKQoSQKuQRTwRlaU3QA/iENT7
in5Wukwl4kpWc/mmIiNoLYvcYKTtJFv9FWv0OMEqB7n2x6PNKnEsGyS9ImfQGmCG
iDRa2/z99cf5RZfGS8hOIh/v3Gthli5lDq1inuuISF3OHcuOW1DTLaxZpqq/0jPK
7EjltLHZYDNTP11LaHYiVKuazf7CXvz0WOpn0WzGveJFLhE5I+rQdvRWtr5K+Qj/
C2e/RyN78+C8dN9+KfGb5I+J/GIuqWwFmdMa/S5mPKvLdeetcZZOKpuWa3exnu/M
2+CXbhZVaHTVuIg7qJ8HkRGU9B9iKSuAd+xSv0hNTOCVVD7Homgz7tRn+etuCOLE
2EAPA/lf93NnjmGjiZaeWD1umGF3IQnajmB7VF6HsRDgKaTlenCFNOSkLx01HlJw
2AYHDQYcV/hC55org5u/mqt9kLw1MMoPskNJBk0utS5MjxBGtIcg7rjDaOjKfW4G
ekEjsbywoEptP5j8IxiTGXwVRsTisbcTKyI6Eiol79/tw9xmVQoNiU/kqvaTqFyg
hI7rIEJUdCX6Zhdfl43rFfphv5txY5OiF8QFKQ53iubNLOVUKRrvQDrpFKKrboDz
j16VDLULWdEZ63tn4ztV7Bd5sArnGI0KVe8lrP8TMOZNGzTYr0OJBc/p1MnhFTKj
CVjVkqOFrLlELgl+BEt83DlsIKlQk0pn6pSH882yL4jyP6DpfFGcNJTwpH8EnARW
Zm/rFI+SfbwYcOZgOQgCk0C8JXNrjyqABdEjwZxtbkk3SdzddQTAdIUSof09MzQh
hixeht91QWC1VBaplFLFl9EWQqQ8vET5R8VQixFkmdvXTXRaSprDGAGOBijsTfi+
lgSPMsOzDBZENRdTlMHtOinrh4d9KR8tuWa0RxchOG+Pzp4C8sKLPBSfBF55naNj
xg9CiaoYLS9tlz+V3n1TH3ue3ftVScdIAuqegIMRJiuzE9eKdv3moiYVVtV8/DKd
ZFcNccl7Mw25uQryzSf5bV1KiEzktLwJCykr7OuTJ+A3lQ5GeGCGvms+x0Mg4aOB
yjXKyG92h1FdYvRJTKaOr64zjIziuQ/L4620U6bCiHkcrBMbFiNl0m1KtiylvkD+
PdB9qh3iKFUc+k2ENwS0QOz9jVB3HzHts9m+a0pFoIKtklkRVu3iGdIASZJFsTJF
PP5yw3Gh5xxN0W6TTmYYCEXly1M0XU4NCY8BIeqIwPgnsUNiH3ubuHHXp5LvgbLR
rLaxywu67m0MGKh8OvTatz7fPZyTzftbVSj7lbsDBNyM98Pnp0sKUQk74Vj9b7uv
jVPzinwASXIQPFKBAvaxCOoQYIXvzh3UYYTrJQYfLY7r3o0m4ofbLep6BHOYIP36
rz83ZopZqzVCBGGkcBoISxizbSk+o+4UffCD43+7hhaC5p1x/uvnTUx8G2Itr/e4
TTt3Vid04B8m9mVQVY4BABPCnuXF/mjheDTGgoJKf7mMsttjulrB/11wSTRLoQKo
LXRmxmgsLnqrzbne3X5wwHAzdBvfPjvQFs+Houjun9RtLGcnreN5TtfafWPQaPgp
MojwbQKn8Xt6iXk74i1nDyR2KwWYX9iML+fNv3byAkquEAtnEfhYnjWIBZzeLrGj
M1EqXyGFk8bNBayKMS6VJ6zql4s3KsBfngZbJ+lTagoID3phKAFe/bdc4K/8HYDd
4inVOTRWduHOlEmQnCb72c3VMx4Kd+SENGDHhoPetIG0977Jo+RSdQVqVY1lgVyF
IBTkgwPwzWlK27+0dbtuk7YR8neWxlKz8K9PzwhFLRTY0ert8ygnmRbRfUbObOuI
zV/uqmSZK+abbHqHEw8z2Ys9F50EWdwW8Fjor8GYZ44yMhq/LobqaQ0zaKNWsf94
bR6QkgPUHWRGaoGf8/zYED4cpvYcrRGWPHsNwocrxoADn/PWYXaV3qYvafCkpOtb
SAwy03bUx7/NPhI8ZuG1pufUXTNyQdVjjvU6u0WZW0GYooO/LD0mVzXk2SnezovO
4uUCLvlOxQ0RyGhtbaxhQ2LDyRXXDjfp2OdD9HpKIkpRpdAP9m+t9A8iD5dV5a0a
/0BrZ2CBTm6UyFw2HjIg73SIqsFH98MFEmgzJPfMhEMeJxjjUA/8u583iUvsrgtm
S16O0GTSQ3vQpMD+mTdKyoh1pIkZa92cHAKkwkDoTzZXuNpumjWG4fz/7dCgoNWz
C37WeyTz7K1382l6bQfGRRuZgQJO5ovg1Hxsr1uSr488M/Y6YkyL/VxhK9lj2JkQ
eryKw2ORggLrURQhubJD5dI6Pmpvwi3y3ClJllkHh7Edbftw8+ZVq+m8PomgLy9u
OviB4L9VWFO/SRw63YpwTbw/hkGcHtItSRPE6w9WOOyU+U127TsrwOha4Bw3uVfG
7gsozebWybrKn94Pn06cYHs3s+YaxQGF5qC3KIMFkFRTxIogaMxZaqOdILRw07FD
ICtjd8yZAn3JstW+YD3BEkUKL07tajZ8vK02a1pm/bPoq9zCBl/cu2XcbOIC44It
1awNovYzIfyMoFMcHaQkRyzRH1Est/piDyIJGpMiNvhQWYegduFRVPBVWROyw/n7
wbEd+AUyv5wsuDnJduSkV/2+KCTdV1fkfZzPIE59FOfPZ/LWdat0lGA0VyDIKGC6
ZAFj8VMz01JAgY4ag7zN6bO12sDKLK7YcvqkiNOBi5MAdvZNV6z6xTHrlg5LliTg
SCDCPAphDkazkeLujICAgrGUWhUVZjHD6fxXooo19kZqxjuHg7pufomcH2vD/oM5
H8/vGMi1TSN+vk1fuWYVKsxDPMwwV2JoCVPA7QmuCCeW/aJ/IwkGehtpkwUDxK3y
pcHVfj9cxRTi9/qT1W643rA5ax4gMqqxoOayAje6GawZ79dylUkafWlVvLCX8rT0
naToVv5rVVmcyXc/TB6ErS1CLjUGGvEFOLaJ0oeZNbb3QEitZjrTCfAQ9sBXaiPm
PzWh4Z+NRYSYi89GoZbl9r3Ff5Zp/4AWx9ThnG2y+FZlPYqk1y5t/hCaZ9259yPH
u+t+WO1or/YI7ydan2FiI1Z593m4hpKMc5lnx8cghoDzdyMa2cUtaCufF5nDkc/w
0mOsPczPwmq+L85+TRXRijL/9rGhijz8EwLVuhl7Tc87qdaIo2d46i+i+zKbZEhV
fBvALETyhbLIKaKKirepY4dRL8jlIC6GPeStg5MoBxw76upLFKafx18tEa4HYn0C
zIPsYnpHj2PNNAaGEatoIMUWNJs+JW7oPzVyPVuvfEUbCxg0kpsoqk3Ll0F2Tg4L
IC2oXtMSgRGRHssVpc2hBUviBYuDo5cgg3jk3OA6Nll2KyOMZxzKlBcrvPd+/u6l
C4eR4718J04Nol35CiJSfTBj8AQXqlblfGHe7qsaTThdoAdbQoELcEdGqQPE35uz
Efuv1bt+m6wzkuXgJrpuvVoTXIA0V5Objo6Bo8yRdPikzJMi/hUgDx/GlKjyMEOA
ePGqMputIb5gUHBwJxS5+KUINBSEne0vkzYTtaoIb31vyqTN4oeYkHZM108lcm7k
muBhRjfpha16Y5AtvOq32tPo75qA8RJD8GqvpY5CMunJo2f+5Z5qBG9Z/E3gBCKR
Kwx9IdQQmAjmRc47TeEYfVzoMTYf2Q4+qeKTuYYCdJUaWnNfKvgrQR3QdiH0ITYk
LloUS51iYD/5hgey6dCl/7MdnoRriQKMP69fVc9VtCwAHFOhtpXp4eNTS6POQ2hT
SETcxRfoNPhampWpCNguzVaYQDmc4bovIGf3iaPBzLlS2atvtsi1rO05Cm9uXtul
KTQyO1D5Wz5oym1ilXzzRt/7Mx9XkOlNGw0dgU3M1GAvzYX6uwCCNOo6shaIa1Fj
SFmuVIqPby+T6dLoMUyO7ekV7WCdDbxLqTcLVhdvOIKeNhOo/0HcfdKk8zFX1BUA
i+U2xdFlsVXeqzZiqx554bsZXxSU/QoFqVc8QkrS9pj4UX1y0lAMNpkbM9lqHQya
WaE1p1eIzPuD1cZBDxu7wruSprhAYxfI2B1Btm8rpBEvjM6l+kaNSAYWkBG9+XS/
pGSHpA+KZdSFO8sGyq7Gi3+j+todZeMgP0cxBriQBGjwxUdJtqZsjbhXytJEYwld
9SM6FYL233h5PdXHhRUIyqjieNCNXJZP9lrA8tQ574We9AJNiDkn8oh09QRlN5KE
9fNsA519om/JXahFEsE2qJuBI86EjbpmjWuxf6jboM1gEbkXUHXcK8enZAndYduS
nW0cjs4IWJXlO1df+awMmNC9PiUl66DFMyeE4pa1G1jLziCEt33nhFZhZaPCf765
wO/+Gxd6eq7QNXzEU6NTyZdxg4vrFizJPi0PemVXL7pkYmnD9Y/nhfrWXw1wN2x5
XjVgjbo91E0pCyE9LKUyxju6bNK/PnZahnMIsJVYNV0V+frZibinmg1HFZZMJwJo
DQq4Jdq8zwEf8zO4HMQ/XYrbxF8RWTWSauEHqU87tEE2lkILmFmhXrWJOT07sObO
/GMWH8yEAwsytEQGM1ExDAlDuyjRFjQ6khHaN2HYv+Wp9XUMeX3J3xAg0X3Nywnc
Cpw7NMcmdGlHcl5WQiUjLx1hsjIrsZw4tPnfOyLpyY+T/Tx1qA3KGyKCRX9OzjX6
leXs4TbUTiK+yHD6GQqpEffGkkI/LHg6fjY0G3fJ7iQhWBNLqTheOYgxbVqa6LZE
FV8ivwp09Du7dk19X5q2fybJCWoY9MUMq11+ZkkYbCMmSHT92Fmw2oWeCLRID+xo
odYlaz6F05ny4k0+Ya3Owi2PAuaK/IooL0M6dXloJBoXXpFsn7J5xWdjc8LqLXux
0RlF1ENtMiCg/7sUf0EZDqhQI8xyc2qJuJzuJrdLcOd8RZF0OkgYjKTInOyZASAL
iAMsLO0q0t4feyriYT8WyKBKjDkFAwEMcNaq5f8VVESgspeC213FKr+6wxTRycVu
EWwe/rCXmAwgGClMI/ETjHkNiIZLEinjjEFTyi2SqJiDfuG6va2RE2j1lA35XGw+
QluA47/EJyylgNBncqrLi6XdoxtLvyNLiX9lByOY9gvuQ5zUtPSKvajr3YXWrlnb
AJAjNTuc2oC5cy1vA1S7dhGRb5Ra7bEGXOu0sZvwGTD8SDk09ie8SJFoQykgOY4G
DCVhRYt+IvYeoobvZ4/PLcuUnHytt6Mpwhfe0SPnmLizKgDgsLFV0r6QZSVcu4sc
gIL3jaCJhM1GugflT4TiOLTSJ72vdCyu7c9mrdY7wav+8LbykwRgOIrtimu43Fd+
Zq02DIulmTJlVYiA+yBerz9Et7jeqB0gH7KNTtVC34OyD0U5MfQ2iG4lwD4obdV2
dqlg1zQ/rZ7dlkZKsfBgTMf2OeEsrFAqmQuRfTOyrIsoizRDGeFFn07rK76EmBwr
p9Ky5uDSYjTn2LnSPDnfYxZS8QCeIHIV6FIwvp1xbunAEXpOSbsZmo/2YmlYTYMW
IYxsbbt9u8qFajmDXdbkuX3RTKOTFSi5iEkIUU1XctLqkQqvniyjzxJuNOzlbM80
H8SkxoLC3Ve7xfJ1uvdasZR0TOdOkRQrSdJr4yAStlVoARCSP7vZbuBpGeEXuxgx
FSNG0tP98DnmuijkgmJEXsbnE+y8mGhDbpD1C50uQazn4mkZf4pahcnORT5iJ/Do
e6yZwBrfhs9M69QvGUVKin8kdMlUmUZOok5hqUsqoyt1aMKhOMPQwumo5NwUVYRq
OV7EZBDb0vA7ykdRb3uEOXYpCnjZd2oeItMowgMSQJVFHGZdF1Ysq/aCy2PJlkcg
rZHVAGlOEtBEFx2Nnwa19kKpLZNaw60bNqz4Vd1XTQ1a3mlYMzL/q16vNoCDTzfj
3h4DUnYWdQVovAZ3ZtLd3TresxKIK8QyiAQJMEWWOQC7mcNfsbfZK4HFq26kZYl3
36RmMG2O2gz0wxlnRA/L91oF+zK+vpcuyQPgRUdHWnTfelwjTNMgz2Un5qog5E8D
OfJ5rbj9hHVkDQmnosK+2OcDU2W8eux2pWy+4K6d4yL7GvaM8Yt0doPuVkvtGr+L
pv6amfBeo8bwCeba+nh+axiRsdpeZl4RvRXcWGmkaD5pJ6QxG/bSlybgD5csXggT
mrq6ePA/zob1FlnBHmFXWyzjPJ8nDoRAP/swpPfxu7UZCSd3aBiatzFhOIng2B4I
X3A83kJvz3aUrGDOSWCYYvESnPLYQpl+zPB1CoK/cKE3Ilo96nj8dCZ9A+NNKiGR
yaCkGUqXFsVSkd8U8PlU/9mMocLLtS/wQsP8Zy8H2boxQvE/RsyoLzbSdR1Km71b
mnCNnJEoM1AFyN+IDyPzWG0Ew9IyQxaIqCGmT33MhwGTRvBQu37cDkZInfTQMsUb
OtHW3M0OiVDdCvScs6otcpsHHYvJoW+xSz1RHerADxrVoO/oAR6wyhv1kYvE2mLZ
21ew9xzJ/Fpfb8xJvzCPgqcR5FHOeOh+Il+V8YSBjlwk9jpm1rgV2qHKFMIO1X5q
0fyn8BrlbdQBZmR9ic+PUIaT6ey2N0m7HJXDh9TSi80WnDjZEUK1OtQkyKNcEwZi
K64eeCoNk15X4K8ti2VBzmTCMFvjxWAFlb7XpfvRNWKFv2/RNsy/rK4Sd8g4cGmm
Hv0kI7NsN4eFQ+ich7tCJoyy5SH9hrwrMu0bqL9jmA01mJhnCv0HkT+9lffzLH6A
nEFSABOSpvl+VvT5vth2S8TOTyphuZRSyXL1y04i+e/dbUSxYQ1KHLw2/mVmHtZ9
4qn3jqMV0wl2fm5t0fp6FIjPOFS5ZX9uNXBslLOrQ4jqYAQKB43R4M6sGRbPEDwm
+yrYQgii/0B2PX/+gA6LWDVemCljUMccRBc6HUlypD/cZQlGdR7e306BoLQbgdaW
s3QXSF25scnDWHeLi9dhF58StQlQ85KUTJSbEa6Vxcwn7MJRRTX8hiw2pvPJSF0u
m15LmSeZ/Mn73XKYH6kUExOy0AW/LIL2zRBkJZBitSvtljtv0ujLvQgip+A8iQBP
3tJWxE+BUZLjrSKs8kOoVasKX/W1iJ9QacOx5BFVaLYsvZpJInNirLJyDB5n0IOS
u09AtZJbc7Sdop4g57/E1RFRzKBy7Vdv/egfk7vpm0XYua5Dhlqvahfwur+y+5jv
+a9Nfowmdrg2YvN3hBRJ7zC70WeLz1RElpxxSuHyVvwF0FJRRCWtVxc2ARGK8X0x
5KsyGV3gGL/bYR1fo7qzflMz5gyaGhPfYV28vqvV69UdstXnefYYBmjV5W59uePU
JxI7dINI6xp1oQzE2kd7hC+wv+N7WJ1kh/SqV/FpjPLZ3CiiJCNstjpyQdU72Qtc
LK6yylFs4ND+MRxvoABFMpBHMsockxTWAxg/JPa4P63JneZIDlv7gn3UsIpIjS2Y
sB70yLVm+AG5EFc7ip+u4+7m9my76+Q2uSAjZHVFzZ1+43UraF8TqiJ1p2SzCpnM
ftAgGHvA9AOSNT6w78NexQU7/XAlqGVZgpjtigbSVaVbi0rMUnn0fV+8jefRb0DX
TFgfmh+zmTSIsbZRN7yAOsHFqI9565vdhVHbvqHYl56S+woVCQvjWAFeEquo+4XY
scpwkVjwbj78y1AiyUhWjK/vsbCwJv3CnU31DP/hjme5RUzhBgnykxkBRxczHI1n
wObya3BYFgBoVFH9qkEXfmlg6nGUEb/j34EJQFDDGmEnSjhrw1RhdqvXAxDnuiT3
jocn+33cXLD2XvkauKuNBaG3OdGSaG0HRu/kCYQa/O/G+TVNAwB09HqwR7lnthZw
r4bQ8wRcDVoOSau7jd3EPxNQKvIQ634y4ZGljByhrMQE29M3/bDurJkQ8SA9eh3v
9ZqfSI6jkQFGfox9sivTvLzFVo+t9s+upcbgZ/TeT2sOdcBTk1NKAFC2K25C+KJh
EO79MC7BKTgUpcfSTELu8+43zfRiC1LwtzJifUQRatV1CaDHpx8pYBwwu2WZ/d8t
sJq/U74DLt6EqgpW38wIN91oWiWGpW9cElMZW1nZGvty2yJVzytl9FtxNT6Acz9G
c+HU+Zo/Ni07zlQA4bd8Wj/clI3r4yqE62mDdlAIl7R6JCyEZqw0s2DcJrsaxmIV
U1vX/n5u7HxuQ+WjPFEgRRPx2LrdNkq7y9Yj7aZtWk5CHMxLvBZMttPCOlShRZ33
oLfYmJpgOb7aSJZTLZS0MDU/0Hfclx6U+LYYJwPlmhiXCsrELb7u7GprWaUMS8WK
AKsBQjq2YsnKnuCKpfZ/+6l08i5Su3EfIryA2+PfJhXcM/KOizODtwlMjuWYChXM
6/7BUVZNtREO6KVxaa28jRKcAqddV5JERlEfEiD0Z0zTeKBdMB/OsvmUDk/YlZfC
qB/MLjMK2H1Nag4DKMA04Cq0/xkVg0+zKJjoMKx8LVKFTK9fQZwfY8dMf9Qcula2
ZalF8kO+YSU/CpEOdDq0+aTu3xgBbzz+w8A3f4GERF0v2D27afCblPVc4OIBJ5cn
LHPGuzl5lD8k2zQEGBBwRRZFKhB2MHYyYT75Xo+7N5P1vt5q2+gJNyNa/TLpKRqc
VC2dXt3X1M+RQCkaPvpIBvJgVxZmqMHZnw2miFea7r/qd1eK4rX1wTKfKSTOIBsn
g3jq4RaqQDPiXu+DMKVRyXz1fvD2DOSL5O1MvRMnux036QH3U9+u5UcFEvCxBWAj
Zcv3SXUM5Wx2tuQ21OvCdx5sJdscVxLX7UU1HgNE7vmvwqKFRa/SZ2AMb32HEh1V
REOhL2Z/sUWx0MqIIXUPQXqhjgP8KEaLLKaDN6oedeXnQ64kuPJBwSidyZTY24qM
l2+d3nLAABXxzGrKqZdkWpfCxtwMpRShVSbEuP17pInhjVn5dXJyF9aLjFkW0Ea6
733myuGJIOQbybUlLnxncARJMBHqzdowbu/wFamYumm8D3TDOis+Vy8kCkOMrqAl
3EOx907+1JdXFViGIvFUFvjPA+z3sqtFA6TgiXZg2LyI9Cx3ALGTi0sNol13BPCX
tax7pKwjg9rFvmy4cjarzvLZuKEEvgWlNwRVI1ePXVNN8rcYELG37Ud5WMCfCqBC
mYkWLElarPXqlJPcyhbP+TbKxmsJiiqmjNpfzJawLF1LbRSqjya2FMObiUwM2qGP
svMV0Z2JO1iCmfVUqEHxRjcWlAJyb/CQDHvLH1G+0aWgmFAQZ0lt+pqiJXLx6WgN
1MySd84qSKYOzr1+pnCVYivbcZmB5AbEQPaTBvaO7okHCsVoKRTac7IPod1OrK5W
UjPLMHTVCdvSlgovB98Kcw3msd3+/ZiQmt9L4o4OFWlNhaWfzTP4LluFrXlijk1P
yp1IAsB9f4CTXIvvh5zX8X3bm3YyThid4ecWSwaI18arDR1xmIAuFJfc2K56mD7D
ZgDQry/sLrTcHnE/zM/mrXcfImdZPWZnaHipWbGtP+XscWkoh7kSfEPt2HpT08+9
B5ixdICWONO+skW6WxA/wKgPPCe2226B2wzz15FgF3rGC2R4S6Z5H9+2dseN4aIz
cFqXw2zgZNLgPihAkevL4YNhbCtAPgmXEiJhXz3Tb4eYTGS7hTKKQCKMf/6Sre4x
VPzh6kMnNbe0rjXU3BoM3uZYIHD5pI7o1dUC/fS2+6sSOGovTP9OErM7v/SstFzU
DObe9Wo9J5p948KthrEs8Xk1pn83YOEn3kbZO6xUmZ4LrBK4WOahlmeUkxWypuOy
JkzA652Th90DyeetYLgIEY+OTTg4oNKVirY1KJSoTtQhIX+JYTH8HPURqiVEt3CG
VzLsEO5Kj79vNRTQzNdtUvOZsTL9E1IStdhG3VK5OmT6qlNOFr/wMG5xLLyBAjQw
qk6R1oUTw437n2xwx322pBVnMTAmbAgjXf4tTs6F/S+CiuQTfi22qvHCz1cTwJHS
5IlCbKZV0qjUtfeqU0C0MMGb9w6Ao2/GPRXbUFnL0d4YF8BwGM3iCz4UxGdhUOfo
/j9kh4xcqKBOPjm+TZi6jt5E37muy7unpHzuVXMJL0P9qA2ZUrPwrbjoVritLp1W
M+LBs4XsiTzCUj+ntzVfqXQSu5Un4R+e6ZQy1fWbdkJBfiOMk+wOA5UGhvcQAjlt
yfwmIFno/f+/gy2lWrbME0EilVVcXqq4FtSw5k4WbLAnqZENlKKFx4R4N/AaatIa
odOfA4SZdjixIsKOyUhPd0sDfh4m4FFqcDebcQeoHBNtfY/jOAJBa2qzYwVB7eGC
wGWe1O/d0aUkRrl2SsQ64M+Z3uSqsS0bsEmHsEr60dB/tzhPtdQ5JfRHwmbi++CV
oXTUwbdF5qfsaBLwLvuUliDcz9BxHRgzQAZRYzoxy1IUPjS6f+r0bs+EOxA0TeT5
wevBVtPSuArDna8mTuTdNAbvccQgbLicCn77dx0ICGvw4iFV69sJ0VJCpJmSPmco
koYs2Jsa6t4p/cke5jg2EjohkddMGCupBNteZjzq5knW06ZfePPVcLhPFa2A2eNh
g8xZeYQGVWU9fQJ5OOjf4HtuCsxUzUDuzBaJMOlcO9BnL+/4lvPUEh+MbF+rgupi
7kUI8XZ40+d994JaI04GHGt6r5pTNv7907VSaMEGokZEM0npt/XgotP0pWKMu5Ov
K697o/+I/SBcSeWEupbCuAl1Aa6RSSi0skV1gDMJHSh01E7E4nmZsqdL7rj9oqkm
I3dyMgQnrh0Db6ooyK4GGmvxRuWtmhjWo30q58HKPy37CguW7EZYgtYSqgBz/sCK
Xk0orf/ZO4ioIPexW7WC2ICUaGUZpaMdK6BuMYC7bHSvwlzKGquX+w8959O8rClx
t9ri7jjFoHQ/cYAi7+CnQDYDleBYiQ7OKrHyjjQZD7C0rhcPmMznXpIp0jF7DG7m
/Zd903akqxcBZJYuFtN6bponW6U4B0j6h3rYYn9PCoqPnmWdyeLsc/EYpg8SGIGN
zXUF7v/fkCWEeoIqL8AXh9okUDyvIwiWeCvbMu+69j5wzwIFHDkbRxarUB89wfPv
mJYSDbVOuZf7ONvpCYEopx1wnuuRUnW89XrZ7+MRaVBlpvYlxMopc/t0dreXAjrQ
G7gXOJWA4OWzuzKlRk+R1usV5KiPyoVQQrCbTNYCYoRCOJ12NFkMyiB+4v+Vn5eM
2dkzcBFAfgoreykgpfki+csUDOgwkar+o56NrNQWDZJnbVguK1CEJRGdD3QYFOwa
JsXdcuTpBJjmagVCP124zQZYKi7+ZP+K3KlVvfUhDJgsT4D2SnTDgXTGb3SHL+vh
YfF6MAUF338s5PiQdw8w8Cd2zajfJjvYXFiRQKg00h5Y51HusscjF+7eksgTifS+
FGNVtlkXc3jQkj5ao8cSKDw31yVxe6aKPWT9vqIV6H1y8erYSCD8OCPQiFzjJ+ds
KgzHiqRYrwKnmzOXLoJFF6R0FQR21vxyI26jJQQbPTjeO91KX9ENh4jo3gC1le0y
VHoUz37unZJUa63ybcaKhkK/35g9sdv2GzU02KHA/grwPG9un1WUb6Vy/UeNYcOx
1Sc72N42BECoVJKy7SQEh5fz6Ahma5gBTYdeesNYQMBGv8+MZmuU57Qv3/OQoKve
VO1ZPMgG0WhXVxJ0OTVhMYMAb8Iidpr5ldWn8yfplPePmrav6cepzO9m3JYoysbK
z2XVkbViqXxPmr6+pUtnSqqpTLAB5U+bJ7+TbZ4ICgFt0hmc25zekJphSD2I6Q/2
5EyzNfzteX3ikjoxIBdSdaUwxIszfwwznHwGib3/7dikBgnmIHu5rAzupQu7Sbdo
d84PI/VWXiUXP845MyAxBwyoocleksOS2DExSf48/CQcDoyPCtyHTyn552CmfkHa
TAP5svesMeRZ58D/8slk/gyTVrll2ei3YUJr7cpFEMVQhTr1HX7C4LwgcEygLyzY
fv8pO57Zg/QIJIrzY6ldODA6pnSTCEWfb8cFYbRDalFssUk7DC+mRucERUkS98ye
feHdxgL8QhZaINV5KTmBGOGIacFpz2Pv5V29viYRfYTotDbYn6MflZzh0yk6EICA
oU0yQ81x5AW/Y7ZMM/IXkltdZgvvDoGEAnYiw9K2xzbC416ZiLfeN8i9IEtJkzPH
I7oS+6TYZ6W19tczvornWjZhQalPDuxFZFgBG7KW9F2re7onc0qDeF/yYLxDWh6i
88Z7LgZRhrerdspDu9TXYhMSE1NJ74XkUMPIBCx3iedagu7YLBkJHaxkKk5BnPDt
st13pWjCJeh2K4bfUx6bGkdN0DVNVbKXCyUU4q+2qvUJmvQachCKfHeM+/YX3zuJ
Vc21sjyG3YXM/YeOGwJpyesuabnd1CSqe9XMifVtqP74k/BzcyATSAJBnyaiWk8/
tOAQyLPk+m4JXgoOWFAzWoBdaPB62KZaS1wflm7WMuCOrDDKeA5TlN/EHgv/6pAF
KhovkWCHAcSZGwdDhWr3/PTdXSfUlQKxy1P5TMp6Jz11RJV+v0OxNKVDQeLZwHnG
NItuGUshYZVuDfgAdKYdPBw/RdltvaF15ca6aC295iYY0tbl7c7F4udM3Uc30/D/
89NhXhHHWArFapACzdR0TzaHzcgXrXLmLIqd1r3pJxi/D+s0z3eFQFlkXIAJ+uxk
grHGNpvOwdv2+Md6m6UurrCf1YLhpjHcvltbrN5hU5ZWIiQ3lmbPi01UZGB00HKZ
Zg1WnSMMeNDSDEVwUhAen9GMh0e64qc6fQcciRHSLJ7jcf86t7dwevsUadfF0Ud6
TALsNPBa7Fj41miuklI1tOoEcZryydD9igqy7ragseXcwNOdtHT5ko0FiuJivW6Z
WGB4FPikz2Q7duCgoLSIYAOQNKgOaYdnW1PdfyTyLU0pKNNLgUxkRzMNRthcjBrV
gdiNCPbDs0CKSLoJ7chVavusAZT9kSN8DqdHQhsUBQYWSNuccsaVQXXiCLoQX5tj
cZSl0Gbi8yb+YDLPFLEwMlmacyiF12pyYihL9aS6ynbO/9+7BsvllIpyXpu8TX8H
16YsS3FIcbpTKk0lrEU/HPS+gmt/LjvuWsMgziW2TxDSNTsYu5h6NcfxzJz2a8e2
YfIooX3IMQFcEClVq4SWBqvE3YQQRYoECKQwvO3jQOYQBQxwVfYzzerv+TMAA0ql
w0DVyeJe2jFAESNTysB1illEoR13hp8BcfXMf46FKW6cn4W0oVvobcflk9WRCzBX
5dYriQiqtlfRWENQb6FBIeVJRSeWtBFLC0pU6Sx9SkLCJavQwRsfJNtQ4/LfyCCI
x5Q2JcU4OVzCvlvQjmBDRcUZ2JdqLMA2Y/9rDu7xovvFnK4PZ5bb/wia/C7rh3yM
2eTtvq+2UVUyhrc6ZVE6vrh1eU3r4kMIIReVrFR7qSlQwx+dYlu26BUyB4IJ9z9S
mBcE+mrWIqhm+M46LYr5DOTMjY3HMwUIgBqvT3jvBi35Je4vdwU+45KDuMFWoGPh
6YhsFA3pIQl3rHoLAnCTVFAQ4KxneflEK05wSU99shUHlrt7eGY1wdvuK06HpKlk
sbZjh87bMZBY4foG4yVsM0DqNOO8BYLdMsFI0nSyG0DRyi7El+DOjLk8zOuaeNEO
po3gR7jd0juds9wKwd3wwJJxO5AegFyxSK0GuBeQUuoYlFuU4cdrRSBvACdegM6T
7KWiZdx+AYPlOjO0+2K3uNVFmIox5P2AAFRJxbLbnZIcJVrlsPTxmBmElYKZuuif
Jq0afHCdgZJMK7RcMxIi2p4CSDQKgOuEn4NowGMiUVEflAXWLigQp/V6jDATYi4z
wkOX/mTFx0W1zKjmcAgmd49U9LiSTDd+slsZS2cnZjZgCn+ja+AOBm59OzWitM0d
mWSiFyrav+YlNE9v9LZMxvCoWjSL3Qk2/upozqZawHfsGWpjyAvN9WrjepQ3A+Q6
0Nk5h6cT/kOaXrRhz3zkCfvzGam7czZwF1k6eUmO5XrDVGDIXTPo88wToWuV7e/u
fyZ+qqkCtZqHj62CiUHNnOpsCAe43E4zxudMw3azTgaGIGQFLKWzIVNTECmC/TwH
XyM6qXYS73hDnIG00dbxHnbqcC989K4HEmb95TZ1DTba4v2TEDXOVNiIWQcSd70r
DCimLejc1gjeBazwLlVEfit/iaIr8MVgfA1MUdkT8sBqFJhzuR2HND4ZhoPoAC6T
NoKUtwLDpAB+hw0bL8ZMuJCjUkdugoxUgfxd05s5lGeXywGL4gAylpICaTmyMmuM
42TXT67Y4nn+r02w2WaI2MXed0DY8pvmtqbYH/QRFGQqN1saBAbeDvrhq9DmSC/N
Hh6ZlMCppGKoF5qW7NcIe3pjmx5WT67CQmSl+ekRRsM+Fy+YevuX8WnaiuW2yDYS
HXkracv/sumgkeeqyTf5AL1I/B/p3bDFbemO06LkMKT+8TIC9sLoMSGnHTJ4zCT7
Sl0l6/8LGIWN7JhkfmHO7x+Qr/FMFLx7wp06dMs1zTUJ54G9Kc/ElecPU7DOEHYN
+ziJWcqFUw80mFr/T7VlGzXSBg1fk2yjBiSMg9d8kQLC60wO/mZ2WWqnbqhUjkVI
PlQi5JcEK6SzzLBSup2Vd+F4HGHXLDie1ZL2GCcWWJ7HK9VrxfIjhywYFaUsWQz7
bffRalMkhW5ddqUL4Ydgoyha43nFn30WwY6tlekiwI2+CZaHGgWsONv5WTCs4GAb
oRRe//Mmlh9IpikK3zH2am8VD2MqXIuRi8msvwinJozawiDmXynxh9SOisDJZKzs
wST23G2blUg1sc2DclfCnWiwdfeeNRXy/BwFTXFlC+5JnVN2guSqrZjX8Orun6NS
hgAO4+IwB9aItA7Sdj1uEihwSbDOvT8c/E1ZCa21Uq7O0Kxfm7dgWuz0qpIIBe7B
oOyYTPQ/zH2ebNSAH+rV6OxpdAUIkVaovHOeoz0uXgNYGnpEcpZUbpzDFG877bjf
/XiipQ6d8YHvK0tBgsk1ZXtI27j9x+Vgssoz1iY5e0bPJ+serrEglpYUv2xFVpkF
lIh+i656Zktf5TgSV7S94l8sXG6jMCM7b6I9m+u7Xti4UTRLE4t7QmJ91rNg6hmp
8xUAV38/USLpXOIhLC9PswBXEOffxJnXMKmTqPwzNef+suE4vW9G4FTk8Sjvo0Dq
e5UuDYqIFhfr/jz+tyK9/qmOcKIad5lcx+wvrkIacSSbMWlU6h9Tc+FtAhJEQqbA
1EsL+lk2r+p0pVmar+SM6KHblYC4vf0Q4c5s8pcFcOFN1XXRys8LMSjzACbzWR+I
lXcNGlGg+WhIg1XWL//RUO8SlbOL4YHd/NPfAJ1JA3HqseF6yzhxbJVzj6IFZfbU
0K09TSRtNGHOSVYtPQrrh0CClL9Y0cOpMfdywYGStvPPAffeEotVo5Zd9oZrHewb
PXRBTXGiUaFh5ZBBZQWmpsWLpYpPpXPUZVfSBoxTmtroHyTTcdIS3WG2Ou2wuXUZ
N+txZu97EmroKRnJoTvNuAiKgLBl/l1XL0Uv1EQ7ju9PCghixnCzcpOnkjGA4Pcw
xAMFYS+47uJfrKWPuPC9gV66DWCJjRblkmmwun/HBTPOyeEjPr3s0ICVyKnRilT3
mjbhyD3p0Y9HgnbJjw08DaGzYJr/98pboxACJDtINAoJ0zfJ3lhS04Ry4mvh8PlP
PjbqLoeLwlv1ztochKRIdFQXNwJwk7snBFsTOzIHio+64NkVeqLuJRp8OIqw86dH
29jbE8dTEhZ7XClsmNPbk2JIPhXunbQc0jkbWHRjzAPxN2dWBIi4WPfZUZJPZbIk
VjG86paWBZMaFCLOdacw3bYBNDFPXk+QWXX2T3Xg+OyXBLulcBRNQ0NUkgpA1szY
3HcGpbBpVvnh08+ZMISWe58oPi8rhyg1chQuc/Sgs6EvpYd62z6uZnxbxh6FVdSh
DCBM2sRxk9Ib9P7+at8xJYLkjxLPMtveIE9QVmcXWR39fc4TAWXuDRjbmeaCXz6p
RT6V+C2ZpuOOP0rBVHn7kXd9oEcXJefvNqgoQpWK110uOtWI6HGInTNRff6WU+qH
gJmWCuN72YumqqY+kUF0GPh7VJb8d+cVUmp0X6QNxRwcT6CuK9AjiP0Ue9u5Getc
S5LQfpiLrB7i5UAoOKwXLT3nmIFh6wGJUGoc/7+7sKb+//qD5sn0rn1g3FZKmOfP
Qa7nK33pMMzPM33z62sOQEADhzaW5HNgIBc1vtt2KCxb7sGwyIHyYsI4pYJ+iiYv
yRkRxrxObmR22gzCixvlYIppiHiZHy4PUpVx6tVjFkbzymJP6eOgw6fXh/TsC9lt
g8XF0ghIGwD7NYGKsiyyeHZbe3sCssQCiEBFgrIZbhyxIK/j0GlukD9EzabLRuf0
95M4DB+uyGKubjksPvvLOJBP1dMF7jqE/ZLOb0Tnr0gnKAtNhVXdUAvaCjDYykA7
0a22YOX90sM6VZuW7xH2+IGtuu44ma4gIkVJyFFsgTqkpDSv53FFRexi+Yk/guS8
qGMczodbbOj+W28gq6Ik/HyY9hbTJlS01/ITI0RuI1GZxGkefB3PXWMe8JIADBcc
zIBIIUMe/uoZM9pb25xmZV1sWudV9rxFwPGccSCObyhzvKigO8IQXlq8sPTHTl31
j0iSHpJYHqXkTHnHPGT0w4XVB9Jcy/Rx4I7m1nFVmcJw8WJUy+WSXIDlcGH0IA6O
HOpib9VnSr4dYq+BE/5bMPRKwiNC+enxamq9r7fWALd8GM6sAJUaW5XMtRAJou6S
PuBcOCMmT3Mms213BaMIUyhOVXqxZnPQF5JJNkFadctpndsntnGA0OYnfIMD5P/6
k6eecCT5MCyR09Pdgakfr3crXEp5/i70pHJ0sS+5rAZpj9KbXH7/cqfTDp0Dvmgj
3dxSpTO8LrkveJqsrsfnlHVAseRX4nk0Adrqx9SSLmbDaX9zIgr6DOQsyNY8JHg/
I7zIAiFdJNed9O2Vsm80CY19xr9vu5yAbc8zzyc6zSoIwXL59enPCNHxFcwoef7U
YLd01VFzz1/OvqimuvePeHlz+CJAyOYucn4FP3eNA7ZUVwJXf7VFumUxAC3qUviu
towKCBmLo9X6SGB1cbcc30usyuM1kBplLvuGCJ4b4RnDNS0OABeV+MQsfspJ+S2C
bSfGMPLP0+iUYEJysbhUi/+OatEw+wlc0OuXa8mkQVz5NVbRRvmlI7T/V+8IiajP
FO9ryPluYb6Y2UrmT/WJUWRsTf66a0A1OxIEs8aJxWaV1t3fZg8nM/8+wxVvsxbk
uQadFKiFKQxDHMqu5g81n5GfD9c2vY3SIN1cxuernpTb3cLi3ttyiiP0gwjhjOod
dMTLjkdUgXmxNnaD/kdrACWoAzKD9DGLrFb1waYFYhtr32CNajQHOR85naYlJCjk
G9537kks54QBrVjnruSpE0osbqK/AzmYujoew/LQ+CuBYDgKcor/S6gWRLbW9qgx
BiPlCEqtF3Zd7etd1LhvvyRwN/c6Y80LUzfnR+fhUvSQywFZue5v1zW+/BF9CnSc
5CZ9pgmPb3WicLFyWeM/Zrymya70rq0Gte/N4E0UuzcGmrhzddsxNTVqrfMy5rao
rTEuYTc77PxEVOGTLwE28VISsVohcK50PI/h6LmdcoX9Jw1izzVcVFnAofmfNar9
bcwlZ8SaQKaVDqVcBMiBjRHosoQqw3UkZp5Xvv015eocndjxq4jrey3zaVy6h2EM
r6wrHz4vE2uLdt4Kc6ee/2ivj/ZWtD6iQfh+qIBxHq90n+HlcHOOkJgiAXty2eKz
jLeLv4LNGG4APpSAyDKW4PM6FKDvSxyNwK1aZXktXTDXP0NNJQhqWyV/lM0WDYJN
jpe+LwqgcR8ZECsI8kMPunqCuZxg4ttmy8dUuaBLcVvN/6EV5n0TOvgy9I97DOih
6HUGquoZK0N0FVW2DzchbWDsfV7TrRMns63NayXwLF0Ff5WtGBAWxtaROeGctN14
ktV9TiY0Uqtpj441VVikRtzLjgQFGO52WXUJKRmcptktAmTwQXGg9RhkG9CrQdXA
hiPuQBJkjAClVnrLqxcpeGBGg6n1g0qUeBea/RvUEgw4WGTRoz6eJUpgU1lIbe9s
rpYqiSaR2j+ys+KoIxmMsu4WtsmA8b1jxCpfAeQXfUYFj1aI/3FaV3EMa0M28T74
J7LKT+owHmt8wzJwAmIL42hKF7rlUlclf2BA7p2kdeBZfLb0gkjkV6tsggUgRvXj
hXRZVFhMC9Wtzta0OE13vCTqbsIVXy8T0uYGJYFzCtut46OGnkT4+MzbT5UCulNr
zC5Ot++N8NRdHvBamEhiwhZfAdeMPN9O32icWUIlzbJ0OHCciJWGNN3DQobkqzo/
9/lxtigMJHfiRMAiyNI6XRmlUqqP0he5UNdVMVvbfXfWaCcNJDRM/eciVhoFrQ55
MvUlUzgM06tMZ4cItJVcEMXf9uRDNKkXN1LEhaCQoDnw2iSQjKTIz0rGBDd2sUKL
5gdD0059ZmPeZcIK+XhQzgZFbKjlNSRrjLz4k91u4GS+QQpctFsp6JpUxWySq8e/
w+Bk/4MuopM+QfCN8+qC//pdaPhHxWHlEug3N1KLQHV8W2TGWJGWPOm5P2z94aGx
ZllBJVwuXNtbpx03L81mw1bKF306M5YtxHLNrF8472mZgQTyyUrGHGA9e7yP8K6z
1H433xI/42ir8NeQ4YyV9OtEkftyJsVnNMh2NaM08tCPRU0B2sPmHeuFYttSsu2F
6akkpVMaefYIU6Jgm7ITdQN054afviEvScRgDgNOfJMdENduQJ5buN+cDQ4Za59a
mYRmkEDJGIWBIIiugvVksWix0YtG4WB8mWdvQJPSrVGTz81Tirxy7+fL4RugIfLi
NE++or2FjeBJgQhoQIIq1qCL4voBxz6c5aRazYho81IPhErjFAHCjeLX+520xpOv
quoj1YM3hIBcsHHNOH4Ozw32pwXP4h1oV6OZY7fiAP/aGa+XFtY1i9zLokKzD4HV
1UU5aYNACcLzja4lW3AhFvAID42h0lRMJsa3iynXvCU1T1naznJsyT7ib0FZIcUv
izpyIkwiT7pImsmuD8Co39262N4DGzPcZsnLNP3mM1++6ZJl62eYOoO/LmF2FeXV
JId8cCnfXimIaagWPWpkTGKHHH1ETZrxIhB9usgX9c4zKU6ltqo2QI+xg1lidcdt
EJYPXY7MH23kw/ekgSi7AAVTkOt4lenxZ5q6f9hHlZMRJQA2+BRvOMv/PtYPrxTG
iefP9y6Q+EvqqhCZU5S2Gi0rImrU4Y/ydXiUNcPKLNR7QvXjYbCBSYhHJ9VBxLlx
8R+9JEGven/D1DlLo0XOFqW1UXJYxdLRNSIJ3t78mY82DHILwcGHZSbSZxD6Hi/L
ivIePiuwrokjqlgqjPyKZZMv927spggQpwJFWCyu6RwXZR13IKYLMjnMDYRwU6Ul
HWzA3EsoBZwDyU4xM+0YihYbDnkIZu2Q7qHErsWU4shh+EZCiRZS6f64bqOzIWFs
k6M8rEFJ5YPdWohM+hZQgb0I7kQ8ZkHVw+w5wFDRtDjwdeYc53iAsZXXX3LCRaKh
JYIhzhqu3zhAvwpYMdgHlDsOg/WjGRTJKd8TxGa8+Ii+ixsG3cUR63IPrKnXeo5W
HCaI3laFdbDOEmXe26SkALqKFILkTkIqefiVx6hc6vxO9g9NLX2mbzOa17D59SGf
PIUhm2jfRc1MzNvYaOmCgClW7GK2VX75sm9J8gS7ilDPrrfTJ/ZWnj2xw0KdAuG6
6+k2WvxF2XEKMwpCkCdkJV1MJtZv3p9J0z+2L9q6Z9onfQHG6t1qufOYhrBPZ82a
V74DYwzc2OWB0TG2MMQ4Ehq3WIk6ihMnvn/KCnnGIVyGZNd5BbVxsYVLwhbzCG/8
ZPypLB8Jcd1hflBWtnVEkgxtGUluuNN/ABVxWtNAXbHHzSufOn3eSxsipXPG2G/8
oUFlllZVUQS6tR/ASU48hHlg+qU8yBJgm4PTdWrAno3M+UGpuBoOFYWaKXvIkMrm
wh1nskMpLZ3/aDuPnQi7LvQAFQLgqhGt0UvsEyxKgFzNDR6++D6sLwmPCIZ9QFBJ
rGNhv41haBS+A8Dvz8neDIfdmVu/IXlg5UUoKlzBrOV77TzDNA+/BgiLdW576DG/
m2IyQa8p+H9yXsfP3GtabQ0+bJxBpDIgTZbX1I4N+sJLUW7kh4sCPmVqRxsumuFk
K9NBUZ0B03m0xSP3+wB9yyZwYcBHt5632yCGIwCy6qDM+vVHxOqhqDClESnz3e8a
0D79V8ccKMsjkEZR1g8WnpPhbALs+VkkHRtWn6AhXYFUZPEOPOqiEBc3K1ovrXM0
z8Yh1egBfVdC5biOJ+Qx7iAckzftOT6BC63c4HVyU15Owk2RVoUslQnts3lQRR+Y
jS4RjeEW3FsRdoqLf/dBf/B2AxXNNJ55RYaxBAAQrs9p5xW0zk2ODsLpYMEZk6AV
6G4XuHNEkJL1PVDhyUJfFWstIplPq5PBXbmSLg1MFliSY9j5enTdo28uBUbR9/Yq
c+tYjVY3J1UFFIEs6cLZl+im4PCUsowB7qQKxPtzvLjTn8voY5yBbC6UrYcaoaxW
wuCx4nWm9V9qOGKKVfuCWabh/spjZKj2RWMiDvdjsWJivBbDsKjWAqMf5+lpgzR3
vkSRSlEfzjCPkfkGvBWgm6PMpJvgIDaQR3E8AQDHux1YKf4f6sz8yZJRNjOpgiEu
AL7jSfJBYEMMZfyaXNDNEoiuS1V/lo8rOE6/9WAqsCNBWpXhKgMtcSQMUJILR8cN
iKN6TEe18DM/CGDRgm948MhRofnwLR41Z4jglmEDaKzwVnLVJ6aVILGJhFE1EAvZ
PYxTgXY7wXvM0vuqwtvywcr5QPISzrNHraflpJnwlrAPQ1vzi5CwHrTbohYlGccF
pDV9IBU2PInf8WUnHa0Yh0atRS/OFPm/ZICwEgB72nzn9s+Ml9mN/WnlFQCUvCtb
brU8Lt+yUWB16k8aSabRKdJkvUMpYUpO2dKY3PdVrEZLH0SQMYjmGoZl37+fl3/D
U+9X60Jh/tHTe0VTQHSbWSVw/jJ+jexARZ/Xjr7VC3BjclkAbQFQsHH8+8ggMKBP
m7ejLqLCI0zhM1BKA+YAdUONQs/vmLvOJ6PiCYOsGUgul7CWgBwLw4ff1ruqY1+c
OV7KcK40zegAhrtu1KY5flfl2IR4Qev3bvYkX5TpU4ecfn9KMfSnovN46R+I719D
OduQAH5EScDQLp9FDCvEIXlS/QFwNT/6mtNhHjd+8tzNYLgrAUi8EzO+Rw/Yfnml
52MAO85Sq1vn1AYvtzQPHSEj6z+PZCSJvojMsj8DTtdLG0QtmF2y6XNc0KvC6SA2
ZB27LMoIBEWfRQcMof/+2YQm/VaGlnPl4o/2dOYDWo1wbokfX/w52sBtK7jqwQhq
HF8DsbUS/MjxiACF8s7/RLbNf7RYKhHq/a8BGQYSlax9hWPjOLhQaY/ks9EP6p5o
HwSdmJ4MFFqUSaqTzYQ/OMSLNTYcC1OJhaGr1BlO4W41H4Yv1mqJj6OE/TnXYSKh
dxgi8mRZuP/MmkKFgumjBjCVEMya2czVK9qPI+8HaTgKaTdplOcLU8g6fXOejyS6
aPhFrMUp8mWhFJ4euB2gswHILj5p4PWx186VFkPO8pKBvpa9d0dYt/TyUDwJG9SG
g3Lw3fFrQ+X/sKQF0EoJ6kPZFtdFsCkFBF/8veZjDcXQcsuIN3Ow9nkB5dSjNuI/
Jjbvbs6ae3OKVtMKcm8m/j0ISGzX90X/hUTttYriiLX2oDdek8Jt0LVr6SCaJsiQ
woUYqLku6m8CZTUOPIvml8kNZFSRXvEtIdZAd2Yumv0uIkCmV48RsEdoRVdB9CjF
tMB3RJ0c34dylfIAZzAQbpAGOOIiSTlJyNVidciO02R4rzeXMNW++bumRVrSs91c
DqIZje430qj2Vx/auDvYwQhoQwgjXGkMClF4QXiBKmiudEfY/HG5z0k+2nbnYCQa
+vdvfHfSxCxA7KLVA/D1hgFdm4UNXydWgFdxd3zhofRcWcOk2yPwi3q7tW9iwzlm
Z9l1LcMh/eLHv9dv7sEqqDt6nuEkqEt+0dDuGs9c/dOYuMBtFnLUH1Owpvd0iyG+
WJKcpeX66QOu+TMGH8ZRKtOEIwD7137FjJRfK34YsfXwoZMk1rZHNm333mlZnX+i
7rkKTovFJsXv9LscMz81waInuZ85Bsq/HEJOUpJnpp2vPLo842Xhwb2jq4WrEuzo
MJkuQgVCPLEfqz23uwM7HusoGtyOF183Cdy8dwbppGWvTHXH1wR6m59vKLxLHuwf
/kVaqZf4gf+HyRUpbMYzTnBTQiMUC5h/zPc7/M4BJKfqFgms2g3+IFDi5AE/8doU
zb9sTH6zN8OpYtFmjPTLx7RupQch1TPrSstBGAPPXyYQ+FY9hkdDxmMxuSE+KLXe
rPg5chn/fRM7YNXM8y64vc/SlVRYPi436m1Exmq7FEAFYkzST0kn70vHcNOSiNSg
A1e7u4yf8O+gbA4V+CHuLPu12Dhc78qVl5I/eqUgxyF3qwllLfd2godVcm2S6Yrk
nkGchM0RNLIdILZJ4wGZcIwMtgUu7eFmr007zbnr6mzJs9A/zP3wCr9Vf08rgFKR
5diNm1Ifm7/BpcZcgKrFRWMVBNZ0s5C/3uf1QvRHKHG4N3pRRDP2wepI4kEUdwbV
0zRb9WIIN01VvrLvjF19hm2KDYTuxTq/pCEgPs9/mFra8aB84MCtNMRwmIFiWKJs
MY2mjFitRJUXP2S5aIGlbgSfQ4/j2ylP29yM+vizeb86rdCHFHHvu8cRvUbDdgh3
KGMDD0V5YxeqJeyJYsEG2YUVsFkmR1wrG1P+UgKpUhqhXSbRHDk1L6OZOgHk/xa+
56DoufYTXmx/QhCCF1cTnTUYH0eKYx4NIDLKt2kgC8vqwVPHZQYmYxgw50l7YZtH
esbQScVx0NPp+1nqHLyW2lCue7CD7Ya7HeK6uwb5ze/pS4n6Doonw4fynDEz1Lgr
oDHTAmhg8Wiu1j/VBAnm7/eDHGDatUsPQfsg0rVNXP3bbvbXwdv+9V35XfbD28I0
Uijt+Sm6AhGB2XgqeH5uVRlPifVcb91xNAAEIXtk9G70O4MFDFprPYu7AMXWebDn
usf9ccvh5kTP7nqAnTsxIDXYTqG6CBgyCaDaxvSy0oLezQP6OI9z+kGMREvWKeJF
n+q90vfwdcwJ2iNPGSa1+ph3akx4LPpa7mC8b9FWDzzhe5HDvoPQPY03bPQPJN4c
n8ubL+HIs3Bhvledx8M7rJrbYLYmR8Zi5eKnhyk4xr5bk84/uMwnGQuKrb/TJVGz
3JeJeENz1gotX7UCqhAwz9wV6R8A7rTNUSI6cbw8+Ff6qxRWhriJ3fEd8SohJXqv
9KZaWVlS8mPmZv/iAT8ZPnJnwGaLlkYGaR5Uk0Ku5zChTc0OKiXtSymla/Nq1sFg
oYlrfLR36o9MPXB5DqVxr+9K0sDcW4+kS/u8NXv+n5ro8ae/ta4kuVvu6iZBSEyC
4xAaIdWsnrGlSPhzJDxGDd5khCjCCCSkyfRM6ekWhhD7N3tF4Hqq1gy/aDk0oZre
po4SKSCEOYsbKsT5KwUYEBTF9pO+XS3YWNYmlRpoNpgYZSu82qlXvm4EINy02wqI
wk9c0Z40roK16VzJhwNO1y17UTwA1Q+QP0wCcpuW/kNSkZ+wkKjCTL0DSRUxqcRK
t4s7Yq5ckz2ELefZrK7k/DcWlGfY/NipI+GmF3qCrLzPfayEIjYpKxXEjcOQEbQl
lzTQUDAj3TkkDDCvgiwysDKC9uUGTCUfAKx73zPydM9ujnxFO2y4Shrfb09j9cvs
Hhzkxep/RlQqBYZBJhRENR9LHiXaeQXcQKxjOmpr0Sk6amRZwjOabyr7rqDS7OkZ
M+yUtCKUHguGewzxd6qjLI/6AJ3HGDeGJo1kmo40aqI0i/FuVGpsMJWNB1IS2cvP
n4jsWIq6hMFqEyqS1VJmtnzUgA60AHOoahdLyeZL5bhcUdZ6PWJkUfqkerhLk5jy
dVfI2AoGER3A0if501qfWlYtMu3iUoC7Gt7gh4c3vqARoJeg8tVsjLB2NORn400H
7sAVrd1ZL5u72+0gNHRDhHCFu/KusBzXSQFZ/SAky7V+qxW/ziyN+PDZl6bPPD/K
YUyjVZqPm4UjIie5AE3evsGcPuFIjQ63ei27wjIwOW/iuSRNxfTD+l7wLS3AsajV
SaF80ODByI4g4bCQypsdPEXtdVt75+9G3B76PEUOmjClBsVae2Irv1tto5LWvTOA
SQIfKQYeH1wI64coWSmfNIwTPzazRS7h+yBuBRAiayyhIDrPst5pWorqoEiO3btb
ibfwYYWcJ7wI4v2zfcylMP+zlbK7ixIvzZWps3wmf/lfNelIAiysSkcrzevk3A5X
sdLclmE8x9jTJG++9Q/xcJA126K6jk5VgwrU9pc7ZNljW1hbi7TEY/ymw0FHsWWz
NVcYvxzRj0MUJ5/tocvPOidW+NmpW/uwFbSiza9UyBc2Drqr78/Crjhc6kmCPiTF
93GLBrRcRcsf9fiB0n+RKLhdKg779GlUpBZCRWHtpAHB9AQISW6wS7ngGtL1RCb4
1ZEdlvFmtYWx326il8hsLAfnkzbi0j3y+sZOfnRxSYTcrA3iBhCQ2QjIgVyLQbPh
MQWKxB6Oib2UG9GU3JeO3SnBZ+mEAJLhvpB56e6j0hqEXbUR7FeeeK23KiqgY519
Swy6eg/bqQPT1hrIOlDnabD6zOLfjBh9u0end+y5pSpyiBmvQY0c4TObMSchZ/IR
yOWEIySuMgfvqkq2Ql3+aOa+ffQJnIzeCp8i2Kn7yLLBsGUwBbH5f3GKPjDIZrWE
TguMl8oCNq90zzM/5PmfGH/XMICScFebRiV00dMFI9QwFW69elXgwiVxz/2Evo6l
bWPrlc3rtJQ5q/lOhWt4mLM5IHHmzKlDvd+D4dH12IYx8OF37fefr2JOybtrWYcC
uWF9FIoTpjrv5C7TzpVs083emwMjvBahg3alCIzhAR0MRM1sJHfbgQtGF9Ykh9wk
Ogw5uklu3bZWtCVseNzQHrXx3Xm3Lboblfw/RaIKx2uP3g7XqtnEIrd46bSMPt9B
HsCva3FXO/aArAXNnVXhtKkLjABR8Cifx0No7XaBa2WJDcTUGAaIHuXRqNu0Q3vp
m3dkmQfsH41TZH2zOyCQ4dROMBT5DTtfdKGumCQaJjFa7qcDNelSAjv123GnyHXQ
mtnBpExPpb3erA+xMKoFWC0ZWGMPTQps951ITBOHHu1+C4qt/+u6ezZzQD9ky5BN
OKHzSS4gmt4EeDzryfkdJZtU03ZuP17zguxletnbf2s3JTXmMswpTqBd0uoXtqJA
ZxszmbMqDDfBewAy2Rhu8V1j7aGzALFqm+ENyyJD4NHl99dZ284PJPfiT/o/ymSs
nbTsC3A9wgCRgQlczpVoJ6gX+f/WFQztzTczGvo0quuGuU25/5Iu+CTsGPFnSRdR
kR8UU1WdPV39HKTmDFTxRFfug6VQ3nX1OaxgwVviK7tarFlXiw+aAUy/9oQfGQM5
JrxmjnnFdUzqvJaGLbfTKknTt/62JW/62ZjsNZl/xFh9bumG0IFn3XPqM/SXs1Dw
l/EmhZK3FRSvmp4rfIYkVPdcSpPe+kw+nQzxLj8fl2mik3RO2yaqCiwNW1Qqzzna
jtVktkcRWEnuFXnIcTOs3BuOZZpOypNtqE5utv2gn0lfnbFBk9sP8cBvLjjWfudr
igHerODNSC314Lz0BJVWi5tLskrFJlSJchJXLjvWNhee4VdfDmrusOyFpBKjzMtk
sUJ03rxtVf9lS7tB3jSE7PPkvIqjJfSRIpPtlcLN8W+Z3MMQnhxWxRXGGYo8B8II
7zSgVOBWUpUZ/nqltj5UA1FwVfG3Y5PIavf7YmTZzAbBRyN3D08AlFvFDV32+wPF
4P68p0mX0yW8v0t1kyGkVbjzGmcjgtJzIVRuGMFqzH1LtPmUT8fgMq+hmewMVeHk
SfkhLUQLcOffmIcBnPXPeS0DdK6XhTcQl69nPEKg38US8QoG5obdq1z57aUkdH7B
zfWuJ2uy+7MY+ZAU1c4jghKjx3tGCPmWuGpY+Xp7+22eF2baMhGj0NhSXJyeXDmA
9niEhgyCWL36fyCntAXxcDPGwGpi6FmEzBgpnH9tHn540ZfhYPn0rN/Vfi+fH0rA
+bjH+m1So0nuMC7vj5viloHx0C8htpR0Nbc89Y8h4F09STmHE+r3UsdKT6m7ObT4
VKJ8X8EHd2KOCFk5UG5W2V4PlcmzncnwC+oMy6DQ89r211YQ4oI9N+/c9/ci7sL/
Yh7I6vcmgosASPs6HX3xfD4JKh7ZsaTj5YujuO/e1e/Zc7wJa+KckARjX44T/KIz
fxL3S7Qveo/VI+WxmqQ506GggDxVCyKcRptMJiuL7LUrK3IVIVY0pnKpQZgayXMj
A1pTYD9vC9MK5Z8xeJYqfi1AomaWsd5XieVwRWH+110Eo5jMZiXr5IMB9QORrJx0
tr6j6m6hRPWnAo2zEBrzsArFUhPYs/c19NN4+M2NxZYocU9+gZIzN0ZfFDhXwTD+
i7vPNLVPZAjHzyg/E/Bvmz/NqCj45JQ8l/e1PjHHPNuA6Io8t/AYjMPxeGmFD0tL
d2iWaWBCkr9WV7+R/Kd+zySOfL7yX/0nTrM/5/p4cXoEYKWIIj/G90fu1lECrkZh
UzjWwdUKKcVI8pg0HgI6bwzdy70HiZaTePH0tFuT0/HHGMS0ximi/7iIwAVUKa/T
xy3a5Q/uqftn3DtcXBMrUFbW1sVma7Gn1VaYy1WAiwhITh1RHG1kUnag1pN8FcI3
2SXeI94D9oOL56G4/lHtQBjXXJPqqYaJbcv5N/3pye8Md7ZV38+JF49g15j19HWN
jGAk8v62ylppcmP4UKFdwWRiv81sqdR4Py+q9RgW+aUey5S2z8LmRSNnFlsmSt6/
PL2+jjON5TwVUAMmGzSLKtvvRwR6blrg8EP6PcTOHmBuBDCDuV/pfNpi+D+S7koY
Gog7eSMhTPue2i8t+sd+Dwj6KlfTS7ZinpMEOnIvhK7Me5ujwMI0jPPavve9CQ2f
IJxCPlmpgFFY1t2S/Y1YH4nLs4GZw8nk3XQZ/lXIvCicxZz/M+6q7aEQp1WWpPQJ
H4SgmGb+MSmmftZfOYxafDRQ7OFdSG0Met/nwJV5yAe12uU5bSZIziXkbjXTK0zZ
zjOJ+W1E52zzIEtFGZOTbNRzjuS5Zn9r0/6BWS8WxP+legy4PtnQaUESasDO6emn
g/hruafj65UiB0lelEBqv+SI65+eC8s4fcjAzMidlAwWDMgjAP099QaPoRlq2XK7
bFGV6qhC85GD3RqBiQqMXvSsbnj1q0TQFR8AyBnERfr0fCpce2vsUy9hFYRjG3ym
Pf/m++tewDWCA7uPGMLoq4kT/FYuGYSD8Ap3mauDKkwU7FjfRTutmOfx4ZNfoZgP
vtUZ0t4F/LtNyvWhBWhlLskqHdcHk6jcTOMLEe1mBVkT7zwLm/FqHxWAUBRuJnv5
+0ro3+Yh+gQCmc9LWK85yeFY+jWdNXUMS2sYrlK/PINjSUQAFxe36cEDhRPWVSAR
+3sNmZGwiaZy+H9Hcgj1ShH0mXp3K2vLGw4iJ/o/AHE+nffiCeS8a1Wv0BSkH+tx
jdD1ZpQsxWiquCzMnrSnd2Tw0E/7eUPgTolIcgdVuzhdGlTAV3PPPHUbLcQGD2wn
pZlhp8bmg+C9YxH92G0+uxnl0RRsiyIka1iX524lJtwCmVnel/PAjs8y4LwWPqyC
q2ZkewU7UoFudM+cT57mXvOHfW+GgiVcxsEqAHz0riok5LUqZsoez1YnJ7ORcFnx
hFJ0r0KRJ6/LgTGYOOcOVye4LBUwg3R3nRr3mz89Ov9HrckpQHTV/4ok0E57h4Xs
RAd7mk4hvnd4hX8OPe4aon8coG2ARLEfLWaaMfw7TjoyMH9gWij+ZsWZfJvUxZe6
tX+k7iyuhiFL6XEsE3rJqNP45QRF1O8szWXRGa/krb5mNVpP57rV5XQ/nOFnUZim
h3g91tSo/BPkyzgdXwjpz+JxHZgIC6akFR0Uh6IXEEJSMZzvm66XKFN/wPeKA0Di
swb3bHfurdia+6dWPOdfP1U7hBW1yZMzSguA5+KlFtaQ+aIQWWARnNEyI3YIcKFJ
6J3H7rjupUiezKFW9Ekd+zswuSqR65s7WN4WLOnqFnwt3mq/vTi3STZnh3axani3
qGJt5tuiv90DwUy5DtUljdkDWsEcqHFdXEgFBbfUiHD+a6x/Y5XxmKlXtbd5cbth
bOZbduJbRyMQunf62fK/M5ARROisMKhncTIcOh9s02T/TeQh92y2nWPYxT0EvuL0
PlLkk9z8HwuWZ+sXZ9v7q6W9H827TJwsndgBzASdFAPAtXO4cL4XuDThhyeZarbW
4W+KNI/Zv5lDK+1JP4B8gfXXTIwFf5KMQK09nNokLnDk1q41Vipw3wye9mo8y+nH
52bx4ywEbT5ETgOl78cHnVFLjlu6xJhPql6Rvtkn4MjrUhQyiBOApd/dkYOS3Yvs
Lbx1vQDE7ikBuqfL4Tzted5ZumFPwvEQCPDEKonkVnxlFjUBil21SuKCLD6wW/l9
ziz7OESoIgFKqdCMZTdugkDXCC8A/O7LEcodBN0YJFp4j9jb1Mrn4ZviwCZ8B2hO
8g4MgJFBCOLTAsRRnpJVWm6XuybYsbNyUiEEet+WlsVEIzcX8+K9znCnVYuUVBJf
arIBrr31/noB0qFSZV/XXIC+W4mjLPt80O7VmghVnZ8dcsx7mKrzlKbBkHDV7+IT
WiNxvNAHE2kYVzzeDQgs5ax4MasHWZzHclhU9k/Xi3uvkWENevwjSRny9cSebzgf
kFg8pIkh37D4b6RHu7+JrbmcXpEVAlxUkIs7nXjHK1WIALC/GpNLA5SpJG8W/F04
XK3Ycnzz+kr0HpsvLXJpBfUkAOiZQIAvWzWrfyQMOk7t1uqvwQNIU89jBHuVVsCb
ygcJ987YqzF2a+d8AHFmD405YEEEWifpm1KKiER6q+H4cAWHFpkWzDjB4QWOCIQk
y37aUMFNxScC6/47N/+b8cfHSekhfpM9qdJeCCz2xIkLB/uVHzoKW4JIy3bm/ozA
Syc6HnD5czpnfRBJUHN7w758Wx+xnJ/YbHMF1nZX49NryHBx8wlSXbXlkgGKv6+g
o/IfFU8GFouXNU36DQnvvJxBxbA+TG39vlHFtQgXZA1jFVZaUvAobqNI72Boh1if
9XTcGSR1RfYyKDMezauW8lnX1k292QOw9KfToNWavcH0fOYZxWKmYcq/76XAro7o
R3TOQ2FV74fP+uouf67ieXsTkhe+JIKyCe20J7PBY+ncdINfq+yirjI0tPOD12v6
p7MWjyYkDl5jozWekkuJ5LeuXxbTR3eXjJNHYVrjGHKDkfyrOdMPcHxJKasy00FZ
hPw50yU4C8HMIhcZSWG3Qcib9ho+7bBusNxFN1tGhn2qIsPKFoXb/xBmtMErBhQV
sFodP64goVzP06J8pNw0DaXjr82uKuJRMh5IP1mEm7EpRasZVT+7tGv7mCHMEGeN
+no758oo8prBU3t8/fXybkenlf7fapBwNRcGzs1SUBJZJlhHToPmigKXO4X+oUCP
upvLET8+3ugJj2LfaqDE5JeITDWstUf/l9ZRIPI/rP3WG71RLRXl0fg9GQG/K2CV
IjcENy48Ys1y/ZdLxlYA0Emyx2M0SVLb6DHyf7bBMFyfyhjlG7uopfTjnlZHy6Dr
EiuCIF5UAXHQaPnYY73u9Z+rzQn7qOMpwYhDXVxsasDW9obrPTBo47CH1xylNba+
1a+pUfV4HX/kapAQKDio3NnnamuiNF/9GGBx2QZTvjJm+5/LB8SS538bjDQKWbnC
br4gE2j4WPK8Br5UAKzJz3puEDJFde1PlOM8Nki5DD30EWphF0ZEiamnf5sUb69I
8RM07ZSI3N9VuLyOY82P4+Ew+UwhrqojZPyuFYN+d8ktZ2yRJ4TK/JEkvP+vT5jx
wsYody4oK4O2TdshVzaqhTGWO4c0eWhF/B+PzWsj/KkG3y289Pw5azZAZBnfvefy
2eZXirkPkQysdCyhRuaZJfkAVgASPWLEiwIJkfKCj0GcgxsH98/hawoH/keudAgC
ClLjPLtBiDRutGovpm8QM8O123jXXKOo0JvBrRD4kJOPfGKzx3o1sa4FhyF7Q88y
bKqphd8V8lLwvagHPzYomSA3NofazT9GcqSfqrMeYTO6sr7QzFU27ZiNdJAGeNiP
yZ+N/fCmitWnnOwCQ3TTK5804Yi3ORFG7/hMmjbGwsDrElswTyECXqzSHvSU/aeu
k6WYY8Q/MELmkzfmqOPgCAPrvzxdzdaW52gJVam+Lnj2edx9YBLzIXL3TfEUJUjM
hOXYstnT1EiYgSTlaxe1GAND6fPbI/4aSjMhS44iF1cRT/WsJhvYS75rCkD+rGFP
Jwzyp7pRfJYBMAONkhbIWIbJMcSQlH7n8rv6qyg9pWWx7b3C4QF5ROmB6T5iMAkb
wUyjpCMXQEUW5FQn9erz82vKWQ4TdzPjaFwFJza3RL+r0AsTyNC2YzUVPWZ71+/6
epb8HkZfR1eCJhNKA0GMFmMvL1R8yEETnxhAzI8KpCXgnSaWpI19tNgWZ6ShM66T
NB2gOcBGClU8efNtqLHTgWcnGAmAx2vOvc8Oxj7Cl+g9XnHs2qPuSzvqNMUtNID0
fW2N5ZupgK8bssaFsLHI7B8WpQFuf+UDred2aLbjDii+AJKkwg6TMtISADEo7EEk
UL6zHq2VxuOZjkx/TaUvBcyMOUGSGmE5LwCdju7QrVuk52GT//8+jQmfDmyv/I7x
rmKuTbOlw6tuavlC9fo+b+Hz8abBhn7y8CpB+7PecNljQqzJnDnpqIbIWG65eQ7v
wgAWrCTlIA8IimhIDCe7sGu1h4fCaqyKDPqtdxKYFNwe2aZze6IHYkpN7hbxFgp4
LKC1O8YeHGoeA3hS5/zopRTNzx2IEVEwzVHZyGAEWF0BPv9HYufcwSYH22KxlGxQ
lz/Xcst1RwhQfBygH1TaA6G0MYteUaMH8k+SBObff/WMFddw/aBEAYh/mmvsVYl9
vdz5sH61aaDtRni5ZeEjtSIAKCohY4s9QzVudQ6x8gpaRx1CUqLVgjzeNnq95+ur
9+nSNxMFP6APoVL60ZLUtrahcOAXaNapGmKtWn3OkcikwPsO1J7atSvvscMTw4d1
trKxFUA2P6SULL2cOdMNqirfDGhdtdI6j4ehB8JDK/FaLHA3LVoEqSfz5ZLf07J7
dmb0vAASulq3Z8mV8D8ztK+d+RAMdd05XHh7/3luoSPqoLAf7Yd/mPKg/Z5+fwJJ
cuwWKQLstINzkTuNjTfExJZlUz8ax6VIwLtvycW1BRnouYQxhOZ8sta1/yfJrTW2
trGauRacHebWwFUk9Lw2ij4q4K24GVlqiMGlQLCJvnzTukI6GmZA+5/c1Oo/awZ1
pZTO84XAhYuaYSeIqbcHue7i5m5t7pLEfzluDEnMGQFb2uYxGfigMXSwkKXyanKu
DUaYUer9ANB1PPbXXQakiYQ6fsUHwGSQxesjFs6FVW7+e43zSGIQUkeO6mH2HrUd
OeIELDybRh1zOf41OkZCMrC19JSQKr83JGuWVFcSlwohMtEsiwvv2GBgEFNqcajm
W390LKSE4Yu73X+YJseEzDsBUWE5n8EPAFwmb+/cTPFC0dDfBM3Jq5XqB0FYECET
mTHNo2dsdu9NlHw8Nj/SzpX+YXhagTuoBLJFhJ4hvu+ifT2LMj4cSy2mzpz2wJjW
Bvd27ew/vYAjw1czzkwsh44e1GvuriAHwoJbzY+xGJ525kFc7qc7955vauN3lhFO
ukgLxXBjscbRpEhpCjYk9bd/RrE/x5ulpxY9RJpoHUDBGQAxiEEHrZ2V6nCqZy5j
I/XCj7tf72H+wyo0Y+iorPx6x5SW2TZy3Vev0PlphE31kjAS7WHa/en07+cSm5a4
+dG0iI4maAnkLcA+hgezu8YXbDOITKow2EQjFlBXD6fQlJ+ySt1I9gJz59NwQHFp
y6vcp78rT05tTQmNLpWcl+huNFRtGhlMo+rDys8VbBgSJERws22dlersZYSvC+34
Bf3l50s2+hnjA0ABSZAkhTPbiDsKCfpVnANNxLCmU8JwsDRxlynE7UJhfVIl1s5G
+tOIKci/JbjeX4v3TTXYmMobiFqmDsqztig4QiRLpxLyekyUvZINgDWl0T4517bL
y915IcfOhbYXuil8QyFPhKU25yJB/H3/uiwMukM9bmRN9wTavsKVZXCkfQjkAv7G
q4UKUydgfwelLAfJK2wRLAIfu91MHsnb2LrLSFi8aUKgZXmrxxPpu0NCZvS5qb5x
JuWm94WfWGnOrfteq+xTdfs79GD6mfVJqpEmS+4JcxK4/kvzbh+k1v+6bgLTkwIx
557vqj+DNJEy6rS29hlLg1RphKlNQKOefnrHcbjI2sqRExtF6G9HOK2R/kH3IP2z
/DDoLMaglYTuNaR19pYyEYUwo4sn93qQ7M8nD2nVjJMp22mhCzkHI212Eg00hrdV
xqPABWmz38TyjHEputWCbYudMMp0Xy7rqldUKHIUjgsd3uw32NhRDIxeigV9xdRT
h0s6yQ75f/Nd2yjgpYlmv6O6nadJt+cFxNPqx+DgxgIN4i62MzpsDBaWaE29Yglk
t4VI+PIPZnDagOvH4VmURZXY1YxOKf/del6ekuc5HqurTan3HyFkHT5RL3CsreUH
xcT7J3dJh7L1NZUUIWprN0VsuUAoeQssxNkrDUy8dai0oSsaKkKMAYLv6O/H82U7
5J3TwTrRmEsUNU3k/nCbla1c3x2Sr/KtJpboo5f3U1XpJ9GimsYJfIoKBzMwilxT
HQaupAK65RuMVnY23zN6ASYriAOvGhCU2RuZczBDMvcthIgREsRPt5No8l3kfGHu
5CkCKlXajUNU2H6j47NfYqyQ0LYWMmUi/65TbASbqW4jt7KAjKv+T3/LMYfXZ9ir
ETFl1Ac/3Kd8wMvwua/nggQRo7Ugq49VqQBJ4WkVu7gOLywktISjV5unZXyykgRA
JTtkV4kNsh5OK3YRXscmAd/VniZkNPZAPXtuCV44M9zsX5QZPRbB9KIwLA5T5BlV
nypFtPCJ7Ny1qeQzXkJB2fc3z0K6l1PJZFYcgNFz0NBK3YQb0pdGG0+8XLxmceYX
CwEGPkxi4khMyt+QrCnMk44BBlpzaWSlHVUhPee3mtPa2V6heLoNMSA6+4+ks1fL
Mf2VPwegzitSicfT4UhwuDCUMVzmn6eJUiQZH6qR50C3OpIHqD7OdmioR++xgTlc
B7W7rxO779shkppQh5v5NOuLcKp6Z4e75jS9ih1iaKosLFSX52pUDBnrXewJJcix
NYV2sfr9ANef8ezBrqPZTzFELWbSIJLoHTLFfwumE/lT+u2QQB6Q7eg86mkh0zQ0
m9YWaCxckJRN2fMWNyyFY+JTsDPELj2iCZFmbkeLWYQebk2RYU2Y4Lmg9HCUFS23
CqCpwktw7KoIUQAjC9oygNEo8BDI8d6Dae6TMSAQgDAniSt8tOFxnuF5bC5ZM5Lo
Pk/PwSrFL2Fbk+A+SgWDz91gsYUy0iRD4Ri+15BTGgONNnZgMyFn2xd1UdL2dt8f
WgWZb83cCAaHbGuw0gzCAGo5E1yfHKSmOvQlLrFRPjlHrVixY6QaYn/mKnmiGMRq
ZEvPP2U7KEgcKBnydPmGKmEORI1I0hmlE8i8rUEc/6sD9HkuFt7SjIWJCUOH2v1W
XmZRdCSizG3HeMgjjJcSCyIV8qC7zT1sf3ezRZkVxRzBaAff2sazpZnqoBbfRm6m
/a2Y3bD/KiLYvbveD10JUH+2RUdfoZfFL+znUELNgWpnBIJDdxXghrYlHoI4jAZ/
Umbko7lON7F6umGb/+niR0nAdOH5bWM29CBHQIaVMKbXcktX/jO11s/09F6hLLvl
VgnZdF4+0+LgLqUOHhQBfsHwUFYHo07whMyPbwdZobvbHPE4LTDw9Dh2mLFJMO85
/1OC9wX7IrQdN4TRjUL365YrHqNSqw0RIimDvMNvkb4HqExRc2lwEc6MA68et/c5
pCFfi0F8xGscSMdxU5dsx2SjuvIwRLPv/x2v+gPm2wmxDc4aJf10apbc4C7u2SNf
RvciQhw+B3fv48uS4mTYeXPvRwFRMhC9RSQnPWIKUNLSgLiPwVZFW09/zXAwfgzQ
eCQrp4puXSSSm9Src2vNq2oANaSpOLRW/tVTCyuIjUK1a8eY62ZG/w0yCXwzlsVr
zsqOzb+WNuTimznTXhp/lxah8Dm+ttjm72Rxm0Y5l+Yd8G5q1FOczhJTZdnZ6JXl
1mAUR+OX9bnw2RIkc+YQl1XvXsF3Bmogkr/t2CDsDqBU1BzEuUp+t5Z9IEiBPm8+
g4ued7DdSVUOVBh/M2KT8s4B0nfgfFH1U0Z8Krt99Ta3TWwyMOIevQR1UX3zmEft
k1DC48X/w9/qdSXVCcvMPP5afTFrJBQfEOLWGJ86eXQDKDmCajzvkf2EwBhY1+f2
D47KN35wRUhgawobLb/uunPyTDJqqHP+8cGMPV+FbjupJwFOjhCIm3dkt2ZCiFe6
icpqk98jsArBpzSQGOwVjJNRugR31H9CQ4hhqc9Nhpb1mhOJWdZebYsalQq0NyWJ
zDGNI1n1PhXTywZHl7tcfkvEip0ng1wukRhJ59GQbUz4j3ByYZLvsGSGMreFPiDu
RNz1B9JC1QFEwju8MkPZEbnc8vKCFI+ciZz/3/U7E6r9iG0PGcqdt3cAqw8EgUGe
Or1SAlkCMyq4mtbptn+ZpeSfsXeOPi3fCU4JwKcwHRZzE/qlytE9tJ/XHkRSATyc
GaRDZ8ueq5v5+p4QAOHbHcc6UsO0l8o5JgEjn4eL1GeSxxDwpGrAOwP8P9RvNUSP
Xreiju1zDex+HvAsInJGv/A9CYYS7MjBhtP8GUIcK+vEaSrfXBVMWVduCXQmBCe9
QcCC4to7pkg6UfF/s0XS0QIJRU4MSt+lBFDkpuErvHC8q/gYUlyFpNbS6+lupt1P
wF8QSvX5hYp4m50LcvPzVWE2vl7hiKPUCLHwa5j//7y9eAN5tTB3Q+0NxsSKe3HV
iHgzSv8BPsGdCNr1dt6AYzU2RQClZyhR5r3lR3kgwy7xG+scNNPJfvpmOiWHJbWi
8/99kuHfE8gBcq+O50u2hoo7RPel+e/g/oqrKjNQUks0nC8OvkLbOSi7/Oe4SM7g
94lQH/a35tKcZ8cgk8ucRdOpnTjXNfLBQrmJmChR16fhZw1frXXaLSBu8meBxDFR
twHCt7onkvvA6OOyNW0GgZ7d9vextjsRz4vE6slNYWEpEob/uL0np5lwErhDQQ99
M0v46Ytze9l8NCUGiTagG0vdCD3OtDxvZAlO7oPTq+syOZQNmP/WXxUpgWeGb/1t
qwDOwj418JF2RZ0CPOtQXk9u3Z3R4ZF6PqWTLlnTm4NbnLnYrYvLE/yTKamraRgk
54jXUCp7H8famNkl6B630M6Dr+kqrkAYFOgYWyKJXw/SaKH0SyMPC5MPxwgFsheP
P/w2M96rbh+VFGy+FMw9qehBo1z5OHBHVXNiHFPwqLvuwRkM2fYfQ0SUldTaN2Ad
02RFN7LhgLpLiPOJmUiUXyqxJMU7EkNfrOcYIFzM+wstGOtnUVCJN/u+Xzcc0W0z
lNlkWeTQ3fmIYGgx0CoU6mxR9gKHMCF6tgM/phDkfeypzPQ7QRisOOpwkDTNxxot
FItkx1VM+/gnxq91MtjBiEkMyF6zyybbbHksCb87R27RJ5X+SqAH0JcbFLrd1UfL
1K/pe7X4QgLiIEnjlBZWCVewzxZsNj9jxjo2VQEpPi/VGgMgSiy4o4wKRWJLfgW9
0nsmhihN+d14+tQWwoYcN4lkHT/kIabmHk9nxvypRAKfBoIpGhuyKXTUVmqhg2++
7vdCQhIByNJJ/f1uoz/9N/wj206GHHMJxMchXP3QLEFtWDW/ZvYJj/fFEn3CX6c/
9/fKC8Nj8Ypbl1Jf+h5zlMKCp/DnPBTjg39ZP8yzFMzpFuoOCpH7Ke1q/jWAqNw/
O+ykk7osxSOU+TXbsF9H/9a2s293o6Ktp+1javy9uAwO+YRb/UEUdIdRg/IMDEU/
zfU+p0xR0BPfsysjVnEi0k1NXg5oX6BZDeENCJrCMPpWSNOMMeeRuvJi/GmgXsmK
Qeuh9pOMIYXLtIRTGdDipDyL+2A6MB3tvxHfUpj2AdRcwwWB1cQgeIS9btqVhxvb
XV7E1DDJnj6O7ei33Hv0XnnHPDEFSeteH+6C1wumEEJaZO1bBZht7o5VEPbcoiga
zl6kVhS6IJQNR3J3gsrEfQEM/Dedtf9HtD1NHQqOwTF1ifBklr+dy2FJQ1/Mxppx
d4ICX9WgCVus0EfDBraiKV57HhZ6oLkP1Hi0ZKLOjSZ7q+vSl6AIAOVFJLB3soDl
Pf08G1PbLKAVteN+8YVfENX+91wdJHbHAt++iafFZAwrTeSROOC2Ez5/Vpr59aG3
kvIPf/ySc8xVzZK0Tl8+MRLZqEQ4dy0vEC35UJxcH8ljpumN7aT4a6wm1HwSfyGm
cUcNMP1zMIIfp2FhHiz7iXWXlIau2ayUc1UYNuf0tqVx3Ea6EEyRpovu2mHDc/6p
bIiqs3s0cq4G7LoFttytF8aT2o7/Kw641AqgpaFWEWmTIcHfWWyLb/YSbr8zgPCf
ymfx007vyyLkLOVAPPKIdmp+a5HILmMYWlHZGbFfnLbDOQiMvuheRS0hFMghRdSn
+OZnw00VIlpQo85xPzwDwPF4weyqRu64bK+scXQqHQsTbPLDmRfe+J/kdihAeFL2
2Jhr1xDqNv6LA1Jz3vFlQRA3cgvwxlaBYFdt5CvsvhCuyVy/GfvwzFNw1EgnOyRU
FxtnTkRP4DUtalFVZrpfi2JhonuvcC6dIsdCu3G8XWaZtduUAPpnHfTtfiGu2+sy
bSq0Z+LtTzdOCYzID0Fd17yjtexiJ2oKKyhCFCuDe7FhrW/gJsLDwDCeIAjEYgdn
QEH1uu+wnpvUfjuaKc6elbSi9aeYcKWCQfzBpugi5P0+4jz6ag0dG9vsl3mQ5rSt
I33Auj3jdzflD0DuODlKUCf23MW5o03xWeIFDhojOcu4SiU9DyDcJiblBQThGAw+
3Nxl8L68I+HgXijoK+nFUz6hSm6DqYHejFocjq7hIa/KCW4WQ+uoKNGdP3D2Tm6b
mGjZ7nn/PYbUOpfvU1yafZwcuOsGt/Y5XiD3oqLwPjU55MGc6/HIeY5YfOd10A0Q
6qBngZI3UYx0Bo8kjkkGmUubq7EQom0i7AN286Cm+KfLGvF/Av33f1BnO/eQhoBZ
qxzwARoP8qvBB4JFE63jdju18B5vkHWP8BcOCve2VfUhW/XAGdXeDLKXkmIs5Zx/
6D1gLhfgaLnihgGRb6jogXkK58Hng5FAo+kK5JNhHIj5juitxtGZHxVk4SS+pEs7
EbwxRPSmxtNhd64IygFZPb/FnHC1Y5Q6Ha6Lu7aI2PRAbXQt82e+8KZ1wBeOV0rO
vjUOaSYEltrcyBGwyK/lI/lGW3lZhSCrh76jojcSOSPfjU+kXqxdXidkEhDuvri3
GGSPXxbeuWFc2fMVrjqVEjg+dbVkVkPpPWfwuYBwprKyjp9vDBM1Nfxn9VIo8qvt
RLgmvpY7oJSHD1ksSdctzThMwIeXyYoSJOf2M0vaHCB772096yevfc8IwTicCnQF
7ebsj7BLjRqdP1NpObZTj7PLhxjlngTCQqGh+JOW3iKHmsAqk9p+kGM/L9btHrAu
T4475XKAc+XWPznq/6exzkwMRZoOB+My9ZEDa3Cg7eV2RE4pLGczIcO77y4raKZm
WwDFPtMk6jfgm3p7ZrSsmnCEWfrshbVfb+cXbCJ/w3xKS74j5Iw3qV5x25b7PHnE
CBALm1KKIWwOwNg78F/Kkud9e2uo01Qca7aG4l44q+KpK6PiqHOQ8+9h8/7CUaM2
hua6S5ia0/TJpGevSwwz93uBzaZyILEDJdCB7xYGK2G6jDwyUz+Qm2EB8iIMsKBW
PI/ShhNVVL5Cd6uxiS1GYB1cTuxyIjJkS7Gc5mMq7Apz2FHB5TAMRZ9N02pLPedd
vuyypRLrSjmOkwNH37wytcwUe32Pu95LOCtzBzzIUWlutnH6EoTQHt0al/GjgMR1
5U7ye4YgTLjlYcAPS9gvDzN6ZclkjVolA1pAfAtcNZ9b87a2YEsWCo7kXhWypbi1
SwUA2wzJHhki4ez6u3K5pQvSq0lPjnN7gk2d5WSQBM55v1kdWQioQ6DBZkcKaNSB
V9g3iraRXF+lTSne1uGMRx+HX7pG3oSUf7liQlF6CHuaDFHCvWOADesv3z4xB1IX
MRE2pAa0Ij6b0BtplIHcoPLZaItp/+nZKAkJCz+cGez1IgKyPlnBi9kwdSJRSgmX
tzG3UR5wCIVSwTFfNvLy8T2nBp+OVI/j45f5HfuYUQQjYxr6MQn6R+ugGU0zdIb9
KEhpdVctMa6aJMt/TX9AW1cO/aVhreMF6xhcdIJ+sVtFHVRKaOozuEBQFVlS8H1j
16NETLMLlelSSRqgMcb8iHxc0vH7o6HZ35ZEwt4Of+QBImI+fJKXzyR6/gxCUix2
7O06dkgniIap2QHBxTXSD116Qv0xyrf3UNYSSejjOPYLE3Bbk/TWg94BRgYYy8TF
dn0FAGjIZNYY0lXeyAg42dQrR691J1NORJ4uGHdOSs9nKfKZKIXaKhapEe1vOcM/
apvTEpejiiZ/0Dn4pEzllpvuw3D9bFKPIA28OGNPE21AllXWD/NHXH6qsGVk9zOg
vuKDnw4dvajuhJ9SdQagSE3NAh9LkylcpcbC185+f8fuxwcya5+t0Jydh/cYnfI3
2hosPtjjp3wRQ8KJfdaEJhBlOU1rzsWeU5jNVvPL2oyYgsCE+vIE34jDXeI+eKzR
MANRA25zfq4rhnWBoWU0agpJSCyrsG2SkMDLebu2DauK5APl0FUbdQ1sBnkIhWde
xuU1VRF2T2vHeF9NRuKkbALU/OWEn3wo822Ktib4YvVrejtrg2SYQ3VQF4bH+4wT
yy2BojJvhOmwxTWLj4O4Wiq7I7l4V1/8w4tK0NARZQhTy1S7K0gFFFfvEX09tapX
c6SPM7cqGLcMrygh8MaeyMVQIM1WDNhBjwJEY8zXbvf67gULL3TTxJRpEDRXnMqr
qj45Ep+EJmkAWQgzrj4hwhaCgbMGgjDHbRzCkYaK5iJp+7m2aIvZ+ZmLuH/qEAFS
9NlMrtFZa0+PKvBguutSZl7ebQpyFeXFzxJBHqr3TZa1o7hn0tnRbBoBVYOMhh0/
sYfLDmWXc+xhMdQgQC7i3vXwngoM8m7h9c2cl4bNUX0+fVuoGGwUNkiGa5FR+QBj
tQoz6llxQyEr2Qx0NHo9iTTtOFLJCUug+N9GWWnjUXZdlNZ4rKcjmJ1dAPuu1RJ7
dCndURNMV/uoejIQHVS3V5ZiFrwAW5Nk+GpPo11p37s91mxzhiWE8gZ9yl8EAqVt
85z3sWF46M8jwFNs0Gkt2C1v18Vyz8NZfc4Pcg2JcvgMQlvS9GnDPnuKmahn9Dl+
fy1aH2lqcLFnZkRNmYKt5ReRTTAdhLKIWoZOxENbBWaB6drn6xcHgUCRwdKWuQMT
x7OGLNUlYkuEpr5B6utJcl5rR59NNCLZB0uZR5vRoXWFXIZl4hUiowKbPmuO/7vX
euPo13KGMkRZN18Sk7TRr6Hl/lss4BP37se+6oX0I+DHTa9gpluAZ2NTvBtaKtxG
h4RD9/H2sc5zG+vfxmMyqyPOc3+yMFQJD80NbCn5dzxH4ouaRLEw6dPUK3hFXSNG
rB6qzTZwrPPf/kUHR4j0gv+tdvhp0GAWHBmJCBr9A6V0YfZItlHDh2A2NNiaEauL
i3149svLmPdo6mw23IQQW/cjyVzMkL7lYfd6l8VLyF2rmuq/LSotIW9/7ysg49LP
K5KgLZa8490C/M2CoQ5W5T5L97FYK3KNS8WBM/AaYkAm8LaEOS0HIduWtkGAlv/g
0i9bNjZGkaHuOqTEaC+8SxymZJ/p+WYTCKV6Xd/b2m5Ks0C6iUu38KH0bMPjdEEr
EjlzoYhbz3peE6LQX8rCfTkWW9+niE2uf3syUrVWiG+lRqFIGchgI/Il0JMKuNsQ
qfoVcmu7diBjD4D92MwH1on/AsoxQH1oCxW7Y4jMwPIREe5LgRmHGVFzILj4K7Gp
SiUvYYRQNIt7MAal/zUGD54lb6ecqFkLWA0tMLCNjjKa3445qzshkQC6hy6iPGGx
rSEX99U3msMVjJOudEeqY64D5acDd/nHEk7W20CuQa6Kn0GjjnA3PYf5laBSPNqw
uXu5kpaOJdxH0qak5AzM/fmPzNLa/qHa97hCRnhEzXCj7c6ke3vCX3bF/ix6csvT
NJExZhyV3Z9m4dTnd5Wa264jNtLSjrDhuDxw0WMaqWSbNEWhqDE5Ve8JwVPyAIZn
00O80UMK7SS8bxY8gssdhRK08Z4nUkHDXTZc46dX454zN7KsFp1c/RDQ0VbEOPVi
djdQfshmsXWAB2WUK1CPY4ge4WHlbe9DZOmI2XSKjRUe1RUYqUWrNVdztMPW8sbJ
KlPAyLazeyGFluQYjfKdkPrB3wTB8DwkAyfo9wP3Biq4XpCGQMyJExpbkOVSCxxW
WeiwBqOxUxDeom1Nilb6zTmp9QHmy8pY/I2mfJufBSjJ9wY3+GMCJkGoXsrY9xF/
i0RuuXQM/67wjSRB8w8LEzuGKCFwyzGkFte7AXD87zkjR0rNWvXUMF2AyxGXWltO
JxfXyTzbtyfauGHOVN9LOko4494tmgcxiNxV1WSdCWRf2Kc9WppzYpvfOcS678yW
svRnOoS1FCXz5gqx0EUgc4sYoH3eOy1gTaWq8Gv2w63jT15YyCZ/e0GfYPUiG3fQ
ERKEw2YYElnNPylymsa+WQhn8WEVa+I4UzK2PI4TWzcRbkaBICiHP0wlAmgRKaqK
Gn5LBZSKRLPW0Hnu/l7IBCJiunQgVgugqPlJ0xGIiaBcCcEX2wJ/yLc3ftK21lN6
Km3CdjeTjPgRFqKfgrcYExJijmNm1eEkL6Qm7ABAm5wAjZBvBvemn6Tzrq+/HmFK
hCBVaT5zId6A35iRDgp3lyZ6pG+VCnBEsXXHmskk9psbQkeDL20SMUSqRiYt49eC
RHVoEAlK0efI8HnDrzPQP0QQ9bkWhl8WXz1nISj9P3K1ssmUQveBWAZydhYavHA8
fueBaOczaEglbhU0jnsuOk+Br3jdhBe0Z5pNVtNQVgzv2/SmOsPX4e0sw9jIrEFr
NW576SjzEzGsz5bgbXnd0+vEyt420f7oPKPp7Di1//RNoPqqDclqdK6K8SpKwDM0
qMaGQe0KcFe/n1auyqDbcvrKJpKzGj3kSdEWJAM+5gsrc9QP0aRiYynNDSLDSVOa
2p9b5Pj4GpOPxwBgAEmwHjL1v7K2xmq4HyuOWzNOvXLg6pol9JXX7m/viS9fmMoM
i0PDD9RVN8ePsn2qhZP2G4idJV5ujJ4StHrZp/x+CzoZgIUNdgBtNzLHEUXNBFPj
P3f9CMTa/umN+z9uMP7YXGLwqbS13zWUSrlJNDqw5GhY3/KxHB8QMwcGopYE8y7x
cOwag6DyzscZIwF1sRYO/bPtJ+j8K2z4mqFgzk429wkgDzWyznCpowQzRf3hULXE
m0FMo/2jrmA7dDQeTyXg640M3kaQWJ6O45NkxvERSG5bcWRcLxrt6RNakH0X5Ux8
L2Gdib+TuEU0fAMmOW4n6EGwnefP8zTfn/PJxYSiSYtxWHEgv1txSmMmL0Hp+M2W
ZO1rWoPLyA+ZVxxaHp5/Ly4LPxnV5b0lYML8V1PxhYWjY/gqAv0TYAwwZITyEc7o
r8N5ud1Atsq/4qLtOr4AWcUaybpw37VA9LsvKLU/pGJpdi4OF6QVBZeL1fOTVcg9
aXHUYhD8ehuWqQRH46mMjutubI46Hi607Q8d7GUNJIGJeP2kHcDHFR+zBXp0bXMY
IxTkNYW+8CUtBItmbndgB4ppyUTKoAXumvoZUUA2LtCWDWvKU+Z0Dh1Al/2pDyG/
E/G+LpkTKTljR5H2tlSTbU5T9DQrxxmXpTpyS3psmIdpd/judNpXPY9Cn1Gi3Vn4
HE9SRWdB0O1SHzn5TPk++uAhe1DsbH3JmSrp30jfRs2gSHH0jufYtbIzdv+LX0Lb
p7jVkSsAZEETCL+ysgHr4UUCW6U5501nIfBu29rcZN41FQddj40PD4e+0Jt2/sj2
Fx4h1R22hP8TA1Dnulxzj0bf6ZvA0IhLlZaKbP7CFRg51tHy4JbtzHhl0Se7zj52
bNiIKOkpYulfPklZ22WZgBHTC420Xa4NVl81/meGach1G0UjijiB1sCZtBbu6n0B
eznMv8UNQ7tnmppxwb/iqDImJxRzGwZNNruOZXiD8QmkRGFWcMAP40POOiBSh7g7
daRidlcOYtKK7PFalQ1hL47OKXPTLPBuYwrmx2TRD3WX0TqSRDoh3sX1s4jvxtKg
PcHo2aP4P533R67awq/J5EKnRZsveF1cAECeH/mWg4wn40VcUiZKq6jLwHzkajQf
hW1+I+oIjdy3gtAQEH/2osQwCE7woTg/ip7ogLukw13ZuJi3dDq5XJGWaqWo/TX8
gfbfKK3qme6MWdliy57ACgJApvcf/GM75EOeD0ZEO0Thb+6b9BUGtwsydDAgdlIC
XsWXz73AiGDdwEgdeOSzD29pFgKkg6MnlbIYRC/UwLGVUkeF01IENSqbBHeW/goS
o1OPFsp4XLHfq7NtySDXw7OmQefpU4645vVZ/8l5zVbXTDCx3Wo8IDqGpW00FhlR
tUWK0gUC2BavIBEwix+P7sJsSpx5bxdxaOUZWwGR1hg/ynlJc2k9OHn9330B/2gM
IAqGqUFzrXEWeyoNCkCdgDaASfvzJjNnGHklX4JvSBuDXP6snTSfiLbwcKOlpOv/
eohhn1IYsej6m+rJHL4uI1Vw6oHk+Uc70S2i/Dkj7JewWEJlSmK0lf3HhKyil04t
G5xEEbzM9lqQSWETi+B2YQeh0oMHX8TgDRdlPsjFc4vW8/Re9JAFNwraQZkgtIWC
Y1BmLMzFKd6y9OPvqM//IfikQbXu9gjSmLNLwBvIm+jxaDeg1/g/iH9fMLrACgVO
WPJ7utzppxTdiCxLrjrtHfV0mkeOcxM6LD6PH7fbe6sm69YNmuFy0jLjCR6Z1l6g
ULHTlM2Qhf2EI5PF6DgqKVqeOMR7UcxGumgmFIgDrs0IqePvS2Dene0F4Jwy4klt
vmCjDVPgXXgGLWgDcWa7M1gWS8/PJolarpIM1OmdbS4wfl8PuRDB+ZVJueUxQZYd
K7b4T8bZ3FYuW8b5vvuHPcT3FEQ2lt2PElSkGZ9lH5nEVOFL7ZOOy3BF8O9tiqN/
a4560sKmste7W6/xiZiF44cBJ4EY+IxZ3NWbArfh5bfvIKofRpXz6HorekOHU5ri
GrSznQbCBeL0dFyE7tOvGKXm/l3B8k45abDRvhDL1jheb+5+WiaBp/y6p7hPbQqr
3T4bvLYQ+cTB0qDcFLYxVaeZ1gZzms+Yl0DBu/6j9SZY54ybObzJbbtiNVZOktJn
xn6NQ8TzSoers+TOIPqCefCQqGPZ0/INVsVa2uY3270Wt0QGYzxFNpRhwMQevN3+
s4szRpoq7stodEHOVYj/AF6/Z92vMK/08O8CIAhzFtt81mK7e4zX0FfELj4n6RZ/
O6y9NGHytM2/TKt819+4QNewEaTJ+WBM3iam0aetX/zR/OLiCSR/0phFfyvb2eBV
Zi0fTEpRmKxisTDMeqYtAEH9jv4EkbNkHc+7ICA/uLqUpK6kgGbd1y4fybjSVyQm
Ni+P+UvjYl5E3gQMkhnn+sz4Hh3EW+6EdNajyp079ezbkcC1vpfv7lP3+agZdyhq
pqN48iycJw0rNqOHG6IePJeS991ZK8ovhl19H4nXaOpWTKF98SVSH7dKAivAVNZk
tzEWe+8EMKvK4YeiOViIjmuR6MUJl7/29IxSYfXso1X4oJnkzoLYlZdJpYDim1my
HTO6tdS5UqzPOU06fGgycdzupoGnQ//1vJY0FRTxfXqmOTkR5ccUm7Bo7h4j6ckI
H/bGY2vQj19gxYsbnbU6oGV/ekrTFCwVYzHNjrPzsUO4yWci81p1CtxDf+cD+X4j
O6rwqNpn8N0Vp9pVYdNH9BhWmIkG21y0DUAfRq4+xVYPR5CFDv2xlWPi0FqWMU08
pnyyB9/J/YmfU/VExJijzbw6Hxej1d0ZPRey1Rbt0an5CkUTNrieqPiGI2fQljtR
YashXjbvdV4OLKA4ApKFsRaASiSKjdGbCfMfu/OUicTDcxEYActZucoluvoz79Gz
ucJ/RRzenUmxH/UxIuBv872q4KP6dHIKy9pFUWGPWtWc3OQ0099WoyNkmk3+yFyF
CEq6GM7neahKbfMQ8H26A/wHxejmhRmkM9k//nOXPivsS0EeT142SpnsNLgip2SB
HvRhXReDGLudZ1PUDHeHy89WyXpXVzElL69T/AIt+C8KTpUJeL9mfzH/Os9dMRcQ
K7mAL7wmbpdQN/L8zBAJhueIxgzRNMZveBBXSd5BT10ES+j4hE2KJc+9EL9o67K/
sVleGNhgETMUJK8h7G6TnZzLxk//M+JEyYNwGgQ3dK1fczdRQjgKJfd51Wo5LRPi
LNVThWdfmHwxlh3IfwW8aG7pMYEQpOoplxKFEgviW4wroXePUUPr+R4pgJzkoMlB
tmpQ9V+v9uXQa69bR1CAd/OHZ9QO9fpB655wOqoHcKqKl9fBTQC2KZK/V9fzPfEr
TdZNk6Kj9ErqAf9eNbSN45dSbB5sCqmIC9qf7gClPyffqUCJ0z8ScgbCjMu8k03M
g2cOt9mzJG/zMvM71fomThT67RNijYm+SAtpC3gvgLnRD00rDmkKtyzyE0ijyDgc
lz8xEB1a78WtlDfRWxUi9dmDzWxvImL3Om3lJwzXQPVFJ3cMJHBtppSUbORjnbfN
xHJphKK06v4jT7Gon9a6Cz+MID/FiJZrmyE3JZpjFy+cvYw9menBxQaSbmK3eNyS
o9pkAcTWkIs6zgkjYroyeFrZyRnKWJRPr10nMFuzmlXqmmhmiPaPP/f7KpnU/uvq
RW5V2JMaeFinQHa+zGHb71fKIVvXIyY8VL64L/YpFWC+jnVBBdXak1lb4ULjkUqb
zdMqv5nHiKJfZz0pzj8DWHo2Mwy+5EdnFISNlalZeRPfReJ0LHY8tbnMWNBTdFhD
sZczWP/pVoGqr1FRQTlbyzmqB1cgSBbE9MvGrRJHEm/S0Yk3q/zUhurmb3hnlZcZ
ByMe39ZcISj+z6xZgFvfcBEA+5udrDcyf7nFYNoq6ZPXveuY7qnLtzuEekgQj80M
QomXMAZwrmnpE8FjtoOK3W2gazqQOWFStfgw52aEhKXtFMdgaAEa23ulu5LVSHx7
qnieasIK4W2nA0Wq8VKhkOvB31+EqbEv51/l7rbXd0LEAx9NtLUOWo+/LfT5xsaL
YqRAmRGRT/2zoNJ+aZ5GUKggDLrIKxWPXlXf0fckoQOZ8E63D4qgJAEY8xKgpEJJ
cd3FVQ+F4vtABjuU4bGGgC0VzGAC5WvoqhvgbBYJHxV1i6P1EEKPt+hTWkLfCA0l
COev5gyY7sLFcp1EB87A6ZkBVPUlD3YN06KgOzOwreHB5X+0FTpjXt6pvjt2wa3j
A/6JK4y5orNKHVqLE1YYBCpxShoByRbOSca5BHRC/dGOQst2Xy2P7UDbYpQ+s05h
VSqQIm4Avwg7FGRL9Kjf7LLENRN3U2UrcCksvaLscsagokRVHgUg9HytNa2KwrnK
AFe9sZY1GmaHehPeqlco69h6xmOP9/HZ9Im6u7F+nTP36dX6clCPkmPbq6UGwxi1
gv/m3FoFNA88kwUqLg1Yl27c8tCIDrtAU0svxV5je+SDjefuSCslQ77hxc+1IfjL
WSgk7bFeMvw/s04P6Xt6zhoR1N2gBGhoZqZnuxoxf+mKB7wW3UBzYIHcpK8jQ5zH
sGvlb+UKM9bRA4b+mqG5K4RtozUhaNj0Ng7yOULISKxiv1F75+ySdRCCXf+h8Q/7
Obb5QrNLKzAsRBCoWXMdlQDDmMCuCTTwy3/eOd4OnADp2MnnqhnDjeotBbNQ/2/R
0HihfAlgBahx7m4AhE7/9y1LB3Bcgds/jWNObwyVMQf+IZEqNo9r8kAWYYBAMghG
g/5hcSAYQSSpFBfk4/wuCpZbgTff/9sOfmYKstEcUJ18sHk5AR7cV2Nb/5G4c01g
kB9PYeKx5Yn0QPZzAeOrwxruHaLY9S7MjAMrrZuHPkPUgi37DPKsvrug0Jx6rfWA
nXMcX+y2kRWhhbb94MUa52wWPvxEPqB4rimKZUw1r3kSfWYo1V8DUS860EmQMizZ
89LI5qQoT40Fz2r+AI21uT2PgUbpS5X04niEj3v5qsFnzPIjbOKzfcrnRGfX4Dgi
idYeJNy/3KhHz/GKJqdwUVnf2dJXh/SGSdPhvbMuoY4bD/bxWuDuDKKBCBdI1w5Q
F1sCP4e20EduospnQ6lo7WAhde0jJyPf0cq6UuxBF3S+IWv23YGsgWIIu+1gxbYr
6h7Ea2CmjTYN2/yaocvlyux835zIQIZxotKYMFGPQCbCpKQiz6hZbuCUEhvpWFhQ
l71xK1iYHCKW51SpJWuKXYNUu3AynQouxz/XVuZj6nper5pqNMBhCulTHwp5iBrE
ectKXqKmqTQMX//ivR8UUn1uURQzsxKBnmJRJO/YUtSWs/9QueWpqAOUtWb9qKQv
s+wkqZZa1gahoZZT/H56d3j5HPAXBt8ITyM3+2TmGL4z7GHWxYTt7QB1Q8o4nwEF
5OyYfJMadDv1iqnr9xDUr8i7b5jl0+EVCdRx3263pkb0PkKX93EDF//RhlNGLOEB
61KDjCVLp5xGgGWBycoFwK8P8AFZ2HqwA9B1Jc4Hj2pAFeYIptdNW/FTVQjFQjTJ
p6rfHg4+I+bq/3K+ARMRGPFA4Cx3M68UYVcIdWoZhLRWixi/vmU+zKEbNPAzZtk8
4/vnQl8V/Bb/dADpKQQAYZmlh63Pv1yH8C9hymv8lVG97kUESXG30QmZF1YtffT+
QhYgyIyoDfHiU4Ay+75jH2udr0onpejDW+qnOJslFtUoiwNQHlgE/OvuZAux9aqb
a32EkuMHaYX9m2y4Wy/ju3m+mXiUoOTVAZglG+G/qfIfOF/1DiWlv3grVtuY6/k+
LIJxPHUWKp2RkQmlx8f1ZTSPqEjXe80qM9dwDOPc1l4W21P4CtXuZNblfHM4D8zc
KdMHupkVDHSR6sfAYBnaFrhmxYdoUfnnorBbNgJ1SzBDZCwUBAIs46puX+gAlAaZ
HIiK2p0iv5a5JfcjQw5XbIorg2JW6VUUM86NmNC22N9rYhZfOfglqL+ooAtzewds
ufj3dMI0so4jajPxBaRcEJcMVP0eer2ZadvKg1V7YD2gIT1mUWLw2dCJPPJBOMmZ
mmiZVEGKFXzrv+kIC8G0+nXYUWBg4SV6tHm+GcCReEz6cf0kscgDaNCQJyRF1R1d
zfV2GYLb5nvPXDL+8rOOc4+t9MHhL55/qYzhwsY1pCZMOGEEikGPZ6chCcn2zqEH
j0ntyj8MM6g4cAlO7KfbsC8XWlONKNf2pvLbcGqpH/xMkMSPkKkOtc9hrlfeqwP+
OT+Wmp1pNJvnKofWIF2wpuecMMoFIRnIkcYI8i84zxpsfuvrtOMDXsNmALuNwZ6P
HyJMqcteBXS++ZQSNCgirE7shYpFDyv5eq9B28J/Xa9gPAj8cvQ3ZArE/F8HIOjG
JnGKyEONKAsHyCx12pWouU6QBLJgqzgujvx5tJozdqjx9/bTLe51/stESKq+xTRH
I2OXXzN+bK4CnYsX1UxkQBuBysna7vKQxyoexKL2anSOcXCG50K1LgxabfvStGKj
vYhPgcAwisylbx5d3fQoZMu++xITYrb9cw4UHHkW6fCdXG6ivA2GN5I4dLn31tLn
Zhm7S6QQgUAwAefAfJTE/uR2YpH5DogR5e2UWSS9CaK1P3IXcMOLqsJ2WLuEPLBw
tBYWlHmR6yoM29S2vMPdHwg4owAboXfCNkXmzt9wYbmIuMCkx3Exzbi3nqRQwk1p
bZB+LcJfYDFVstKMwiw4pNQh+SbQ7P7yb8RWS0ODSUcyO/2hpFYWqhJ7foXrrFg4
rGju2h6RIrVEFaLFfCrf+8Fq4kfKxQS4sWccejf/j9ECQc8p61EuJJA1wQdbcvwD
dRJxSjPmfIJQh2arjrcr5bCus4/a01Z4Foqo7dYxDDJLpYBR5gjwwF+7TQ7/uOPR
rimDjY3FwGvmndmqoWyBPIvjQmaGIB+1uYjrMZN9BHKP55zbEalqYcPR1Yl3mxPO
zzuUDXotGdzewxvQzseSLBm/uUmtChrHdXUEYx+3cAm6LPZs9rQwHUSBcCvPP8l+
l0Qf91LUPmH4Hmt4WneXBo7H3QpG2XjNgabohC9rgumhdTFKhQv6YoSnr7+wWYlc
Vri+SBZz6fHCbv54q1BVnKba5oaCC++PnFFTl1CTyh5kHqYAwSvVb7lwHD/2OQVM
zGvvSN0FE45w9XUTngTHUp81+4dGEhGfaWLEUjii4DIqTqT6cmtf3/tBRp5oCXhp
dI6oFyUTz6yC9v6PJ888TKQsRHrhiJjrQBIQzun1F8UgPRaEIBlU64+9kniKQvYN
98PxOzNz3CEFU1UXBlkPkC6oUJdAIGOdYDEcTkHEdrlXPoyNbFIWBveVfjPkc+dC
HZTlwvx4uc1i3jA8n/QNQGAtU+BBQn7am9lmQJXJHafaDWJ/CiDW86gGEebUoYaA
aTvTF7ZPKLizgEQbYDRbUR6SJSpV5g8hN3ecTUfVy3Am1TPabQGxrro1pq+oHSGN
hRQFFoDnYkKTARf7NDNTSwSGBXcv5ULFP5yjBKcOqR7pYUoL2o3+Fl/xyoMDiAmD
SNIfE/8sOQpcMrsuwduhhtwzm9eImydl8L/7iTn7ufFoEcHqNes0nzlp+j7ceozp
8MRPVQY+4DRxyLM0leL93s6thL5lhp9dNugaTKlKIoDqxMoEmYHvwvQxF3GUjaIQ
pVyFiaBOxeLadXU7wTKbz5vYewrJWdBsN2o2judIsE911wXIL+HA/bW/IVx+Je6w
tzWuJgFySfAtPKZr7Zxl8MzX/XyNzEMbfUO7FFc13rHMPIZ4LswWOALaaTJKsdgR
PVodZJBUMhVgU3wiMwE/6Gp8WFqqS1FhS3UE/Dix6ltYWInz9v7Dnb7SwQR1GJGG
23beLAwcMCg5Uj7kBDvI1QMvmn/3hiU+YFzhyQXS5YEpIb8bK4OyiEnLI4agD00Y
Ad05nzWx6Rg24LYQthjO8PKBFYAWQ13STGCeCIuCwEutkD3HLM020YYgRAT18LqD
v+Ms4KBlBPO23VDmusJVPuYGCSbLqYcncYB99GWNqladVYsS+bpgGIs5bjNQDLjS
QQpXDmnoDZPcg+6eqGQJVaY0SeyBmRLpkHx+Om2yW/xXAcFomRKt0dMBd0O+TBai
Ududf4hDsuziQ8pSkhzOnDwFPM2Yy0PC65FMNf0AXdpe3+9sbIHIfG46r5UqF1of
8bVqOOUlAsrewLTrC4u1AzgOA12A3e1CktCrqMgDfg0d+JinDYaV9uCOSXdtmvnz
iAXMk6qHtpgMJThWipIM+aQfbQcD8DpdsvFBi2xguyA0kFIkNEeVBZdbU2BIkWru
axqOVUWIvBSaKQCaZtWAcfu5Y5zlSt9p2nwhB74BU9Qphgn/lCQGo28PYL/+Ow51
VZQVe15MXZYdMj1oPUcs//9qeBXsj9tNaExNhGRbwh31rkEcILfNjEti0Rg1czk5
Q4SsPItgjoCCnYn6/x6Y8Qng7fxVIKPh3+Nn2Ao3MwwHmaBeKL8iGHaTfzrj9EKl
Hu54GALpzR42jGvE0SR5+QZ5vuZew7ZoopgM2X6TsQiuPpiou6nxf5q9VLTj4Iff
+EkhweNZ53Vq9LBW6OiiFdJnsYCDghgLFxHpnxOjiN9Rv0UGRjn4ltVrecBNee5/
zTX6yL6XeCTlLDZ1qAdJogrPojQBR6TJn8n3HD0VFfZPGhcG+GLkKbEi/a7KCRbj
7I+4PR7S9/V3eLnlYFv6Rb0IxyCmbQIedhlJaruW4efdpw7MZ1mOiHxsokaHJ55R
kqoGg6o2GEqG/B+goRIPc3WUxeoesZ2AUY9SdtPj1JmYKQ8cUsb/m6cygiHFxm8p
KcgvMgI5ykgdUmDSwlC/xq22GOPPKC3APmGIoMaxn/kBITnDm7p+n+rPDVSDNvR5
up+Fjo330QrzUQGHovtCmWdpvOW3TByKS36ix26lzUvl0Tt6RZqckMFgBaqk/Yhh
2R+wk2lsdjXl42BMmHKxmcLMbP/8tif4AHygCqAtj76bF8AA4AouDC5p12FhRAUP
h2X56UmnwgnH5K5jFZxmu+L3cm7+WeJgOLeXhTAweGyf98AxfR+LDqA5+1jKz8mT
O6SAVq8GRb5ZdTJXm8HBKrxf3DBRtexqdYyuyxAJlmgp3CXPLqyg+yBjGGPXVVq1
xHC5yZpfKwghjRwgofluCTzQZtRdhw8XTrPpf6Ntf7MEixSpwvRJs962zYmBuRKr
vYZsNWCis5QPgUGmbq0k0FKdeiylWizlh2tP0czy3hwlOuRJfblqmcFKThyfOmc+
IZrIaL6s9NK7ujSLhZYvvC9Gpw7oP2/X93DIELtFS90fGT3qMJrAMxV+tNr51DT/
ntiYjk0QyRBTkrYYXxHP4ZAttcFPO0hs8InO4beV5GRtSNir1M8PfrEU+cUEOWbr
uWbcJSEpMKFoJN4RmV2VVIVGMZD/EB1FeC0ZBFlrVA8cEX1YE2goQtyqgiMFDtEy
FIG4dstBpYwkHC9VDF8ZFIpicn2EQwuyoOYfIClSEe9K2D1Gm5SDhiedetm+2S6E
G+gfYctI69XZ7IH3M9r2xoWLforqrfaT5F/lHZUR1qeGhZHiSAvs7MxtX5rPCZy5
H3+QrIunecYtCbR9OWeX8LtMdnY4bfklRRgXPXiSVtao79OIugeTv5lc6J5VKg3H
iOLnO0JnGznHxeqC1fFhcpvRc7Wn9oiidFVDe5Sti7iOgQmEW2xEW5nw7/ONPjVi
DhknNyD7Gf5bb5JZpZiq1IjPns0G+lmLdyns/A3lT+kz5crFlBpmbbGIhjNAWL3P
bSnja/OceAt3AXlZuA9lkI9o/+7y0u7u5Q9vY1VzkejkKA/OkGYLuv1cgg94lAYP
FIiIEAsjRNfZo/nOQqxgYyw/PQO73oth5W/xOC4soL92QCRlhdl91fIZQMDkixq+
CvGfpPr1eb2xA3Ayem1aVIQfIx/XEY+MqfYTOkeih4FQ4EUNU3JHxsd8lF+seH7j
FdMa0Aq1DsGtBXkf/8LpcpdxKnxtu5FvN2WGUaVsmp6nZWvEpsiE7YqNg0s94MQy
e/KNUYYvO4ATSADJY+5hr0ycK6x0yvXsh6io9iA+75aU/eNxiKoktQx2ev9CM2yj
/k6EmszTrLUHAJpuwViDTShpvHZMH/wheM2pi+pE0JUXJi8ZfqsL1QgV+aUnCJls
vkob6jpp3SQRBkEfQUwuF9AYhOiNUiBI017l/ZGT9nw9qSqQLXTrgtQUAP9AkLdr
603q/+zI/WnBduLW3Kpr6vbsDaUTf5Y8227grstSd7Gi44/0SLhbS79eU+5eeYWK
MCViEZ6ZO+gisGsokYar09SffRNDLY7ma1KtdDtQ2w2K6s/qP+XpJ82rDAW7hz6H
t1zGR4LzCv8ZKVM8d4vG/l572qq3gsvmydsNp77w2ULBQxiMMLR4GlkXV/1U/0l+
AxBsm+3POi7wJdxNVAbE3jANVvBBXlMDZN+45tPHrtTB4jKUInwGCT46PEyWMBun
dMKv6/A+gkMMaT3P+Ud7LNJqvia7+A/i9EsDNh5KMLGpamelhjOBYryeY6ADrYI+
x3W1hNXiONXhCkdkAgRplQZDkhywgJ8WV/TPhkgAvAdkrGitb4o6ylhAM6mJBSQ2
7bkJ2Zf18vODKJ78/XsTpbDLLcN5CnCACUcKUIz6NjDRr+CWiDnVPDoLDKLo5a9f
8yRx6zlGfMMZiHLIzgljFDrrVoUNIC/2LdJnI+ybXpyr1D0eN5K9r/iK8LNBpziV
zv8jhzlnXdTncZ+MqbzjsnOjQ9Gw2z1+VRIiLp/KfO+ykbNHlezwisSaGuV/+9Bs
fnyZH1nnPZ2J1DMSoyS7OH10H9dabGvK02RjPPmu5UpVS3Nh4QPd6CPfsuZyGffc
XfFEKXwaET7/3G/0D+0nYdb3qpNw4u1mOI7ex6MkiftmwBWu2y87Bza+1Z39g9FE
r4dIJ6d8OTpdwW4mxY2V+uffwf3Yr2SwnJI6yZzYC7nQPmjV3HppcdNgdv+SjhV6
Qt4bDi25gVgW3ElYNAxYuLFVlDmia9/dNazD+5BbdY61brzTCf+WxNxvUg8ZFZN4
D4MMEGigOsaS1qOoBImK1Dk0jwo5CBdVMkKXkCAPkVaJIPx03jFNAd7dB8CePBaa
fBEOz7vq30Nxc/HyuyPyyt4runRKW1qREOXu1p9epG+wT+KOXNQyR2UaO83jPQ3b
z0+4d7Q7t0ckFpRY0MkEJRSuM564dEgyiFNvZPMEhT2X2E3T7AFgEoG4fjBWwj4L
E/wg99tO15V3U0U3rAMnMcAK4M8OxhheMFC9uROa3SslOk+lt3N2kegKLOJPZaDX
6ooXC1/x4ZT8DMQbCE4JkDDScLDUMSlKLOE2JXzaArKJVBICymNwp2O69yiY0FKF
s2hV8CqmovvcvzsxR7CGyk2FfJglS8UsDQdey3fOR1lXpPsBi+wcy6GCs/LxI5Mm
mfZ3Sirf2XZecmDuNl6BjrvSdPdUOWRV9rNS2VcHVs74cJozlIM+CoucwNRN6sfI
50mZhmqHatjCJn0xkDH2Q/BaPRHhvQxlkC8sKb12i2Oz3wvLhRBFxwalBV2onQ7V
RB5Ya2SQw14s8Waaqc6hb4Yo3vWda/544z2luzAFY7/Ks05OSSIU/AHNjjc7WQE6
L/bc2XzkrGiaqFMJSqB/rDIcVkzAO93LVP6WCR7IKYiYzsRHCdo5mLRs+RvI0X+c
deT8W7hSIfccr23ltMFFMkueLWtvGtbdUd604siRz2kje9Oow5I5fyJjL/+jCOVx
YB/ng6lYGfrsIOOvT3pWf7XvlMjAE6u6xcemmKMnhrnF0vlHTaCHCmG4K2z0TGWQ
3+mFlHFjwvmRFBilmeWwydfe7gt8ghVVRDu+y2an1oBLm4dURo7t8QKZTxzdvzYF
oJK1RVkdT9CtPOptb2Nn9zzNvLIThh8Wjgl2l3zWXznL3SR9/ePwNZRu2A1+BK/i
Xe58ZXiye/JByfe0eGm+pA9dAUdYFYyf3LHVokJFOX/x7M1hzykdG4SOVOzT3RBd
e8ZG6vQpn5rC5TCbwtHiJMrtd2jl9JT3CkATpGwu52POf5gqfirsTW8oUPlRfSv5
JAx9PJAy7YKkIji9pY2v4SMk8Kdu45NwgNNSdnLw2aim7eiHRllO+OvDLhYB7Lr8
UlOsy6nwLHpR7S+m1OtGbKhXpiTUh8ULtCR1nUpw6tLzO+y7TraNvGPAsLFr2hLa
ndd39FIFp5ttczi4rxeBzIlf5o7iFfGPqjd0KIN2Y+1LNjDl9/0PRr1oLk4h0NC8
2D1Cfltp6gA5DcFfPm/xBXpfqNO3NqOdcxr21zuOVb+4mLNgsHV6KaQACst16ULp
gDFALa3RKjtBawkjgKLpoRBS3R5KhJiwQctbn7utTHJWsLr0qS91PbbHSukLQ+XN
OspENuLsuC5O98I+VziSw8zd/QOhc2530ohQWZ8zKPMMzbcAS65enU8TeIFk55eE
3t/JiwK0G4vfm8T7BW07mhb1oxvyTKvyOLEwFHUPFzr7lJW7vKJck+HVdY11jk64
9kwrMVaZVZOuplLD+iNnyEL5IzupgpkSAARcsc7/AV2THOqHCfXvFMHi4leBGDHj
sN19/zBd4dt7jvrkRsNbPRqf0IspBJ4dOZm3HzNq7bc4w53drxCpFdhdP02WA196
i7QtmGbW1PItzlQSC74bBUqWrRu44VCPkZbA/svpPeyuuSC23dMr6sxQRx8r3FSb
AP8/M6GzKjMoPNPcOq86lyPOrKqnO9kukeA04nG7jk3geCa/Zt9Wmg9GmJFNie0x
bcS6h3qU4XDWHS0mTXsE9jJTKK8Gw1Tqnsp/MHwcsIpaOjZLLcVtcaoR93Ihvy7R
a1EUsXaRIsR8kgeiH82DD/fgtbxH49bs6rQGdfYAMbOMq5wlel5P/UO4LHdUfvA3
PELSNjk0m2Q09cziHzEdvXa3nrusB1VtoO3f0XoPloLtQntYnsQ/Dmkk7K99hJKF
7LU9gXiY/4YNI+5pZSZv991kkoJxjFUrDCei2AjhPgJphZ11l9jfFU/hr/JUqnyc
oEHYDX22LLPu5IFnQ6Tb3dc6p4DuGb6qZtWYbNBxggCmjp/vLIiPE5XUF9vbsQn4
O4O6aqmZ4EHOHz0yse2miD7BkrvM1IrbPJUDKl+/g8FadUst+0INmqdjP4SQK4Rk
bDjKbdfF0SsCfpo23soTSQzkdtTaHgS0xqhfn+IMtGGYkwMK5wFLmoRwgJ9Jyqbv
r+WyoGTtiR0x0JNFWJGsXl+Ag/zKPuGyeY+ztyzASphPckm51WlRvVyRF+QRmdiN
tGW0zndW0ovfUnjlgK/FgztxtfthOhJPqHKmhQwjxlcbJyX+WK0BaGF0nMvMihXy
91zEku5vXbBaLCLGzS6FK1ua/x6sP41CPjkId3jRl5rcSETHyfAZ65XXdMfyVx+e
YRTaueO8owPNSEIhsDY3osbKkXGUH2N+HMs7ncQa+bEK0lGwdi0LMCMykux2UdIF
YwgwRNkfF7NhWnmUGPrXU+lWNdEz0eKpv+Kw14ke0wqpSl9hUibnNLiXpe41uZS3
XFeRVPxxuunOsMSOpY1tlCkcXlxQY9q70Rj3ZhcM4EJrp6wetIiGHPyRXIOG1mmt
HQ60Hl73S2fkQjgnDlHrfDxCiYYiLHpA9bBjV7+yN2YZFIX0qkyMXJCowkoyDM6P
0n74/uBMbW6mJsGVr4ErxkeKRu6/Sm5+ev0K2hqhkAdbXkOZ/y7rcaPR6ZadnYIT
MNhAcPr4XKQZIu4BuODlaNh2bhd5r+FK5QMsA5RuEs0Mdn31fQlLuCV9Ap8jyT6c
bxlJbb7FHWG/GznKLgCuVpBQbiMehI2uTAkCTYdeIdLMtPYURbGxtaD9hVyCIQhr
F8+YLB4yueZ2/UCpB2BfAD8gtsunM/xK32ndbiFzbxZBE1RAcFuhkU/ZPBzdjtZB
AQRBXq0Ag29iSHkFi+DSCP63IWqrCpQQ1zy1sAuU6fKYN4HzdJWDHTh/hnhB7gcs
mn3rpFeXwcxO3hcLn6hrkhuvNbDaN2VmvUy7OdZ3BnndM2jrlnDdok21XUCUFhIS
DvAabjt+MtHYCQWo8xXVev2g/2SABBGMCvRhews6n+E1gdFaplmCPR8pveJz6LWb
ZIwyF6bGqZ+f4sgljjzUZaxmBANuuL46N4PKN6IjlM43RfV74m3WQAOQdpD8Nkoq
JC4Xgp3cITTnk/BUvJk8uibSh0j9hMyczwoDdyXAr8hppzG+fyCG+ZNJWnF7tkXF
/lRMfqhE1yKI3KWQY2whk1HLx67OdrSEb7gcblAdwupsEWppOlG5Axu7CG5szad9
mCE5ptnfmDwWwtkWIBPy5YALHKzH4ET6LU3Hnq55rHxibpXVCD8H0KDKmtEGGCaO
gUCm4EyV39GgF5D1uVUe6bseCOsLkdzPXNuqMGFdHgcqS9DP86c/XF8FJyFcE8PD
UkPnQumzx3/QtiB6jZujon0ZuqboOPpkySOMmmi1HOgoSLk4xc9AeHbQo+Gt+Xei
+LMbiEurRzrfi6ceWxeDfM0HZak/3kMPawnkuvHP00Jy4CAb4A7Gsg+Sh4szrnRf
HqovJn1kK1Ld0cF/pQBYN9OnE/tGWG2e+SADrzcVUXLfmsvMXfdnISML7kAq4qnd
cyUdstBRkyw6yyff3eaJQ1Can6TyygkYIlL80tYMW42+q+8JKT0CP+qnw/V85bVH
c6a7GijkulK2V7AD9rF6wB1aTBegl6U4zQrQxX669+/oHmxX3/O2lHpwkcXIM59Z
p1UkonrjbnuNDkhqqd4T+7T0Z9bQxaMtxomUFvcP4geHeAOu53zgIpwg2ZZgdNly
uOA21V9TiBbMJCm7li269Fyt3Ldwfzr8+FcsG3j1DGLIjHM9h3GmN3jb7NLeggzk
wiV6wvbTqWOAaN+CpNA5F5DO8w0jgrkiWfEJLDp0/KZtOVO9IOvGnB+wL1DoIoFy
rkh0wjJ5dUMAXZ/FTwLOvcNMfWaGL7wwMJoycOtq8jZmaO2OnpR5aNlcWW9+TYX6
DP2wlvN7dgPddrklPl1/mlwfo2dWsqjoTWLS3sSpW4SPeSbUr7rLi56T+o1QAcxG
B0xKrcew1JKLqOpKhkpop0D+ZW6iZx+sXNon23rEh5HH5N9bylsd4vfVD3TbrsLF
KwvuRZiWJGTY+YrOQmn+tH+8xlMmn6VLbzd73iyOi7KIdM3IUsCyQg+qLQ2vLltV
xref8BSkRpHIAPVzS7F1WcevuDct8k0s81uRlhQqN13ZLUZdDbg2Fju0WE0HSWy4
D+T/JXMr4wcdrU2rswEeH8Zi63ge4S9B5MQaAETVXVY9LtA5nLKLCJpx5CqZ2HgQ
KsAhC0Weo7HtRuorGFzKY4mRiT56wheEgzLh8L+4Z+sLb5IRJLqOc23PIVtAnm7v
IE3AtKkh2Y8Zl8E7Wl0IcrOdb/UU4ANa2SQmVHBek9XAiQnU/wmuurIfYs0mBMF0
ne5HX4w1go4If2T6T10/3IzBzRiCB4sgq4aZq3DhdJDGzVEebsgbdTzTalJDRLD6
rHd15TruoGngz2VPD6dzHW+lnvAPre37q+TtkuCftedeVDvL3H9Wm86TV8H59zMv
9kmSGLw5ZnMhr+GhjH4EFWnlo3oHZW7TtcvuzM5Ayc7m/oclEHX4Z2L1G+97kYVT
2CgnziB4KsGpFO6/zG1hvdL7oIjiPcPHeRa/kOlbyjEpGNGx/eiFhlxatXGbJa6l
EmeGGWev43e1P3aW/gQEViHQ9nQT7TMIdC0t+akeKPl3dN+syNHtEc9FNaeb6Sso
AXsgLXcXUNvlvyXumcqtLvVmJJZwkHqLZcRgfhjfm8/djWiJdOviMhDUsOSoEkG7
K/wzWPuRzmcyBEQu0iLM8ZwEJaYtAWZZT0ytR66xk7EimYbql5KR07DGYxfj4dkm
fsK2mlMnHC9gCGjWZX2iCfJQ0vLSWoHubcp7sa7S5j1PUQxSorwLpAeN7zS+kTU1
5qLHbMnPrrQgdSBDxD0W+H3Fj0qoflC1XMOGaJi3ISrOSFnXmSVEO4EhpSUbAuEW
nv7fEqQ8XPSddT484S+RHqSLfTfpsSlNK63rT91Q0MeL0urgkWIBQyQTz/dB1eYk
0Ge7sOPoMBPx0rLdV7rAmW92F1qwg/JevHcJopqR0NJSl3nvwIDbDIYuZ85Xb5Vq
oI+frwwd+TuKGHUrXfztldzPadi80YpCQLousiOGLYYRRFFUp58wIyBIheUbZ4jR
a/3Qi2i85OI9//aX70PelNERWrw+QyALmejTh9L//eUjj+0PTxbDPWg7gUbKOGWF
RhthN9/HN4aZeMtj6Kou09R+p42e+RXbDWwFwkpJnL2uNV3Yl91NBJmrKpaJv4O5
yEd7vsxA83vjIc15l3/Ul6pc62mICMK8i9EIDds0Gy3KsnFZFx9vwjMzf2ZLqQaq
AzasMz8WKhqQnSrApN3ofiGt3z6YiqOBlVaD7GT3G13OoSOe6tu09hs8o8Bn1Hvw
2fu51Fh7+BNOts5HNRqMCfw2M2D7CvYnrtWqLCc/pAUqyoyA6G6ANMzj3t4P7Q1M
jna/MsT1YAPTdhHpe/Xn39M0UOszBscVTgg+7pCfQz6fcujKLg4thetFOvP+lkb6
gc1z4FjwdZqxEWf18sDERQHzeWPDYEEmW8Pen2oED3/KRFUZHOZyP+na7TyUEJe1
9mQ46YW9nq4W1JLW8cbUl2gH36kxHoOTScrkLpsgCNXnPy+B25Cg/xHlGTaelcF9
o67bAVrAs8Aw14VlbKVoSG4bFIkDBNGGhkyMlJimqVw7mithqjvssJumMIr1vNkn
yPizDiNokffcrrqydl7O1nl/rvpUPGosDVeDm+PMsPFetpJk1rgiMs0f2yPe/LMr
tdJ39yXGQszVEzovAg4QSJwR9mo9b18U5crnvys7cLN065eMu1qXj14/r3EMABT2
oqaollnDewoakGfVAU+TSvr9eh1EXdEiSdVUR3MMpjO6SxyXsO7cCj60XEAVuaKm
Z6ePTSJHDi6gHPTWrzumZtESxwKYVV19++cAcsyIqyJ29IQG3fF0+UTmCKTBZk8D
eORwaIPgRCleqil2BevQ4Mpp1T/b1b3kRQJL55+gvOh6YXbROwhoYj4zn4mccs0Y
tCA3K/1IoLGfvEpFZW/z3FdvN+g7mwdp0FL+4T4U52b9yzfksmb2VyFLGSbK3NGx
NvMngbnKdT/zawMnUzsxXfgw4zyTEbML1snz3f0E5Hf7LCjZAm5EBY8Z1z07iHiD
0G6e/khYcAqmw0KXd5k4Ew+moxgDe3jh8imJC/GhWdSTTYc8C0lyZz9rQMsl/Mnu
xl5tCOGdzkkC/FV+GEfxmsgbY4KEbiHNYzsH/uXO0Xhyu0ASUPF4IxUFfWWg/BgA
Txj+cBwK01YHP5FX11BWP/ZVprU0Wtdb98kychOWHD9WB8Ue5hwpTOM1/9EJ/Pqn
CPNWdTaYk9pLJY5Oztea0OS8d1xD1gbFQx+A/eukZUKbhPzpP4cn6yb/7s8IHL9a
/HTLT59eBMw/Vz6cg7x503zn3Fno9zSmxr3qxBinMDcVPjWkFN7eLFNSP5WpoVfV
jQoBe98zu/SwlYZUYd7uQQADUExhJrQtrux1ArH1zE/pAFPAYGhWajqZDlqrRphW
/7wkKnHhO562/hQtLPv3CL9qI8/jsSTi2G9coYJD3jqEYCVm1IgJZrAA16edSufo
NT/9YUMnqC0a2s8+fbhmkRtusXRwug8P9bZ67EPScjbnNZyLtco8hZUnhXbo2shO
C7JrMmRgTdD85uZoyG3utyH2cIgN7PCdeS2p24WFwMhQi/qPmbLB7GUrX/sH83zR
WnkjrnXq5cuC6R8bk3grQx7VW7Ax4h5LSifhwc1Mr4g/56q7VRopCR4KiTrAg9c+
nXOxpEezMm1s5nuyHbmzdvTbMb9eUq1CCHy0buMde/1uZ53b6zNrUad2CokuoZQP
PT8EKR2nLX0JRg17WCsM2/tlAnAqsJukm7qVFxaNSuUjpkhs1OnYQKKf9juzKDpq
2ZraYB7dlpsUyQIFi0ZHculhZz9xrstJTIaTRMWHNzhxelFWw3PboLB1E98chPz2
UMb//VbhlUU1e39J4IwEThDionMZEw6ZmwLUFkKWeTJdQX1+j9+iWKjOn9m2bOyU
yLBEB87koggP1sjQMkc9QwOezYiOTgE0/LqJjKDgWmPatypGpGFZHXTWPtu37uo9
Dpv6+Ui9djCIFXJtSCei8jfp0AS+Wj+BSKgHmn1JDDkrD93AZ+ZHZ+JsA7+7wHZh
Lkfc6jctwkt//JMo58BLGxW72S+f8rnaTGKLyKrNh6oLoiVafCBbNX/awNPW/umL
CXccQgw3bz557DTqAIEyUDX6rK5ya8dOnDukHfJZWIC/BWWIsGP4ZUZjiFkmZ6T0
Ff9r/eoKfeARQxKugU51aS0CngaxfKxr25xN6/KjzJgl2aPiXW3HlAA+OOAy5+Nh
6pQ6c6fFQzoHi/hy5vqtKhxYh7vHLQIdaWqxKJNoBUczdb8gifWIgJNR8RGefi/C
zfEA5mdc7f+3eGFX5o9Yl1k4/4fuig+ZMCJ9D6V4zV7Excx5ujqPuEsMlSJdm5Xp
kzyV1vvU/zw83rCnrHUxVle7aNsrxpOp4+B7fMwN5P1e7+e119oCiaSnDnA1xm4y
Gyy3XA++Melc19pZkT19KxvmhgcTPFaOaL7rn968mk57+vbmuB8yJ29bZaGC53RM
IWwz1No0jmpNkUKDdht0MYks0izfJjraoIFz8uDSuUle07956PooEYbxj/n9F5V3
uA+nYftES9+v0nDX8Z6p6ySiThaZ+jj1/gEg5ZcP5wycGKtOdGOLRQbBSdwGFdzJ
lBZS5WYNwIPPEM+ZjrcIo04irUAcQbn+esUKBxTOX1Ub10/jfs3Xqvk2dSJhP9gK
J9xzBEVtUeVm+NSGkmtr+vIx90Jynh1vg9PA84ntxFESq2njUXgcXAIORFM4z1k6
qb61Z0XUb9Ql2dOn/pHbgRD+PFgZIGHSc27EW0F3PkphTSOfOWMd5Ou2qou4q5fT
ww60qu7EuPjqy1XNv4FwIVtx6ngDr0zIGrEY/lnSWsTE65OAhXIGvJ4g6FAF8HZD
ncB4vDDU2ZJS5luLG82p4aYfCv/pRnbqzJ88YEEmcaVjbTpeftxSeoP/HwaBZj2a
edPB0RvML86Ten6vecrGmaPdCAk5aZw7N3gC9nMCH4XJqge+uWvXmGLEszWYw6K7
GJoDGyraN9g16Zi72K5ojk9ObVM08yw0n7x8MQryHMeUckDYVu9fFDKjgmVkiq/Q
rCzSSRk7gtjc0sLEQKLwYQ0kd72dVPG06o2J56IJFpwM6B12bovk+B5n6Ksc9JYF
3hnrkLnSlHiQKBh6UDDxgH73cwJ+Zx5u/qNyY5jdNsT5+gyQMDJ31uKGogrPO0OP
nmOGDek4lhgq/BoJU0CwmfHTt9seoT9wdmMnW8jBUmqnwXOCGERkeSCei1tPpHk9
AKvgU3O0HOhIeh8hNHyKfUHW/JByGDhQi4jN95jI9pCX6i8IvvFfLIxViSDwHXtl
XNo69OCeAJ2bubzG6tp1cOc8mQDYlvPDlrufJlQOQELQh2eVf9KkopnYmVdNorJa
a/KYpDBet0wJf815LDbN/bnsjJVRBJPOPIqDdNeuh7VhIhxkU72C8994zHkpnCUy
kkO4SXEGxtWJqpKooXRUd+9AAGTcEQozoVBzHj4kCF01ESnE7gus74z0VaBW+Otn
Nh52SAqLLOaMP3SO74r1jZF4yAhDfE3ql4YZl5P48onimmXxuUskfumCgRDE4HEC
hB+YYqzVMV8wNAjmR9p7hKAd+k8Xd0lKqYtPxqa+6D2ouqMk4AuJ6SwhnCZOiszp
R/YN/y06AOYBxWA239ShlU6Z1CF2fkwk8C+SyhOObUUwOl3PsY8Zbi0cPIx9BBmj
ySXaAaQ8BaJIyXbkTxxeuk8cDsnvyIre6JphhkRKePnfANeLyAxPiwj6eFQvGFs3
zechks6FU+j0+yO1vT3f43eIoevQ9GiVnzCeUBnWZPbzuUz3+e0p/XS6XMZZ3nx9
ewRBsPybHu8MJfnVUzDOUlEZClvpTukDKiGW4TzhpRyvORcd27LokPKo0UejF8NR
Iv5dYm4wKALTSnFA7I2tqQ4dAPBVgcrtOoEz0AWVMsO33jzJ44ugk+H/gPfmHrqV
7wC2B8BZJI1bLlPyqX1hFEUR5Oh3AR6xsgroCssHSMaq97A80U9xPtSDSG8+FpxW
CKdhFN1QKt4gR6Pa/S62TVcdCw9qI+PqIg0rocNzdeijjEJdb29Wm0LqL0Gtvvmq
0jkYBG/UTJfgguzHUXeqTjE9GmrDMmwjn6SKQh6M6iTN/2sKmSYGZ8Dm6vW9YBpO
QOaBqTFOwwNilKkhMEYIeiFUl0qZYR9PwkiJoO62RN6F660gpcgP0K3zgOnQfs8Q
NsGT5QaxVGQ7z0/e90MwROSo/D+OLZmUcXC/F8PV28FHt5o2gK/BoGRTVAuxMnMZ
a5w+ivDcd0VXoJ5NBwiQ+dzbzdvQB/nuxKH3Z32Dh8S6ER35TBXsyFUoOHWcfPjQ
4KFi1SxxOgranAR/Jb2Mz3XrhphdmiB1Ajql85R9zoxFcW7TjuFqnvXAwlXUL99S
2lfPK73nahtyoVlR6L6/p+788PcoGntaElBOLbMjzMeOUggEF9XsRaaplD61eXDF
TyXAOvnfiGZYJMJSjQuGicYIJCOT97XukEAtb92oT3C1f3Ss7UzvS04s8camvboq
PnHSOHr5l6nHIci/cI7zH5nyOetGs6bmt0iQIQ+MQzrOfDlyYyiOMNtG1V6hXbIp
6cfwE8PvYipYR7qdGasSfhpjHMQHvDYCheEWnvr5SYz9ZsDoL6XNEE3vKWfgefcp
MnSlZ58tKoQskX3yhCGDjrVfhS5D5nNnTkEpJEdAOmeHFysf1H0t94Z3qKUe/eTJ
iFzoK29y6mh2zxUhpyTBX42DWQA+5T/dzCzUKdoXFbsK2lPufNr2SFW1JVRxMX2/
kix7b6Mg5FkW5JusXnEa6HdCf3EZxGXmWjySlpgc/fifx4Ab+KgDQ8F80fM6rxuO
HQr00BEXsgeJd8TJ6N0FNZ1GbXFvddKyx3ZOgqgM/6nhn5jQ0iNoEHFAkQp4A7+Y
yMUz8rsBTNADcU98es3Dq/gvP2o6b9Nd9ZqGpXr0GKnYymHeH6SeCRZV9fUI2SgX
lY/2uw+FS65YBSmVNGogBSSrq3YcP/U/gDUtL4ixipjDRnnQ6EGph68GwTsTRxtR
8IYAXayVRf68lqKmV3RPJCjXQh7rwJatXZbxdNvHQ/fShFmy5YydSz/Kz83T6pjm
2+BMp7XsA/F3jr5QqCGPGyz5aa4GT6FrfiHy2S4HmUHyadBsc7O0KmdR641e4Oys
fZ1bpT68nMAD/LIgl3Vz9GKtUMBPpnYxHMTuML//caFDFYWe0sSCMIHOQKJJQpLA
AGZnJZVGS4h7ljkbOjjywA6l3+4PLz8igPySVqVk8Uq5Mcen5MKLU8wQ4YBfIrec
s8dpH8Wbr4gTh5MhLWw0/0zuBWRHr8RwkZ80A4L9lPeypIxOkjFYOHoPSar+FZHd
69ARmpxVwTTQbpeu5iY0Q5sSWu7ege5R+roci1ZUxUXjuNn8c358fpeMirPVOX6n
T9MVOw1/rnf80KCnY2PvPKFNAtAVQemnxNf0q78YPE5XzK5OwPJNKd/xfXasjWZK
JbAVNm858lceUubj9hub31rpL0kit7jzyITny7E+uPDevAgELmzpjW2KAiCcMo2P
pe5+tiPL3v0+KW8vJ764O2C3Hq/H1Y4ynzqu4uQpFx2/l4P8qADJ8avAQO1Z3dRd
LaEhwO9OleZjbAnBKL5KD9iBOTuJmc2nmLpzeXDv2bzoHDzBBccp/raHBaWl9KwJ
VwCec0BqfPvFj+DBOm93Mskagq1gYsUXBCHwimgbXmABQfc0yLSy/VQmvhlst2LX
Kth4mLjG+EObooqn7Q9Ii0iaft4AS3YMRSaSlgXDx/Ubf1Q01+rpo9KNu391lUvs
md8hNxvHpIRD1GMMA2CKcomRarL/SRHb3x7/wJVsLHeH5Sk9dGYJFnINjRHwnKdc
FGGMHUZ0Ptp3Tdz9kY8bOWzetplb1w+qByS/XPsKzjcvORo8G8J7SPNTnXWxMiCE
IpoedIIj05JKT5Uhq61kidFeoMUUuGI3vcMlUnuSITx2xefokyIwDRthjfLn22qJ
YtGbr6b5DmqkMZr4jqxgUKO9Nea7xlSxWMQg++8OoJ5h0urUluRJ7i0IHwCnZAHy
Q6KgH3b4kDgQmmkMiZvrQ0K3GV7pfNPhNgVXLn27Jz3H3XCtkok58zQGxp//SUo6
ASEu1CeLqssJB0c0tpcG7YmMytuqxNit2bFtlS4MHWuxn9C4VOImtk+orDClsAPg
Lui2cJtqZLqnfyWfi4i+piyM+dzCMnpjopfIfgu7n3b7c6WH/ejmpUHaoXJB+v+0
ovTJithDbgJa3uiKJ60eyEHxMdrgIBTK+Y2OLqL4UXCvzgr6oYKMyrCyZh7+Hq8g
ToUnLakt0TsOTMNG4PN/wyjRPNy3Qqrig7oC4Ykq74SAZPrE5iJzqYYoVauv9aTP
IKvtxjiEtGbOPvO32yw/cpyo0ZSaiOcNVXk4vIUPj0k5ZvjYBIXetmdKJURkyfhC
RH7bCCKE0TiU288YJytxTZHhLFnpsd5DHsnXvyoC3iNa8jgbDlBI6cuQEJVVw9pN
N3+E8s+7GFDegrHDS6vlxT6TTJRs9XQ87kPC7ugBJvwMqRbkm6GwxuRpoyfVdDSZ
gZqsioDjoQCTdZnes6oZJY9MxJ4HgGYjxjBv7zrZ+CsvmdvkFcnKMiMwvB69wts3
20erVJ0BGXahHmUqC9WRPnLX+K2FYsXxEfBp1Jn8To0cw7NiEY0x51u/UwW0DKzZ
idDzbDwm2mtGKBi/O1MtLF2l5fXaEPYV8f2et3d24nHNQTJAuWNFCPTP+qKh7xTV
0fFRaJlTEL2pu9GGaOzaI7tTBz1jbLr6cIQqOveBmFfDbyxc1RK28Cc+LFJhjZ7N
RALS4kYSpvdgq+2GJoxKvlESfw4Ny1ROvgqP8qvQ6ihI1B0o5amT7ZKatkF1omMx
IrMnG72hDGkPTwbHZvmlfO38qS/EWEOhEkG3CVjBYieJs6sYS4MGvsuJrWWu+PKJ
vSt7hFe+GZzDl6ASEBzISYDuhug05KQZKfzqw+qM7PwvBEyJKi/7HoZtRFjto4QD
4yZBv8IjTR/nHlkMRUtYDnSRmPMncL8YkkU2n4f8c3uwiSvx05Vhw0pBUtnP+We/
xeblVC5bM/yk3dUpx1QFSMg0OB8JIjQ282hm+cZXtpoIjsXwJRfYKOTkVMxcl0cH
t6O2ifzw3x0zdLznsN9fVZrHfXjnMe7jDgx7aFX7PoiEfBHSUoTx3h809nveD6/h
t1xym+DPsLk679R6ta1BMiM8POHBJRg8dUmbn1SpgauSVAxyXhTCSkmmMvVYQx8f
QSd90mQF9AsXZbWYUq0tExdYkTdp+idJ/ZObttYIWGJ1EmojKrXnV8p4wwYfHRdV
tt0nUdBAnxsYmAeHOT9+uV4AtTm69VRUER7bT/zBzd83UlQ/FsUNqQUpYc6Jk02X
Xolm0aom5VqQiDsW+gPOwHO2QvN+T+VaqlCMejYgluZ6KBXW5zwAzR5sivtrzCd9
wCfbw1k1KKJ71DBD0Fc0z4Uc6cqTwAIpUAZ/FYyrClx/C19Fo7cS9GvWpy7Vyp2u
B0Tzeg3EgbM0HA9t6fuqJb4v0zxRgQAN/fgGx9rthFR4nhXrNljvUkSk0d6o7eFE
FirenOdeg8pj0MTa+/Brkm6bmMnrfQ0sw+q4Im2cfH4x/BOf22Efvro5fhvXX2uq
wE1/EV6RjiSo90Jo75sXKSB2bzaFY26aEykB1UUDBaJvkz2IgzVju3MpZou9zbV0
egqk4VvVTfH3eprzdEuE4v26+3nk6+Np5niVki7mAmKg9vlOB4TxRF5+Z/MbylPa
EqlsFSLOJ0jjdyV8vw6D+yjdeoTX1ZAcuNnoO4VXuR2tnljuD/T/AQ0Eb28jKhbS
7p3Qavx6oR+3k/C5X39NV0xV+pu1jkRCvlH+iAv2Azq/u0Hs7R531DlTp4G2W7ro
Xmd1E00ZIDth9VmoFX0fcfC2VqQdjs8uqZ1Xhg3xN/2WIcEhKUlRg0c8Q/VwF7qT
Yii0XolpDoeLT5AXTAXkfX0H/yI8yevwwJdL2+QMh7OXBa4So8VS81rxfH2XV8ZS
kVUl0gn/vnzaFjAYsc0771vGn2/9cgUR89tMaxU6Xx677yFQqBrycmHlPjbERdu5
+GT/DnCieA6MLrEiyWcVZdXEJZubp+VPWdKklYSRPHU5BkZGDzdOQ/DWE7oGLrNj
zmI0n8GYhxGjzbDUZPyYjKJx+SNgs8erOK1Vmqt5aHZ+WOiZr9hGqm9PAFf6UbFm
iYMhCxkrhGXIoYUMtsqRVui/iC4veujT2UWPcbS93FPAFqgOlM6/GLq7HBsGmn8d
RcqY8ethhvNXn3IiPf+3kUZY9HkGLchzsmIqu5/KS+y5S5Sig/uVnwMyiWMSd9st
Z4jce+UBOmEygz2iteCe8N9n29x/OgE2RMxIbrMHvtjmCJSGGR3u9S/Sd+jv5NQs
pz0KrJvn52pCoblvKZyGPRmtV1YkSx2U+iQAp4zQwXL5kvfSGPhJFqwIhSWGke/e
IBMjqb2AW8a8NAEsNylxYyrh5p619CMYLRq7cGyKUJKM1DdSfJhfmTnKxK6CfqBy
4LiyQ+zKiNWWJcq0TYUJGeAJJCB1uQtUEBedHSZLD4RMH/sNhTTlv0YGuteE6p14
t3J9ASqBl9IfZyfIjo3De24u1TcRtCISsvlTW8Q6qyJKoNe/TJ1Mvj2LF0LSYzRf
O+WxU2tyOx6wxT61b0al2grdSab+V+MmlbTY/gbmZ7RF9DxfLq6qqdzFLZ9Ni/Ge
MNBIdLgHr0Xzf+ZWKFrXFaPkL4/OyJBsDJ7sxZZnYKjrlrOZEeConVvROEvy3Fjg
rPCZ7YXTj/T5ZuXDeb73gPYOERiVLU5blz36tZAtIgOxgHuvtKfO2azH/TDqTtRd
orr8NLDRJkfJpzYSv+sN1/EjXEgiBTbsry/BKYounh0zfnmZPYCeVc1Oq8Uaa3Ly
HcAm20S61aOqfwUMJsor1+JUW67WJewEMtsmQWCF44qDHQeXK8IoXwQkt3UwRS4T
1sJXB9R57q0PJZBTJ9C0C59m0ZY96FHdo6ZO75mhQO4eDbyaeYrcsGwZLASOsRvX
RWenf7ba8h/sjAZM2pwC3/RieAGx6vi1SrMdHfl62nTW0oepnZWCfhwuXBNBE6GV
/bucGzZpCUBQLPqOLrsY7oNrdQPl88UF0NZfPdistweLda/+f5HgXpeSdqu3ddcI
NAxXNb6TFGchgw7nI3wreKudeoILvO4vayFkGjlOABSzK00Lv0cYNTbsQioli3Y8
e51iqWbkL+EdlzWNRDyRJs0u99s5ssTzuKKhkBVy6NoBqcwtSCPqRPvtk+dT0gj9
1xhHodSEcm6oJ9jdOBCv5Ae6F1p+WhTzASq9I+KdnHyO06YIfbIMqzppUHH79lew
fw7rkLKHp7OfZvOsgEixqEW7o4WLDF21/AMyRyBw4MCK9yQxRo9ByL5stgARTSwY
UuOzAz5LO/IIIj1qadBkdY7kzblud8ZoIDR6maNSISMkzbmc62/iXrtHK7uOcula
nHFl+qpETn6brykh5gFNCJnsydMRPaIp3rmsZeq+ZRrS/3KKyMbSTIDFvo0aoY3m
CLP7t3dK6On6uq1WBQU3dktwVPIB2czMAxJ/V/eOREqWB+SoyqrIEdnD68SOw+9Q
krtlMGEbfAaKDCncvlhJozETAo9IsZk8mVk3OOze6aJi/HOonE7giITqL92Yw6YZ
y9O62z+QjS5cMxP/WD/ALzYpzad8c6PrlI3RnjpXLfof8hMV6M1C9PFipTPzmsCT
rPXte3jU9BsEaFlI8IMLIq/AuxSUA0ZngE9hn48BXog61ANl/i2Jjty3ImAQDDNh
6fVZJis6WTCsShHge1YwCFAP8JBVT04v5SxKNG23UdieaczzMJT7542JLG4MIWQy
yJvMBonIY2/8vr5bZ4jPLNtBW56ianzarvFzRtrBOLHAkP1Uo2jHi4MCCpv8fhLE
TTOjHOVn/+kWLMwjTEoebtzLYxJTeX/EePel9WOFgbqAsHfUtzIF+E+1Eo5mz04b
e8cdvNlvKrD6SdibjPzZELvsVtfobpaxC2/++xxZ6I1okAxSqav2K0tLrryXnU+3
unzRViskA2hsJAz21KP9+kQKEpZ0BYRypfnp8pTLH7x2ki5LHDf9tZsSuqUUsI7V
OGejrH3p8yylR+c8JNS9tI99xme1AlFYWhMUNGuL/2MWYQ5R/BX6N+LYL416UOkk
gjlsWdbKcUNxl459eqhbb7b4NXtpdjV4k+1M2mQp9KeSYPeArkY5uiyE3cLK1MiJ
LhvtHDJ/FufzY/Qrb6X4fP/roEhf6nghs6MliV16mOA28qGHMijTNPcBZinlrtTG
KkXQYF5KWwH+jKDnEMHQJwyqB+s/mu2FsZR2T368k+tmb1gW8eM5A8e5gZStxShz
ACvOzZ4OlSfCmPiAg3pmmOitjkQmCk1HGkvLe4Swli4pZc2nNyMBMp8QaeCjOzCs
nwhg62K84sOYTmuG/qepT5kZgs3fAEmuyjaeiMQw2jHPxhL95KZph60yizWdl66s
JoCFJqS6VFhi7+uNob+mfknwCOYUoD56iLsGjCOuI9aKHXknuFMcL8SGZjDSzWiL
0Tsut9weU4M3UAhVPUhEK9VCC0jk34ObtBJhaGMAm+WWMxcx02IiBKN+qYie9fyy
h1sEVgUKUT/nF8n2pAL/skIcDSr+CGiNBEn+sfV1u4BoUmQ193sX5eFQwktq3J/v
q943sid4WAro4DIruVWJ5k75n7MkLGqa8GNMxiN467XSi8+q2lCVlwkNWMR00lEB
HVVrG6jgt4u0Jv9KnW1va+WF4LapscpWiVOWFeCjKGlxZwGrx69aHIqfEN+D7Gxi
92gFewJAaX/U7L+YMEwz/BwTR/xnc+NW3k64ZtZ9PKyPWzJelB+EjeoGk8kdDNxP
tXqq8mGLqtvd/no6toN4v9YyEL1BNzRVGvWRlczoDJ1X0CyAgG9M2FyYKtM47KFc
fyKtGq1oPYbRrKR8qTgyTmlalmhC4BTwdiNNa5tJsCouE/x3YoacQZMrDT7yQR4s
R561cAanxKLaWkXasks7XrQNvCcL/aGVYbL4I05PTEtyhD9ZJ5KJBbLI6DA+rVDU
QhpbKoRiaasfDXh2I5V/UhgwlYhz2YamrbRoNm5ujm7PzT3ATvLL+VyH0HpujFdX
YLIXC8fXJ8P38bm0gUbd83b225U6N8zBn5ibGiOzyTw6Dh3mhUgzIu6SGmtgvT8B
wHktpIPmniPzwzHOchjg4VMYfZvRfxl8M+m6O60BTx/O3E8GQJ/EyfTBVMh7D4Zo
w1GugwHrAl0z/9lgW5FfFKSB5ll/mDj9bg+IdX9NRe3Nq0A81jufazSpXHwL0jCc
P7MSxCcB5/gAevtm7s21yW0KoJMNS0/XZxpjmOdRLu4+CMvdQ3aniINFjYJy6Wqo
vj7ZewxFV2h0xRxtS0J0kNejINAOJ1j0YWdpJ2e/L3myLBueFhqXTyYtZcJ55BTe
oVFk/Rt44Qh+0aOhnDpIV+d39iJLzgk0CJUWou2rXDA5doKQ8ReKJcOhkICJkRxx
v7G/ueGJDXhFLmmixA+8SfwgLOb8gOsUDQNgNx8v06JIu/e5pQamgC2Wwg0nRr/u
VGdRrcCnirpzfZgjdSDJxNZ6COTCz87w0lf2mWPJNdPiVWFDzhCZFtpRm2Gwa234
3ijElGGuH5AoT9NZE8hgL9GoWQcpsYPqN6Bu2EvO6nQLy4Vkdko0QQJMZdUWCGEA
LEGG/wNpmjOffXoOxYhYeGEOxATuAO0zbuJE7ZFpNnwxOFgz2xTs/3FYLsa0MrKy
cxZ8TwKXy22w+B9Pmm59Jw4joEjmMCBZE5VwgP+WsKbySj2t8A3A3Sw1DFqCB2TK
UHQbdV4lijrwHAHLNgPK9tzKrOYZ72xzks0eZH3sFv6LyudBigtjLTMLR2cUGRQX
K/YXOLovLum8RDMcUDO6s9V/2CtCfRuR2YPmvcjBbLDPqagQJCOeKWX73/K9t/vP
MJPUpncoXG2azBR+TUrevnpbs3vsa9JIybyazxLuGcZaYbQllbgg5wmJfbpXGwD7
12kG9AYHPil1gcFlevdW368da1YwuDuN64XuEuVHMVAl9RNwC2m2aedI5o39Na/L
/aboU4wGUjgtWJUqp3+c/pfE+ptrMk97Bqhn4TFsJZnGZesHIof2Dp3Ne63f+4GD
QcA8tYHd1G85n1pHhILGqYJ11jAkNcNTe5dLr5TbfcWF4r0gioISSDQrAi9UVXNC
ypk4w+UXlDjNoRottx87EExkyJI3zVlQq77vqfHYfQ7tSh9Oz7A4asBsTOu6sDGD
3dHi2/jyhql6UqszjaWbTIVN+LKFdtm6NmTxBGJgwJmcGD+fQEAUu6oJVX3DQsPO
lkVPV27KiKxIqiC46fhvsDlS78p8lsAo9eyrqv65+enO+KcOdQLNztscu8F+CQ5q
lrd2Huk4KVAD9E5PjRohlE6TQgpR4zHgUVRUy5Dl2HHVf4aFB4HnrsiF+KXq4ZFM
IDPUvYtREywzVOj8at0VIkBeHkD+P+1zfv/lSUmFzwNaZ3zShxcoMSew5G6YYGLJ
DwxoaGkoELf5QAsd67uSQBrxITENQRDVzVOF9mdCUzXSYHHMaF6l8FmI+J/8REQF
rcyR8O264FY2IKCNl8RYnLPEgIUhqR4Dub6em7C8OV2bRrTPTsW0IWLiB8qB3orV
moT8c2krAccBBnCqamkk0IxUpGMyiYp/GxpH5cYITWRS05F94Btg6ErdW/XmlpJy
65cE29vwUd7Hgv44+yqFn8p18w8CLA7ymDDspkBsZbuXgy4bmeRzGDD4kB2v8NtV
U6p5zSPoXdtzcqVSrE34h8Sp0hB6v9aeCl2CsHZvUAPRWoNeXAHZBJeIlpIHTEj2
SlY0pEybqXdQVWOPziEuOMpSZ9Ff8OU3zEquz515Xdg+xUkttLzeYBgCcXjGFEWA
QE1A9FWUVucKtaywmjydZGxb+3gS79q3elc+NowklXbc99xY/PkysiuwqzDjTVfI
j32wpAq9qNQxAKw/UkS0A9SJVFOPcudYFQRiyaeTfuEjAERanmzCn8eu6qRqyuKq
c9kyHWNnea95n7bFm89/FeIi0DX+dWOBTIKb2PcE3WyWqhBXq3MEAn7SCCjqKdo6
7Q5eJE0CTUzfUpMF6agNpKtxueUxnXPnwzOsNgW5c9xGjVnXy1tmtImVu8mw+XE6
KDEnxtrfgl72/tJYC6IBkLv5WXepTqZBnpI2li0udb1qRc+Expjsot5oWQdLOyvb
Bhlj40aAC7MEZ+BcsUXphwYDL/gEQagChepHW0CmTvHjvmkeKWzQToOzKLQJaQNu
5f68JWjR2q5fz8l40zSIvtVavatj3JVhKIj1G5OOosUhiHXQ8XYC7cictpQtzbeO
Mz9IO1hmAP2rJBiS7c8Th0XFIvlkPjCdd+tbbqdv2FHxkSptwQ1FFq8RW8Dbd4HU
A/0lJpe2bj1yyJo2ZCPXypsaJ8bZcdwHwwLj499mk0nQWEmnYdYxKNn/Vx0glvmG
K0S9J1xfq0F161HWgufCgPqkQUTy2g5on9B/DCS5IpPdjag6TxIftZG2o5G6W40f
JW+ukzG8bJ02MjgEO7bTYyqBUmYTBy+Sc3haSADUuCMchXw5X1Ck7P9FP/nYdVZx
nwXETsuRsBHI9QbVFsLnJESaxdCvhabHJRMe4HUJ5cTpS51jCfZ9xAjVwjDO4uK5
JmdsioBQFjXs7Fj26vIcoUucdIOB1wfAlsjqeBg8li/rlcdBkKDujyrszcxDz+K/
BdfaUO5MGN4u3NtpAdtBSZ2tK//bhObFVeIZu0F+zVTp/V6fY2+mAzUh889c85tM
zvZ9Xt+Bg7g7mOUGQ+zQOK6zK4VMMKPMex/3K0ymEGljHXnW3mUJzUML/mlV6mNa
ty2kYn0w9MgB+XL4/ifSUvRWrGwyQvUwgzWoJBDkOcOtCEgPQITNpMG3B1GhxVqz
S6y7CrC9mvrITdEgir07gMAFT9+687hr7AkR6rz8vD99HIHZhN28k2h2XbF3BbaV
c+0hPsDu1VgjJOynsNFO36HKfUFpk4zANm1/rCsFDDuTsxKaaLEOSDhpZslHe2+Q
7Tcqd9hBA+gAg80SxvczKeXMWQKd2/sxXpTW/n3ZalcYWxxpFaQ0XT2VHCQoi35U
s2e31k2oZEFtI3Gx6ID4e75+Kaj5AZ0dyfnYRs5JSCiXh1X2WS+kkXzq3GQi/dfO
CVKIu0D883JnxtoDz3UA9xDkwsNYULhGg6cAuxJ1t5kmOyBfwDkuKwd/CM3hbY96
zV1nCycyRk3t6svPK5ccGUkMMfXoBnG9kTxo0UfG7jlgOWWhQ0gHQSA+xXnsaFKl
5k0oreyj82ftsFwvKF8dPVQ8x+/DSP3igm1AvLbDQtSA30amD39i3yOpCCGoLZH0
kSE524nQTc8GFoXIT3pGfdkd3FOxARS+42YIEKrr+j9B7wd5gSEvRIj7mRToeXZG
CUPjT0490n3oOwh/v69hf7CjwjxFbHrBvVVjiLQuiQDCuODnzLJm94PwB3Kiox8w
Xx6QqQ8df1fOqItuOEzvQe1MYcOsH+BPCvA69dnsiJCsmETvxuTKBei4+GgmfIFs
8WsFCNgNZUVSzLmEJRHDSLTJU4wuNl3mZ1Fk5lcuHbFFvpfa21QAVQtEsWE6935X
eIGL//4GwV4fbr8P/dXUsj/0EB6GT7Go5+kiO9cJycbS6+WOd83zi3bGs4shDmcE
/h5+ZZHxc+8kbVlF9cWa76GNVzPBPbP+A6Jz1s7/6YtJ+llWAdAO77R10Vwe58XM
piNUobeXFZsKDNXsEnsOTTRbBY2erd3iAkIVeTcVt0YyAp4046NHA16P8JAfa/U9
9hz+TvZM1+QNQjqYLQ7vxCHCiTm2Oi8sff+6ZI8C/W6AieBRj/8Ii/TfHYHzrVlz
0TWe6Qh715148/t94EL2FZ4FYglFQ9eS+5YF/n1hLNCSJPylAl7xVS/VtlLV1y6P
g1UYJdsVHIg5HN+SMTMeLZHCQ5P+6sK+GtaHkyZHgUIu1D5DwDV6l8WJ8h/dax9n
UNfSG9dAkllkjuo6M951UGYwh9DiCaGaJZXeu0uO5Y5oXS+iQjVkxIj1tWJ51wfp
LvFThsITOAH/6NFRASuL9zydduUTRJffbWG4hwijgAyHlCKaqLW82r4ccaDIm8Et
X55OsJ/J33TWKu+djLAUoHT3LXhIdeCRl9xzQGWXIb0XYoN/xe8EzRrk1OYOcm6V
EQnVwvYtYJPgiMibg0icUdelfUcXvsU/1Gv9Hlam1JKsUtVtxzQWff6nd8WYTYxA
of+R1Pkqi4Ckb8Ju3gTDtSHgFe5d9SU8vXMmPbusxOHCbj0rPY3Mj7fxj5Vqzbhn
6LNL0VRkMDHFIN5XZppK2BREk7WJvhV7HjI4DVCZlzlM0lKqWITLNPBugm2Ts8OZ
QKYVjQInW1Wc3URU2Vq0Gx1Dvi/5pBt4gi1W/CWAA3zx/t/lfHA8IoIVAfgEzhlD
j32c7E/5Wf0mwdKljY4nkFGslCtnMvtXpu9XFu6GPZc/tVCCco30uEAFE/RLfZER
LpFlEIRkrFP/iDNOln5mXk5raYk9txNRaMf4AvEcGLtqQ3UabxtNdx8MtK2JUve+
IUCPel0uD4HaIhcbL20ft27eVYxMMP0HWqaSSIlXjenRbYbaELfvX+JBCbqZiXzh
hEovh/fMYLGg+mLv9dKeMOtcVNynJtdPWeSDbRuDmOuATrjyNhFsf7PMI5XdZxsM
jjWZWBtG/hZc6TOZWHZ1E4g7WBCRwx0tqJAfQKUgjex4mYFimEcpDvrO9anc3PHd
f6rQx3Puot/yKgjY0jcER5HorfiZ2M4aw11SH7pCAJdKKbecV1zOAikbSC5tgFF+
jaC3kMfS1T3ZlvifJO+QosW083gKiP2dwAtaCHS1MqWZUn6clX8mB8KCEuKtn4mY
9vTwaMAjQygGZ3GWR+AciDfCadWFYGSbG0MzuCbnoN2P627l6Bd/t6VAskder3Rf
+4a/h7KCVjYFVGr+uQXHjlkhTXz1xb7uro+wsw2PM/fXoKq8MwHKUv+l9xvZo0QD
Iz41LNquGh4Ae2ZsymkrFWyuoifd6BPFVQZk5ZZ+xiRY0dZAwGDEvcWeCtgh9mgw
yeLKuudSPDdXzXpSEogpfW7OKfY6us73M7v7CA3q0Prvi+jlCNTdWnw0qMmghcmr
LP3n6IdU0L2KYNl5+ZwxYfU6g1GTDmEIGQqU6DcQM9LiE4b+u5uVxrevVdvx5cGo
H2V0YZmQAYZvePnVXQ58/Gl74rxEAmDZaQSmGYrPAFV9OHD095oVn0cY4enDAHme
uZ3inCMCzWRNBgDLDRwp5nRt9lLZKXBGGMyh3lgTPmcKsObYj9vz9qCosVTBUcEa
QSKPWO24rHQ1vmmWKgT4Y9cYCCCTly5cgW72uCKcxD2T3QoME7A5CYSMPS0FiL7e
FnoN3+3q4JsJT46H7ulSqEVLPEp9HP2JXLuqPINlAM6ey90XuDC4eF1EnovoKjCY
C695lVo/ZynR+JUWS9OmV+to6uuDiXaiDcAIQHwL93E2v45xhK05DqC14VNC70AH
9vAb8uTtCBA7vCBESvfTZYInqXT4AXNroyugyFWI0IxHrI2XMgdFLYmbd5VHDHEE
wnltFhpPw6wW6bDsxnbeMsAjNE/XIUZAc2fQPx6Va6jSV5Qt/sMQlMMmb3C6e7wG
SBlkxrZMfQIlIhhNP3klOPXbfZ/HaJakNquqCqJSMR+AEOU9Yucizh90QZjjKJv8
jwsSYAuFgyVtTDPEfvw0Iv6q49Clj2pb4DAYD6Y9Dp4UddeV15btxhRZb4GiwFPI
eWviOXt9rT++3lCWy4OUSzYYVfYh/V2E3nVEmV3KCPGzGcHXj/jbPNDZLbc26jv7
rJJnpjUHVTSFS12E50jAvO74yUKeBbqnV608+Lc1fV3OSsa0msvaQFowDalP+UJR
g7qhMVWkpJbgVjBV8Gk63uknsVc0e+9F3vGV92ylxyMog/3yryQR5Y+4/F2GHi3s
fbBfAU+a6YPKmsoiXID47hl4HA+eY3209Lp61EbYdqt7UX64hMJfUUR6Mf9+pNdM
qH1iIh2qLCvASqpYxyaar9lnIu28uhpJHDtP2M6oDmH7V1HYozR21VHBDfqsdc8t
pNr0HmZYS72V3OajtUDNHX3nEPirnDabN1qyJEyfFpG4vEVrU+1qCPOQTMtVJLqy
y0omTScdyjFoHutVriLNoFVK0JgmvE+QDrabKtIBcuAQxg9WxnbDMdr9iwUxYC3I
0YBLApVkgrLT+Z5/SKFOOARAMKIkDC5lLUEC0xHq+HcCvmFv0cjAPhzn7qMpk0E0
ufU0mBBBKnMmMYKWERausZQy6h1U6tcufUOefY1MWCoaLao0x/4LwsXS1Pyi/6rv
aYDr6+G3Hf6vo8MGb67OCY4JQmheH9d3Z2LCVdraEKdk3RjBzEkxhhPgCPc05COM
E0oaQyG0pUqWNDeCE2OiewGusxAZusCDn3EBs58PiOrHIKU78tWeaaspr1oEngDh
u0w82x488tocgw/QAH8y2QP6gHwLcLasMp8wmy5w3aMyG0IcVk83W8TekEMBtmCw
h+yu0Q8d1hkSJ3X0h9dubqPfW5DTYXqRINBJJH89Insfj01lWKF7KPgk9cNRSX9T
miNM+oIE2kv7auS3hLwYzaANCYQ+vOw1C/T3cmkY1htNebiUZj9ciBPHrIIxV5ow
L76h/ajHwN9/74J7JRLU9G/jNhtLyPIBB27hG3u5bxgyrAQyGPWgLBH47QZ4nzny
KHY/cEkYXxeSdv+4DGDkcWEOkPTGmZz2Wkg2Wb3yU69HjbhaKQzxC62t1V3QH9Cr
JRpG/PlxgoxdhKXxfmTrkOw+Bfy0PwfIphqPXP9tpY6HX/cCZLwCYNA4qXv0m5dP
rxxatKcOitjqC5T0aZ9K3j5IEj6nAK6lvJjOsTIWktoT8GtF/+pQrIanJJDmQ0zc
tq0FW33sC2e9KV2RiF7sUZl4hoTK8GF5wbNHbYad2jqfxFZncfIPvXS8yUXfpBzp
I5LbxiTI4i4HWj7ZPjl+ysivJ280nC2GWXVfEdpE7DrOsDpTU+CQHk6Ud63G3fcf
ECB+X6p6MN3nziqDBXkhTcXw9LJitjO1/oB7TdeSPT6Ml1/CbuacqYVgEw2DZXYy
l7W9JW3wVbztfnR/BiELlxE+KpExRl1rUwxeaFA8/5XQUMOWfKPCWHp6NnuYjJYF
8X2qEgIA0v7p6d79I0N1UWSeN83zOKcKHPRKSyxp9OZz88YoXU3y6pngqgfuK16A
Q21EQhVwQMwjo0p7GTogJ8YoxialkSzI4rb2fIrTMB0qR0iE9AUCmzU//XfpQTJi
yOJdG/EMVQxjrr4zoQlyd3JiEBqfOj4DofJ1xR7wITy8RN3dxsniI34fj/4yFFu9
Er+HV9jWv/edvWlovIobBwChTbz0TEdc3eiH7zHQ07EopiPAGRCQz5Hp7l5K3XIN
5KylHXW+mphucrbnSyZLTzAlck51ZsQJE2QoWUriAC/bubtth9j88Oerh83jLib/
BxxRB3lRA1J4S2G5DmaX3+JHxE3tEEPJptDLAAM/vJ0IEVlRiKioS1EMJ3+rkh/k
QL1hrGcI9qmjsk8tDtpdQGybJozO1taSb8PK3q/l9vDoLyPyp53JRrpIAihgBarH
Xnesi/d22DgHmS8qObFP41awoKNIE2N8nKsN24cpmaXKx23uEpxz7VIq1lrpZzmB
46uzLjyppXWAvP4UXGu8/Pg5yEZ64agZxHnmgfCHl9XJnnTgGDtfpenqlaA9YXWN
NzalHH+uP7z84Ny0IugID/VW/fLYMrrMGansu8Tbw5boOrSyksDR4J8pQtlPtpgA
IhPSD31sXu1svlqzR1NXeDC9cMalyCl8ZRxc26oubwHqwZycNGt7zz6U9llM/H6A
T0VMrIdcWQ4yom3AJDHo/BuxbIcRXH4hiA2LC3oXelvDfUw0DeLOfDwV+3ZgIKAK
xYnjK/1LhIL9BrPnIhrxNmHHK1qfZA0oS9L+JtEClWrxnvOA7MLG4vxYRsXIn9LD
BVnQ5rCZ1ot5Di+6VJesYL3A7SurYRytjklDLx/YtezEr305neBU2Snja8tYf/MJ
9SHoZq0+7hRyTurGnoL6X1F/9rue+1jNcPaQPdn9WAbHlCZ596KL/EdysWAkzVUI
K/oABcWaaAphUoe0AfzVLEZEtSYoJr6nv1Y8Z2hTfXojDZXLs4k92tQQzvaj67zJ
lXd54mp0K9p9rqTuf5YDbGI6LjROO2devMtAzUojlP/xyQb/z559j/I/EPMhytVH
/5Wz4BnEgCODAps3xK7QGF/8h2tm+fItohT6OoTeOKEFdJbdA5irVfV8W0cnNJTY
6W6xULbKDgSwOOTm3H7QIRhIlFEwz0mAx/+p8KJ2wkxU0bdcVTXNcAUEUnR976V2
emPoHsoCcTBPWdIxt0uuYunBTnFs+SL7V2GzTi+/Qsv3cDA2A4x9Netq8iqmk577
JFOeaUNyw/Tkg4Fmdph6WT/ScSCDvWP3mBi9L3s42adqVW0WL8BS20aZdhA9RBwV
mLUImKXFGaCBMyQDxD400O1JiYtTw4PG2rzuCfmxas61jcEo0he5WFx3NYSWbVpB
GHSFzSg+Ra7mPMt3ekKedN7jjBAHlaoLN7IWGt5QKAWDpstv8H2jqdZfM3vs91lr
zEOdX50HGGIrL3xyCIxfQr3dUXanz5OBJRf7ALtqMjcT5lp1+GSqX2iNkdaB6aCL
BYg/F7kP0/7+g4h5vnKXGnuGj9pbkZCmuJHfmqF37B6EAEi1TA+8Uyn1qWF/kFh0
aUsxeJoXD1rg97g40zLxFZe9LgHimFxGBdC82MXpNMKbSWw9t13hKuMnb1hcj2QA
YMAHw7GnSHoHbaZXtj+fv4jmJf7U1u37ZRV9FAv7Z62onzo5YSIphWbIxBmG3NK4
eplzu6ioxIEs/Fr9chAOVqs0ayCXBg9gqNhrQAwdOJmU3hJ/3jBpoEDCSRCl7ceS
FDxB79XlxRvcWP1KetmMQTrBX8o6tKhA7xoZYhAJQ6zBlBCwIeZlUlpnAHHAtuh0
z+cls2fJ8Je/NbC26Sb+7ihTnCykjxj/+pKcC4ryIfpe40JyzhbGzQEVp4i1S23y
YHR8guhd4U2tG4W2i5ptW8fjyeKLd8S02x3VtnGU28Dpc4FCiPch/AMyP12tNoEf
Eddkcd0oX4s1ADMzHl7EGLwas+C3iqDvLh1E4oCYExASOrAAaQ5imja5I0NnsRuV
19P7HuFVyApoPXtJF2uXCjI8nreo+8ekyYPW3NwtyJd1Ts+qmXms016bCBS6UhxG
YzZ+Om+0MBxdAta1reXIestnp4C+vWB6xCgTKRMDOJAEzufkqVbdy06jVLWsdPMZ
JxKwrEpFphvUGvqs2DQpgQyjgvka7AnsVxpkAfmAwyOXoL0OZHyCueu8xThqr8IJ
AJ75PQvcvon5UECS0/Wp3u2xo88aO/jVC/dDoqRaYgbafG/SIbCElLzSj4bBgh2/
b07P573qBgzYNZNThzEKkCsWDJbFSdPBtiq/CE7itTlaN0lEwSxTyYQnJikXIiAN
VDNCKvHrs0ZpGd1Fd7BxrsZO05LVvjblYo3Y6Qp0FoSeAqox35iuYUw6duP8gtV9
trMljlF+iilIGbVPulwD2kLLdTx6Df0TJFzrPafA5Zpdibqj8PkulrBRJ7Gilx+4
mAgKtw1y1ZQRUffZG36XMZjsHeiE8DtBnUGY0oZd+w4Cd6z8RCSkJphG2pYeNo5V
ktmQ+b9ui3GxLVrQOec+aIjlzlKtyIrL/INT20wIrTm2JYjQLVBT5zTok7DF2kPM
zwBj8z3hpH73jTnbOvPOeS//rSWotrKMlxNJqF7hJnJgJUSYckqW5XMLXFBvUOMH
EpLXORBdge9KSyG+Vtux+ZnrLugj8jxGCxF0ya6Y/Aiq7bo5+iczYddcEAJ/DJMD
lM1EgrL75ZQP/aWW2OEbGxtpeYvHl/X+fa8dO/SXVoZxuMks4ZU8b20KATYKsFb1
ORgL9WxP4grljd2jQPBGMqfb28NWTNfAfub1mY5iFmoxiYDyPKvpUmGkCqZJeic/
tXsRS2nA8xA4W4zUnI/WLyfMaY2DgxH1yQYNy+4xnxZnqv5eaHbO8xF5xeL7fE7k
fMrIW2slkNtAJnQeWzBsRFCJt9y/VRWLRyTnFzKwQBpKzPI4xuniTnnlSzOROYzz
iYlRp5cNbT9TWgts9nzJDMe1AZkHEe/TmsJnlPxQAeb68hS5YsNnyk01cXXNgj+l
yFnMdW3TYcovnRhEAEXODm4Nyrig38t7a95DyT6+ZrUPH9rXZjIvKXk1pC0DBxwh
YJcOQynUrLEgUYbl3+Es08LdzyUuAwQGBbmetvIZpf1m5LvEEJ+i4kwrNze65Caf
6Q4QFG7m7nkktuVMV5oIU69nhggtuu8nhvGo6PNYfMU4rbIkYznkXlSRgCsyELWW
6B1ufrrpvah9yQNcllqBrbG7rQMtqmYjVjgyHZorFyKpSt7s6MVJFrsxnWwZFQwR
r2nUBIcrhXZv2X9OlxKSbP1H0EtWoo7duGRoPgQFyb1k/p4E90IcVWQkdo5UR1dk
JY4d77KO0EsD7I2yjN94Y7bCrWFt3a8J9DWLBup/87/h0/s0Cb/CwiesW7S16JHK
d/O3h9kaQSJ2yalxSeAEJlGZsIsXI1aKdBDRpjmlG00ePXjziCGwvIVMYHxBngQk
XOLdCP2xtaaJ1w6yzdND7Ui5KlKzvIADK0sWkJUM0CjZGiXEqLx12eYIqkxx0tdU
0hjNpnKfX00poSmUTn+sgybkb2PNSzqbevgKmt7PJbmH+GV8C2wbnMAejYHniI13
ohkk7GqwQn/7WZWRmUniOd5FmMja1+JZw2nSg43tu5NNryaKY/T+pRwZ3qX1tvAx
6in9VzRDdyLt3G7b+pGkcjmsp02TG/6X89eL8Cy4kZhSG2kyjOOT8/tEPWFqWZOf
ZzlC+m8verimsxm3/zgCGTE7sxlEljUP/V6A2ssFkNuvsxXeot0RMU0f2K2l5FGb
O2cF9iM6+dCtmR4oMRnmE8vLpOHojIN4YLXSw2j4k7j7j/wfKb6xpnvrbVX2p3Ms
oxqddv781z+TldRW052UurC0nyTNmGNpT518YWk/GAqG4RxVftf5pJltFk0IIsb7
4Ye7O9AR3WHuWa5WJLuI+LTRlWFLpCIzEhgwRkR2UaVkaKmbSHFXplEdubvWaz8M
B8MvpPAGgJz/pzN8sh4weSNlPtVfu+uXbW+daVGaP39HmsV20YE8Rik4QPbFdd2A
AIe3tVu/A11TY6UhTIm+Rn6OypDCsFeB9AQGMPk70uwCq3s9dX8xAboePAKRGev7
9ILbR6WUSL1j59pUDadPAGyT4QT9pPtIgb/cWjTouOpL5Q0bGT02Zik1LjzlJI1E
K0rPVRhWCnQTOCZEEuYBj/Zt5T8HgNj3VgLqzYZmWJ0IFPXURPjzLWEUhYJ4xDI3
JhFEXRYpgPlRx/cOdlsMB7amA3o1dPx8a5w84/c2jc6ZlRVzPKQqdygSAFaQvwFy
hr0t97t8c0PBrLPYpC/zsKSr8vLqZe+DxPMPjk/7xhbJ+/WmBcZT/1utaN+y1G+3
X38TaUxWuV0bvQuzZuUXWCfjqwS0XOY8a0nOwEbXW6slQE8jRjepxQxh8C1TEfnp
7ac0ig8Y6wVT7y89B4VFXqLMHNQxUmg35SYG0+l+n7YDcilw0BRIJB8KViMlk89M
L5hchYzcbzC3xhI/bl3QeXlgGfXqlYbLcUdFU9z3WPNLml2ofTpImIm32x2w1v3g
9G47JBt8vHyjNY/VMuasNXuuuC553ii3i2kajs6aAuZtlklonfCV8BfEZ7VebZnC
faaWKDd3JFVPrZKQz0ghjkXVDB+Zmen5qTRfd9KZLZIkRFudTHAYSEAmKbBQVPAd
SXL7CzPP5pJD36ZGAhfBwPsaUbAEJrfsBBiWlJ5TmW8RDMiZ8VGXJwKKwDGqNdV3
58SyXiXYERSSFiB+4GCZd6TjdvFhdUn8ynYm+8Np/1G2xgCjYRuiQDPIsqb6nApj
wtFGo5Pr746B2w6HMrXY713s/W1E8BxlPWbvaYSyqNAeM8Q/tAf6aI4MSyjBWHRI
0NsRgounAC0IOoh3Ao/CS4Jqb8ANM7O3wNh3GArg9wbO2tnIcjWoJaHws6obxWaT
+e0p3DFpaw3CDnQi+JBJI0B1sa/tBxdvE2GX/gdwpc0DPCWDBKGeZp0VWyOP+OJy
9Zu5NgxyI63EyZ1GHyALRvyTZGXhDM5p7ArQ7YE5xLfg6iJeV1PEgWaqONqJghT6
Aft6wqaillf3x9rH3rWpIhfnTYr71iPkHdnhuqYrdpfXtRTfO2a0U0QC+OGZETgI
u2UDc12Fom4oB6VjVx9nECBER+u5JNziv92FqF+iTJmPceD1D6CkU6HfhpZ1OiuJ
SU+hYF4KhxheS1Sy7r6XWMLMqDaIVWbhGZ5Y6LD7b82NaQ4vFK/XQatd4FYufO0T
bPAbfEXDXV9XbTBb+N4hC4QemhkFbPR+Ulz71d/80RJ9L1A99fzUo9EBQS0kZFS2
4QygcZ+STWhyXzUdWgKcCBZpkeZjH3KMjOgr0BmuFI3EP4+4IFOMOQuo3BRYBtBW
kr6FLFM46uwsFHjYeeKPZEeBPzOibFI8bLFbfm4f8HhlahHbgT8T0urZSQ+21E2X
jimQl0N3AowAzGp5PpM6nby9Z+7qtypgmCj+9dUq0w7LE9xcmZ5h2of3VXLX8FEH
c4V4DZSM9C5EXgeDF8bGdplv6LxFzYobUS2iDF+DvlBUkVfbkIV0oZoLO+U4t97g
RL1T4OCbv2YpKNOfHJk6ZOk3zYsVyLJ1DVww/yb9M8ZFgqGcb3+37e/hLJp20ixV
l92fihyFN7WJ/s1Kohu6/8aaswxXqd48nFRCC/xyzHKGuqHiA5FpDhIgwtHUZGTH
rsWfkPJPAJvtdEzSljptRaYSjxWni/r/j4rvSlO5jzy4t/JjNgZi46fE4zKFJw8z
mKr/S705Dwf14UbXi7XRvsh9ZurNS3Iphan5BO1bdrictPxylAkDqjq8fuy9DWx0
rSR8DgyPUqrA0aCr/DD4UGpYCR+s1ftYsqwoUZkNqrU4K6eg8bz2ntNtzfUc9+Ae
wDqJLorD6MS8RVzym2EMIpC1le8QrI7ow4zRPt0UkzMdqUDs2ij9SIr3wzL3Vl75
2N6IYYzeYBoUqw7Rofn6TMBuR0AJ220Z+wQ6jot5uXnCNvSNr8LBdNCP4ePKOU94
vXW6vetghbHLjEOwBLJUREWydR4vmY5iDZaYPVQP6ppRuJ6rOSUjMYtkPiXGEZmL
rf6eEaXjO1yqA4vbSgJdODMBiXrx7NNETKh1sy5chufQP6wznL0sRuNF2+zAsRgi
nzyUS+VeDK5J3paeZ6+VsfI1vjnvjyF0yvcCyFiCRhl1/2QSA4a4oJa2AxyFXh7J
VARA6ofJbTNOpMCq2BUGcCzbZstMv/HImoHRCl3viy63xpFYV1MtnCgCMcGEC7Im
0XjHwY7/4q0rHhfYe3O2s1Yy9qZ3m695FfCqbLSgoJEeXujLH1H0vft9+HT29STV
EOyklY0uEb8y9eLtOO+IgyPCmDNxu4NTyI4/BavmdwV9d75Fq8KsnIpHBtQGNtk2
vPwyi0SC4+sQZVPe3v9i01C0fSJ2gAIP3+EXkxy2nL+0imuaOLoNm8nOh0198Lmd
A0/sBiw1N+rS4WVrShUMocGW/d4c54nmRooAeZ7YG+eqGEWw2zbCtWE54Zf4wuY8
1DzheQDLprZoJon3B+lFtRZd32RMhkR6gL/Bm/fesForQw+jIbr6TBICld0xTwPM
8wWcxK4iXsBaFH2tyG+XCxZ3qkk+fqVYyeCQF0enOfAFdAqpl2fu2BYINbtO+AkH
WuGMqvCgUkwtdsaReT0Eswg9qy+6XtpPZ/fd/H1nacQh/NgrkvC6A2ZEU6avTp5W
HQvSA56pp7l9vMSVmF8gkXlv9456fV0RdSRw1zz2mBZOIsxtKDZ0UVtrwWPHG8JX
HliWI811n8r9bSHRgTC1+yJ1VsVRLrWDQAxyQxnoz3pa7FzM+kapNKwgF70gRQZI
DNJsL0nU0Z8yNuq32FIqjOXoW0D+LLffCPcloJrTlQuuDTdPxQcuKSICFUBabwXZ
vI0jqugoEOGZkz2FYuoxgeQDwTMXJVa37oT9H8i/dcFddrDvsoLr4bnketvfSAP7
g9NU7V0j3+NZ5JqLAEW2uiYHWO/KyBNXa8UhL5aDc+sprSFAuE6ibUpJFc2dKahf
B/sZkO3zjyuecAHpe3HSFhdqFyg+22hmLXY/STam7oI1k1STURguNQySkHZtDH6A
SCWZyA5EAoGBVGpKdDAWg2HYli1+5HmEfXxmPkvAdMrNJDFCFsdsO5Dc+YxeHDOF
g34R0PmCXOeJjEEboNs1xb0zVz3wXXfrQHO6SE/aMdTzOQQZldFPE+46HGiUe2mY
mjuJ8YWx2fDmcn7AZlASAHiNz5QAZr48tPksg1wMfqb42W102KHGB13jXj7rkcKp
yPgeFvvQnf4y3e0Dlc70jElFo6DaOhdJVWn5Dz7IolubBgYutTteB17NIIVv6H5r
Ad1wdr0jx6Hh6NpppOxKWoilWmPOYEn+uUATzSK3eZD4mDxtoGX/3d5scTL7eMIf
nvHkPBqPpxHsoae1p645UMxpArnzR5OZjtr8QJVpycg/4gM4E8Sq/VnpfJGuP65n
QyUuhsK2gsydQLCtKFX+1HkN69m6jcgHDAMrCi9Z+jiWCVX7xe/s04YGNLG46OIK
FB/IJRiUuqyAvoMjdzlddVtK3EM+nSxtI4uUzo/zIYSeOgTP2QoGgEOebBm/b4tF
l42S6JkjuXVs2s8tlIPLWR5GDlsTlTU1lU9FLT0MJfvULec3zBvmOgx6ryxponHr
GmX0tYAbAuIRPOMW1zTL2rBP84A7myLxc3fIRfoY84FB+SUgOAxBvprR8DR4Q3Yd
wH8lstGW7R2CKtOuVuVZmgPT2qnIVrD3PR7Ivf6pD51Lv1DjEZHDvg8szXALcWRS
w1yQWbDqd5HxIH31hdXRm4TlvMrFPaGVGgN2iv8iBmRkP0s8xwbxIkTfDFB0AtE9
s61k5xIzADjFHe+Bn27Dc9q9N0BB56IcYvcLjnb+t7AAzc1Lbi+bLbyO1NjjnGHb
nlRIgxNHfDWkGwAgZCn4W+5RpxCkSXyT58dt1PxghdVBsTakdDPjIlb60Cq7Itvz
Eko6AkPnskLrQhHpcsA59f2jwCTdO6fTBFClwFYWSiYkb8YyS7bFbiBVi2yjEqoX
SK2FcVO4eDYwVqNBO5AzLjJ1wvmjeNG5ldXBBrN18sXo0bVJggnrxU84csCo1Aqz
whgexkmNtyFdTxzOv2te2SOAyi2fEsTWZ/4mT5KLiru9BBsoMfgMAabh3lC/6XnM
UlNmaLvbj2v5WsWlv1rcJoyYiwSi7gsFBv8RPJohNTE6Rl1IOD3XHC7zdEd2FyAy
o5ThoWwEdNM0p9z8XPfn91wp1Q9HwT+ZaTs/Lw13x48sgJR0vuKFzAMHmFvyqKAY
32RUOKEqvskxlFNWdS7YNYOrfXm8JBkGiXpvKhCcXdDCuBn6Vxa9jCsXNzY4EXqa
cCXwJyp8jRLjBQoo4IcXfXxY70SAc8wKYDEuo/ZTzeDmcI0TjEt/6gTJYBw5ohek
exe0CdtOKjZbxGEUoEmKFJy8fKC3Q3P8ZIJJy05McCXIbO4/KLz91fFymltP+jmc
ea519JH+/NO9wjnCy52atAhze3poMAexy/ktrGhhRXRC2nORX1Re84ytuf2tipzu
e5B04lAPoXPcuPGLalhMFQt4pjkrEHF1QysBgRXIyw9nvYCA1YeVPN/AR9D/WNky
Yyt6yFdXnQys3cNd/6mOJlw6at10Iqbcu8tYXyCC0eazph4koFBanJRMnkaiMXkj
TI40bNaSRCu5hcQshv4Cufn+2EaAKtW4DBHkJngiBotMDUyPHnfq2UlQD7lc6Ec5
poTm9RpOGLURjR4tzFmmMthHvdGNo/YAqewALmv0aa9CwH2eIlxE8O1gCExwH3j3
/7jWPuLmlrudtqbO4Urax/MsyffRHWdfJ53016TGb+U4jUYmiGKBPXypX6Q3kfPG
Kid2CAJP71e9n9Qd1EvaVeNFTMYM2H+dixmM09gtB4oH93OM6qpi31Ia9NSO1+Eb
Zs2os+m0pd7hqyww6/FNb9QBiEgt5+lQcUI+/ElF0gSiRnnf+sMnNw2O8k0D+Lr3
EZSxomaHQITlx2+rYYuNrJl8MwXKa2RDeOLsuCLZDlXm2O0IV5iFtLJcfD8WRm/a
t59nfNGDMWlTdrQTT80ILkKtAQ81G1F0HUTR4dRPX052yxQyWIXhcaozOa5KDslT
YTw2fPQ+CERMWnwApzTstrzM+PjnM4jNYRCgbrAwMXrfPMTfx3dX6ABVN+MEts7C
ynUnLkP1QD+ayxIHupYUKfuskv+zPief/hOonPhJ/yGETnXBoEH6Yyu7ixYBzmpX
xi0e5/M0i2JMorVxmAZbiGGQltph+g2TVvSaUeOCzNh2my1muEcQMTWAj9kTOiJN
oAKgkwxRBNCUc3bSv5MgA4Dbmj3N0iytp7dp6uaVjrsaIWFKXna1mCJftVuYUBSD
BYPE0ie99gRRAfz3Hr23Np+06ZW1SEck6dfxTczAKDXYX2FrZDjseS/ldF7EZWzY
BkcZT0gaIyiqT7oKM/VDI0l2EiufwUtG4BM613KLP2ifi3y5G2sFcrEuPd5loQ4j
iu6e9iho7JndGmzHjB5QRUbCgjjmyfEbiIaoYnz+7CmeSyS+u0Uw5oxyzie5X8cA
NH7TybLMUsi85MT4EY0TuzMdWNTUIKVycJRtoPs9Ym5kDwyiuKOE54F9wJbdzHvi
O8P1nWmyZvzfmHwjLMI1+HBMaQ7LY7qdtFLeYGNqp+FeNmi1q34Btf4LZn74cKwI
fJEWehApHfL9rrOyGh1KoujGQtnH0JJEVEAtJEyTap0KPXIbeAZsh72XtSK+CsJG
gqTzlwzCnYBwRQ7xnB6VdnCPSv9KhvTvVxCq67xFI328TNRpqxIWFzQjkyKvmyNi
x92bRvw1AcSXLxZcjGfgMD5VSFl4+7fwpqL2mQQb1Iwjm9p/vmlHcAM4dfxqIDli
9kwdYzltFrcddrL8MJCenGfrMjUHdXJSoYQHJP8xQwri8yxsFpsxLREVdzXI5Lo9
ETeNTi2aWr4vTCIuWvfmfVJ5Py64wilIb8ZSqdliTy5BKpD6hOs89uRU7ZJ3DriS
h9JDct+Taw1KZgSCp0SzfISxtcPTXHDnw/pb8746BNXkuHRaYUecPfSDeXwovjxa
XkjgK5XmXTEATZVIHFE18Xb0zTjN154pux4xBghjy6NutOLIUnSJ1+jX/JXmeFT8
VZWb0LtxwLCfXWQjseB4ybsa+EYPSksxXqzfsSmuWZP/DifZAhn89dhgzx4BXMd4
Q9Un1XQ+f155Tsd2KRbh6rwWEvJEcwpB9zSGox8780MbtESv2UrwVl7yvC8Jv7rr
Sw9/+EHrlkKIQX4xblzmHQ6U23Z4jK1+tBL3dlpbyWczQGu+3RSsGj7XC7jDjr1q
qpwNdDhAN7r5TxSHByC2a7CZr/PeqopsT4D6U9R4FBN3ypjlBgfYTfrsQdB1CLCC
TfsKYwrHjyNNfpgu1m/TIDHY1YH4O4Vce60ZU8ChZIRoZvKWfCNGCkbunFMqjwyT
EO1hhtEZoszdvuV98cXqvNOmXev5rFgyKSmQx0ZvIJ26RTdMrkOjOBKE1zCgh+Lf
AsTF1QSRq6jRNxBhQco/jJ4nuqDJsq2Bf6jherAw3Ixl2wf18vtz77jZ5qS7Wy01
uk0pmqjQsEoTK0zv9hd0lsLsXtdErUvexDYP8eQcw5REtbqQIoZv1jl2OmuzQGNa
toTAw4OFr0JbmCAaS+iD03eqmaGInvj9JENbj7yTYcHBzedE9bGlqWhiQnQCqjax
nySNOum2jYDC+AbFkh45WZD77jnLp4evKdWUGkTnG+FNHLbyI0qpJuEKCERZ5KPk
7c87Nz88P84sC+VphdymiUKpC0MkoXp7GP7NPGqY0pO7QewkTxvQa6HCsvtQXrdT
cko1qeXGWHvstiYjosD/z4DGnRT+6oFZHHCp4MP41sCYQmKhYDVmbZxN7WvZNahg
gL0IO+dI/HUgW+3sfCvkokQuRVB9fBjRLOYPi5EOHylKWsFgwco4JrGzUPWVLBAE
1WHogbQ2RpGypQepi12e1rnpPdT1eUoHD8Kje099qjrKgwzkLpMEFmoX0ww4EYXp
Dg+gFxhdsryCU6KOBC+lkWs8P5ppMXmW4052iTY4Wy9//AEr6gxoY9ZFDIknaKuu
vEiEBV85ofzGY5oJg487isgt9HjkxC7HQ5pNMENn8+gajrB2JBfxoM2p/N69unR8
6v2A46TNpGUfAGws9DhZa3jnTd9EIT7mxhh8CCNSe0iFHDmnWInwviTdu2BoPfY7
FNK0ByufJ2ZpWyrwueorpjW0yWqrfnXvI7Dt88p8mDDS/IA09dIwH6sLDm72t72e
5AiAzYfHaQ5ahE+2U6bRZnWzS2ijjDOL0Xp9ZoOBgvvcHJKTYts+ntfjXqkHTOvR
m6i0qKTnlTY9I7iRphl+qKTv4F+Zt6g99+NJMTnNWq1PYWZVA16jkaH5+eG8fQ9s
zkfhaZWelbUB3x+PaWyrt7sZqQiT+ET6FVvc0ApU8Bl7iFQfTGPrBoLhE+/jwsxc
QHESWbiAb6uGqLqo9jbm3uEz3tnsfOrOrTOEAtYBGybbamclKJuar0UKCJTgnaZx
pC1x/nEiBWnQwhxVabuuHpUb/eMD962bkB04TcylxS0yp0qokolZ1MNhUvDfbzaj
WHrezbhYBr6vpnkc9JiYQUgbeLYZrP3Ge0VrG+d+yg+sVnEB8ONICLesN2NAMPK7
jhO8PdGXNdj7quyS2TjxQAN9tXQ7fHO0rjxlQG0tnDSTei82fKJu4ibpm1fGiQXR
bdHfZmIv00TzUmpF+JFGe6UJoPvN138Xlssj8ysWIpX5ukAcPBKG6eXbI/fto559
p979Kkq9hOcBuQWdn46gDqNwuc5t1EsBPgq+tXGXLi4yAT/7llKduUMLw5jbaEnb
yRnRf8uxUvvbR69Nsl9K5/BtQtLjLOuUVPO3ezPzEiecqKkCaxFysS68kRNmM+Fk
LbJbmQjc3M4Ih+BWPJ+NKswTCLSjsB4UBzWRnu3FIc62O11Fo99TL1NuwkAhlEhh
VqiM6zKRwExeYU9mw3ewnU4NKCxhHi6ZD+H6LTq3z7/5evjN0Gfz9p1xjBTuC4h9
OdWTcsHA3PR8r7Uk/rtGXkoQJu6ZfJDx6PvMydq7rSZr5+izhcOWibA6gQt7u1V/
fEczeK19OnPNRwN4V3i0DuG1k4qMlTJ9KD6j3+O8KEA5ULYjWljiW5vPo8vQUI1X
EnNFiM+Cd+z8F84mHtRDtXfFDsb3LM8Ip6VZN3YPJscVMAmIat5Vr+50Oq0Ljrjd
pRoaHqUEKlFWDHHeqOBNFgFQAjQHOxHB8rPMXoLzl/BSRAQyylzHyerB7FbAz9pZ
rPkoZQpNSawpCaV+P+shXrB1YBe7IkXctYZUNfibCJMQjs14lGdkB7fzmpvSqJVH
IZ+pvl7FXouaUwWeYZecj6I8BFER7QH6dHeJCoV2zHYnLMfYFXkzDup0wcRQ+LcS
g79vVQLLxyNUoI3wJBD3DmEJtvhJhSoJzoyZdySAgB5HQenlLQfajEGgAa8CKgdE
SOkpIGcGA1LSCFcNCKXguS4dAOjAeJouIH8vhpP8oe7v54slZQNnAEceIWD1jAsa
jdWfFt/XEqJk9oKFDXqb/bSvrE6HWZ9AE/gHvKb+ZOQRn3d10dE0xfwQ5FbViCbJ
jEFuKG2KUbSb0Q+o0E6cRfsHSwgprnxuz6j78RFQ8sa26AiPmAmWkaTuh+idCY2G
bf6KBVh4Lbk65JJoUvCBpgRCpV7KIuod2BJbtGrYzG2DRk6aqQ4Y+eXJsVbjTcmg
dvNiCmf4ggSjfv/pdx2lH+wZU5SgEuz0crcUba8WiGLt+hLZJ/xfPaYNXKdGOjy3
saJdGvNLwFFQsWf8nXMXKZFqJnOUYFaAm4hAn715O3Hdl+hG/r0f+0cfouQFMhg3
yyAZDtvpVrw6GPPZPz8xd/1BPtu7+iz43SziRh3Jn22L3v6deA0OO48tAyg06ehS
42J0sQ0PoyfMXtpDLTgRFYVliYXqbj8vUnFfbVjkCJMb/tGaHSjbYFSbVBQgYvGQ
wQ3VVLHQvceB+TpPOgQ614ya0vku9m1nWLEzPIV44Gnwj29Nqr+5P044s4aOiCLm
EsMIT2zPzPh0RNENkC86dJW3yRU88mWD0tKMjn3eVCsj/vrFcd9Q9CEnYhaBZ6Xu
pWzyniVBD/1mNHHq+VxotULWj89jt8ra/3Txa1hYpKfVEzLEsH5xwylf4QK7fHd0
Kcby87SU1ONbo5phdVbv++lIF86xweOQ5mMat33mLmkcaz1yzfHJk3IZa2B51+F5
lUEnMwRQFA3jfkb+sgROqPPCGtKkYYER/2jxJVz5Gwa9z1H1/jSgqT+rGLd9N4iB
L3VQJip0ab/ClgtEmPMF8mWodSa5nTpJEMb2TE8F85v3FjVW/SGY6GMSxelS8U4S
6r/Inq8joBcEAbBOFajvF7gAkkcrGkAHFh+8I/B8rCWUcIUj91BDhnCNsCAI6rRD
53VZm9rqbw0UxRlkahKZm8H2D878JxnWPZSXdJiDegvWcLSDDQLkzzYmT2uKO0XN
Idga+OvDPkBIMf4Ohwykf8Qc1XlamzQHEM1DqKMDBSdWBrZ7nrSMxM1vLnrHUko6
bVWi8m1+dj2bEW9Ar/RPvv63LUTaMXgzhZ3Lpl+wjmjLjwkItmU89L/8ia021Pnp
PXyO2mcIlcqptTgJpAShjyKvVpRRLRFvP9rvpugmudSHxahZyY3PUJ//SVnKGVYA
QIP/WIX8VAvNeApPC3469ljJVUvrmjidnr2/Cph5IuA0kQWQkm1yhETXrwzSKwra
/ebcnGQttCjU6F4mmQFz4p6jTYSdA+rJ1Gl66gDQTBvKf2mEBGjQ37rDPS9Qrh2G
Ci33LGp5BrJZlEWRueCZcSKtN7RLp0G0owavZrTQBelTjq1U3ncAe0dD/EUzfHbD
NX3yMUtWnBDyXnW0/vE0CqgJiwWRe8bRk7LwyrcEhPeIue5Hd3BgGApgaZ37W7Dq
LQtk4ZJnVpZ4CII8w0UL76Wax1nO3DlPy5j9MU3BILu/jRLUXhg7aceIyRoue+SV
izl4d1BZjZPQkhUmTYpXQbNFAtPsOA1PYISpyHnq49vAYL7MktfvTZ7wwWVAHqC7
QBaUHSaa7vxGivF/viZf5WjoZAXWfg/W7mO2y+2gNTr+NGc1+KW4I0YV+z1aKPG0
TCX4PYBknrhujXGLnVcFazLjJFxmchOt+/Qg9rIFq2jbus1L5fwqVSwaLZES6eQE
9wKhsa8WKrxIbQxkYWuDoh+v5W31S6l2tzvX0GUC5p/Z4Y9bio7/YK2/AToIOnQi
NpeT322yZeQptoddNwPjUAJ+EFapBhvDZNH0GHFEHR4Gyhd2X5xdhhovu10+C5yI
Zwj2uHMNankBi5NlGvigvhrJoqkZlbc+pwPbZIJSQdoJTJu1LBp0LNnpL4dyW7aZ
8v+mhfnahRCN27yYsntCQ8+Li8SSzQ2uDGmKA9Wgbdv3tO5aayOxqjx7yrAac5H6
pfwxCFOFP+lhdky/4XF791HzkNaeyBWVBQqJsuTFoLhmhsKRd3c3DjDF9TYH5AWJ
rYDoG55TO4qieRXLurJ6Kz8zN6k282gT5nutPA7btl36BlFHmQi94YhUjwb0vUQg
Fzyg1LyZEv1OtdMLKBXE5VuD/xReytUmKbhr+PGYBlBZR1JErrt8Kth6DL6ytgEu
wex324+lBkUnLaiByIvKWMXlJmT62NJaJEXy/yLLwuemxrEPqRlNFTR7++VvEHJH
DFoZ0gnoDZaHM3/Zye8/LrAgx08FAy8eMonUHS1L2XqvY4nUHCYH9WC4sQX2iAhm
0jVozoI35lr7RhNYXXF4qfpqTJ2aPvmYIOCacE9ljpgGTPMdoa2X40HftWBtCmM7
U2LUuizzjPog6nY4h0CfbFRhqdMhs1i/IEJ2Oi/60vc7IPpY5SJRFyiXpHanTH4q
G4I1DiS6s87647C5s16sx+bYXN9Y6ME18SZlhkbHgt4nWXuyw5NisLjMDlF20mkU
VqKKrPDVpA4OmfvigmEyZ4H6n1otQSQt0fayrzh+43biO0D70thYKRPrTRcF7vr1
h5IDmYtxFS3kO83NAlqVhhPCPSS5D8wiQVpKWZkLJwFwy4IqNnjzdDBzCk05xzP4
4thTNolaFiaWNNXRp1dFPC759qr+8B48CRvgIrsXDkO+9CWr4kEPLKMFoovnFWEH
VWhWftR7udqTzQXvdx1fb23VpB43dkHxEbbQCHe4uL9lgL24eqoLAacvM0+69p+Y
g/4jcoGtqZDI74NQww43iOKFrvFBpRydAuEqMIcfWZlEvVlhNkbSLDVx2Y9hgDuW
P5f1oro3NsRVi/8ndQ57a6Me+/GUFWUIKtRRg6hwPJyBbw8fxjqURVyYE4udpDE8
QitevOGRA/onRyXH5jmOJjLttHSV0qKHaDbEM0f5DJPpsJ1/IvWdOkxt6lfD4etS
Z56bHOS5qu+0B9+aYzvr4AT8u65JFqCpj4JRZ8lwZ9uVqB5izaSkAjaOAw9aEaNP
sdlmQfovd/G66gTo+UhkEsyqPwjzTk/fZfkr24lVCzfaw5dZ2kkzTlFW6chds3Hn
i7DKj1XeEUlKQP1FJxLIMkML5g0KDaRk8Wrk10IFbIP+n9C/2gbV8h7Yn9RynriZ
kkEU5JLo1tCEPiTUo8MHsY3wXHwHPUdfj2lw+/IxNFluvuFcCRP/0RNMWwMv38EF
PAqIEYfvXb8WN7tgruVKUgLzxgIDGUWbIPfeTR6Gl4RTm1A4mO01u88dNfBKfVaj
KX73X88KQXRw7hjza3DQHnRs1unfKJ/2qKAPHskWB3uTZoegY6Grz0Fx1H51KkFM
zNCIYv3F0KVjlrGLdtqKJ/8Zac4yAnp6Hn5YdS9lKMs4/KNjvSw8M+WSYK9g3i/A
PAfXCV5Lf3Z+tT7THuzyHxV61ou6W0C1yvhuhQk/Fl6xkxhtWdANGN5QbHKhh7dT
g9QrAD3dYJ3brPNL+/oI3IoZspdw6Nga2kO6PxPjEqxuOONq3dE8mnypBMHToaHc
3XnFPjw7wZjZXXd77Px2bQ3nI+UnuEB/6Lj0iKgnVjhkye537CY3FlMhr4w5D1vD
3rsF8gMVUXKk/ZRG+E+yULdwcUYmT7wkBzgdu8OzdqB8SMrArcuxX8kpnlXduWDO
ZV+PznFPXH2tGmeiqD+q4V5c2DmuqSb0Gc/8nQMmZUhAUbBbhBhkYfprgr+Umfjd
n5JPiEW4XJcF2R82S9iAKFpvYq2e8hw4A0UZqZrwzFacGQrA5VnvVXWr1vBX9pUr
Z9FJM/gyWRWbsi8E0S/FIE8BLt6Nvoz4HhXoN8SCzzKudbMoHzKm4lLy1T00ehUk
KPhYenMsACldW0Oae4xd4E7+AdB5/S3ddxh6wS/HFRq7afe5Aob6FT5/cRHWwe/d
n2an0lqFA7TyX92/FafZU1LTIKRSSal4Pser46+3Fj9KKCeWNFhtcdpnIlJ77Ucz
HF2dY7fUZ6jh14bkwah0VX75PDdiIe+QPs2L/rG+1dvjKG9IwElGf5BjkxVpquwu
QnABkmTX61KICm2XrRY3Y9b4B0V2YnrMGcqK8o72AJzNB95JApbzK+DsrbRO5ixi
9ZKolFJsMYVeOvv4FHyh8+aKVz8LHEiEI2AplIbnzq74J7E0cdl2335mDRBVsMKR
TTKD6xVU5M1OB/AL4ItcZn8o9d2aZ/r7i7I6qTW5lIQhZmNyKNir+6f0tcFF9KEK
6fX2DZdGrTTmjs4qsVCxngFYPgv/tz9QWbaDrQY5CjsR4s4/IKdTIeHyRffGcPUk
LT1Ixuwt7vIaOFhs6jS1JIadpwjPanTYCP/fj5mGHsUC579haDhN9xuwrs/NvTK/
Wt4iapQ7Z/CjFJHIDwEb6+vzYrFRC8PTTiObW59tGCu7nDzdBXoYIu++Y3XnnzoZ
Zns5RYGG7G2u7fgxbmo+AMHty8ZFVAfMXloLsyScgIokvka/LR9ydM0GG2xlhLU1
d58foy3g7x9o7nTSbiFGSZgMUvFRp04nO7cTL8jWS5EvGusL5KpB2PJ83t8e1b+B
BLuL4HXVbNZXLaQ15RYoD2CSYeUzalilU3iGS+EC14UWwJjS5pFfHcmy/s3BwJjE
zGRBHvgyKB14kxilPFQhROMUIIDuoAeZTLirSwCKObCLm8D+xM30n+WH5nD7rXkM
5DatNGTdprJVFi+NHYuu7UE5k7ybj2VIckf4FP/KXcZ327X/h0GkSqSazhOML4EM
/XtSY6bA3/QqhNQn/mwgLUnjmC0Vyqsp1NZA6/xc9+B0LVFsN8qF+F2Vt3nNaouZ
cxVjSG9caprvcTnn4iOKQXuaPFJ2ZQI6wSiEnzTiMyz4jbMFVdvxdUbrEUSsjiPe
u/BcUJ/Erud8hcNyfWyJGbgiFEm7k51xrLmFvZ2Lr4kEGOJ4A3zQ1qaHxN9PBabs
SRAZSLBkG2CwOBDXo4U/sB1AiUppFTwUbM0N0u7rAevETQqHvaexut9iE8Jt8zk5
8pGFkfOC3HgVRrYPp5Man9oHRMphtIftqQdTyxtvOKqVNvVO9x7stuQE+K5Z8D68
m1OxQxC+QdIlCX577q8yk5kVlnaZpTXZGBZ5XNQB2eIYkfx7+h5z498Au1B+/u32
pjlZQwd+GGcOB2f2cZ6STs5+4M1kyXvLPbWal9OokllKYSCLL3px32VawCkpuxWX
gwLzYOpWpv2qRHFr1a2CWf/6dA1HDueIt2xXipZ2djKt87t+VUgRHcf2w9kKQLmO
op1/IFz/N7gM0e+zMa2iQlC84Noi8bOY8tZTBD+qJpWgIhLSRE726aeoBaXt9Az7
mMZq7W1sDbjzK2vKBYu1L83zLa+EO3N0N1sK7T5yrf4vw/NEvi8mF+77FdjFVyIm
1TdTHIfFXiotXSOJVziAlAdcYWDbquZ0K0bjB/3p6g40GnJwh+064sAz2S0ZCGzT
o9YKJf+reRm61lYpvUZU+5VaenIK38Ejg9umJjhTvYEU35sUUvPCgYVsikI+/kNJ
9zqXJNGcxExKrnvEfFssWCLsAAfCkuI+39cJKeL6frmMuB7RjzK6hbAlmyLVGsDR
Nk5AR+F/gB5VPFoeLRJe4U6E/0nJvYCBoje8RDRhHsDRWG0sxQdjF1hjskHmPFpM
xZaDN/+6KdSMZdGE4wk/9653xdkTI4ZZbRM2J0F7dfsBuDcMld4q26t9bHieAnU2
E6u85yFVKNUijKVC3gTp3emCo7RuNh93UH7M/xEDT1R7jXRcyxgqpFIPJFydFnTD
h11o5x2+ojaQivG8GwWDWOD8PVaEt9x0pmeanyQY3DsOujJAUnCs7fQpJo3f/cz+
8L8WC49xHteUbIuExgRSGhcHKkgL4ZDekO53sBLop3PC9DfLyLGEIs3iGXOMmzh6
3T0461HezE3YB9LWWCCI5VbC3GFLI5qk4/g2V2BoEopYdbPJJ33sdMAWXdYjoR+T
E6iA2dKGCHg6SWsBsug95WiIyk8E7X/5uIP9Pfeiho3t3XuJLDHE8KGliILSXxu9
FBEJRna1r3w/HfoWYIa5HfGvuxKM00JZD10YhFUtc9HvCFtBoJM2SsPFJb5fpyjB
ZO/cRE8TMMd618/5led5j2iMn2pPJnyYY90bgG+xot4VkWnlOqWgljKJ8VC6ULCM
EPxlLjRxAnpeBZBwmQt/I1onf8cAz6pioBow0Pcigy03AaM8RzRQOJhN9oIsdal7
3HcAIFcO8r4pd6uA2q/+/FAvqdEKfWFyntfJAQJXLzw8DDF3t68ERlDdZzmPrigE
fEFT4UaDvv3tVuJ+UkGQhDxuSTA4Bx6lDjbwm/ksuN+1j/aV12sIlUIYVoJfk1b8
4L2XWVT4IEe1T4pcCgs32JV4ru1lYtS/DuYu68nxe8LG8QT2ag0QEjBslIoPHljR
lAl7eaEpeXeScrjVswBNB8/hYHNsNevhAKMm3wEI2TfwHUJwV59VjVljjqoOFYiF
72xeKZMp89QuydFBzIHCcCXcKj/Gy9Ba6SbHC2BLaKOzICYWQGEDVfYR3ew7oyBy
RYS3KAOGG/qODFvc655A31f5N7aRz06Wt3DEaps75vkE62qbFZwhPr7/yIRDsTgj
KlSoo8PJLlrUJx3ILbcKkBdr76Nmher+r5MUeyNv5TReaw/HBLD3Ww2tgJLu1UA6
csV8NMXeFKDTG1BaY4iU9Os+nFLxFdsYIrqmavyB8EUVEkd+2Y4abdQOxWQvDSJx
qt3Jg27wZtWqokqFg5rlx09v+ELurTmC6KC3WwPX4MwblU4kKc8KEuZvuHLp4xGf
bSmfd62nhJV++/fU6f+fFoFXBWnGJJlv9t6BnwzrH/74tAw0gjQWZZyZ1d+d28nA
aVt15Jeu9B79ws0oOz3Ae485khA7SRzZZgF7d1fyfGmIpiai/Wq984s4dma812hQ
m56gBSTrB4d8JehzMl2oMjxOWERd4Hm4Nk0Rx2qXPTBmECwLiMQPae7wN6Rs7v9j
tgnPlsTz00FpyKG78TgTuFyFsJ02OeInN2gKBZR/m7M923aSuLStpGVBWxx/Bjn7
xgZvVQHGM3qy2XJSj5/ZwkcNwicVV26WCnrwksl5aTaPK/j/QDWbVXEFnCD5T9R+
lZYENFIaLktVT6+n8M58AGXYZuPttQXCE70GvbBYnKEOpd0YdFRS8aKRBZAeMrZ1
QlEcnh4OfML1SJ39OILrHPQn0pDqU5QxY87MtYVf0pqOv6hAKyXQmzjrJw4pljyW
JqMkm191V+YzKC4kwbVtzcfbd4KUq0774RJqaDEoPvi/tG6l1bOvglERe7TAZOd6
evwX0WROA/gIrqEn54xys3NI1S+tkEuE62FBuXXAwulIQhPLGMFASbmmVXvsMekm
UjI3Vr9qMTIUGAlLSjDZgdTPhBFnYeqFQRSeDB6+Z6uyJF2uOLpnYrlWn8CPMIFI
rXOFDXg6KBBTrCuKvhW9AoR1ypLju3vN7al1MBi0xBRVY4XWPfGR99HxaY+JXkOx
eTGEOJIHzF9mn1fNzQGAfsVch1f5KpuzEmELGsSxn/LBy/URXmCk6UVMcsOjJVls
wzMoietn/Upy+/4Tl6HigmI4tOFJNn0UDQCJUg/SW+5GR3K+8DxL0J+ujiMiJjk/
xu9X1+WWpAigdKVvsKYoa57u/qKL0v3wKgW5/piAnziBFSD+39afpBWiRfwm7WA0
QRGgSKL8CUkEC8TwIwbAIbDEo/BOWtKbeMiAQLAcI50hVCS2wfRyGRtevSNdYmEU
Yo7cTXTrVgUJjZ9zbUUBAXQDUGKOz5DTzswnBINS9k7PEa0wS+kbolePtO9klumg
K6WaCB0f2Oyn/+GUTeaOFT6s1k71mEVDAcjLpnRmap6OuYKCYYRmGW+s2H394fmz
Xktmjy56SnTNAMklf1vgM3cM8ByodSUmt9CiuGNJIhaN579bXQKyzZ7XeupTV8Bn
8RpxH/C/mL884sogDuNGEPqc3HGVVbB+lKziBaVff9ciP2kv1lck7oW63C+/tqCP
RmAbo0kCKcFvxxWeyEa9USrt0bKdQjFUwCqtMif7oZ/2rywRwRuPCz+AbIKFPaol
fTm9P4IwAIMgLK0jsI2iu+YOmG+lQ4aSpVSpkIq0laclT2//Zdmd8qv7HMZODl6V
HUNBih804YFQuoZxJh03qA6WD2NLHo4T5nr5WRUj7V6nknMfe2a8/2Gt3dTWmZKT
rg06aPtsq/hEri4+FGjSIFzC/22+ZUejnkjt/qfadclAQPXML+mftH+GyTAvsyUw
hzJaECq4uqrShcD5Xbojf1XNKduXNkioAEmVuAVCElZ0gq4wbNzJeG9bL24VlZb4
xLc0vW4ol/wijdPVEh+Mhk52Nea7yFZne6hInEiiY5fMe5cEVTn02BUIoNOTx54V
m15F88/CcUSIviceFZSi5KiCEWjjo3FAEI/fGUFvurIhSEwStpoNgdogUx1wukC6
tW/nlN1ysIBn6U/bIG2I/3VidlRfeS05fcZkL9k6lQrsyCX22pZx3K/80t+r08Bi
tnpTzNn1Gr7GccrNYhjskD/ALb1aPOLEQ6YbehkDq7B7eWg3zy2zA40dJua/1mLM
2gjcEm3bnuGx6YeqraRuyA24ZhpJT4sxNbL+dxKJLBaOJQ/4H/Em2Rl/JBNEpg8R
2/g4LLMSIDcX78+mJjADF3HXsl53pNZAcByV3FJKg0wksbftg5LxTc2e5B6w7kOT
MmoH1m/mlhYQfk6YrPlMkDX/h7vJG+KxsVJCRF6uNHtfE33je8cF4fANUIPGj84e
vVPsSrKFpQqQFtbugt9Mmvf6t+2hsaBWOPVeyHaMEg0sFl49ekbGEu+X2cSP2xnB
32W/hSFy2AnBVtefpyzn4HbYk1DF8N1xVax0wFyDN2atyAF4vafh3ytn5r0oSHR8
SBOdD6pvF/OVxZqG3EkWhc0+2X2oP0e7LOD95M0qSJ1Rc+AxSfV0AGwaryHk7mz3
ibMxnHO1fXReUXH3nub+Uh4xj4c42i5o+Olk3zVX03rGrKdA/e9InEwj/rdv0sTD
1wRPGDI93MZoJRbZPyAQQmUVmm0mBTYfifeizD0bMNvnh+vCa/zS82Jh/vIkBoM5
OGw/mPmIObbiYRbdUmA8ZHLvwJmF8vR/BiAktdUVe4v3Zv4RA+PcCucLJvukxbNB
xBjoMqembxa89jA3CDbvH0NS31tJQEm+gWs3xT70QjcHJAQUE9zWG2nJaMzkN1Wl
NtxjqOGa7YmSHaC3k8DB8BK4E3is8yeEuQMjIdaJsDhr9FdBPD2+n2FmoPwS+gbx
RfEOcsrUC9dzSlnvxoKx8WS15slcb5So9Zn7oQ0ov2nyWMG+hZXbK/09zY9dQa8A
Z8KOm90qWluHqmD4SV2sQ5J+cDp0KkycLqFAgtns1evTVsSs7N/UMDj/1nb7ZSXD
FXhDgts9EyUJlEFh7J1HrOrA9E9WEkRE9Gt+zmolHBp8Rp/31x0BnF/A46HfZeQz
IcHtgFX0iSLnsWo5JfGmTR943lbd6OH+ixRdX0n2IfNhHips32Ti+MlI8Y2jxNOt
qTwkA1NxsXbykbZz64iIcDFvzKFDDS4NHM/UrBN0fLcoPTapgQToPS0BjAvLlrJ+
8U0yrJLRIYmeZ/F34kIHrfGXZds6ttwp+bp9Xn40FNZg4iwvQrj1ZSk01oQ1eZaP
gSe3N5AoU6FENv/I87iDwRX10POPlp5Lw+E0lypzxvmRvSWGJ4kUvJkaFrhx9A4O
YzrpkVZ0M1Wdf+Uoiq5VXxcmFe9lacSHlDU2Mp6oriIDojW5lLadms1LjWSz6iBe
XZsn4c1rKMWI0jf42RF1il0TBG0RxCVeR3bx7Q369TC8qT0tRxkxzmNlgTsn6T1j
e1q+Jwo7jspQY7kbvxZlrwXZVyziPUbH+D1LUr+ude5qkm6/p5EhrxO9U9CW9DuA
zxiCqeecr1DJCwu5WVAUWOwc5IOs73gJwK1NQa9b6y7KmFZB2PgPlExkafJxNmZ/
+C9tZ8cGh6CY904z2IATl4cEmkqvNUokKhBG6jL/w+UxsJlqLMxUt85vwwWVh1+N
ZM/x7RGQgW7n2MPWEU2juKWJsennTDreI001V4DoDyvY60GJmlvJmLG951Cw52fU
IhKl2Xjk86rs5tAGBjhLhVLt/tVXKqDxNN+Ok8ww3FoKRLEOzu7ZAGad9x4aaAzk
aMDEDPEf9efHJs1AtBMeYigDy2gVpD1tUSjR7+Lo48uUWGp0Xotj4tETWdqRwpX2
l4uBuqqXQpcGZEJkSV5L9yANTLYe9aO9L2jTKoI0gACQispMsaIWXjpKkEy2mVis
i/MVrXv2L1rusB/4SeGQAM0Nu58gT7JozAodWoOEPqyCYEMEXVXf1t1wEihehNd6
+avvQ5NoNJGWGZdzAB8Rru1v8zzI/nOFeDwYGbQRJGFHARZYYF6/RQtZioQEkl1w
TQwEFImeTW9wndTH1B/fOB6+hEHIiGfJn371xWvs9inBsOZ8OH2Pdeg9I2RfXROz
uZObPU12A4Kq2WVfXxG6/A4ZcVYr5DZ6QW7wSuLUT4ig+fm3eZJKstHhXIe0XeDc
8dxhuvMN7IfLW+cdCdIbu6ISi8rXd/XNjE0AYIbkVlXtt+WJL5vX2Y8P2ceSVAqr
NmvuTd+YImuOEslq4/Y8Rat4Ei1sOnekbi9qWykja/L3YcsD86f/HGLzO187H8Rz
h1L3scdiGau5Qo9mylefcV80IZfF0KwHyyTK7d78U8JOzdN3Kg4fM/PQSUynXSDV
agpTA+ThkhPLzS8FjeoxZNx35mgi26miKGzxINnkJX0rL0KdB+Df2ySZIFEOFvjq
ON0pOzyv527kcH7XYPb92bsotllaITdoTq7q9/tr1fsd41h1POfsCkUyRSpeuo5r
eurJsRIQetDDlvk2Ovybd9a2pIAK0NGkDz6QR9CNmFLzKKdq+lyu/Eh5EWT8CIqj
BsPKD6fmZ3yf0sS/b/CDi7KCEPjHsWvyt6XipcP9JaXemjJoLA+Eo6KDBRTCvRwS
K6uA8CO05p2oO2z0fCqtT7+zRvE1if+Pdi8HvyxO/+hw5Tgvqc334TdtBxZVCeZC
7ZHYlMxBdWZHB+FsYV4Ytf64a/Ql4mtmRiTbpeFlYamPDwmspy3gG+g9Cat9lj0+
am5WHFhbLHEsBR6DHtamnUYEc+LJMpO0zSBnyOsYLlICUG6c0Gg66hBTQhsVXYOs
qZupSqo9iQhSsG2n/giKDpStVG54D8WAg9WGwRtb9b8BDcg8bmjf3Y6HStHOskPl
35kmIRUkttpmv8sDsqE0lvJnINOkwnvlFWUKf8qhDefodIae2WqttTlpGNowXElE
fe4/9DX/0N1yY7M3Jd+EQ/WGPXvAtGANQTB5q5Jq2DqKLhOUkiv9CcbP3+weSOCm
P4vhC2r2/jLdZ6znEV974mg1aJSWv+81NKlkP58/+bot3IgV9vRO1ekJx/mXJr8V
RUEQq+rJ4jPNu7GcBgpWtwAg7tpLeTCYYrS+8o2neMDlBOcFuo4kNSwVafR87Wek
eFNMeEGr3Tc5b5WuEgBMWQy/HLs2Ox/wImbOdZrOs40hPeOalQ5UUodGzfOWb/x2
yPwD/K3c6Va0s7QKjz43dLliG6AEvaUfOCD4bmqQ8rxz1URYJAzRHPCwYKAXiJux
u7OX5+YKe+MTXzdH+AFwbhi/ArwcIFS7sQMs5+VnBf0VMSXsbiKi9/YGazS6gcwo
v3q0atiDfLARFErzvVgkLtmAl9rn22DC4RoIi/Arl1kEtN9YXBagUSlH6yKrLXJ+
WFn2k0ppMVFwyGhKDMdmX523rFH1qhEY+0n27Hr/0ctkHP8u/0f1DmCfDz1Lt2Da
5f7CjSx9fb/TB7TqlS7YBSmzgYjJzaRapi75LEroAYw/20TqQ8LeGLnXsGr7611L
fc4RKi/I8+hPoOP9XIp8vlr6vSKJDT4V2H2CnPR/hX/agMUrQ3xu66Tcgwt64UXo
XbXcW3GfUcLctSI9LzHwi4LHIzANyWq9SCcnbNPIe6bAsy39AJNYdL4PygMmQ674
pBFLvliVjUEVPXXAeqyR5KQ/Ft8Oqz5akdSj+rouJXwztR1l9XP+h613UtxATA4P
/ZEOVPw6cDndjM5IfAKjkr5XoKSW5VHwjtVUqEQh99ZmNp64boaGlJ3+bB+ANk2t
5HE7tx+myI/t9BpnvJT4GQpfYkQLRlrCaOTQLCui9FfSTj1/DvpngRpQimtrThyC
v2Fd6IN6txlFrrTPCoiYU0lnhkJfRLG08zgQFIWF2FAf1pVLGAMTKIvUTjGC4YrH
KfzSuR86xbVNXsEOdEZKiatze86wIF1GHS928vIrVT+/9noe/cMTuH0IMDHr9MSk
p61iDdKbZ5pcSfjcdsMtBuMvi5L98pyPgkBacMnhUCYuZg+hyeqViFOD99FruoJ/
iOpQu758khwsOkgiJFXXl4nNFReEEmgehAcE2RFPSOTQTYXkTqu3pnSieRzfLbOq
pIkcIBnxI4M4xXjeSVPMYYB+Dl3wpTdddbDteZifEGFN9/76LusAwUloIKZUob32
0WBrF4at0V0TRPWaX+LAeWn8GH/AorFwJOiK3y6XEM6Ebin6E+fY7zVZDs8VFfyK
V5HjBiUhirzcHSkODDkKmCRgyO3yO+5mgn0QMlkF2Sk9W8hT8ib2Iqqt4HZjtvfs
HsQu5V5O/LixcNLb58pp0prPBF06a7u1KQRm0NUS9Z+1ICdGq0+T7FFzUjgF9P0Z
+twUYRFIhfGTd/iMusrnYJxkMgzqHUZ9ye0XihYFT826ktiUOL7kj/DySYb7oFEf
8GJhgVpue8wfl8bTKqssUYHOGeQor6+tLcpkYGBPYH9xgIUyzKnpNv5XE43BPW2L
i21sb3GNANzcYusFJfmKxc9ylfnpjJWVkps2gfjCRt620NMVyku5YAP53c/+otEV
ysQ/ceiYzO/q2tEjaAhXiZ7QSgZQ5Eo7E09xmrp9a9danUx6iC7SXUnCCtnbXjYV
g1EQF1DLReTRcK65Scm8/BYT3I/oInRv9ix+Md5nxTp/ODQugSLrFpUjdmeiHSFB
7BCb5Fha959oFFfSe43CJqqtZqh5++A41h0YQlKUAnrEQbNfP3R8u/DpgaGzfPI0
vMcBinvgiDGaLj497aa0uqGjf3GavSzfLJGlmpzfkOAWJ5EdjilmK0rWJu5iQsR1
YZ8vxh1vZL09r931jZU7F19cDs+dzjKTqgLbwn6cqWn+VyJkf0ey/9nS9cmEBF0F
f5E+re0RYy4fThCgYUILRN8r5ofHkJy4Oh9heR9GaQQRiGRGaTVPZtcXGV6j18J7
BnBi1DnnxCAUwUzYcz5LZNXEzrDkSijN1ZaRGubO8eMUHJR76rvAxFv4ggqgx0Cf
4N90ZZHNRgtiVFeng8A3zxZF/lFN6vBSfsfOXVGgbOCbplXZ+n7o7bvYwE2iWZDX
AG41whG/oOTbbZG8RGWMv3IIQ8JpIPX0JMVnZPZx5IBsSKnu1ljFmQM2LutfzW7C
TXF815BhrwB8obaNdesnvsJtYl9MXzn+Rh1Be76/rOBI1MBnRw7UA1K6I95pYAOs
4whQuANVso01xIjI2bBzGUDTmGLra/yIlPBicgWcJgcDsQIzS/dx5xyUTSnn4I9k
uwfwNtbXvlhEpQs82kjw6ouZwQFlSVYr8FWrUr/RJlzQLBArQ7sLY3VCInkY/+x0
pcdz8S9VAQEyMScfHdYyR3e13IaB4qXJByHCjmx7eiHxj0lf1M4j1qczZcB/Pe6r
stVqPkCLatgqbaMZ+urD2clkJWVwwTvKWBBokgVEFpekkcyQQrqL06MDjpc9pGhb
LJ4qWv72q/+NH+TODHLp8bCBHcRIaKMV1OnRlvdyB+q+dfkG9P4Bj7VECSI1qjph
Xtsi//QoMoZu1Ry8jx3MKsbxW6CRZ2NSucYpYhQ/h2WFttxccZMxLoeLupESztHi
9kzpq8hGlV7t9x+09Q9MRqd/1l4MUGRPaaZ/eK2fQuXi57yMyVnpNImxMsRwc8Hg
yF6AOoWbgFQJttWpZS0BAeTUGRg1wf4+d/SEIgfpxAhlqxcZJJLlp7wwEN7xfpFo
UQ9H8CVbxiQgcrBexR2TKpojhLB+CkTixOuLHHcw1AkRxW55/s28ZW4/f4e8NCqh
PB2R6WQFt2cbQs8phDWqgSymbmVQMi6wP/Daxwaqvh/ljC134f9LkJfKM9ZyLde3
UJ9j5aSHP2BBQUslAfGvYRPfX6gWj/3bCURM0fI/w/kUySEmskm6g71nhrudXE0S
UzDKDmXiW9ec+IXjzy0VWejydH0kofJ7ueOfdk6ai+JwQZ0Stp9i1mKrtqMiT6qw
UJ3uoPNubQ8E8a9FXzM1qHlcq/ws7mGBVKPOSApYL4Ovk1dBepx5kU2NR5ZvuURk
dh1O1NB1CeKcL87tfK5foy5DvkZuOx9GRxlm/2D6BTrhx0ocbmojKXWHFKa0Ho64
+E2M7FEB9jmqHVt8TcxkouxnJEFRx1dX4/pYOqC6bKTtXXOnH9Z4XfU5JtuJ+ytG
c3gBjXAtN5yesDyXCt0hH0J37tWhiD3+qL4n/YcNXKeVx7pTJpdkz7/ej0lq7SAW
dH/VXvCcv27pKHTBp8Sh1KUaMYKdFghsehKfNNDv2fyKvRdFfreXLzpdQlWIq3Ou
I2Qvrs6v9kMnq3Mbw8QVDMG2805vwW2EnpaKPBUsBgPprOTiEpdQNDVgeGNwrbOi
vnCPMHYrQMgnNhFxK68JHWJImgC+tBZ8/hkcK24GGa1GNIOHI0REn3txcAtfPOYB
3utqN61g69k1irPKj55qdC81ugHOOxfkHd5HE5B4g83qx6hsLiAQRbcb9AF4/ccN
lHjMuyWJf9XLnxfoV1fu6S1UErFQlpPS35KO6cqHCt6NTKgq+3hD3toV9N3PEEil
uWQ2lXn455Ficbwv5enTiO1OWudP6bpHnVyVpACM0IQBoiz5AYPyk/Un9m62oBzD
vzXuTC/2T1zLMIx0TFPTX1X9xsZCT988D1J86CR1/kXWIi8syWvy/ZZaXUT8mTv3
cMTlVVfMl10eR0iVBv2oMdb8wFmL4hMA/SqAKfhQl8QuauYNP6Zfb123KraIo9cs
pcbpfF1YC2nToKHxYoTv/fjoKitzSR34PLgWNLhG7wr9p14Ven5rvTwYgCEPeGne
J4Q08kivE4Y0bwCsXlHPLYZTzfWVqc6mx0MXK4Z9OAolGZ1bcD3Qe5ZhMnrrUTV3
elnCLiNfIpwutM2ku0zQ1MXF4ymClB8yaYCc/+3zkZ2QQuqteTuMKvXu5DsI0RVG
XrcyfH750P9S6yw4UEbfwnRpUviPdxQxM0KLHmvHnMr9s42bDKQ5toO8ntyEN4B8
275KpTjOA0dmjPeOwmmCPUAp+E2cI9I29tOXTwMHqiuqdbu029lBj9g4ohu7DUvB
npKHXktLccn2/HvaccmAny72huXKIsFoAPV8e9NYM1byBAuN5Jnp9V3Ln+y3UIwl
9fj1b6kojRs4+KK45ZuW9bNgp27iuDEcXri1VItFgtUYqgP8rpkygGFr6medK8zh
jX7FvYKb4eHIdUpaFJ/kYHst08TM3+lNzNCmi396cHGX45OMXTaoebhz449hzDxs
iNYp0TXZ+cbGJ4O10Pk6X80M25j3SHwJT6IfxRj5yAg8rx0+xJkFH02ev0Mq4pv5
6B0KSZzDxgoJJajuelXJfgyNAUngLVbPgSPLuH1iAF1z6BsHRyJmMs24LBMBYXXc
oTtoVU+KbLBD76TBwzyRAXJ7FeBT46NRiKk28gW1ELxdDmca09/kDqHheumbBesA
wEc0GrGBUELMGaVPvRLYZyTyrdUY+1pgC9JC0WpHQkCF7uSaUEoPzk+IZWGUeU8B
IEdeWqHJnfDDHm25d9afxH/TIhTQGZ/lDA4Zlu+v8WbywYTjshYlroV8humf2W9B
TYdEwtjvPqUMGXTDSF43/lQqJ6L/O61e2POVZ+OSrqAbdUYQ8FXMt2PJY1a4Itxm
ZSYvkVvVSt3iPIeqm0ckXRCqEfKSk6yC387cGmNvTRTLvOiX4gNHMODZFQRLEloT
gEeprGVT2zx8kWEUr0eJtuu9e8/ODR6I+fimBxQHIgzsGM2fGaRj5U8Y9On/Hno9
uCuHRvQvg6pf3qJNeZwH56wEpgUqZjZx0pJvW9jCW4ASnSePjysaDOY5MY2aQWw9
Vudcy5NySIO+Q6jn2IGq0qam4VXpwUu3jog0BMwopnjqCDPoILEmxydL9IbfbfY6
eumrYvhNo/6eFOlsyaWC74/zkmdFuU/R5yoWERM+hEDCGpdEa+cSjFioZXG6rh4B
kVfXKbUCQiVCvl3SpybE1t6XmrjsGhWAaKOkinrhVNEUUBqM1YSU3BAFrX88yEd2
LTeKqx2AyIvuBUACJ6nuvg/aRwOWGceuzOZQ1/hNvr9b18hBNkCBSoBW7J+e5mLZ
iOwOSAUvnrqq4nogE/GFXL2moUmeoAt0yoVtMBI3MauHUM2u9bmRWyzyAOBFPTnz
l6+v8hOWd0tssPDmITNZbJmcKHR3IovRhd1+7LsepunaYz7zetIhZMxW8G3/gZuD
EH/Uqd9ILZjloLXfD8fXX9xKzjipkvpl3XV5k5hXPnhpDg22MK3aUM0uTd0mEF7p
TjRXZ6m6t1xrDPYalZ/3cp8bOf6loQnmTXi1TDA+1+75UAAQgN3ZYXzHOiMswXvg
7XPU1H+UyJ6eRP19pGzOPYOicvNhHnnCdged8eX+W6QeAy74xXmJZCxWl+xLTpwx
HxOJiZ57TH598KfBXCEhAvFfFqRrmI9L9rT8hVTrDF8k+MZRDyiQwz3fwTw/OZ27
ohzA8lJ9KkySv5Qbv5cDxogJ91lCQl3DTr/8fc2ZF2Iw/LajDSIXS23CGk3miP0A
MYpRJF2PIkZu9VizhBwfv6nbKHJ1zxi7mPm6EMzLMHfqYy3BTVNTEC8oIMg8/MXA
u0GVrEL86Ut7VtoDXu7KdDejnZpV7V7OeIx7exPJLUFCFfOcaQR/tPxkEuJRvMzF
FmSAqNuDF1ipdIvlmdg1wTqRN+Xsrqkx0csrISpUqzag0XQnrP8PXl+Yj/urldve
YZ7LheX3MuyFgb7FV5ouiNatgwyzsT8bRMmc+8ZuWfCRV3FMGxFbrb1QwSxI4hRH
HTmJ/WN9qNTxfeQ8l+vFf8pFZn2ND+/vFDJVvH2vrCASQ0MY44YOKLwgWL1Omyy1
xzodWfLEoeSaewkKfngbhmK+EID1sGgJ90gKN2qSc9GQcdqTSk3cAL28aGtPErrJ
vr8tr8gI3Shf7TJGXvd+0oTAg9AwUi4kwVNTv+BfdZ3mCloLbbkZjbCWJ1jONJxZ
Ov5JTq2HOkqNuh6aBnSEHtn/YYPd/LZArqnhJh1yzDczauXZUvYmNcBI02YF+RPv
RoH9pUQX/wCfVUuCJ+MFF6umVuoQxUOquvu4Ehbs5GxcswUQ3DKoNZjF6okQ+NO7
+KJJgIcLNtCUioLmVXKKmMVeCPq0v0GpDnfFIerW6LzmSxkrQggW2WHmOgXdGy+Q
7XYiE6sJlG8yZ12Z2N56wmxsYB6Sql+3SFaHeQAgsRvpJrsZncGY1YrMOgQeA0OJ
9qWgeHU3bmBDt74sFONzQRmuCEWm0EHWzrRzkono7rLsqlVzKI9LUOlHZOC1GJex
PTzOYqjNHthhjM6lFrjF0cgjkiMYNeD6elolIDI1XdEqKo9TwVci4imcNlMY8CPr
IuDt2/fBTw8kiTT68aSUoihIQep2HGhFzeSYwm1Uj6uYbUgaSYZY0n5dXSmfdXwl
Uj3EaPWw+Rn5bH0s4hsS8AtEaunjde5X1D0diYMre+UX2t+zljV4dTnBj6R+w5sW
9jHp6GMihE1cdmP+OBFt+uDeIGnFHew1Ejphcs6sSQPRf7P1mNX6AWjt7p11WHxI
lyzd/buTzSPfVHTvE7Ha8wmqyNU3vg0yfzrYS95e8s9oq6X8xYD3lPsEDf5mO5+G
HeE7jYviaE7tXjWXeb/aEIkJUF0QeUzjcDTTwqkapOfFPSLDEyC9WjWfMRj7ovJe
k7cKysH70wrJRpql9o1YA9CBTOtAB4XNGrh+8WNNLKZdYTjDY3ASOSLY/v5WrDuj
g1z9sCk7fem3Ni5vYEIIktCf334xhhlOSxYcz2zhw4djaGTClaxpS5S7rAorep9N
QykjAxeG8UbEfM3zbKSI4Vyjkeid9Lg8v3ZZ9M7F10W8rWjCw1tCzccBe8WYcw+s
/OxFsg0gmKxAVW3zm08HXx4dIEwG9wYsUj/gFU92P9/2nbeiOJCFqExW/YMePTg3
nRF/4AeNqnBHEfFMX7kzpcWXKaWuKWIHsscRJXDAXekgF7LVsjs+8eazAbPC8PCU
IyEDslAQNbkzCOtKE7gZjKhHu6OzdMuWH1MGujh+Rtj4fMqtYFYN08t8UyWsi4dp
zLufcmhKCjWPuO9vJep7qXcWDF2uD0Woia/9wIw/TwFI5ZxbelV6eWnetnqZpw4n
AkWWtPvfhxhxnw4SCeBzz8h44XWFCjMb0sz1oGQUsMLB8/X3pqilBsiykf+fZui4
l+ijS4jtoeawixJV4rZsswJKoDcQtQTEBRo/os2LWftd4VBR/WfODfeyAUAQdaqz
7gg2OKnjCSgbCunRzS5FylCmCQ1+T7U3TjwO8uP41cFj3ZIWVkCEXnUkURlC+OLO
1MvkFFu7Jlea1Zj+29WSYxdQFC/MV5x+SXDfxHATq4U6CAADKGIxrJiodmDinUv8
tciNWVeFXLvaOtJxPgXDQPfIjAD9c3zbkMWNzxCbj65HJ+C0lJGMOk5hEZbjjGYB
8zagd9u++skPMxPn48jmH5cFwnomJ73a0Je+9xjb4np2X0V+y4w+BuY1Fra7nbSo
uWaKx/j+78liz5rpjwTuDLi14jex1oH2ZKQ22ijm1FkkO0PA/z1ynCoveRkPUBeX
Rt6ftLhmcRDTWjE+gsveqWI1m6S0I3cn6kS48TwiI/H0MwGgaI5/JRx/SRqWaUCT
mUlDqKmrV8Nl2w2GwWMn8H2HTfS1VR9JHy+8/WNY2ssSD97aYDpTmgVuaUZTYkc/
FmZKBiWFera+J4/w9KfJskowCS/IFSf28xNsi6WnkXajCbtoOkXxZdRI6zqN79BS
o9P1i7BIEIN6guoyM7cq9+/0tOFQnzl5QfUxZwMun3jhDa496nz44Dehj/RZLzK5
XNhFYH6blxWbxgAzEknW2VKn/qRMxPezRdP/hP4TW/1bk3v+N2wxZ9WKrcGD62wj
XPFsUfqToumd5HoT9O5OnKk9FQwWvEnjuC+iHPLVMrEDGCN8yAC5SY3tzYULfaT9
jNmbhpVcBrSDqw6nxVOMGPh4mHB+eMVkzGSA21bfjPPPfmbqmWE5ieu5oxDDKBoi
W7+VLtP1BsbBMpjicJb7RWGeZuzHJpnlOel/X71qg9lnEodQOmZgpOwxYZ9Jr05a
f8X3cnqlCXRgFFXgWhJuiIRF8jRKl8MLKI6iLy8iR3AL2SnphRhGbyVcF6VFjvcV
SHRtrUGzgJKrS4kQsXZatRVndNOaBsN2ZCjD/0eijhbYzgQpOEP3vT5iOMEBDDSy
1jYNPB3CBTgurZeUUMl9Oil2cyirx8NiHWkInLaBxkLrAvbFIakLgn2Wd7g8KJKU
Dpy653yQPNtf3+rH3+Lhpx1UM3OxMz6YZXPRiIEdHq2jblJw+sMb3oPieM6/BKIM
XsfmYa8tqWSTNKc4iJX639EU5AtSr/BAoDu76OYk2vta8jTRxtvTmnAh9eZFJRFV
wIIsA53VnupVEPS7d5K25KhSf0bDthe7j52GshCJAoNlRmJfONQT5KpbwbP8C12z
V9jOeud78kjynhIn2DPl8ij6UvxMULQa04F/SePAThD78pX46KNXL7+MDR5b+oHm
SLBM/uU1Kdi7dl7ile/QRzmueZD6AhKy+4oCD4GnD8IpGOFM9kcFUuNLY86d9ZZE
zOWhVySJo9wYqnMEeOydKcwJXFT0hFIXQ4uF8B7SLU4ymaavLIcnKtMYS69PGBJd
jAAXKr/ZSmXSertZqnGU/pUzfEQm/ykRmA42rAPdNMdcgTh361R33RuVVgQeMzvD
9sKyZTxZeHnxQJjwTYGyw/A0t2REJa2Pqlz3AeA928ID3eaDBIlrNPIfkfl8oxTx
UuMoH2kzEm/3ebMYP169i/CNQItlkUrZgj3BdsgTCo6X2/7CXE7mmSS06flQmHfP
dd4ee4/OnM6oPC/G61HIAWHFvjm45CIqp8EecCPTawtIONb6u52UrYo+aw9Josr9
rQ1wYgdhnR6mFfGFwWEs56qAmp4gyG5pn5DlXP3cVQhi9RIDoY2Mw5I0t4qqRrlO
D+cTxoPz8/IvRn+VI973PNTlYFR14X0v1pUsArmDeJWhD3eTIGyqMXk10eXBEBxj
gktqY8sXqLhX/hC0QvVXDGXiJ62gTgChQ+7JTSCVHfm006k6jXuujM+r2wKYjbsr
ToFLqqXxIWgS8DayhfERMKV0YiDeCPcSZvewojTLgGIbxu/uO2KDmTqedcsdDbpl
p5gdz2hMRKOx+6z3fjWlPnbhWlWGIqSOlRNLmkFZkE9qKodeP+Wydrpta4gzrUnE
rtb2DIH7xXVs7SDLjmQDHZcXhxFELmokI1vICG8OuBjs4SgJ0fSLeH0ncWgyvfEY
wTfLwBkNrCOoT2w640RcVzybm7XsRl/MTKj1ctDukzzpbSYqBPjOb+CWIltKjwWj
RKYtah4ahsKo6J558224e4OAg42hHinD6MaCZM9R0L8TIDLuSZFEA7g/fN7C2Oq6
Iz+4RqcJxPnY5ELoY5EQ/qNeN7Lv7ogsmw5BTRy1Uxz6HCOPcZpZkyslIe0ahXPw
ll7dalXHxhVDVmdYMaJXPxVZqG2CjFy1vaNWMOUw7L7WhJaxs4klaBkDQyt7MeBj
JaE+3IzFgq+HAJ6l3ScODtqKKnJvG4pB0fYgld8tVdZ/wtgsVX+xRY0/EE+SA7Vg
9FrqHboCxJdKoV1Yb8x7xpu35TSaI67uZiiifcHYCbQFSKVCqczZYSShns1oP/32
26qgOoK0IAbd9uFht/YhVVC3eScaXdq3FHML4E2AZxUvcJutHlyJBdu8bL+dOQkc
svQelNZSvfq7kXaQHcl0xEctxoVv0FADz2Y6oKh1tC6HrQZJYiOjHP8mowG2HgES
IcO8D7x/roZ5Pa4Im+6+uxPcSPmQ7Ukpwh1WN93pH+k7bTEOjqtdoweuZ1mJDhpD
1Ax7k4CyEN6sDgYnVKNjnz0dnSBFS+2V51iNJq/QAlHEXaBhrddvEDbaa7zaHG5T
k2SyvaAYaSVZxxOK3YVC1LjntSSmkH1+D94+HKNE23FXlsMDd162US0ROnX84mF8
Aw3PU9BTrv+gOy43RtBlcvWowGAB7/SvkL+8vFlIkjfV2J9QSKikWRTAfq7QbJIP
WyHSzbwAexHYEYvv3JwxQvixRCdVCk5+waXN2o7Tj3fMO3DN6f85MdwJozAjMXhC
gz1XYuVYR+HEhISadgj6+m4owY9KavfDXlcnJuFLkQsP8yWRdt9A2hPy1MVnTfna
84m1n7k5vQYCblo5BvO3uMM8T2q/KWaFcZpYDCEiz6AL6tZ7vatMCnab/7EUKGvp
UcoEk4r7h4B3Ujp70kqp5O89Fom82rBCh1+v24IV3zewEZUgYgsqyHFgEzoPnsjV
wdzTNCM3Yp4JUIFTOxekGkLR/in7RDud7toVYak7MJPsesDYzhShQa+THLR3t5nD
gFZXTua2D2szjNiBEYqiQ0Hjz52nnF69sHvF9IA8DVTpKNmnfHYFj8AAcalFh2KA
1HFl4ePKNuvRdMeCFYHCrV+KlFsHAUs4aaG8l0SaCMTcWW2M3uG3I7OwCkzqQqz0
xUCwTy4D12WMI2NF8f0L6LVSskjvFJhT9VuIuVVTFS/AN0+1bjRldZjsH7CnUhEe
RH9Duykl9jzh6s2vPznr3LoMAvmIFgTWZKgEmp9dFmlq8RI4gbb9CMoNk1BS2Vov
lozqsz6KKzhJR9LQlYRoUShF5FdBG5LwFbHDM/pLr2bQGJ0TTOaYSW226x3MCdZH
mk6aHnc7Pu3iFVEf5CTJY89sNrUxKKi1Wyz7aitYEp1PRYXgDNotEv83haglEYTP
IbsCxfdKgU+BKUWp4TmZUWMGkmDSrYmS47/CNnpeNsnlb+Vrxk2f1GSQJx5cGzSK
evYnbHwsn1WRpDWF9YOikVxSIwOsxtb8a8n+jps4OXOptNc4YKPnHmd54CnF8dni
4r67taQyvanJo9htMaq2gsFPn6BLR3AvSKZtFtrrtSPhDN+TljyB34MSVVRAOZoz
ryDp0vU1CMg9ayB1GaVSBmXKmYPMrRFVq++ZWWMwmdfaNL3eL5u7lUEknkPLrduJ
DiAPcxOcK08YxcP9zJrIoFl2AWSZhpjv5kXUp7wCTJWloU3gShWFXUvLX4iBqf9a
i3u64Ydkd5XQJgERXu5txNRaS1RAIuGqdx3h6+99aGCOb4AUYRjOb6fXxQgzFrtX
0XheQhPoom71EstZAxfy6YJICiS/UfC3qmWFUukwbfaL8WhcfmsXOY0YgHM/wR4G
9CUWW/juiG2LjCqc0DkI1KrvMClZlaYczqe+VufPoymchc7C6liApwSJi+xJEo2o
SFzVZG8LEo/adtuFgu+Dzr9fqOQlDqjWnmVvCimrEA77P9gm09SlGMXkeVCpBVxM
ujJsKBkjiSWSPZYgggfXurPL0Ru6xialanGeyZL9DgtWxCTNJVmjrO6PoGF6dF31
B8R7SjkrXOZ2dezIVppeuJDLt/uJtKJUlJ4GEaZPF8vPqm8NT2E3JFVlpvpNpk4Z
gl0XzNIz/4UpL2ABvBnsZBmuMq9yLDgHxuGhLg5OxttV+bcnFu1s/M1BbW1HpGKn
xhRFX5MN3rnJ7WcMgdVg39YXgsn7QsIaBD1lnXxv2tToGShD9sQNZbhQzttBlNpr
4Tu8vaeu5ptIX1jdtLW/ne/minzLKYCRWxu3LYwB/U6NQJxYcUUh6SuyGVUEsQB+
ZrTaeqMA23fwaZWI58KqPmotujvjHo8JUjFwLga9AIg8sFlYMoEkjMIEyZZRh4qX
iD2ATRXN8uRfL/EQ8FS9awvvf0T4f5k2DLF2KonVpPoUQCtwiODs4GBnXI67gIPJ
3HJPK6Wv5ONaHzSuUkSXbL3Jwn0dBpO6ou2DUkoWOEQeAn5hE5XlwaGLIdHvMDiR
YHUE/kBj2sSgBSKH/vcQtGj2J9Rwy3KKX+1goTa1w9Mzqtu9mM9zPwNgU4FGRtcL
Kyg/FB8xdqdTJARF3/Fed5QNkbmN3keL3e5w9tUjkdfU5e9k+LY0++zonqRIZlXz
iUPQ7hPQV+IfogKRl3msNN6uD8Yqp/QFMVBmNYfErXsYuL48AjtTKhHaXxxDB5Q2
Wa+nrhyIAAbzyHE+5vxlKT+zMUi+rxfY9Xfkc61xsUmsujBLSn4DRVnoBQFbhp8X
otpzwD2aElDZ3qfGUp+tEkyvCA/igPD6ODPyyUPfayTKBo6UicH5ekAIe0k4jK+V
dLJlLLyelBjQviPqKSkkhK5c3VJ2lSUD1C8aZv4PGyq6HLFxtyd4Jt7i7wq3jNeY
Z0qqLqvShWz1EAn43S3nTGSne+0Fb/8nmhDmtYrRlUvksaD3tGsXigirAJSr/JMY
gprl6KMHqiHaBoSMj003E4/T77WQWb2inxMdI9LbSCA4gMomF74NWlFbpB+3rVD1
OgLYVZliG2F9Y83TUMq0GEHLfTrjM04mwbgi3B+z1jAC2d5kIh+s74WZ3khTS0Ku
zMBSJZ2DTv5bdlufvp1GEdugv/GwG0pO4xRtyM4I+4JA+Vq07UNSdgOyuOnVVYyb
iI0uclkORVTaPveg8EJ3fmYLZA0s/9DWCg+s7p3nOti8Z2dmNSXM+YXrgG5MXr6e
JF8KmQYIfCzIVf5sVqTjoV6rZthR2vnq8MV+BoSCndHVuND2QN4OiR3C3LdFSKhk
3CLPpmgd7HJvoLzNfT+3pu6p3bV+TlmsEkM5FPgAVXQUO/stmJooBQAHMNIJ69/o
kjzYPb3PXdhsjKrcqZfgQRo7D2cC/HDSyE9gzob3rxkhcnIlm0ixmRbpgV4JpQNk
5nf09k0821+2LPNsMysEShh4plU3yEopwCpmxcPsIU9kC1aKVO4NCg112QLl5Ucg
OhEpQNntkBrJ7uf/nt4ukhx7Uh5EmcqGJRL+ZyoFFv12Jgl6gTJbx+Z+o3DiGutY
NajXSW2rS6tHeoLPSQFyWvZPE8Y7e5SXNz8H0HJ5niE3BLdMfTi56RPjrYA1LTk2
1d6aAXPYQrXCxNfyyVwGi84fu9dMn9B9HR/G6pVrj7yaGMHdo73NzDFFNkGZYNQH
S+tbn9GrRmYs5Fof48yfs780a6Q9hfIT4o+Ayo59a5sfs4dOzCf+iRnS5/vUUEr9
tWEjFRGepa6W0M4Ohva1bzoe7ZG3sSuw+4ULUv1GRH3PUSrwDm7xncSlHhNUjqFT
uMjIlYS6DWH0hfyz5d3Tp+ZWB6tO0jDrVgOTl2RzJ4/qH1Oo1QwxM4KOC7CEm/0U
i7bFvfJqUGew94WCnIWe+ru37yQK65SRMz09sB2bKtkCAHAr4n5dzAbjtRgYHOjh
zi9yZgTECypGIX/7qmnvqWMK9yo5kQKRP6rkMwodOPkdrmZLVnsRvYFoCSoiksym
c6gpHfuX3WgjMT75IPakYbRN2oZEReYBzGmZMh8Wvdxhe0lHQ1dYEWZZU97ge1Pq
wnXkkSqT0u6gfUoooe/fXkMsNIaCgEXmESu6HmYbL9hlWxtQOXR0s403cJruEXUU
p3IYXox9+XwlJRlX3hNbtCHrs/eu5ojT5ARDxngWwkOmvgA6bjYv24/Z+2FeKeNY
87Oj5t98L/DVE5t5qummtXDGfBUn1HqUz64fuTda70tX7SmTNOMqMl+wYuwCJvCD
TPxs37ISlEf3pX58gZvH7JF9jF7UhBfj3f+oE9pWXQMIQZdqOn3eqKQGCFdkcdoO
cHrN8eXcVRs06QwoSSXmPTtnyvcplxYf4A+liPuwYj4paHyMpiHXIsuBqnTbdScN
eXkBFXemUdY3nEgQFSnJ6hGySYEYWG5C52j25/HIig7NKBlVQQBCP2lg4Cwgit+R
B9xf+wVSGJCJYi0b9SZ93gcOBX/oEUxt132OYP1m3f6LZU8sq48QvJelGKCu/VDc
F0uyGI5JPDC3ypQ+n52ycuk9lpUbTgFG7yMQQ4up59t4X50VdqGTTEDQVVLFPLwf
g1RSWC34JaisEVJU3lNE96YFHAkvJHbH13gYzDC8Pc9Zok2TkS319hhI5BfZQ4+N
Xwu/qJBCwJJED6wfTpVjXyc/sQlOLbHGT+Xip+6WOVv4tMIq5n4LwVEp4eUAl7zl
aegyeF8AN1YPHhiswmOZTaytlckNIZN7/A0DoTSfhQmZ9KZcXUnHslO5Lxkbx2aC
Uj3qHWsRjdB3uaKkC3kC9aCvmdf6FG3ZK0sv+oB/C/69vLPBR2R8wawpgARYJkV8
KhnfRxxMNgHiq1GTFo2ri3pQoW0wD2CkLRTkNf8joTaemtr9RG+xyB2qK5b2Isqd
bu65G2LSmo0kxSOgKicTKZ4dnzphNG9bhWfBr1bDpMxFfiGvqA8zxF9FMRGZynpU
6L4RfGLcJeGrP1LR1S6PxmbYfhhLmvqqCRpZt6KFqucynnc2huDmctLJZVzWyFtK
vo7xpgPanKEWk9DZMmDH6jeb+m6Pc3rEv3CCv0BYYTnaoMVcK9VXSxlpEv3Xx6u/
Ucdf9KbUxK3v0vPUVf9aKIddy3EQe7GImldzX6RVnHTOyfRNkiAb8wDUdnhedu03
3Nq9wX2WZFURJ06nO7UrmA8lpwrvC9YWBmZWaBjaIS+47SN2BlqjMJKe656jGr2+
HsgU424AWsyvtblfqbBqqM5qzy3irWy8vVgtadw8MOdGL/80Y8NtQUAro/4tmZ3s
xH73G1Gksc34KyVHFeN5tIXIiBNJo4BR4cEW6fqi40jn6eguWjTAPxHOtovkLUkj
TPhUhb5bweMmcm281bVXoFZ09yH+nsk7kx+Q1hDlpYoqpLDJQ0VzeKw83/6q7AoD
DxWgnCjZ6sH/qxh1Doeyc9rPUwlE7Wvvkh2oIXsGbjnvLxXGjwwOuyDU1uK4F99A
LWcN5zMU2Y7n0C6qC3BItrumaM42DFiQt716JBA4rfnjUlcHLA7q7U/9VxrA6XOg
zX0l6K5sNsouJkVPHaC5sIoBmLfSjn+BqX90SvfA8006IhM7Mmf7HOm1r4IAoYvq
FUEX5FSXshIZuUyExNR0AH9iiqk4xK/s6vUJrcGeULCQdJODzfvGl2XUnjcGUXnH
phRVuFEu+zFuf1ytgDTqeUlUY2VGSmxa3OsU1nFXD0d1v47t985yu4IsgM0kc9jY
lti38iuobDLfe10gjNDlfjyhW9my3+JvvCxxBQ9zrD0GmHxbdIrxeWeCnVdeWUHv
Jr1nGqCJhOCwQUubTg2GkmStNygD0nFW9mZ6mUE1Do2jJFm7GxnIIbYOWYa4G/a2
nV898fwn3IQVeNNErVDx7sPOg/lfxlJszYAr1v+x/fRjYFA4RRvkeu4EsKNP+73u
qG/7IAmKTByiSpERzj05Hr1+2x/1AP19cnnxGmpGK4GJJ4MguBbrChCZPyuAwANd
WHv/hRGwBYw5FTpqkkRKlZyjX611avdMMMPjFC79w3J8yrcOphkMoSc1N4Ya68Tk
/UVOAijAsR5j+md/V3S5EAc0+BnkvdIg/UCjCAOG+KkS1CJ5645T1z1fgMeuseEb
u2wkWYlFpXWgXSFJM1xJZUvySq/tNWpr2EiihQuGXnhGwUGdL/X749zm06bY2I3U
Uq3Kk1cI+b4pQqn0S84pZdWDmhyyyusafxUt+dhScr87DnwkAU1zAyOXporgzO0n
ouiO8Y8W3/V4+dHKoEvIi6vguux03WfgLY1xvsbUJ5SfBc/ziJHyn1bR7dHDpmry
z/VxMweO0w3d46k/EfgRp3jWcRNfFiBiql0cn/Nz4HGZjCHFmCcgZMSCMbrt+pYN
UO7USq7nbiui6exn0+jcvN/j8r+Bz7V5VK2EIbP3Hw8QDUqe20Ey8yt+ZCyHGj+6
afIxD8mQwtQAmNs41Rex4F+BX39fsrvl/Wfrg5oqvHipMa6FUSd0QCUJctOSxSDQ
orThuoXNlck3HcgD8u1pqoGpDbRT8tFfohQLkcuDkdQditPU3QZXNwni5fmJ33Ip
A3/FvZGqNbgthERqPSH/f7E9Hcc/xEiHftu+8uzzBex2bUV7JgSRoGH83CffsyqC
1Dhb7yIDPedja5pJmvsli+d3kKIsmf4Sc19U9TxTiGkuTyC9j4azxe+jC/17zTbF
pbRSdLBndiNN8od4hfGE7aVEutL8IlMegR0flJZoG98EJ+hnUPKEt9upjxafCqCY
dsTc1CpbSdqFzEiqZx5h26w1G6x9/9Xe2KbudvQsBcX29WxraMfViRdhobxEG3GS
NgQZ/eLl0itvpG2g7TwmZNr+NQFuRcePXSqwc1ClrVrjurQJSqz/DI0fZbGLYsP8
cIqSALs1RVZ1gZijm7T2hmEj3NoZafi+ST/vtY7NqGjuZWbIiIUUUk2JQMA32kKd
WKElqPCMiFvknD7MebyFudHzUyhfYyfxz5tb6EbS3IPqjMO/X2OYQUOo2WRpDjMv
kr4NtA0+aLHkpnY+gWT3Hlxy2htcO4RLaQithrHnNnaHl6aJLG3UJ0qqNw2/rEN2
x6tbyTMF9Jesc+QV49Z50ZzDbmQrnnP4FOGnCVdH2CPVL4zvCtvHikofff0wfz75
eIjZfyMNw178a5wTPlhQy5yovM4c0QDVaHNONvdvo9wTZDLB53CGkChb94qdDKlc
OlHB5qwS/BQShXPfbY8D+Ie6GHurr42ao/BciPI70z4qeEEzJK/banXKh40Nbq3S
eIDO2HDQFFrltYtCs5eBu1cn57Q42+eg/uIDekJOiL/LofvK8342wxm3E18uFwoY
qDtbfvvAE1Yk+ntaAl4sTw6GpEzf4Xs+1zMofUZ/V/bmFY+1KYCQgpLeSMUrylW5
IwCbz4mjWnHNwHh7EuF8Bn4fuYDex4BI2R+scuwhZrDxbdV3Ot0skzVTr3sOhq4k
I5B0SPUtL5RL92vXpJzZEpY0Jj08F+psBu/unmaYCRtc/KhK8f1pbFwc/IA/T2Gv
j14FxNt1Dkbp1ftrmkT0ir3JoQOLlMiRiG7W+rZ8mBf5uOE23NRDSeT7ZC2LG+wA
vJmVkpLeAz3G5FypthwluH5EVd/QVdZ2a2u7GZz/V3qsnQ49595a2sFT4PmsDT3x
BmKFe0zD2URvGxdKZBovn+m0WxzAeuIrvtbD4E0qFq56eo++Md35TPkdrnDceUtr
oCmX72IkTnpq69nJJWjfyzVOU7kDK797UNoY4RzHnDjNHa7oMXIqBV7plR6RfYR5
BeTp0VGUn0p98Ii1yT5e0pJ4O1tBRQ0t96Zzb0vknRihYXCSTOQWvufeOWCooEmg
ApImlgDHfYLZCbtzE/vtryewPdGN03nKXJYzFyCmIwqPAFHkg5TEjkyXFT3Ciasi
VzpZ/J8QZIDsk9oT5nyozflBpKrVwTABwLAAJRk9o0B0W+FCB8/mkQz/zH1Q4e2d
4TXJOvyWY464dUnqkCRx+oP+DuhDvo+GXMMoU3oWGX2VeiCLxFlWl3IQWL6NbAY0
4hckbUyIrwe6tSdxf+o1b9dO7Yl2I4jMVQjk7kj0OGOn3xC30VlX+QrckH9HLKhM
7eh/7rf8ZzdTXcDWFXA2+6WNuNB/Z1EwdOHsefn1cwE1zBJUs4a0Dbr/b0BPSa/z
MD+Hgda16hPj4XMuaqi+spIa6YDuzg05SJsRDjXNnaaTM1j36dE2bl1hM2pLhV9O
YcoqaPKajrMbR9cIpelYy3mGQs9GJQwOjgOaMu4k+6waY8+UDT2y6sR7d8Nb/sAm
4NfS4TtoUFKwTmcJEA+2VI5pRWO6nF/gFnn3r+zkHWY+H8cPcgP+7xfbvagSSpXi
eCig40v/1W08Vs6mlTyoQ6fkjF6oHvWnx5NTE9lDM59TWYz1qqi6CKBVZKS32XNF
o/JjZZVgQrTNToutb/7nG7YiQlMPrDYU3mgUIEyajA+RD7aRxWjFFhqYiybU7AIj
8OllfGJmSZddpaxqUsSpes3GbvvfestpUt1IuXiKgpFyEo0R2z4oxpfSHbPM7wah
ShA3D5/sRj4jZzI2p1TPCDQLdZOlxafKUOHRtyvJiu7oeXOL5U6/odQbpYCHkEAw
iwLeWnMOiaJ+45TLOhMgrkzFsMuy5o9rbtAzlfSHTuBRgUr/OBVpU8nTEKCxRfSb
w7/TimhzMuVAy4l8wL6axSKNlhRglYKC/Aje3CBjy0QYo2y+sW/0iOitv6t5M7ff
gDdA7tpVD6sZOwPyBKmLOcEwGBJik1EHEeNgklMeBybMxCnmtITI3+MZIRUu49n/
mxYl7BZItmIm/IqcGLAsnK/+M3sriOhx1RkB7CpE/IxQUoFZLhhdqNrlJWKpazl3
ni84LiStSXruZwFp1wew+XH6NHwzAsGkNT6Io8kvmtFQRQK0VYWT80cd9Q4C7xrJ
208GXkX2d+jUzwNLvPXPCIaLkYm4v8kcd36Xh5jBk2z8GfXTUn+Dkkg8M+1J8vUU
D77IqQNtdJ2Yl8Pvrww3cuAK2q+B9wrxN2qxImYowzoK7av04wSFD2x/RSjZncw9
0ez4IoH5L+LymS6VpiaPqAM0Jeu3hBby6wjVDQEfjcWpwXRTZwyO8cwmS0pJ6Nke
YiKr4p8yYJUhGmU4Zinm4kY4h7IE5W1tY8sciVZ24LsqpMwuCNvuVQCoY6CBmt9W
LyDy9j5WbzoOMekBBnIwIOM2AjjVzi5gic8JXl9jyUGeMdNJb+zH8yUTUde1qnO3
Pf3NIz9WVkV3ZPy7BSzL2OivEoQlr7FdK/B6M/Gv98kHujHGTp6pe4YxaWteIn16
FkDkWIFz7UTdUpjpY6G4a0m8wQHdrm7DxPN3kTtCLnCBoWr/IPJb/ce4ATDUkpP1
5rH44vC65w88Qgxme6HLaQNYlgWNhFAWfbJqKfhSx+ivdl2mmVF2jsCoWrGSl7Qz
poA58ySfROYFy/4rnXRq3f2AkvQvspG2mUI1nKki1t+CJG+YMN23qQ78TtMLyO68
2Z/Iuxdg7z74mvbryhXsw6jGMn/lsWCxUnKsh9wQsXvDQrscbuq80l5UbKfsp3Ap
vLgLD6UELcFwynWC2e9RygifmVTFTf1YtkeuAQvZ/B95V+NOSYj9d0pcH613L1Vt
YaWf1c77p2MSLzKBTC+qZNYzGBHiMPJPq2BCMtWjr32kikxWXHq6tES0G7iMsTit
fjDGTM5fKaSfuAJ8IvnPV1bzCuAK6uUj8h8PAaHqT9fRaZOtP487uqzqbeGdnV89
/AwKN2P1DZ3ATDiJUrp4S2DBtaqxYZRwYaDgCopcd8LNoPTlW9ND7vpIVjRsbeCx
gcaWxcB2wi6I3vAU4RImuIk4H7pvx14PIjs/7oaWaDSPwu7tlA7twSCUOsdTdaCe
apbT/KvzIGeOD4Kv8xhda7F94BdVC2eg5M+sLNOIZZYiATkRuipStklLXGzluPFi
G2SSwZRTrzmquslzYU/OrSdn46DeCNmqOF8O9IKJWehTjQs2AH2biYuNP25XlZuB
ifrq0ila7uvPF12uJvlR++kNmOX5R+7fzlVILzgN6/IQuApCJtE4yCrnNKZsx11k
+t7JiI5s9EoGvP3jYYlSTVZNEEASEDq/hDGm7+Zztef7CCX/83jl+873tLAqwKaf
IcZZX+7ZOiyv8NbOWZaLTqiJYAD+zUo0govFmpN3R/iOQgfMQih4S7Ph0v2v8MPp
w4LDQuTEgUD/o0AJCGRB0TzU1Yp8NzA6eWJi9rXuyf1z30PUidG//nRhEeRbWeFV
rYX3D7OD5MPyL8y04lQxv3Fms/ae+PLQ1u5B6XO2AZlqZ5C44uaqFP17OeEWmePL
C/e9Vtwt4EpnwE5AkkGkpQgouOr3C+chSmzAgELS6JUot+lPKo0Wpr3OFgp2+SMy
qcgQquwoKsjZCgkPqaFwRXamAU8eiFkjKBIyhlWzaPIK3ujjaLQvc8u45Z3pNlD5
hcusem34WH3sG7x8QtWoZF0d9RlOqX8wLfe06Y6C7HgeEpO6TvVUwFQEv3swNuI4
ppjWi0c1M7iPq6J1oLFYX+7SGS26/eEEqrvf1uJ1DcbLCk53OXG/ypgCrRb56Z5t
IApYEBiT8RZzOUmP81DdsRzLy7G/LBiA8vBAAIinby3zzzy9MRfMZJ6mS2DcbLo8
2L0MsGUaJN6jbMSVJfQYbr1eNrwGyLgEuDpRb2e9HOaO1UwxqPvxHbYoRYLxwTNu
QRdr0mKkt3YJkFnMjYKzx4bGuuQLqU2/5dh/XYqRZMtfGCT5TPQft6hReKHvMn1V
hOUNR3VvVR7HGCezwRUcyxbQEYnCvvLZNmSQWkiT6OUl6ERqNz3kIASgS13xlZat
t1D6Eehoqwji3kky/s28YoUFiyTnKwXSHRH1FTNCAE6pMlrxt6gkKcWS8fpB2i20
2nyK+1ooRBTvR/033i6PfMg21Fj/ygkXMJLsEznRQIeGlQUVUsgyo7iRdn8VRcou
F/zqu9kgg7RVH7jDj6MnWGjnlB6Ni0NpcUIZ/lQ2kjctXg1wy81pOims5lhFtKYE
TIKu8+Z3zlotHJCQdf21N2Nzu7z69bVvCE050t5B7ABsp5i4hK4h2AdnkxPme+CW
kPXThDSKScDUBW/X9Y17vJXfvfGTq5mUuebOsw+ygic7G3mSZkLLG1TqXbDseFGN
IkdYh1AAebr7FZK9SSoJlGHiONvUoHMASZf5IE0X8ELCSoWd698P5migSPNpaIjn
SRtxBgEnjEhzg7rdBfa78SiijXFFKNJgNokrdYji2acAbem0ZD3qR6UCa2phCYyt
gd8rBDxECCX0XVHYt/ws9xkLztDD2fIL65aQLtJNKqthhgBdj4M08jC4fFzyJZP6
MrxA6OPR07s8XKtdKw1ZLw4+24k2ZMzYu73usUf4bfG6SU0wIRUHuYdrdafNZHyJ
r2DTS0L3ejqYODx1XoJtnOqVtFPQmG3YvsXQiy3kzV+5kli0WCUStLqnbMQHTwqf
qiOFcHHmUMFO4QlvOnJ5yI8WYz4/zEFgt/HroVNfkAQUsTORdGh0zs+li0W2wFKS
f1EB/dhbXrp/Q10WMPHvFTahm4Mbdb86fKJZMr3Lbdg6M/zydkVz1mq4yFE93bUl
xKTuvKWtQMQOyJ73cd/fxrb+CWe4a6wVOs1epR6acvHErYC3CKBnPkpsw1pfAh0I
4AcmBjm9B6mgaAhTL6le7afEFTWSHtOk/9fA231iDpysahpoagosXbOmTwnU2kcZ
3RHdl4Cw3QhiTvcSGMBsbqCCif3IkC3G8GlncO7fg162qnDB213M2cJvWpGuy8XP
LDh2GMpiVRpivEWDj42v2FCXkfxQa329ohnFn4XZH4SSZmIe9Ua21lnVylJ80IWb
yMV5+eJ2pLo9Sv48Aoy+KpIhxqNB469zW0CxUt8mNzvmdJkEOQkEeoBzCaFuohDL
ekoiUTclgH8gDPETWaMSi4TafVYBXJPc7oLl0fRP18GgFXbDOqzgwXLe9f+5iv8m
D6b6JtrTweV3d1NPteh6mioFfgtZ+Jf80Y/7NKbiVmgMYFgZCTP1Af9D5xArr+fY
2Bddo94pq/DKwR+pfXKMHYQLtnGP/E82sHq1qRu6oPunxmfUVJtP9yKO2ikBs8ef
AX0EGjiZ59/DbSwPfWSt99nqBd/SO5kV9sWZd9mUGiOShQ38pijYTBeSiKDaKOsN
yDjT40Y+9ztkfg7oxnAL4vK+ziHE3ws3HN+YUhFqI0v2df9HXoVsbfzLgLLTBMRt
DpAQ0ZXZeXrJ+Lt2i9mI9Et8hnwF1PEBP0uU32GpaqzdFnuDpKykr99QiFJsiQtS
RutBTogKhFb98PKq+aGXFkKXYpZDl3rXXf3dlqgss5p8MjHDs4hc5r0aO37dI2BJ
PdgX8kNArE2RXJikPaczN8txYjhKAmPcDfeeUZFZlOYN4H4+Eurydb1+JG+Wf4aX
rkk0BC0Ucr9UUQZlEDnxVVMB8Zbwn92Trfo92w0TmeB1zHVpuTqV+EJuOYEoY48b
mveUOiz2JEq/f2R7rdfDSHgp9DQ/+ueBnurOKJOLDieugBSVHmU1hjeAFyU9y81W
e4tUIRZ2An7GMZfJz7hPunGt9siLV5Aooi2QiJvYmNSdqtHCAU+RYGddISH8oRJR
o6PqdSYkFG4N43NNqmRB5cN6nxzukQmfc0V8ATGyrDeHptUCopHBWwi8UhHd/2oj
QLZ74BV2ryEcDXINuyXEFQu7TUgpuF/jovtRV7m96DjWS0QfrSaZJTm9aBfYiiti
A0hSyZQ57lY7Hyhgt7y4d23tJRPa4Np8Yffjg8S5VNFodYxXEPzm6LVR/Swdhvj1
TGyBp5awHqKGOps2luIbCxvBr3/ziDitz8uaUq3QPz18dWafO5a0Bl14nai0vtNq
XFLSVWN+rvwYMfHJNIHOLQq5SAKuZ4pVXnkVWPIfqWsEoAVl6Ghat0tgK8nnlnzw
ko4VTKi7+f5jij5cmXCuRn3U4ARWCGy1sPOZ8jIa6kCAkaY4lBleLBFhBuhh3t7f
D1PYv5ZUZuvv7Wc5Dti6jjI8Yl3hqAyNX7AXSpTfhkUemIaKJvEtOrljnJh5QRzV
GRQI6jO0/9wa7Q6va9jI1IDYB9JHrKFPG3hCwDUi8TWwyAnu+rWJ2fgxb9ANkOJ3
1bHceDnGTByVS46jxYS1It3zTLqjMhSygVZBMr8+Ro3TBDPVxWCySPkJ2AILT+At
Zi6+YGyO0qZ9flYl16/Sziph2edbsEZ7J7r1evVaFeuVTLI0WKPdvuP++0V18zIM
4FlxuWGcskGiKMRt9Gzy+TnrOAx201dfkDZyA1ZHCOfBar66cDnr6xfd+ao/FnUc
oQ3j3fOfYlGD9XO/htGkjXMSh6Pk/ue5+GaD4n6sm9HmGUyfog3e6mELGMBHptH0
19LjXnsTNGvjGI6keQO0d4H8GGnNDGKPrV5wusjECRBRoZoyuzKPyLvDJDy8EgoP
L0S+1NY/XImJwJtOPHRi8rsDBSMFr49Cfymo7eYVaIJqLqHmSqt5wlWRxS9LbbkJ
WFwLrq7XarBGjAZ4HEjQKzD62wTt32eVVe1a6TSANnNvEivsr5m9ImHhF2GQ35Ic
IRKGmmIbJP6cU19mLw//b7mmYnFAW0/NXliOoNakCY5bJEz3ZUiOSODWJJsAtsGq
p3Kgu1BYIwgXxqMVBGybitLoPd9A0V8/yDdblFtGu3zknFguEc1Lm+CLTyfnAoCB
azL1V4Z4ewes5kSqpLO6sq0AfrefNtE5SaKPi1bh0XTPxIKNI/CeH4S9JB0LVl0x
g1gYouaFXqA+QtRt2bTZVvI0TROzyd0MOPXWVCFboW3UHHPvm2rCDoUpvbQvPIFX
rcRU38Q2DX4jP1C5NIHMQE0A8od6Rp+YgS/qCaY9I2LtQQ7PR+wVIfcqTtdqFNHY
rTWjrZLrUXJhnGRNVvAKEYX1MlVRYhU+uvV0dcbNQkRQ0wm4r6JWsE72S4dejGpE
/aNga79S+o9XJMMfYGK2oKjMpuI7hujZNyOP1ruLnSlGcM+GJeYCHQ6qJ1hYq5TN
b+x2T+VaQ4L5EUPZhUqAwe+kVS+3LFHHe12V/6U5O9uUOdRSM4YNszK4otAh430k
1n4QotF7YL0Vx/RpwM4tQUQCeHeR2qJFLwaKgf3mnRZzGRXT1kt81SJHWX1TH2OD
tmSiulT0oKAgbJpVr+uDIMIgpDu2BxQLBan4WHFxGSG/o9arBCXsAIl+u+Ru3BYl
8ycIsAtqhuhgkLCnMfV3O3/VrFkB+Sm+n6L/iAlny0qgj7+AcBkoXhE7+fXIveD0
nBClBoet+oZd5G8stcHfdQsDN6tdClTnj2hXxPDgcESL8Z7/OgBuF8tB+00KYUOp
0by/xzQ/qn/NpxmnDhZ8tsKZruRgavHWeYpP5tkKL+T/e5J+BhLKudXA5eoVBCtK
en7lAN7q1CPXfYGssfu1Z+T08h9t/b3hravyDOIIdao/olHNg9ML5AXh9lets10j
H/IUpDlKLfcj+kEV7KGioal5qFaZhfzEG2KdqtJ81QdTHu5RFydNtPrbq1+d5Hev
M62z8ATD1C8LoNXGX/gkPj7t5GPRet/r6/tLKlWRhpgRkHdxApyH7dKX8bw4q8Bb
U0H6du1XZpU9ANfPm2fZcVcQFslpvaEj38RQ0faOS+dt6kPMwXFy2e1w3nfWxOn3
4KAYS+IKEidLK1qFPRQjDUuLquSUK02bZhBdOXQ6OEGUFiLEHCmbBGLhEwG00YkQ
UO9PgUBORZXaXryo8f9Z1BHOAkD8NXGXmT2ipRlj2T0prfTxdQ+/vom3eGo3s11H
427g0McM9022YZLKMIFiOvg91kNun9WzFwE/U2TNCHj6UrKBREuqSJFHgneifHv4
aL2dNr6B5fIrwcVa8v5SwAshi3+GWt/oKZsiC14yKVkCTwhoxT9Uad8nD8Fi8i8C
G1tJ8ZvHkMpbzqXWUe48MWfsTLmOdV3kXkFRgjZTQmh0A8iZXoFmM2Xykjad/of4
y5Ca9jl6aXsAuJ7hKkkJBzXIjR9KTZTPDcLInJ6cZ8ds8tJICMtSYKwMSaFbcHVC
YcC2tJslKCjK8NFc8a7D0sofEL4FLapzUOgnrYrSt4uc7dG5b6sNlat059/Wd7hJ
JxtOy+duP/INhVCyxBvC/YOliniJdMRhgIhQ8XGQrtvuowGzYHcBlWUAmKwm1vT1
mmQUb9uiIAGr4rAYWcqAA3d2lEh9XBXirFym50Ya0vvSxvdWTkzaKEfid1EiGJuP
Fhe6IUGvwpKbv2WcnEhbTL46YGBxGj+zLTOvU+NYqFc8neSRStDsITe7KtNvk7e4
gCpkuqUKtcfGXjPfFDHkXMoEOYLwPWEH34OLpWCTJhoFuf7CQvdXHnvn/AJoT6Dc
hvzDCE6diw/P9QdtppbKqxuVVPIIuzonoW4SqwTBW4G2oHOOr/J54HupNdJp0oal
JEknKZoCVPrkNEfV4u0QHsKQsgd8kiUA6jR+RZSqgiFOxVY2fgxqOSU2ctWAd4qA
doIoOwfL/JZ6/TbTQgnrZWlVuCDh0Oo8754ucMhupyFwPfJ/kH9k/hT9Or7DxdZ3
3fVUovaBf5YV3ru4HERvp7f8SuiIKdzyDxXLYhLsy5IYFA/e1evvkMmVeYTJk3o9
1hQgrNIv+/74jp15haAgqRtbK16mvFWuUTERUByVM5vFEyRGNZzDInJSIdRS32cD
83u2r6OaHAB0dvCcAvbpbQ2ecnrzYW6d/doXRqwT5/28zACQgYdEJHDYFJH7iEuH
gYroMrMdpxnlK1XTw2zJA9DJ8iqWgqeLTi7hpLrbXDwdtdKxlb717QIba9Q1/lEy
5Lk1vlC9CWHNinjjBlUJhEoIEwWHD2SAiCN/u2UEz/XjII6PzLJrqqajLnlYAcgN
1xtTYD4KzGw51aLInyd45930ck40+80lGtLNoSw2IPot6ALy1fgCywEbc1yp339o
4/FBAFZX/Ru8wdwCikjy/f2v9oBN8HvDsAUwuoX1UC84mOV9DtxqKmV6DKVYVWpM
W1tyReiM5LONv54+LsJwW7h32q19RreL5UpkSXWGQ5fHYt+gz3w/sfLU6tnZ4u8d
FdaIk/lHKuljkldaNti0cPCctfoOHyRJQYYzFzgefsSaLCixA92BoPq2PUJAvzal
N56LTwMl15sEg0hySNPY9ssEQK7tM7Nu+q1eRcwZUg6XTqK56wbxMdOH5ICdMHrp
GQoScm+Ne5bgLnqFOWdkxgsbvhG9pAhvS7x9RiBVi6SJ6rg8Xqy6Fyn8jx9HcoN/
HGW4VdizcNUN/XYh9XeZ3TvWQ+QOb7Zqoo6j2AsBhxzHTxHqZRvgXI2cZwLfKGWd
aqTdpUDzPys2tPuUntBw4v5PWkbLHTQGf30MLLAuKW69VGUxuTnOAOI6FMFS6y42
mdLLawCGUZO/zACktVZHTLM8FPrmuKHtObAII1pQHO8hUJXPagZgruXT3i2/tfBP
HDa7hzD+ser+DyYpBst//xB0X6BqSO6OXQUoteLhIFmz0B4Cp8SXAgcbGkeM1Dc5
gA5CFjYFoDT7eqFXDVmGlSqV67O23ywyVnJIeHHr2h0Yd77U5VaVpK95xRUytf5G
AerPtHH5EKbhEyjBJn0cZZYInsmqTEgfe8QfblnPU5NyMjL2X1DSAoudpHlQ+rqp
/mPe/iN0z/dRAGiRSvNx8tXoOBZbMSfvgd20A/+73z1YUjhPAz5Yme1W95xZTG7b
zORf9CnAyfgdM1vC3+hnyQulfIW/4sr2tP2u/QVN+C1icHC43D+fHfs89vw+/gHS
paMbcGmjS89Mn3nITyTFCCRIXMsjYQ2ODIh9+QJqHoIWH8zVzjntd6VzFMV7uwtf
MzOUwfsmi0vIRAIVhxsUJjNZX2WUmH4oYqX9nyCssdbFHt9DwNA3mQ0+73hH+A0b
kmFY3mROd8wRT9M5WL4xBQBPPYM+JaIJYLcY0NvdNyDSwX5nJS1VF8RoNWUPpVgK
TvNd5HgtGqetSsFWF/aOA0tsApAaDdf5Ej3XyQe2fzq2AwZLxBncO+n+4H/lydgd
+WyvdUbDzHJzXhiVv8AfKTNOjsR9sVEY806lwj+0DNxsjfbYGWARLVdD4s3KEGaW
/aTmGf7IB+iZ4Xr97WvaUGYM5w0Yt4MP7+Mfd0y6QkeuVHXBO2+YuQcpRtk+slRV
9OgcWgssbgalRaMc4VHX++3wEXOrjy/Sb/1F/bMlvxoG1UlpeVjWIo8x3I0Qtk8X
n0aRvcXIGZn8GH8MMVsHRpfmLq5ngZHw43tD3ULY26PBA2UhWjDtN104RotOvosu
vsOuHgIiLNOukNLdkCtM8RX3TN/qkz2mi0oo3E3dHBDzGHh71LYx0sanLmbPV+ll
QxG4MYf4/P4FCwbcrllahe4hfqk/ZuQ78VaQ5lC8QTvvRSepiteqfMw6iBFbxqIv
ZMLtNyeN7qt+OX6rxyT0JO+owNJS7mxp+V/gSZx2bN/QqNDT+9G+6CrCWloAzQTO
JY9UafiGgkf1kGxwjktTGPVm9ruyJNx6BOxeTbMBybb1iS/kmeI2EAQ403yD3Sc6
GysKrI5eJKqUzTLZhYxiZw912T/WTPY0kcsKVOt6ohZxIrlFbmBJGxFpyCD9ACU9
KXWohKDtr+kfFzhc01S/iy4d0LRC96T6+r27jK8AKC+Z8LehjRZ2O3xOBWIlp+CH
nyAtUoiBv4MnzDlSvWd/WRyeE+MZr9fzlKfAW/hlm8CStH6yiZw8uHZ2z2oHfMu4
dttXxSQHBOlrWGx22IFNaI0Wd3FuF6jVw0AJx2iy0v3rMgjET3xl3nL0oVrY1wSX
TSyI4dt4xmH4A1I+tcM37bYOMGEtX983nf+AWrehCKj2OW6/iH6f1SOdTVoJMsTE
0aFPVkR3keZ7M70AOvZ/J/Lghp9dOJrKUn9WQQfodXaRDbS20pye0PrX7ZKkJ3Rw
ZovqrR6cXs8dCvInlAqUjzg6EvsmS4t3QLR3LK+IrZMMiPCr93yfWOVpUtA3N7LD
UOZy/wHYaWLdToMUifKh6HrLRbaS8EwhaBsuT2SZM+B1/58QCCs+AxO8QKFGfE2T
7poFuBN+KpdtVgpGhEQb4IayAfexfGkKeqhY3CZEzU/IH65WECFoUtpXTZlNgPIK
GMWMFeLplO1sINS3KAi2ECFIxfDwJU29TqrNcQkkaODJoySeMumovBzsZdPwzCHF
hR8s3cjzYcQ63CLbIoocKV+wTgcL7Nugv4UTrn1lI7SAkb8dhTRmEaaeXHXoHSBo
r+07fsGGjv9Gq4L2vAVAFUKeA1OeLobnkmpXfXgpK164awsogPsWPHqH9bApavvQ
r8Nvl4CxPaui2eoWefktt38zZutYbJdgGowGUeTUWCxP38A+4TklYgDF0/53CRIv
2NCntl3HR7PbkGsxEHFiPj3Rn1Zo4qkC4o/oQHeuTksIwGLnPYzzMjoSgfKICfAZ
KF4/22q5ev7JWYReawKJNnWeHSsAyIxULokDu6VOTmI7VaqD7sUFQ1QMHLRPRNrs
CZRMm2/BnWkcpp/DKb6QD0EH/jrR59GDzK0q+F3iSlUzZ15cKG2D0BP1ecTTZjW+
SwpPHW0+Dy6+HklBg5sxLHnI7/uDN5dxBNeqN3mKgvCupgQhj9N47RXV6Rid8IcH
iaieHpqZwvC2PvfQkmAQGxIMwhP4kAJvt6IN1NkLEXDEjQbvJNTiAXfz/ytZZEGi
+L7KUZ+DgEbBdVKdHB9Kx+PwfbYpDZDDLzOoT5/VR82a4JuHCmx6Cy2UoPhQujns
1SvPNBcr34CrPiyooCDyHjaY1FTkryvTfRNqVu88QQbmCcv/OqLRcRt+92gvr2Wf
abYLoDMHZLxgAU1NZgYwBzHXYo7rIYQxgyfj9AzaDxUPYF17NDd2HCpyMs9dIgvV
C/XYwfgKBJ9wpOFK/Xh6Rs6WutzzVfgesJJ6KQxafGt1w0ls8uMKs3HZnlqEbJ41
ncJQMHK9dmsl6fmJNsCfDeyVEO+0CEjzWFuGV37H5+eKb1QmDDeOAUOp/fZNQjjc
K1Httn9gdt47JQLXypXlrVHzn0K2bfSx4g+zU/XkyZ4tr5eUWWIWLCB+vMK04HOJ
syzZ3ggyKmNVKq/XfjEdoFnbw1QjmLg0y1xyPsjWspaNdDcSQ4hmmoWKb23iTv3o
bV9Uj8LELqleUw/b5zlIe3FhtHQxeyZF+ou+GEixl+/v4CLP3vJb5hnhO0+B37ZD
0STUeBiYsxsb+Ek+vZ6y8ffh1EYRZUP4E7uyCOBtsDg2Cc/ZTuRoAIsQ6oi94PMK
rY7jU3J00TapnVnqn36eYJnDdiEwxv0YBGhCj3AzGp5ly6j2cDWT4L0ewTGXB9tz
6uRCQXh7kziMAmgQzuD8Rr5jQR/XNZDV8nTkcVc8kBJTphD19opBi2lCjm7Oqq6N
1WlVFcqDOrgs43CBp40W/JjrQMXR+v4S9RQFcufSv8LbElM9NkEKiB8Fm/6JBMoz
YnO0NKUA35bztu0U3fpEhNY/uRq12dvGUEsBiZuvB8YgAHBV/HWZlpSDxYmWDNlF
T6GzZCT2qiC2iOgDnRYVexY4JuK/0cvu5ykQweO5utt59qnf3Ia4YcO3FepAVaVB
py6aT+T/PwQLzIcSuab5vU8ktBaIYZmLgKwYL7j3jfTfhhqy/9OgSp/9fQMAAUy+
3+M8g/7BwVw7R6Ihd+mRxuETFCbu9PDY2T15gndj0aSLrLbFbZpiqODoQBaCBMtK
6Gb9WAqPALop2RHXHeF0b+gB/8yFeamX/Cz0mGmVOLRhmdmBw+ZXauuQ514TBNPg
PbrQmbd4vfxJp1oIu/L98eXNDO2iU97yA7sN1KObmr2wWlh13fhTNtiiMviQ6amK
4Ao42tl2N76HO4/3HpegdTQ8ia3wyDkrFw3w1byjZCmabioSKbc+5/HntC+2tLhx
GsXCMFzdiMbm+DmTa33qac90FynrE1nbHVg4wBd5G+gcsQjTC2KOb1o3jcV8pbp1
65AiIrpnoG5lrxH7Kd9hT+9iuES+FJeWJlrmqdOt+AzNWALgpABq8PzNNJXrqDzO
kR8AjEI2dTc9yrwsHcLtX61vhMbThEGNH2/JrNCO0rruC8QYH05zC3RKdbLKHe80
aCnrHnBG+Ef5j8Lt564YS3ed8eCYHkzmSMpB84F9yCIE3/ht+4AQIkIAwj0MX9VU
BvhYWLFJ7yhfnLvNYLcH9plphlVE+ZJ/hQdAVBbPtFs8X1T0J4vFrrAJu70JfUwY
QZC7M+cT+Pz9c2m4gdmbRAfNcm8ju9Sw9zWWHAwz7rPkXxKGwTtnGjgQgYWOTPZO
9fREPHErF7gjGQaUrXER9zJLGwx9prLxGqmBo/M2Q6xoS/oyD0fLnWgoGgJPvbBN
KCc4g+4YhoSGDWCZOJqoyT0wpsds3P5bgYVgcBYeOpCXB3MzOYTiUwlGFGk+7CZS
V/MoME1mWA7FkQQW2e5vW0py87mXQY9NMc2Rk+v3FpiQWc3Fn6SCMXuay3MvYoTW
UL00RykHUNnf3Fe7G9Hj6sp7+5oLy9T0DTKQ+eZLL22+g0qHKGDmEQXzaFmc4Psm
B48QiddhmEsqbsC8w5ykjnANutJY8gdS2IWKKGe+ejx0PGuZtdiyICKQgn87eadr
fiTWoEyTfEvtXgMbUsjWcPv36Mjg0ujoOaj3kTRr2ZPIMQmEasPrI6YftScImqTQ
/vk0X7RHTNncMrtQWxHJw61mwjEFo0MCdfLC44qXZ7wPg+FSVMqCoPkuoGNkPmC4
fR65xN1JpTSUVH0v0POnPLCL1jxLUMX6WB324ZP5qIqe+GmAiWg4YhRLxMafCk/6
YmAdmE4TKQOsFJ2x1kcRvpTBdEX+sHSxtnCljk4NeVEElUkuNKwdVBbN9LB8ZTy7
acuKnf80c0+x17W5aOe/r+A4uZIx2T7eujNtKfcvHn1MrYbkbJvedBdpE61u0eG/
S5oP5nNhmna7D84Mmm5rrAzVLe5qe27enZ+MmvVNsv9nSrdQjKYfqRusZuP6yDFK
x+MnmbuOpSSS0Epok4IuGnsVhCJxDiIJejdrJAe+w2GUOa5FBYWwXSPENVBRV1aU
Rz9u9V/3EdsAP2U8kpMtHMuQCsS/CMht5qygkHcfS3dz2TR+VAsU4dbl6zZvbrih
ycnbfUXnMUJ1MvYgck5Ibiad4WKjPr+PD38x1rr0oUlGJsqOmxZUtOEbxgBG79W6
KYnl5HCbBJXb5lls/YCIW9HgqQosg3J/3Lstv1WXDKi2YHAybgr7VIoMUNyshprl
gOZ75X0fNTwZSzJ5KaaW82/JcU2mjPSaxorqv7xg+EIHz+Na0EDyYtRObeZhwzg2
aitF7wYfMUZPnyCZx+IbYRUEghHIk4G6pZFyMR+qo0dAQTLLfrft3i5/H2zPzv0g
0ar4GGKk9r+XVkHThL6kfZat0EnpKCCX77yIB/3TkP1QKlCopmvWcOlwNTaDgSER
jai6vPgxvzFT5QYluoYut+EWk0dIROXWDFO5Vwwa8P7EYzqfP66BX05NDCvYZXKN
CVxcYIi4uhjAESzFP+l4AiGAXP2rAuPk0y9qxktdLUwKjJx2uuMkYZi3EWE0Ef1Z
7plAuyADs6K/DcE3+3WZnr2Pk1cNM1jHXl5Yev37hZqDdC0FYnjREdT0H768207F
8K/1F2/souE/ursS/jrvNRW/bHFU+zBKqOIUjkJ2KrC1sa6oHtDkYepKc8sENyi/
LzmnYSqyBgB7rGSfYsW3BfOSQc4/lrXD6mXC1oGfMDr02SoSUAp7QfQqJ1Dyx/rX
tKzuIwUWFDvHs+7/+7hrG+hgAk+DKu5VS1P4oEijtHIH1QdXzYugrXQwvv3SUo5m
YIcRQ2J3zK1TYQW2aFWAM/r8GOC9RAm+1EeCiAbErjHCUayLDdELNpVxGE+ZNFGq
TbvpkbvX9kFi9+amM2owQChxFweMcbmRNyh0gm19eSQUX2g4642Ik0JkOtIXY6FN
HGgjYPrYhkzcQ6jWVwmEZ9m5MAJYU0DZf2z0Pgbt9eYyMDzX7OvKSIXGwceWIp5F
1k0GcTmF3Hl6VEL7e3uow/FeOc3kD4dEKHSJ0H+klJZNoV95N4Uz6WOHrlcBXl1E
WE+U3U0NB79hpWVHj7DGuzKi0255DEuKiLdTTDPh0NquojGKTDtcBynG0NY0Quhh
2yXbLt9rrCRMNB0zcC5FVYk9V1w/lH8pf8FkmX7ElGQ8ehdh1v5nj42LL83rjLgS
WwPLykqilRMZ5KP9B3iXl5rufo76pRTM8Y5jhxlnAKoRSU2SUXHU6as8IyoM2eFH
FrhnXv1j7MgsYLe4bKlTM8M8jdDhxCaKN5CkbIBdPDM4je6bpqScIr1H4KM7a30/
+llMHuhAc1IVlSStBWDjavHptdWhsoIsfOujBhr2aaUG/8XOAHgBReVKJkTXpKSG
zIo6I1GHRjK1BYJHDBjByCN0Cq/15tUGT3+vv09nc5g9rAYXA+RE9GMnsoec9uZr
rtbUR7VH+QfzXeDaYuTjpWNmsQKJOQLBEA2QsjQ+jnqpmY0lHXjpn3tPKL9H3sOL
I+hPYjrKLwU7poq0kJmw8LGfuZIPzunVJjABkDj8g0zK+jC6Dl6fK3+YLdMQ8wF9
SVAWuu3cvwncKZgfNtH4c0jHx0O5Vv3F8BKMK0vR13U91vFEwA2YrnqDrxG/LyHU
fMD11Ez4n+iokanSKP92lDQukBRZkId1Z2r/U3+lpLZsAOBNOSK82P8uueJ28B5R
VY+H6JKaivapz5GCrxw8hu0Q5ot5nGskqEDjXHDpepdiLKV0JV9Tc+lTs/Ntvh2S
+7KtMQY4eZVMtxRkShy4Q6wpSZ/98XSAjZwbtL0Y6TsWU63aK1h3FNX0k63Hsnew
9+cq2A1ikhHRfBhuvXSoiPw/a3tT/Gi4r9MS87FMXVId8EkWlgU1s8diVMz4bJ9H
bbhKoPKgfGvDq4F/z+UFCN6X65ZocH4LdWmTUJ9hGySK7C4P5DFOuOiF00iIipOd
IkGjuqMlXqb60Y33C7vQB+RsiOPCtiTAkuMmn6BZzYGhYFZnHkfnrObtvmUPA3eo
TEClUkJX0Y7p1bBDwtrIFmhObGipLgNccpos8e0Djp05FlL0rdYiDm/72dVF3FDY
Pwt861OMv7PMQRhStaPWSsbswtSqcsR+oFw5TgZsFupY0ej9LJub27X/9U3JtOfZ
VffUXPqox2rFoH4IkJieT6KTARyebbBvflVS5PnqlURnuGG5EOxnQk9VNgwAKO1b
w4kkPyCDZkyY6PGHBWEGcqhGjtHS6nxbYP/ZSfqjzVu6Uh7TUBEZe8ap/ZPBKkts
7Lczv9+zdItXpHdAOrKSj6e8QH+F0rL655Iy2hG3vgkyBrQdzqys0Iay2V7qneBz
eZjK0zpkUA4sr5RilLf9Hum/5SVccJ8g+FhtQLatXCzifsSNmeduSGCQLIiPipoI
cLarTwidDYVDaX/E5C76IW43kWQoMIIBK/Xua8qZjAwkQ0S2xR3r8SpCpkMnf58u
TT/xQIm9+s6tbBfaoXxo87/c113JmD2O6c6jO9JU8wffQvD/Ff4iGRO9QIXu5cOc
uN6z5Bo6Q/KScXGMQUiQWS7lYgZIa0aPYQLHGbgIPph6TzqxkYR8JOxF1K4XkrPh
GvGZ0nU+FwMd+maxw8ukJ8zGH6Etnxjn4VoZ2fmJWXKSilZiNgyhl8NIuSNtk2GQ
9/yEsiNy/CSbRF2K0tdjBoWUVAPbAOHh9wFzSukX8J+iE0qfhbjgYiCjgGZDCYw+
mCb/LZjgZIWQJO4HE2topFxyYop0dUc/BTF8jruGCrWU4ws++s8CLdbgXhO7suSe
vMSRRexC1jz8gQnzkQmmfQS+QLvaOkYv+faL/SkOzj18KJTA6dr6eNIHdhNYaVe3
LW0gfJoHEZn9Pnbk4COPfyl1yn5PSqrNUznkvByB4xLSqqbDkf75XpTCePAI6lrm
uFAUeRdBytS/u0FVldZYnaXg2lNLJNyXmFgZHGrpjeuFeDn6ViO0MAS4bsSujXN8
UiaQ1sQxrXeaGyqDYz+mtm+1WpfTbPkCQ4Rp5MnBSG/DKu5FGSb702LAyMcUcHYu
WL4zZpqtrVWH14z2SCUwiVN07YD4SofseMZe555daefdwIA0SbeTviyKUTGR0Nz3
CxUXqG6ZQjNt19br42sfYV+ykU7gpyC643hePI5ycp0ZS67azwg5lrGZQh2qSvmZ
su72ETNg9xIrL7/tUP+GFyghNIdDli+ZSM25BGFgIc7XC81YNprnq8hSS05koQne
gMKRMg9eWqAzwDc3qC7/0SYhw/YyIc/CpcHWGmRIFWQjbjndDpSJiWnpvS1lD7cu
7v0XL24HKikeg+WApdH/dY1dvdII9FlvJfaEug+3XMyYBcVPjKI5BtepGdqFzmmi
c14GUnPgoZZwiSPPZZvJ5RIpXxS2sh2HRMbsqGv+KSuFiUfjyCakM0vBEqyXKBPF
4I0oXqsgGqXPGDmgUewMRdToCK1NlkBOsK9rrPNdsZkunE9uTfk3DNY/nI0RCvaZ
9nITEkQBy1xl13RHFq/p5NnRLBeuFNbB6JmROznmyiRm99VqQFri+yEqV40DqpwK
v6u3b5/YlRyIVAzTGSd3KTGDVjZbJvESx+4LqGfD0bwF0oS/Bn8/XbywoQlVFjNh
DWAHrncoX5sDrBicVXF3avykeGuk8OYLcOKZvT2/0WTWBCAd7YzBkhYR9deQeeBZ
GGpMjLeuS7ccIQXJVE46WOymjXWec0qoFHv5nJ4xltnI+dHOc7b0NO44wbshYgWn
A0pBtezHm4LEO/gNeDTKvbZNco3WvWhQZbYpOD9j1jr1dj8onMVgHrKAXwflg93u
lDtsvqY626T1TqDr/UvTxRuMYtj7hh2wRadl/3v+ECz2f0Nb9tpOD6PyWvG19d1e
lyP0m5VaSYShE7cRuNPPgGMRUddH54Wdee4JA4vdAlkDi++tMoHKig6loxWJ2+8F
nucTqon7SmYVkUIjyoUw9aiz3zwqz//JC4OfBV5XjQqHAy6QknaHVKXBzcsJ/zkS
zihGTwcJqGrdp1TccmknLEKTYLPSi9t4KeYfGjCW/Bxjemp+LFCpcWD8BJoYlW/W
5VkcjGTX3Ws3yL/bgM3HZyw0kwdvo8LqKXP2l9Y2UxDQa7NKEGAX78iF8UjNpdw4
hGCisS/kgnGtuCsgUsXHfITJal1pGR6G6FpBgcN2NCu+1LvZrqM5bilikHyyT6aV
0QOpiYr21Qhhn3CxY8bJ86UBgQAGpnjsKTKE21i02qjmISiwNcTgN1XKS8NXf57+
9sgQIe2BzXaMY4ZhHO3O47ZBY7iKAkmOaXPWzAQTuC5Ajk2h6/NcGvxhNCLcUMCm
sV6MAOvH7zp2oqF1SSBitmLnEUIoMszolypP4RcLpeYD+wqX+eRb3vMwHF7IrO7Z
n7RFQoQqITVHxedpjAveP2Jh8VgzeCRWxgE7ewDasn/ffeMPwCo71PlSJKqYFBjB
Ixu+tsyajqLLGSeZ9dXbhmixcZevl/nzx0ceSfRQPwear3fptzoduQskdjJ8a0O2
E65zpiyyzc2CEcblGFrj481wfFJnpDH5KSSN6za4F0LBAE5L/iNrV4HkScRbLgbd
aFumeZ3NuWNWDx2LPOFcq6L0GDR5fyXfiKH7pa6xiCVKsTqxRR/+PlazGoE+JAV7
zXO5+0x9lFuDTCmArkmQe1pNDW7ODWa83RaYyNOw5aNkPRbsDakRi0BUV+5eTW/B
1AVrDizmrrI5JmYY2p328FQZBjfQCC4eAJAgaGnxssOOraC9TFieuSe0XRAwFU30
KwmkwViTpMgbqlwiOzqOvgSSv5uJyDrqPmMkfKHXTfpNIXCUgvjbSV8Ppwe2in9R
2Ug8XWiV1LaWiKYtplUyzfcvp2pw0zUH8DuyEzEic7Q5b2ple5ovVNTqL4KecOhO
rb7EZfTAUY30Pif1ZMtuDZvnIhmhd9xejKavExeQaAHbjEwZ40YuDj805wZiKs3b
of3QmMBn7mMYKXh799UUWPJdo4KF7AddgRHdqOIvCLsSje76u2U9Zn64fXiq7bxa
YV4Bu13bSuudJL0X4R31hL563ISvfHcSvqGA78vrozlRuX4uOXsLud0ub9EHl81J
1igwaYEV9hy0uklRytWM68C8gxwXP71kpR/xgaIO0DyjtyInT3lDUmDZXk0Uv2dN
zsWUenz0+rYlQOk32krBsKRit+2Ae5TNfSX/rVgTrwybKec9lwTzIX0Ud94DDso6
On5ZflExZ6ku+Zv7o6ccZSY9i2LGjQWCsNAsSRvQdYN0ioJNI5VrZYwoeMPzbaNT
5eRH6NgVAOCpnYBpN4AWysdMm0oVPeMQhq3t8lsugn1zD97/VYqypf0bdupnWnVw
Yw+00mWkPedvqgxU1WmJKij5fVRm4B5yKblTZoUj1khGxHcJ11StWBGyjnS79tcJ
UNNSD3PeZuEd4K9+OG8piXZ4uz6jQ0uHlD/J5nAFSJxcPIILlr7Vit4ntyAEKv/E
G/2rM0zpSLDMms42bWH5zTPWD2idFMTZLrlx0cl4HlNXY6mPhNQUfpnO2UOlxq2f
ANB5PO/09R09zbp/4HlUJoEul5TFdwgMNgsAr6gbcD9z5Pkob5vtIrVn4DePShwW
rLuWBICir1620JRjxVNemtncYNhZ/uioNPkkBdwn0qC+SMG3pSctZmOIWrYd6SiN
/GNH0+X1B2KocwtD1Kh7lBxFsbrbMYrlE2eg66eDQnuWmV5JJd9zieyxgJ9ZsiqE
2x54fgsiqwEtsv7LjRNJx2EcwAqAmpU19ykc2yAUeCj8xee2NPpAw8rjjOxu+9Zy
DcF+u1se8UwqXRfH2yJ6Qy7XrmGQxP0TaJqKLtcFc22y/CwtgysyOp3rBzAd6QcM
O24204+P4W0KaMAR/wYNdTfiYLAnQcbQWAuEhWJRUHyC97pfUZvcstF+yJEoRocN
10RDAx1qMJgIhQJtwq373I4iyuNdJQzIS+akSGKJes1ANbhzaf6QT1zuVYq1GnjU
IS7J5MlrSgtXYpOG6kAlnVh5ZigxDIS/LrItOklyyg6gEPbZa7gteukLxrAwbVCC
o9aTlC5UWBPUEZn7Ewe8YrYBLU3d4qdsCJgktXFOsvUbIxCsDy7lXDQSDXlLHuck
avsyfr96OAI3u9RiijM/xwoFCcBafIl2YbiYE8jehU8yoJ+kwI30UO/+OhMtNCol
37KrJGNKbMHGJAs8X1gToiOIw1GIvAJp4DCea3M4GwDVhT+Ajnhb7TLWdP4rQaWZ
vfNOMr/A8BkxzRadzfOZufziRtFZfaDOEGag3eLqwl2UGCz0AnADJVFHShRC+azl
To2chShS3NM87l2SpkxIhfRoXHWuzjUa7Yi9IH5AXiq0BDkgp1AogtvtBefgrPS/
qxtxsXZimifksahpDdfpG6Q/nwo34xsGk5mo81FICvxPadB9Zglq4ykftdedCEoT
VkxnLp738H8JooJfdTBXGBb9t5+BQ/geYRpzh0bsOrpKcmv3M4bc+pzOiZNWXc2w
1vDFK9J5cIAHGbkqSf5Cmcze5qhyIc1rBryjitz5gBu/E7yYpH6zThmA6jxhCjuf
mZX2JEyW9GgxKWUOdJ3VU6jcYgxXVfa4LVNaesxl4zobTvsuwq3OOQ22mYAe24s0
y1qxPBRDe/orqNXhr6WUtnQSPPxi6E3c9vIyoEizqUfijRFyustZR/w6gdShUW5G
RcdVdMM8iptVMZWDWw+tPEizZnAs5s/6G2/KIaOldYiDAacJlD4q2rFT4AOoT9JP
9geC1QhMjGRvIs9LytWaIQUoI7spziwKW7bhbrrSq37mzUYJEpqHmVoITL/DfMf9
stzqd71yuxIFE0IjkpjJXLYxhzjzsk70pj3ZynRwLb163awgpYKaatBAPpaHCEbX
K/5QJEwBxREhqffKsajrxWNm7ASJA0gZHEJdPZSQ5/Z4QY0jMhN+yP2NNkuNC2Uc
iKz7HJMeMDdYPvFF0YUGCVSOQx1CE2POMOxNw/QQoPwGA1Lp4fhUcF+UGadCCpub
VUBMlb/bjnGhUbVopieYTvbNClyN4iavRIrynRP8Idv/yOFkvg+QyVH5oI8ZBQq0
fWCRU69cb/F4ENOnVLhEK/j7aUyXlJ/9Jb+oJByvAktvOF7fywos2fBaO0voleeL
z9DcwIqDpiFOVOia/AFTKKi4LI/U5j4P0LShyQ553wfdwhCvt7JtzUm5ujEQIuLk
JU0BW68DQCD7vo+xofCHxqD5CRYFR11JTZpTgU4Wow1srRnesIgbKIteN2IDeFZD
sbGe2L4z9JHNTiiSv22xPCJZskPDC2rrqe66jm7xnt90MtwVKke0FXcpliukAcXw
KGsxqb8A01AguCROJgWpzoFiEy+kIHpfX3gOCI/jmTxNBNhu0JtcknBZOxFiVmj4
zyIg8J9V+CuMYfdyzWcevP7AG5v14U3kuPSzeDqEEzdK0S1gBRsApSWia/5DZyum
8eRVxbnFif2zEQmU+mekHgW5MAzqUFvK2p4dMEcq9aRRUKwcNqJA5AqBNKEBBpmT
gyWvOdLP30kANAK2OEPlqSjFLXTySS2lgn8ijEnajVuRRGrd9P5zgkP8fCq6z26b
mK3Cc+1+sLLgMdsyN9anCnv0MsTXY2tla31ntgv+wKqjqcTTfXfk3fKFHfcyvD9D
zttmXn+i4eOZvbJzM2tQqXzoZ1zuhWeykhaqHlwMg8CzXsHaTxqyQeuYaLQb0jKq
6mqVD9UhJlRX6FPlzBRwvcTxyntM+HOJliDxhYmEzGAgD7TmRJpZJuNaw2WRarLC
3hbf1pQn6ls0slaSeO+JkPTwRXeWMapaFresfRr9Pt9vN9EpvYZ1wlEajoZ8l7+7
d8L5+Mdomplu2bqFD1LQ3NJlrq33hNcoFFm9fS5VX69bjgOXgkhyL8aJZ/Ty5PHP
itrO3v88bSyuYCZ2oeauHmDKlmkeB7iQb42MRSQgdRc3c8LQ43jOJBrwCw8qKMle
wrysrRveyHoBv+20sXT097AmOoQ3SHsec5r/CycnMmcS8ZnqwJYWh5fWqP1lCMfC
i0/eu6iQ3BfewM6xLQEPavvkjlYzqtNVkKVC6TiFccl2lYv/q6McvygQe7eRYdLo
2IAoTw2xzZ0gjHDpjI1iVCWHMnLfU2bRrl/agpOHlPM7nYjfHyK2W/uOSoFyAPF1
UNAC21qfrxgqAipj4CGFluYj7QH9mYe0waUiuTpEhX8x6yxDETAqRqvZE1G5oGwk
bhYiFFSzQpp7fdGPv5UQ+h8MB0oXTzhxYEXzdf24Z3pOiniVVUs8PhCVX0RKm6Qr
xED8ohoxLrQffo4FGWqmA5cDNF7ISiVMrC5GyMCdsH9iIXIc5D6H4CHaAKBtcZdT
0McLcthq5/pCkyQ4ZeTlJ+HMYFWyX2gq1RtJ3nun4ONRS4CL44e+JfMT8syzuUMW
G1MgSirt5b4Gpp+TH+/1KpMdtkXeuk5Uucy5HhStzNnxYzOF35mTzaqmZLBwAQXv
oBUDW4xHcVL+oF+5Iw3iVi3eCI+1ztGH9QlN2MZ3k/HB9KrwKUZvAaDQ3qXhd3Sw
gtHhxKwXc+INElFlVJIWbHnCrLWmto2EMExt3pnqQjNAv+FS7q2QjMfpqRu5fvUe
Reg0vGupGSwJMq6qIkYmcnEIZN+I1rNY7X5an2N18ttz0isLoJfw7li4cPs7bZwo
eat5CzmqQXJuvM0UuSVRDC304mk9xRdDIk0SFN7yfW7gyuyfMEUfQnV8cG6lUItF
hkjH3M83dA6AI6e8HgnmPTfjhqhJg1wHJI6HLUBzLkp06LLWeSwj5GSr9fcyLkIU
QzvNilD1ROrqkBDyVbqjJKL8R0AmcpST1mkCPvZtM8aAu6YCDeEQfk6MIC/n8VWz
i0hf6D6FFpCSPEdx8384jz/7y/DQ4YlZawbLz1NIKsNbMQdZpFP8L8taplwTGwag
oyJSa6qzVovvr56Qy3Rt7rr2O8GY6/DJ9sIQXm65WdoemlGG46LefBu02ZpXK7pP
xiQYmjVwTd62a9D2o64+LuRkoqAzzHBmMWya72jKSpGkSyibV4aS3n2FoJmctmBv
mj2rGWRGAq50FAQJUYtQD+huU2LJYq0bjtN6u+T+MjHtgtfgg90Gz8I9IJk7gynR
RHrXiwtE87hQIBUbSZC6j8EsTwZOz2gdMka8PsAY5qBjhaMRCbFF/+L0YIY/17w1
NjUky2z/BWM+XPXeZkyK3qHzM0HEdhtkxhvhht8y+rzBbzdiWI/ewvu/liyeMPJz
4jzBUseQUfpqIDJKCox3GBjAIWqRulKPlYSl7x6qc4V7i7BVSSCWWVK+L8B3jlam
53GYxQQZYXLtVoaXHoZMrsU/BTjhidEIUrH2gLCpdP+Pw6okWFcuHprqO/rVAjzC
KBAWsVuvcCA3nNvMrFgt55kop/ujZfq7mj+FjTPI/WolCOFa+1j7QPGWv1zdRDvs
82qAptGL+s4MrQvwx5k9zBXcm+cUFV+BTJiHY0hNTihfqsHmD5UtkViBJ2lMjK9F
Xh1dP2qUDHd01Gfv8cGJfPyeqCDEui9Jk/3ssA6JQnbmtJjIhY7m4oA4zBs7b/KK
qThjCiVyJ43l9wDLsGtqpJ5VSv9Lf5IwazDnSRFBjTds8GPmOFSoYF+QdL2yehpi
cHNooatI0EnX4ZxKppToaRw/PhLbfU5rxmJUkfCeojfsuHKCkflecbWCJWSoKk3p
0O5HDhUb7Z7XMoTUQOAtJ6zoXOrcWvDB5wLpvLyt/JQyZx9w9FgyRE3dzyg2PG6r
/E3raYEy8YTHak1I3H2dv3K1WzxQCPidXVn4Ip+SyId9hI2FI/ekcq9Jn9lEXMRn
VdJu7RoKkxHs74++2NiDHuS6QMdmI9rTkVjHGrp1OqE8EL6bWuYN0dWW/CwEXpwf
u+hZ27b1kQJ/LBcSayPRKf3SlqBI2ZTrVb1qPJe2NW7jDJ5YCQECs6MypnFGD7ur
uwXq7GiUYi3hngK+ed4yAR7JTJ413VedxARBqZ+aqR0ea4lLz3HyBEyUDvHGtq3b
sP1cyV30as5mFEK5OahPnFCQvK673rvwH91wxeyjrj2ETclWbDd/e8c66bTpTX3w
lG3tusy9AT/dnSJJV+EYLMMUbuidgDUgK2aolR5oYq9mK+VpMHYp7WNRLe0Q+WSU
h7Z6XTc0dWw/2LguHxzfGhWdbzlZ9pRHf44lWxbmvCkRMebBo/ym+rCqTIgdDbI/
/msuOG+Civ7x+hzoCaHWugSPfmi9+kW3zUv5jDjGntnUVMgNSzwHyrLaJLFoo09s
rQ32RVsD/cnfSrfJZAHL1c06J/N6rmZCnGN5vPou46IMTBTaQrH8BSwmRM4YMIeh
5DDZTAd55QXjXTtdsxmRFHiE262aE85V2VKPRETMUyiDMMBomugdh9FDmNNvp9PF
K13Vb6oouclos61tGfm6AIhhH46Meij8+iWyJsmHdrTZ6VXjbbecxZi0+ZX10BfJ
gwQQJfitv96UvI2aW+hIPEWuofIoakiriWiJ9bqX1XdLopD9RXt/oBo9skxVIXdG
Noy16aN7zu8MTJz/VgR2qlM37/M0t68m0jbDnEEkk9O6Q2pB6oc9gEG/xc5Z/cUN
/NH36eREMKrP40yDT0HzBcfWcpjSbKwmh+IUbKUaPJzDF3fJcvDvlwAzbY/mp/BE
hXKAlpY4GSXR+8Ejidokj96alE4C1ZVhpIvoH17PAJsf8P3TR9yA9Rph6wiGyqWy
KepK4GZJ6poiDgfj2r4oqmmbqfQWucCSWmhQ6mvAQkKghj90PIK/hSyo+NjWi296
GqHHobJGKn3kb4zMStDwkG1+W85VUGzS9D/4UIwEMg8RWo6Trg91h7cUfItOcL78
vjHLfb8phkp+xYjgL47OVCI1+vnIau97y/sAz6WcZV8DR4Pv7Mz1XFzYGficU9D6
SBkfPnPkYm3btK+ZoBjcY2cUisU/veJjbBErWBVxadKXyuUPhBPUGNnBnMgGO1XZ
3bB/XUlNcUJXRb2RtVjpM5JbwQ0sv8HhmfcfIUPd7nENWk67MoKwUWdWKuk2NDTb
UlC3niIYrUhksf8Aj4Ov6AAh/wAMCOdlm5w1HSc4rxMxu092K/zmU8OgvEbPh7sR
CBkZ+Frqd0YX01ArrZiwlj3NduGiVpYKTL3qd5gHiWpClmQF8wUEbeSywHGn90Il
Gu7wficwIzgd/iRJr55olvfcihLcVQI6a/HWjw07MqUwX0ygs8y7kZEb3TANCSIg
Z1s/i7nkFYibbm+kFnjBS+9Fazzdz0htYJLYYwP+2C/16wqbQykSQB4lXWWek7M1
GK0XmpX5prBPPSOx7GbqptGIWiZyd1bEIfm5nG/Hj9o1vPLmOH90l+E1tmzeSIEM
aSWjlGRDDMzkvgCxF6PoZE4DSLLLyFaiTExd5f2W7NR2qOQ87GJJ0/eUSXOcjqYn
bsTLRpQ3/sbxhCSdMURFYVmhTFTa80YOZJzeC7PKO+FlhEkh7HiB5TuI6xUyYL9r
wcWXeJjJ4+M7FYF9r6Q6eZlrJNlPXacoCW9U1ro0NriwiHUlqxlwkSsNRZ40hbLh
QX8DVOwoOqMFfCm7w5i14jKiV2NXQNGGOG3T12lAg+0XZsvDW59PKcPMHI6qg+1d
QQ0MIC408nkqyAH1XswuF1dHLUqCb9yLvhaKgJXp26prym4JN37F+gM+VlJTTSR/
DJ9HfdY5wga7uEU0KrqrzCM+rBhxjNfq/zTUy1HY0xb6scsXCjIOGBr+7DGZy/8U
dsmrnMVZe3OcsmYjLetDaIZDn+KdfE1vBNzDdwdM0kMhDHTjA6Vd/wwX/PfVz47U
OmWER/JYXEgoGlyeCdj+VQPOGvom8j1Mp4hltEDtWULVpaKvff9UeyQShbNhQY/K
1JgvDW1hwBvZY6b7QcAdfe4N/Us61dKQRf+6t4tfq7ZC1Q+a90mMwyDPDY4ihHkE
kCbvo+RVhWgrwFcY9gFS1O1Ev4megp9GKOyQ2/2zx27ClKH1AS0cOINSGgP5iv5d
CqE3XQ7BPuX1hPcecp44O4WX15b7BXMON22CN8j6J81DR9pZ+U0aatevUtoC/494
2DvUHf98YYr8tmYsuhZpLby0hsGAc7z5l1GBVFpqkAX1HNmXhBwUpiaZoPTVac7D
jHbBFZN4ioF7Px6rvXWpbJZR+eo+/DjsSPz2AhiLaUFiU21plXmZRUq6wSFwf4oK
pOtyLQn389o7vja4YuKPQnDYvvVLmb0/3DxjfFfERZTdWGripzZg6QJsSWCYz+Zg
5yxQAbtO8n7d74oSjPMgosFO2Rnq8Oy+EYwfUZ4qnifXfKeOrz4d2ENr19qz26bB
kriNT+5bULAnQvUwoGLBBBKvX3sD35rQfL3ge0+79Mw5suSEwSSjcDmyQsiOTukw
gcW8oO+01G5/NDPLEI+ixgZ4n5+TuaWx7RqDuq/kOXzwq8fKyrzjgJNlgkiBLKOA
+HobEVwkF19weM3pMG5SQ2XFzQqXz+VLjg2AWHVicd5EbCZ0KKzfGxLs5zAkN7TJ
/E+fX2UasOaNUVuzjVFQvQuc3WbkODywgs0pUkTngJNzdOQ8PC2/xA+10qslhFop
RulJO39eVz6JJO4lynfwrwO+kuyUckUv+33vH+ihM6cDWDPA10gHINs0x476igzU
CTwaAUJQVFDmvJfGsj5MlYEtxssVD9FIP9mCOSzCvORSsJhiLTxEr/OnedzSwa7D
ocRxfwG1J6BGg7UwAaicwuBo+d6MtWbU+Ary76ad+NFsP31Gmz3XyrFmo0lGMyEq
U1rHwE/P8gLzoFKt3l60chW3jcfGRx+vTMKooh//aPNsUmapXBsBkEm0mexT9+qL
ZZ9jXj7eEHYJznNIPSDUkmk+dF9FtAih39s5G+1GEt8efqAAfIr/bvBtDpnnAt2X
sw5yNeA23DLjNWeTWSRZVrEstZ8eqH7Rcas9KjZYJ/V1FLyiiWjgW2bDUYFRNutK
TMVMVhQdgsC32KK15PKKbe9V9nC8JTvwcSpS2rq4l1YgcmdzBN9PNNG56vqOb+82
xRp9tlkWWNOniEA0SlBCeps1ZHq3myqhUdvYSI8SMEXHWJ+le5lYOoZadSRdT8Cf
5cD9Mf/Xe8cHE+Q2NMQFfAKrRsOl3K1wyw0dxKeti8v/ohbXVeJdfdrHkJ7wfoa7
ZDlsNmdylhtBJG2ANPucqHWZTcM+3bfmvhRLhSzjQnIV/dhb6V0hlIF7hY3icpuc
/CSgkrG+rhQgpV/aLS92OfSrZd4kUv5h/Kw/8rRec8Gw9bF+CQU0p/ZzVkECad3b
MSIpY4B8/fXoKcHcCOFCgxEKrBxOz8oiAaigbndFlSw6ghPAIQwz1wodaROgEVEz
c7C6fMhDTY0X7HveHwDkZDypUwZ+YQlhWdOcdaLPIihO7lezK+cjr8K6nO2zJKPl
SLpTlQt05KkOgK/I/Yey+WrgLPlbVtb/MEPJ1FuBQR6IDi1uGePXWFbqyWJwRoei
niA63bmtI+Xxz+MUUhPZXEXASyRhNl7KsiPiBheWorCRFe/NAjMVDKJHgoVC68dl
yD9o+JzIYAnSLPuXZO++rbWBsuIGU2p8v5vXs1Q6ZT4rtWcMRTOv8AP0HmNpF2Cb
8KuKwb86FwGiTCC92bO0PZjEWL2HBPZU77j01qQP0X0F7mXg9gO2elMqwO2UnZ+k
mUw+/AaaEmQucrwVhl+Xv1YY0Aw+zJotXPKfu6/g+mlsdkKv6aByVTBFbFRtvZeu
BnYuqqqv23WZki7rsVezgP1/q0F5iYss23LqATbq4s6gdOx8VMD/JnEfeImPkUt5
+kzVk4gb61xFVPEUUFWD5XV81gjaRTatieEgAp5eRPbzzAlgSotBMkIw8io5b9Il
MQ0J7wuuO58nwDUiAKoofrKNuAla8KUgncpU1iUze+95nPKj2UIOWnFx7l5KjFxk
U/NeWqXE8wPnOdw0UDDcUQHN27k+T6kcPt1jFPJSk8G2/92v2OxUfWpHOaPVotaP
OZT04r4Cs7lo4JEkEz+7nF9+qdoxyv1xrvvaL4mjCq+iTb2hYtzlu3PFppOxM9si
Sei98H0l+wl7gkaCNTAG6/0rTpmn0e+eKZUSeQpqWwV9ZnlQURxDVx+RYh+mq4sF
vZpZbAuUsMOJFDaUfeJ423qPkNYPVZL7MAVP+LRapYVIA2OjwSbBCJpoWWe0uJxf
XF1Xweagwm38FJWXix+H0Uu+6X5WJQQrbIljMh3e8ScY2lkgz+hOmElih1awVBtN
LwXvd4tF/RLonvKf2AibxfVtojCKQNMu3pD8SIjstLx3Z7aXl5EimlAmwooFj4ow
KLc2ImGz8ZnAj5NwuEtHlFcb/hHzIfBJDpyjiWoLZZUjvdunPErtkxKGL4kFEYjF
h9GrRB+qp92CiPysMxDahutepAkRKwyyuUBU2FxhgF8NxWH/xEagm7i19C0PG79r
7cRXWiH3BgKviYQjt2OaleNX868155fX6EUJRgHrGimiQaRnLmhkJbxDKmxWMHzk
2t4ALIxGNElPcXMVmLpxpEpGGYWeybz8KeaASxuKcOclA12i2Z1fB32mZRGNXvyC
FUyMKYYHHGJYag8WXXSCYzjDKZlfI5cQeZJYbs0v57fZsulC874+MTSQZ/2HhhlY
L2OlXuPAeJhJ/84Ow0Dxwy/LNEBFmPjNKZ5GFIZqZu+3aHAync2sMVPNK8kLvQtw
OiK9HgEZPYUgTmEgFfMsYjok/d/D/b8c/hxQ1YxGO9ItPqattV45YZmjvjZ9Ougw
CjwAIgs0wO2oytHSXNHfG5OliObnuyT2KO9tN0fKFR37JG49M6BlZu9eCIfnw8rJ
NpQLNS2/p/KXq9KRUWFgrGWTFlRkSmx9XRDJuR+hQfty1kV185/zYKJnbglahhSl
1HmB6Ovzu4NqcO4R1kWnspWFxYkZFUMvPqmWJxatlsZ1ZBCq8//qgDclprRYa9tM
AZQ3ZUSN8oxqSmLv1V+GBClAiY4B2EKzvcX94bb1mNt0M8Rl3Aeg83+dzzZsJr5E
PcWCUMfjmSOdQIYyFwlwsRoW4sBzB4WcCjU8Yebh1ynwhyS4dJwFYvT6+O+YjLLQ
kQdztmXz0rpf1pX0NZEvoB/a4YF9imRCVeoJNkiQTi/uCRPKpPnsh3VMHCpMN6Nw
rbpDMsETRUjZOTamwL+mNV8Axvm2RRKJx4MgNlmZ61g5Hj11/EpyAxYxCZ+U0XE6
B53UQPiUlMyK6Rsm+TorZm930eld/4af/IJFF8JJdOMpRg7Jdk91P1Kywpi4+/rU
7JdliQnRtoUk1TgopsB0aNMRuyHJs4K1njq+SzoeRYLR/reAckwTlSZTqoi/G6kS
+k7JHg+orYJDG7LpKMEX2L/Z4uJFy8ew/OWcjSm5aSalHP9X92lQ1ZJVLeBZC5fy
XNbgh38vt+yKjqSqxnwp2+dk+jT0tbPb++uBFZitsPPqwVIkca2Vb6hJqE2WI3Hn
MDVXdQ7xlDipKrJi45otUL/YGhN57TxhNmMXWTp7ZCP+X+TMfiaYLz0z17sK/1ho
bbxoWInxjlvpzG7UkeIM6+Vlwro+spCQ/0oXrf5Bmpya0sJBs4xO80+q2IYNAn6u
sVp/rzFG8vfaEPc/e248fGp1Tfy+vAKwrQagNB6hY/raKIUe4RSY726D0cccJqya
fRzEdKt8ndHrknS06isxe3Inup3M8S/jBQ6bT5YDTtI6b6PpTQOaLH+HRCBCwvWu
lqpCsWcLlsM8IbdpGFu85CGJbM09kecqItYY4WuMypqoxSUdrBtwjSsh/fRTor/S
UAPI8AUM0js8Z7m5zshnz3KgOX8Wm3gFTUgmO+UQ+TdJoV4YSNXhflSjhAa0Q9RZ
cp8uHHKUlZVIwe22KehfaT7O/fiYx8fwdWVrzkoYesPuNQ0E2si9vegxNUBd9baK
K8+W/GG/zwNmay41YoazV/X2tDtJ+er0v8feRKoLcD8rQscXUNwbqoYaHNbjI4X3
4/NFdlCA1ujp04htZPjBX7xeChw12kg/64sWAYTLYjNrCPHZWAvK/Bty22/yrpKz
d661hPpUoCThLDwHRzX/qKadOLPZAzdQM9GGDU+RNRsUBUUXa3tGgntyXRjh0t26
hGLfNzCcOHa/i3XQNQMsg9QgAdCKQjKFYwvETY8dVyUHLy9DKlwjRfitGJ9Dga8X
axUDFYP4YCrhbJZ3eve7ABxRWSCx89pbzcVy2PReoRq7zn2hwXGeEyD5DZxnVLal
65RGGrEVgG2Q6nRHCB9j3dgMEyHKMAlbTxVk8VQQEP7rnly2MgzMD3rmvcVby8Gl
CHOAsS5Md4P3DqCwrpF6ELpsYMc6MT4HsYmoCsC5AwlF9lGf/HmZiFk+89x0Wohg
h8uqDBlk1XDiHEYophKeKUhBJRqEMZMdM6ffMd5P5SBEjrNR80zGC6JzLecubTU6
DTHoxBdyUI8h3BEsQBnRJCz3ycg/Et832E5edvunhSq3IfsV/TRejG4thgNHaJmN
HskYa3UfjMDmwW3Zv3UXIR0cA3LB5lwNwzSk7zj8rFIrHFe16gj5MHkAa/pBkguI
jxx7U6SemRxbjhxkrU7ktn0hAlvSeANrKQy5Bx6SdyfqjUReID2SiaMOBtAiDxiW
kbdfcEGIDAp8Z4RF+m3A8gUIdl6b3wRmh8tqTHgBbaxEqeO1DkSaiUweVfNV9wwy
sMLWxMCwTeRE/PH9WLdTvwayF7jP+7ytYJtiWPAjVbI3lhWAw5Q5KySvk5hFg4py
fvtnFq6lquVvvPDdgs+Xce3BatJVirJZgFRQe6e/L3s/Mf+bepsGtdVBT+Mc2Hv0
PS2pEVDFUonhl7/q2nfDbO5XOblpQ7XlQUF0SHOjrgGG1aN5gtOQmHSYH9O05WbE
qaOdwXOaXin52OdIzdUEMHQbAyjCyoXa8qVm69+VsjC13Ow4nMAtwRmpVAScN9QC
A1I+A9vyMyWiwochG/OkUUg/grsYibN1uJW2iJNDYDF66zBGTM85vFWkN5hlQ2zd
GdfduURD3cynb5Jir2TXkmF/3fphQaVynQQGvggvVOsxhVDrwawyBB8IouAMknvZ
+S8yeKwK4lwWA3WZbUOBNKAxRa+A+0iZRsPv7s9HibkH3rcerSxu7GWvpvGz6y/Q
U7/b6GXpVrITUFPtvaQ+9G2hA+9RkvqEQFQe1n89WksJm534eKmmBZHphmPXJaIn
kc2WOZBBGo5s24oMh3xCKxriYIUGoEGl/QTaj0fcd96pOXvWvuKXF0g1DZ9T8fT5
qHd+XzvwaSOLO/XX20MPCxEBOb1/zYGelKJTsazeRHed//ilstL9jYYeqoLMjpZe
DCFyQF2Eas74aWpfGoXvjtrjDaqW4AhW4sQhMXNStXsCZ9OlIhOTt7+sunc9RnYt
3OCpRr+bWJTWwJAMw63WqSgHLWboBCywBbBRAigqZpfuQUUCvvQfONoINPIbGryw
R7qPgX8craf2IwtRZwCSXnw7b8AbYRgIebkcWhwGPUGFlsF/G0aj9xvklP4+dhnX
+HKvzaoOYWvMMHWZCWkq4/WbltBxDrH+/itypeV3yh7IdJ0KhQvuSNmUoZzhu639
80j05uBU1pyhVvJXsP+Rmn7d+Rdm1c48fk1vIe3iRsZTVAnihh0ZhA7r6q+vS9/F
tCZIthzkAjapkbItr3Bz+JSokT0NDFOQ8Zhx+tmD78cTorTB70ssi0u360xq2gqI
/EVKLUKDhuvqSGFEfWIIodad9kQeXDYDQoUsVL7wsJ543IHz2sn0YuCwFldrIr1G
UEji2FI71oFFHpoWU50Z2UmYHpa22+YuQAjm05ujESnND8+FwCr4ZtB5IKp0m7we
KMKZ87m33exd6durgjvqkvBIggg60ZRAtzhVWh8ut20DGM1iC6MwZiRJmdQ/YeUc
yIy+nhPc24zdJVnjQ9WOpLtGZHYYUFAUpaIbfmjgKuril9XQ5vfDytu/LYXUPIG2
rx9YY+oQcGHVQAQGqP8t8iV/5veh9gjEQaqdH2L6WnMl5UJ0FHfPbTArCFqOq8kR
GD8Cq/85uFTXQS+o2AKrSEADpNfch5simPXd7puuk+cc9NuOpxgcWdelIuCHGCfT
piDWK0/b5OwKmoCVS+WpvKiZQ4V6HMLVzrREulJyu5aN5jA9XRSysd1bT9B/gagW
dxvGh/DtNNByA9CywZ4ZYGy4IU62H5NDxt2IEFOvZQ9qNP0QISZI75ka0v7/v+Xy
DUbVt1ljVJBtXf6CiGXSsxIyvqQzgFZCXQAn+pwyHJ+0Bv0LNvpJPxOxUdfbzC/x
YKfmByEIE7o735BaqOfTGvgeB6aOfqV3jpVBZHpMpKD0PMfKXoHRhrIzVLHPTb9k
gmzGh2MAbWfQ2ZFby4NWjnlYKTHXD6cpnHvUBjAoP06wvahHF4Ld9UOQrZx4eC5F
9w0ZBo1q5ib2RnjL7lJY/Fh7NQZky4ToN7EjpYqgsd9hfRpVsSjZwuzI7C4HSb+e
OvixEAWT5LygYuIlANYngNcAEKkwi+GzPHEqDfruzFGYk9ykVaFGowf0wmbJ2lvM
MurqVtR487P6aR7He82wVDsvy2gXvcD4Q69nRsppoE87tCsk/CXgq6/BLrneNw/b
ci+LIbdnjBVvyUPK0gbiLnqNt1HqRcdk1AVQt9hBN9R+6mVMhTbyPkh4nz2az5P/
BJGbmN6ii3Q69lb7ICQw7laIysWiu6wGDOWkB6dq8/VDItlEwHamPkRd6jzqBdkk
V2RSp7MgPiFGRjIlLWaUSbAl8gKPHfp9LtJ0vu8z2pyq7WLeyFAp/MlqMfrvNaIL
IGnfN/tx1aqr1+KJjwGR65RHPKFvpi9d6bd8BI8wUcm0XoRAPmCHQ5T6wFeuDl+O
WZ7oSWCQNJa2olStihY4mjmnDSz6fR76RtOHt29AyRme1SQnH+EgLoDcLWVFWTip
jIQ31rWZUwE5fjGZpX/SMOWrLZ1bcDt5nMLcfiffHwk6GRMP5Eng/HpU+XWQhnnm
uu9Q94O+q4FAwjoRFPunyzEG4SS6ccM055MRpbftRKepBuQemeX4ta+SkZpTBhPH
5aUfN1hwZYUDprSqFsUzAZHqkFYnb1htc3NCVtvIsSMatvkETfcqR2Ma3IcvrSnt
JkkO9tCZXbkX76tC59wjDteFykarGY/VGFKKFi8uTcjr/iHmDIqEvtBaVtf/u8yv
ylgAqg7JymCFMFbd7ac4pR91vAvMdAlyKzj6i3zz0wmv1kD/Z28IquRqV/uZ3B2Y
uVhkesCSIUivfRZY3TVQ878gh7W29Gd394ucRqmvU9/MJOM8ekUr9qYZbvlPEMQa
7ZwR8fPoZHQuhl9jjwYjxmq4yIMKirCZ7VTsbuQqiKXicxQfqSB/34IzQDjxv6f1
WPcGd4OwlOCNk1Cof8+OzltuCcr1IFer04zpuBsqG1Pe8N7E3WPv7XD4IUxeZ8Tc
p4UD+2P4tlKOdTI3liNukhBn9Ef8EZ8jZiAAdu0Eof3kfQa2voL334V9fsk8gRNn
kKVwdCOjOmJXBITbnGyMbPgJ0j3DAJ4yxleR7qgWHKD910N0jjds2C1g0G1VJyeQ
Zi4FSQOHuUx35jUwZ+Z/rHkSYdRS3wePplfgbPJa/WNCpsRVInGCiKfYcKDWIqBE
PhYgBtMOXqf+rGKcnOmwPrm8tnhbh8fpf/jWfUMfsv0tIUvPDwTcWyEZB6OS9ej0
PxcX2nk/0cKap9wPlmR3e8XVWTL90NuGEDuqDqocs7OUWN3qoTl/R8xwEJIIuLS9
Gys3ObLliWztExDhzdrb5YYWp3RXOn00BrK2fTCC4v2Md4TnEFt2iGmnBMfTI7YU
JXUHMDLLVaOCba6EFHH6FZiEMG2gXTX1yxvzDMJ3rx62n+V9iOqGaQ6gUNyaCALG
qHmrjpWnJRcWuxJKf/3B/IvYS+BHxova5lx/nyVoP72lQE8J+4FIJJjEWY0GwTLX
iREdfqzK+IJ4pt/iapVvC1utuUs8nMH78Cmf4H8HKL3hC6BmmCdAY/uLfQI89oaP
mGRURdCjN5RC3LWwG7UpXtuESCLbmxQMuYGZBQLrC4lYWBIHgcNgbfjEYYNpmqrh
gc9CJSwtmhWhuE2bX76nlYBR2hYp1gZe94TP3ASXwADrT38KQnjI2mWEOOggRyWX
mXJCMXnehlAhFZa1LVzlXD3gfztlSXDSThVXHYt/SH+7jb2p6c1E/t9egkRsLDfW
vMNjn/Yn8KK773SAbwgndM7E1iyrXpHwWH8vy4EaK6VKo2QQRv3fpMrbMIMiMNKt
viCYi1Iv+myjLQx2KYnvXHGsUOooBsd8Os83N7+crFJ5PcLgTa9JelfCySwwGgx+
PRRKlkIltF4nVHaiZeLz5lW/Mw7FtSjnnbMhwVILRKEUgCrSvcHfhrcQ17dZhKhQ
mg+gJ/pqEPT8hytO2AfPzPmLUspC+UyRxnTGzmRnCV2C3qsYxEzmxAMbc2DnCHki
0ZV/ZMbPS0l60yiwLGtErqXbz2elQT/vAmq/e70zLPalIr5GXKVsA3qd5xGA5P3w
BcrxdINjDX+BG0CM892HsFAhoEVCCdukouJKAWNzBgbzR7HB2i/yoIYwFDNkYGUP
VUgSVgbz99VJ8bGx27AgeFDD7k4Hh6VcvQ6jhtOR9aqv/shLkrBMy7u1mAO4+4bS
+5uGwPTm+leGrnQNpzZ8q4lbvFPyx18SgVuHLbavOcF8TnWmQkLhxosFO4EZ5rOs
J8zkijNxt4kj6TMjpqS53n8MpHtF1ySPCATPHRk/KeHg6ha/tQBdiwsvNUndVO7k
xCXnx1SBWXkBpboP9z77HSCdGlrDcrwiLpOSsBSRJFK8toloJGQFA4YjgFtArAY1
oX2LzrrGdyWmpIYsf/fLxrZM07/7Gcw7T+Dee3fLUzYgEPWBzzNAJP1OpOyBG8Vk
LI+AkEE1g0c3XMGXPkZ2I47WBnN8VENMBMmTZ48SlT7EZkulKWzHvhe2QG8FjnB9
fnTAOO20tyG+9RtCxrUjlRYuR/CWwiOMZB5St5XosaAbQw7N3bqrHSlocwqYE+q+
JiBIEDYpHvTlYlzE3+CXWlKREXNtLZuTU/fKD1dEmAFVRyYrlEwMCmn52y3Oo+vo
PnZwsjT1TROkMWOlPnoLOjJlSa3TtovLGGO6f0guSyAMLS0xepcyTI2TRKANdQC1
dI3Koa+NgDLYyKN4OzCoshSe4jtX8CZP9kgIpvutm3Oc/ldhGOguAjgPpU/HqrYP
k0+q/Uw4oj0x411+rKZxcHfHa+xo/jk5iZJ9beeUWovHzVu1ZfrDCXa3E8FltBdG
b5KGv/jAdfCXpGpaXiJY86sNAne15rY21L2/6NxPxK3jKzp4SdubrZPYDAFlf2ef
iogqMh7JZawWeibfyiRJZouLhppKFyNXNILwaIQOoiAUcBgxL7l718Nxzwyvq5GK
NpnZ4jqoaEkzfVDsmcitUQjtMNt8GavQP9b1CSXyTmwxZIynxRZBceJT1gLc2WSb
mlj+oN3iGSzMG45kuVrA/R8k1ZdcnV6OxPxIrKxBnnPiteSuuE4XXmWh9/firQDX
A5dFPXh6wjuf+i1/kDZ7wV0eZXAYnMn7vs3wvlQlfrfi2qQWZP3j/xkE5g7oz9/1
pPcLVZVplHQsujk63zR+fGScySFmlwubrJsiaMrdBo0+s0osvWa3I5TxmK0OYocw
wydT3Ud3OBGMWvEEJzWYCqTzNFimHcViYkn6Lr/KmVOVUsHJymSKNv5ps0q9yUic
cASCVyUDvlpvY3HvtnBTModV/vwcEzuQhaQ7O+C5i6DysZXpqL8i2EK9NFwWJwoK
iDgJIG2C0c4fxjbp3OLip1PSqWgMzFJkg4Uz+ceWBT5OY/HFzwWEDVckwWjkLUhR
O69LcjpFyfuJB55SuabVsNjSxASvS+JeVPCiCuw1kZf7YZZnhiG6cEHRFXsUIq1E
J5pxDL2yas85zJhzWwBwRf5uIqF/AXbK6zPW235E9sniLzLmAbA70UpOFgGouQsw
n/YITRY9e1q1y15KQ6/LtGBlIbVIA2q90XpcfUG91Wap/4zgYtJxSzHstJNxEyfY
DK4D6DKrRafzEDQmLD0WC937a7We7fWwr0uYbpx5UyQdfQ5/9uggeNigaGuHj5EO
u/WEemsMNveE+qVwK/TQYeApeOcdwWE06qEec8qy1MVt0RpS5PSIeKtDgGASno3i
nCW+GgieoO9rq/8PcR7GZmCn+6KD6fCUxCa7jcAhJcjLVOQCBSltRqBv5Nho/iF4
syAS1XZ6nvckMpMKzuxIRlLHd21DmVcw3xFzXWsJYJyDks7IH7/34nAsuQ6ynqoe
klnMQKRdMr8EPlkJ3QtCcUJN1hLjCCJYQJRNnLleLtNMaMA1o2GahdO2gB2yf0wi
Fe3kKkV8ah0EQOGlNuC6GsvNmRTD3SasnfDVm1YPjKrmjpRCJkiYzDhbvkxEfG7l
0xAjsfrBpojGM7rLYSuKcZ3zyQ7Blzm1fhY+SwoBCJRrUZuXsgatWVMNw0UR3l2k
Ei3nUcjOoPbCneTetAPGJ5tLfPaiO+5OSO9wfE1cX5vanwA5fsLV1NWUjjrxuG6y
jngGsrzwHehRPUewwBb+Oe4FEDqnkw0FiSxZA5Xf4H1EXqfR3N82jDGnEmhHAsez
JHROhr7jSKCJseBSpNJ+2rexBFm1huGwxp+utA0aNgGzDljzYKjS/OrWx6Jp6HfC
AuKHT0UFukwxGy1GwY6AO9/rtdlW4VrwvnHDgGoiYF7WEf2Z8Z6i/ICUTXT5K+gq
Oso5ivkpWFup5tM91QcXJ+UYrjVmI/oMLHpIBRwKaCCv8YHmVdG9gpxcuhJxjMax
T2SiF3IDioGHIkT51I1fDmzAzoBvR5puJ5L9JPCH2CSXn9db8yiTjUVXglsqYJuC
0VtrAK278vq4DxiG8fyobDTD4sOYrLZiEDjWNsKXSi8tcfp++w6CJeWuOq7oR0B3
N3QBIRD9A/QHgqAMdBGYG19XQrIyyQdSdDHtRJAGSapK+r+RdjzoiWSaDL6gFmP3
iwf3giSF0RlseSjnc3U/zSoq4OWBk1z+OLwdWemSr7QHL1HTI+1G8th56fRbuV7W
MUdoj7Sx59ysJ7uy0am17v+WarXBQjwamMWw9qAkuTt24lY1pU3NLr0P5umYTQDR
rZdum1RpwLTawBSuE1AyZzdUexvGoTQHYE4+9roAwgMhBsfbBnEvoqRP1rg06jpk
62NTQVaMqocO8vWEfuBpwa967Yk/zanA+5AATSrlPYwASrae00jKKnbmymLcRhFm
bQ56jgiqh9BYkp/+ZbMD7NJW2WEbGph0N7WprmX3+PY1tJYz2dFucLVM7Yweh9Bn
00fTcHhCVFo1JmXorwxpGqOSfpENHZaiAmU7bERrY8te8nK/bAnXBn8iiUN52xqq
0GU9z0Xs/5MhJUg1HuWvTTF9ErhCb3C/LhtIZVsZ2oax7mF0stJY3iPmzV1EiC+B
Uk7uwNbHt/HY6pqhYy7Y8jMAmvqZAkznctHQbqTSyYXTQ0NTn1B3nhE6byGtfIPS
bdNsQs33AJqHUYltFo15JfDjAL+EaC/Y8LHU61ckAccDqYzXyD8UTXZCAWeK2Uyw
F4uykBD/k0NAVR0Jab5hAg/vzDC7Lm6LTbjPb7bimEPKYJacW0MLhS5XrNmUJJfv
bh+yuDwxuCid6kuEsO6mG4rz0MqCVDTpToHvhlG3HSSxutoeClrfJuNYcKoB2FjV
I+rmuHFLbsh8U11Cs6XKhg4sFvQ8DLVrl5vx6t2i8ZHTz7U03HeBlkfgaD7E+YJA
k0yT/6C190Lm/0ZVCEUQvHA3Q2APT4TEVToomxV/YLFfNba4oppHAIM8BC3uw/jF
it9Qo9vArWy7b0P4WYkTeoOisnEf1uVAco6paY9VUBERn+0Qhi/SEU2J5RkiM2CO
QTESv2vbJ9M2jyKguhEitK0+uCkmOz37suQ1+UHfrqlP7Tt3FW81YjBzH05+nl35
Mkm5izZ0mZQpus6z/6nhamtHQHdWliVUyatYnQ3kaFytxeSq2py4KJTg2ulerJxP
cbAqVo42Rqp4iaxwkUaVGm0V3FlHfIhvlZgA5jVK9kdz9g1f1jH6CCEv1j0ixayK
GqMdw24A0tzRrvyLHOSrOSbHy248B04lneVBmkvZ8UUdvvE7HEDkvcQFnchjxW/c
ZpmMwzbydK2L+er+r08g3xnkxYzPr3IXKK2bVTJjIJ+Su3e58TDazy8YThB/25RH
wEZE64eiUZDU06mkzCODE/LX4Kr+qbsVt7NbcgV0oC6TRQOqXip18hSVxioF85em
aXWpPLaKZ4FTkYwzX0mBBPbur/S3kEu98INgj9mXA4I3NNBtaUFRB0Il19VenbCE
DL/mCF39F+HtHl35zMpl196/hkTOm8lLFbsc11Q939uyseyEIui92N/I7pOxxWX2
rF60P21wvLRG0aD7quNZkWZ2WP1vCROEGtTGRage9YXLOa6sf+3u4DDbIB19EdT8
ZCcDOmw4fXIHjtdp83RA/5TIpCkZnA7ksHAO3EsAIi5grS9nZPLbptar6Vfaogyh
8pBBIIy51QdUB5AZyNWFrLOPyMRKlsrTw/KhrlRwO0zw+4ysCUKqiOacQkIphui9
97LEARa+Uan8f1Pk42K4AavRrAZpYy3/kTE/B8si6FvFM6a4a3DzIY3C6HbSk3AQ
fZ+iBA2qaIBMKhJltIHHuegp4ikCJsCmDGIJ9LjrY7M9+8pEr8BZhmADsCFTODbZ
tUQVKUaTP76famRBgBumZ0yTOMrTH9KIFWj2BposjN1RtNGCGySZi3JFbGgD0Zs6
d4kVUNlp1F5ScZS2fUKoRvGuToy9V/tz0zSfrd010n2FtTrUmQgDdqfv5qK+VzCF
wherCRUFQ1br5HtMbvvBdqxGCJnlUjKZk7P/zwu1kSvE2A1C5Lke/Pybp1LME/nN
iN59QuNUEaJQvhO3+lgcNP+zqZXe63VHC8txv9ynZEyt6VCscGqXPoLSzwIKL7B7
5L5SFZvAIY0npgHlHfazJx0lzcJWgpyOVJWIhjFLbX25QeioJ6J/8Pj0F8nlgPUQ
ro5oiPfBTpU0eaDlGHxLCubd302SoyNGhqksNmD9CVctHoc9LlRKE05e0ZN8v+3u
O7LzfGQ8poTEn2mxooNoVa7y1X8rQvNIsMvneYnuoKTm0CGfqPc8DLA+9+IYYVix
mjqx3MLg8wmKyT512lSV8XntDSF6hv066E8V+3lZqysiIIJJgt2C1mkQDypx+hV/
zkZgO/251N66j028TqsQxqjOf/BraAgM9Mo5oz+SxHMiINUuv/xxE7v26wxc9RsN
0c5QELWfuW09FRz5EuIqQjdzlOCRdTub9aBpCLC9paexbfxPlTc1lbkFde69bwl0
rjZTyU+oszmeEZL09W1e4JfyANju2MmCBV71VqoZOHAhux0LhEyZlhSoRx2uZ3yw
dQGdEJ1NWfI7QVl7aOGpHM/PdvTXGCvH4dnAz0j044KFVouGM6RObgDlnT/HJFiz
09z09GyAGpAavAXQKbUdnxw8+9ADSncokSvUNc44vtHGdxEsg06DOhXGLKIApEQr
dyDEr1uwedcCoIn9C3TZlK9h0/IJc99edrrp+1PrWWaH5KaR4TqDMYu3WtZ6JOrU
IkwOaiiOzCV4PHmtbljnMXAqi2D3/0v6v6O9KGOfRPwHMx6qIlwo2FgOdhfvFoGm
VWRpFFzlNsqFBgfIxOPK3/pc/ZLjV/lWWAYWfegACVoRjn2wzTnhB/o4KA8sz5cn
wBnz6Z0sbYiUiq+qOelzbQYCrG6SdlVQDfdIPCsG8a8mOLcjfwGWUm+INvrI483z
8Mgekv8XHN1fQeqvorgUDu7NQeh3S1ZVqbSBiCirOrneZwTN8S29IAxskD0uPcd3
lqk3Qyh0IXlY/oKO8V78kbpO4oxrOi5Upa0cXyXVJPNY3ipiM5BCu7e9VShYwsS+
n5qBayJfrdypsl4vg528pgDXnv8RSvbxEMysslU5u1qRX5XJdjaKGWK5er/hm3Vg
AtDtcarcJkGjs+N8dlh2AdUMIMn00d9cXptdmSOXminkVgGNFjlS2CZ/c099UXiX
nvI+PB2vjEsssGAXvlMbZxd4DF81YwCN3Z6Nw+kT8AVHAycIGRawQSJtKP1LerrK
KxB0PFDkm/ZZby0eMJZzU6wNnxNfNU5CZ4ih1OZbyajzKrxBylkKFPetR3SaDsl2
LgO5jXgHA3ibMBB77ExC4A8EaZuu7+xDFxYVNakky3Pip7MVXjAlLyAyjkEl0POH
sMcWquXA4SbsWAMHtJ8zuaghTaQ0NcqsZmlut/S0tohct/T70AXEYk969GoUcHdH
ZVu4wb0YeIaROOV9MxsrHwHDBosPU6FpnzQ+YUB6rEwB6aZ2ickTR6oraCZnOOFK
IeQYtb8qXhTXhJ2rNyRkaaAEG2KVlcVdS5smkb0AKIAnPNjnpmIPA4Lh/+gJbZSd
pSbAG/OKxrDdy4UzzRclEk8ueSiCvtsVcq8Tg+Fj/Fy89Vbdx3W2HwscutCrdl6W
4quPbqeoQ59iWqqK53mNnhor9afL0ZDAsIzVBXLsw/6r8aq3oBULkqxC64DnD9q+
+RpH5JGafKToAnUoGlxg8gFtT89fhlBFqk66vm7GZ+VQHd3K0B2wvnLRfEb3CxvU
SSxLzWAofd/QbLlSJg10KQkZlnvLM7xmVInH0U+n++2USvxrY7xBhwahz3wm6U6T
dqiXg4wL7g9Wx5n9lJDKMkBnKsys+bZ/IEUUEn8fmKuHrwWoYIHq/lm3YRoveBP0
55KwU+qYwQmWTTOdA9T3PvB4RFCqktFxfG8TIFWG1lG3hCJ8GCJ3bi/ZqljpmBCl
x38XorzfGAEwSb7Asmnr3lRSgCUXEHhdEa4jwS0OuzApzxnrT1Y3zGQiVcGaQ386
toPmw2L5fLQLH0n5vLV/KTRRua4ywd/kDDPAj7JoEZaC9VHyWMH0D4QDhYjlUXNI
dAlYz2IYW8GlZ0q2ITBxnofYs3PdQ+Y341UfZEzBWgHGi6P5nVzw5AkR4fNzjNPd
JzS79Pp6aUDaq/YODn1pAD2Q/7yUfbmIAk87DFemtxzu0T89F+yrZ9Olxu1hwL1S
clkhE9994PxwfrVZXfnjBxPlailQfITv/CBbIyeyB+M+xBLH/hw8JcTpRmoWda6f
Pg1wa9nXYOe7xxM1pr04uCEuy/f8jVqqQghPUfzrgC1cVKKRqmPSwqwQDU5U2CwA
lNx3lBa7vUsnNKOWjdTGh74NF/U1dvz6UawDtzy1k9Bsa5HulmGXLXaJogPCsooL
ZsEKSF7c0Voc+lB8l2x7YfECFQB93OwGamg08Pmbs5U+FbfwQ8GiET/UP4h/BV4p
MTjK6VEqOrZ8GT/bvJjhBMpo+gc2oLfm19zosVFRsFCpbCcZir3WcCmAJWc5rZHe
oTRzJKNbVvOo8kAoI+l6RLEHmBE9LYVGd6h0mwM0JpJEty9SY/HqeTkuE3+7vFJd
hcgx6C8L1PTjwE9/F5AuGzalHiL4+NXFfoNdx1usfSFldTJjAKetOclfgegWzXK5
D/nG4OE0FcxJCpGh0IYgq1C7rcgd62OsYpTdjOlo33TgYAX8iKb6jv0+yOlXAkAx
p+uyIyl3E35G/LiiehGhhNi7RIUrW2doxF+yRoDqRllpJGllRcbeqbreuAWxWRa7
C7FC1jqh9G0I8BsqXoZ0oAFzG2deBVvk5Ut0vzbnGC8jRhETjKIdssDIpPz+CP+j
PRFFyYfZKC7w+pJo+KgzmsbdyUbe/VLKNwtWHNE2vpTdB116jjKdh2q8Q8d5Iumz
iefEvQFv8sEqLb7Uj6Vcs2m8ew5RvqY6zfmWHKLTM5YIuDrLcsKDAhk/ylz5ebg6
xDbGqShKbU3m4vbMe6cq0KQPXkYMJVreEnOX2AtPsdOFPGXBwYcfVH33PWdqMMJL
T0mypVvrj+w8yHu8Y/Q8o2791DRxGbqUh8JlOjf4XJQc4ZasH3IrCfXR1Upjl1O/
hgLbnS0Tztfx3vE0x2AaihYevpoqrGjy2QghnOyb0yzRMT8+lvCrGv4FYsFvYme7
awWmbwLhF25Y3N0ct5PhewOhClglf+jZZ0KmBgpP31x+lMoCFRFpiNvMPO4dV5Iw
acMddNVbvimA3x49RBHeO8T943i2Sekk8NYXXh4Y44BOgQy2qNedlirYmjC7EuZs
phS9aOdOjWa/NKjfNoHeWu4GtuEjxiE7yH+RrcrBbm8TlxsIu7ZqPrFBv5fyniOo
/ENeXJifDGK+sGIO9MNynG00ekpJq5Mzwq8T+TaTqlly3FbtoSFt56DJXnshNxGB
7vZ/W6P+YAXbvJHMVQ2Rp4IzcKqx+M0cU7cxEupXpFXfT6VnBlw964Ag54q7E2Qg
MgiF/CSBvJhhvCSx8vR//isLzYa5F2g3IOdb0c6uOSgCK9Hi0fE/g49EuApYRih+
aXknmYkfK2GM0vS03aHNV4a2FQXYl7gDlSB9TSDLtOt9D7de4xfubGhSM//U/DTD
BXraNyD3q3RRs6t94m2cSJGUu9E59uZSJP3S/O3+Qq41wT+kcRG7IEO08jAEuW3y
hdEBQE8fa0WMcCUVU1hPZhaAapcpp4amwWaGMHpOs/5NVwpGMJNmdd9UcmpE6W8W
ZAqbAaMZogMJnUjMIh9C2cepfSarIJJhZIffrkpIkiFZ1mGOjyJV/b1bVvLQgymR
sm7eg2z/h1CSmbwIqk5zBW669rqtiKnH/PPw1BBsx3hkZV6HUgxdqA5oHu1R9r/v
fhZCuaDHSu1kN724/R5/sOlbDbpxR9gNewSg6GSg17v4xPjizDEfjXOwZymNlmz/
IgIHN/YxW9GDh/NroZAPxUsKZWxteDyI8iMXKGmsGdSW0pE2Sszyv+WIVBN/8xJU
4a1L4uDjJChwOvoUAZEmHWh+Tp5tj0FkzTcoe/SF7GkEr1GM0ZbuTgD/74kgSspC
i3xYR3Z4Sbci8TCBLMtUVNuFASFaYduLt3Mj6YHy58xQbUS8girmmhLEVYstVfoe
K2eRE/UsS9mnBXzfK53hOeas8lYIvBwvIH1cbBEU5lEByMe7muz4fXv76dL0483B
hvmcUPWlov4BtvTeP2EsaBSKPj8v6vaX/XSW0mjJATmkeoK5RTH73Ct1eNyBx05P
0tFr8tFPjJDoqLB2YItk4r6Za104+kkhPWWuI0WnfSXqA+O2ZELxzkF/Rgeac5sw
q0JRxwATCKEqncYweW3I6Sadco66oME3ypD0NGVXl7kIjKTOld8dlSTL1c/1p0+r
B+c2OHOW+8D/7sfsXQRzPZg8Z9UIcQTou9z+z8pVgb+pIxsP6LEJytq5wHFyvodR
gwetGRRWmsE39aUmLbnWhZ7IgCIp6eIzPFTQLo+NN+3i+Fy1E6rZpGOozJ2hmXVo
RmS9O4ll/JZZJuVfe33hnsOx2jSqgFKtdgDcsWROBBAN+ZWoSABwGGEI4kLf8uHK
PyCtB0WPK4Z7XjLDjRa33XiE8/v1aYRQL5Zgx6Ya486CbVEJJ/ChNyv3zzffJuwW
X1IGiw08ztEo6KMsCK8Q7iINP2eLzSbn4ecTIyJY8d2KDzRPf7oC0wXZq5A3hA9p
71QvMGtx7cHgE6IZrzD9gY8qaRQsy75FSH2YqA42KzgP8VhSxNIrQW2DtfVS7Q6J
gbvSX7MVKZvqv6glOJeCcB0BobR4LpkbGvvf+XKxkDVDjqQaezoixLqb137/v5dN
DJMZT15fdawt4FEUkm27r9L55tUMjrzTeqHqERoRnwLd8BNrgZaHR7SP9r6LJtP/
LUzC39lM8x2RRpfQVWBie0TBxE2l5WtqoeIEwL5iWuarrg1dpyGsM1/IhLYLVPsZ
6gG84TP33fTIh6mhcD1ZHJLU9lhPTQvqM8dv66VaB1ClwtTAGQCJhip8x5PVVBJg
PdbA7phbpflEaRE7mchrSVrwKvVqsXCnIUjJzZjOtlYamVS8PjBcmSLa6VjkDNuo
BJ1MJVezPhHoC4FAApu3jW3/GnPUIdSK4VTJZnudDK4wa75uPhl8jME6CDpORNox
29E/kCuIY7gnpEw/MrHlTxRkkn45PXp+wCg6MSVyuBGvccJ/6Ta8S/s9y8SzlqmW
xGEHyu+o0BTnjf2pwh9YUYMRBnyrG4tHUMzyyeLmzfXUcasgGXHclLt8yswm/b9/
OqH1ERbBNBIKQh5jCSr84VLzi7mUn8SirYQTfsWd04CvOqb+IU4zL88i1lpkVOIL
rKkFvYBk9u/IMwKXrJk790RStXdZx1//5nW9phKf2BZLUv6gsqn5nWxnoNIHB8oI
VZaEBf2tNG8B/Z2F9ykIbBjVQoTODQLnm2qmJ4EpdjcM+FUDkxd3ltEr7tZL9O1I
dooEn+S5rvEQ57J3ZA/p09p7TximMZYEyDjZeZWBTF/XysdjOPBHGLLrL7fGTB3Z
gzro3LGSB/sc+A/episL4NvL8Kw6LSt7cznovPne2Zg8urLlaU1cWHYjAhIoBdXM
Ys57w+c4JlWs6b7J0QqjPw7G3E5QH+32+5S/1y3bN/z57LWTws52rpCZdv6ROfYL
VQF26Ayodg72TLVygiHYw5mej2QmW8MpDFkhnKHrxEr8eZohsBr+OW5cErA4MzMA
mj4iXQR8QHrbCGq/wmQSXEbcL+c7edogCnG5JM0X6Te5OP9UwwCWDiogrT6/05fv
BSULpAuMmobKrNHTLW+TcGfOOUTPfNVWXpU7Q1QVTM+Ja6vdEtnHm4PemOuRhGgA
y4GsamwHvvyzG/aSb20dDWQfftVV+MenAR9r9G12PrmV541kDhxOnoVu8AwjPbJY
J9u31+yn1i3JLdCQqu8/BMlKE+V+Khz0Ua/xYcSjnO7E7diI0FJcLKWkDVUzfMtt
6LX62mrhsxSSdYkKH06yX6xG9IgUedySRrna41sg/OYyjZLbypWK361hq4MJoMkD
kC2fxob3r5GcGIv1aLCryA6EB0+c5Y0bqgqJALFWw1jZ2MQ5O1QtxBBUPf4eutDi
SzD0vxRtcVcUn+BKJ/vDBsTgN/7C4x1CW1iGTMybsJmD/b/x5RFpD4OfDlhQPCl1
Y4LeGdBghQQgA9RI7PmdVe3v/n/GXdiyIKoI8s4rBU2lr/dobOwG948/w9cEIF8B
Na8P1Lp5zTtxFbgNwJik3LgHAyF2Mp3jTqwRyZqZdn+YhugkokWIG+thx5pCG7ge
8wGldat6HsINCHLl6niBjjIJM/JNaEHnI/yVjrv2e9qqKj+jinOIWSLl59smStEq
f5Ol+xhh86oFBwKTdHSOFN/YN/I7MywOu7Qhv2xGHrm5cmVSWB5pyUR0vfgxCIa2
qsk6ODXt11k/F8VfjnwR4deQX2cTNpYVclaJU7yvm4rYpERG7xZSFirJllC4LrXU
0+ucf3BtNV/l1fgchALuEbauN12Gtnq1poNGaZnzdCDZr66XpdiKy4ADLYmtyktM
AI0FoRXmRzADjok6O7NUWpkMDOvJkwXbR6Q9v/lWXF1tQ7b/tSK1EfrRn/GO39vt
pwTBnFwHB1UD264HWyxfjz2LI81zuVxtWoxoQqIfHvONrSFeb3IwTciPIN1gLea3
PPhVZXGy4GDvsj+bbNlz9QWpsTeSPoQt5YaNMjAZkJKsOZvPdhsfsj+QF3VwKSg6
nyT9B/KVCkHOfDvlrG/dL8f7dpEJlJd45Zulx4ajDcnDYqp65uv5CK9rQbHhw7uQ
E4fXZhOaYyiFgFRn7KSxg1KoA6oad8vmlumZU5OnN+VdKGYgG6jpfEbJkKBQmDqj
9ZmyxQLra19lp/6VyI3e561X8QqtVRPNdw2EcO1HpYKt1ZZCEszETkTWY3kYEzA2
q7g0uvw4BrsCoHckm6hkMZ4Hlr6MiN+l+Pf3V7ulYDhknd4HHwyQu24hDotIXKwR
xWio7oKuexOAxli1D609WrlfxEGeBZO2rwFMkf6+PpfzsuA9ec060AHtEFFx/MnF
yQuaLCC6X6r3ht5xSAHNWuArzQ0SF2Ksm+8ZJ8w5FwNCBg/i/0Zx7e5I7TPWELqh
m20h0d6IDN0OoTHNpdG0W94fQJjyVhLbzquMvL7QD0RUrseubge09VkgS4Vfrt29
yk9pYTKZrrtO3vYpTME0MQ+MR//DBr+osiLA1m20b6HZN2SHlS9CXWx6CTbkPN6Y
fZrioBwHXQ3+GUBwYYYo7Uh5BQsNLuLNmqQzB/tnvmbwCQVndCTY8A/LejtUTirB
HIO5sHtdoKKjuPs1ySYNh6Ww5snY6jQAEFPMyNCgst/fyx8nYsLWM8De7AZeDfuX
3kbHgHJSl0jzc8hR/KNUWRp6zycPNqYePzhNi4DqhR5yMQf3n01oRq7JXwG/vz7D
6zV1mPYmtI4e6JcXEVL0JdRt/aSsB2NMshvLZJEWbhrzFGIstp7ABtESnlYe/oH6
JuXTyjmKY6MuoZnOJGAqrASqZL1H24Hy6EQ4/ksXKB0nvCt+eE7F/K6S7FtHPhk4
uXhdiAiRqKOwB7SAwlJy+dwAKzy4LP+Wpb+gslNUH2nDtTXgAKtyg6DzTm7XLKET
Yn4w7XzZouFCcUwre82fFQ7JZ0tSCLxvRiggktICrrtptCs/q7KMYDXNwHLT5E9i
Qm6X/iREgkIZ54vacE4ParsnaYc72rkLAYItjDbQRpl7s+piLhZfOJJtN68hhBW8
hI0cUVS0IMcCC73zF6bsxL0S8RXBDq9M7MxyE0nwI3RcfN8KzdPDncDA+Hk9HWLw
HiHrfw8GoI11WE22fIXo+DO0HY3JS2XpPZtng58oxqrvJsgnhcz+v6XM985Tk1BM
vDuZN8trz2UdY4JkeGN/DsHEjf1+HdVuzeywU+0S6DAer+dV/2DHFbfzLeWrccGR
u8aRWo+GvaqOiQ2QoszleLXqV2U6gN6PYSFl+ra4DqWhaGIN4OoRn0QigaOCespL
B538Fqpkl6iOgs/sCguPqeMn/YPlyIP6K9GibF0VJRbA3Br34JcBPHsLmlr2t/Yw
lkcNnL87MTEQYSEIinsIlDBpoFwmOnJqLMDNR1y+6FNvc6wKw/3lQAAIjNDe2nvN
ikfDGWcmOL80P3+GFte0T67Nlwg0rVpdObTgIg+CJR7XfkbW6gFx9Owv6GVl+n3e
piCFnKSLumhBeB1y94Z5fH+w0HZF4xTbVUL8QN9kHNuHAursLjd9KSeqlLJADXR0
6C7MDzWijCh98Fzzyn+GTMTyAq7Ox1zymKkAvPbkYwaJWJv95tjvYatyNwUomV7E
GEzCMzjImI3JtKuPEZRU5fkAG48EZ6DjjLp7gqS70WmUqI3stm2TIYmevbCRtUgR
YzDDhJhvl8R+E3bO/0gkmsCKQfOae7NKezN8gmsas3Vcrw+0LNGJ5XJXevj6DzRr
Q2jxPBcqqn13xq23hw7YDp/OemsZ8IT3h7m/hnAldAt02xRx1POrKste651cPWtN
rmnxd9U0PkmiHxzz6cq8M43nqKo+EL3rty285aYJc4u4WJQdIQcOHwfqQcmaLR2x
aZ39wr8ZMJxiMbuaa8KzK4ySe3RG102X+7zjHP5zsq/i5jCzF0oVclNucqoTvqnH
swn+chcufx9CiiCOJCFvGkvI3jdsF4OCzxVnqDTPgEHX5bUEEn6akycK2S8FGQUw
e8WoXdlFwy/rBSolpL6fFV+v6xlXLokHFV/JrsXQBBgV1kiVwrv5hNluxWb+dq9v
8rJPiyCegdJ+UMLu94W4g1QNHanAFQkSgX9thl9B3IJKLCFiksY7kaZYCzt5BH+3
AtQdfsIZ/cZNnTAESQJd37i5m+JnMxZ/vgel3hacOtdiZmQp+im/pInVwhuD01n4
TJVxEMREOTlrNXsLk6zOKyyY5OnhB48JASJ902GPY8YhTtWjOyFJCtiFaycy6U3W
7r6oDKEQZJDCaJ//dIk0oyalWvwMNvwlK1WhSkIFvpbpzlH5/95y8Xti1akk7o/Y
ifgjE1KW7M2dOKKdWT/eR/u3+YWDDvg9ra3iqJnYvLtHEfeQihKu4Hbq1nDKwn5R
QpDXhOwxR/PeQkYEL6wddYdeVkdAWkaWlIv/rSAgluRIpzK331Qo6r6OkMPQs+zu
V4XwanotaslFJkk7zuQ1DHYGBXr7mzUsb1Lc1OuVsflxKoHitLWZTKsAi8tNFoJP
lo6fdNPsgMfTRgq5rNIPeROyOhIQGs4DlZu/vX9sU59smuHQxGRtUQ4h6VEiv2G/
SpjyxHqQtqaJqnrWwZ2gWBs5k4efN6AiR8HqmddORvuxQCSaUAc1orToUe8yL0QE
2x3bHGOhkMGCOJAl5aGnD8iSNvGnbMQSAW7GgyzCLrr+zrDINJkFjdKi0h5TvkxF
ZkuJKmTmMOQNxgY41VJ+pP+XUNfUk49MK+b/wZ1ef4FjrSYnoStNtYPKOrJlyS1B
LPdirbvhEU8Xf1vGD+ot2tQGBZtbkbigMPoseEP7foc2syeUwl4nqrsnCShB+vut
kKfkqW9OIB0DeXTkP+JPnPVn1/cTvqpIXHUALcdb9CzPQ8lphME1TLWYwL4sfOyj
wOkWDU3L/X6XOelV0TTqW/YyG0HtBoXrF3LU9q8q6NSjPz1lkKOCCKSBdmcTPzWN
uaxLgOlYGDOxTxVF4weuIEuMOFDbB+avNsFSbOF7hwPkp7/91mRUkm/H/z8wkX8Z
rVdXvMzxOWOITXWoGyawHSx2ThOnWplwGoBkqiMkNnXFbUnfOB4vgMWo54A5wKJO
2kXbSYiY3zwlkoTJ4awRU5Qnmj62pzbuDyv60f82gD6Ia2d57MjFdZttfIpb3pQ0
T4tbhqSUSCdvJ4Myi7MhOVA4vgWFU0/s0YVNewORd7oPrbvSVYLhk0H5pA2g5w0y
ksJYsfl+Qp1Ccde9FtV33x4aCnEqq4tGI8RLa7iz7u8EJj+Dm3Ns6ylpX9VNqXLi
DLwyv78H8VhO9I07W7xC54eNteJIcBUaCO9Ec6ppvbPCGRP2ppmyV6BezydFoml5
hbZXvr9olEEGai458jfBjYxvqgDI3u5IOFlx+qriGIvRG4Sl7LEPvERCPjRHE4Pc
6s+m/7k5QE10vZJtiFNAWpOBUr0hJDJ6w7nn8dr5Qb1pemLM8o6d1fsYxT+fensr
HN63kpYoo4nlQIBBS0vUK14hyNLBEqSBSLQvcRaF2G2E7OABb75b+WKf0jwFV0+i
cAaweSrH5NS6RCrQgHHmYH8oojsIyPuHTL7fOrfiVtTjW4Irg3Y8QIt+zeoygN2m
pjYkGdsevnITntuFHSdFlvCMdVXw9CpmYUXFsxQYwlPpusd96pnBCfqlb1R82WnV
V/C+6wKULC2tS6lCigtfGuUmQi8JELFB2pFqRiJBBaFJvlMJpYmT4lGp9SfkgMhU
qbHGT6TqNZxVfIYTrdzoEWXnM/SZPmfU6pWJuQk4nsfBrffakpafFASqdy1VW2yj
vt/vCR56wmlfR80sBz1YXPBfpK3gYIUJC36NlmEXxqiVqMd+Pqk1qITrSj5fJ1ID
FGjr3F1VnzAoY8CNVpE1+xIhGneZKVp4nh16gckTzaTY++b0bnsEpq75EZkCJmvr
wtJNAiVFdEbrwkMnj/wJ6GqFGZbyaC0kKsjTUgbhua5b0aHv1/SxiDsbbdeKuNjV
ZKabKKFBH+oFrXDtBQ6Y8p2nMkP+5xRhjOyMxuwTbPiJ0M8e2706C1sjqOS2xCtk
m8fcTM98wc4ZFGx18OqR55Xws73nOqP4wTNBbLcY0M0tyEDGfpFerV+CipIiJHsr
RoXmi3epnc6/RXCGZpYmIOro4nm510QFIq5WMheUh5MG0JUnxKW7O3e3m2OwY+If
QxcfERzam9gip++hdulMU/pcOZG59Tva3vtV+5VopSdbbQU595zd2s0BCe5OEsoy
CK50vDW5yDkPTWjG+lZ1EwLCbdpktZX8S8rJhXt0fyFAAxW5z0GFfPQyzxPC32O/
qaw1TAmb1lBVsGRHht3gVhKrX3QauqfI/bNBRD7mTV5LHIGusqM6U7IKZ3fFtrjb
sWdHMKmWxF3D/Y32teoheyGKkdGY324xLspaWGFrQ9ZIurufMv8c7hlJ/HV6oy+B
K5HJGehLJAUK01gi3NXZJaY8XSXrbk5Q196jRD9aGYKTSoe2ATtHxce7rnl7P7I4
N8YfhHxLGhj4YFwDY7PQJdC97pMZImeguZG56+kZZKLvofQsyQMlAsz4Fwjhq99z
wH0MWNhcTff3QjRWr2Vu+mGL1jvACTU30qaMHces/SHY4bi5OMyzH22oZPM9EkV2
K42KOS2K8tlbW78h0BEm0e8M9xAHMb4reiCNZwxGfFiXnMFY9P0U/lliJ3UURpGt
0D9pEp+SeX66fcHVhkkNbXe8JLqbT1++gIVV4FgpcFqEJCq3dI1bPTNxIaNb04cy
S3jLS7tUyuAlh5zi71m0Ew6b+V2/Qx2+VXK/aogdaeAXoNOQuJoeBTafnm56TFgv
1QUelvIWnVvVjaz2/KIlnEZXf6W7KwPcDQEfugm/+GSLa7hw/f6Nx/7hllmuON7r
B9mwKIR+ootbdWHizStsgHPG/z+zsC/Vh/rX1LcvJ0cO8+DOMTwhkae/PpaRbRVh
DOSkxEpD5qviaL86unQAOnZ8uBoLWe7UjFYv6CDz3OSnlACODgtJdnUftJ6+4LIZ
qQKbg3SjNAP7FA0NNq+7H92vlCM3jQZ6+dg5r+0QePaZVePXDbRJ9K+JACvqowwp
IjmLS4crXPpMtFfgJBoBcX/ZXWSLThwGjdz3HadU0O8iabwgo8p38rOWVmpIkj8G
AJVpdeeogXM3KNoeEgg0eCKGfaJcHK4SGMo7UBh0KrUmp2j4pd9Yzv/uXU9ST7yS
yr1P6RYeliOrkrBe8IdxiQyp3CeHJYgHwnYhhyK0wiy3UpJSrDXS4X5FMcurK0Il
yJeDu4DZvbaPg9lXDK/q8ddTyT3gIu+hDsmcmY39ak6Ql/ZnH2Kb/py7r/MvlTXL
Pyvug9NHAzWqWuneKrUbFSUkzm7wopfRCr+Uub44DAnGfmEY/T0gH6+zyCLWJURy
Y4XURuGowCNyahUVERSJ7CqlyaTa+z1irZHvbHyHZq3omYPp6+RiaSc1mpZth2l4
Y4JD24ePvlESEUMoXXsAbkrhfxTd2G3DTwy/YgXNXl8PYIdGrvb6DNgLCKAmUH01
Z1UqUPDbZNaBEbgBxBHILwWH4nIKZXNJc6M7rup9027QKtumBYJt/FooqOn3+ZUE
OnD/KpNMM/3OQqT1+3mLlXfJiTnuxOke30vX+QnpfUoohsCf4lQ8wMMb/8xIm5Er
9wZbKAL+vgccE+HlhETdeFl1PRp4RveI8b+/iTgOFzwmlsR3YwO22rlrO6Dijo3A
d7akDSRg1HpTZxWRg8y/Svbd5hiRUDH9yXxG/addudDirr16SZUeZf1O+d3JFRLm
KJeLBBNxdI17/luWfw1VJBnY4oalR4VF6MpVkaJz2MhIKSr6mTN4Y2eDh/SsEzqi
jbA5USEgVPjeDPprqvM8xRhLuAp6qcNrujYXsWqhLPyqemtHvqP6bkWCOHttP/0s
ApCkSIcd4NAYUHDM5LmOLzton4GeUZfpz/bnblkyfBemnuuFceQ/212mQULWBESc
C35gWxaW/MD+5VM3oajZQ1Vbvrr3ON+C3ebZlnPz/nFOPor/PsEYqJsvSd0mX10B
Ge012C2ALTSLV2xNPl2vCc1xorkUD5wFL0N7klXNNE72u+fa2eeo/O9TiNjAvIZ7
/O7QLG3pA5+vR/ygv0oqUuBP0gGLuHhA2C3aHoCbOZf2gb0keP7gdN0OPI9SbtEu
l+NFi3kFuB0/lhnjca5/O889+ob21zxXyrf97vLYFYU5xtqbLkQi6+f4E6PqCZnx
q8Bqs4TqWNiDfRS2YPmcr61OzF/GlCyjJLJV9E9yMrbPzJVUFG87vFjcNdtJi0z/
aB6Q7UHMx7mi+SS1uduhe092GeoQ4ltpUG6s6plHwiA+ds70CEW87T27KOhWILob
nyL/WXIaBAQzUngliSdZPBxB6lVFeyS7tJ83M6EJitQ51I42PLtlVvqO/qXF3aS/
PI+fQktkM/FFQrDuiJmE/INIo621861nNn1MJLh0nTXKmahMA3bwKg67VCn4ID8Z
IczZFYVmcIsTx+hrX702uwNBqoBFAKwP7qsLtuV+c3a7svaFqAL/iXSKlczkmnFa
3iui139JjNPbwCItSdfAkR05gtFu+T8sPz4h/w/0s8ZVUc+st/NLoYexF7qXqNUh
698le6uDEe3QLqsYH+/nWsrnj125uGL5x+kF2WxNc9nbooi+RmGmMEHmP2O+LTkT
NBD+e+zURLmEHU1pjGWaHRj2pTW1oH826lqYYCt+IaE+wL6cIQLRDHMldnDh2qET
k06kAorlqllTBUvMa0n/d/fF7ej0xdQD++hSajlX1LbWUvqkghEMU+uNVQcEf9AQ
XAil5Z8kvoB4of/8wDQnmFh6sI7ulx7ev0zzRPebI5xK4PhBB9PO+1xtnR8ymecc
tv5bNkRT6WtHvQSbcQGMjbzGtJxlclBw3rXG/QO0+alv6rJ1P8DO7/ILNt6rcIF+
P2yUrjr/865l1Xf5XTitMhQEAMVYBOndgeLMiyzp/yteMzfboO9vME8JRQRv8ZrU
813t+apASY5IQC3wHoPCD44qkZRNe7JQkdOm2yuEu4J8s++zW7vRk8cw1nkS3KD4
JHyZnxjCWK3kLaCuFX4lDQfkIdH7UVBazcyzPk5XhWRShjh+iLP8FgVoUF42e45t
3T/jNb1DETOd709FbNu4Q62ZKr/kaKiPE1K7LHRskF/9JVASnMz+8pN/ZxZG3VXU
fZcGWosgbkl6JPuNTdDe/CGX9s0/iap/ZuybwOcIvtD7w8N3KIH6H4e45uJCrvYH
U4jhXPj8f6Y6vbJYiVN631N1QyWGWd4+eWRnpmE4ifpkGsKlw95kI8mL3LfyzcRe
rvy4xIUo4zvpJ1OQ/5S4MTlStswiZWih3+B6ZQRkMHsDmip5Nl1FcOIBqzHfJ08O
JBZ+k5+5G2M+hNc/fpeXbGgyCXwCyxYKb3n/+BWpCAI3pBwPBzk9pkREf1uYmSYN
vgqIhXwEY8sWKcWsdG2eJFiW7aSKgY+1wguOJx64HFBndWblTjUYI/XSPRm8UXNs
pbTp+ygIyBI+cvJuULIo87SEiVDdO/4qTgmp2AWmLeYeTut5Wdi+fXQc/HVCvfLf
0qQVsRmCffC3honorHxjA4yMy6yamfWjJAowumQ+Irzd3QXEGZm36DqKSRWCJqcX
c5vkbQtV+wO+fg7C1OoMzsIm/1Dc4n0gYpJMjHKy7iYGpHS8dQWkw71fM1203or8
aP77mlhcL0pJIPlp2ou1LrePnBYlB043xO3RdEyjmWyq9pXomMjLC66bJqkb3oYl
u+nBCYfHUNox2DrcWYWpZ6S0I8ISFDZhjg8aN9ALIEK/Zm0NugqUZpfo1W5CFhOn
1mMiK62jVm/7/cVtImD8MtW5jVceLqxef0IMgoUPJUTnfmExYDh1qWxFv3hRpzIJ
W8P6I8k5KeWjNDxcH0iuM1an1cZRHverUQM3fYo7NJXowXyMx6Fc0G8cQTGYC7nL
wwnF1A4F52FpIGagMHn+L83M77BG86L+z1dSYuj7jC3LppF9KHfCVWncs/VknNWm
Xf4D99gR+IJRLY6GYPC7rLmlOM3bYHuiklEboY/KTwTRBqjaLCxjd6PUcYXo8oK/
/G5rUrIffRSab7voQZQA/vz/YD8GuolVjf3ZieZAJhspnFm2S0mSBf8+JhZhZtBn
sfm0PDRK4nGP9wAA69lHf29Zet5hJ6jnrJ7/crhad/e0ZRy/Lijk7kyhp9tkPfR7
mTKEq595N9DXtj111ft+6/JWLbzJ7XTZS9XaYc6Ew69bPAwLA1aV/BWJQXi/ZjWc
5Npbv+hiOOJ/Uy31LM33mNrtr7UDCNorMMv+uZOzXAEXk0JvTEUDN4UqMZ/TfHfF
dT34JJ+wYhbSjyEu6NcZ4+haMy2w2gG5ncvFQ5nLUGOYREVuzg/2pFbg8DscUhup
xQg47TUP5uH0EqIrMXxy25QRlcgx9N5cbt/1vgos1d+ZvyycmRaNB6UvgHwf540/
y8NW36zSD9NmimPJmcYIAuSrtGQqEmvi/3fyu7Fv/fq1sCeOF+cHxskv/yKrczXr
xtaWBrhGS40IIMsYiNoIw9DBwBQovtthC214FJZ3rf/QxLoJUp0+gYj+Pzbd1gYQ
Ctrc3yUPtmxdVoVrfGdnOpkY2+yMhOI1G2CTDraWWwzw1aopfAxuJcYSefaHg795
hTwWjnLTZJrUbhcfX10+vpE4twuavCGZ0fjdK6fnqfU15AWedK70a0isfRLrQEp3
iPZ6LH8YwVc7P3hVsSmEYgxLK6qX2ZNZaBOgOng93LCyjM0AeKPfLCBuvbbS5ux+
y0BROHxaLNOPEuJ8LRgf1t/GKM3+TNZ7y5QajfOT77djHCte3gcxjjDLJGObLBfV
YBJL7gDtmLd36yaMkprzFWSGiuuIRLQ+Dh2AZS94d2KX0EtjMvRDLpvAgecV8sgV
Q5djRCLcU7Ygixm8+okD+pr9LaRQrh5pqJjAfTWxFw34zhqEQ/6Ugh010L2iwp6/
RPgT0oJ0lW8yQKxNYAlA4YWVckrOamUVqoxnmTKIoUdei7rAF7afa5Y6QWyEQu7W
q8z3muDJLt979EK3MLax2lYNu64yjnaJenF6a42JLFXB/XZ1fuFHEX9L/3lSAMvX
0hNgQXxRuvhLE2sw1ncCFwKDp/d9247a8XvgORDvCMk+0ZsSx/8eM84uTFuD4sYa
E2o52GiDTISRweqNjEQ9EDUocrrjlhW8Mt99hjZjD766MX+18QlNffgDI4p565qP
XXx963dHibaYrrnouSR+N57GZ+XKDt2eTV7p4bJewrHsy0GHNgwBWVG40ZNGWQ3t
FEIOLTyGv+dy+tfo1VTWdkfrabU5/9+CAyG4R6S3jxkM3PPHxzsbSiEmwF2Z3fVt
Z6MJFYhNo9ClTjlxNBkqOL/mICauzv0oR1n1hbt4/BLi2SKA/6mfJpgp6pk3p6En
Dj4fNlSx3gblUitES9Zi7EBU1ZAJCwBYfqD4Rd02GXL3d+eOPDS1Hf1s629/5OBE
9+EVC6u3hkS6MxuvGLrFVufQrot57sY/voJbwr50IXZWZ9K1nJUmUZn7QKr9tafE
4VHJNuVi6BFqOzuJIkmncKvhRoFY/SYvPKObj+OOAeLorVqdNKSwJsKE1XT2Z2Ef
cRFscpYlBpo+whv/GCrfCTJ9mGFW17txLIX4EBrtNktqinNn7RgQPQ2iyLQpMfcf
pFu4Gvq/lGejoSkf0OCVd8ZttuNrYRbTgPfR0p6Jvs9w5uX0AAYCvVbntcEVjlqR
QICIU1hCu/L3b/7M5W56Pn3Fs8/mxETG8Tl/wF2a5gviYc6u9gD5qtwRILtwZZ8M
8LLxDCQSgqnBoTxtUzxHwvgTE2VwNF/eaCevRnePMtUvesrjHlke1DnMndIbMqgj
AYMCBhujBdimeZ0F2oOdmulClNwdaejKi54Espg9GhN8pQyD+Ry0Y1qUWDenr7cK
QbhvC6Qxx8a0je7KzcyqqpW4k+81P49s0jbS2d6LphViZ9IJ4+h6ADtoEz2wTJhO
dVDwnxWO4hF3M9UA1KFDVB6oIHlBzf83svPKRQWUmf6szEjA5Ydsu84fnZogNq8I
HnSwmPtWVARjXndbnc8U13GgELWED4w0T1Pg3ArTYgF0buduD5gYQ4zf9DHOINdB
vRsgV7eozqYi72iJhQa0OoUfh3MB4nkkplK1iPfXRlMm9vf8Zp8te8KHFfh+1UN3
qnj7gWuQODsoXHfrM/Me9BMu6YMSeKFHcFk/7oHHdt66XbA6+xwD0r8WJ1VN32ms
0ZuU5v0nzF07w7m6IRX1oyJ3CkKHgNS5NoOS2PS/ztZVQUSiwAgGFZI0Ahn6IC6+
TOEy1yrrIG0c5zYaIS138/0UP+M+aRh1GQuONNqCNFzm8VzIsehXSCklBgR2womw
Lc7uSKgIuj/Hal0XwJ1iVaqTlK8bFqlrWQQBXbkMvlnTHEGpWhDBGcXyVGlTNv4E
EgbszbpDeIuDWVxMcx6KCRKJWVOSBu8sVxpUe6x9Wc8300BkosgSKYZ9hIOs3ngD
t8wr5NBR/DsOz9S9yIWlqFCsJVcAZfAa+JkCS7J9YHX5jt8oLqMz8xdShRblwqXN
Hitqt7sQ7HyTovIhygJHzI2pyzwwOTjkJmoSc+znmeBNNUIm6P6Nvv8PEVe6qZ6p
EYkSyV9T9XyRjJYNSbhSGj8gO89Tr1DvAV7qucuU1HyUYl4BEPa6M/SVrEq08Yth
jmX1WJUwTPrndgBvM4CRBIF634PXzwBEZd/FQTNQQj1SbHx2u0c9xCqRXo5cO6Ko
6ADuDB82PcqoYQ/6HmlORp7YlP50j64hO6wBXKlmMDjkT+7KCgBOFFqH6FTRClVx
yoD06cPHo9mxLuKdzjzls1yDaTpx8l/P17ZlFO/ieHRt/Yko4rM9pDYhpkAxqDlc
pwrIGt3wPcjnaWnKVVc2T6gTGiDvQV9awK5vtD5GrMytI4LOpvGhkgoSq+oXB2jf
co6jar9dd5eBmfO6IAV8PrYcD5/r47MuyPOkqtwoH0QNBOOnTZabbyZYR+yzWZUE
DG7o63CMJgDpBmrdW+W7gBJCU7uPfFY7ZIGstl4htWwxGGSEtfHagwmHD7vlZO3J
rEyM0Ta0yKxURY7RMwGIm8K1Si7paHK52xnZza7oUmbv4t09gWbzVmjhuXG2SEYe
Yu0ULMWSo1zgbe9U3emM3XYlJZ8kVIYqWLn8dOjmm6s1h9GNoAy78fLPxS4NsNrt
s4D50ou3VLF9I4ivLQSzEGHQ5LB7KYB4ArQiizi40nSRCXvA5IhnyszmpjqqWqDz
yHioAJChv1TGM1kMr31cxoJeONN4hhtmApZxLK/1byjPMZ/4VO/+aiwJd1UyA1j7
rx76DRzDDwKq4j/vZcoNIApRayIqcFEFKG9Tpp2Y+vmlGfDFno6LUmCKdal33kR7
as2fTF636voToecppVefhWMW9GkVkPlxfwPYtlkQvRrQLwJ8XhBo018r0FjOel6F
ASP4nH6qD7wpEgIyeNLcLaucxNVM5e2kk69X/mN4ippXF0DEHc9mNJKPlUyEPXZU
pI8Csb/LpkRRHKywFIWY3863RULfYFD9YSHu4apBxBZjqv7eA+VnwHc//+0LA76C
chcsMpKgzRA4aSgRGNw7O6shXnU+dURs0R7Z3ivx+TmJqsv38xZQ3s3n5nXbODEp
mFWpAGDeY7tMrwkLQZiUOrPhqxTFfQXJFVRbF7Q9XBJZ8QvmX+KL79GuU/eiSp/9
ZxhSZCrwLdMD8dpi+kzxtvSl5YOT/8i/87l1CXqOOUZltDEi/SJY+qb5Pmk+lerz
Jyp3i+bYLrxFyXWqyXF3vEze7xXHYU25t/yDm40mo5uZIpuPgW7v1tH3A6ENLGSg
+uUrr0yF9YL8/KvhMyP0B0xicg7bbietDvKwddQ4MtqkpRaJqyhWZR0q92CQuosB
6B0tleAYixWghRqxiAefLGlSv1Fs0cUDHbPqMkLOcCdGMMcZm6bEBXxuK3lk1ojt
rNFvZ05U7Ry5GsDhnl5Uww0/PrxHcVoK0eNF17ey/hn8sTAk+fLfXK2XLmSxK2yf
pbR54lV/iP8E8MuQwLhZoxpzrPRu9f8IIqE1ehG+JwbDH1WGGTve7Rqlrud9kgjA
YLjgM1Vwba2xrAPmDemxB/UPvQf6xgC2A69xWfCDoV8SvID5wWygbuAUoRn2ApQQ
AGVlCszIqb1GglKiVmNIKNHT9qRpC03nO+FpYXP2S8CIoG3lKt8cvY9ORMhS6DcT
D9OFoTuIl4PbnSwjdOK/Hg+bn0YaVYQLXBYfkF5zhiJzOPmT0zXKBr3Qz0HFYjwP
ACCCPmZMBNJXmP2GcmOnqXxSnOfXKTKGYdRMGGDk0fwojPrubiF6sa0/2KPNQQtb
ZLjz/dg6wCcfMV1xp1NdYN5Ys45kXdXjb69DzzgpXHjQ6eygX5eeAO9MVVTQ+yln
M4j7G3bbalwnQzOdJcaqtyuaexM3MCSK+G6nxkE4h8c6wKAzLZPECjrNdZMpRNMX
3LqjEPB365pEqHmsAQMWHheCJXKGleZEpfhBX6V1CJO9xzfaPZo2feVxzmKbIrjE
h4/8ab08YZyEFSQ6PxsCf8Slu7X2keWpUQ0mhYLkVw488upFl6e7I9U28K23AKpu
3WTyYjm/+fRI9JVDDoIPz/B7RpQbwq3PT8ID9B3nmPU4b5phVktPcJiQrVFKSAgj
xKIjH0hsuJ146pMASR6qAfW3Ux4T96jBIwmFk3eFgNz4rZHIERlUEk5PfQUZTycu
MuCbg3kVEIiLZFUUC97BOsKzlk9k+Pi6EVEcnxjvsY29FNs8pPrIIwos7rJ7N6PC
2uBrZWCGFfR+0BAD3Y0s0jj9KT4MZUmLi+4yOwXScqe9KtQnHqxCs0mGpyQs1DSR
fNYTCKCugz5pmF5qyFperffXYen+O6WJKuMyMzWvAObXaOC+7iVmioTzlWCZFBVJ
llf0bTmwOA0yxANgdRwTHoLOeTh1lRDMgMQJnjnA9D5R1itbqvKFyeJ/4+vvnTTb
D3nkw73nKcC3iILOBe6feVRyJC7bFlH+wlRmf0L3hCkx/el5pk0sxRIv/CxxBK/V
tLDqFrHQuLy28XhR48F8s4ECcW4zJk1XtTB8tFdAelLHBbkPcLDaEUYbEx/QqJ1z
5KfXxSH8MhO0yGv5LoJzUmQoQYRtQGJkXPG2sjEL1twjKDuOvWcvdyXOmEqACzoi
WFcLFbChMkteQ6wqWhReg0oZDEzS2iR3OCeIgw9NcUaCkMLlS2Tq7L5zELV8Vev1
N/cOaK2AhP9v40wrRTa3cCtPL3qAM7GWXXgwZoMzmk0Flr0mzSKXGJy4HzXIWKyw
0r1lfXXpoP1gmkAb2CM3PGB6oL48Tdnbb40MplZKUsOJYq578VlFsncfjVz2TFO9
s8xjI3gEQogb7aXsvyI7gxcbNUAaHjj5/LDa8VLVjJObyTFhppDXmhYlUyjF85UX
vt9xUX4xeGQ88MTKMKiwnCMg9SOQeI+QmSEQ7VtdLbbMmhMijbPK464RI0276B+s
DcFW0E//TWxIiVtCCrt/h+V0RV0ERtva65RgfiNcAVqxtFxqvJ9p72gUQ5OVrh06
YtB6QSLAtoJ9vE0+9sD8Pmd4Xt61MiuTCpz+lhwLBSwbjceiIjvziaTzzZ9HtljB
YWbtopAonlH1VGHtHJISYbysoRv6G3BTV9mhgrNoy26e6C0ZXdcrhGahvwN+mCLp
B4mg7hswdmePPYowvRd7ac8Sla4dQiGE9xQEHrOohosamP79xzFM74Ex1lT6sXqJ
fNGCF+i6eEnqaxkUwHFkEFEuk5SstXIx4Bfh8h2Em/hL+JdC8q3+F6auFo6UdR/c
ia6ABgkoiVPgE6IA5CjnlJe0Are+m1+Anky9bVkpUSim/NADEH8vOCPjWPB7LeFC
YcAhVD/cMR1ZVgT38mGZq7QEN/bQ+WsDBiXcU7smg4oObaOhDjLiZQn88uq1XNkA
VeafplPTQVeu+PHHuPIsHr+FVqUayRYOLqazElBMOK5ZsQ0RnUjW8L077HDZ5tcZ
wZAoJpTn2LO/ABWp8/hOL94Qv4e4PnQwRw6qGRgGX/QSNbTEIVukhEIT8KBGypEg
Vf5adLx1cDzLhk313fNJjeZiVdMvyY8pIh9hJzW909muHi9bkjtv0gG4p04+47Wf
2eFVU9+qAWOFePsKemAari6h4l5AIQESuk+3SVfRxSIy0igj/rhSzyWtT6d9yHju
FuKgiJXaATivqVFnEA2Rrjfoin4JKbEtaAIaGxaJh0H0n7MzB57XkSUunoJ9vdVY
udUxlMLCpnJ14LsF0TPON8I3w/7Aj6Nl+ShMQ1w6qF6Q7fVjwZ2g1cPVuCZ+sWyT
00SQ+8VpclgnixTGNer4Ht3rR93UQ7fCeopuL9y/CCcETBX0lgdop4PRrin//feO
lzd0G7O+iuFbRrIfvGMbcTDPp3yRrOJ1J8I6dfwR1LAx6cFIXhK5pv9Sw0UnWRJS
6DcQ469oVhBoQcKbWYVC23sOuDOViLCorh3UejsFfpEW4UZt/6kVG1FzW6KYkmlW
94POCKsAWkJ0dD7mX6a/Dj7cm07DrAZpKewCWKHbEjhXd/QM5XgnfJgvuS1R/cPd
aygBNga76USB5YiG3rdEkM4MHeQBFTdiVhwn4LjbdDJ65MUG9WDU2eXZ15nLPDE9
KGepp1oOBsCvysmBZb5f6oO1LxkWgmjV4hj/L8Hy6bVedYK55j63euNXkhFCV9EA
Gtim2F8Q3LRAaIiXTeTfA28/REiFODr+88lHsrGy6v1kByGmPqphJ26LH8+tST4A
qUt+25S6yw415A0achoqKmC4J+hKkAV7OpoNLxqdkI0p2WaKMaNTd1TLpEIWhhNT
qovhr9jvnSpHQH6TN3gPcmjJanZI0aj92mZj85Zp/jlqv19w9vrwjMbg+XUqxdFr
yIFx8SBnXOWZTppFEyWfQ2ayYl6JUCjnm2Lxi7AQtb52FdO+QAAlXBkgGs7+HpuJ
Rc16PzrvIlM++9igoEIcsv2F0o87gjPqdjSgz/1/BQPJ96/8hHfiC7y7oI1FUbhT
31Tkp1RXGpF/0oewMpYjkQhLM1lgB2gP2B11iItMdjjBbb+5Z/5n/9JW5S7r1G8V
bNNqtMJr0jeK1Q4AmMvmRJeb0wQZJa1cJ3KNw6rFHrl3+0/hEZa9bYLemURcwKOJ
K1dTMx1KqwwpGd7urf0sFtRiYX1caSJgPDH17i2ZIum3CGGhJe4j2JlYAio+FN/F
aD2PsiO9ZeGDR5Dz/xCz7BdK9EFBv/jHfMlTNOpNiEhNMXVnAcvbU6MGRKwW7gLz
088bUAlkAP8iWn30eYygcEtMfJMZbyCJ1Qe28pGRhDgYmBFiGcggQWY0US2gKC7Y
g9xdB1BHPH7KprYQwxK+3YgRMHoSMlJE8dVwkHWCr/bmwpDDYnn47FvvqUzESpq5
9r/8kT5CK/x4EVxl3f/Y2QrgKA3zegkwSHASaGLto2MXtJP9M9T9bY3rSL22N90R
auRwlkB8FlFuZexoPrxMJqQrs07Xu7aSF6PHPyeQ/PXz4iV5+WtNXCfEKNJtdRIF
v1ZeD7GaQhwU6n8NIGQ0vbfRPN2zrQz3UTXOCWjSlEo6MHUNspVZiQMW5icQLKnb
LnHxJaw5YGeiTdIuEPat544CRMZgyB0e6kb1f8KV7WS0OFvVJRA9MVyofGDrCKya
Mg1/vQ9502E9JZyc2KTyQzr2fx2NpNVzhJ9IgISVKJvpLcdScLWts5PIzphsb6Nn
H5NkxkTVA4BwQWTnP6AiqDWK2sUZhEM793LeTtXdww9cL62p7GReJO5ubbTb/uUd
rN7bF1Y+aE+d6UJIY5AiQ0X2Rnvp5v34OU+ciUCBX0mBXhfIBqNqghMG3diUA6zO
9wUpoc1V8ID1awGDGE+di6KrnV7hcyUCba4wC9k+Kxwbx86yA/Jx/y+ZTTLXJyHn
77xYCt7OLgMqbDLqltVqF+EhsbqOxGlBbS4Sj+MVlXMO17IbKFcYAfc/m2eK2u31
m+6YL/7i3Y/GcId5vjLGlkpMAJRRZ/Pyig3+7OCeZMRpmok45hbmOeS7etPkyUjr
toEhrdWpFU27S8vEzl9PBD2zToDXJ5fP59Okx55PmmfpQTXfKt1vPwT2oxLZ4Ry/
zS0xIYq10Kb6EsRDOs91VJRZQ4lnM/iS7/VYkldk26zFmyIj2zYfsnaGJxH0H6FL
sOuQSLVQoVnhnetckmojsbuPue8TG6v34n8/AqS7ChHiP9hkpyMXavWxGBrCKITK
f+InJyJOgbzj7nSCUJT2CkzkKMn0Comv2iJNO7Yf55/86ETm2uLmu1sWr/pbsL1C
qFHQatv1n907k0VacxjJu5GqyJY3CV3GYawCNG6kG3PnDJf1BlSKBuR8f/zPYPoi
7TBtw7Ab5p9oofsLotU1iwitwm9cQzqnXqP8scMybhaw3egfWz9nv0wXPj1m7+L5
xm1tyFcA4M9alLLQ5z8GkOV2DrA6/1tOvLn5Jw3wlI5ifZN3J7jzc0iz0nUT2FWe
DOcmTzQIvnOkCLjzaMFlARWWBZwKrem0C9q6cf0bNIDskYEyc/A+ZT4y+74v59NS
E/Ve36Vhq3Jea2h+6zY7HtxbkQ0fzNvUCcEehKb7bO6GS/xxL0yfloBDJIxwzyNm
JS05NEX3HDgvaND7uuAAxuMgKpAgJfChIVKsLs3tLNsehmFG3W40B8qe9SAzGNVE
CGrmag/eWW38UxpnUUWjd5Qea+4lktobJ8qQv2TsVbGntf/XGdvXbsNbIa0SsqiZ
iDZfxxpJHoH3SakAOZ6OonZvX+HMDGK24+KiOGwATiehKP/36itCOFBP4VLdTFt/
qSuxewV1o2sTggvZUUqiGSXt6DDWpPKFR8WNjSReeH4BBXX6IX0heyicLnDOpUFL
NCHpBZCT87W5qDsuNHckLcvymj8IQVcqWBET5TBg87DerRwIir0TxZoZUtnmJB9q
z5b+firNqF2Ememi3c03uWzFm583zBcg7ocbLIs22B5IbSk+AKRm6ANdc9p1LuHb
u3CMn0ourVAstyn0Pr2E9Ylj5BCospweDDU/bXOM+sjqqhngEJCLcAGDVQ/WQ9bc
fvBg47/jLxDRDh0XqFiuegpdgLLYkjzQ+idohASdgTP/OSENq4RGqdmgxs83uQxm
TxuK3fdU0SHL3DQbfUpmP3LPhMIM/Rcyjhcqp/rtPd2XNJnSa4dCn9dV+tnLSr5Z
cBIUBCc/5ZUVQ0CiNS33ViizwcHga2BJfvBrwzzbRwxfgvtDHnH9ckeilRsDRrg+
8zjWYoPfKi7dl35bs2cueQupAM1nE9r46EyggNkZwKYFNi1yJoQ3NzDIJQY7G9ix
YY61yUuyATnKceX62rpwFenChh9bsx6Kz7fqITBZ0CivJVSh77Tk4wvwyPVtALqQ
O1uvoAt4ujTwvplWy69o11GjFF1uTXt7pmnORQ/j6AfSaRrKP5P+d3xrrDNudv7o
TqwcRxE1HFBaUuKKQE8/qc8bnHt1bqmBgpfCP2W1XOmeNdrFd5VT9TZU3gsQloQD
Znj6LzTKvEUxKrR2eCihuVwZaUt6GQvLJ1k4K0p2Y1sy2F3h3HGYhMdGVmyWlUMA
2e/rVQPViyYLy4mrlw4yMQ19T+ldPkzhddLjHM4VZMqkcw+Wt7pyWQFcXnqALrKA
KiF8vUipcINQJwSzmrWwrt6BrDmqtr9y6ezWoVcjzfEisGZ1z4qv+K0Z3QEKxjDc
5Tb3pdki4ZWoPSXuowU45mEcwAByVcSQcPI85i2I/24gJICpT1q7I5ZSiGDZPtxa
g5C2JX/+0yy4BPAY2LqoeqUi07mE+K4mq6/d0MKK6knBiLkWmWdlzOUfstks+wa2
vWYERL1zBFWr1XU0gjF4VSKIsJcXd1UFR1Lhj+hbw1S69f4DswDEufTQA6ATFezP
J09d5TVQ6u/0fwLkwY/UnYz88MKOxa8W2oKZVgzAEKbC6Tz0MraIKtbRHxWKl9jO
I3xSlFUj30hd0dtG3E5BiHAbiX305BNJpSDwNR7dODXOSuLxCUrmwOtj2U0lD/ZN
KOByKGjQc8RcF93dMHWH+jSVFp2/M0/PT4XFGEFXfAmgkKya3wZtIxNfgxtv3XXS
2O51ze2uRzoGl2pBcuUv5CbxfG/iicwrvu+/Yv6D+IS3sGZGCivmj0HKOOL0qR5w
UVMh3gTroJf+xA4KpMeWu9fUFpVifOH0cPGAx1ypzGRsDn4E9oliLkmiAs7WDdv/
Xa0ucn/IlP38Z/8hoVUznqxmah0ZHjpWDkS/kc7+D0SGP2NGxWR9cIzRNT6PW+JL
Wsrh7Dy94kC9yC2bLHOA9zHZSJxIDd59C5FbcLMtFkH0FRkW8AL1Y0HoX3MQUFps
a0AKz89axnQsUi/YV/Xmw9dJ7T0tIec9ONRbakdfpyzy8mhfvbZJ4VF7KVbDGfvW
LOyVN6xCusvdsAayIU2fnu2PLXWcXCu123lZNsQ4EAP9tHO7SPoUHgPVUuzfWz9O
g5YQ+Vuq12EbqGCFCqCKUHpDZy43ND7wYtghcPLeiqTYjiRAqKgA/AhPAmUNwY4v
7gYHIwrv8t7dzBV5B8iyFawTONU1AhgdFrL7YFOBc5PjElTRz7FWiSOxxRjuTGUJ
QuX19ewSqJ1JzHJnA1GIaCgmP+NIwpmzN+9/90V1urASGcBwoHVabrn8Ig7Il1eA
ObfeOTrOAA7SLGgZ4XXqSsMP8jzYJ2cALsVzgPXMBMf/t2cekFMiNh5Ghi5jEu0z
7BVVzbYsj35TwoDaFI8TKSL85kY+QTFepphS6YRSHW3CkZ0Zcwo7zfLp1GTLZXIk
Brq1uckMvBoUDcWGGb7M5MgIkXBxbmsYryk7B9cjvRJ7AxTN16BF7VmRyrlVZcET
ugp2cRXT7LtY3bGgBwc8QrYWnInICGM/Jcbf/Cp+9voCricMX5ARK8Ef7bT2DTrp
r4TXQ3MdmJxYxduyFPLDxcsQ+K+Y7jbHksViBAkyO6cyYoQeEum8i256XmqDV60h
Ud1bbKMmBDPimuPX1mgPw9r2kqkvscMhLqeDFK9NOpAXI3YW2J5ZC0qMkZwH30uu
bmM6qu/jVIyvpxvNtcOU9E7WrZCUfhf3pzvGVbfSKPoNcZ2OheJqtHHPjcO546gn
q14kNIu3biFy7dhFbTcBFWIiw1EOTp/1lUAHr9uSeSoQTPoU1WAL/+gl9rdriofw
MsSUUiY0UWf7axB/UnonWAl4nAYD+luEN/g3+HgNur1nGTiiEahYPCX8jKO+hs+x
GXb0asvKwA+XS3+Q9nsZbpieooqF6e88oO3anlArTkVEF/MBYAejE6B+d4eK+u9r
r1HJYOCAybgmipgI6TwDRkWEWDJRUTuH/FpEuFh3xSYWSwRd2+hxypVbHKIJWlQW
IVBL2jusnApz9CLYQJQNILGgy8/KkXINVejVFLGHjNPVulEz5Xh1x7jYSG5k0fn2
ibpGroLDeN5tCMYENLzdQzkY1irlnKkk8K1I7QnA629AbGtbK+N2i3yEHnJ3fW3G
EKYG7UPeUWj6DSOQSaVKh/m1NNr4LNjDNfVadx32fNUDb33yeCZjKcQMEYKNGHRy
axDL6HwkS5xkZTbt1NgpKY9JUxDv7IPTA0SySjbnMNtIzy+p2ESc0nEL62EYIj3h
GiQK6uX6PoaEqbQTIMY7fl3X9tg58C4tySxyhwDmZARxLWI5hHUvKUu/fWd5qso3
omUZJt4pZ+a1yzdNS8RZZzyMBlyo0Rmupv/UkXxIp1b0GHLxX9FGTyn/xmsqMSFW
Sg4fF2qdyaTFdkjdXddN9h/sxY9otHfTMjQRyQbSVBM4PTvofGH6/RBMFa/A/tUK
5jkHPlwxa1uLdzC9Mv/+5aYYhDtsrvfly8BdCMHobkjeWSmHx6c4yLSj2ImdTFBu
yTATM5LPOjhAXTfdW3CgnIWqVW+v0Pkfqz8m0qP1F0y8G0dBaLupAvOrQvwXitKJ
ndwRzYI6IbbLtuECug36x3FXZOiOkfvL2gQOJU83KNG/xQ0hgEEcTGxY58Uk29ie
hjtyqWdCTL7trbHQEUdOMXUXTz5RIdxG7IVVc1aqtffQKU5TLOqCBfz7v4VQaaoY
6gA2qzrWJojbtIUzlSH7F6HYc2fcp9OvRAWVxonvDIAOazEbhvQLVWLFBlhibZGD
d5m/2WNDo4B/8LK7cRCJL1QVzL4AL0kruximMG+dM+SGCFDexayb//bGy8Fx6X9m
KuFEUCyLQ5v6+5NAzZOt8FlQFIdv1LxqdavxyZU11qjqeiY5xX2Dz5ew2iaJeyh7
vCLc7iYl1lKu6Zm15tSHXep4M1n4kQLN2HKJTd8bXT4qPBoX+ArUTXzO6uc9GsNR
QHHWTbd6YmkKIHeVpKvejHMjYrYMlJo+doxbO+BpBS1n3DbZC/r1dnCNR4eILfph
Ql3MF7rnjbQULTIuvFpD86e4o97a798s6PDtdPWnvEDDYWepA2xU+l4xHqAyZetq
/be60oUtQ/PeKTiVjQbZ+DjaUbGYAzKCurGYmOBzoan+HbomAmw+AjnAmVJfPOjS
Nk//eTupNUDr+snVN4QHI+1qYsYBwCkzd4x6ju/vgDiS2eMGPmXQ+pvJx0OHvIzy
lhaqyIDRZ6D9mDJjBdfJQeTo9DXoaA4NUShiZUehodJwst5OUEecYk1UTgHboS03
bNQr5NdgYgf4SYbBeYg5x+HctNCBEY8P7qOnQXYyxr4se+PGyS70yC7pnTzA0My3
qGje2dfBIiNNjd7hJb4IYMpCaTzZ3QPrjZKBbsFQYQO9vdY8uiyDkFLRLBRkZ3gl
6HBNwJxpoom2Yik2Gtf6E2Jdl4RZ5yIH1TvXtBRd3SCQD5DbAq8hQ78Glee+1REJ
s0Sj3+u15+bnO1wKI/K93054ia960NGj5jBafS7U+hkh/z2Nosf6/DkAAill68jN
2hgRaKI9hvt0gPA6H0C2SsP0PlOoOamjBgi8C2wSiRwFytoUeqjTL6s+GbIee7xJ
rEE4JBferOePrjOZoWmGT4zDTaoGLhbsIOP6ADig11zK8eqawm3y/OtRfwblnWY8
XADls65AZmygJczFmjHBKpBluA0t6gCuSIP8g43ed+D6KiDEH9bYXqBFoVXDNM2V
MQsG7/jauZDvWxHCKWzTuSUKfeFKq/rzC+cAMxTXVrhHxDTOKQ7kfO90l/2VW+fc
ONJ+0T8NvFN9eFNxJ+Nrmbi4Y/laoVQes4i3jgVL7C8R3jjAxWIiKJz/8+jlM/dR
TUXhLQLsrpgJK79bs/KbTn+dP503Q90n5ZItF/JM0J0AcSBViXaFQGezajjKWO71
Inf39+A/dhbDPQVv8/ADcQfHhyDetUwcpytxEOvmNbzeUogmTja4Cz3f5fRsNaRd
x8UJMKMduRJNOo9XktFrWVkcvMxj/Usqy4zMEGtS6iK5XBuuKDNMa8vfsRBWMAWh
5WeKu4R3RzFOs2YO0RRrrMNalpoTygQCjZked7tnocmPZ5JJSsOQWdy8ZDCxvO48
Rds1hkcSqaklL3WO261pEEJWfhlb+c/GZIooM7XZQ0TUOhcb+/mHIBJ5x8Bz4G2h
ReU7vx/o0vWE4GgA/YPSBidt8qb5ypX+whH5568FY8XTb3D59nVJhFQ7yOLZ0Fcy
ByX3VEMzqMZFpUE+V8p7oFfyvRas3/PU7r74xEK+65AxvLpx9fmf4T5k4G6FGnkn
zbsAYsyVohYvlGxTfkuuxKoSVY3LgltNoLWtbcWZVZXw6l5upsn8R+10IhKs3O/t
sNL3G7PpgZdsOWJx2hEiuoBkZiwaOSLJq/CG1TV1PVslgU2bft7pISWm1nfjnVNC
Bg4U92cBeP9Mo3sCV7+9MNfas8d9bMTtzozaH9Scr0yuNxqV050gS19YE3Fm4WwN
Pg1O8M3yyFmC2zlhPWnai8743FPKWg5Q7+onjKoS5AtyJ5m15RLcRd0kbLqpGlYr
t8RXSZezptekXtLnJNCYnM3/QDqykdReSFgeGLws9MEvsTz0Igi8H1cHl0CJWkIB
Uv2LOB8wD+4SFpUDzJoI8FP0wUSH0wVFwcDrBoGIh97nwlZ8JurdeBpUfJ0bMNsc
NEYJnCwyeOzUkOIDHBn0iBdVF9k05/M5snruTDL+YDbrPAOm8sQ8eWTnC1QNhHBs
VYMDPYG0YVhXy83iuKIsK0bSfpD+lNqcrn8wstA2NXmLZhhPrl/70HvP9xojRxWB
woFw4k5B6qika2EfzdDBlWxjItV163LLSZoV5ejNhmPvhEBvU4clAb9dNqz4IrRh
7Fk7bliZJ3aOWdhNgUeO9EN0AypbCttafjvkN6Gnq3JrWSWPWCt4Nl9K7af+8pXc
HGvQkTnW8k/HgJWzKYK/9MuvdOwV4VoImd0BccxIkH+Gpn7XRyLz96bVKL0CF3aj
xNfN9FRra1TdyFEi87jY64hQbXbj/gN4xN7kUEc1I4t8QQAkyZatL5W6yRQGMGR6
ZCRbduhoUiixMrgqYAPblWnLvwuzO3k9iZiR6cH0SLsEj1PkZ69aVRP1W3fHkPIi
VO9pkB7IHeltg6A1WeinAuZ7nSHPKJiYa/IFsymLkA0p2EzomYuXWD4RcZ79et1k
1d/bbuUfYxMDiivmAXIYP1iE7c+utPjGD1d+pGAntSOQC++e3SjcOoybVNazS1tQ
Ke06XjyGGJWjwIGC5dkFuQ97oyXufQLy81c6NrtYS8AyQC+E0p+RILsa6gttf9vr
vTVO2n24GQ2sjUM8rQQkiIkI2MVI7nnKMG9WfFSkYPbIOkSInJqpSOaUyUZIjNiZ
Oj92+bhNrMaAitYEAWrcrBNuCpl8kVfcq9j7k5n7/BCw/m11fCgt1kVrmSqH3KPH
QfIao8WG4Dfv3I+ASWW806Ju+uzbrmrT/ZNOGnZWmIIQk9I55E+Cd6XIzBsTaCIS
mzm9eMf7YF8aCTbwk0GzGvzfKt3ZMD1YKkpwV64y/ZYrEmjryksJmyLJLt1zH0/y
w/74R3E3lvMIck1yN/jrbHG9Dxqk0TpaVxAXLPeJKP1Fcr9Wu2Ya7CSXNBwdfMDv
QlpdTs+qu6aT/7SLOhs6izQjkoU4TDeyrCuoW6khB+2wz4gZn2xJ10kEZ5HJgX00
5xwozbk2J1ls9a8h2Pl7p3hCs5DbH0ElxuLhCdvUiUPU1whkl5+YL7feaskELz7u
nnNZlem3bA0agtwQlF4Ua92SY2Dh4ncy9aU188e17KmA7ab1gd/sH3E4kV6lyhKk
GK9ZqS0Lre74fFRr0PE3OPd1pIuZjp0+V1LmU1n75n75UOi0JVFOMvC5KKvP1e+E
xMqI2LoY/6H5L/ZKmtMs+SSP3tOJGlSRS+yfC5V5/LFicP8kXqigReGwu9nIKGPh
nyeJ2qDArSjKrCHJhwJhh20xxBw4fXU6LQ4DHxt7JvSzUi6orwi4+pBxu8VBcZb0
kdfMnhlL/LsU81NF6b6KpktClNUocdvil6UNIFUPiT+WDfgaum5DuogcTjUKGtsb
TAzMmuQIzIJR/NU1/K41NDAR3tbMFempjWaNNh7GcjHgtAI/oj4opPpFTpLr0hhf
kuz5hAV2B6qk77eDHoPOwY7xf0Ks4mu2gljltiU1IdKp4SELd6GU1p62zvx04HIz
HcV99nCSamYgbotjmtbRe3iWkVPZb54EvjPp0HHvPWyDLrzVNGiDwWh0B78R7XGh
DBbSyegNGXtUobwml9Y5sMgWgC1bU9mqARkzMGpL59xVDn4TUjdoeUzKXxLZSGEJ
xTgTA5L+rAUEnKaw7kGxveooUsqLPjrTByGqZhUWEerV83gHCF9K2d3dZLbh/lDt
kmfN57F4H7ojXIDp2Pa9cRZtVVeriOoy0juycarcfVtL04IY1Li4ElglWfdkn3FU
EdsJo5wmCLftDsekKZ0o13bJaVh1Xsf0+Yw45STfU2LXAbbiT/k91XnPcZS/AhpJ
AiQCr16alGeSoULUZINGiype4MOYXqg3YnXSVjm105BFkhqN+bY6uUNB38bXOANG
K2DNfiiDctV+5VjwQh3zAIO6kpynI3IOpfh96icOaTaQNcPOvThNXIQKXZxTsVdX
ymobBEJ9OJU9DLJen6v+/kuDX7ef3pfwAHp2LdZcqZH9K1kR0pKZGQKv0LBImnoq
MMbpO/W7ueKZXlj5UcdsOTCxAnjuYDAmLlDp6inl6mDcRki9bcVC/NnMgUzWa1wD
clPRZCtE690mLjR1/e1xiOE0J1NhmEcLMgaa2COoVwsBwGgAsOqOIP6I/OvRwHT/
GEKf9tPutRuQn9BcinxRgSH3hR657kbA7jRgESVHDHF/03Hibi6cxtEDZRINZiv5
Fc4wALA+Ac1Qtb6d2OqyxXsPMvzxdx8Vlv2H+wD2cmbKrgE72NuFqjPWZtdg/KU/
TbKN3uQsh4IgirAw4BF3JMATTf4DsTtQQ95+c/lpqPGGr1iGjcVhr5sfbL5hP2UR
jk/r35eg2wXwRJRWqcZKFqMFHpx6nifRFA+ledqkiMVY6KOGe06Vbi/LL2FvEblB
HGOLbdgZh4mh6cG6NlFEyKGcfM5Vkf9tl3w9u3Rpnbgf0j5KolJoHsmDsXv/VqOl
+v8zKtFsRzs0gbL/pNb5qQl7ajK42IUMV9QILr9BQylFJ6B/WN8q02U2wQ5bK1qv
yWcahNBTrzWVWYVUoIc9WHfHYZIzHlpKHR50IT2m9EKNZme8p6mxZlmrQC0ICqwj
EcQTUzdufKUq7arklnGEbLEPMwvombNzyaQulyudOqyETKGkSduFCmC7jCpmvs3q
Z7LQirFoylK1qVySwBNpmJ58TnHazu69yzWUDsXvcU3KNx+t4Md+PG0uerUYUyxV
mJpr1LuqBYGg3Q0XQvR9XF6vsa0l0dIvERyJcWYXs8LbBOTtBzzS/AR5KFt68qNR
0uZa6479r7P874g9EpeZnKJe/883vRBIIqKGglnQltfK3fJxkngdhMUBs5mDIRDM
+TX5kAGrcRE85ddYtHoNGFlUKLn/HPMCE78X1PWeL0NCRiCz73CPdrOCq2pBvjXw
MOm7BKFLwJN+vx1U9/Rqz6P83/MOQui/r66kFBDhqU7dZNWTenAMefs3mUxA3DPM
gPtPbnr+1gJ22BlyTS+GY5M+ITEIdnc6MDNEKs9LA84bBt+2Ybmw9kAaNmoIlz7Z
pkJYBwixyOT/76YLdILnl4uxUF4VuCOBq5qP/leOIrLLf4MfVFV9JPsM8Ab9jlj7
Wd7UQXSddMPHDvdBznlaFz6G835j509ycJxFxbGY2cQ+UV7OHI+to0JIau93+gPU
KWWb0GrvFK6EqI3h6ifIKhhooWfNtUe46RNMaSswzijB+pM+3bkO454xiajRFWWa
KOhud4ZDo058VCjmRCFf0g6ZeokMau3BBLFwHoJ2MCfHavaEizaNqn0vtaoYyvuf
9KMPumSxiH4LB7+GPwrwVBWj0dg4Ffn0qtvmuEcQGbmzYVBxfdXh/hAWg71dJwGn
Y5fwO4SFY8Lw5dHHIqeD6fLKQ12SHAz6a35lLx79dKyg7MbDdsltNNuBKpdVVNE0
3KpSKV6DP+h5RexT17+bVb/9UaU18nP81jFMou2sj2l8gRwVerUx/Y8N8Iy+cn0V
g37cZK7tB44wgapSEbvVXtTjvKEg0Zfif1X+WU8CjVkONo6c/TLsKmNdvyvgMK70
zxkFvTl5kWKxINhhFaOm7BYLxaxT7oskVmLsDjSB9jia13oTC9uqAkCWdDPIRPf3
Bx5OHdJ/Ei5CXk+njQ9Wx0xdCpHXNg16k2Zh43V5lOWIueKDExt28PKsiv78/Uas
cXQ2Jtim8ewK22lUdnq6rIDNTjOUbkkaZRwSUr6rLqgV/yxB2JmyfH6RwPDm2AD2
ewTMiZyE7evzIVcfoRiPmFmPsLA7RDv3JO8mY+bYgsntC+8+VvN1/CREGBnJvR6x
8poL6jvMxchlco1jX5fQA6hNG+e5iB/3bUgaDNNhazgLbLl2BelIMaIx25tZLChV
mDGzJiBhwdY66rjk+O9WYPSN+MVrFlQvvlMIPnUDHOvycN5WCFOh/IZOptq8mKIe
Ny12BA5HeLH0qRQ66pNbAqfPNt8oFylkAfW0OMI4q+VEK9LfLcw4gG843zurq+dw
3XLeqkit0ypdFhBT2bU4aERv+VCwwiwI8UhI5kmvP1Wi+IgSJ/J8e4QN4QGd2iNd
oZG4tw+xfqIxaeDbPuFB89BsWRS3SqTJg3VegzDjdNRkR+U91iVhPB7/SnGojDNV
54AN0x636EHTvBoFPtZm+2Gc05b+LCGahAWfQ2yq2NwC0bzfR1Fx3DlOoghwF82a
nRaidx7PSa97PRVrbyyNCIn5aQpumsuLJJnjFyLNrQw7iekkD7AkCmFzeNZp37nJ
SlmPQ+PVZH+s2MA+E6p7vALnM7GHY0iEPLcob2vLz6QSg2Yjlf6eQmtcNLqUDXXz
opBOXgZ/ZTDoLLW213zjKdzYVN9I9LP8PCdg2IkDd35EJ/g6k3pviVa7pNgJGPKg
IC3Id18/ObZ6fyvwbYC3P02gkz4QoO5W+XJmO/GGl1S2hSOP8pbd6rXJls25RWQ0
a8dcDaDZTQ2MTqQFulmUMN5TbHNSyWvv1+zievs8ELlIDeqb/eIV9E16IHB2Wj3R
0niT7pYcl8PNFqbkekRXNSXFJGjBjFmmWf/xs97WoeX1jEaYyWXOlvAJ0XdU19zM
Acvga94B8dtpiXGrARCl04+RpRCfxeR7r0dtYV9SE1uRo3xzytw0/CoyfthtQ2Mu
AWO6GF9xb9Z/3rKIYpm1eckOHAJ+4jliM3C0SLpnE18TcBsVFvy3HIDbixPYdu7S
MubbkEPvW0kmZJPhiYybHsE5mZIg3JX6kA5BZPS6XY8ig5WpeYtFl2zPsisnhyGL
4SCTswAiwlbCQy/ECyW1r0asc5wI097LaDfBbX8fbUG9C6KSoTeMP6Z/hA+1jxzR
BEk6pi9hSS+q08iIlYVuTU0j3sFccXS4evCIawqc7SPtQqDTwohv0ZlNaxXsiLEH
hK6v8JhjerUso2mqiezcgcO5ag/0lS/Pabe9o3rWZaGZvXrYkEPbPgUIrhmClgnL
cWltZRGZR+VDOkkls4Y2pw+dcqp1pGrdTlWyoubY7VfHZMz2/NNK21bHR6dGeJGP
8rd68W+uc3UhCv/fUqvs/R+D/eVxNIjB6Uz64BytyR7A8T0YsE4I2xeh2cWszluG
LVWDQn5L7kmKuz3gBgVN0uq35RQWAi5tLpopfzFPq/X2ppQQm591M0fLhCoIlfI1
GqRt7rDH1xxs70kLsSX89WMSwqZl1rn3OJ33pYJx/mVmxANjQDSHTQuVuiZuKmJb
E0NgXeFy69eDldmVNGZeRfZlv/zcakshe3lrMdQ5VQQv9ynPzNZBTaUw3felCTpu
6qx/9vSqN7y85KoaWW1dDVVbgY0SMrqqAHsd6IqunwzGKKlBLSfpNyRcC7nKSlPM
Eax74XZjAcqdxmC5jUYyQBCEBRgENmRGV+dY4G2pFImFbG/KVl1BUY1XWnj9x1gb
42WQY5gDHEY/yTo7Xkn9vdJGyOPlKrq1zUEs8fD1E66oETqiHGzU/0+YCjP0u3gk
3L6m7L2324X21l4ISL/xPfwBpEvLsC4xTQjYXx4Jg29QIIiMirrIRQOP2DkPQQ6C
EiLQqW/Di+50H1+1nccuhm0zvbIFTpD81++ZnYMAzA9gZHdtPNR3ES/kF1SPWcfi
G/GabmpApj7wxvl8gzN7yaA5jijlOVhgpBfbWSTUHgMIqWoacKaRxxrFc+m3av4c
PshYqOxe6FN3mwPNmkZ344A9ZVdOc/TdlnyhoTRs/89gR6myJqvz+UkUasCqwaEq
zq2nIBuuJ4icAi/tLFUFNphjSoiwAGXINp4ZbARdwQuFRSzL8Gx9OKbLXARvzxPr
3q+Xj8zvbZFBqvnbppjxtsyRU2caKil7I6ocgerW0vgzaweotxpFBiAbCT7fqrNI
7yN5m1W2Vt8n73chffsgOFyroSuCL8Sqk/9G8byQA/zULtI68W3qIiD/ALVYg4yk
V708Fr4M+6srVHRL10SPvAIeEo73cH3ERopn2Xm8y5n+kjv18tX7hEQ2FmKyjsYm
J7IEdP4k8mmukEmJ/1RvjF3FjHhEv5dxlHPVv+CDjpb3oO/2LR4K9tCLOEApSxIH
zKugfygn8mMjd31vmmG+SwqnnoLpqrgYPpOsAUKRLRFwfI8DFKJZAUpXvMV+qBs3
dEgRieotHNdsQEl72ULdXDtAKWHgsB7LVkSaM/QfaNtPfDsoy0PuFvWIgBoJv99+
MYcUsWmcXq73kvuuk4VzH5BLunkF31cphIHYO6VJjTP8SJxKBhPpT6d070/Za8HW
0OjVFPnyDIM3bqqrMwJ2o1bOcmdXqdlAFTfajszj5AGYTEbGcaLKcgj0lsbn6f6G
+YUOEwVtwwYom0iuPt4efMWiT/9SwsL9FsuY34OXgq7nS63XwWRJb5k2R6zzMwFc
qOsxvPZFDaZ7TA9xXtsh8RmaRC20UjFwfS9P/PvqiAZzT8TF0GgV8HPcFy1A8lQO
u2XIm1jueqdj8i33ikEcAkIn6eoOlT8Vbfqk3uCAjCM6mClt+f1KFQ8fFmIOPCLm
HPGQIXOvxBW5osK+V2HdL477USHUIl3pmYr4K3vjhfPVoV6p1anakrDTwolvwXYL
BkLexZ+PaLGQg1u1Fw3vpfeDr2hQLcuhijW5Q6ddgX2+euGlHU4a+zayj2Bidjwd
/XhJMsV3lFhObl6T6MdniLTQMIPZrrnqMh3ldn1L1a79MWU1xic18LsGVSWVXUMz
w//vg1V/e3ee5G1aWpNMnymDBH/7JCNv1rpevomm8+eZFeRK62mXRMe2eV1kxSCj
xsxlTjV1LV4XSf8+voa/3gmojsdDnHEnpE17xIYbXWEDB3GhY+Z8nCb0N9JlzTD6
D52cymHAIFsejIgYd8yQDymYf+I8H63WreBk7HILti2gp4fnP5ltSDE1z7gAq07/
gz202oFhuA4Wp5T5wRcgjAy3TgrLAQCS71jWPUPDL5uk8+X8rreszRVHctfrq5P3
9rAl5lFsuVcHP/P8ecNNijXyrr/JOOt8VYY7kdoT0hiKqGsYsmP5mr94AEvNtiEp
0EgmyYGXIhFsEtVeT4jl/D9D9mbnmVwN53h/LUBclTrsf1p671aBQGN6H4d5RZnm
rTatg2rcnbJ7d0t78C8yKXhyTZKO6E0A/LRrLYh6B/fkSwNPwdggsgdOx8tf4h5e
fZT8Nm7zNvn+sKqyXx1RfnfzOr9opf/c4rN5sbtjDwjHTUkpepRC0crOLy+kyIRm
GOMgIpGC4NJ2fHGnkTVnIAPycE5BQQmpeiECoey3O7oSLVjAnTottb1+XAEKew0m
K5j8LoBcJwQpd5HRfdcUFC16GaMT8wdsq05kV5KSMQZVjT4+SqlUQd7jEHmh/Zmb
IblL10A6RnZGFw7NDtHjoskDwBMELGaMcih9PAVfTJk2FDVwi6fLZyeZdO/Uj5bJ
l6SOooONdYakqnMvkfPNRZCGneMAZDdfG/8oo0WozkSTjWMPLr/3G/e2h7qQ39zs
eZXodOxU5pcLTzT17RaDzU791U+qO+JwUqee/Doa59jTyOABxkiDtiyb1IePq8ay
aRZKl8Gz40USas+O1SYQza7LgSJj/WzzwyGvWsgH1VFmpAdnI9/FwlKomm2AaWN0
Ei7tJRCCZ/P2JhDxc48tFPZpq8Jsx8+xhtsuf4oSObHHYnLSxCcPNGczpH8b/0RA
DdZjUW9BKSG7VQ1czpFVJqmVLSZTVvvvkiQQg0Mg7uMfQXRhtdWTe4PgG1lZ/uKt
9PqRZaiDDhAmenxnv++bkue3+P7CRFeK4No9isiiOfu7eVdt3H4/E07X6rBaMXJp
fdH/Mpj4/B0npnxKBqVJ6psy4UXEaqcWnhXU6rfiMRswGqnoirDrChX7FAn6cKIS
92lFiyM3r+9i3EoIZUZGfAzX1J5mlUQr+j+U9rhNDPk3xwrN5c/URxPJ/8ae1Bgi
Uu9uc83UaO4KRTvSXhYB764YtG8c+1q0A0KNGl557aexqcTZT3FpfE6K0VXEJ5pv
va/dL7yati2ulUKOb753R/xBZKwuTkB4/E6P+ebPgMAoOYSVxwKiOsH4bk0I+SGT
upGRqRC9+dqGptn1MWgl0dA93dI1II9LzkM0lbfXZhNk3bfA1CqTaOYRQife1LjU
eWZLLiSYbGddJDk8TK8guhB1KmwhUCvEAexBppcRc+KGY3dc/G5z1LXUUsJ6RzAu
CpanUpBVQ4QewtdbNJ1epvSKcxqNnzVGDDgFxVKDdsy42vXDYfBkUg9+ol2IHPuf
orsKacV1WVoAgIg2lYRAXcNzCPaioTSLgSuqiXws4+te5SKXaRND3u4S+JNcopbr
qW4RIclUJL2GQ2HjVwTufdSjvW95/qS+U0rxPl0ZJqOUV22n1aFChldKTygKSLBx
OG4snDZJI4a/5BlTuLV2QsZLonMjpFYZUbu36PBi+xlqr/TqIcWC0L84DhiAYu/D
JtcbFj56SzJwQZAMkbbn/8qnPyBo6lXfSoGwHv/FmY4bit12UDaLF+mOmXSFT4Q5
h5varXiuWDgCZm5JPkuzwmmM0NFgOi1iGzDbv14zOgpf9elMtf/2AfcCbmJyu8B8
+MQEGrourmh8wMo48lRFHxk5SrmIWixx7W6l1Ob+GjTd6aGIlrslHmU01YoOT+9D
X9zRotnp/UYwpPJdRuSmP+bfJIUEc0bmAiu6E5bXwBVmNGmIrDeG+mrZer2jIcDY
LU5CjypiGx0gmTnLR1Omuj5wJGzsAdmKyE/yH9czWs1aAnwGfgL5vL73x6o3PI2s
9Q0b1xy1bSBFpaN7jVmyhHhnaNQwN9gNX+bj3hxAsL9TnQjh1QBuaBwByG2VTHIt
dK6VHa8WwTAP5JRCy6Bw3rzdaup29G9EtrzfT8y/YgxZ2+Cw+dizLZcD5peaXdCm
TybsS26qgmifKIM5mtib6bqnIfbA+RaW1ihMIbUr5LkOV486ft4CmYeVqzrIYqsS
lt/Fbqtskq6m1d1VDI1a+Oo7aDB5qGDLmvNBYvR/SkDrxjGLeteIuXMpnIFby1hK
puM3GXF2ZbtXHLNL7bLWZ/u8Ka0oeYh3D8ZSGihUYFwo+lVIuHFNxx1ACScAcVWr
Dzp32YJ3wYZctqV05QdESgkWmAKS5CNGdt0mng6SeJWL50bpprLXjT9Kp6TxXakb
WKNhz6cOATRVUIO6i1zZ874S2vlCAUt00hRL3J28KygB1odtyzDl6rwAPdfGPqA3
wkqiEGP1XTefoxJi3z3I7kx2WVLRnZlJCt28EbAQLeFsLqizxFZp2DAGv8tB99yZ
eblaZ7dLeDfo4j6xmAaHw20ztXxQHM4N7Q3+n+hJugI5H5UY7qmlCbAJK9pQefrC
s+H3nqewP9nxWflsKyi15EgvvVem53evsszK+uZrKM7/5gZiBuoTvdNhbbM6VuET
tMnAR7cmeaB0uSgwj0n8b79wuvmovKwmJHP1FC4amMx0y6PXNdv/4dMoNVwL5LKp
jPGtRt/zWrZxBnXDKSQlxq2BJvKuu6jaF6oph/TufJmK+9tsE7YTEiZP7yJGgO0d
zw8KqAtkIZjWpfrVEjqZ1KxqMEVFe1xafeDjs2cxCXoZr/dOgrD9XsUuD1g04FE4
n8I6vQLm36q9cC7L4ibIVCcamodLQ9RmPHHzrZT7Yl3CsPx3vI6GfEXcU6FmX7ce
W1ZMgRWYNPXsRWknY6uCys1AMhUwu8Z2q8aNTvgqG5j1WmCDAiuqKiuvkZjbt99x
wCbghNcKm/b8cPNX47aiZnadh/DfEGl+tsghz7pE3G/hFcUYZRAqvh9y4SNbV+fT
mrUp87gvqw9hPWS764TPy8Ghmb708q+4zFAVdJP17tgwp1ovYNBhUEmkeTZ8wz5E
3FSdEVo1Z1jq0yY+C2+Y8rSI7s9xFpVImHC/0ldO8RKEZ/BsZ3MqM2juD/ctEGvI
U1z3Qc2mVCIZo9WuoZQH9QZJMBybXuC/EMiEfRy/K/TyFvoOlZRmPfg4kcQEm8Dx
qL1UQsQZoMS8dtsffEy1enBb1PQUbrQHho56SlU7WbmmWd2mHn7+YIMhciyMPX9T
rKnBtphs+XZEC1xz4KXwY7rZ94u6JSDvIg8VFt2CrTVG1aY/s2PcALd6tZUn7AS7
Rz8Hpa2TFRJJggKuGqp09BvKKYnvS8+9zfL7oTbPda9EiwfrPCoP7/9WsXkuLlGh
tWg9GbUq/VGmIIu7XzQapb7PAEiEucEYlYvM6a0xXYvxl78BQoH9PuvQwHQM2Vee
eXq78hbPwWFEgBx/loqOGEkPyrFqj3TcwNgixcA9psIXm3Jlwn2pf/8pzzUTCQDy
hgfuwR/E74unFfB+s5uXB/Xc7rFMBVG5axFxHhhEivsdzJzKAyCAB/ZLVUVriQNS
U57LycmGV1n84pAIR9vyr80llcH5uP1ZpOslgtrGdcrBaOdgFwtovlkSuslZrFWS
HBP/sOrWkxbnv07G/F1pg7mNCgSpWrefIRJm3hLtQCq2w6isVYvjbu385Va97Izp
/2MvKrHuSA3ZGPCuZ59K12AqFsNLkT8FTRrCCxR8FtlNN6gzy1tZg+iwvGfIySVs
bILvGYeALo3k1aovJYxxtzBJyN/CmZ3si6WW3t5u08jgmOVcFnx9I6P8rSMUcSC0
yI9jDGytPqfAtKxFK3PZ6c43DufCfXd4asu1fQHVHJoAFuErgHkXSgBatp6/aH4z
wWeXgtOe7XY8li/WrygBZUkn818SaDdAWpzQpSnyVFEbRFA6wlJlakJkQ2GJgzCW
39xy/LzI/tsQRWg/UIAnfpKzxGTNaGge7oF4rTjddn0Mfk3B55azROa+Y1+XMFJg
eor7eojaXYecg/m7vzIXSVN1KMJm2P+l8VERR2mnA63Arh7uQqaiztOsrIiwsfWN
hzOfU5DLIZM+MiGZOWrCTyNCK1BDlu13XqRX7OkDp4mP8aj/cp8xtAEkUSYps1Mf
jqX/wkTfDB/aMTEiwYsCTVTuwe+Ildpv3BF0MYNOPchm/vSWjpXgc4cBZlttGZ1Z
OJPPgXu4BSTFJQPws6Fv17feJPcGS6hr2MT8I+hl2X0gctEtm65L1SIFtxchiVgv
rEG0TTtidpVGpK833npFtN2EAxSt58Ou8vYxYoHYEnmAignWO2iV9vyCtKMTw+lN
AyWU6ct9wFlzuJmgGRDm65TtB6TCID9Pso5jXp7zu15dmOeD+q+r1e8SRyFuLv1T
ij11EN+xflAtL06NlxNZL9yz67VO6nR4/dtcHTLnZKLDOOP7kiu/z38yDHJLbFVu
R+ffB/3cddgLQ5XR6W7muin12lERVqyhZN4VpV1K75pPlYbJiJRQ60775ndcl1tX
dArPCppdNB1xFQ9dwoYsvCQ2DbpuSUHo6100pghmmy0BAuy1rJGDaO6GlU1GIR5T
Ey0Ms2619rYmbVa1M+uRLVJscQb9ddbZ+SyIjUGR6ThVYEe6ydbTJfa+DihMZmJZ
2We7H6SxeAJZ9pmB0EMTj/lf5vJw5PMcqfnPSqGTRXJPUH0/jLoUQ+Hw+rul3O9Z
fc2TSgJfA3v6eVwakaQR31fJfdDTkUbcj4VmYPo5REgXBQU4gMV8KGMd4aQ9z1x9
enwbZf86MsL6oRNRdSaJHWaaNVzoVYqS1ZJO+yQh0yv9Lt9yg2f5qaYVQYWaMjvZ
TmrVR0aDBKeShny0ojUFdLSkto4NFLR1u+uGvlbivS8d3FBMKaFtCEKq5wg8Cbeg
apQjmgrNHdNBiOKL6VCazKBYff/1JfwUpaG95QyMkZj7dXmqb9NHtwHZHxdqP5P6
wL9F53SykTZVsNWVM+R1FZqbBETrOfNOKN0OpT8jlTOtYW5tZR4rrxyhp3xC1Sqw
k0HFxwjlcp7PkE038qEAJ/rvEWmF0pBhDKeO6xoKmDnJP1VB4Skt6em8PlRSXxkh
8gHb/KZ2REIQZf9LRotohrOWjJuv48cYw+oF0MkDw9Ee4d9B6dmWtja3Wm2Ey2Xy
+/qZIkR8sZ22JHX/uCdhJBsvS4kV4TI34NPqtL12YpmfL0/VTnPj6THKw9oc4SeR
OI1/emukUViKdZHYvWXxikAliBLljHIxJQWxn/BvCBzoBdXPSuAD19CtO0IAtNSR
x47Q4xQbWntLIcR32wDl/Z4oAIIDHM8hrDKlknc40/lLx7NWT8uKaJ+2kjoDr3sF
c/U1RQ69IzBXlK1SnuMrwjBq4/Ifh68TgMCSwbK1socW4vEZP2Dp7hcLPys5lgN8
O9fGIchffcg3ujdJYfivIm88Ivx1qBvrrQBfDUM5WUWJXwrlKv+jIG7eHIS3+CFu
f87C8lczoXr+BsWNdqHFiiERwUARZWF66lqCbHVZ+d6gheF8YOwuOQ4Pp3uILbQR
MmNoXtMOLleq/AN4SQexhpb53wRduOuVR/E62BrfjzyHj0288g9Mnl7BEjjfMsvb
sHSUn78KjELe+prtLOQLrDw2aUj7l75uRSIDDE/zGngqeaAO3OX636zf69NPeE0F
8zcNaixUWpqDKpt5IjM5DZvVuJ89eZzvEo8nrewViFciy06JZopUPVpiCmpFPXdl
na73p99qAzWmJpXWDcqtHdIY76ChGNfi7rqgE5fa5Mtn1tUik+BSR4EuoxSu4IA+
CEXestsy4yay/QlK+IrQr1p2Omov8RWbi0XOBoAkXBETuYjgObjTmE0ieVz0RxnF
My9bvH+/WxzL2NvMxkYxoGUMAlQvPxg3gRNvRZdlytKtSu/hrzg6imJTPuUychwm
mfPxLxO4tdV2TDsD1FytgwldQr7wanv9GF2jMRa7haue4MDMj833f5G7SVsM2FL1
g3gaJDlHdHneT1dbmJ1ajnnzr0t/UQVaTYygZ1ihmTNDiDiUIKxsN9i3VBPwF7O4
3ow8W3AOUIuD/LPUrCIxO2FKQUi/JGjrgnn7Z84pUkYt5QsAkxLqHOetGfIdoSbu
ZT5kPMZ5uhrDkh8i2hju4Lzt6aAOs7YNq8W2xZYbEQ66zwXWcMyaLtpJrTK1NtkT
cuoVweNvm2BBmld8ejCYg+qPw7WIWfQ7ja27fb4/DLIvZHSx2lL0oIyq4hPldjCm
631MTrAMJV3ELFFq0Fu8+ZfzN++fsessCRjPd8KKswnMVX6mNJHvNTFaJ4FVzNKK
67SpgzjN62AEyw9Nydw7kjC8KCh1LtvbGsYGBSZLMqqyGCUNxE/2KtTb/o757anM
uoz3up+OjDrdghJ9TygVQ22LJAHhRr1skRVAzTXA+nFUr7ZK4tBJhKP7psWrIzBI
u1DbdYewED0M8D8SQH89mkmkV0ELnfOVVJmdAcEOF3xvcJO558nZ3Uy61xUkByQa
G4gIoHGzB6+07LPrZn9d+ZNmdlMPWJ5a/GiAwQW6CE7Bjep5pcEx4ZbZNPIStvXf
pY2Fn5964hGc2m7AoVcbV62IwVaZD2e+kQytizkvY1SCcVGbvPF9PInzJKgUk9CU
u7ZOB1nEXkC7JdunDYHRfRnOwsktNWOnBNrnmSnyBJLgraa7z4bM+AQzEYIW6qQt
bQgi2cIO5AYtMoEoeJYuHeAHvssyH5hp5Nmhuj65K7fD0aky84VzYSQD6setU39C
zAeokJkMKrBT+Y9Pg2dcqs4qhKQ4V3geQ6rBWmKbNvIT3so+7kAUl1yhpkaL43EN
zphVwG075rZUYy4GEUJPRjWUoNWn3dkSnikKb6z55ufXt7Rv+AoQIT2mFUpvjF3J
B7UzLsPIgIi/HX/yj4iCh77ZX74cPw5Kfwj/kA75mz+gwE4wzOCtG5AyAfTlJCQH
Bqob+DgAcrl/umWrDZjknmBlqc+BdET/8proHUnDN6vxVT9ZpoGlx7vwWU3vcBJg
E4hn1kLHzHR2u7SJSQBxaTFriAiV/INUotprNntfv4Nckf1JE8yCipZuFq4L5mKJ
SikFTQVZ6P1odQMI2Fe9aM0oYjNZ2jaVIehlCD138YkTiEILz5sxh1uja92KpUF2
sEmbKbY3vWRZEs3G6F03hVOhnJrhyU5VaIkME8fU8RP831vXPKjZ31nRspN+g6tX
HCUCzw5LT1cXiy0v+2jtxBPRsNHBt0F/AsVvDrj5a4Rie8olVawSJCdvbZ9ntsOj
1R4bqd382arEqeWX58ZOUa2QHLPkWeTS71mQ2huBXZd8smUbSw9r5W0ilzvmVOIb
i5DY4TQj1PsD65txAqc92rER+XOqeqG30JsX1xf2xHhEiIcxW2KFsU6aWepF3+E5
3JsP6FdzOfO8iesg26rkzlFm25/hNJBjOe+uRrnQ0q9v71f5kgDS6Ih8OgkW3MBW
5KZr00Euo3S3+xt6RU1/a4S6UQWr0yrSWZJItZ5Wn1pjzfBA0uLt8C1mGvW1Ztot
8sfEzYzdzw5G9en2hcsLGlbFoZCqgV+UOL1vL8zIp8v9C5SNz2grxduThgThemqp
Oi9BTcPwYDM5IKTclFIQ1QlPvzayJqxnfKsB2s39PgxgmDu0BuiVMWitJhF56bkN
eFLxj7riOzbj2oHJy/M4c+ehFBPLlP5UJpO0jBdAcZbbyENeucLoYmQfDZT2UGRD
ao1/gtVSQbL6DtVOcQyFd+xmNdCBfuBkY3jTiTrjydUcaiuwmIVoOvVDj87o4kXb
I6YcvQXOT9/sfQJGV6gkAAprXGSyKEOkGP/unRntG5iUCIFVci1RCLhlCzqCtlNe
035HZDWPARlQeMm3WWFEMebxe1o/KETQuohI38VmQBLbchRKhEduA/j8M8LziY5/
1dzA6IC3cu1MZm2R0zvmrUeoE0fk/CyYwq9viyMYzbCRFqE3QKYoFeTpnJ/VBLhf
1Y/7XvwbelmH2RFcLnrq/lhuxLPJ1HDCbNzWbpqFP8vDLnFyMkgKmBYNvAjdQncp
rHAKSWxCcDOWooh7DsevErR/IDc4Fa3/iSUUN2mp6J2xjfYsIa5O9yBgveRsLo5h
VsUZ6luYqxDST8kkfK6rfR0WSRvXft3OmQUahwoHtVoZBB34d7Cy/TLt1VBtbiyb
AnzOB/toxRXzWLu1saW6DAs/0wROn1qWF5wWJ7PIo6pwcGXIDJDOVKKv0loReMnC
+Qc/ObC1pLCi4xXChU9viiO+hNdEZWt7ZwCWAz0R20wW8OeTldIO/G6PKzdWu00P
OAaDF4RJ81Rl1d+VGh9LQoODMCL8dhY1gGazMokbXwGk2vHEYxeqtUxhWlrI1XnI
Jlsazu/qZn52uCF/LCZYfv9TXEWIPL8XWEOm8UnHd4EWRdsXxB5gX8vi8Vj+jgv4
w0gdshp25zW1IBAIrApsiVyaZmawvb7zxlJM4REVyf9bi1h96eiPfOUq8eZX/7Ro
Muw8uEfPo3akTUpNPJJx0GZJmuTMNrplZCZK0HpQ7XvSic/24iN3H+4i2CFD9NZY
UNxAoqoM1VMG1fZhovgBNkGEXJcWRLosYnupSiI5Qtb8Zm+94jUwIw5FEfhR6J2/
uRBMr13x2fymh46Ec/pTXKe43HnpjE12TNoV4+uvt92M5rgBwBYb7y9ZX+WUQl2U
uaykEVStz6ahZqd8UMPn9aiwufmpO3YD+/2KYR3aiFqsOnJ8cbCu49mZnw0YaVKh
+kmX7stj8JcxAmDt6wfr1ffhbgP1qLkrsuNKMwODYOLWIZ576uu1lhuMg3hmUf1y
Ps2UniaWMLs6VRPjHw8CZ/UyDsmYSUyTVwBfYZDbOObDe0eko0iocHEA4g9zcxNF
GK64giwk+uGywLhGfdV3IEhnpj7poFU6CyyWdcfGO9UZOxmDDqp1aNztqeTLh+Gg
InFQcwelvxQN0fx4w79PBBXEpx0V3OOkvDkYw2w1+QgNDH8kR3DSGmCMUY428XUW
HmeRmwQzBbsxkYGaBUW/mTnVt77KZmfcWW4LScrjCuMZatRp2TzlquYmzFGq9wzP
rd1icU/A4N9A7P/8mQa0aLMjnlD7JsEW66VvnnMZ8AJZGBLVaA/sjX0fYJB/E8KS
4g6Cu4QA8hOS2YzEoyVYcqohLl1VyUQ19giqgAEHFZldEp/w+fJFPt84x6R59lhS
RypGd9eLxl02QJ1cglgaKVYnOwEmMU7bYBKxzm3BfFbqALBhjnWbNE900LmOftsN
9J8WWVk25L6EpFa8fe/3OC06Q/cBmJq26YldGGX1KNAcz03aGBd4qogQ44rzt6Cg
az7ODgwQmNtXrZ55TVhOIwk3fyGQup1UFqJXV1VbZ+vK8IF9DQq0dI/DNx5e3QOi
sjx93pSIeMvv45G1C8Zg0GBcurycRowSEQLgvuMgAg0RnF3sol82QekWLcEb+E9D
l4xZEb9ZbYTuOzfeaYjxoOF6o1cUqVGwgiQ1nw/ss5azUHUf5Z/A7rGultKPorP1
M82wwi6jQNhueVV90HzgwCj33PSQ1O67ryR7+zwM++x781fnFznUeS+EvB3XZXyy
dV55Lwjm7x0GzvkM/PCYrgj6u0dZK8sYOK3ZiMmBGy2OeOlO3HR955tfbRypgz96
Q9KCUzQHOTTIZoNPCyAdGIn4wp8+wk9gAkixfYxaIccXjXER8Q3bX5B7DMLxUetS
YatHOJCw4In6A81Wldl4wJGcEomqjigrKqBijNghdSKhagUE11ti5ngOML+zXLsb
gDmEYk5sKpQGvmmNPiarybDZGj0Wa7IchO9n16EqpWMo7OtuVvmsUFSatQCpOHTX
4wb1e+YchExy5OD37eBrk2k/f/I+W+xsF8akWechCHHFmUPLEn5fWi4AJ2V2Hamh
a6YJ+BuDfXUfkULzEhPDpGfCXehwChTBQMBCrZK+6L9gXolBwqgZPOH5kb8aL0cB
43o37kc1YKU/TyCXlgSwC5Xl+w1LGIMXH76gIDWaBP2fkDFTae4Q2lrmGAKZVmyH
qj68d95aKxGps3nzHL06Bskk5Qqzo1WPmfKfYhFrqWaWLmnOaMoFW6QXHlpkx9bF
KyKs1pGXqYlb74Xc1AcBb4+o/V/kGYDVwQL8iEGJKW0jUFp2P69ILozSK8hVUTOC
GiavlJ3w5ivVajMTPchI/ycjvNe+coYJhimB0akilIlyZdiMmnsj/VHbwrs8noiL
2wFTpUX44VZqdFey324zXDv89UpJo6M8ZBSOd7XEodT3CSIyKOUqrKMDVa0Mzn7Q
4+cHdiiIa8aLGuxcoajXX9MdFNw+JU1wXBrqbm+WP5Unq99wM764UyUCBZ5K6B+A
emRH+Z3WgaNTEukp/3uDuYcZfmyaf+cG2gjEMa0QVfEntV+DNZM7TU8akzq9zTb/
oN+B3wkAd4aIwW+KCtcOyVzfPqmHaph+ic/7NyOcROcGlGUjkU5QyywEaS0qq6Ot
Nl/DK8jlTpQIa/xG29dyClR/tzjTE7/XqEYtZEEm/obonaS8VqeGkBVb6VPC0d6+
e7QnSndxZbdCD7Qi3KzC26INOfLuOehN73PwkZAQOzcH5yCgk0qD482cblnzQ1qb
8PuKl8pQ/nir5p7GA7tYp1kR3e9WvOu2U6Y3VU/jHu6xKpwMZ9ctgUMOSV94Ix2D
/Kxmq5mzkQ9E9TLORJbwUB+uD3vNZ/KuVispEczPKcBVceQtnlgYKott+WMh8noY
4yCw8e+N90i9EN9OV2XrpgV1gt5wZ224MKULsTnGZ57vzeBTuXYdSDQMTzjJ2e2o
d3WTQJas285c+z1cwYSaiQdew2piGhi50Uj1mGQ2NIMUjR1aQ19xUzOMegNLhquS
4RMvW0lheC23ab7ywrzFh6kZ5FLDBIRK8ubToA7FhzfSWyf8rO9UDHZTn1XEcc7r
gD5WA7/wjCYHZWzsHVU9/LDGiS2eeOeRTo3W0Y/JwO0knodLmH6AIzAzJdAJB5fe
NpK1zcRS6MuR5J6q/kkWbMKZtP9qfFUiRXs69fYaRfkSi1zzcOULDYgdlMGC0vFz
kIdJ3OjZzeNpm8MEdKehOhk8cfNCAVDnmoSbIspa/ZxQPnufXWyhvj7/qoMfCo+T
hey7JGiV7NWPlJxQlzqY4ID8TdRvdeQQYgqnEG1aQ0Ry+R6uc92KbdhhquOb+2Z+
It6ffcDus51Xp4pkwrgQh8j8uX/qm5eItX6TQzdxRzeG8a7lN+Bo4GOOsYfvMYM5
u54jsd0N2jt7pvrHruG2BoZZwQiXmpACT9wXZJVaal6YbryiHTabbkUsKkdtpfJW
Id1amE4Xfrp6B44qYvXFJQuEF+8xcQhIUU+cJncG4NO0i7935NQgjira+fO622ZP
lsweYd58c98P9YWv2lzKtAsS4twLkOINuXfOscOx4+JkMCHploANmnK6YHe5REot
yOpOcnUBc94Jm8FG+yqXiFDi/XHf2hBChKarJtw1JiraKC7/AyiFXTIV5yn1kyYD
nvr+uyhD82QAVcYq5su97QGEOlvy0enZTXhsGKNltF6uQwoFUEmOYtBEfs5IMC74
TW757uPVyEt3Cney4KgoVSUKSWJYS5idKAf4TfkEG8/Fojey0EEyxR0rtKh1FfNh
0mdhNre9+j8syDxZguRNVb/sXZKdGD03rNYJ2SLPDMto2U7uU+mHv4CRRUkxfQXl
1Y/il/xzt+h43BK78+/vDmBh3uAfxb43sexVtt+wqzxh27OExJ4c2CI1ORUlPFjk
MARqesTaOHMSiypl7Fm3A951/YpwDr2A9/jWevX9hr2yV1drydfNFZN9TTsCJMRd
e+ZXIx/+ZY4OsJNlAoFjtIihNhWpL2oh4voPbRd48qJUWNb3np+SZrWnKr2bV5Yz
tHlyNgPsSa6C6VecYkbAulkMMwL31/EaUcVkU2OUURNTvZ8fDCKSqoVn69x9rhEK
fHZ06JtFPWUSB27fD0FSoTwrdQVyyUmMvpsRDCOIxagVXZXTX1LEtXiIUZ2yggUr
VI6OIQsP3nmCDojVGJjvKwTGkHq6OiVGM3fnOtsVmbefL+N+GEaavQ0mPvc2s5d2
IhyRi0ytiB6qrES6/BVW5dMet+Zij+23Gz/4nsUPx0CI8Qe23QOGHP5l5shJoC/3
7SWlT7LBIQY2CugkKlfzE5XBO4XJqLbPQGe+57CnljW8bVwm8Gyz6KOLEZwc94vD
TxGOYcUKRAY07UyB28PkJV+JCrNLLRKlnF37nXqlPMjgchU/NApTJakE0ekVakdA
x8rABhshvjoGqHCedMkUxXRGZGc9Ej2VEKHie5vZwWyN34/HIPdyixT/hTyd2HJw
CRa1q8xF0SXkB9QMFr92ti53tbnpRTBpF1EYLYDLk61KN1ouogMpIupdtQRXYrUp
3cgGGNs8AAVpUNL8dB1DuS0kvzgkg1SaPUyLNG91PUSJOdmBOVaB7lKoYcuXI1zr
mL/oYvhoWsG6670/YdxdT/4v2qymYFAoQVAzIC0i0lp200SIvHxsuf5DlJ3il/Dn
0NhwZD+7ft8slHoQlXy2Xmg21hS+ZpiridKCmYdOmx53rAei19POrlM2JAjv4UKX
gZIV9sYur/dD02puZzyXHDzwrlwkc94+loBqpEeEHSf0urhFr9ooyueoOv5ycH0f
3+rBxoYNVuMwoQxUAFaPAP0LxFOLswsxcGa0y2uFbUeHk6Oi56su3+dZ2+gM0FSC
XpnkFCP1SmDIZAk4rANYstY2OPypokWfX6HR0tVjU5E/Zq+JzPd8sFbUFmpIh/KI
M9Ria4OOUFy4YuSc/l89GmNxiXbboVEBvy1JzNIG7EKjzGlGSoXTsKEnzS2awrC9
pzOM6Nnjiz3VCPrmeB/mh8q2F50s8leNWVA35mTX/CEdbffTx8rP8JjCVg18RabI
ZRp7fCM2DPgW8bAcB76sDLQ7da7ux/qcEGlKRLqTFwGbEYE7xANhoL1MIfub2SZs
pNgKnObiCdTUKGGq/lrjp+B/T/xSv6J9iX7bZWXkvvqrGzJD1SH07dEYhc1tzKpY
EhzZfc9auDP8VdqOUOIUV3q7bd6kCJsQk+cvd6FJ/yuR8+grS5QVQsnGOEUQBrHA
q3ISOV77nTJnpLhF0Lh8QtooRHivyjOIwBhSlcRMINEjWynlvVKdKXSBjKRIbVGK
Ad7EfQYRs2T3D+LHiUUNAToeqr7JLIYWneY01VfWMP2DcSrcJ0T8wl7SSW87SNma
NMflRQIW5EOrXHV1OD4gjXh2EMndcI9HhppmPQVOBLuHCUkfs8HGaK5UisI4Kgl1
Sf5OcopWIXFC3Fb+l29t+D8KoTlTBfcBlcFYxioWbubyms5bhb/mdIK4lyKyyj3B
bME/S8GxIdZr8KinUu2V+R8uqUAx2K0T3j+kVPZRmSxuuY6uCXPMiRB3LyJ6CyXQ
kRPkrCd8dU83TjSdZncZ8m0z249YItIiYytWox3xsUKuRoa/TrMyCaS8ysjJ/Uze
QBTVibMZ5cixjeWZPQgPjgLYz3RBdjDSBzcAzH6WEqBBCbe5GtmkYRnG0cRJ97zI
N1HZhjS4JovLVxY/XsWQNJN+H8JAw3zTHwYWfsTOTVF1676UG4o/tNuGoxTv/mYC
EJsHQoxs4WleO06Mu39mbFS4WNn/fjwOK8SsPQ4MaJBswHS0DBQbyVHEdwkhFbmd
QfHBZC0xCc30T6dtOa6PhYJvCfE+35GIAG4eGJmZYoCVx+bLDwwfKEh3OhGI5DBC
C0F15jgtMiiBtT7izpSlizQv4otKPg2qMZoXSx1Osp/hGM6c6i1Y3dty06vf8JzZ
ZdQZKzHgznQTwjzaxUChhjFS903o7QkLtAVXpX1AT4k01cGyipCpODg99/Pc1Snf
3u4/2dFdnBYRsWNxLkT2Ox4/y79wXh+jgaHTxsIes/LMlJp+ejHzG67oMXwsdMr+
Q8ETYmShG93m2kJgqbzJPnptRVC+ZghTPNBWeH/qBSrkH0zf5Lz8RdVTY5de36zW
+GNpkFNwFQY/XnRa6p4Y/r9Z+RtrdgJzFBpqaH9CnU4rVp6b4cjsKGd/6jVEEPCE
tAhYPZH0j2nuHQAOf+ljZJ8XSfcLGLlYwnLzfGYAfw5Me7u/vfVOi64qBEnt+lek
Y5sFnp0MYcDGtzRta5Hi1NUlTA3CDBS5erTTAja9rtGDk5TyxjY0wycG6WSYVWxy
qOEwgYcGQOWLqu3SIhBCBPoN7Gk8p0rADB1z9gPbMOgAAzwB56wHvDOJUAvFUga3
TdS8Ln8JMBnOZyi13QdkH14lmufK5AXSlgUBl6q35rDU/ytLFznzwjVvg3yGFuNi
KFOBe/tI7oOc+pKrnuDNq8iQlOw3lksLUKSmSiXeBRvCjbgqAdo2UbBIgw9Jfixq
OrTVAuvoJlrAfTnDXt4m/gc0DiGl5l/zptvfKB0jrXfIk4cZrHnC3lDkojgEEpyn
Xo6ZnxLe8FcteoLLJ8unP84rKI9dC1+iTGEVp+W5IYbjaGRq0sa5UlHpQTr01Tcw
2vS8yRp4h7csCIRRUrZKvLb8vsGnL8YPpKvxdcHmJyJmbfzew4BRy4hBflEv5hYa
jYFxrVRgfHQ9wHBMUdRptfFcSkJZEB8kpDxxMCwNduUEmT63lbpERhJd59HOZxgQ
42EfXTJQmigJ+mbqHfC/wpHdlmsIUU+LAqFAzhRz4XJhIA+YYFeasqGBltcebzdV
xd4HnoFhRP5gCpvO4KahodpR0fhlvVaTFgsei4bgBdnlV0mvkvMROf2dQYBC154l
WRdGo7qub0OKEF2K3wG5W0GG11QyYtJ4g9tsRbPsBb2rtg7WV6GIlYFotPFu5Yks
kyE9L2ryGRqW5XRClioDL4Bh9sAa9vpMAiChu2QqDZiVQBW4PwQgOtM//cSOj82u
7JXIseFOACTksEt6Uq561ylJl3Q3mlZ64O3PCS7dGVcIwTR5nCzU0XSXzPpxN1tt
suQ1CwNNZofKBdi5FancPblJZa5L86Kzg25Dqncse09o98M0R72oQNd1rSNAb7uT
rwrg/OQSKzybJ1ksB8+PKuprtI2f6kD43P9j2oB/L/nxo3o21z/4nOuoS5vnHFqa
U3iE2QMMIkn/oMpgzko4aI/XvaWvA7qneLMGh/lWwAyoG8gKWyfZ221U5csKQRXT
57etK5O2JCUb39+cxJ8hI+tdOeTLkfsSzX23NMBeFI24LPkA/ZOgxJomIGYAZ32y
0hlH33KsM1IPBEQqSazuLb1o78gDTA/G8lUZbkBEzReVlwib3fMGEzQxjKSRy+4v
ZT4Y+G1AIYPFcP5rNzs11HtRX/XxlBmommnuHEcgJTvwVNEQwWqMMpSFqRBVCepj
3aWiAV4MUuarQ1oC/3dRWzD5/AIJIEM3Y33oOKYpw1eerpTmHsdEo6ZVP/E0UBRp
AGEBCwGhCbEtpdVUBtmGNe95Ug6Z7CsfDJExIaal7n/xtAyZwRvmCSoGmlii5WAK
N7k6nA68lCtdpyAYKYorqrhR+pD4Np9zzQxdNrTn9doBJpFmOmT+w/qbDhF1SoTs
j7DfAQOT95EQpU+rZV8vlMofecaAJUYVEfE88leDn/p+CxdzvIrMKevyqtMPVV/N
9HZyHKHN3b7p6H+wyTHSpYu+XI2dLyE/LHiprBFCJ7z88+EecHnIRny1+FH40tGd
0esCCZ+XYglLtUKipDUS312B7A91CSpArCbnJv6OoBFh3EYEjQrST7NbhLSUt/or
WbR7pwalK/f9aDGwwjTjlirRZVuaFrL0JHNt+b9LfOZWeccB1OavZgt652pg0NDp
m0ec5Y4gunoCPvC9XteYlzoiYm5EOLZAT9AmMmaWIEDyNbMILDbXvJMeHNVOle5h
Xqs+DlFgTSRnRBbibm3tEKXN7JNTlHlVUuD1Q8KxUQbA9JFyM5RtBhXHkIyOk5z4
i2/7DOioDh+bnY72+/XTf2SFjwLp1Cdu7wf+ayEpwI/RFWPx/ERnvrdzwsnMgyqh
FkFOGKpAVUTki1vN6YWn+HDaQRsJhUV8Go0o8QaQIy0vS9V1bSfUkCDjNAIF1G9f
s3FGAnKg/Ek6pzV9+toHMyWpcxJsCIOHDr9vvgVbdO6kHTxXy2VRMOyoyy+cnVnS
xAGWDyLOpc9Pvz48HAbzHo+N14570ODUZ3+tuD8szVkmVpNtf28vLeNj9RA70mzr
THLJpfoE1MctyvXc3UUPSNMEXs0UJtYeSpOfLslEuFr3+/XHUIjE0EMa885AfbSG
l/YLIIchMhH9I2NziGY4FG5HNbORbvTw1oFeNkT59Tp6xQ5TDEQrHFWY44SnosgV
2UAsCWwS+EfbwozcITuYtlPb6BFAykRvOHANHSMNvwRz4UogSVteFUW8EK3kGNhd
gTAoS46jo8Y5/Q6esFaseB+GjUonAew0y6/QaN06RtlVnRiZ0uG61KdrPms6n6Vl
XUUDwoKR68xgHDqPQn2AziZFO970efCZyQn50jgKHMLW8HvbKZmhIQmQnqHU3FcM
qmz+GisR56u60bcf8alpTNYucqjT1uHTlE9ZYgTLMPKcpvlWbx7FZb//nTfkIcWo
KOD2dGl3L+NenFHUZjvrl9FpKp6Cm/VgJKQxD609qzZULaEEO12emR1vjJrw7oqu
5hGD8GF88gyWcImGfX0Lnv71ZZNA7RVa8Ffh2sbtLMzpfbnfqIKfPEJVyNOr4FTf
hZYd7448F0jjKQovWQxU6ONr9GXV8ZdmMMYah5IG5w77Fa7qWEkT5yPZyNPup0S7
ecQ4tB1QklCmbVSJpwT4Y1JO39eHEb76PmDK2/tFHtnjLAY6qsSl1aE0MbuoF4lE
jHoWdoBNI63f0F2w+OqLWj25nlS9Bod9bFgJ80S8S2qu1ZpYwZCS7j/3Mxz4rpIV
WITMWB5WkbAttUR2sIkpXN6SX0JIU9pwQGUz9WICzLt/XuUpI3DaNG0mRDomWY3Q
id5Np8+sJQxa/NeFUC6/BvESDL7TsBlJTdTN0BPFFsBxKEW65JtOAB3cUU40VMbq
l/D9dzRJ4pQMn0LBhhwdCt0BYaW3IlYdlJmosYh1nPRC834/CxRg142lTxSMUXt4
8fJUxmRo8CYuGUAQSHGPU7fIVyHum+fb5vgDxD7qdTMe+qs2eq1mgZKaSuSbk0ct
3pTB0iJLTNbZD34MAOLQ/rCNq68n14cJhJu7VNdn/VhwgKs//7xz9WMiVgZkKEX+
hmLdpRdnopzJicZaMpsXSFk2VJSbHl7jq6fnw52KT8nSwlte8HcX0P6KOwuAMjql
H9lmPiVnZqfTYrrk+J0VP7yxZLEMc4LGo9C7xn5HDeCvZdw9tH31lZntEo2ETALt
YXqt+WqCnH6KgJYmjyWdD06Gt2ehB+wziIRaAYfSfCGPGQrSbO9r1594/pup+m6U
Qncupi3l9Q9UWvXs2SrFdxmVOuoUyD0t1FDxbHXmXhiw330AqeKc+3Akm45d4Msy
nr4dlPZ99+knoeSb2M/klXYctmEaSJePgbroroS16xqstvK2jqg5sD5PJK2z6MvC
mXMEjXTXYmA7L7St61w/jY22jaBkf6CUIOzsO/l4jxPmqiNkKCsWPXK3fhZ1TR4H
qjxjNXCth+9tx295M1ePD5fZonBpSb5ZCrqLtmVLcVjBsRwU9kJAryBQe/QqMRty
ddYGOi7jLKAe00h6VW0q2LFbABhgzdKm8guk2OpJBNS0nZqS9ctgfLdrXLvFk1cs
5IwxK4g9Ytv7+T12IZ0tabe5VcVkkM2sGgesMEGKe9L27Wys7ds+sIhjK8KaKNEi
tw3hfECUGlpTc7iQ9NSb1NoZ0jmZU2AASfbenK4IafyrcKQ2jsbOlxaSpruuSnPL
GnzxYd0c49i8xCzScgpeNDRw7HB0AZxMfZlwpDVsnfjtXsMkt1lLuw0bPEUWmm8g
3yqIAE5w2kn2ZmErXec6I592ruUSXrFdLug/tjEUYNaRsR9lt8nSFi6Z1uZ/L6y7
5Hl+7FT/jzAuKpNkypZbf11xfXiC6zw7Oiif5z0IhUEDolJ9sy+Wg3OTy0z8VBhr
dCahA99tpEICqGI6G/QC9HrcraZo6P+b3tVegnlRb4pmg9qTBoq+sDboc+PMpjzB
J89kENoXTJK0BMwz7HWF24PqiKU59xRRNXv+In0utEaBZ/cUPxLXVWVl7EQl1oKZ
dNHqbOHZltvOYXOshiBATOLESBqDdnwM9CSXmr/Lq5SiyjZ//ChvdHOT/aG32B+/
ENOXyQsQvlGj247XSnCJuUF1q4C0sCGeP9+V7gKBHUj9H3+mXqDwpGXunmvMwQyw
UClunSv5VdDdhp3nA7nimEdYPLiu13YdelX4t3pbmd3oJ3i7L0AdlKFrpgCoMg1W
UUOsY9UWS0xZ43tVnq8kgOUrO+A5kOSA36EiYC+TznoiurYxaaUwQ8ze67HrKkzm
2AUQ52HtvdCvR5pbHUUDfvTvCg0Lc9g2kNI6rbfNr/kLyOqTuFU8qINkyrzNU3vg
ES3edXULX9gKVQR2R6dx/USYAFln1zwVR2llx+TuVBlqTfCr4+vslxtTNvhL8+Nk
m7stvlVyc+APdm5OIUyJFFEoTk1JqEMGPt1fJnSjkX+rHN4mbTMY2VZcmR4ewtw7
cMNQu8YJ/yLL/2wjXbQsaYug28L7K5/uvwnsNNMsNjmXvh3zAQtXmxkk9KcSwqhy
r5GErbeCAmEEC3hXOALaRYQW36T/GLDzyqjV+bqgx+0odLgKvrzUFg5c6uIgqWGS
Y/gJVCxshsjBW06db4xRg2cexDToTF2rtCFKgEVjXqeN29TUgvOprjeT8ZxsI+HB
+MArg7yYYfvXc2gfEtuJUY6t5TKo4lwwlcXf5valMY76jHDxSBb0ZPRt9zPlW0DK
SyjpEMV9ZYWUKeT4pu9aUoEk6YyzmMVFLZywRWhSC1ynarwqh3I//j2R+mHQoL8Y
rUOcPTNXy8Udd4eqrPr8D172nLqk2yHLG/mkAOj8XnEbsBxxPYyTVTxEKnETStpj
qpILyRZOZ4jz70EVckmXoXDxoW3TEdn6RQA4bxzSgNVqaUCC8nt6rZe2rnpBaweJ
DarRrfY1WOaTz75aOZYbLzho1GxQmyI28LmZoo9QEhTpK2s4B5Dh2ak+641Nqr/h
x0rtKK1hQ1TZJDfzhRGWhVXOHJifmC56pcS6mKjWdG41O5kZsLpkTVUOEHXYgnJ0
4wwNvlS4ETQ/ZstFidTA9UbHleOGqvDIa4QtBqPNOFNexj1EbeaFhH8Vbc7lvHy+
I0d0RmjmJPdr2gKyyFMF0Lbs/jKrrvJ1LZEIurBioakQkE/YIoEn4YmFMAr3/ox+
/16PA0QmxAUAIJRRSup7Fylj/RtoseWfnzfRw13JqdgVyKyUGlV6jXKgEwqKpkp7
JhwuaxoIAMOs76YJAsd7h5geq3RXUkEOO1pHJHX70iyMz7imnKkC/VR5HeZZl4Sa
oNpNlfvzqGi0xKrtL/Rgxv41gS6l1A1dA9wZuq4Bf5W+uGTU1s8hFsa9+LEXf0Mu
gSoa2zAxv3+LvrXP0KR8N08zIknlQnChserqaUUH9Gka7BJ6i3ccMSFqrtbDNta3
P39Gjfx57zSXrNTLz4UVp/aH2jylYSb0D8qOPGmEoo8tOgLg3SW0norh5vpwbUGq
bg4TOLYZGj5UKMqrwPmn7SImCzQouToT5bkTQkL4O18hrAQtzj8zhDUCE6N6tuFG
JgZe6gl1EwUguabGAOdAp12NXKbPkXJEYeD8/9Qj3YRBC0hVlWRdg+WYS8JYvwyj
3E5Ct6b+IyZXkakv3AZfeqYofTx1MLp25eqatUX9aouzsCofQ7j8cdqQajYF1X8h
6tW+j1alnP0L5ZfyZY5qlXHIXtLuqtuPG8B4D4vfYftb9LMiT/MV8S7VLQnpB2uN
5Cg7DeitXg7yGbRIAuPFhjW8nfS3QpVmOQE0jqjMGRie/7Hk2FyRsVtiY19Vx5UD
j4XQOq4RwxerF1ewkMtoNXvbJDdBx8sPicFIoPB2nBGXBOxD0KqVtPuW9Lfjijrx
JwdSTalg1CuyfGMr7zQf6JPNnllFojTvKUC6YUTrTiTZBSciCu42/7EOGHOUb/gj
oPnwz2K/UgPxCtEBVFnWSPnDTmycm/OnfxSzjEYCbC20aJNL3RSFEyZlJ86mPIqP
6UfurWnfiOkiU84PuVSPlpDnBBgwyKC83L+LwhRn74It7nYKsxSru35X2b7/K+dO
j4aomHNytL+zXiLoz8U2fiJUubM4YmgvS90ayck03FKc4kY1ys2RU2KHcqovk8uX
tJvsN26T6Lg3GguO9XqwMeAu5/greh1Qje2xyS20V1/oHmwFT3hpC5uetmSOGTIG
2rdkC90hAM0ZUsoZfxRsQdhgtv2FM7fODyFpoweZlgoIgBkb/8dUWo1OUG6/I8ew
fjaLobSHGhHAbvBMdfSC6vNFYFfZqVaFlEc4RN81jK2sqvpfbJTGccsW4HN5mFfD
8/89HOPy3E7ULAoAVJAWf8n4CfvFrPq+IXmwp3RPnv/Yadr2mJVfm6SZxI7Hrt7v
6A6sUHjWwz6Zp748xcgUf8gEigjhedT1XYb/05dLNjBnKeJFdnZno6yR7olFKa39
2aQgpzRzBaD7is2okQqrXrZBQrymQDBG5D5cZAWwuwJKrN9DOqCq3ca8cj1WeOac
KkINbPOHbNY00bXoqDoMRXuyaT7YvKOZbfO2Nhfayapz9GvdbI1FOhwmpk2BzGhI
8d4SVZ1tUlkcg1T0yiRVk/1uLVYzsj0eZw8j2m6osi/S8qAxsVxapNYCqhFoJGav
5anKja96a1NYl9kvDPGCFUQhYDFBcsZ+sB63lgmT1YkYwBHper2CzVKDfu0a22nY
UG8gCU4W1O3LhXnkmnIRNdlWczHaZNsEwpk9yNIj7eEa1T7cAlOmyiHC1lXklCa8
UEDze9XxxGoIIkYKt8EA2Y6Y/QGzFN9+w/wS/wCeM9qCYbPGeqbm3Dt2rPjnhUuo
JQE/ai+lmhMzE+bxR9+jW3vtaqTZQb5yhzispzMqPH+WkdqmxZtl9shD4Nt/WS1k
1t7a9UrSupVq9zMtKYXNzcA1VJBXngVFGARM4ODbM3ru+E27tUhxJsLNkTXvGDdh
oK5kTqoRsGdpcj9xeNGKVKRD3NWxNWMbQrcmaA0zwZfkrlX08pkLnngTDQPg2DaT
y3mr+B4GhTliBo5OdUFxcAMkOJuO5tIC8wDFWUI2+M0sosIXZS64gXabQMkryQBD
KFUTGYsMfUopT7UCQfOD5bMjX4e7VR1CpAvYLtZCNOkIBlmS2m0IakWxmkEU9uIJ
ZT2uTAXIlo6hE/B7FiKgGzJsFsOXe/ZKLj5BqaCk6RXfpWz/WpCDDTWkoREZ8XCP
u9nvnLNY0X1gPUC5xjxXzm4FvUa+VpiBbT8e94OG7NpolEFwrUqxfB/0vJRSr1l2
5XUih3DG88KTNLJkpIWGbf3aGgwdDBdG+/llxWm64L7HOCD14I7RqFZ5piE+/Wqg
tSDu0pRGSKEHBiKhssU5e/8X/Y2OcrQIQeBGBlrG7dMfNSN74/RVwIvkkegiuQWh
KSCmrpqJl28JzG5A30vpWT7jj0cpFyiabT3mjlMrVWkGZJHbP44Acy64Te7/pLVq
bdax581rp6R/UE8vmOiT4p8oBqtqLVdXs899FYdYCnsZNKVWejk+N+zt9kZbeo8a
c9WH80tGrJbLAzgFyonuOmC8d2aFBR3dAdxMsRdC5zOlLRHrR1v2SrhIgV5oPePW
DFWGmoG+NKOiQfUO1GeskFztgPW3zxqsmuZQlML8B1e42vs+Ueoh4x2WxCvvGT7b
pT6nxHNEAfSO0OgNnVI8QHgICfLnmVCr4XFOzCp0ispJpdVpPx1CzD/nMBhQO6ZI
Bp1QxURaYB6cOQ5twDKAqHAwZvGR0sBzpnI1sKv6v4MXWKmXTQUi8uPqy9IiNNI9
DLivUmwBRmEflw1lUqdv+NHEUC8Cz/7Ahj+WHQKbXSY89bjoBZZDbv2eMhUfin1Z
dzkczIR23YTDmG0FOoH2sZJBaF19pF7dggD7BxzWcczl8H3EBR6QiF/2nxzcX4Z6
SmEfPRC0rvVFVNADFzCTjstYLGjF1NF7Zfs8TD3B3EwWsIMk6yj6oiFby4MScsoI
ETvrHoVZMPVinZ5XOqnYLWFyjG9PQTqpIsHCrYVzObwMR1xF9XTrlli5blHR0How
/9bGnxBJR3kuUDDP4qtDtVjYPC8xkJL4bFl+jbGG5DscFB9rDdlM/FpCoB/B10+u
wL4pkbhGhe1BXfNWWj+o/ey7f7RUv4iERurVdTLL4hX0yzhxbXsADl1rnMRKOL3M
mxAGV+DAHcEcFpdgYKOxbt+CxnXXX5jvLTlYS2swA+rsbNA2uR6+h0cefTZcdzxq
O2qreTLY0mEnBFdsyK60ZQMGd5OPrSA/eGUNNCDbxQN1pzVUeESTNULps7XgF4G6
BHf/sIXPuPonxtwhIa4flB14jVULnCEMXfKlutZGbHMTANaVHojUEgCuarJaBgO5
jt/xPMyfAoPSwQp4N6Jat8YNaKVXAeC5b7hcNshcuoaGbb8hILsEGctwkjQ1ILV0
nveuyAiBjrZgN1ypuAIU/t5+waLLiDK6w4f2r7wiysHdqlERTBTohTosUPWyNquF
+yTjow5HocxvW8KEK1FSj+3He+zdOF6GIFJsNt66SMPxsXOYjv1Fhk/IQtYQKt4J
hY88EpjFU9xdcuOoLBFhZkDj5RLtC9Jy46rJa8m010nyiYV7CfkIjSAjgbJnDjT9
B0ASWxxsiDdwSIifUaPgczZ5aWg9tbJCQQJZNItnewyBd33zgOjrrOXb0VoJYbgk
f6GNIDDR+8BRZv0+/hVeI1TVPyFpYhp0XQRB1/AJoMSJx72rlQ+jxteHfrZ8K+6G
R3YGDeHQb80k1ZK0THj5rzUKBsGazJWzLxZVHXk2E3zHvP0B0PGbl4uTsH8GqZQu
mYQurctPY6d05XSnRkjDUa6ILuhmbvueCtMP1M7LAsYt3FZ/Z/kwQQ0SSAe3/Qpa
IVpaynMJRE7/u/bdm9MB4TnyNPyf5au/hMik4ViEsiW1osx/SFB4V4VYqsiRodok
9SUpUKXErkpokIJJu291INPbhr4rbDDAKTPgL0dyUSpWbxHfzP30q5kb0e2ObXuC
81hSu8pF8PRTucl3ZF07VEKJ3E0BZ9UYkFgG5o3JwEt+m8nY9Emu5ndlPBXIEd1y
rITK1vQG9aDLtllsP0MjzvVDvP8PPKGmCj0bggvWRq2oLT4kMJuk6P94DkvKItEC
cfdihBbBAwKZMe/TqJmA634mJ2uPTS5/whcEleYk/mT/SUAP3kS4mtz2yZaiWB9t
NnCx4YDdrc5HkrwzBM8ov+v49+KrT9VnauFjxGitJiAVoz8TCP9hfW7b6C1abquJ
Dm0bm7egHzTICRu2imnp5HNpbk3HWUVV+AMSlfDLeD9QeYrvDuSYmvkg6mNlsYSi
sfz03hyYyMkzTv8jPLmoSobxYZ3sKI7Y9lf3sbo0qMyEHBGjtZLCkn4pJzJE6m+F
NUqU9gCtE59XfA+5495GNJN1LiQjEJ8bJ1Ltwdmi/BF161iSgNV/Oyra1tqN+Nys
/8QlzMF37a6vS131LpdjWbBjNrRwYSTBxpshdZz1tNgqGhplUiLe/MX1gMof4KKj
EJXS/6DYMP2QgUFklGAG6obhsjAK2MmN0ysuZJUT9HzBv5s08mUYJ2HbcYQDG6QN
oM9ByM/L0JAmW8VREY8ZPt0gNt7ymaqO6zkDGLU/re6WdnI/c0D9w7AgXxfzocyB
KVTeryrFrbGryDdUFrUtC7ccALK/2BD5FefjU0vEcYaArykvCSq6NxDPO03u1/sE
n5T4k/jORn7CwxVVVgiBNDxXn1ZJTBaBEagEffLsLOcnyeO5cmnfBPWJchTKpgfr
Epa9FzBMlpWU4LbLj5UwKoe8S5EAtI0Yc8F9mrpiYjSoo8KfGiiwy8HjgZX+JFz7
lJqjzTSHzXvXpnJ++pU1yAtQk3Mg2hsat9WoVXgb22yktYa+2h03ZvvaHPN0J6i5
7q0p9kfYnN1swriYMmtNFkn0Q1wg/zFcZuK0In10xQSRr53oQObqYzx7R99jhtcK
9cbgYfOOLMNd4yxQOgOJGDHivIK4EwsgxLnN4B+/QRI2Ksbv88UeBOJljlIMTbDn
1Q3EdYYc1+9WYT8P0PESwpREihqcbOvLo6hYrEcuV7gkctS4k0bxBUXPx6aCed7L
KEeZgi1Yp2xpFB8fbEqO/Jav2PDsAKLxgqf4eXK2fmCUrtED6doWeJvCD9kQKKgu
4GcR/ZcscatwFFWAgVDCO6KyOx+dvsweIW+oYRqC1zVM1ukXtKuofXUSAOwA1j+4
RyUaWIfhsabW/+m4yiQwFOVTY191Svr0b+usVqZcbWfKEVf+ktddXM6T/LmQfsb4
iosMg8FVB9yeTadi98DrCkwsp+8lRPa3rZzfmJ+Sf7dA/PzebPlNBW2Lv0rB/Xmh
Ym7YUTVb7OMpSvimsNxDBH6RtgAkW5eQ7/kST57awwGvl7qBPw5f50LytMuPlxmh
hE6kEJWQYYxqXcW0B2LyXm/P/yjrijE68bsH5QLsJ7iAeVIDgDdGMWlV8cL0Kr2H
sAuJgDc8nn+nav0ecWRwugBNsOHg/LOF7E3s+P0KIrGBbPsHiQ5IVixrhaQQULKZ
5wtl2xfnE9JB+VjA32IJ2GDS+jAe8HcNYUZzQwlGC6OxN2Fe/0AEsi7MgRjzmBE9
lyLxkoa393qwBABEzaPBbwR6epebyIP3jqbtsp6Avwd/1+nB+TbtSiDiSsoSsCHP
GGj3e8GTol0VoDW9zGRA4NQOfbNWe+SStfSEJ4BURmfFG/ROsnBz1qjggpL4VNRx
iHUdPG8kHR6vWl4PKdK2XcVCJ9XjHgir1usR5eSvRw1ywB46v/nrO5pk7739OgaS
Un1oM9Bn5pU7yGZCiVmxNgboMlSV8NkNrTasymMg4pWNPCTv1ID3F6unLRVZTjFh
uyItvaD4ak/G1Dbzgq5Yo22fL2/ECVv3SYATMtzDMjz+L8mDtslK3UXVwoll1s92
dbmbBDPL7iB2h+4XDQghDGNfuYCGyBKiCtYAWQePBkIjyLiSMwkzzWRz8zLRqf41
0dDY1LDsu1oyLST9YneH45aaAACeLODUy6ckv9z8K20qx1dGHyXLnpob4JWReVSe
T6pS8tFcMIp8Tb6FyMpp2eVazBwQsTipJvrCzjjLtVaB/jqBplaBMHa0eT1wqDvw
clhI0Q0U6WoX2U2ZOUYuSqewbobPjCmZW5vCRQV1BzZoUzOGsCysoZrpqYRhorCG
T2U5Ur+CpoQHuyk+GEXED5hIRRxrrAyLT4/PKEEdhTGshcZfco/qtYUnGh3ObE2Y
Xw8xR627WjQ5MJq4hQSBWfBDLCKsFVhmL6NzddtbkQL4EADJPPz0TJ2sR9OmyY4U
7V0jBl3GmmGUa3dM+HLn0Vu3/dC/Au9Z1BoRstyyML8VmxZ3NdSb8xd8ofMbx93C
1em4MmzYzYeTTYtCO5JKpy39Vqgyw7X8tbt9p65T6JvoZKVCe3FcivfJSRBufh2p
JyEcSYbbAaMjw/Ln9c4Y5qynu966/013C8PphFGXHjKg/PVTlUWW5An7VK8xLpKB
GA8Z/scmhCDzp1UCVhS8OwmuBRXaB8nqbLzOkiwg7Q9DNwoBtpz/N1v+IjEp8nB3
7bjjsharX6ozpR7hdA1AbeHMLh4mYdzUDC5wYqt4uTdtFQvbwz1fNHmoB/lMMYT6
aXgEmVngylNREHjLwedVXF9fLFCh1xweNWF3/xFy4OjxODyRMNqTAUZxFy5GTnpF
qedHn0tF+EUakfipsY8KmsrH8ICUCRucOivhHwRkdQ0FHGemvatCh+iehsPOZifd
pAYolAlGf2cJNKY0SNDXJnuZcwSA/WoVAP1zdMjgs4dJ7dPy7M4ck0CL9Y/8+Ie0
i3IqYLqULCHa99WnIeWvW8+LuCmKwJmB1uryw+UDAygMRurfmTjUJxmsq1U7L08C
Da8fNrabMVygX3erXEhwbdEtbTk2wgVL8OgjKNMRJ8EGrmRTaoDgwDRSDc0FpVZx
dpQO6B5BbBzJSUEAPq9g55x6fIvsRVxSP/2ET2tSFA45vPOwDmD3jM9mXi/caAhu
VVvF7r+uxYsRCReRYtqAce3u2c6n4/U/ANKXGLbMD95b13vDaNPWjPqQ9fSLReiH
weqg7rkxgm2HDTfUaEI3XE1kjNgIY3bSkM887wXs7lSYZjgyOS7h1v6F5o3RwU9V
g+CECjuf7AOR+qkBb6PwCWm/3rY23HQroxXFCRPykAJU5n0wquCHDYwMkyyELIA5
3U/gmBUuzYwiIRh5c8Cvulbml1sQAzGNIA6AUEztb0NcYQrVrETEWCbgLDp7Iuvp
+23FlVIXoiG+I+5pHtjJ4wXxvzaFUergmnzTx7IyHpdkja59trscHwFOt1YrtuNs
x7z5LdzwKwmxNrrVPD2ziGcJ420htEsCx4lTOf5tpqrLfHsX6a1UzvghkmcqHhwB
Cl3ObBD0VR8rUGobNxtc6Yv1znNyV7TMutzdmNKoAGyZv+J5SfMtN3XWtawzPtdO
p1ccG4h+3hdDBGqGiSTPuWm9x+Jof5Wj6s5IRXzhvchd4Hrfi+AEna3C2mB990vL
ZeB+WA0mhjIUxO2u2TrpcBGyx+p1VA1HCI9divi+ezHSnsu5pKJ8nMzn6e3MPqQa
QbK4EIPzAJ0X00O9qRqV3FCvLh4vc88J99ew74fDSUOej7ze7kIgN1jU4Xo71hLB
8FwHtUzYuqzONN1lUGNX9NI06X00FDv1Nz1/xKZAbS39dUNFxvBJEAraVF5sANQU
7KBuen/iPu/b1wunmoNKhQMLsi+5u7NZMxnhyYHb/ujOHjjJsPvcMSgNhiPJR/q+
EP5UzdInEqFvMuaiJdHMGrShlmV5bKdf5E+v/sdqvEHwmcxwe/mncZodikS2OMY8
Zdw4m6vsTEpN//kiAWFowiMMFFmbaskk3z/sSx0jfE1+t5enaahnKbWlHvRZo2oa
GU5be9wW1AAxpoYG0g6tFCUfA+fzMqKnxAGQfk69yKUN/oQuuoN1cfo1Wlw1sXYn
kA1qozceU5bSmBFAMcMaiKTbP72ifd3BCLRCGWg/ql1FvvTea4oGwN3N38s+vx+O
xw+uEa3+KCl2yF173/6qpFKNDetwMYgtAKPJHumOF1yh7XfL0nJp17Nqm4JaeZoe
S7HZ39AZOG4eG9TIRMWDr8oo9Vetlfv8/4MIhNa1AOs1TPnL0WziYmFUsq0OlZP1
n+CeGWQc33Z2l4TG3vb3roKJy+2uSRm9/noX6SsSD/fojL/bNU7ie+0jm8rNzNzI
kcGaU2Z2sC/L1vfN0OVZqKEfqfgo7jxfSxHsVs5ek1a+8Lg3nDYFn6P0s35NNN3o
pvhFgYPxA7RDjM4X4yatx78pO+G0QSyRYHqNRzJhariJcBDWTqPPf4xS0HYtODrF
JKepFqhVeOrmstTBfLvtpyXh0Fjl9YRgH+oLUfMKU8skc87O6121Jmg16BK/n3Pu
NnfSLP9hNQrcYNkeAIYhQCHkZHZhlo3E8USI++1c4WOudKq0X7lfM4Ht/ddeLBA4
QLSi4T/q9MJ1M5alz8Au+1wa7u/37EWGNKPT9Fk7lKfHoiH5Da5TWwWlLA8pStSO
vsnJw2E+IW7pDjKaJknnzmCe6QGGRfi950Yj3LRZsQKjCE5i4gG+dfWyJkBW45lt
94rcQGThg6vMu9JsjcBFcQvEMno95GrUZuOk3q3h5/lCNxL288Eo966uhGrjNta3
I9hKbIFcZ8bWDXbAMALwnLjNVqh7GOLHAXSoTEOv8CQ9zrrmgzhrNbNxeX1ILY15
4qq0CJW/OlbsYBPg1zse+tAvrAQPn0zRqd5G0haM1BV/coP/DkfnTQV6tFPDn8Bn
c2fY6FnXdga3pRhTsdW+QeKXm+8XZZ2l3jKxi7gRy+lK2Hb7jURjSW5NG7qFZXWU
qbrNwloUlc0RmBYMyqzd4ULJB10xSOmh0sfJsWwA4Rx07XpP2cXe2UjXF27291CE
s/jwfOrxc9Uo1ujvzTMAUXfKv6KCi5TUNIQgmGdRqAtzsWjbKLMySUGSDhU5cyV3
CXnwindhXNdfhYpWbPD1ewUAYGkNO3lVdhvK8J1e66aEVLgGB8/dY/KyjdfPeU1z
U7OCtpg0PlPl4NNLGXj/IYX4AXYBrAvtOf3VqZuSaeW1HawIjSNQKZQNQht6DXKf
SMCP+McVaiIS7LklODY6vjnjpfuwuWNUBzgbYeCxP5JaGfJSuKNViJtq10l99wxM
sEJiWKT05Xvwfbtooqpely3GNWVZMKqipNPBvwphx/UR2r5HUtUjck6+myo/YNFm
vHeA23XZTZy1eeoJ6IGPDm503qRTPKN2zQdFsS2DiA+QxyEHgxSPE0SlD8lvOCLh
Fohsgtaewr4gcDuVWgm1S5oSux6vew2vkZdmwhk3mDiSSQuO1v9QRYEd2+FPFOhd
CqAku6XuYTJ3Mk8pbD2QA126cBnvV9sdgg7k5rKWbQzn06LM/CcHHPyvep0paAk/
OC29Qm9CPykWi2dbPzs1qoDt1m/zBvTgyNu+29Xn94vVjrFZAmRFNYPmdl5ITMMl
Rl2hMYSKevFJEotEmc9i4ibtpTKNeEGqF2qokP3WR0d9T9NHAsSVuzT2fAin22wP
zWcI5I/sz5KfRgo/r9ne7KyJHuP4hR9QuVePgfR7xyzZjzJ2QQaM0uQEo59WefIC
J+e/JooZomqKoUekYthiJt3xSn7m/h8f8S0AElGK+VSeNaNsyCTVZwjIs5zCkG0Z
PEctX6n64/AY3czJbLxCvbVAZWKrkaY9uyXqOLJqo3Auv1QHfYCb43lN9AzXoUqF
yOdFj8PQE9sQyaXJXbN7KAQN8an8+LzELQfe6riViLacN1GBxOEdWgUiymdGDLK+
MfTb36eun/+XRx9nSJ7F1qH0fjRwCQvhCrbUPZGTV87TiK8ieREaCpQxNUc52El+
4zytqZsOigdgQIBF2QgzuJJt4qZ67t+vbMeTJq2g5zJIPEvPku5XdOC8IjjPL7xQ
fk6l6+kh79+ZYpjaouwUzIxhUsYWjZywwV2c1AdKa3Lg5yURBiXkLbTqrPR/u57M
dMhb0yQBTucrSFuc9X5LRIrfmLBJ6IA1oEeHlsqwsJTSeVil135CjguEFkha7Z/o
xWp0OGPumYBuCIBaXg/8zA8hPTMjiKfagkGxJS8jXRrBtwOgZ3XXDdunx53m7qzn
9Tfi7VWeRdMl+i2oyZCpUuqRq7EHxG9ldJDBEMm+3xin4tdSbREURjKuzXi8nvjD
q7Tr9Boe6ZQSHOZhZQyRVo8M/gaLhq6jWDxwhb4b8U4I5YN7p3dpH6bkwJ88edVi
P5u93Z2IvwOZr1CbM8WGsNG0o/F1RAyXafsTEtsmbO6ZBrfTM+QPf2LnckN77hCy
0Vd916OyyJcIVargXcP/qdnQx8vmpI4Tm6fl5SmkU5mnM5VzV1yIFXjL6g/WLVzZ
hXWeVtPflW60zCXtj1zlVbOYuCZjoc9V+irBS7JAOzaWqDT7913LoYIyWy5pcC5N
7T6oyMSOGm2dKgz6k7pR6/E5emIhwztZ3Q0J8+ja3Wqjrs86NvOEpMkSycdUs+6H
uSV7ghkdroYb7BQ3s+2IPRrcvCGaEWoQAwxCEXbyfKMOTlsZHn/ndzc/bQKto7F8
qvkTlTRrgjzC6YbE3KNkcZYOFk56djEVGCbFk8OcPp72t2HwMe3dUqbKnZIea1VA
YV5/JQ4H4TnsHCHVBAR4bOBNdvcA8jxfi5rmYUZXGVyax+ZymuvkXp8rkuhy46FD
f1tYSKZAelFPG8WBbDQWVklRpznwsOmzZepn0NUmxm3FqRxo0J6ijTI7GXqSCTWO
N16/GiWymoLnGE9meqc7E48TUkYs/pLJJximS7uwQxjIDiPIcl+Uv2DIlWyRivaJ
a4aQf3TDYxtnPg5GLdHRjBHqClZJlCwQB9uHhM26zGdMO4NOimqPDgogSmXLwMdi
dztBwgLTVVa74d3/h3PVa6t9E4jflyZ3tgsb58/kMDzvNBB9J3kwqnxRr0QwB24/
6JGoDErzBg8Dd4mhW+Le1FnVqGnuS6cxStZtgh6GM7yCFWAm2ZaJmI75K+2tJLC+
dy02D38zp/wN0wd5VPDRkvdxzFGGgoEf6qj4Qllax6s9glZF2ivUn23YfzA17+lL
MD6fqJ7GNhpbPRn22Z1dMegX+lNyqppZe3qfnz6uPSSiqRVI3hxnrq4CipuNmWRJ
Tcg8F7ZBqYQdniEHAV/FwWMsc6CGrPIo77NBLFjl6BIgdGyOTHpejeGV0ro4z1ZZ
h50Y7uuINXytffWwGSvoNBJ0MHJWUMUFS2iXFBJV71c83Wk+gH1V+NMgmSCpoB64
TnIDB9Ii2I0OB+YjzsjN3IdnDcAJy7U37vVRzy0d4NJ5RQQqvR7LUMiz8ixl7M8Y
I3C6RoKEYFaqwkwq7dEi4XdLFNYbvtNAQ0rgPwIx59qrp+3JP8fMKak2aC2dZRCV
S7JCo84Y3n/zXZNi8gGjgdSLN0QlflozrK3ll3qI90TmUt7VAhQT7aW6PIN9F4wl
C33a1GVe/+OTDBYu5fjgPXr23UArvFMIHEC9eg6x9sVpQL91WCnvjF22ZYDqc6L9
sb/JOs2e2gHopkiF4uHnIaWrh2SHOJTzkSckKPiZaSilQhDzeTtg+K4FMAQomT3v
62qY+bCj2p+uE1OW+lxvVXKCTl8sQStnu5b98DkINt3Q17rC0K5lXxmzb9Ehhov+
KM477bp3mjglyNKS8fJzn/BZo/HjFiKrfaCFWCwX4egvxCvWxVCTNxH+xzsxT4Ck
J+SPEd5AvTo1B2yU+2xbmVP30awkWXmUNxqoHgFGZq1ZHYBwJJV3kyZJ5KjAxE6C
EHJE04Alw4FrZlUQwPd7GNdMygMcd3SxGD2q2ao64cGWBiKj2dXsmLXz/rBTnv+O
FqVTn+v2EoV0cIPaepZZVu8ULfpqhNjho8xLAsMus5AF6NNUcGmOhPDHuTN9g8jw
Upvx3NaUyK4t1q7zPfOiDW/VbFFTxVwWlByhBc6e7d3+63NpoLc8ipd7zEc0YDTK
SiwY6oMD+c2gfKr70lHGtpkUVQjpH6T7650Xr7Er6gwW5FyYoPll1SBz/wd3HcLk
ZB4climEYtkyqJZ5F+L78klz+Q6tMxaX8bIYZDIMdrv1rFwCcuXaOx6m/ftx35I7
cmMM0BD/h83gn11Tkh9N4gmjP/seIOQb9JocNpFKerOE7BKPePlz41Lnvgs2cQTr
T1cFDHTp49+slDnPm/UqVN7ZT/FvpAoBPLi67WaFN/ZtGPNabK5XkTGUF6F7sL+v
Wt0NY2VKitukir6iwsVg3x8gzUSIaEcvDSHUkhewrKIPOywKpEHRzXjATev4KOyv
i1t5naZoJvpCU0Nv3pNnbu45c9v+9q6+lE1u2F2bFQwrUowIl+kK0Tog22kNmL4h
nOMCQNpVD6eSSKK9+VW8g3+MWYhzRPcciErnda1ToO1gkrre0CzOmdj0Fv1Rak9W
vI0S6o6YC94n4YPoQIyFu3u6YEJ/5MjyeeUDDd5VdocSaYOlUnLeGqnJ9ZihE1Bv
SAp6AuS18iIkVKgi5izcg2NM0wuAGvP3LMwSO0YWM+vXcsboXDCbcRkqZyjxDYNA
oa2YATq+B9OJwvo4947TPZ6dH1ohcwnLBCXp5aTElb/il5eFgzX8Tn7UwQkXEUee
oASMWDaXTbKmxGG4XuzQtVb2uPsqCNaH098E6OwEUj65fZ5NtjFnyBTp7KgCPpvV
cXt3ktYEKtjPMlOKTtSPVgENMdQ/If3GeJzJxlVWaYu3pr91rsZ5oZ1uDojmHnLV
TDOzlfE56lh/aqeDcQ3P+negqiEEhCkmL5Tw0OQxTQEJxCd7YJ774b40xi1XV1WP
KgEPBMyyxwrLx+SBmDd5LJO29GYShEb5QO3kZ0qUfukYTi1X011Fn4+31kBBy4kv
T46H3mYF1+/Hp2TswinQTl3GBcvjETYJYCvznEM6vFvEuwLwonGhfm9b4uh8AoD7
7j6xMOrZGxz6LTl2gM8aIjMlU0r9Dlt7EerEU72AS+iMX14fEZuV9oO/jTXa84gL
mmN2H8390BiRFE40YfGlgJOIvMEYsJ/jIyuDyLO3gv11iXcIKj+FrlFpDiZjIfdr
rHzZMpPyurrENCTArOnq3bNmxpBe9uKS3rgd66uE8EJtLL2832DxkVOqZQq0Qrtz
aOv1a6NUAy57okcgkD7OvBG6jyselp8azanrbUmn9GBAxLyqfjnjbL/ZoHlr1LR2
HxE91r7pU6HaLTgf2lcrbtPbg9CW2xcUzuTfcFyQhLT6AC9vnBXz/S33dZdIT6Pw
GH0WaTTFZd+vmuv3zO3dWec+BRGUt2s1XbNNyNZJzb4JXGXBS4wrRNXACL1Ad0rs
ULPoWzcKarSQc6TDq9LBc3hV+KF1rzJzyOyd+XakTtP+S2AcR/4KPU0eQpgHK3Rk
0RHwbwPvNRfTYVIXckmxsICtnvu6mssn8QcXbmnbMcRUHkbaxDjW75Ep+ZhIApen
/7MiE+gPZthb9TmjQmdRybRfB1QSNvGAhH4NOEUQ8y+M6uoG1qoRsFsBx/9R1Ojc
xM1QLoDzj2hpxJXkba2JCIJLfQSfASPNAtGQDk5ek0RxFWgzPc16uJP1PEuevtqE
DX8uQdx4Se6ZXASKDchq1M+A8oG0W5wHY2okbL1PpuRFxKgURSlXLu2oNGIdF936
gtxcq5oYsVZehq82VnOaltiNJEpgVNuQXAnnBHAc0Pn9+mwrYcFgn3gXXzC3T3h0
/D8CHUqV606H/5OtTQTM17DQYMueXcsibAsc88h+SQBy8XSmFIfB5Wxfv0BdNLPh
3lsUq9R4PcME+p4GmYIThivIDP8LGh26fcQULz3BlLrB7aDue4dLOTHPLqmgG3Zs
X3SK2mihL90MKlC1LYY4IpIsFMUN1B35EB8dxx23jis1/Jet46IUIvafo2A8b+Xb
pHP8ZjLuFKuHb8yOvXoklfC53NME2exVcNghtfPtjIaqUD6o/k1d+hEAgbI6HpoT
YcPT1+/kKbQSWpBGtHadO19dl0obZGumrTF6K65JgdXhFkygIsh6FwmSFNzT7ZHR
w8vpvWYq/+Xmd3Is+xgqo+1K5SYxrxKIx8FE4aufLX/M55LRTpoQIHjVavR05BlL
KglM1exuwfZGUzz8yeNIeKVIRuqRr1vVZPrlPn015bXNYnIQP4VWTs0MrcD3yjVw
84jnNLMCBQLz5+svoM83pHuvwCbwE/q7Qx84iZd13MD9AarQFYDVcNrHkC/7x5ar
p8npPIG78DcdxaNjkGBZ7dw5RrmKyXoljzCXGluwoLwWk6c08RmYsnAkTQtz6OlX
q8uYd9Lx/1zeaAnMlaK3rReyYZvaPbF8Nah/n2TOE79BMkc6cEx3sT+tqftefe8q
bF8o44DbEWtftlCd9wFf6BUywgR2VIPt5cKG/HOxkk/De5isXun7rQmAahGhBqvK
uN5TKGIrJ9hOHQyNhmVMlAevtVscauF24yY9p4rm69MhUehvrAhwhQlDHEtoUMA0
n/sjJob/h+iefvTfz4IKY2H5slNgNmcMtMlBnn3/97O027UP43auMwnzwRDBJkzn
3HhTFLBYadhEqR1DnP2jJRxA9Ta10O6z/8lYfqfrJqEga//Nu6TkNlEneoMMkyry
naZkwoVPq+/wsd9yWb1kJB+/afa7THpC1KHN2rzQJKo8SoVWqm2B2KC0m/5huhqi
3yP2s4Fn8w6yNyY0WE8ND6WlMvGPJ4McHceWsVvpIvCN9X5HBMvOT58DaXm4mBNm
5G7LX68HpyAf4YS0tYqb9iYX8ylWTrdEdSoNSIIDA2/tfVZJhnilP7Gz7BdNLbrF
Y/6T8iV5aWsa0P2EmGeLwqNr9pPUZpygUbFx5+osAat57RN3yRZ6uy0K1EOXCZP2
sgMZz/dx7sVbzZ1fp8G+DUInYzpP0zp/WUEtK/sKb/o5MgHfSx848d5KYyYkpMSA
3BvFUhMzOYYt1b0EUVrPH9v1MZ7cGYx6FUMVqSbeb6Krxpl2dYhdFMu7DSjqn7/z
8WaBfxAQb0LZHbJiWmmvUiU+DqIo6uQ4SM1YGvKrq0HBTr8t26RuR6q93WI3BvXW
RlcMFMiGLEI8CiAiVM8JrLDc0tZ5PSOjYoxo38zBg42IXG4gKmP5YwgaqjX2zjo8
M6S3Vlmiphcj3eLIbZtPGxntOjWp5BnEbJY24KWatvTLDzQoj2Q7bI3G4eED4Xxy
nSuKmIVrDlWT/+5dih1/9ZgAqke9Ts0ekwYBQ6W6cnXgyJOKuoomkMeOzmh/ZRzN
CHohIIY1J3UMSTx+G+DaVUcSi4BHwuAXN1oaa2PUtu1d+dr8jPDEQ180tnW3Mnol
MZScsu5uyPOIhSzQ3lul78yCdk9lUqtUwwqoW6KB7Z+xteZX3wQoXl5ZWQO0v2Wz
Fs7zox4B+uTQ4eDMmTzfUjDfUEmHbziJMs+Wa4ncPUWrHcRRt9pp261eUs2KG8pP
vbPUaTNYGPZwY5NNPJaymQtdKjW2S7tOAod3NzVumFDnNdpEWundiloz/UyxXlYb
GJsw1mxLIfC61bLztHEiT4/8hopZrZ/JSnSlHlIxue8G6cM5/lMus+ZAjb40asAt
gLFcCgrsgKseRJUAcwgDoI8UlIf6DU7TbBix+hGDZ39ZX03xQmNtEpAchXlDwTh0
wk707ygZG6jQTr1tfM8wD/l9oFQbYAjpGzIgS/64qV1K3ec4prRzhjROCuwZrGWD
cbGUEjSR4/cKOdP6HXHYpQ6iPhpu2fyrSlHbEniN0VHobiuVciVCB9uHy3HwXU3k
5lBQgZCbsK8OKQeD5VXdQ7ntEGcGVuTvtzZzJ65MKPVCjKiMLxBEXvaDiDnUpI4A
Mvl+gSp917/iHBPvc67u7YwkbiwRSnxRsORF3/z5ZsxWOs20uGlyBEo3JK360lju
vtZkFiUNIxPHWyJ2Lcn/I6vhQtZUZVgJdjjWOxccPsyxLEzus8SxpPEN/hZLvUCV
xwexdiL/4swHExJ4gOaKjCDrvTz8pZeiRIbPXFlfv1Hvkrabai6+bJKwO6uy1g3+
dVRQ+N8Tmtf8O5hLug8GBKko5ZqCvDo/EqIjh71uOXq+wE/TiVDsQ/giTma14/PW
wu35Ds2Lk+AwZT3Ke6/GFZSgkZS4rSaqUXZDz2JPAv6KCDD7zsHmD8Yv56dy+z5Q
vzkALeIdF9mt5t13zJHVjFZ+ijJTL1N6AOpJD4rBExFPJPn/B28ArzY+CMlSQDKR
ZZY1u4j/VI22EZfgEANqeGTFAUwQd4Wcm4jB9MTF8hZci004HVmzpycqvnMTfraC
y5HX0tjEQhSCuapzWMyR4UcNr6QxhJWe9Qr0iDPQrqwd1S5k2tF8l8JihZLQPvLs
BIKFxL2MNPQLFdqa6a+olQ1WBhJIli6aw2Hop7vZA/MgLefFE/etNTnMzZBMbAru
lzIQLg/0mOJ6QljY91q71UMBd7qDJkeKIiHicZ62CqywbZffA5l00wYDKh8UTB2N
34DStkhfXAfzfT/OAjDx1WZl82Tccxw29wkgP8AiQo9CVLv/sn8DnNofK3IVaLIx
wG/02Fbl9ESgPcQpBWD50cCMSpC1ok+6m7yGkG6WIfkQHVuQ0D2VRl32Ajtjz5W3
UZcWc1Df3JUcH5wPvvYCkyEoqDTUtvahWlNWKK3A9nlyFdvC6K89fHE9r8p6c7+6
xrQ3+0w3GOBfoRIMjR8xRxWobMa8VWaB/mJCElVXp8oBmuSdkTuaUKpyIzBqcEoL
zfjQhuUzOXwB37JDLxUPFSAkO7LJv2oTI48VNe3og+uXK8qYcRJgnRjxsY9E+inf
1WU5lPZ9SjidMvfIBHJ1DAWGgN8kicYYZJ0GkKOQ3dU18CFxrMKWgGUvLNhiXP8w
NA1HEuMkv68xU6gmeFc5y6rzz77ZUPcp50T78qZ1sbYwYR6TgFWfrjSH9JVRPaBc
tzaaQrDU098w39+MbDHjwBKIUJc2J5TOPGI33QfWtp91kE9alqKHmbx6DFK8/a7o
OUuqw+2x87EZKYcRPUh4DMF0QupgppTA9WV43wtA2yZXuCX/bXre3bH9jGVZVi7H
sDEPy4DrJBs9Wl6Id8u0rXDNZ8DWic8WJM/l3Sr/flbnZ/2x2jfd0Fvn2f/t36h+
IBc0CSDzEXPDPz0qKCTl5SW/O2cKxFnD2l25x5DIWwwpVY7mGfAdVDFk+BWEDuGz
/BN64WGikxaXK4zwDgxLuEtBRGLyoDiZIUAP2Xpe3eSkS0azaIg0NuBdATHqs87F
suLPxyxYbhw2JM3HufjWDyjhWLLdOYiCQh5vuwuXRFN9iT8nHXEym/BtqPnMvZOV
NhJ3jclo/ouuXcWEW8aH3lcY8pEokMhYicM5Q49ORgzunerL8cSR2Co+y8wHF9XI
0gpxxJ042tiVLKwaKPPPyK2FGq+zic5FeDFk6u4Zpe4Oj6soW1q5fp1lP7yqvdKl
4I9bPpjK/3eIx3JQUm1aqYV7gPovx6xL6gtbHjj67wKHVMBK3hAC2VzH7UcRKhSs
BOPUkStT3yPA/VzmGfWq80q2yhTw8kjgyRMnmyJZcFI0ynVQQKo9fczzekNunEmp
EBfsquhsDrtK1MPVo/EuzNlwDAqeRya84uaL05tuhu4/3x57svL1mLuL+OooN+FF
IP1LmdjKjk+0/IfglmW9WSQie2JTRua19kgkeZEACM9PxuB/RqMHQRvgqoKHvCfl
gkpS78H88IANyKv0RQkk+NVvGt7Sz2Qvn5KK06cFK0usvCXKrhv4Dbo0n6xRVtwM
1W418sY/EysIcqFRshhaBt8oUYsSdZhjoYCfXFRG7SZs77Vx3GpLs80GAYVmrm7X
kOXtR1b0y3sHhD8k/X1znBj9g/MEoD4r4P0bTaKvwOwJ1U7+YyVd8xX4XxSdytAe
LJ+s3RYWhGohCsk7TwGof1uTRviFYtHFFuzJEKLLSlfWpc2APPHVEfSATG+sJywA
OuhY9U5M8G67JCNy5c9FkqbqI4NBkdEkVhzEBKXOxlIiRLTf623S1X+Z0/XIk+/d
ojcrv2jbnLkkH/Oq8L1FJUmwGlcEgTXuOHl2Kf2ZSi2emSl26i30hMFl+U70q/t+
bhmu/GDF4EzkBb8XSjiIj31D6LItwPgXMzjxOLYzeHKsuTuCtve+AyMfaIyk2ZIg
2/vvW2STvk7s9KHEyzuyI9k/G5ifpnT3D+9t8+dMfZEx0DqQI8IfSiFoF9as7nlX
Qf7Ow9JKoK/9CuOtxcyx2PD/rfLwTUkhLOWuD5YYL33qre2cEz3LfvyXso9+G8Xn
ioEy+oVTHIIhmDSWh73K00zawesGUn1Ss0VI50gCJO4D+4nxIDA8v4Ok2CAsch5J
soZujnW/iWIqEZXikYONMccZW0KrTagkfqT5bA0c40wuiUxzduKjGl2YThh6ToqF
06yN2tWD0DbYHJ2wINk441Y7c5Y+az5oGcnd/SOy7kdGqUV58Svu4PlRc+MoVPxJ
9y+BVu3hwc46G2t0DdJ4bY9lljKbXVcZVq57BHEKSyT9akL26J8MPEOPyvLJUOJz
OypDpoScDpOvj4ydnvKJFvg42tDe88NFqjidBCYzTiSCvyvZV4j1woEJp1ZNJ2hs
mQQ8RGyFAgXEbWoMVZ1GkeTi7uFpmnUoVgVOaDRE5GV3l6kon9gs87Ckks8wPHYj
2efNUw/d18DKTQl5t6RJLPuqzJJBbi3ojAqPOh48T1RQLSTvFcyGaKssxY1Q87VN
Zmudi2K1zzUzNkinQ4iVpKHfbjoJqedw3FoPnPTbqXBYfcXqsQiAXCKgGdRYi+8k
dbAqoPdctXhjw93Oa8ojZFoCeSSicIc31+zYkjIJbpo9UrQrZrAk3riRdi1aFNe5
+/ab4ekcR7+Fb4IhSGjgcGYDSw05cT4gWGXVWggnm3NgUFfbH7eU3dqL2c8hpB3Q
yYpc7PuBMcFrgasba/NFsSidAL2QqY6FzzeOiB6X8n09FdaFrSRDdpor/bVCsq2q
/aYUz01Fn8t1cl6lReYKIS4p+wTEjoFtLQoZPAGrgxbZfD4fNJmqApMfLx6lsZww
0ES0w9BlcE9Drc3hscAF+I6e+/SSS0EzKCM3b8kg8f3GtfxLd884Gnc6TG1eL5rB
6bPDmDpaLtFSnzM84VhRF78reIIw4hKNaalTajagtxej0QafWNXUuWLjKB4nO8CD
Dm3upzM3IqlGFxKOiJEdhdePxnG4PqS6fcBD9RUDKVUJJ+OWamjx+1x3tek5bSk/
GvdVCOYjyFyHWRdqXIw43hWlupt2veyhz3rlxA4fTRTaU/D1ASwqzotEmuAg9BtD
0TcFA//Kq+8lBqUyDHav/268WtEZTZZyYX+zrpE1tQxUbAW3tECsvVLPTQFC2V5f
XlbvGSfF5/Tx8fzF9Xs8R9eeoYPc7/5vvDKRtA17/z93RIu254v2a6py+pe920zR
jFyZplMVPMpaUhl05JSVdQ1CKsWjRPdNZrWlRIGEqmRkByAHC/3ncu6lvf8x81GC
fwsbwaXaIhymgPqh5CFUY7mXYQbETyGfaJbbZthH9ybcvB2nOey36n/f79/CX0L2
yuHusE6BeUZ1MsTPVlBfxZ1YYExVDZV3WeoAH2d6cMA3IHrWsF2JRPN1OxIK6E3I
LzdXPfQEfaOOaWY/NOu5MrZ5qVNc1OLp42qVb92ot3HEqR5wPRdS5f/Sx09o/Nwv
vF4R7rWBPZavY38Iasng0UmI8oKOCKecSm+LwqqZ9+C5lQNUz5nFpTYZaCmSq9H6
4I2ZC/d45D9XUain+HsTD0lpoz7rPxHhhd0Bmp5gI9qru/kxQSwr77RGRN/JT+R+
K9pY3QPxRWpUgDkur+8mgtTthA9WBLegXeaFGUjUb7Ji5bonanAQ0f33uABmQdfT
SNByfcNklLAP56R+cYz1D1/5RuvcP/otuG+l714I5O50mvBL8vLUzbdM0yELY1jH
Atopg5zA3qkV8y3o+jwCp5rqjWlLSdxle7i3+FE2istu3jpOkmbDlrANzkdhmbXs
RZEonDfkUz/RC1LnMUTpJLYYHR4TgD7+YWWigj5oWoiOEBUuAJ0ZlQeGV+7BJuKQ
RPUJaeEUT2W/ZWYXFCovei5gc1sXfPgvoVq7Cu1mDu8+0s3By1rCh8Q8gmUfowVY
VbT3Lwv8dBrN3sB8xeMESZzgaCg8x28DjGJ7PNWUTmKhcMN0j1lkR6w8y+7kdvdR
eNIm7dF2/KD8DPmx8cQP+63tXQWOaMG3Q5sDp0Wgrqkh6EfTxpGWXSIp8T3lxRFX
06mlX6sNJ/hdP1bJC2LYEvuCWQOrMHyi/KcNUjPNRvkeAyv7tR6hiUGD3QdFOGp7
cag7Zv44j2/wgdt4lb+G8qA9CZ4bbaF73BGVoTTONXH/UG5rEt2HjwU6auGDPMrI
qoU4oQozMM4wiqBk5604iidXC5mGnu7Zs4wtH9bngMnfq6FQRc1N9cm2UMGxr6R6
iJ7RY2LNmCNab9GQyYhQLuNPZNNhGSpgIxeX9FJO0s5N9fwxmchwExKy3nW2CFmL
csB0305qaFJhAJSP7rmP/oIqmb1W42k7bh+TjvBZBffA86Ir1Z3cGX8TwlT2BtWy
pujiKvao7l+AHmybGRjuw0RrxQ/1AMuynm8v5UNWQN56cVjrCT04z3c5qvC8o75e
/k3g+bnF0N9/VVkedsEh4h1lWx5CFrYKXfauhOj9UAFEnzOz0eieKBxddpSnzHjO
QgCNI3ofmmJ59cY88rWtTr8VrCWnwe4rkrbnCyt82BRM1XvrygDG7SM3tYdwMMN6
T1Vvg8Aoe7JKYMH3hk2U3V44BsukLxdZdRERoZLUL3LsIeOn9BJbD+o8Rsf3Wvxk
xkFu58Yg9f+Nydzo+RtdTy9iPBQJEVXsW2+ZqE8wJQSi3Ip1sNcz1Z6B8SpJddoI
cB1e836/hSrpwZelkiCZfpZ8K57j2TSFl7p3ZYFB45I7BKFbIQiKCZYQz0JzW778
P2+cPFXMFRQRRksB61SBdq00L13Jjtvq6WPLga/kLD8z+e7KAurgIlIo2JlL2JAc
YzqhlzvUbPsbftGTLkTLJ/5Cu38xdLyFlv+3Bqu+dB+XCxv3jVDXQdypo6J0lAMC
ra0pY9VS+4tFFV1TK/iHbVLYK8SMGPkgEo7tIdQxN+ji2usJ7PcUMuPxg48zX7gL
MdBqxJ+3XI2eGXrEhumA5ONUH8fph3FC5sVrQhEcn9MFcZyCe5QN3F74XEdTA32e
Yoswp5InIeaTH/8QFSyGyhqIH2pr/wWXWSVlxwYU19SYAvKRLwRTNO35vy637ERF
HVRapIvYv2HHiObtldiYkmwSX2TKXLP36DOzaXIy/CneHeozx8Bc9jTBtEXIVuga
16NSh2wPT59rISL/v0Ql/zzHtFVEAPRlUoAsGRvuzX6rdJEXauaOG7SjK9zCiwgN
D1zm39OKk3eirqQmBsmtuancXHlx1pZYp9HuAU6tAchODzRs3x69WkX0YgOQpt0z
uKsIHs5uJo4BdjQEJGNucd717ldNRkmhzn3633xjKY8BSyTybZt6UjiMJcweaJJT
DqtX6NE1eE/fQqsJ/IB4bcz+X2obNXwRg5KGbT//7OpselZ/S3vOrO8aNBisxX53
s5dXFy7gC6/SzGF02eZDVYagTgGY/TsqzSmv6NoveVa148F2PLNyTLq/Wp0EdIRt
YoIvT3AT0uaUcWLfZPepnVWRRRPznfY3kraY7a0aM909k6Eip4Xxc/nc853Gzj4b
CHcrcNHbI7RZh5sXhuHeZuZLBjoKQYwyTJkoIhDAWtUyqQglSa6JAXzx363fjxvF
suSY/OenCM8/P211Sx9rxtxe3kQPSUx75eVzpcwUXle3i1FK6/QbQCZ838thPXnF
rUiT6x5Zjqsdw71OiRJpuXuuBFVWpNjafX52tc35HkIPv0SxKOJaWzgMNXfQJrX2
eZB27f7cD3CYIcQfeZoghci0pNpDL6h8DS25NaDkAY/ikwhxo+Cgf1dofpPpzCqa
yMnrnu4Xy8LuymUBVQ5gT9fPXxlAUom5ngZP4vGLk920wQL0OmFzmgf2TSGQf+KQ
abJQc7PbOdDwGFS5AstWa1O9PpNrd+R66YxETTGfRD6rFTQ9U6CV/6OwsMV53uxJ
Yd36n9rggYBZMIZU5FHtLmdrlRZ7HnaLk9Gs97drRnHZlp4v0fM2ay7iizXbSDUV
pTO6pyDxuAxyPFlcaPzF8SayVq/KkA0snkRHOA7iJCF4yjxrk0zKi/2DTB01vIWp
m28/HtRcfeWHQW/YXnmYOGBYR53FQOTeSCZXe0Ke32fcbhcUZfozqM6AD9CSlryw
lJidwInUlG/KvKEkvtRuQgMrpfUcUlWj5OwJO0bJi+MToSjJHqLTy5n9vXSKwWIb
C+1ykNe8wHWuVjoNqSuKgSCTH10qk5bng1ys8OESCALxAGiaUnyWBRFWGNMsOS3M
msLu3jcVerPRtQgyOJ9DTc6fv1bjlK/cpL+teucrPmsdmLFlSMYgTLO2VHAGsqqQ
PLpmRlg0Mgujo87d1BdVODZ1EI5/V81PHk5cV8GMuxAsN79GcC1tM3xyI3zUC3Tx
p8/1X0vZh6ZSiLWpnKKAk/k6viOhZ/TowLITK/bqNqSJPgIzRxWrMZgH/Xgd5fZC
oziJNtcaj8N7G/2/4tau4GOsC3ewdC2HgogEWmZMk5GW8iGd1o9g8uAWvrN2U8Os
ECVBYeonzyUGjdLP7pCOZeYml9L5EDp5R4QsqVaZfUOk17Xt9RyjX86YhMWq+0Lr
iA1Ellu6Gli9zgWecuH9hThSLnQlj0+lg6xg2DB5IVYM7KqrfWwV0eV6LSFAL8SS
BPjpHL2c6JRvordtthlBD6Ai4Ds4w8knTEI0oCgxpg5qeiC/w/Vbn+1oUaSMhWQM
TAqs+L6YoVLrJQcyfa4Y5wUPQHTHnx48U9rcVAzeFq7YN/lMFiKevwZorbZ7w5Zt
EYBQjvqqcg00CjIWSvMI0VjnnKHKVTa2Isz2bvIJ4LJ3YAYX5bmMfA5H63v5VkdV
+9Ui6+MPbA6hgXd4K+mvvGvO10isyM1Q4DjZDzUBymblOHTSw8ASwhIcDxHsID9k
V/sCfWjeEXzQm2rwsBgy75LOlYtfk6H5K+FUIOiUa7aMHxNMdQqaCL6HFMj+dDGn
HIIiCtK2vtOoYpfU0XGwwp3E+3YetZvh9M3qJ+7yy/j16h87Xfbw1daylIuzzkQP
jO0qpOaodPlftYwbjwW+s96WHLynO6uxhwWw96r6zJzdA+5mkSdkNnTxd1mKgkND
fdTqIRMotr7J68Wol6SyEQezllhmCFzCuAPK3EwSeWkkWhFsuOW3MVZmal2ukFTd
CeS9v695u5W81YpnodRiW0Tptt3pjtqxWNbge0/quO1ZHQOFEzbd6NEPKmRIGTmP
NM7cezY2kOaJoP//tuvpN/MUiUajfnNvMiSNZmm7sfZPljPR5iaO5tC3rU+Hi3ob
GmsvWOVTEHQgLSDeFmnH8ITcM7t5puua2mb0u5Tq2uhspVSNaFl0GApmP6o3zqkn
6L8BmxE3CWX/1V2GGmnzFqH2RwZd3yzdJXHnqx6fgButTDSHSKxMiFlJt4p+knTk
zB/G3PhotNSEboYVjJe86Tw/Z9MjcpK64iRnXwtmd0zwYGknbWwOnZP/WKYH66Ve
ZrpHkcYZfs+SUA5CzH0EgHet5k4XZX+QttgjN8V5R39OV20EzWTObQEXPA3FPnO9
TzlLFowosvNPBfZdpyWO4mwZgWaqBOCdOh/n3hT81yo6sN043XfPM25HmeB456Ag
o6zYkizcNQY2ScRMGWZqAJqLAhxFc8I8Ze01zO58EvHNm5RJN00MSw6+VWFE1CAn
oHYnhww7DN7hA0dOnCgVOqrNYfVQG2kZ3EllgvtivtvDkq+sEX4W3zDfqPXS/lOK
TCm9iX61WCmR/pbdzq7L4lFrjjVkl5LXxdmSdIzoV9A2ScMun35xfSk/zL8Cxieh
fznNXdIZcaeLNBrJzxiN0Fylv9hpJJR7/hGRfZQq3f6hFUzq87cLFrRdXuHK74c1
4gcVeeNTg1Kkh8I+JPPPHpxOnIPJrH6ye1BsK0BmKwGtHfceMTn7QS8dMbGk3MI4
X7LpAdPdPL/PX7yESpYAz5qiyChhzIO9qJ+VqlkvPsEmD/diPb32FbGFLqjPKD7f
H5vFcc0GUn7rgNiNLbAGOxR8+AdXJQJx2UG2OQp/61KxU9UwSXQt/kCiQxxx7AtP
DagcfzqHXlglfD3/GaFObUazT/kpA1JoUA2uvf4DYp6GQVt7TeSVKVBVn0MaPsaO
NeFwYiglwWzVro/Peia5Krn6q6OkcXQ4IB2MYf3E3t5mKJzsMhDM1zo6/C4LFfHK
ce/zNsNDI/BzdNk213BLRpL4fXt5myuU65+Bc9ABKPkbPSgzMtHFoimT1ylzY8X8
OQW8lVIpDDtSmCg0SjtJmM5eQ1IamfRXAG4FAZDflVvZkIg7/IvB58QKeKQg1Ahv
QsXbPJ2EI43jW5uHbvJX2UKYkjj+RstHskN7k0bDJ6lVAVvSyYNDluskOsHgNHQt
+G4ln0e7COR9clgwuhH6O2BGYjtHJK4+tMaWkgfYawwZK2253wi/ePmHZutgwmsp
gf5Pa07k0lsifPbE5kPwKGZz9e3wHA72/dPPjQYxGLy6u4o6P+CSwKOQ+otjFpBF
xmX5qzMUnKb0M000kRgZVd6W5tYe3ajYzbmlsRWjHyoXxtVxlkcfRXJ4D2+Dnbvm
NcO1SARFleC9Af8RSQqf9dIlrRunKw0ozk2nBLNBfTwdkMykIaMSzRp2eG3IGlyE
4ZLaqz4bjsMkhgEvFzESbx9p449wGXR3gIPXywbZ3QButFvs709OUSfGAVH9jOZp
Qvz9DTJtYxcyI9oFVtyzS1CiO2wXMsRX5uNquSjkzDZllO/zvS3Grc2VB4X6c9Pw
d84HzLyUVJdKWi26fFoGN8qT3SO3bXtCFI40uyH/fjy6zWqKLd2AhqSLG8tduSKs
Kyq768xcNFjSxvKAyl/G7ZSuvDzorOkfXS8sPGPwM1sVZxjo5b36EMaxtbo+OvPe
IFpXwEOD8/ndn+5efWbgvVuKPdX/0ZF6BfywbrLaE0EjgYe8DwE3nCBz0eUIwY4x
Kccixi+2aiQr139weOKhLD/QuGwARKiaG1XGu6IUjs8povtmwMVILW0P+Rv3r83g
w9iZbfYNwe2sWdopimHFO3Aoly6LdNLVQwpm6t8B/mEMSjUezirtufXVyr1ndZvv
lXKxRka/Tv3teqEdk8eODbLnWSmpceNr6RKaF+F65EW86vP8su2LJ/O7GAv8csFu
9lMerhuV5gcdLrznuN5dJev2tVUIv/g6w5rXn2FMo67Qr33mk6xWOOlZ6rzRWoVt
TaaeFwTSczln4IdSJDSlH/wigTUSPq6H1J8Pd7VnTYa9hWVDyAADtRJNsc9Kbe8J
cLRu0Wgr5Ob4Bg7TX5wrQ6wTX06aJ32iaGBq20HZYfn9Msn5lTTFFi/cQ1fGc9cz
mV++neLnjYYX3GPu65bJaguuwlQEDVgRMVNG1074WXdzh3W1kTeBLvJ9NL2ceRxk
mWDQwDryH5kBik9ufUdf9sCNPLxo8FgbBA1GJTtWJ70x9RcoksrK3Cs+IXvwcWUN
A9VEzOk5K2v8uLfJiQnlAChObnVHpihGjZilxOK954zA7hCN4tM5YhD18zxuHreJ
dWevNzCf/ZqM0bho5aazQlcrKO/86HPBwchKTNQvLUNVHrszdJUEkPXodIDDIuKH
PA5B5PdQDvwkL1uXqrsKNR51j2A1rs3/dOBw6UH6Ugcl1+yDNrQExIFQbxoeAvUL
/qLrHahhfSljMKoGuETmXihLihJf78FlhclD8XmtEqXINq14xf7YYcM9Vjw86vn0
YXanG5TP1cjaNJhU2gkaa8J6rH7o1KiAkKAKB5DvJvoCtvboOmnXZ9vkv4uY8w40
69KguQoy7kHsbvAdgnTFINqvIgXBVyh+b9MRDAF1GfYM2K23Dspx8aUVOmUrm1QZ
OXKrjMqawaapc7qfeH6/HjtLxjCFrJb7ipwefN04rE+bik42Laenz9VLzRqVu//p
Qec26FHq+owdnLazRGTrz+H7SsLwzfhp+xSQaDW63dzpm35aLFw3Vazy/6+LRNjc
swL3cGauS2yb8En40uMJyfccYcm9cYvvYR+VK+cuTzu/UD7s/HSxl5mGdTrRU2Pb
djVA8Flrnu56J6ME8jgiazIIZZWhTp2tPgDbqYmFJZp3ohsIz7ojhcXbU9nRiPd1
Me4Pn8++PQsWv4Dj0c9Sch5QO/Pgih1r49gnHyTg2hh6djnPxjICj+fjUWF82L0T
d9wijLMtIsej3C06bidmasw+Fx5cOw8s/n4lRl3gI42syKd+BTSQsZbt+crjW9eR
IeudGAwOGkbq4dyrAOUWVmaUFYEgVTa/wu5DKoFzxrJMaWhrtvEzYCsJZAtQ9nmm
BrCeTE5fpOJJhY4LC2G67Qi1x0YL83BTjDPZBl77dEHlrb5lMetrGdVGNUfZKsgx
NO8UhmDWoyUq0CB4jgYyjCN7xCZlmwR2nEY3FUeUrm7OmZczZhknV1zZ5haU1rDT
N/wOkkEcF4TxM4xoDxjCB0Xp8GY7F53SrCKQFod2+cnR8rduufXGUBXLaaKpuhH1
b4a0cqKJM87dHIftXvOGxh+CclAMHQ9o3KidjP1MMQO7JPg39apCmhIpCkzi1U4r
yZcrkpuX5Ajeit8do05BOaGFToeb2BmgYbyBRCFIrNEQlFiQvI3x/4ri3/7wqIAy
pvcYbPyl/rmufinI9tZsBBVOt6WDv7f43f6DOBKXpyQfVTkZqr+Wo+PSVAzW571M
O1PzRVjn533tDZB29lhNgKEM68UcF9XDSDtCWSt+VAtI8xPr57F7xhY5GJtre9Ch
RCbhqeggj9IuGHc5aJrXu5xFbxkNplYnUVPS3jWLiIeMLM3lakIdmjZ9VM1wfX8N
LWtgMAQpcUff3IsqY5rQMlrtoRC+GRGeBLGy7TiAcdUJ1Ka7pC3/T5xhPrZNF9Qa
yM6ZWu2bZM2jsVclekIiaVh0EChUNZW9hPweB2viWFkXV0lr4MakEvjpRq2BHTKX
lUau8R0HyniBC3PqhKppkdPQezPN1u+fobxzR53QpRGLe4eNYCfwSS+7DuGDQCFn
XymM13pTQFIG064QoI8DcvwJIwGsYRuUEF1lE29bQLRRE0NFHREf2zvxo6Dem1Xt
ph1c3qIxLz6qNib5bzDkQdsz8hB3xJRPPB7KZFBk68h/HYqnFxDkJT9KxqVye4OA
RCEMNN0T38kpsmZ6YybLpVn48t3jTlZj8WNh2CO7xZjIFDBSbMnhYR9hZQ+Aj3Et
CeZHt+HfN+v6fFUuZEGGEOegebGByTTQL9/H+H9XkRqaAl6Edthk/vStq6ap6rW3
sLPt3i7lnO77LR05GrMSjWJaUUMzftLqI533sJ280oR4oATj0b6LvhVlGBf6v0Dc
0TqyMGUeAN2OZZKJA3YOREpnHSsoYAV+FD0Ynq8nKbpT5ulL2my9FdUjr4KI9qbk
MBYPN9A3ROjhp6GO66XQJSq9XdEzcVgpT9T8gB/M1zv8pj3wuXVt5vWuzD0ZjUjE
NUKEFid4UZa7+jCaNSN/ag/Jk+tpbssiGPAxoDq9lxDyc7OcACZMNVaMsxz05HcM
9vPFQahfnf2ZllNvMvJ7tln2SoYK349TEq3E3ouxlAGz5ZpA+jjfYsZe/3AnLklu
7mHl81li+ObjGOR5rGPJ7zr+poKVCUT9ZjxAwGVrXUZp5OhXTQcBQ5+t3q7Cz2Mp
PLnUpUX3DJyBqTWddydJQEGq96EgFZN98lDuEF61r2tKV4IIUSN4cCz4taIwfk+5
IOrCP0oK0ER20SE94Pd5iHbncRZAJ/bE7ykeoPgrbyrfMntX/5U5vafPtYK5HQ6a
Y5Bt6O4TKnyBh7scSDSPPDcIo0l8hLML4u1Wo6ysYQA2jvnWqGOz/YNhlPyVzEsy
8B3Tkq4uUApglOwj/14DCk7xW7ajZ+S6BUETUv8HKG2J+ABiYElgQUx5ULkyr5NZ
PdMQmeBdH2i5dCbBePRdzTVC6sPp5OdvJdPzrBWD131rx8QB/YoXcI3EXCBh01/v
OWyrXslzQZ+Fqjw8tzLFn6Zvcctq7QkLRvxg7r0+gijVo7AJRDuHNmo/wEDb8rN+
6+cIJNmrqdq9UZX4grL1bMtpSHNETN+j1JCs3QdnzI3m422TMvT8eELDoCrlwvgx
5B/rqgn+b8GpW7agnEolCgLNuFuYJyv7ugzNrgnX8kIdMqO3eVEBrvSWkV7dKIE+
GFDs/hmLDFJ/SEFrgkBZ33G2LcE1itMUsZq8dQkJeIGUcezRoo+xyadYRhiUnaMd
btFXx00m1OVon3EY+0ti+yE2v1DbW9T2pzSlpV3+yFdykxWXFU4qjW+TzcsCqhkR
hWU/s39UgobCre6rKZrOWoBhOMBfioznPBb0nyoTvh2bS8XFCXx7nyI3Kx+83Hsa
INU0Jw9uiEZ3gKx+dRtfHDwS5fUPj2f4d+pJ7GiPVks4XAT/QkrsR8wcFTOKQWx0
K7d1MHOun0K2+sZ37itwcUb7weO+SVUroeRKWJ7U1+P5JlVY9dji3lfefKLbiBYe
6T3S0DqVnRaAWj3daWTvQHKcfjDp8rj6Qn0EcFq0yh8sZcfACGdHuD5MHO311jkp
R++KETlk3H997jrk4HCRUGTqwlxHVAOyL6BLmgRBdb3hy5ajYdTUwVHC7y0mNmWB
VOR27BhI5VoNsaZOFjASL1d1Tip6xFsiuBZdkGrkeE2/pA3Cn3/t6GTpCkvYtGPO
y80JTl49EHPaMGJd9t+STTBH7Srnts24S5cE9VuJ+R0selC9TCkhndKNQGyAo+6V
ppu0ub9jEZW19NgEEMiGGZhhdTS/yTOxUHJiTU4NgymgElggrvxRfZgyMkHiUi0y
Ds831wNnvkbrirejVuzlk9XS8EzKqmT9weqmRX3rg5Ltg3aWmvJN7vq3BNX55ByE
9XbeM+nahB2figqS0kLvQFYZYCYdBpdAlAo3kI29//XVUYtWSmar6zht/UNd6PjL
sXfREm2DSwUfPM6k52/GImsx6GSuNWg+ZOTH1WYnzAJ8myio1pQkNsP9130j3uP2
wbH2ktk+cK/5pldLLlXe46OseE3bK1i2w22Y6RYdlLSK6r4D08/uttv5SOvTO6vQ
UT3c2MVpS6OcVJdZHMDR6+IHAYWhhmnWQnPDbKVohjxJWBOlegIW9b5Ay74vGgIz
IsCk69hUg3G2cPTlcchsPGfVxtwDZaoBGW1Ol0wlKm6kAI1SWNHw0xW3P9trQcEn
2fcZ9E8DmiU3j8f1Ls5ulHNXf5CcJrHh7GDR7tWuS4w2ONpkZuzA8SWvL9W3CZkK
JfMXP6RY4N/5899DzBF25ekKv5GyeQlcHi1pRy+AoCoHL6H86PHbT+IOf5cu6P7J
nfeHRBBF40IgNDRv7PJ9sA1bM6a2X959gGHx5JzB/B3vNd6nh3tUxwB14oK1wuiu
CzrotG/RkeXXggE21HAElax0/1bJXm4xxrEMatYKcNpP6BsPD8eJhnvaFNaYurzt
BKicaVOaUniNUYg7Hy0LeSPP2hDLJrxOx0rPi4Mj55gQAYhoYKzx4ydAojoZCvUN
Hf92dICM8uS7c4IRxnhOeyYfUmShv34GF8cLg7OEEQQdEe80jh9j6lnXV17JzLif
3n2q6C0e6T/VauZUO3xTHFc5uqE8ZGXxc7kPhN7VKx6aMjFCUj+GskCMx8OC6CDA
g7/Bzk8gLR8PqhN8O0Szlz1dFVZZMaydAnlrO9MEKfK9NSQF37r6xm58ZJRtqdny
V/SZEb4ghpASUPypbPjk2NwnhWeGcN4pn/o6MHzCCGgKaCSOXUL97mekXlDreguM
B1ATkGX5Ukes93KA8Bkw/wYfclFBkampAm21TDJkeHIpK3PshrvsgBTLndm2kOgQ
RcKyvu476IitSv32NnHtkXaVtCmEFJsUdd7xlZ5JhzLfFFg9Ltjw/9FxZ0BUCfjw
JcBx2OvRxzw0Uj6FygHb6t8ezzG5VuQ3fm47hl3CO2hr6A5Z48EGi3EENDeeuQuY
2kGND+VFH5Amz/LrhamrU57iZjv5FWiPkxqsYzgkX2EJEI1UAGU8sXvIh9U5rxQZ
pQ6W+bUJmBqmEdTv9KyTH7Xl/KJj3gFqiDSfQmn2PTEeErQZElASU3P7dAWqaU+E
DiVJnWZMHi9HG3ZOAzB4JSeK6sPD+M3yYKsLkhVGtK3oPaMJ8+EIhTd/GTrmFCi5
64ufYXHBfAa75AGZI0r2QUryNThvgKfUn8zBwS0pi6MNf6gxv95TYhL6FGe0c637
ROZ2S5DzuYRxfNLDfYLC54boNmTDHgX6uOivkPeFG+S4DC1XB6dejYiBTkm+wmzw
NV8/Z0T75h9wguh2HW6O/shuWURDxLGXWxUxgTFC+GLKqoISHmIgjNjgjhO2bi4Q
nQPTYoGRnZHndwoqO1gUieguSh+6wsfzgrAIFPzVFs9WmW6/cYjPLQR7J+216p03
3XiWUUZHaI5nXL3Sj4jejjrtbbXireyapBdME0FcckERS3gyxbIA4FpgG79269gV
LDnUcXPcVPlA4j0Ti+u6RFNfySmo4nENcQc1QEbJyJDv2j5avToR3koaFOYy9gBJ
yp70N9gr3mg8GfjnTBSLclODJIJU0Wv9Lr/sBPtaj9o8QpULz/Yf1j/HHEC+3ECz
sIJGnnIPDr8Itk5rhKsm3J0OCv3/CQ5tqbYwVnXvLlFHRyeayO6FBuFQgm5dUGvn
QOgoV+yfO1e5cVkhPR16JIXK59Ii8G6E69WltTWJAp0EsrgsUpltaRzHdjsDsDic
AKf+3wuOOsCj7AQAuV4S7JeOP5zjDByD20UqEBf+I0jq9HS27Aj3gMRCE5XWDAiP
ECk/gYpDqQvCCYCp4DhAV7g07jOaBstZ3kJ50xqzYkRMCQ2iXWcEtvMoIi1CRzQu
CYWMiFM4xni5SBbV0kPPrH9ZCQpyElzZfCNtUscspBo+fkYIOHqZ3B073fKuks5F
emcUEof1fvrdxSvBO922+1+cJwWGOZfq/Iw0+ypkI3OCKKkqBcui3b70IE8QCu50
WUtD4QX0utWdtICbHtymXJOUZq0IHW4cNswrCjLs1X9WuNKQDapXSnYQYN+hRXpw
dg3RPu+4Jb4IJ36RZ2xtFfhvEbUifDA+PI6rMsMTuiRSyzzLxG1/Zpz5fXfO9fND
b3mNNfakna1xQQkAIhwp5roEW63LqcCO2jFfQY6OsNZAM310Cw5stIGxl5vjJJON
8tpFUIffZz+e9gMdtDx3M8iygYTGeU/Cmp3cGpzkPT8XIfVi8m8ON3ZAnJF+CoMw
EvIcfPD1z0nv8927RWXdJShEkbi5YOdQuGpIZjOjQb01k5qhd8YU4gsaqKDlVDBL
L6W8udJG3y/zXzCYv/bEbf6KUXrD85FwIgq+wXPXUHowJPeJ45zDDihU156eCRhU
/pz3TBWKX67ogtzZoCg6Dj2v9FQHby1LRVL389us9K/NtqaYItSywFG2TPfPT/1G
VwzSLNrTv/RyTXvL5qI9gg2tYqjmrviabcslon5yUMgF5j0LsnqizduJBugVrg1d
qjGBZrmEnetP0BhF3kJ0NEWgwyPO7qKxbZt7uTWdgkzR/6Zr/QN46fkW8G59t61M
vHBj5XapMWhRyYwGnU3tBpTgZyk9lJ5hyCuWUwO4rE6oJLlITKV3mXCtCkfFQGaN
BMmZV1UHskDbxrh8sTJR9EhFiydG1yYmQJqoEUUbeCas+HmPFm0T48FsjVk9jq+u
YYw7O3s5q+NI7aeD9KVFy0tdrW2jLldaLHfwBqTdRGE+cwlmrg1TlnOnb3gZOVDe
7cDYHAbZYpvsDMFND+9lJlT9q6VNZiZq4LcOGUozkdwYNPdQBn5SW20wg0/vZrZv
drCxEQvR4UYd5i+coRX7EH3Hud2FBxGIX5j4czJToP++JnN6b8PBHDBjbIslWbjB
rrcW394n92AoEmO0hAjrAWt5VN8t9BMM7TXOw+Alf+KAVLBTz6/kcZbRKlV4voVZ
jcbK7tCT4aFpn+1h7kTpqoKJDi6ZQbnsIQyam+P/loe0PM80P8mBP7WGKz6tHUSB
d5RDT4vSznPiqzzaRdYhIe+UsFnQWDW5E30bEOJ1GOvLyX33wz8thtWG4s0rlAgU
GtwNzXKpebH/XGWLv1Wex/+mbX2XAljMWHjyDktee6GMn3H8teFK3p3S0Ixq8+yN
jMB7x5AlVDrRfyZay7GDkOjYAR4ea4NDNTHfgtDN6Mho5PFyomVY3itGA+B0FXjo
bx6sHJnU3noLW23HK8sdiuBCewCwJJTLdVyy+NRcyZspyhxMvirFQ/QxPkjZ7hqe
G51YTMI04blHwMfBi+iDw8uOuQ1v+nVVD20PwM/+4TbUwHLInbcznFzwgyv8/hGn
IMS2t5SsUYj18A7ueWRJHTXpBTx4V2QgXAjdY5rEQEXWAlVvFUAjXuWttozfmWe3
0+pj0btcRsUiwUvQnS/mueJpmJs6Z4cNlnXCnHnuUm/7jfVoftWIDOaezm0hiaBH
VmGxY+lQ/DZpNKEwVg2iT+XlfryUDvl7JbDPuY4pB1V3OX1hIAq04+/2J29FF05D
bvR2ID+MTbbRJt1Wh9EEracn2HY4ilA6eqgoiBhCzhITKS/wcw+dHghqdajyGRPc
jjhHKCceMl0Ps8xowwnDBg6DFEQeIOMc+7uuUyEB9mqQ5rL+Lf8pC6n9zI9SdElX
utiDRnmP/Mt2PwUl1p+Ul+caGdj6eVFtATF3woZp/hCXgokCRf1M/MiCj1RplT3w
nvYLtZ23CA4jqMmjP+dFHCG+9Dciyg/3p6psZZojkKkkmsZa9mVNJuLoBO2yDiXC
+CgRhQ/ntMIqoYfqtD4YVdI8mE+6CQj85ZmCK+ss+i4H9W8BYApIT6K7geJlgu9P
xjTRQwMaywpzcKNNpzlCM/+4SK3yUK2SVxMMrVuFHB+YlU3MLm8MLDn9fFERtC0y
7x1GFRZuLR6hKCmD8ZoGwbrqGikOPaoucmfU1q8kEuqDjUpxElre90eejMjbOLjR
kji/799uuTBTqmBHwMjJU4Ewj4iwe52tSvd9SobJu3JnWmWbxs1ii0/mtF5oRpGp
FskNIg+Usk9EIkuVuTDqXkYas1HQr4LlfVjvwsu3kXfx/6wumedMsLYGTbiCBcOw
NhlizCwNBPjuVMSfghFDyG+QeSHaYvSQLRa5uBS95Nm4NJo/7Id/GnHwwj7rBPv9
L2fKN+SdH1i6d73Xi2LB9s6pnWdYH1Wa3E9ATeyKVeVgw08paFaa7mPyXdsmo3rp
cFu6DebUTeabFeSPwAdfoizrbMjbHjS6y95zHBeas+15RRG7Mu8iOzWHEoT9HyE+
H+PfIIUf/IittZsUpOkAeggqBB15P1maeAoD/SQxE7yKbGyFVNmJ4VzKH7KhCpko
3kwfEm3HVg/pCuyX+r2FFV6fUAt5u/mx7u/c4Ek+k2jf3LajkQpy78JSuO3xcAqK
8mOJ4MgvH/9AwIB4rFWt6Q9AIroEifySCuCbXqpVRKIQOowmAFLjahco7Zx8BWbq
5rshZJQLlhwc2Nvw8rydg0ccXExyzu8aQ1ycnL0qvQ1zOigAYTRGtvrLvPNQ6wQM
Qo5PjX0slsUa2snF1yvvTE1RjqOXZ/ayOXFplWfQpWJBEi94LyCR2C9Q9RNj0H3V
ku2ZPPmbE1nNY9S26jkQp7T2brr0PntPD9Pf3KCKNDwW3xUIR0hfu8ut+FxDYN73
DKFFSoYDtSHUgL16bIObw/LK2Vd0jPDAVXJMNk81Lav0ujAXzeAUOM6VNzWAV3sj
y5A2YrA/wFEO5q/zuw4o2y8lVTKAtTnEpuqvFWWxC/i2HDB8j8jnflVOXR0OMs3E
M74HTiYzYEIqFW5lGNm7Pt3ZzsQO8T+2/dWiqO7+Pz0fkMK0NaVhAQGg1bdSiAlL
Eb0JKTkAVZVSGt8SzNtoPMRLkMNnzqlhuafp+AjoxXnycAvfxZoSk+3i/4Ta8CgY
JJKDcjjy18t8YoxpJbE8W4JoN5Y8DQ+EDZkjQw+HNz0Bskh+M+WhM7MVdHYDoa7m
hUp/FBoF4uCexF9TR0v6MQIjFfa3VZ8DZeeH3Ne6UdO8R+n1jTa4JoOpZjuS9OaN
aB+06tApVO/uSImWUSOzG9CTeHnTGeu7Q7YPz+cOLyx5NSRAaKRRPaH2I8sB+7X1
K/yslF0Hw8HlKTFBGPkFIWKYsYQzQowgDSDmro8bShk+pYFSaH0XbNv/B2NUcChF
YALMrKYWZHUm3anyaCzvKeznu1mnNUUBczvMNRJ/GfdENVTSI8RY4UitpVXYK7aN
ElakHmeNICe/sUqPN3o29t8ewV2b/UJm/AeR4NI3TFMrMaXh86GyMTPaBz0le6t2
PCGWobUZ7lQ27M3i65ztp1BgCrkki3iliRrdd1Lj7PDohGIWjIB8w7Tlb92t5fAt
IzOPKvB62GVDAbuU17/hH4RIRAAC3hTdm0+/NcStkIeMFgwyh8heXRTWjungWaN7
6XmoMc81HIXWia0SPInjzhULb6sLnr7MZWV050ZfRFktytIDx7hspK1+0mq5liIF
z9wyjNOajaA2/05ZMcc9vjJPDp83DNkzY1ccpYl0JEDayAD2grA9v4pXNmqo1cgx
vi3zcJ6rVXBipc3Xk8xyslQv9/kMKiI85iCfLVnhe9dms3LU0f6gMA714HdV4EyH
YjGwBMX11KIpD0y0Op7rmZkKYQ0t2llwzCjU7ulSIimIqdfZsceSCVqCGMyTcYHK
hZNnDXHdvW2w2YC+TJPZZRd8lWl4PMJo9JBmLmlrd76FGnivn86TVgYvjVV2Rtfd
Pp4dc7AwLPUqs9wQCcluXKD12QXSz2G0tUNAnTL+KuISXIExra885QZ8AxRH5UFg
3XlvdX6P3pjI5m9X4++jLVXissKtAs0awc3/B5cgSnshvmKltWZXRbnE45GGnn3m
mjbqesT8Kur/e1ywZ9t8yFg7QELbmOXvFdmMvajo3V+ZK7sgy80GGo6mupL1Snu1
NvRaq1sxF2wvcV3fsw+r2tRlh+6M8hD7rHO79J3kUYtPAPe6cCZtAd0k+zDvt91q
kErTlFXPsRhXEkoThcWixG7E4OnUEXB/Th76KPH6+9c5vTlorYvbcz3K66x1JRTS
RKwm64cWcVxaAk4shLCdmufeZOX4S0iPC+dowHUqa6Gln0qvZx7opSMHgo0C1CMU
eoRpy1MdHJwN7VcLy4LirAZsS30sAQjMkfakm43MlOpfl9sYrhq+9z0rKintP7ww
BlCer67oLZzfNGonlZbjbyvQuIN/1iSyVWyzsoQDV/FTUUIsoFLyov3/n3DNN4kn
xxlPmqCvFeGdaCaZ62s2mv2K7tBZcPJ62JJ3Qyn2GuTVBu3tky3bPPL/laVX9AKY
0NZssC5Ou2R+Tb+eE6rahLT0uYqR3AoHdR/GpempxrJXq9bZVt7OlhGVs7ZPjwmM
YpeQ7c/ifrWteHOsdVR4jwSi8UtTiLbvvmIDLU027PINti8Lly/pqxl0de+puKnH
ZhuR/PG4xBSo3CYfkmsURpDVRWXX/JY6EbWZPuRJu8w3MjXlaQjdDs2WRwKDC4xr
v9lLFJlEAHSpr7Buduh6B5ZN2SUvKsp5x17mkmoc3duscGl4iSNC6sJDPx7DJXAd
inddNdXNDTeZ3dSNbNEPAp7/w421AbQCd4//fDPuopgof+lpk9zE6P4tWgSrQpcx
X1gRoP2dC/eOsVOK/VJknjYqku78wDDvuemN4Tj0WUp39HPB6br7t8TFBGQr378y
X4g2Du32CCl3itmVn1xf4EC1upp+LQsTO8E8iGpRckuCLlXyydesUjTZTAyZuAaT
FxS/Ed4C18VmcetukzZCyrxZu6G2Y2q2f4VxaUAv0SgViukTp411465JIAZwgk2Q
B2rOaG/PnWcnfdX1Z3XXfEfuOqZWP8ATcVtMABWo6tCTPWC2gqgnfmEWqEg9s8Of
CPjQjHdlxzWxH9kTW+Gs5LQuzmOQcYKdLPl6P8OtE8dTMjKw+V3CwHHfB3g0rorR
RiAarv8bXx7LkH3z8UR+LYyDZtd/mypHLpHpsXh1MyNaGz/cpDMu5cQ9NMzNcfa5
/F5TUSWjJlieYYoY17JYXzqULNTRTE+v0nLP5NxUAMz0ngOyXHWBb176o7quzd4X
H+qnYT9mM8MXtkXd2HwHoh9vNr7IVs/GMFKvqSbHvyx/7s2PBqYILhpkFq5DRsKn
waQeXmxsg1M4pISSLHCKEY8+LdFWR9Fzh11JzK92jTvtieV1gzMd2ZZLf+NjbxwI
urJcwUTrPODKd3XXhhKGfVZV5/EYgr82dwPiU+OUf0gHEtnFmHkKe8jPRZE9d6Ul
vlP+us4WdZOQyWItM38F2kwd1/87Pdf8YRvBUy8pu4sWbYLCQ0qmxB8je0t4h+k+
Vw1xnav0gUGRkqFiA5gTmq0oiJzovC0x668rWG/34/hHyWn93q22+Hc5DHJ3S6s7
6AIVKTekMGYkCxVAe7elxqgmUgvM0g5KN0PURAgNbtE27ZkTMZJtqpXOtBFn46XE
fbH0H37T/o/ipf68Jw8z1lde5WmBbRjdTbba+4dUornedayqedpb3WsL2EuGRtGX
KGqOAUPFyNUZNDx10iUY8Y+9ExxAvGfo2Yg/UaLsZLJX+uRgNgPqPB4APLRWkxFu
FmgSK6oofZ8ox32Q3qfkzL8w4dieooN2BAkITA2rbOgHuN5iizq+n53yP1h4jKKG
bQ7M4k2R2k9nNK9PoWHR+PUyBLS/xxZA02Y/Bw6NjolJ0hoJ044K+7rgWX5B5RRx
y990XpsN/YynXoC1FKVlPsxlSs9VCmvfkQndKVlXnOVnQLNU5Z90McuaFgi6NvVA
6W+kgBL/YqOJF26PIksyruXxeZJLHzctc7ci3y0HukP/KFq0rKwY+lSjXbFow9Kt
UDSZYTRvcfYMUe5psQe9pzV0VLMf3tHWbzc/i8ZXRlopCngJs5GpT/wjbKhx4JZQ
64Vft8DiGbQQkWc6csP+7E7ouRid2FxznwZpP38vcZLZMR0MpJtRj76wgSOsqjfk
kYErVBGb5K671JaGlOKpVYUnOk/Ox0ie0ceeLAGVQeaMegdYd5/fy7NEtcifZJqU
BcFgnVmAwGS9wZO7GjjhO2sCqPhNMhoHzeAAhc2LCN/Bba3WRnDIFRUmyxcUJrUw
/NQUTt9pgka5KISsRXPU82KPtIcONH+06g8EM5hrIUZIFmtyq3ftW4xuWWSFEGyg
PZVfpIcL1QkytEvH8oKCf+OCK9CbTYJc743lym8vxd93Ag+ZwPY36QHxzvCBG2ER
5Fl6u0Cy555M9i2H2qw6uM22bDUwwym1KbaDdGtRs2XwuHqO4DMpwoQVEBCGsAlh
8dLV6SG2WGc87M9mj+6iBsg28GjfivRcu1O6TsBzmpVjByMrO5ZQqLkPGpfWH9P4
WqeIGkfBKBbAFkuXS4hWgOBeh+Ghr7ZzrotJFnjN54tyk9aiWbYIaxyg1/gb2DGp
eGrp59yASgE1zQs0yt9m10q+BoHgTp6tD2jzKajZkPDNLuYLHg8f3cuggI0Ir7Z+
xcRnIPwT/hgwfday3COxHVKAQFCXj72sp48mx32AX0m7Us1tX5RDJtEss48pf+if
XHOzUhMpEUkolf7iaHGjYWUdlu/j/5YgmqAkJf7QDC1tFaC6Qo9juzZ2MIVFKPsE
6Kt3tLcoZZVSedrHVbhUWOxuc9o0Y1RS+mATOWOKHx17pKe+xZaoWyjcj9nlgGyk
txwXQou9V9El03gu8SKjV5AsMEy0to6FuB0AM5vMUQUPeZnCRUTCDitSNbOm8fl3
l3zWkID8hl4R3r0d71SBE71YefFOrrR6Mk18UmDmubIKToMBdWETaqI2KncndSIL
GO1ezg9UN8TAWiX1/jxjAgUpTNZEfLoca255OaZZiTkzaBaqCN8dpElzw+iW/0Ye
b202m3/nMbJN3Qa2jE0TbJwJB/nOO4roWZJoG7WwIEodzDvwI0E9qiqIF7Y/L+2H
7zyGAvKFwkyWZ4aEIF6TnWfN4UAwx6Zd/Zxc32z4qxi8xZKgwVRjDZ7Y5xS9tfWx
xD/OfBBJ94d/EuF0p0KVb9K6qn/gnLywStmdOsza7Hu8iUplmAQ2BGtiyIX2qyXp
41jg0SFa3oJGqbGwOB9XDz7U54S7B6jzUypzU+1O/qBJJoFO08ER5ssVFmi+OfxS
ruHdSx0vSoVLg1eDF1yFSU9dLBOT9BTTRWmHL8GRVFOB2LdrA7qT6NDkY6HT+mZC
X0bUMbFL+dkGr0Ak2n8TBWwJ80uEFE7/+ObuGNabv1/jmtqybn6bALa/i4mnbv5L
E0Xd4UF7hLuEl1pGKL5OQCYyGBmkIWoSlTIe875W7nfQSIbVnd+jhTN9AiZflGcM
4YvKju6u/8HG2uu9F/V8kQdRHToJaO7fZla8cotNFwVTENuMJb3EMxGc94LJNjr8
NN/CF8sz9N27BmQRo+VfnD9ycVop1FWl2aOhU++1Js+yWk+7Wc0x4vh9+c9nK9uG
a8ei/fqHt3fZeJqf7iI+PYOVaL+43AaVlwcuBMA+gMNjm1v/60wzcNsYyZw+6YUs
GXN2opHJVA/CpBv0nxhmt/zHZMQMkd7NsUqfLsJdC8x/d7dF3f4A+Pl+lb9kTYY2
SrDwt4SDS9vo2VifK5UE1nWlHm7vr1f9HIMbBH+A7kcA1vX5zXYkJRw9FE/DNDbK
GmBJ00zdy3l2hyfxjSzBpvGsE3XCabricB80wGYI4F9iEiM8vOQJGWjx8e0lrNbZ
zvNvjwIRQsBb9mPehlmO0YYigdf5w7kqlaFenttubIBb5O7MTIxgSKDKEXMwHDBx
drmd/8P/RnkbGB+YNkoJbLmdYVuBTg4Wa+SyvsvbShPTWJZtx2VgyQSxVGhjitDm
jxOAzC8FLJO5zuqSTqXNCPA2ee7ozQSDRQjSmtUn8IfCEVuA6BoI4QI82eDuzzJv
C9S5BicYXEFlj6kgigEV+3Nj+BcdLsa0VlHXkrfs6BALYJAG7n5h4vuQtw2VF0Me
khfSUTF8XNGUu65STfL7vTcmx2CYblLK1kQkJsYvx8Ud+ZeaxjE4kekD/VVeR06F
NCR/Gh/jOeK1aKe3w8PxCtL4oK1D6lmxJ1m3r7u1E0wi/TIzRTft+RsAhpmvZ5PP
658K9Y31o3S7sMpX9xOEZWb6JCmgSh6dmDmoBAtUipI68trC9/SIPyNNkiM0uDk8
YwRSl40nyCZNlxSEDnIujvtv6BwTarYCqfabD21cABPsnV19e/SuwkEGlhZ/bp90
JTPXn6aDK0Maz69Ru2kLk09CyIC0cKL0cOLiS6kXK9qxfWhqIwB7teVVyGviiLyg
b77TMsrc7KWTge9IE4t+oA428tcCKBE6WBt2JRMlg8AQbgFaqTTK3SrvrjjuRFrv
cXd1FHNBiM0Q8S1xB9fopPtW/8qd4toe0wAwlnwTuzb7EVqBvzmovqKzHwWC40Dk
VKnvoWXl7G+AeJL8AQIVkFHolUdDuxatHbznWd1sQIadezhQ32KAX068Lldcc9nE
J05OagdERf4qz6+wnXx1lh/OQYPBiis1wOKK6R364Bom5zOt0+l05lfqoV08gupZ
kGXcwah3Q//d+DdyB7Fzvkzr4KHUoPfUAMHN7PUk4RgYQSCA0kfNYnOMPCEnzf75
xfwL757My4RY6PK4KgMMPIfFSKV7xTZs2DzOJW+m+AQikgfxcr47ziQ6NSB+U0nh
yNKfLAsN1oydEP/HUVMtNcUcOSqAyNB+Yy25CHBskAjGiywCCB3dAm8v0VrwAJP6
ZR/ZVFB0NuNBt9rVIkd6S5a8xyxlskBLI0Qr4Mbf6bItfqZ0aZVi6Ez4UA4xiXtc
j/lpjYmNVyq+AvxcpS6J6ZbzuZaV6SrpJVNBwJ0TAHHZvKLH4rZdpB0DSlkZ6XHs
rnA0PpqoRBWH8+LrQKbobBbOKFvMLvXqliuhGl/Y6ykgk3Bvgk+Zy9MOrFlVZXKl
4eqhGYPrJwayaxNEMuT+D0atUpLnQRmKBaQ/dmjikNJcxTIOTOiRb/KaY+lsKAkV
iL7cc/0fslEVOdmPAH94bGady2WCslt95py0ul1L5cZ2s5vSWLPWiPYTKHdwO6aM
VlUlJlAKQfdNMkFNB8dwiB370Ks5UKq0o9Km/Xpv5thfAT3Xjk1B/kbUmQYHZddj
cd7tXZ/vRmMXw3GGaAsPFSziRxlfGrh/hOlKVdUNbNw9MB6mtScFe60I3M//wquT
E6VLT5RmTmFmORNw2xQTgEat+QDlnnhQxNqLOUQzjTPBZ6kLhfUnzhnOOALVikKa
1WX61mUqTN7OClvOe4jQtXZhJtqkdolLogvr0MiG5KqnwUFCKrLjxwa79mTyWUs1
eb/pb4FzngQqQbmtSDErKxN+87zELD/Of+Xnr1pfQMoQm8rJdM/Fe4NdmL6SYKDH
fcxGrxaTipCs1PIkvZe6hqb4vWAy57FZnv30Ni2HGk0J1P0KQyIz41Ur0Y9DcIhL
O/6xZj7wT6H3lUVbWkla8gD84aAPZjn6w5V5CgH4oetKG8zLy0wGtG+lND8ImDqt
8j/amqnQZYhrbL34b6ZPxUtDLbSDyKXlbNb0Y8bsoUwjDxS2DjiY6h+RiUotn/+8
NrcfH/5sp5QNNJnDOJfsbb31viMeSAePr3clKn7THd7ryi2z58T3sssGZKtYsi1A
di3ZuxUh53sTxD4hvLewZr8dPYx5JzcBHe+KHVGmRdVFMOSWUMxJrAdQtABViwH+
cb2RYfqbjm6mU5NCa/VME3DaPLd+UXA6MOo75n6md3BEFg7sd9QoV+AuawnLLxX3
sZRhyJKvdVYvuUIelHG0QpcL1QH9DYXUg6M+cJIxBuhzLayCXJsqvflQiLN+wSbp
db+chSUwon/IvSmnwrrPMlS3nwKetW8QNDyQzHaFJBJ1gI2XJLX+iZgq0KCtBezf
j9Lsir0wNKlZYIx6vvkomCcWsKhi1ovSabZJY31XCYYoGpMDZCXiH8NXvHI/BSFo
lsC3EoNA2b1xyLZSuhMa82C6Tnyn3WOEGy8jXguLdEVG9ofAOIN6/QZEXZX/ryap
uJXstwjoAiB3pDMtzCCfDw3TZ+jm/e4encDyuW4bjmmcBHTF4XPiW0po1ZF1NCK2
RtDovVAmRUSwSS3UDklXiXR4cwHENG/S8EY/pVRfBUnezrIaMSFb1FP8qGFfBPgv
G3IEIu62SOIw8MUiLKXU4cEsJBoJTSZzAEQ8rVLAGDsdU4KNXQLKvlDLLGMeP6ky
WURsgG0hOk/j+hbffrVxTh2n83W0WzK0ih29ZBaMZyi3/MiVRNr7My3ehc9bVKZM
+mpBJYF6Ji5r1Ucwr1sEMfMbaw4TZSEkWiuVF3OTOXCjwUHZWLwHyxakqW9jP10c
RVafOQ44hYz7Qum8Gd5lT3ZoI8MRCwfVpfA0LW7sv9sQD1Z0KTsux9yFxs9D9mjS
9IOWArXqnFMU9jRE3PJbvSKvIyWAtQQrjvA7XgLbQqSmNa+ad1mDfVspj+stn5ss
uouO9cXq9xmuS6HO/xhwnRhebGn2XLh8tBZ8Go0w4yDOfUqeRC6/vGmGSbj5W+Lm
l59Q6gTi7d5LL3FFG75XE/F/TvcMFhzJMS+OWZoIMKDH8LmvEYeTm6Oncj7a69Aw
xXuCDm744dI9qDvtp0I7F6Q3c2yhiqtyE4p0i+QeNCBhBRJbY/FvppiNR60hAAeX
FeqAnb0zzm2tSnhwhYiHvLDw/lNWTqgxp5kbb4GfZhKMHiKzOLswOah3/lkG38Fi
kbezxT7+U298e279tsS084U21rVVlYeaLb0FvCFhjLe6MMzteOiUA13UHpzfQ+T+
Hzd+79a8YMY/1tmLxW9rPsFGxpAXgXoj25ubrb3tyVgXSKVtekGkzETd0NYO5FKs
C382EJao/olxPhzYrzlys2tOktSPl/iKRcVYEvUIofsTtAz8sbGDYNz2wQTCuKTD
gER4Z9EhPIfFGvItrLDDHPupzaDETVc9zvieOK5cH/Ow7Xe5xH5u7CumLQYCZQhz
GpBhcoxXU/Yk/kcs3dqN2p9nshfIkqdyvdJ5q2lyubVxHGwpzfMCPqNGdH3B9YQv
TkepOQ8kpWAyFU6dSrAIyB6qQHhTq+UNYNz2NCkaIzSZ1YvE3o51Kgm7aX9VnMCL
umRglHlG2zpWeKofzsBQKViPc2fp5FDq3rlCRxbRoLFHqDeuar3v3KDIkK+dEZ1Q
UudbZjHsyJED3iPScX14kG/WrCEsehy6y7f63A6LD8tkH9y5pbMXj3lYEXqCA5HX
TZZZTvAHXbYMHmfsj31aAEV++vt6ot+IVyKHrOTN2/1MwbcUarbvr1jm7CSknyJG
laUGAGr/2zNAx9m8ydnpOGFuZnLMyUTJAQ/FYJctccr/Dh8kIwemMGtr+j7p6oj3
CinnDL4/fp+zsJ36J3jFIuYo4lEusRki8b1eJqsgmFgVs6lmZZlGGZkFIRvmdw8J
oqEuTH2f4m44pMPUfE18nXm9Kr83YXdWPswNTMMLCCuO0SJsY6O2/PsjM+g6VF4H
lbr9Jm6/7nWaRg0aTOEA0e8W3KsHhbuvR2I2jg06jkpzS+wLwPE6SG/urc8V2rzH
sXeidZ7xDJhqEN9R71HvKHW4LY8UzUqAE7KHFyIIWqw+l5XH+iHUCAARr7UFiLo7
hdiCcEnRirr1E1vlPZfkyYbAtng9Lhjk4t4S+nQl2OpFJaqBnTo89mWUUuezA9n7
r/vZXpo+mlWlTkO+tX5+rTzUWGuI2bpfH95pjitN8esylm3xFRsoHQUgHI6BEH7c
FuOLBPVlBMk2onq9R1lmCqZdRLAwLctuaD1WpQjq4ERZwbxAt9P0QUk6ztq/VZVx
5pjU5f3U6CUlPW1CUQtsiNH+A8xm4JSlu3dxBtaCOtQScAE4bwqMM3sB0qmYiX6J
Hh5FAeC+JsfvoouTDgLeULZ0cOHpqjXqxJ526WUg3hvApBLY5U9wwGpscRMqxPOu
NQcTpvuc2i2Oo4rABEgi1DCGSMtOC0+3W1oJHHnvk3c7lszHvb+pEQ6vSIF5sbXb
+2lr5VW/oQ32ukwQcumN9fSdZ2FHyWPucqJoazicZab2hAoC3TISMCseThYtmQUc
/Dv1nyH4bCf3fjfIQn4gfkxfuyvNqbbVEzSFVLwUsayyFUZpLmSwKimXXa2nIVwa
F8Ef/ZF6mSDn1QP1IUb0b6JQUxWoL6UWBHDIhwwK7R3z1BKF7pKM0U6MKexTozv6
IVv1/dfyK9gHl9rDJN8vmTGrNPUwocvgZK55E53uMOyj3nAu2NT3gb332r69jE1U
XDEFWLOMgZu5BLxB2fbKUB/UCH3OIIi8xzRm+xKS0tAZ2CPpbyTx/6GTlQTFjiDh
Xl7CZHdS4lkA7NPbtMV5IJnBmcVT4rmcpFfkYT+/IW8c62UHynYpidpYowvb9BXG
QTRwTncGyiqWz1jPcW6yO04+w7g5vKKrea+kAuq+1SC/6b/EsU+y7x+OnsEmHmtL
F/wv++PzMfVQ4VIS22azaJgA5yDfPRHBFMZp2o7pcrHr7vYL96vxlWiYaOr7QmIL
nbdxYekk5TUfmFZS9fzXIR6oZj6foywcUfeqbWT88fgdhEaoAnjbnE5JIBpSgy06
2kOaycOjcaLmU2ZPQjeIkWEF2duuz9ztXb2Ojqfhgrq74Ow0EMfzOFnnWRoizzrN
bIq8qpj5JznmE2gMmldSHmGGYYAptdhxEm3q9LE9T1GYWKBK8OjZltINmCRQ1v4f
OckqrTmtWY2Am0HcHedwm4DzySDgD9PsbVA8aOAa2LV9HYolZwiiNG0hO8Xrdg04
0w61fVmHs9pLPpizmoEUgesFz5Ehdkmf3+mzpw3gs5V7j3fa90NPlaZR/VdijVhf
5+ugaZbkL9xM0bjoJ/j8hW5IxZqqsXFBVjybqi71c2FneDu/EYa3rw3XQDtoJFp6
Fw15yLcg5c8JOaJvtZ6CFljiSr6vHgYMYQ738VBxK1eJthQby2mDlw2HU2cB7SKr
hPEh1RhkXgB3UI9BFBnCHyV8zlNU0jpD3hXEE4c+xUrd2M+h0mx03nbPDdwx5An5
OwCw0O5B/lQgV90d63j3gaHWVyd3he7Bpxq27WLG/QZdOzUrcM3nbpxo2lQLAQTi
r1epb+RkIeFoxGW/rUowXOwdYSi18ahJm9t6IuK/g87iBL+LvxZfY5iIbzlozySY
QJlF7YKuZkgVQYW+qH9ka5TaVNS3g6mYw+wYybx4U/dj6Y+D/63067mCi4sv93K/
bI0YPxt8AvEZ2mbQ0VrC9rczyFevNwuGgp8rXNsjIdnCSruYEqvJqOyQuJoSlukW
VITml6aXOxZ4sT6peZZCoc94TSERaX+QQzpdW9QIHBneDENMr8YVFGGWVxYLeBgD
kUGuXDhooBzQFxiwDvUvIXxlo2D91Qd+F+jmPb05yLtVcuOngj447DowxGQCikhG
MJiXH7RA2TIdimP7rB1F0OZ7WzcUOD0h7HCh4hghk8/rgG+cYwD2FSVD0nenB3Ll
4/1aFEzbEMc+JA+QV8lXl36fJmBIe4iL6Er7Bz1gt+nExNs+4gdRBbwB8BpGwKs7
qWRtGUVa3iE/2uZSZ+KtXOgCqiHcEYh5u7+Nr0pr0cL3FZGWTwGLZ+8KpBx169gl
TIlWFfh7QEeA/JoqCwcgC1ED6q2ShZPgCOkLfoK7++t3yxXDgRESRb2SiqbsnycI
Zc3NdvUrCZtkBtZMwJvY0IvV2bNIDv082MKguhK4ZlObUbHmzVB0TI9Yfn0XuajJ
xU+uFsm+qG4XeaUfKm60P3EM2ImgOkpy4Z3pYWltqxswoR4Cllt54oWpzlbATYcl
3ygj7BdKqqKaCEu/P6ZSA2HYqCWlXVxKSY2BTtQm0bpQlkj0zg4y4ANDYUVN+zBY
6f8B0ls5AWnMh8h0JVWB/8q93FQ8p/R4aRTzMvneKnUUHD1O5uuG/u+UsA0FUtIQ
0sM1kHbPw7kQTRDuoKbNHohq4yl7yEqjI4ufZwG3P21Kw8WTFVXe6Nc5Cc4WW+8r
oNFcx73GBo4jSIWMJNxpirwInq0TSVRj/ItyXzLOQPwwndCDOOSesdIfOTYcK0SR
oLItIJdjgzDOn/xTWfQuR4tCpEpDR2ZhqsWsJTgwUBngeesm6B7n/jSQd93Ewacq
LlAhtW9RyB/S/MG2wc+vOquHvAhJ+yOEISuF/2wBr3FiySRII9Z99SmHKmpvJdkV
jDIzH4E4zLCu+aCeY5akrxZ4Dd5Jko51CG5kKQNWPBZOa3zZcGnQ1Uvx4c5no1BR
hfHsEDJV9N4ADxMkKK00leVW5oLFfz0laSK28VZKznaPTxIxMvAVFIx6bvnlavVK
tskWK6K7rDrrUS6JEk2ywGTUStSwG5c7lbA6q2maOLCVEodHmtynwnxpEcReM81j
aZyMsDPQ4HI+A9f767UtRtpWUNfnWGmcxtlXPythaq+BYCbid4Pgwenr5vXvmsIk
7Mj9CCmK9DBMq2OA7RdcF3omJLkwm5txWSusqviRfdgVkmZZfW0oU30EyFRuhYAP
ptwP7GNiAmBsSJ8HsBa3EnLA+BMUZTfuqpcC6g4TH7mb8Yp18U2yiPtGgoHtCy3P
GVddlVlvT2gczlyhHauvITC7gFfYM/iY9liN5Hw3dJgtKs8rV04S19zfkQF9T4oV
KRDTuQgNswc0vfEgmZVqAsVn//+TXkOucX9+fUmjHU2k4n7FbRj2sxsiq9n4+sCt
qwE5qqEjNNjOoJVM/qThisj6mUkjQeIGNHtiJM7LsF1Q8OJ6ylT1pIDu/DxY3R6B
PmvIlJVKGvCmg24LTUMEG8CSV73iQ3F3jmVdD1jZ0l8dXxPNzl0BjNjSWCS1Ge5y
LxkXnZKr9jeMr2K12fWmWQqBpLCDf3pjDKVT5sSbdCg2MGBZSGg+onV5Iro+VeAr
ZKngWfBjmnMbtWQjONogRGqXmHaJaEpsNOoSn488LRKms05i9Od6Q1lW8BhNFRLL
eb6imCw1Q3Qx89zHVBTbonqJJeZ38/SIBF4A0fhNdkKNuSs6nb8Ce9gEcFVs2ifD
2GRqpBdlxM+54OdfsjbG5N3K7Eb9+F6K7RqUWoMLGX6GOy41jgS2r/HahGmxdjiS
1oQVsPzFyKz+aPjJgvy/yBbaMjiXBPJeKwnLvTmH9LIT6o0uzJwd3ycpiegxb2ej
g6a9g4greI6sFDEgo63bTK/9lV2pdwXKjbvvheL+lQrbuLgv2ksgbYdAhEujwJW3
+i/5HuVOYSWGjF2SvMe4YyAWbzeA5kSkm1Ja0a4ZQQqmW4eS2VwcJbQX+DwHZ+bg
6qO8BkSxiVAmset7qhpXpjKqi4sZ1P6lWVnZCqbX2xbbe8NEVr4rSpcb5Npvq/ae
bSCdriJhGKWkLCs0mzAPe7/aCvau49SVCC29S4IC4f9s3+GmDftoj26F/AinivUw
uAiqQDnfi9+xjJNsmnuLLc+Uf6X2Xim6u8gpLgIN1C1d7ii+8xTTFQ7wUsQH2nfA
5HF5Ara3nWKn1ji5bkfMAL8E/FIkiMW1oPl2E+wHei5i9FvnniXfg95OKHXTrooS
FF4gjM9TMgGosbdYfkwqm+Ekbkdt9tyLPQCVEzQAyhbJGi3n2K0uywn9YlSknYLF
9XEHj3B1M/Qsbl4mu7P45uQ81U8o0QEZP09s1b/ZYu0+pDASKZIwCiPLPEyf26Iy
knID3EnJEnhD2FaUSdAcVTbpyw7izA0wX/FCbMC+ZIN8LldV2S5+8sWM0P+PNXD0
I2V/+dw6zmGtFkUbZ9UPfSh9CHU5XUIkpgxuvtnr41yFuW8iFXEkj7w371gJ349n
+B/5W2BR54BqaGr/B8Xq4c+cFGnYSUw+AyygVVdNQbvFHQ2nGoZmLlgGfpWyaL9I
+0GGGYgCB8SO6smeW2zjOKWpV4vjbggIU1/2HI7oxruXnw/CKBkok7uC3j4HpoiL
gkE3bVUR9fBG3VPOT22VEd3nuyiepb9kOqoW9wAOjUSKMVhpqulUJSKv7nKYSiEr
Mjtbbzbv3JMyZV+VbtF5ytuDU/THCLmxjbolEQ/vAtPPm2Zt3S9cPgo7TDv1nckM
uwV/bI3VKX2WEFaXQnuVrcCjoPykS1aoiai2owQrS9BD0fHdvSyosv115/286l9z
GQGZib8/SgBTQnF+kuuDQKcJGOJkEXP3cwxkiBVF2kHPRx2XrFKl5LFjw8cPUfSg
/3ikoGMfDLwmIth5psk8k0hnX/NsiKfa6I1gTD35kSgUauJWCALwrzCLYcIX2Mq3
iCQJNTIMXZSwN3sGsR1mUE1JmFOGjky+UzegiwwCk2UgEEsil/o89/7b7kgtQhMN
078/jPbw07K1RzpyZMSovP81Yth2ACVS+uc96MbHZmF/eaoDTYpsOumKp0EtS9uO
57HR8EalgMriJUcDeOF56cpx8zw0mJ5Rh/ME+0/yqZMap5mmRgjLQzVK4J+mGV6G
Zb7YoVwJQrWo7g5ben03s14FhWoao5bdK3x0smSTUSKb8Wm41xxYlidd1waNBYKj
T3tiynfvUd+pc/6DkSFG6vjasxDkulANb7tHyzmcsNYtxSuXid4NDH2+wNk6wn/I
nxC4FDF8YDpSTAPB6iLnxLZQsak3/PxD4iZ2mc4dYHZFBudcCXYYFxg4b7p6Qe7t
JN2PZY3FZrlwSClpws6341PrelAjQC82nZYtDyAF+VbPvV579Ro5VQb8jcMINduo
eSbwggSDznI5jwsgGwZGGvWyQAzUyZXaaLmme1oNtbBIkJVYQDxaUisJNmTS5gky
6MoJRzltFBr/eS3jSc2IgDLC62k41IG1t7yc3PHBfGut0PAEnECg/YQApjtKg6vs
Mo2Xdp0WKxMC1GzB78Oh6XLN3umOF3oevRzIBB1P/wiZClxd4chpHnXlbpmftAf3
CatYqw1gyc7y5KYD1H5Avra3Kte0dYUxwSZV7gBZ4I2qlYK+McZT2CzPSFKiRDNm
DN8058hSbNmRjx4EHSrxjBLG/PhVBMtsLIg+S7EptwCRflhj0xb+6CvzrW9wvVp3
DlIUWAjbkKG+uc2FWgvGWbVA623zin7GWHn6SRQVxOFYctwa3tUat3rC3G7v1GWC
QOWheSX74gD5DP6Ec153p+YOzt6QMmszdoDSDen5U9VwGbcir93a5hJnugIdHhBA
wMjaNDiQuv8+Bc1FIln7WxsluykjdHUbBcgGy2fiEt/0Xz66R4ueCqrj41OeVKw3
pGC6Y9iFprS4kyLrC6dZDqc+V2LCe1U4VGKTq6XOIKSpk+6DhWrbqpCqCoq93unA
PnsXqm2Cv2aBVFgv3d9DAks6erdkkxzezdl1CRpdtC9DPk+GQIcQRPPdW+ePnOCK
nUhCUuW7zbvsa2EMdCDl/0eeua4lKjnyP7Nj7EZgJt2LZnMt32QGiQxH9HkHtT9D
x7Z86Lc0mFPecfZWHm5LIUKrqMMNGq2ZIrH4CarXsFHlon67liP1/Un4y9/CD5sl
0SMxHv+l1TcWrxP5t081vXprJOAl2LGbBNjddSXG9775m0VYvo6tKobFk5FkruBr
Yb6uh6jc4BmuehmsmYyXk/Gsy6OjF9y2hu3TZzPlQbQe2VM5LkIvgeSoIMIzuu0Z
dk3eYDvKqvxCG35T+nQ1lzuc2igJSr3tPgIt/cYKpYssEkGVQO31astOyb9KJU7b
oW3HBC7OE6Jix0JATLIVKBd62akI7y67D1TGHl5OLFfAG7HdUnwSVQtSaeaflICM
MzjesnzPxFplct086pZ7j7zufehuPuq30ikxP5eZLhRY1dx/h+JfRPgf3kIzgRMv
5tG1NPhulcTkLOZZBHPPNANrkpYNT49QkUlrY1Oe/dzkAqTtt/ERfeHK/PkN/EXX
t3NhONtTZIMUkfyUU3o3iggf5YTezAaKX7FbCF8SuUiYeu9a/ahoewy44YEjoYro
xeTZ61+IP24oy6TmKgvdIBnBOvjOmLVOW2ANYDep0hsii8MWs0UqJY33XYHBVQNq
e4o5XW8rrQ5TUTlx5sexoTr1BqgdQxfFdsmB5QysZFs4YPSUR9/Nik7sEnnKCkHO
SGqCJZpjldgHFwxiCGay+D1ThbXZF5g5HnHsvVvhGJ2YiMuLvIIVJCUzmMMY5vd8
EocA6+HTjwcx5yyz8tjHCm2mKlV2o0/uQ1e8KLHgsybXGXAaDhEzU7DCC0ERSGnR
tLWjKnwB2ymH/IcrEp2NJrlcj72F6wOUE8zjxBd8M4Ij6apNlnIuPNCFrIC+Mc/2
Rn2NA9FUhq+ySuLwsUvWEriobF2xcnlOeT2/nZL/Dd+78UlScbZfs3ziOoAUXmjN
qmqB+y8GY1v3PJl4fU8+7IPSXFNQBBscBpGyJzgeUv2kc2q7X7+/ZyOBQPid6PKZ
+IjvBYlqHF9LlyEwpB9VDkXe4Pc/jpCrDQkoRU95sApeQJFWf0deiaQvTX9d3fGx
Ca0Wb68Nou61TLCa/cDneKEM5i/UOiXkUxSZFDkvZoWQx6P70BLnzqwzqXyziw4p
O9vtrYB4ws+92Dox+lEzbfDCv1Gp0hN1X1Z6LtdulXrv1ogcsQZxtx8/SmPz0HGw
SjEaZrAx+oBCY8dLmJS5+r2HLznOCCaAWLLWuoDuItTUs7VS79rgAkK7HSoHFBs/
oq/EKhw8sZojFA2pXBTOfdzpJOH2w0Nn2U6aC9UPWlvw90B6+VQ8FCgAnWen0pfc
VqWwkZs5BpJXPQK6e1OsY776sR3RIsp934MyN0Fkv/Y1qi6VQ7ha8d4gvryJFS6Z
PxdQ8PfQSPJicTfZaHUjlKr2LzyMCf/krd8vxwNp+oUO3Tjn5IZzLPxEt7MkUZPC
AMAlOI2C1YUsaYUsLJMc9mTacqgdTVNaQBMou/MCORHVcidEz0Y4k8S2LoT3+2kI
oZ4RYwdgEqFDFGpgSS62DISK5dEB7aDnJKgIYYB1ndwdp56H4nNX/Uiieo8cTl8x
b6F7UBiQW/eBl0odHMkogZ61Zms40jWvfRN9xBxkz9naREImk/aiVBMpvT8rger5
S0fchVy+niX3yr232ukqMtph6QIGBFukhVNK6CuxF9Uht3hNZm4AoXmP7KiVLN4y
93uGypaRg6z6VTdseYudEow91aQI6FQnK3Yw6VSlg9ftV/E8EGzrOFM0MhfWsfzQ
IwUuYtwYs1zfv2J4p92giFB1FRk8gd4gb+LkJbTxFVO0ApKUqitxCiyhlyw/w6Gw
bVi7XIeII+AyhbvukjbK9jTswZk1HTBziXBV/NBlgakDlyl1SujRoSeezZd6bi5i
zYuVT0AeQSJ2/Q3nm03jzDTeTsjqg99XbOOd0XqGyqrODXO4KV3pDBT5aI/vbFqE
2mY4VOgkavtZFOvUcgJmgHLhH03LSVtLQnLWvh2QwfxTtDH1gXxONFNLlp/3du3z
gexRUSYDzjOKF8+nvl40yPSLzcZ2EL43qXCcv+470mg03IzMR23FYQ6SjHYWhmRX
iugkpl3zsL5L0N6oDAEqa9zNGbYdsAEbVu3ylEC2IoJq2nsQEHXYRLDiKw6+KzVm
R4k6mBoK+yTvVXnObTIGDSBzOquJttCv4zhRI9UB9cTymkZh0XfdJFZgHykvJs1L
24trPT4hPW1PmZCEIlq/G+HOGBkIkBtY+r+OYPNZfBKs1WDlOxnvQ2uUUhARkxp9
QsXlKt/gP099WJQ+1hlfBL7JTLByiV9HiqwP2Kd21Aqnd/mNA2tiDLursnCGj0OH
/SpqFAlA0IsFchFTD9vUgdMame8UAnJQIVwYYVMuMW+T3kBSBNBEmCJs8vjNDDbO
/PS9uHhntTzd8cvb1WmC4J17i9bbwHkgVcCVZR9h+CcYw4KsDcf4PQ2kxZc3PK9a
pJGgg4YNBXLBRLPIxlARr6Vl/8yOgLOH8Kp6PWPJbmI8U8b4EfurzWsPAE/2E3wb
XcuMjueBjRpokdu8Nj2tmiNwsmEtHwtUhIP3K6LAnw1NcPnFhgrvZV4/SCybrFbt
GKF7bHalVoUjNgm0sYVscGfTU1ShmHS2JfpiKOO2tjAfh0/dFpiTzYqfZN1b2TKh
3NFTE/5w1zWWtqtBsdV9P7ub0rr7fSaBrQGrazYdA3JvCQgTM5SLcQ9qvFDqUl+l
P6JUirMFNlp89GuaMW11ebqfpnQuaP+T6XHCB5tmPmK+FCOS6XYUfwB6rNyP0prS
PpElmJPgN/EJjYjOa26logdguCb9AfXcEBTBDeYtdFm+penqsseF0PsZ8R6AaKsp
7OMUyarrlClAxENd+w+tqZyHgJ0NgEtrYwNbUPFWcD+X/uhddIhfKjgBM4875dbI
KmYb8UZ6ekSnKp2Fa79UCJyIpH7KFGWPD+fzB3FS7Gxn/VElkmKW+p17CWGIqqgQ
Q0lGoyWiTrmW8Z11eoZy0ab8Qnq9hswr0NNkYmA7LPR/+O/3p0qSxhD+XDlyR47I
yvd6ueKRVJ2PklFaH28o3BsZyrX5AtZhGsg2rHtGfJ85gNIKX4G+ryzW4uazidxk
qwvv3KEHbTFymEEQruiQe8N3SkzeUz0OhtGqhuFWH1VYuX+p8oH7Y5yv/W7pCoz3
pHNwhw91pEE2e5xYleYAmYHZih31mW1oH7zteNfm9mKvmeohrTRJI2z3CGwGS/ze
JPMw+gL0QOspQQJgit6E6qc6v6/qPkvlQtMVShr662JnR1VU1cdCLRwvo+1bv4WE
esu6CKOnosEX83QcjrGlZEjpEW1HwX7iCuHA6JMMqLAtBWimEzPS23gn3zzROJ6z
2+PhYvkOFD4XLUGCIYXOytiTkx1H3tmqbJoMG79XJ7nYmIkJp1D3HefBJb9n1D3Q
mPccoX93730rNG5/gE3mUGy78th5/wHfUUBYTRrfS9WbLlGT1+0ps53SnUqKneBg
UUq05U/W9RQyZWqq5iv/KqL/2QzCQ6T+6y5Oz+DaTVPrbyPaleEu8IgwVzbuAISm
/0/YjjQRmYbC2cPVUc7S21P4zbKl8mGmIyYpTy9B/W1Stp/BjDqvzMaD/r2la/M5
5AHo7aZIBX7OCXBzxZJIUAAuk+DsbiCexM1w2wlYV0k28ByHJhJp5hKQbQWRhG3/
48pZuoEbJ2fzoxULJ0/6gd335r06JiJsnub/A3/ISObvfc2/qjxZX/qBk1r4tn5p
ALFqRIGtCHkqRSnf2x7tICtFA0cGoXRctN01ZGkBf3+RKONwqo8pJSoA4E2T+QKS
nMO716oFoaE6Ci9H5wni3zfXU6dEFUYd6n8EvnI9PzGTpFzXGRJ13qA/PHzGKKTX
ZEe2j57Z/pKvpeYy0BS7srGsnqKuNLVo6pR6IWZ6M9MWL63QpE+YcKOkdKNty0ZD
E/QxliIBKez7ByPrKbhgVKFKXKnSNhE4YZWAk2t4/qorOnpHq5ZRnk5HbJHpRqSV
B18A9MFFAlqh7/yY4Eq46eVwMGnrHK9s8ZWvoFRZ7aYYe1VO0DuWXQVKYWKwKpJ3
ZP0j6DNi5B/9/VQo5MtV4MqdN7JR+LzqrL2vhjxeI/BHfyR7Gvnei3xkt5cbX655
iKOzP6w9PpqQTxX8Xr2XIz1zIzpgz7m+rXFTW5d9n6SUym1ZbLoqzWdnNXYZ2MsK
0BI2VK+ZamvVpCEpdrCzXac0ZGpBYL3T050b8tRgxPR2G3FzIExjpRi3QXHSwo3o
3R9RELrJ08zp2OuDeLz9uMT7+yfB+qsWWRMNco9nVy7GbutMeuR+SpwicIr3xeAb
oBsHUOl0a/bSQLnUa/CyluZ1ZofTHKirnt7RpA5ElAEbEyhGw7F+KP1Cvf0u0g3b
qY4ynL2+r/7QKONve9XidecTcfJct433w1ECQF/0K2N/U72QWhuCkeWeNkDGiPiS
mef9XTdamdGM3Xl78ceOVqcHQ3R6fmvZgn5NWE9DzwqzJD6D5RfptLU6KbdvwfPX
a/uOKjIZSusofoPHkgEP2a1nT5M/TRl0JAcbReNHywoaZ9/Cof5JB394YuWxdqKo
gwYgPR3mh/re+pA5wuFqGri65u21tJN3kzjZICStw3l299g28M3tr3dQfLdZABnb
UikNQcGJ/2wWpbBuGTqw3mYk47akIa/7yUlBzen6uhdYLHB80mFDxQKGLq9eIFgG
OPjdDpczi8YuyumBxX9Q+PzTHs0BvOnvJecQMhIuEPXrOio/PTipgItgVLyfROFY
FnH5a5z1hEjvMap7pus1mE4c72vnv+xLlRfcZoumiZzvttgSIYtxuLBnuI3sn033
tz82yLkCJ+HcHjMqub096OnqN4XB1SUW1eHPW4lCR3JSYAZkjpLHQMvsnLAaKJXw
7iXBYaNKjimspS5ILJ0EPTZJZZpTH0TMlucT+WU6EJIlTUA9/owR5m5p5Z4g1hNS
jGazl6HZbmCy8ohnkYHa2cUaFp1bEOkW7CWqa2SAAQOHk6JTtG5PTu9nuZOuCiZC
GEQ837OMoi9msr8W609fDUo7wD/DX9KE3VqM4Tw4GV02LfQb4ioKU3LX6x7f7liH
1wD9+N+k5+PVzAjaApGVZ2+dXT0mHnpZBjFs3QA1E7Qb8tJZJnnhpChv7BRLi58c
x6trJ+Qn98iJyJq6R5H9g3dsiOyw3UfKyDDl24ywMWnPdJVH7ai7JpCIl1j37xel
zhwRI7zzETbBtyiXYSqFKjB57JY6vi7ByndkQxE3EVQV401D6nylCrG56HzBPWJn
gEOQcqhHOyMAFANzcYpfzqgiWL6eoGgt68QN88VcrPcne7jd5mEfE8ORB9s04qJl
KfG13IW5Lb8nhwL3EhDNck1qZntyGmA5R9t9CvOs6h8GB9mqxNzHictNhVho2OX1
+5aUGBFcdM0jXPZx+In1qX0Oz2moKTa3Yldaec8ocseH5k8BDFX0WxN5tPG2kjse
YY0ALQl05/6G3RwcsZ5xOh9xmZzlj5Hdx103EY1Smp9xu1ocBVrOHAmsLrRjgGzC
VFz0H9jVNhp/AQUFiDqn2EpRvYfWQkf8pa683PycoCuqJ8TZQjbUJdGWzPaAQscY
+F2+7F1Kk3WVdsSiTnC/i8KnOc9uB0snrIn+v0YWaEeigQ0Jua/VBrXoiye5AMig
Z6S+jwfe8xcpaFlfCnH5UaPr3DUTf59FvCrcFkK1kP2qJBEV5XerxNEGgqjVIalb
dUdbhhiCcBZwBqKx09paVwBFtoCeCVAXrXg+QjYnH1W4RGtmbTgGLCXuVPmbTJ3e
j/ZHuVCBMXLyQW6UKmXv1Njcdrlz4JNqr2/MAuoYEZTV6ZmVie4cVUWuIw7j+We3
1OCvO5c40OgKbYtff6j+lE5aNynbgJpEi7y6bBP8whA53hCP2GwD0HEc7SHv9W2L
Qfx9pTY+CNIOk3CMUgXbvRfTsU1gA1DBlsVXwlATl/kToN7zJ+E583DhKY03njFU
Z5qMN+QTA+Jz64qJeKtiszge++WgCBUvzS7ufCq6N9T+VzTkY26EAJVuYalkIhXS
AJ8Jx92bW/i+Q96NC2/O6+SXFEwznM05W9s+x9o1ZVX7pOnle/WSNW6/m4d9QbTv
IJ6CDLZcsdd/qi42qcMO7k9TV12w8qm2LBEx7ddjw8J333oPHbOjYcLiTIErPdq/
X2/7Law4rO2o11rjzqw8lwv2YdiCfUvVAmW5LQtRzx06rcjCYa4VrDF8yk4LqRNP
Td+pxeTUV2xhv7AOF4HvaxXUg8TX6Fo+SnCwdIuD6VtUs4Q6rrZLBxNJLvDhX2IZ
+TdRx7rZ8LLPY0K9+nxw9UEFZXoa/JK17PSwoz9WU2O3Y/M1erVHmZBEmQ7patxF
UscylBKlqXmwQqeSEBB6J/gwmYQbJw13Fy9siYNUHtrLAcJCtpS26syFaM0RsrxX
8+VDrSwwZQKH4KwLpCE7X4gZXFMZsOYY0Iz0QKFSiNAIhASt+3OVfNbfiQ5J1rbj
xWtNEpV7gGDIxSb+7Sfy4GNaCKPz535RpejW4wWjFtoELQ/zkVdkHYmvugxEdamh
fjc817/kSYu3hQRcwVp665LswDVhknan2v3vWEeepSJAbdeKrNtXWeczalxVqvf2
LZfQOOZW7O8DhWtcmz+2nG/8j8h4zxx4X6uQxV4+rEbIMYrod7TbPw07iIZRAECa
VNjdqZmtXuZj36dQPJPSD4rrLoj+euRh18oLVlN8qXVasBEeBa26i04cttmrvJf8
hYY8rrRajIOO2CfPF+G5TdZY8uukTaJQIhTGgGyMFYBxoQbWMP1xqDxGwZAiNJv0
h9Q29+2vgazjyZ4Ey06+9BjLS2ETAkIqNCeDd3QiXBBzJjvgLYSDtLzVq99b9Q3h
S3yaXL2GiQ+uzL+6SNfHcyFuqNipRkd3MNGzmGWKyGZ8+hYuTyvQpchbAG1Y9bCW
osXi0oZEcDFqbDr5c1ElKr1ZwnltyGmNMk2K21MLp1bjq1K9+i+w1N9pq9ISAhp0
W6o8t3veKOYnu/gzrFnfIQa3YF53GNlB77wr6HQnXUmORrjGNDx1Ma0IWR1zmQJn
JVZmsKwEGxSAXSYTKrQ0Fmhm3yeBQzrbc64xWa4Meg8egUexzLyZGe9ziaHjwBrZ
TCS5Py1DYmnKcENTegZVKi7LEPk5RjDjt+kNTXDCs0lNhuuGMgePELyqZOeQQ2sl
wpg0nbA7bEM+QHgbQMH4TKGfgm9JldKOTevefHdjvJNoAFzJa3mTq0VUG2F+QYpe
t4z9WsmyBqNK41je2EBMjCb8UORga3Kixq7JXXDLwW1FR7jOFjP2yV0EKXbZdrau
r/gMq715tb4H0j47etTf+6kj3l+udKUhzCAfJ+WT5fHJaJIbaSU8bIPFTwMMnr/6
hrQaY1KN8lhLgnssyCOBgvpjGzrS5tgz1C78VFtWb19Lx/AJhDJvoV0557EvHg2k
kkQ4dSHKM5T1lvdxGwb735PIcWFmVaVwjyi997++3HNHUROW52rNE1l4GwKgG9Vl
RN5i2evhccS8HR5NGKSem7FpmQ2k2+9vPKMH6Hk0d4tzM2vnGYJWQGlxgt0Yzx2O
4g17PieycNwWEKBis4c6gEP8fwrIjEbZLtdPt9PKujF67+XdfghRRYJxcbol3O8d
fqRDv56dIf3HwK6vUS1gqbdBXfk4aLA1zRN6ZSOOEeXtWZcvpNHfmSDRcSixxkSd
eZ0Q5cqpU8xrRvBNSU2jcg1fRvmTI6t+cvxui6sxHb3p/7wjXYfGwFkGAwTRAAdZ
u4n/O+DZWmlU026lDpCrLPdnj6x5vouzJyBUffoQ3/Bqv4g1fIatEa7yqw8bC/9l
JIDlRsho2m+9GK2vtAWmCvCz7Qa4s0Cswt9otnmHOHf+H0HEsIq6rNnlhdHb9gTv
bn24mmDR/SfOaecCPAtI6i907ENEnZ4e80GPh9X7Krz2j9LzcYzYxaUdUGfx8u9u
apjJ9goWq1/gALNAVyt/wILcHX8gwccbzUaEy2PdKddvgdRx0FU5AuuMTsJfRCeK
kdRouvAOdU8vIDEYTstGr9uWQEBNBrKHAAKmKwtWxwbMOstqHFlQLt/0M517b3s8
MvPF+kKJl/TDqYa9I4b/u3JquflLrynF182VnX+7hcEiiHW/lTBIbCm0aNLM6kU2
Enc+yA8aoYxXlgFdJ/Ji23d6URpuKm/NqwlSTQc8v21szQPVaROewohxI7ZB1kLi
9KaNQXe40UzTp8Cu+q/2iIKgaYpp8xt7zFP5nAEYTPfkPB+92qrQucQF9WjaKfw6
5D3pHzqNaPXs2sKKMnP277IRbwUXh+ANPfeh37+S/IcacCBLnsrEpInmVbzZvlfM
JYO9VHH3+CYuvq0WLh5GOEZLhi9so3ulRjcADrc1H12FJnsLby1C8anFCLyQnLjL
QfmDe4qp34OPtc3WdzWj7iSKRMaTjMWkFHtv6fkdhSgcSFIdpGK4iVmgyGDWP3DV
OwflpYPUhQHhyNJF64Y8QOo+wn1JKwiXEJTEJ1+sN6Fg7KGuru2c4RLW+YH0I0Ut
PWsUYgkqCnGB9pVZu7Zztgv6ttwg/8cE1SEaAZjRX6Ns/+ft0gkFxNMbTuAqoiKX
atF5kZwdIKcb+QR82iNILvS2l+jrWqnR8JzqqJfSnRNX2PXmjtlxJYjOgqL2yDtK
XJAj6DF3kJVtPzpAiPO6iLKKVJbTB0RaRKuiuSl/BkB3oMws2UtlnvpoTzyMrgsg
CH2H6Vp2TwngEkU5gIW0WiN+qE7XfAtcMoQiSdGjFqXoMA7T8c4ZaB/HM1FBod+r
/hgfLvTVPjkAPwxBAxdG6/81kkERJhf8N+Lq54SUBfcP+wwkQBZVMAvzABPV+xqi
TlG6AKN7h3BcB8WqkhfzQ8q1jxzQbTF1DSsYywds1AXrIqqq3GZDQpCpONnesyFZ
hEIQBWOnePbLcwAECG6lWF8kVcUVKe2XMWwCJsZ2IYgUwcmcbuQo/pFRh4Pym1VK
K6hBhod56EfPcsV0i2/xHsqQZft/922d7lSh3T6qBTCmHHCa7rif3zUdl7Ig05KE
nVqm2cLHmTy2FiKcJWrhzv/kdkt5Ju7CWAZD4CruQQ6D8sns5D+4mURxKF3llOGc
WyS9VZErOu3k145NY7d2rQXb/AXN7UO3ub47CoeuWXqGVFeHuKu1Ut++W9RujHzu
/LMOS48j6dPGui5Pm6IJwRvWFuKa7v8yv320ScCekO1yDAfdRD1ZGM8oCMU5elsA
JJsbZEPCBjjKBOVW7Uc+P6pxanVV4iMyVMdLgFdFNx8rPNzSNniZDSJy2bb4MyUF
ckkwADKqUBhUYjJDkBnyjDhf5oqd0T41EEHUWr48opjwAqilpH174PkO9ivd8ZT+
aGdwWC50L0hEZcirGOsRVU6o4F4PxrNr3xajEWy917H7FKkrW8JpjRQg/4R8qFAb
bgmAtRy/ip742LC8RNIjDWugf0IDTouOHKbuq5fspu7uc2+rUTHax7UlfoO+keua
JWWBfhpgMvay2MplnEgPS4T1Mecq9CCAJVMwlNDxDXRPNAXs/NLbyhZlao94IROv
XeqSsLAeJqyChGYLkZmXDcBBFD101kzywd3oE1aiO6mT+dRX2fefhTVcfxg82Gy1
suRfklIwTjQrk8V9YZUgkBOf7PCBJuU5WBdCM9/Yf0/ifDDM/1sNErSsyymXKSWj
hFEaXe6qPavRbBI3sWB1MGfK05S1nORla7WNY+FaKL89Ny5RpRI1AnPxdjOi8KWP
Ak6xzHIThBI8S7Y45W2jKxdukljnjOyGvsq4fiEq65scSMftWTYGXScgP0Ual9aq
SVE7oQmwRcWsF6dD1RwO2sARbFTBDkIwt9Y1/g6W/ELdsJF6PTP2utTDj6V7IMHj
b2ZVj0kfz7bhs4FPqMqQSLSvtAGLDOgyhHAj7m9OXiEMDZEGIRQKKUZaUnhGiyGY
5HfFxUmnDs1I6Qs8DStfQEmvkkey9BZo9EsMcmfdwlo7iRYP+BprgQWVWbgyx5LJ
pJmtg6YwIYACXQ/athOnsJfq6lPnjq8qkMWLb2MVnDhefumhYWPa/ztqFRO8n4Lr
nfn1L+2WuGwY1H6NGSCme39Dx94rXkhB0URJEAdG0zG4TxWTOnuv0NYwnspV72zy
q38glalN1KiPwruhA/hlCYWMYKAwBJzyH8kF15sUkQiMKwfSo0v+9r2XOJ/0kRxY
jt64aYJAGxrL7jS/tVyhgZCPT9bSo8QluX4BLGvq3yUc7HFKAON7b1G3jfXKkHJj
HB5ZBKKm/ptE008Asn6zRpvZbOQ6KzQBu1lgaxtG+rH3d2wtdruPw1OgpVHgcTj2
JqtX05taQZkb1RgSm/rpcfM9GdE9GzeP1gGLiLuTanDvC2ADwwDHEF3su8jCnxj7
6r4RbDzHNdWi6RbxThPmHLGLLkxlmrsqHtSABJt7ec2IQ5MT6kZq8950Zw4PTo6C
g/W3MlYEy4qrraHwn8FYt5fCDZjnl7BhcII+3XQCg9qUmqUCm24KSIdcdg88mSVm
vja5NEYAEMe8RdQnAaUfOsDq4drSqNdbS04DLzxg2uE7uxqBSJM5dXOiwA1xaiEr
4PqiHcFltrYt13U0IaZc+uMtw9sNIQqoxbOFEXG3P9ADGd/jiaLgNEqS9GbE/74P
Ttfd5vilBjWCsI0YqM+v6+VxQmNzq4tDl3vz7imdMO81R3YKEuNRoQAZKnaVDwjW
RaQInaCF5t/MZTfoGd8LdTCc9ghUggp8q+uX5lV7CYbpOaTL0EYvjKa6GxRz6w+P
vbLhvAsQ8So3mYSpuA5h1b3SxwcW/Y3aZcQdlQZpvbuo8YGyzqVlPT8luFxDF1Hm
5kpPoaq2HuazEI94xPS+LR+Fp1kwLP8ZHugg5J6iCdTsII4uWkyjbuxZINjUS0c0
ZHGC7rgT3k1p1kzNB4QWTsYU/yyuYyNod8W40IPWNFoN91VV74TiNvK2cyn1aeUa
zSWmTm4Ao2aBabNkXa/YImxKGsYvYoPsst75feOMzowfE8IEXQlGSRinx6YFZ2jA
YteLPXlKSHxk9Sb30jOIDgpyNvzTCZZs5UJkrqO1pVSxcVXtec2hR06yR1EBg0BI
/Wheef8asil6fxhGEk4T9iV/wnfd+FCn4Zzzupwnnnhkb9gJGUojZhEzgBQpzzUD
b/w4BLeyRk7tkZg/UiKMEi9eNEdV9nwcL6x1JbHVbUXgLp+tvsVIBwAYK68YG5qG
we4G48tqX5xgLY10f6BliHa7/nVaxJOfYz2gyVhDYRDFw34O09LfgxNX42T6Z96X
W2h7oG1Yx+/BJtwn7A+sXiz4v4M6rwaqRoSarO1JfZNVcaymJE/c5Y2oFR8LV+/a
T9L7IYKli2oQMrmb3+z01GhSfm32Jcy/PTo/JxX9uJH6vw2tlgxBz5Od1mXF300e
5euYa659sCdtvuicbFzmDkeJdigXhJ+GczJjZaXgZ6pyKjuR+LxpzMPet3+nym7w
rmFR+Q5yXcgGMQrCGzI58VeH9yjsWbS3zWZ2gwEvpUKLxdNd3BXd93dLFEz6H1/Y
tzwTaOBDfQNa4qdDM6bgThjDjIHg/1GbeZmHh1KdfTUDueyDuV6ilTst8KBMhAv6
bXAQOOBUvY/klt70rgYVgUrcUpQrum5B9KIWAk70WA4Psuf9UYpimTmx0qgoI3q0
yqBkkzHz6a+xEV/bEwI5EYXWpKTujLKAMM02AwjFltm4NZnbJOj+764nAn/nHw/Q
+IotbZVAb+N2qCuHnI18TkJKop1OcPkjmN5Q1lUQxCOOQKqIX2xoqU2Iw1vm24S1
yorEmveVgA5YscLPBOI8nBsfeGXshmXFVr+WepOsyiXLEMu0rRQPQ2P1+eVFVLFQ
mQtr7HlbcPCEVTUgDCP9vlCMGq00oojFnFCDloxu9RxSiHokPMAEHmlfdAT2nCjv
3Ok69U6dzCkTAge4OcI3PCPr9Jj2tNuVX5bgwO0lsxzFmxUde56uhQOzYJwR4sOb
DetebHsT+ZoOXM3rsQI3FNISlhBcqT9xKOEI+a9wWazu2w1/l4wJJRL4l1+nIO1T
ijv4TBP0FOfUUaV+NSKrWGBgpGByhciE1dbUCL8zOSB1S97kvoEpSA6aJnEgkk6O
VrXaEJfUVQTbuoD9ioeKqKjIR4VzZj5Lsw7Hyu/nG9JxcNmX++KtOFdpB9zLcok6
DHOszZL0+jYjWO5AzGN6ysViDzrmUb9+aOOc+KpY0n+Zo/iGvx6r5xK1RbVBzis4
6gf7U5lVOD7TwTG6YaWuCdo1ckgZEJfTZchg1APHzkUcuhEhZQpQ7JYqeYAQsvl9
RmSX2bHJ+pwkRe2hz6UpZxjjIe07Tu3aCtYr9s6jBREnxQsBS6DULDF2FgZIvoh2
o9t2Hkm1asxNQ6DrZXmGLzt7Gmt6FhI4vovESHauytpN3W6019CsIJAfvUCwDxHy
XOpZfk7uQLGHsyI2zdnswjUIb2qcUocBvKJe2tD5mP77mmP4EB6N+pLCLX6XIWjy
9zXQiCGJoJJrfeUgc5DsjsU0//Xo1w2gd/i8KyM/0WGIcQG15wpCyB+eeqCt93xM
uES4mOGrmVCEjH9mbCg6haRs27Bt2H1+ShTW3tzPTDNoPvdrPkwQFWviC2cgr884
NPpNB1sLW5L4qglfFDgP53LkaT5a3pRRFSWWeNAYfstxVeXlTvCYkTkeq8CGHZIJ
E6ifoqGl9iNsUpR2O63jXtgW4ijXM5S7J74Dxhw+YSyoRW6gDcSKidhvIpBAiauJ
pzlijKu4djHzvAGWI82S9srPu1f6gPO7CNP4AQQ0PSxpc0ucm8PdtAlocdj80Rg4
SKp0vCq4VL4byNMUHx5Uq8hzyTDI19f9nm6fbB0iJH1JqQLO/Tntr9OzJuA6DWKi
2tbQU65H58nNQkDRSLcVxO+cj5Vbfb462IEBlAEpZQdlcIZWuEzqsp4xIRFc7cHC
2DdzN+3XjjusAka6+dCijYXZv3xSJN4bdc9VVtb3qz1EYPMXn6Ehru5jJY6Vs/oS
Bh9x/ORp/iVl5r0Db3dprCGOmtlnUcx8JfqFPZVrm82stFipKgnDD57EAPzhcMsr
de8M7TYyo4cQJu+H7qyW+3JlN1nVedcI2D/GX4bjveo5UJGYrICkGqL+t1EWvK9m
UdzDI/5GShq+zWfbf17ovjaQ2+/1h6KFHuyMaYEmeU9BAX6U6bJTOhX22VmQ+TTv
ykc683X0Iw1GSB6S2ob4FG2A1X/YceI2i+5t4Zs21e1r0U1BDYTooLjqOuqFbj98
KVNe6AHhN78jp7je4x1pVuPbcJ31zTF39roHsNfbQBYqQHwjZcLJRW37//vAcXW/
6H/NhzAdNSfqQHZaBgZRXp24yDbuwdJxdRcZqLGBi9LNqU+Qlx64nQNoh1Whws8l
JFvSTDBBf10149ZTY9NjlbTGW1F/I1tFU0BBRkU9lEOXRxdF78cuyJuRposWd4/4
AecTo07EQ5qBZRapgs2YUnmhCOEB+1DtV6gsgbH0LWnNLdz/NeV/7fJyykLe4uK+
mhnVcPo3DIIe9EgKpZEnrQl9nvsaKyfVKxfq1/Ke0sa9SWq8WA+5Sx4fKbsedxwp
TWH/uJUNElKEV98jyeGewb9pzokyqTfLv6d68YazMwIoGBUPgFf4qchocGQVa+OO
CmxSx/kF6Jl+6Z4Rm+fsHJ+acX1TRj7/XPG2/iSQs8jMyYRqwL+Sh4z+RWYxOlQO
+4KaOUFUrnpVO8t6KAq8HtQMPOTwJ4FU/MJgM4KNXQqWLVoR7lXYNsGTZPY/MRU0
2nGcWL0O7BvyWgBhjtpmfW5JHnSvf53BtPOR94VEP1RE7W+S73eG8Zpfa1ykU0hD
W2HK5SUAJm0RD/298V94Lg3WifjiTGbz1UFpSa1gKU8igLvv1eFUvgbYtoNFSybj
B2VQycYVSD8hER8mj8MbyLeDTskMZh2odAb/b2lAjK+QQcEOIfrTqfa5E9ODAKtn
n1cjAaFQq89Pm1xKBD3mv3FNdjKChYb/EICEol700qZ3NKgYZMLJa92JqSNmo7xn
PSq16/05wIWxjJ3RotwWzsPl2pbcStCIoj8u+W4JtyUNZtIfU/cZ3bdkWY64TgIe
nw+eKLZLaxQS1eYSF/LTI2/p87o3M+x8MqlZ8ZBQBVxPlOtvXaOkO2BRbBTA2hP6
8YdSMdy+cTKls5VW+tiF5qAAud+Z4jPTq6NmR+qNLFPV9Cugrknd08yMt1+RigpV
RU8o1nKdItz1YLrzRhtqUTdotEF9Ubgj+N09ESAdEQAVRb6hwfqTkLRS3owA0am0
6/rQvOJld8pPixmey06uxiTwMbMUvkZTS0cBi7FQcjnppDuohpELQ0V+gP8MVTCV
TKEqVX6YDwGNwHlkF/PYBXcpv21IxqA6+WOyZq/P37wanJ+674+5GHgLkquxFWvx
ZoXISyTL3NtfyH9yHRrKekLQKd+Wo+yhu59/QnowBINF7442KNcvC5CrzoDZ4ndD
CRHoicGvOBMHZIpQCwTim3hni5HqNk8rnXXNHE85r1CqgTK0COVhIcMVEkpF6IFZ
uanYwo8qcim7HXu9FhViM8lxaRRfam3O+0dpAIMpiPm00uG7bFAgbLchXh0qIPza
tDmfJpjLWW3G6c4274sSKNoPDwiyXqbF9wVSWjZQ8ANkub7p25kqMvYbW+ddL/n2
vFbmPs0cOex9vsrxBfFf+U0GCPcro3EO5ELOhYewIi6KIZavTiMjYv5yJLMb4OjC
Eols2azq25AUlqHYh8RNw0Kd31d3qnKqkaMFRe1YQwH7YZq48ABUinW0VEKSFqPj
QIpJ6ttxTdcp82K/p8ftcdFYgfNfIXXfEDB6NdPFhRpNSWnlSudJqGpQJNkAwWJj
CPXVq40sDqcj7VzoGoWEaWVsqaBesk6Xmlr+mcOskWjL7t6rVsEqjhQOH57lqRiH
yPHB4TsAuAZp77b7SgQdCu0knfPcSF8CA72TzUMhJRmX4B1QTk644ItKWNenOdTh
vBkX3V/Pn+y1rEHPayb4nlI9YEJmQclIiiDdXbSwNYCl68B+UZnSU3cMQb9xMVCe
R8sonv24RzolKfr3Ws8w0KfNi4YD3QWQALjPXqfcjnaF8iX9zWeW4jg9xNRJJk6v
cpP2Bo9dD2T68/i4b3v4x5be9BOwLPFB2fB7OfmmOjogZYMOA0VvNiuj2EUj2T6l
Z7tB7+lz8ygdxfX4/5wrQKW7lMQZiXiGqE/JyXooB2So5VklHwv5NryE3XtlYOWe
NxNW5uVIxCv5zUNq8OiAXQS/+KBY8T21+bkYSf3K8Ex7Qdorw0TKef5YvZdjIAtC
IxWOyIQJilMgrac4AHiafyR+/y7v8O+9GD5DHdpljtbjWBvqCs4EngI/szAWj4xQ
Hb3IUvzl/igrdBspFWKSqRfIKTdjZP6gP/9SY5dtxDI9MmdWrYfNbooAfBJ5cq0E
usdWRw7nMqV5UV6xigZTLhMhmWMJYJtD1SFQY0jgb78ATy+H9GAaACD9ylCMiEWd
L9C9YxeIxUHwl+rVqkFK+i/j8Hp6wFu0l+909m2W/iLvxNH+GwiiUjui0o86fN0c
/kxlCSFV/3l6+U3nwouW303UxM3CedROueOV0LbeolAKTZNuM2WPc67St9sgOMHX
psYbsWhis31u5ymtObPkNiDOIkG0xlEbDLCVkTLupyQG87jdbk09CYRYobVYE1D6
irP8rmz8eLYd6Ss3woIGkC/L+z95BSPiMJN2ubRYyTnjwWPI+VlbE24tZSWImp1c
DZBWhOnOn67WWMcClW6JZ1s1EoZ37PMnpCeJqr6h4/hNJp1hdUls04mjUIPhLmNe
55stvLha6L348Nh4qTr77kPiu+kwV9D2LtdjVa2omTON60/6bpA3Hez5sIPnnldF
dZiAlSD5kmIXtG2vnUK0x7AQJqFtvaTGocjXsJOk/G7FxYFrUn3yQn1IR7MJrhKf
UZo0sUITB3j4IJdHF85l58fAAEUpuWjV8fSXAeHtiIM0xZXWUj8E2oju8w1yaffs
v1fx7Ann8uVSU+4mvTguCrCvkoSV2TuTxBG3HyivdzcgRMzlzTJOXW+un0JJAQ9Z
A534/V98ubYdx8B/vcPEopNLz/8rJdzz3Tj5+4meu5nQFNBke5Xha2EdfVJyX1WU
0dVFp3091K9FrPcnsj6pbbUC45EV7yLWhjvAXeZlLZyQIKOYnuKdtPCnkSKSEyYJ
dT23XVjE8xlJ+MTENLVsIuGfcna12QOvPFcO5z/8grr95KF+RCfvfQFUQMao7F8n
lF0UhFdGpA7MHMD+G9VDgPaDb8doUbWZsl0TQhRpU/DtUeyv/h8OMvsHJFff/FFn
x/DUFqkPVf81QRIzTwtSIICFzERUtwgh0JmfUGHSHxRcQIPHCv7wA2psr7OVgLO4
LPwX4SXXc3ShQUf2ZAV/4jkkRgOuOkyD+DfEg5fXF9ixESJcKEV9XudBxycCgM/D
E8Oun7pELVyoEhMEhRXlxso98bJkGkWVO2JLJpeFg6ZXiFx3tMNzJOlL8HH/zK2f
7h6rteaPpoEZt2B4EXJCWoPMHxtCTqfBSnTbZe5lWw0gvhtQ5prr2Yq2cfdC+7F2
pghlg6yAjenVSvhF+2EHLMW1ngg3gvYP2wVc0RXoHFhKm6CrE/aMmEntkiJVoCBQ
PCZ/etvJrtClTk9bI3jEV5ScKfLp2ECPsdHdncytoXQHlz2s4Qh08w1i91HNmH+V
jZd/X63NTlVsRnDRAVwO9kDPDdPi2luuPnnWzF8AzlIgfbyhBvQDeJ4kdSYFDXNt
6/thvFszHv/Xm0kDg9bEee/xFh8UEZAP2igt+JXhIShxx+q0wCsPvJzOmP+O+AHq
m55UV5HsQJARpCQNjENCaRRGK8rbg+kme/w6cHYWoSpeBhOPN+cScqZE2uX8TsOi
Wjo6QfqcehNO7GbyfJzfxqTnYeJ7KJ9LH6YD49VWaWjlj7VPlpiY5I17xgkI0pEi
gbCyoii1uLmlywMtFIa5elr6hqifE/re1MvKzHURfq/p2nNQMn/qL/PTr4oroS3H
GumYvwJPtqz5lSWwO345JUcxrtsCF5bz4kx8AfujuVW21xDs5U4TPPEbH7t8ioA8
UfIxN5ZNBXzEjENJekVu5xpeAUSHtibLvfNfaI4GbvyG+5OVzqxFJZRTRaqJZXYI
YetMV/1bb+WQpyp5bQYFb9RjDI6g5dhQpYoCjAMwX1yfioLTvh0l3wta/C6N3tU+
BT2T1a9QKMKmmG51lIl60dm4+ikLpU2HeNPB39mCOms3wNzIkE1I2RlbnKIutVbL
ABeRDT9ppWdc59G8BsYCP8+uALrGHEbbUUmWckM7byjo/bHwRi5fO5hhJLwKJng1
yshsnKAkfqLiOaRL4ihqkbj2xoXETI3hRlx/x8VnieKAMWyy8EdNQGW4aNTMxAGK
PcagFqnT8U+LLWU2DKulMpElCsDqLl3fkIwu+h52P98vBiheMI/WZqBnzez3G0JM
vq+gM2cwVlqm6Rw+hRYv3RbjYF4zRhxTIwv3NMxCtQmI/xRbVJDR+d30YSIJw3Z3
bATsJQJn62Iw48CAVvE3Noko0eEWDx5OSUdAeMLamzBcOSFeLjQT6BTROCDLZRvM
QnA134qRakWL6gP9bsl3aDRuL7mHo6Eu77xperDcuXuThh4ALhZBJWZe+4eSSA6g
mDvC90GDnc5s/hpQcblfAc2BLXtehFD8/4peUHbKr6vJHI/MGb3675ib1MbGUeUW
MzUkEzsRn8dsq0CTQvzeUb/N/YSZl0QSgQPXtdQGtRalZ2EMwgxz/Ntjfv2E1zi2
HW3egR6HCI78jEo8cljY6bS2F4q3Js0bjIJqzEQDgKDHJvSZJxqntU9SFkcRTEyk
g31ATtp2KU552Hwou6tlNgyoaHfAoMgH44MGB07SJtPRDFUIgGh+Zd9UoP6SnP9R
C4laJ2hunfiQ7abPHg8e/ETO0gCkk/OH7Ngy7NNBhahBSFeQ2Dj39TngEMuyrYC7
rY3W9WvUkwzXayF10KzRMYaXZH+Q4dJZ1qHO9fphya5b4D/1aDHSn+zaC42wHHC0
iKYjSM9ZEtcgq0eGBbJbHOK72HHxlGYw14ey4jv14wjQ3jTc5/lOi7bZRAn9wQko
dqf22iIsm9FaDCo3rtYYUeea/S7HpPHu2yCTsXl1J2xCIwfFlw3XFbzhMh839o6u
j91yNF6T1akzwD70c/czRGp6tvpBUb4+3WCWY+bTUP9r/BTc27/AWqoriHDHvX0b
CyoakWvFQ6sRUFZNlw0QHyPPAbGOBAGZCr9O32vHU5pfdvhkLk6oOJOOPJv/6ITU
kUnQuZfhN4T6VorUm/uYY31fgRITdjeSzy+ZGu033gtRV972YG7B9HvRpEA3MZ7L
UI+CcQlIMo6w5NItxPldHKspeg9hyjMnXBEVQ8TGCqOduRVvnZpLOrCzSSP25Os2
M1B9T+/kzv55Z3/t2676R6OMoceahDs3K9RJGpP+OOTE6SUVKy6sOXCIwKoOYyJ3
d3AM9miLBxUwesVpv4y98GA8socmEH2q8Jd8Mql+UVGYd8lA+60f+3c2BPU6u57C
TV5PeNRpzlVOH/ZYsREDlk8/t+NOuM28QJCO2Vda1DdU6wt84wsN6TfLfutYxEvo
tTfjUGwHOqN3FumvbuzJe60ODjX9ICkUou4ZHE2WOh3f3LUZupfvpC+CmZIGkC/k
OJeGA0udKc1ackvCa1kp6Iv75L2HWYnu2oYRvAVU+nacWXAy8RR07pS+HAlgasxC
UpjiwAuHBQ/p88GpHVZ7MxeiehmrvomAo5vytgJ1bjmAB2fC2HOkBTGlb6VlSsEF
sLIJ3W2PFHKyML3HG2sV95Lq7FG22/grHYN8aX1kv9I6LvqciLoPs3UELFY8B+8N
dc58iwUDUNAGnv9O2Ho9wDV9FlMDkzYPevgvMSd0W6IaCls6Zd0SUlzLSxWy5Rn3
OsZ18MwfMLdxPpEAL8jOX9DpHhPsPooPi/zrFdpYg28rHuWuDD2DiclDKB72Io+l
mvepcg6yX5Vnfqv3X9AENHWOiy5tDAXXpBzhzZ/cZxzFfPK0QtAKFGD/f5Y5v0PU
5mM0OTuYZQ8YOMvCZQhiNk+WmyRiYoNa+dn6LxeXEHvmfXCACm6N8BSN5CXf6OWN
YhAvLsWqmiu3+5kr3ZwosdIAa+w4ZFmzKNlDvcAZObQ38JV3VOdC8P5o5iWX8SgF
FOv8fN+Fz6XpTa2SnLTOx21KYxHUXhaKXABovShIKOii1f3jh07mjB398lyfF9yl
GtocWnaQHUZwZyhrg1AhoWd7StXVnUeMd7jwM11ZpH4M5yfj4/xv5psi7lZ5zSml
rHuebbLXmDxRZb39986Jb9+bC6Mb4ZxD9tD48db90eKw/w/oQ5n0plHSDaoj8CCB
v1sEkslLaFp7xW+Q9hjYFcPsWlsRKmJaNqfCUsU9XjIiQcLNv95FSoks/r1xE5hy
huvU3j29wkX5J7uk8yxjfJuQzRdvAek12obQ42qQM8NuNbjEntOtaiIRCl45RRFe
wAQPqoRCZwfO9sLuPwFlP8/Cwcbcl/+qjWM/Mi0glQZMvdw3I0ZPHTtBXleVMdWl
JPmDxEE33dvtaLi6ftLipFuyyhRfo51stJz200Q9lnfj2Veghbb+hrabQ4lfsvTv
5bNsRHR0c1cboJYHrdlCP27WYBOkK4+LlKO4ImDRHURxE7OiEceHM9BUrWOx3VPX
GAdro1ZaXRxs/QjsjgfPFyFEHcXDRQfThKBvK9Ix9BU+i56wmzU1Alof/NrNlCa8
SefX2/BpZG+lKkJu+k0YhJbMFNmD9KhBIUv2/AHbfQlaVIodkl6D6gWtKIdSSql3
srbcN2zPWVOEwSGaiyS9bAp0X6bsGG7Q9AymobYtlYwHcCpiRtlBkc06rb6/Ap29
rVUlCJN19pUawhZTURLCe4rz2eC97aU+JHmoZ+oJeqPDYFl0iy23F9LTv1lzfLc/
DzyOYiELmZ/Uc6j1wrXVhmTJlUhlmNRh42A9ufEAhGFYUcU/JV/Q/c5gxiuZkzBr
PfF0pWkh6MBUwsBZEzB8a7c6Mh3Y5FlwTFpeAb4QRwkFk63SPVV0yQG6/FnHglR7
jTX6UdEZ3MqXqksXpC4+q6Gt8TTEjyGQIsevwMcUWU5klXg2+OsHNxaqa4D5lYvM
KLf4Qz/zaDpHhF3LCg3tB1uDs79lVn9NzKwQCM0UEmIItPNVxpnx+cG0n7Zsqxvs
uLQZuMyXTDdybxOW6r+7h0XOnuZLif3zWB50ROeFWSpeCADsX1l4rWJw/ore/bhu
+ErpXX1Si8xJ6oslJLUUPQA0n8u6KN+b/W3u3MiBO9Bc2jcYsAvb6zRICoynnu9Y
LBopGVZC3aRo8WsCJhFkJPVgbc+n7gwgeh0nYbF3AE7xPxdPhjvKYQhBjLnBIrLB
4SaH8HUu2ts8dDh6p+5JUx65spqCXN2EFfWsgb0EN2TyrbT6awmP5JLKjxsrMlIo
4MovZO6O7R1MHrogwVcKPVxf1sP143nJCgNfiBtdQed6rw8IYTovZkkLud04tgXR
hEdAoqIPEhA1ybYi0OdedvxdaKInsHXe76e2yXybgwfBayPKyhFSS8QQSd+BmYl7
affAg9VaO81g7Uto3R+KrYlospDrdgygqRtxLwWbtHyBv5AYqR+tPITA+/d881RP
wlCbxH5wONwgeqvia0urMiRASLSKunzUfgvKY5RkCdJ0XhxhNqPMRUyz58bCDndY
a+kNWy/D0V/nppDrbXXRKR/QCKtRRoOB/B7XGqN5oOctKiR79D/vb8hz9hT91N0n
s+8K+nwe1hSyPLGlJIgHldpUPgys/TVPONMO1vWr8Rzf4WrKCBQZiVXFqW8Z2hId
xvmGiRA3uTN9qRmn+z3FCCmtWedm/oaqWNkEthEp7DZQyP3sI7DvCatNcKwyVhqj
Kg0Yk6u6goo+wWBOb/U3X1o5Y3DajGrSyoovwHQLx+cz3BPuZZ2MHCeKYBPpno1r
TOCxjXDGokY5hHpYEvBKSEYyrs+M26lhqiD/NWy2O7gETt4dpmouUCM43CjFI23l
KuMhUahsOnONimlPw+rRfHsh/tRuU9xj3hCo1PFWtPcTLhjlLRyUHgbTZZCWuugr
I9zdBpELdmK+mY7kMHpxncPfBCs6jLm1JKEpCtgGKKHV9ANE//siApUJRW2WosvY
QvkJbzxYwNIc9+6ll420Moz3JhYdAcv68jEQ4nxVKBRruEtvFkiRD4UGLH2oTltU
VNNxpYaTHVxVcuOQ1FYi+BOsAlM4y8BuR5rX3pI96g0aqSDgaqQsGQEewZqsphWg
ZkJvfGOBVcU3CFUz6Lu/kplxkT6s5KsUvbDJVbvzioEDiCCU2g6iZT4R5g+GnqGR
P42HtZ91C8slXmbAguChRrqS+9aZFkskdQQY5xZ+4WZ2rH3c4rq763XALmeeRtxA
EhN8Gi/kA/G/jRrFFbQ8bDGlMBOec0W92kqRDcvsU9DjW0DJtQ5yX/4QRvR0gIzZ
tlGn5sIUF5lS2R24aXaYkaFrv6wAJ5bt1GiNpQ+f3zHeO4DjyiaO9AG8Ox1pehrE
7xxM4/Sq09NesouoWJpqVoXdHFzK5zKLzNCZWg3Dm1+S6PTThj6z9JcCsq1I+me8
SIIpucw/QRmsM7g1eom7M/wmlRcFca7a8fI59FGL4olXVZTGakMhMa8wEMaPrjIJ
cmN8JTmlTa2sA31yFBbAvYSDG90TnehrRNMtYs9/c6q1IPARv0r3bmuZy7be27Rk
dSvshS9fTMn1jElS5mSYe4cbHrdH2eIX/r8RGvQYapdXk86rSz8dShxtXOCBwrHb
w00kl1N94FzHJ+aJMgSEdSBOghgL7PrlZ4WkXCyxRPwmSEBQOARIqBE7AjgWQYtS
zpdN+TD7ciCvGZm6ZMzpU/sBhFXMmxLMbi6KMboi29GhqCo/NO8c5HNHxr7dTdDx
Qu9pjt30bAyWGVDfWHfupHPaeeAcaLg5NA2gCyfkDi24Y3W8di4H1q1slj1TlPn8
ZozDloMTKdDXBlqAJs429TQnSquqSURMLLqXGIst4dKFSI08oqLnm/mJyiPb8fx5
pdgLRJSMAnd/7vcpqDfV2ZBZRJJLG6NbxVaqGD0DH1uWNJ9sLF43pZ9FgccXGubB
YBlhvEpMdYG2O0AY2K+tLt1S1uFgJG9PdGQLL7xDmvOY4KgAra7eYYPYPCboBQsm
isrdKpv73C/2gmUYqZcoBK46SZPgyRnBm1UDgmwiHxO8+2D4iLs9eibJnwwoZSeK
o7A72KJR6LhD63UCXZkZWacodh2TLHDm6WKIslWHe4t0llq2UJy6xc2VcM1n3SMx
JXJXZ4xIpuZYqXGoM8QRJ9xDUKIK8DTy0rBcMoPZOBD+BDTaOT8y/Y4KH2jicDQG
HU+sHKOe0p9ua2BGzNLFEsiQ9n0lUxqm6/XP65ZK6TqtlxzpsGmvQ1vvvoe4lRSW
QHwmTXxm9wIdIWulrYdrPPNyJQFJBzDc7CBl5f8JKqdzTTfMZCRT11T09uu8u/+l
j7cpK5/6EXQH0v1P5cXmX4yTOvK1QyHj9HctPiab4M9QWNihlg1Y5SoAsnsOwyw7
gFxr7A7agRGmvPt0OAgfd8Ea3HLub4vEvbc5F/YuezSY/sVL4Id+DMkMIgOL5PrN
3CJyUKbJFTp6Umu8OFPi4GJaCsrgi2S2/076AXDH2ZKmPt0KIoG3Inr9b1uvgsho
Wg46O1M5Rjda51WQvrao1lZDVrwONYjovr/DiYTccVSi1jr7yWMf0uCYTMvyUDEs
X1AdUifW6o8JECT7+EsRgblTsrS31GeTCM8d4DVeRuhbEcl+JI0easPyQdvvZjmp
lT+AxU8a5JqjnuGJYWYyCeYldscop1051LnCmYIVAxRzeJviKE71BoRSaym3li3h
rYUXZacz17BpI/XeIAjYGBwduOqlKgkf8q9Sz8nxA8QmXLmzk9oVwEZKwnFd04JG
zjXjXyi2ESItk/CDE9ciTPMFF3HKmJu1NHTsbKHcNBHeYD2b/EpUZw1YsEyeb8z8
+8y9HfjJobj8g7S8SXDCnu1T+HGcJxeHrR59tBbb1bMypOLXMw9OT/suEkhUQO77
YUvGGFd1y2EAzdrzthHqjsRI5GCmXGxyokfZ4+sED9vqcD7JqE5ae0T5cH71FQGK
W6VvKmwpCgAxYu98azt/6G1GI7qWaT4DxAWDvAq0Oy08wuYhNjemksNea17kaWKt
zjT2NMDavcQ21/0ELEM4dlM/epiM72lw81xrvXZS27BM0zE4j2qTzYxoe9LvnU+5
G5zYXL8FJY3KxFlnY5RHoEAmOI/c34/VvUFfgGu6e7cppuuJ9x97xWh0PQOhUxzs
+5PGNFv21eYLPHdYrQ6dlUP5Cb6P6edIK7CJokXZuO3cCwF6xG3yXbN3Lm+spbYl
QIJrd9H6npP+0u8+OjVclj+cgGn0G1qNpWNA701jBJFiKse+sk3WaBRVu8DRb/a5
gRK5DQP2apa9s46EuHSHkTJpq2TqzSiVorQEb5ci2AwwPpiIRb3dzP+UxncshgOX
u5ky6Fe6kgs3elSc6D/SjNwR++hVsIZfLbCCcEcpBrt5dr5pYa30mRLr4G/gYHcr
X8uiKiQHXJp3bjutrneaPWsjiMY/PcJUzuqzAiuTeYXOcPs4VpZopIB1mAJkE8Kr
fDvxiZY4vBMFDbzBIu59Hvk8m7hWi8FmFnlrUEtIgZ5g0f4knrN3qSbM0P2qt9Lp
aWpWJzqiw7ST2cmqOu+bs5x8CgsdH+sk4WFCEh47g19YqX2pZQr7Dm4gdCgbgkKG
TFqKwkbIUiCrUNQYLBwye/Zd8SZ1+HyukpkeAf0wLY5UXafnOgrrt/CHIriJoDXv
54oUkQ+UtFc2xr7MXJ8OC/VHrVuS+mSJWifTE75INknYZej60Z2eV4Ue+4uoqoNX
jwbC96QMNt9wh4H2z75Yz7M19iMATPFZF0w/lmRm3XnkLA/mBJOz1/AK1HA7Bj5D
SdeyJ7mnn2MOV+nNnxlieqYzzecy3Xig9cFb33717HEPqGbqGqMWewN2laH29rHR
IUsrk4mD0dCR+VVL2VV9hGpmHt8zgeVAdZD2ofiOL7E8iz7KW6cRb4Oks4uXyLwb
rGhYqbIMqqSOQObzWyKo58fLPP5v5BvSUBzTru2GgBSEz7NFz9Za3ExKWRP1ndQu
zdyD1Qfan1XX+EnbTXKflhlJDWCrsWzDwxG/s2t5oKJtiIKiMx/7oC0GCdYe99Po
Nzk5aSq8VIjJIN1fl85agKv/QBVzynotVawBr4HfpaxqT5gHmgZUtBmf0Vo6h6pg
RiHp2B5gNj9tHwd92UPodCIAunugyXu4/wKC/SqnFUGqVd1fBiO8UcTg02LIJRd8
e7H3ddcnrJv+8VzXmOLEv6DbY0bkVKcbHBfeix8PwzLExXwUsmhrTAnnYCUiL+pz
72NohhydbK0ntPhdCXlAR2ZTcpVPNiR2xxx+MdLHM1GFD+2DvCgR1C4tlHeEMIph
jiLsk2obmRTxtsN8tzQ2Aj8iGKtaEz71NvYRDDMrBRjy8xi4nXLzo0NfbdGuoH2m
L0uB2bfxCRod6b8bklYmP+r1u6iGpPBPoABuJOX6ViaDVRCTC9dS2XozCuMafSHg
set9QQD6VDKbxNVXPm+8c3RVnjp61AhDmPFpugZwRpgULQRBXveDbflKrZoaaGzC
BzBM8t02mAeTk+DP0uWIUzEjVgVt66Jx9FhJuPIY2sKC0MjKoyghGBbw22bmJU2h
kRoUh7BOjUYq/+1icws7JyYhSvC9vnazIq+3V9M1yKG4Jszl3YmVe7kW64p5JPkm
LZVNc/Xa7VTfjP5ixzlWZM0bU0DULDcU2bjSeVk8BeOfncwJ8+1DGm70tvoFSMwg
YyClvjidt5Hwoob6IyiXoSFfxuoBhNRTU+T7HwvD+A7D3BEv31PqlNlgEnlpxB24
S479zM8aIp5GRKJraTX1Rk702J2hyfplOWKe9SF8EBt/81S4vCXEYOmalUXVwk8s
Ma/aAuFUhdfq959/tVYg2B3uk1E6BazQiQy8qNJy0JNsmk8xa04P4KIvkSLq3/iA
qqyIVCtbf+Fje1x0MQsn+bL26VyUGrszTU04jiiB47/mJQWeELTb1131iUGQvBz5
cyHB7ZBp5E2ZH75BTk5sKkX+U0SWF+cCt9PZKvQoQ26vG6toId61I26mwxRLa9Dq
24aKMKMZLKXibfwpftmhIROeQNvNeRwl+wMixMbREsUrwl8qT+Q65FpVuuEX6jI9
Hb20yp0iIFdJoJSBog9XkR1u1DrchEFmrBBCSuFDQdTwnUIwqJq9pX9xmi2yU+ZY
kitIi9QgSXbsAqUzAogtAbD2G5VT9RxmOLvKdSv0c39E4EAjgtahELoW4whZVVSN
XX3izpt8zeS2b1nCFIPrGw3iZDgxULRTk0sttOtLStP/pAgdkrI91YU1W4/3zImB
DoWdbO1QtvARHGPOi7hSQe4fItECLrB96v3G1q9L4RQbkpenqu62GiwO+7yXQGme
YRoiOHF+iQ2whwVpPewYcwze3zqyw+QGYRZV9UmnA0UWN4hx3/+lKRqqUKYOjFkQ
NRGODnEGZrU+DwChy7rVBOjS+Kj8TMPldLVZLbIgBcgzLdpTC7d0ht5+kglTFx9L
AK0XQl8jrnezTFp34DbPvm1pcETgkDywUAc2MvLgF4lAkKxrRHGNdMRv72i2bAdv
L96BMC/OmZWIIUisNjwDY5y4o6lEkXUuM2SLXliKQvdWnRSaXrN/kAm1Acqfa0Os
c6AuhVE7zphu2U8ORZ3rILnXvM9TVlbpFtrGULzH5kRtcOsuWykw11VweTBy+3+s
B52ZNdnIno1iYBBjlWihOjeRBnjiSsjsGgkK943yqGifJ4/TpT3L9jS8S3xt6Wot
1EHqHIUWOWvExdCiySbnjgRVnW63POKTTSDBK5MoqHzfNNBy+HdpkI+VFyAHLH+T
TeKvcDY6UfULe6hhW8prvrbnWHa1f1fugzuLxy9tZ03jwYRRxeLy8CWS4fMk9cZI
Nb0KHBgsujkdiYcOrCh9FJ8QbdsL0gfQfTwPw1QK6vFF6Z/inbL4ILtfBQRXxNc4
uS6zcB9zBZLvhu5rxZwKnUUxwGMawnzoTuqGpkauPl7DvItMjkm14upTdrmgDcvN
rVU5sWqrkGqwVVfMNoJ1+uVwi9av5MezsdGjiQZx4jWyN3sWAZFUSBqL+BnmaCti
1CqLQ9SiUsbC547TuSti6CbLpCA2xYC9GrM6AztP+YyzjdkMD/+qqCQAY52zv4LJ
C+5JoKyZMYXkGchADCgnUTKGOw0emM4SFhXppHfbp2xrpreHxW7BoNS7iR+tQMQe
XceVmqyLHqVFbPc+Q5O3ZOLOdnZEXg7TFMjghF6DcMQ8RNRZDpVpzT5t42TnnJwX
0cMDhFUvg2OD+FjWVxCJa/LQISKo98XP7keCuegiW42oBR3PPGlle6WPGLet9T3x
Br2SwXKypsywLhz2F5n9d8kMBiBqu0NxQtHThx1JebKo9CsbYUXps8Ai5lyXy3gj
gSV0LXEzD8Q4vIJpaFqqsQt6BKBHLTQ4AKUDEDBN1eMchTdFQT8J9fl1QiOL2Wi8
FTBx0OAd7miHY8mQJ3PeVoXTkcKwNqtGyeIi8ob/qfJQ7BmMQReIkYHTzXS2XSWv
eR/weJrpDZyVc/C8DQK8b8TYhrHUNNsJCXaVhs0leH3GgM/mbTsTE5qOWAbUd3zJ
X+n112z03M6M323gi1B+EWCGyxRF8cgEv45DqsFEPvpWWuaTZG/LKdNCjAAdxqNy
Chk39Gfhg9nLpo4xhXwAcUuhj4nwQgxyiqCtrO3iPXMbAuvc7NReFXueDaVYRr3E
GyxbCj/5vTGtVhmum6l2mknNfBsLmfeE/a31D5Kt/9U+UgAn3JgkdXXzq0Wu53Fm
+MPjWfnsZbnSSZTllhwHjjKRCSLazXotZ+axmsJ9NmcnxIqmQyxDySER0I6GxbGO
e0hHOo+PUGzQZNdTczokdyFiKYRBdW0pFFfihpHERulklKP8uWCTdTVgc/KQE9Xn
h0Uk15K/lUXPu0257+wAOBBdc6OL478dy4PGx2qGicvbP5qR1ZKATYqal0YVgWR9
P28yen/8C0NAQACOU7rDuDPupSKLNAtYoQ6qQm64htQqfcmA+w1UFzid7pub1Vwa
xLvYiweT+u1IR2/tZfbyR9rETFHy/xdcMa5gHFMiQ12QDMSxRkSEwqU0+0u1nHeJ
8HXHuU3iE2tChe0UMHJcNazKu9QyoTBsqoNSLZr1LgTXukAx/BpWuWBzIbSqHEZG
ro+0MXMIrRd1+I45Ax/OaNpV7F9bBTIfvWFgufbBKQ9mPI0HlaaLY0Aw2bdVM3bZ
88qcI762YXWbXiKQudteHLijGSFcOVrlFvTHRw21JI1rrW1um8B/tH5REh2zWJKy
0sno0b9fblD3ryc26gDZJuQNlS2K4ozlyv2W/fH5aLvABlS16bIz3bPZqskp7WUN
rRF2nzUYaBlzga2nt6QX03S/oxBsvJiAuYZUk+0KFgbx/Sg1QvSTgN/s8J60ScJp
w1Mk99TNezQHJPPsr3dgjnjX/7ObGNb7/dVJH4GrFI2Q4ncVmyLYGnhNjViRIMlc
u0jH1Ft/C98fG/9hYQTfJnTd/DffV7JHs2/eMZ3+AUx9yUOBQKQOqd8N6Vb+ocAM
GgA169NI79fXZb5hpyJs16hay/6XbOHnmttcrizr7xzfWVToi6RURcOgq0p94Cg4
4IC6Z2Hcro8gwXRhnddsCpYW1RIFnl7bOGZqCbuifnhldkYmND7alciWxZdfMkib
7p6eGAzcdemEGZ8+OAchkNZVgoY/vj5SjOUmBXPeATYMVmAojyAccgAK9wTnhEke
wFm6e02cvW1k6A1MRvaGyVV+RjVsyppilnxr6aULL5fkynC1mniySco9HEEZdnFq
ptJp74RASSm6pu0kMmQ/AvKzzyTxj+K7ZO4KgDg4oMnMt9IXe7MaqPhJmBWJHRYo
LEkp45v2FlG4X8WMUr8x+qP6bfI78rczVxmbfh8PX6pLMu+UZs48b10fMvILnZNg
sVIPSvtdVtOK67yiTTPGh6F1lVh6iTlrEs2XX4K6U47JycaSvHjVGBGs8GQUyh5j
n8roAS+JAEwZB9qaGN9oSFgURtYLm9Zuxw7WdPLkvJu3CjPZLoDfrpuhSyyDUaov
bv3xhnmT83G2QV7E5xETIJxLtfBfC7U6Qg7N7lT9XFXjqMXZrgdJwAME4ijzoxpP
jHdXptTfmYjv46LpkEJG1bhBH5Djeqj0wiYz4glNcOoLN3e25gGYOuPJPSl3Y0ne
9wXYhlmIYwpKya0ks/U9Zn+oD9ZMEFjyMhP4OtvbD4Q12Ut913parfSXbMg8/PiQ
SyJoC3GD7zICqeZB2l4+pdd0MDsErcQtOUkiOJT/ZEKnPJSMXXibgxHoedtDF7ls
jabJafREsqeoE0CTTWbw0yCCgvsgkU8p08pcUbEvPyX5BCB3RNSkc7rQzNnDeuaE
wJVVvbSj6rKC2LBEbqUmkfwlqs+qeCirlLp/tviteBgHoNRFn1eBdlFLfXEOOIzD
uSDzF7+MWdQQCMdxSRbPQMzycRMz8cxqlpy7hSLXTJ+t2tvwpyNYDDEN70i8YkK2
TLTiiQANBWHzRJHX8OcKU+rvy2Wtb9aKrzHNCWwCqmhtxGJk1R+cp9L9HMRQQv03
1Ntl/qQCbEI/2Fc1gcN48OmZrEljoDiBdz4XCHr/3AL6g8M8qeniBk15fkoulmCU
ob4x/EZ7xEHUCBxEdptLo64lhloonHYF63rhO3/HCEuWYMfCXkeGofxj3dY0ePY6
ER22HeZ4ErMLr9zld0j3eJ9HS7pgnk94mZjjbT++bUw9ZgS1rXNlqrUkMSo6LlLF
n/Z29znyB9hAWnh7f1TfrHGH4XbufZoa3Vs9ncA3E9FUiuar0nFQevuu7s6n1Z7c
ORDKHjuQPqWFrJ+DlCZtsLkZ25Rv7cxCLiurKBKk28ZImWr7nlqYoyFhlCdsbiyw
H53a0IetohEHjTcuaEzyzzbIsLLkvmcacDG06z+Q/ip7nA6XPU93a8Sp65PLMaFf
WxRmKrH2qy4EM5/fdRlvIXMBFc9IIjQTA7qoaLagGQpbR3b5zNM9XIO2KozIH/l/
La43YnucShIhRQgea+UdN4kQNUQ5d2kxIrlLixpVPmRnE+7COyI458cpxuF4gr15
aXRvettGWZIOiXIw2qhtTpdSmNgjqUbYcBpFaVL6jwQwN+Bdx4Om9CzhHRI2/uEy
Eez7Did3bzqXv9nnwdrXpz4p1yxjsmG8xB3HZsDkvlSVu3c3EP50ulk4gha/9V3p
75wTci/4HXVlX7ic2Q4rxWBBJq+Q9nksBeT2BV2nv13CtF34LSExCBRh/UqG8nGd
k/17HGcfuvlgMnePrImCX2ryWKIET190yVP/3Ssv8UrJmTyKP0BSODS04k2lMBrI
nUwaSWH73C+CslqAtZn1WKTrA1tS5TOXK6XiCvgXR/T09YLjD2VDdG9C1pYa40kM
vUTQbb7g2QweobR6Z/HJ1Y+970xT22CS+HLg1JHiS+ZbAEKbiqRTIBFRdBh2eMzS
VbFAXTg4XlrFor7wuoOU/tPLK8hYVvo95mLPMi9s7N/3ydvirTGKjx/lYx3Vf2G+
2ZYTIIQ0S1f37CK7ZA8K70bENlmFkxfHS0gefba17QevlzqsTxRWRbAgbjJyL+rQ
FV35YmK8IfcpoXLMPYa98J32DtlPA0c8lWLQoEKwR6sm+mCm6/ATeZYAZM+NqTvN
AmP/7N9ypkfB8qxfCSgGF9439kfUc03ClcDG8qHHKNHLdple9FCitFrzgcdm55qB
VDlDdb4uHNzegPM8Ym6LUxg5mF6mVuGCSX6nhLPacVCPJkTROYkqmUz8bmBks2k9
S6lyp0DfzMtd/X7l39YF4+MK6oM1g69jYmlSFHzmBEW7WHADTDkpgSRw2LtgbL61
TFrvt/5X2jS44HsbmUIeQiGMc0agrezEU9DBX0/tBG5MkfK5yqk83O4YXMkO0tP8
Em5vHA963elyEPufH0OdzEeiwcMbNIWsTsQZ5Gt4ZQUBuHmVyK59BQMTgnmU6qNE
a8qAd8pOheVqrgKqEJVyVGEfxwT9yteOmJJy0HrVSieWAL8nMN/TrO7iT0fC7QqA
CE/243vwxSDyIvAMO3kIdEhA6c2Qmbx+NsCb10xMsRMWUY/CTZjDridkcZrlzFGI
CYPNUiT3qvtXAfFu55JsXDiZvxmSy8t4G6i4t6Vb6IuuCNL65TB/pzUFwuF0I2DW
SPYEVkQUojtOUjHZbwvXXZR9DPjEGmqqmY6qmNTZbHoGyF+V6seUK4ZH2VpHjyrj
7NtADc5v3pPIaDqQ+BlaSND7KwgTW2n5sUudIfo9FEiBXU2/9a0UzU/f98JBL/Gl
y4iLe/YAQo2JwoMp9yIk/j7Pcc8J2M42WAOUPVKjNZt11G+sh9lLi2PbozvaayzB
VuA5+ZER8c8WibxkVtB3djrlHVGxJWsnHX4LDTZxKaW8aBT+KuazyAk7o0pEQy05
dLZGUs6nlOtNPCUGYtaGq4bEuxJ1QBljfulf4iYC+NZgUhOQS/cQu8aJBzmb2iXi
BdOEpyieoO9tnwO0BdMF85sL8GSvmAD7/FoxqLEWj5gLb4zkUzklJ7RWGiXOWinK
eja35aCbddlDOV+jhy0lrSopilPnNg5ecAlGx/LDQV0XtxsJXr/kKKI8WV26vwbw
eyG5PhBxM4Wb7ztYcyDpGMAuyWDbLoICO3zIHPYAMYaROJRjDUwmFhBmZkhBFD4j
H0ItVwlCAB03QZqnDoy8dJV3AfyX2YApE6zSJTvfIBEEs1PZj7pNjk4xnoyrl/TY
0ecJ/MdX32nF73h+70BufrP3G1NylIyZlJEUVBAOV1jrz4091LR8U7siq9bgE7Aj
28tSeVCfw4OVFnYHZDPQ1ytKN6sXp1Ljh5ZKPyVdheeleStXhMVaKTIuzcbYEMi2
dEvpyLbyMY65hE+1N3K6R8KrM72IKHIzvXCMw4AGW0obI5a8egOCi3RBPJgUr+XZ
SD6ZdkmnjQNXCblop8vL92WURleE7aHGd65iODqitdP9W+I+4ycIpuMAmTksFZ5N
D9z4c/1rSyYmspf6vXGvsacy07mKVMTZPuDkQGkwHkLRopoPeWL2QjRp5pkCHeg1
9OPehpQOkHWhDWo4hcdWa+iVhKcM/t3Ncdx1NWCbnKlyEn6x/5HE/EvDKwzvJaId
AUriDGq5HlyyI/dF2+ao895VEF54uy1wsWoDnTf3P4ZiPtg+yH5BM1qDg4eLA8fE
YCB9ZJ/KQwm20f5mh+5QA/y9Jo27vdZasIoFoRswOu0LQ9BA0EGNmHqFa6yVv4HP
3YSD417XPiVJfx7lGuuVfM4lXH4NTsK0DflvF7nBDWG9Fcq47NfducBJvWQxanwp
BuQczwaMRZ+McYU3p9cU2en2Oy4QOfERUFbHTqJAJqoDkHPQRqa3ux2DygZRU2FY
ruBNMwtrzw88Hgl9arZElvf0SxPQL7qFHLra+ELDdgOb36ldc8yIeXUJzlvRog+I
cHD2hf5q5rQEcJB+nVquYpbFovjNBe6k3LQF66giBEPI/oVBq+eOV9LjU+w1y6su
UiFr3IMHNH2/TjFY3QpHr/wnLc0f+EKWTHkCa2uiCTG6nW48x2xFZuYFjvlLnywH
sWKqa6XP2wuA58SuqHde49x9lmAQgB2eX0W7YNM2Kwxn3/SDxvqO/HNOGH+ZwO2o
uuG2CggXD1LvLzFA7prqeorDv4TpiGUref0jJNrpurQLSa52sciE2OoC/MCJyadf
mJgDVoGk37mpoVgFCArX9yKOFPyvEybxzV7Rlw5Qm2+da1ciMSzfOpl91vaYSKHa
jijc0w36RYlpnffD+zmUz3Pe3vaihk+GgJO/YdIMzcRZie+FbskxaGCBoezLoRxW
b52I0BfjfKMoXNAdllMjXLbm7SQYADGdOz76lAV3AbsOEsccyudMk/fhqH5dgyJJ
jZX5KpXqhx1Ia9oY++9kNCXiDsh6GYG1qOi8Bxw6ZubJnZMZsBjTYG+1Q3BzQN2t
JBYg4NTyYLD5vOxTHlRFtBC2S7WBgCxLvTG3EZxPT9DEpBJ8ZmCSrIpOHPazTX72
qfUvNJ4Icj17CfOuFLacWSuBRufIKibiY/8Z6ZhLxT0g7WyoCI2uS5LVb2/qh4+0
jauUebJICgf4KusWrxvzFS2+Z+YnIyPrT+KH4/V9YS02MEme+YfCf/e7CGoMdbmj
w4Kv1zrVUgofiIQ89DiHbT859m39O7c84WVUa9LjfifE+T3TuyikJiJJ/4/3IJMM
W1gvoBUWzw4pV7smQQBB9Mpq8d1pvtRlPh2r8/RteIc/pfo/+zYjkOjnA6h8eFc8
XBZdvK5+O5MFRvpT64IFVTNqTJSOldP1IXbYTb4MERugZxcMvX9IHHrjsKb1s4rW
dh41xaxu1kYmCPz+P3zhGPxQd72+9IOx4b4HfCVJRNXfknkP6fnUTZi+VA55B5Hx
jN5VCG7NiVp4I4ncedO2mYt1qQXiIPjRxXlYF3nEY465o3Q0aGvvNYUlX7Ch9K0x
c+rg2N8FlGa4iZM4kehsBkkQnac43sPtBKHrC9dwPsN0Dc4MvXOFF52SHKb6CH0H
cdS1AHY0mj+M0D0TCiBmBW41vJ8ARQ4+KsusdnZmALDtw9iUrNSgwmxSc8BW5hOk
sjXHPCIUBMDWpxXjWirOAuJHFuooXyd+xD6mqW7jUv75xZ1lNxgjw6JOOFWCTsAW
KWlVeZUZaJsGx6Tibq59HrLOM0bJK5wOCgykMCnEsR4yyc1tPN9G/R6j9a6gEc1k
mBNZdC8NeXEjpO4BoiEBAwNGMpquiAqtSgzLpPSBffOC7WQhx7v1axQ+SXvWdzeM
Rp5hIYJnFY+NQyKHJmsfuejw1RBSN03mjPCJYR0pbl0jKfcS/RMDjYNe9/BkeQze
xNJmQtsqb6KbymeCYXv808HrQURn23Y3TnLwvWItX7wZrjvquBmu6FEJ48g3ykcS
LeQK78Qh6KPBT/V7BxAlpRn9z8RO8+hFn/KCab3MQHNy7EpLfE2pMX5S3PTjqJbM
jpXe17KAf4IZpk+ZvmzCFjH+8E3GMxM/5QhHdBgCniTZTWMRxGfR6U/1Ch78sTon
o1QdzEz2/1vsXKIUFMoTBH5cgbhbd3fdr/eSxOzT6CUfCFPayw7ExjjJfF7urNd4
ndzx8Rvj8fka5XZgEiNfSMdCkr6XYNbHI6Sxq6y9kdCs3Lf0FvuJSVWkbWkq1r0K
oPKuj8h0xeopB2OZ9UGrsAmvr0xZxz4UfQcu8WO1JgA9yndw4r4iBCBLoT+I3ZN7
3j+5MvWXhYz5a4QrX9hX4/fD8oEP7YoDlsrrq/LSC7bL3+YSQ8+3AOQRYDALRaMe
7ak/2kMTmFK0zXtO65n/uuc0iZu4rBNkPzBlYugLxaVf5Jdevi9GaEd3ABheM3iO
e90eTWDRACJlm3+7RQecK+O1lTdSrgema9Tei4SfQjBIpp/8tLGHI+eq/pHcgcoJ
+D08EOb/f77KhHg04TWQCMdfcwLkxniMCPMFiF+gxUEpLusuG49WI9XgKaqO/jev
ZfIJISVKw7pKLpWW5PRE6CYM4pNXwCHSIjWSFDFgkyPs9UjSOLpaXcpeJGqrfmVA
lt3J3nbjaHYnJCEUXGvEBDOQTL3MdDL9IKU3k5bsESifEr2bt8mmzOH2GZX09Ef+
7zcrBMtpXHA12Xc8d5dw7uHnqDEAgXyq6957GhgL6iviZm2H7+jifMwMi+JSbMCb
fsFxmmUAjbPzN9Zsn8M+27UjvfT8WWzvI+pMcRaNYjcNH6/LMoUZE/ecHfgREL+C
Mmb7Mk5EFOIQtq57tpkP2rcxOnwMaVMhxZ/Tlm4iVQgC3H11tWdqdyAXEbcyHf+t
nLJVj+23jay9UKuxeD0DInJKJrBoFlG/uYedyZhEHRZnRwB+2Yfk1OqU/8+gh77A
sLyPS5Oemx3SCekSmPj5lbeDXUJgZ/YiNCr4M9zLfFRIMkzIX4i1ZD526MDH8+xs
CxExK5S6XO+yUqPZhugM21RZPj0lLGjX3B/z+PJZyypKAbLCBlmuRVPRipVHwO9x
2XikVSZABpDfTec+u0Z8+/tNMA+Pb6+Mcn3+rAR+x6JELtjxIlO+0hv3MfQiYZXt
mz5+kSh309fHh4i7a948PMJNbV2Auv0mGUY1oTi0ljq3xhz7aV0Dnq+1+XeiGMJx
WMBua1DKwbTAuHw2siROCiqe8gMqDW/BSt6Huo4tj5QvdJl4x87fjA1nDZimbylg
BMw+NjvGXpkdxatMOS2hXVNnY3kE5JX7G2X7Q2Dk7RttbonyVSOlZ2oBp2MMFdhs
KwnIW032QeJhaRvJDgYyes5bDkz6k8RaG5buR6/RzaxhI03Cg3T0LWwiKPaazmsP
ARhvfZ1wCzlJy4uyLjhMEEsSmQqv2ctbrzxtVxxggNbbVmKYGpx1nyK3/BfJul1O
BiWE3op/4tr0BBP2mlVtY64CFhgtLZvk8zkZI4NzHIT4UnNwL8nUVixjIhsVSOYT
ol9ImFK2e0pOWf8n0ie4MfPOUHHPXgjqcPgk1yFyZYhBix14u4UqH46z7dc3OxxC
Z6Vbz9MRoeO0bCZcwsbO5DdI3egs5Md/sqrx143mr8A58c5h1vpXRJamCo/eS4lr
/3xTx6baM2XK9qicLbknRc1pDo95GmZPG3odhFe0nPzuky+GnBFIjX4dyIEYYdl/
jHk6zyuvgK/RPfSql9yqro/paBVXpWMYnIhmNV1eSRW3UGQGr76VjwaKpHsvO5R2
HA6K6kpOSkB0TsDX/bU6HzbOPBtp9f+lz/lU2v0vGe6V34gmfJwmynV7tbYSzieW
HyA2vRzySMRY71wlsJPmXU75Py9pLrwwz/1s2rUwRI8LxJInuuGn1PyP2id4SH9I
+xrkUY+r0H32DujC947kbQVPTF+y97Q+eDtYr1jFOJDj7EHCnCO0PUEJyQYc6MRK
KMN+takb8aSBxVdIxf21CDOfXE64wq7l+o5q6S7dVS8Oduk8Bkj/5g/C/C1KQNCF
EqCwFMO1Kv9gz5vtaOdZKjELaN/zYa1U5t9pGMUNngWgHyX2Fabya2FNfXQuw3mm
IwSe8ydeWE/OYXdNvQT6Sf1iYXcIpx2HOc3k2XEtVMoijvNIaXUZi6fPqO+7ZrEp
DAUbvfUSUdKzGzewjHSjfhl21jKODYTnaCXG3T2pN9bnZ+N7opoUjKlRglr3jaBG
oy/YrmpS6rh1oz2yx6vAN8wz8xw6iJR7jTyRio5YEXiNaW3OwLDb1S4jaJkDzXSd
s6C0E9J5vNMDBa3e/FSYJa2SKBnwBwXcH98R5f37+R5PBIt/59dna03dfUG+eVC5
LPRwcKZLASjG4U9eNhHq+iCg3E+QZMaHFZ9f6s5FyNhU8uolzzG875WiXRHwqrDa
PIYEZNy85N+aDCfZFDrUUZxJ1MPM74lRV0GjiH/oDE1tS8TegNLrubpNYrtQE0H/
A6xBvn5MFF8GzEu8bRUvzTWNCY/MgrOg+KxAHXtUr5/c6uGbVc13QgoUeLexY3bg
wzaF5XvoFIyrIimcVFy+gdzhheaHDcDZ5XIuyuTk6IBz/NAm0lUCYwnYgcw/Wvui
ryrzI0EbD8GfAdjiw129fBGxMKWkPWoy5nC9lWsXnT5jW3kepgbnWNn7pAeX8KFW
Ylk0b26mGE62mo4fFZiRI4/+U8siWh/4mx0rHF9riigieJiwzjKfQQdFsGftxU6L
7Y6kpq2lvovrNsitc0AZmszk+V5oH16SU7SlhLDpIvoR8a4AYV9e6iE7RBXDr9Rm
X+Jwt6vaqCRdeb+UUxWvVO6v1RJlUUMxbkfQK3yL1GqqXmytezumzyxoj32b+Pu0
AX+xgacntYckTYIcaiFOUDhZKd4IrCfQ0Pd/nJabBzHIjUp7NpRp0QrfwUTcYNuF
Cbbcn/eM+XYs+easdkQcVg/GVPCxTrsN7jZFcAxUMfn6LQxdQ8HmThoS6YpGYTHu
Ulz3QJH600QkXUaB0joUua+TD92uHkDMmpWn4bNW2nqo2XdU5Hf65TKCFkfYWkNj
5RpkLi2eKrJ3CXKRaiQyyytRRFhEcI1m3cbQyAqKPt2YzISitgVuvkFVAYJLKbo+
4GQNf9MmS9cq39Rkq8pEyaOKMHh31d8OMC5VVD1RwAW+dc+8+C7TCGM08j87Cohq
1qBlY3R+fKjB7OMwrTPtWjmvDgBWc3nqlkR870/MPlD+9Y1CrzBlb1QkdqLn8uRp
Ktw0mIDi7Em4Zh7E1AXpKD5ii49mz1m+Gdnlk2rT+4QFVtCqkXGeTbP+rQ8SDIT0
Clgj+L+Vlj+n7Iqp8jr/nnCnYm3d+8XszydwJ9DARwd0tvJhGwqXdCszIjeC8Zj6
lbXEqczjDH0h7g3nc5IB8mbGyKr4Tn/cj/vOSt/2lQKZ9ZgLow4O3//bqppSUeWO
v1SW+AsgNLZuIWHTSD5hxDkMY83zmo6woTGIkevukpDUzrM6Wo6N+O4xIaCK5z7f
nKlCaeTTGPpLMcDCU1ZFJUHDQ/3tobL/cenWrE4AwecmovwpuUGWk7aT7ObijLsJ
x4cz5AgHarO8r0J2knsNfPHzzKyoxtNC6z40EvW5RL+SVeb9ylnqezAGHz/1PGWC
4UGXmnxv0UxXhlzVZHM1771d7N/K99YzqJ5/H4HYg4WuPkL0AfT4jDTgBYiXBXdE
4sN94uFtGaWEDJJs6AD74fdBKstet77WPamc2k9VV95ramQouUv8DMMDlK57uXPS
aAEfsauA2A+YPyFz0IvCB94m2HB54ysVAiQlG7T9Cvi7nOYiuwZ2R25wQvlQSCJ6
wTNi23J5VarqPElmx57gj3+KOM4ypTLLOF8dU5mbNFIZdEcM2KFcoNS3z3vAzs0+
SRiDLn94LkulIUrUC83EWB4qplkUY9K7uAO5BSxtHNUBfLESj6LYnnSU15mGmY0M
zCP/ermq7cFkS4qOaUmwJ0vtLFoX0pDiu5GtO543jeSOri+TOicSLGGQvYERJdKC
d7IoXt4o266G79o2FjHN6PRpdEC9bfYHRLA42sSaZH6NrrEaT9K7tODSk6YwzwK6
FRMPtdXx+FgrlsdJMxB1kERevcfCXzfLzvxeC95G6oId0StH5mvCbSYI43yA5jcY
JS27jcrReOxQrQ/0ANqeozzOhBqZs7m6WCSzBCsSko5XSjeZPGKTbCgXYROxmvHK
JOl4dUXrG57UXRFH+t6OaOA8p6KuToVB4p3mO7o3hK22HfliMtacD8fgXhQsQ++S
ZbDly7YZQf7aMwYtcwyQ6/2in2neB0JoDKxoBXhEAm2sKQ4bLX0733MBxNK2FbTL
ckcZtVIg/rdlQl5T6XggxkGYZ7R9eNuXr3QqQZFQPbl3AYM7qJfENzq3AYp5LHiD
8qmYH6h3tcOwlk1b7Uj6c7cp2GjGpre5SqAK44V7YaxXsbV06e7a2dpw7K1OMp11
nypkEtorteuPsVQWrmQHmyoM0B6ntKDN6AtqAkiMGsiiN/M51d3ZWPbsJhKo40px
mFwn/6Qct0cNKoa8BYkfUDg5sYEsPaDDHQyZyiVMK4yI6JoUgx2xUceKFRNUwfAC
fCeUk0YAI1Z4D3pfFXxk1DlImcmgQdGJA1QJJJ+wemoNWzMNlT0Nb3FFY/qKsHCn
Xrub5EFnzwDBrvV6FLeW+JnYWn0sU+90a3mYNaEVi/Ic5bioecOiP8pectDSc+GM
jXUPQwU6XhY1+tEX+/dek5H46p3XxhVe2czjoGGQ1j0YXfJgaMD+U39Qae+UJOz5
Ui/qD68bSI8v/jD9vGbs4KiZwiXy+J8u+uUeiASuYJTEMxNS7YLOjwY4kyZDgPQm
5qc1C+Rp0ePewV5hOMMmSNxxNxAPMCdYN/cJQ7BvxmcV1DKx8pdncKb1zFXhshAu
WPyLw0MhGyKxsyjS21s74w4gn//xPXVN1+9hqygbQ/wL7Jsq0ohR254hNmH0nuo7
q1a5e0yW/Tm8TaUHJXobRpugKfoL4O/9AbhwrJX2IDZPAJ/4FTR/nNZvTKa93K0y
I/0Q6GSpKOjMD30E3KaMm8wIopEuaD11X8fEJCZRyK3OCL68/KAqwc9L3vayzbpD
g5SfmUK35cOWsVa4XHUtZfPjsv+Cb4G5T+Gvue1hrgr+oDVb50COcWTv8EiYRliD
Yzqr0MCpmSye6ZlLj4RJiQR+Xov19rIWHJggWtqXOilH+OQuzsN/nVQ6droxduMh
1rDJF/3wE/gUkvBC/nbMX3kpJa50ZwjGda8kQJaaC2pRnnZdjzMYGuVX+yJlmB6e
8/YzJPieVjyrJuAXR67nK5dB5q/DjQU8eD1qtHn9FtxliduM1uh85S1iNnmhgs1o
bW3d39/CdpHYmYxq7kLs1Ju4LBPNMAg5H8LKNHRu4JFv5eFt7iSgpGwbdEoFroma
9boKVznG9Q7nhKeAIl8IM2uWt1uPhIdlgkY9tf3aV++BNGk27/RjcPF+LXxceIEw
WB9gfJXbx/+JyP5fU8K1NgYbtQNNuE0cLccGSDtrqBm2pmFhgkmqjiqe6PybkaIn
MOxFdRbt2nACM/Vh/w+jkDQXSiO12RmZyjbHclTfBP+tP9HK3vdFL2GddJzHUr6j
dBOQVS14r0NP8+CzSB1RlSBRUDaE66vHJJeM2UR1MxkJq/WJPInap6UPL4znNImu
AtxwfWm+7JsL4zM3A5l76QRBglUO0nLq81OFR/9u3C9VsWdTHQtHPUL5GN5xmgSs
SbpgLil93hSZMxYrbLlMO/kOvqxD95ipecgdlwu5DJODEbmk6NA9n/NTQOW6iM37
BsP68AbelFx/FA4c9AkLd3hSUE2feTrSc+XyrXomIBFkIlI1mjTd36iRINvSivLM
t6Pq8Dl8Uhg29/oYTqDW5qRnF3G7HZjIb0/vZuHvs9p3ix5HQ6Ydi7pj+Bi5Ablw
VGv2qZhJnBH4e/N2fGqTj+6i4yw0ltHEhfbOCgwxS0Dp4yNIOWX86BFFEkRLls+Z
lMBxUg7qw2lD03loccvMeuBj4dUkjTg4/QD9ufcejuITR4nf+owtnnD5VtwkROMW
nV/mZuVhYaMR4K50VxcvFUT6jhHt9g5JS9B6QtCtKPiMn5Bf4MyL1ZGiQry8mbr2
ztUurSL2gK+eVMzL+rVQkOwY25v0njAinXkc8qDcS0ZcVMYk8/8iSBZzsI9lprMd
BPupCAKGRIraXu2gkxBd3gOku0ZLIe02sMLtTrBF544RiBMYdjeoAby1hWtp07kT
k8KFrG7+aPL0+C3vAf6Oq0Qgy+hCK238bB5GYIzxNp3789CkPLHXOnmfoappukIi
2kgG3eZUVZB6GBDfS+RjyeACQZNYx60iK2slTVylnWPU7Y1/h3cjgu1oucOVFrs0
fO2plXROitUF+aWjY5ygNwsXJJGK1uKHMl3IoR7qNLL1N71R3CMUm4DQRR2MDpfP
YGYp55c6tq40xNEDbw1tPGHOK0pi1n6BXEHvH0VCmqw6IcLJwSwT9VERekAPR1rB
O1SljX9pmmtz+LZw+BpyUw74or8SHmJkA+767FoocRPW+vB4ZjJ4G9NjKahHCzMo
xKq5dcRlT7Vaxk6oSSM0vacmSRZRrI7JkVYGofUN5O67aAoEKFj1sahhaUiWCzU2
yfaqFEXD/w+yKIikRFolK/Q/21IWnAvO/4jdFNbGDIR6QDx2mnDEnf0EcBLdL1jY
5r6KVP/Lxn+IowZrwFYwaHPCTE39QpWQuFqCy4xUcPSFu5QzbEPBzV7Uz3pzMtsc
YpHcpWORUWuHMrmGKqYt1mhoAWVM8vo98XWIg3SvH+EUNsc8PTpo5EFUOLtdTKJ3
pgMPnZnJklVepozHBW/0Ukewn1QeSkIXLoExIcCIiUveYohfC6FwUATO/W7kXaDs
7CFP5kRtYvVfwFvjKG1mr/VdDer8JkJeQpsWnOAv8+6vh9WyhBY4NNzWPt4K4ro5
2SgOA/B0EMC5HTiKIELClZfNcOYftd0yiIoOcLD/WCgqKT/guox5xyDUP4ChvTUL
UF5QDSmIh+e2PchShEGDC3kxsf2ZJmtyW7gQ54ha5kzDtjPnK1OYKFahuPFge/aW
Zt1s/FLkngGXJIGF53fCzZ3SiAgJav4nYEF9Wq/H3LLAifVx4o3w8bRY9V19SW1G
U/X5LoNMV2vg0ObHo84Cc2RipqKXofJepPOpPjW805PoCNZIsgmYnRXn5g+Y0xlV
EDCUUORudG8p5tv4Xhi8ZiRuFTPfBIW5aYgkufW5ixf3/2rrAW1HUq1JSE9eqpIz
E0HQH9UmGnkP6lUJFEIeBHsyyHOFxRoho16n5Wxq6t1NLxCxd/IJqxHnjBb8IbFQ
IxXxYJTRLC2XFl2jWDcli97pMTfm9MgSloo7+8J541KEkjI9jq0vT2ggWkjHFr43
0U4vMbZLDh0MhtrJUip5OQGz4VwKwplJF79KL04719kswX7Qbs57uNV4ss83A2Wy
3s9ggqVKJpcn6LWEbi1Zm0iScbBYQbwWfrtHyOfihNQXzxe1ZpCx+40/0647VU9H
9C5grg07dfAvZxKEx7FXIUMIYGcAzRYtMKecN8uENDKtYI/6qKv6lDPOv2S9IP3j
FUwOW6zKcbDlmzZ7Wj/EM23i2vhKcN6dny21uwFE0/idpouQURciL0j0ewIk88Ii
tuIJmb40+uljcltg2w7oSGP/W51X8qpSV+rKdro8Mdv+RUeQZCHm5PyM5aHSgkKu
AaAchr3ouqmF66hGSAyvbHXHC+uV46YrxIRI0B/dLvwcjTrBeKFQPZYSenGR1kTZ
PjCRb3BIPm8cj2uaSTGFC0fKHOwnpcqO3Kmsew1MQ4ITdoIKZokUjkyF2xzrnKCb
4y/M4upOge57lNO0cd2RMxpGmkf+FSNflta1AZemkZ0EaOztnbTSqSDRHl31J9pa
YaLxc3WHBU6JmHBguxLWPbgb49kpl3+ksAjEJx8PjlMUDmukx2mN1TDSn3FDXNaN
9oG/rvC/Z+875y2TY/ZYAgGEeAjvFjy9qk1fkLEDIuIu55/0cQLghLTFTgsLbsLe
jgDjk2rQlIv1UUNevWhQ297L0+VyzeEr90i4bY4zQE9Vcz3Zz4piBwy30sb/qQ/v
mW7PPQGV5AkxUVPq4FJGoSAhjc2C34varB14pIhkw9j82ebT6I+qluoFpKNlQNNO
cHvWHVWij6SjrREp18A2EH1iW0DSXlvcKR5NRavgbjdlJPV/dfqOqAZqSb7iAc5L
eqisA2kWD/DpT8TE7EEoVeIHuwUVxrNJpkU3XvD9jyocHItFK92Qj/ZRVymQiArU
aBx3snI+2mvpXDd6wRN2HCmFqL/JGTtqqIcalTujofS3W4DfHQTvh4YgLo+Rm6ZE
Y3OY0oz5VEexA6tL92WGOgCeCHeQpizXpubROXtLRUFdaZxg0ArkXFE6uINNMA0g
0PoUyp1IcvgXB0uhYmV8EW32Gw5LbvARDpNbTbNzSDFszZuGKgTkN6emtiQoqaJy
Jn+ruN0lJr0FJFN/uzbOxhJiT5avkVY67B6NyWJBorFSfURyqES6uyZCaYyz9Ccg
05FyVbjOMhRIGAMJ/vhSDbT+GaVs8WIZgzNL4qjhd55wzBq2MtiDjzcEJZ5qXoVp
GQ75vyNB1po8miJbL+c5MdFIhmU6yMLejPRE9yc2uwFqRQ/reTQsXK3mVxF1lO3x
aoDLHzVOGK2wj8vTQrrWEHYZYbHw3hT+B4WEYLjVnAx928mpe4Cqu3lGn9B9iL/G
L9p3wj85vJVQ5cqagKhNgw7Aw+D48hWP3wYEdE9yhKi3l/xIyaae49vYN1L6uigV
eDq/sMslP73Wt+hPxVKsNDdktx1Tk2VxGAIoXvRP+gAXuvHYm1VtWjSLUvNqow+b
1PRLUW4+H7zK4PBc3ulJHPJOHV18nh3Crij0NbvpnmLhZTXpP9fE8EeyA61i9pj/
EgGkbtKdvGAZXaMtS1T8KmkUenZC3dorm0u65ykL8BpSwseWczV8Szp8aNfP4iY+
bk5jo1XrliwAa9228U2rFiDTjHDQkxWqzhKaSL1jEDZn9dToeMpPgHFl3KkwCfyd
2jWEPpHQQSwo4/JJIHiaCeBsaYgey3V9vJCEFkQkTRc/ZaQ3rCmyuFaaiKBqt7cf
JQbES2zd/rfOy9HK5juBt0B50Rsqg4hkR612ifSeK7Z9eYLsCsItC2On2HQiRgz4
h2vUXzJXfdZ9WjOYN+2xnF3zwDX76CGrsdI30vDRU7tML1DdZDEjkYTP4NyawBMB
uV9NYdBGQ1guWvuNm4oUSH0pyyZGAGaUFKvK18Y1dSBN3Ry8BXuQDDXv54uupZwF
o23PEBI27LKXfEx4TL3X2GvtStseAFqYlpc2R/eKtE6i7W0SXPkG7h1TnPkLC7xt
PQgKmeGcObFQ4XyBfzRLU/e0QUwP95wjIKkwLgN7oiKKjxDE3+/x833cnf0qntpt
CtcAryunexETaW0YY4cMAcek8Znc4l41F7owV5vEcNU3zE+dAhC8HCmXGdt2G0/A
Q0Fo1QJuk1SAlyMgRhbxCW25T794BJYExnaG71Gg3/UPAWc3EUJhtKMy4HhNVokY
j6f1y5HyV7e8eckVEFoKI0hNrXsD+4bucTlAa0oarhzq8jSag+US/iX0n9bqnSpL
rOR2CXLKi2nPCetqFP0shaQG0YWfcuewg/WSnkKtIrIjsZYdzUCKHeuk7kXX0bkO
/cJnyuwebEcUBLBZZRs/0rLUQzjIWGK5/6hA0IG7mfF7/ZUO2Y+VxnrGq0SzqcLR
LXtAopAJH5Igq0DcwQ3F61h2ebX5/v1nKFmSXqX9LBPHNbfYHUkWSqLnIA/3Eyy+
8evntCWYidMGSHQI4G3KvlkVfAANtI8Uw1IakZ8GEaSFpYd+PHDiee5JBrssq6PQ
kbaN+/9Kv7aGt4xJW3g/6WSBH6jCnKpWEG2b6aGddgM8i27V2+4nAAcQXglUNyu8
ijhGEKYYoK0zOvW615/VNGra1cLc8TBKI0zzNeBPk+UhRkpHJw6USa5jnp8Jqux6
3t7JqrksnWX9a8Sh9CWFyk+cPng04LQBohvq2eU6hWKsVz93JjenPRtAu39byo4i
1AKT7WjvRErW2OK51cHzcTbHop62480bqzp6WhCBbQLcUlMXVhIRzr5apxDnI4QV
lZSKAXSGyRqyGlrIRB+RIFh9gFQG3ebx/CAlyxOkSek7PQnMwYG/HstaV7fWSRYS
59Fp35cKXAoTJbuBlArRmZezDhSQj8nY79WK+N2rrrqi2ZNXbe+WB91zG0xqNCvB
/cHrep+i4rkAiLczL4+XsMPjZJXKP0aOcZlW/Lof8Ezpg6fBZShwru5KtmMtcrIX
mAPv294LB2iscZ/MFZvG6q4iblsdsi2lLghExoa9zTzJeKrAIWBIPlluDMTemnbt
rO1Slj4SRlTkhanOZ3kE2HnZ4oN7aDCbKTplAG5vTgvxIz3M5m03ZEhltMIHL+L+
ivPBgY5PtramUtAa5ycIgcTq3E0J/h7c4KMcJy0mgmh8wLKIvdO3dFb40fAkpxcg
NYKkdcbGbc4wxrK9nJ1qIp/srpihGRDtJ8F0sbThQQjAapwJgWpviOT4MXgdaT13
q+or/AbeAY+lDNnEB8JnUjmxiFSkuOE3Q3czzlvUd/YUxQXpLbF0+/lS9Ln+4hTO
5UCUf8xfGrcibayXCrJ19nvpuC+Ge/1LJb9BRtOpGIwLG5heFPHQ3m4GQM+JW46t
v16eb4zNBgBCRgO/JJwZhwvl9n6ozX4XSue3nXS529WDkE40RLyM+u6rDb21adiN
UckBKlSdaYyGlqFovnb2qfoc3GmRJ6ehgiKx91NiYvz/G+eDEsyLh//25ACqq88A
d+44fea8fSPMRO0rOP7OzALPCcgJbHpA//2cdMBvjMlLB5FdE1WjBPzmZlCgrdKT
PsnHxeXcPXov/4SbLq+9KQhjsJ5FI0uGS317YOGScxV1dC0/YoFCSRwRBFKZ/V+R
7V8j7/qJA1umrqxP1e/MqLpCKn2miCoGX22uiEE2QiJgj6ECeWdFkPmrfU7xQkX9
AcgqpeeczEhN7cG3MyXT3308W9y0ncqAu89Pf0DU0jCH9cHek6vAWfC6ygRbOKDy
KHfUzskfuJO9J4fOTbv1/bk8aQ7RRCUDVtaJFZKvZHmjnYkPYgP2Dlbb/Mw8LIMx
x0HYVTQ8vWNSFHTxqlrqj5792q7bkWBpi/mabEoM77A3p4QZNH3FMjvGclGQ8iW4
akbwJxY6qSNLpODYvdXzd7uwb/Q+1zIttis1XNQI8eM7NH1EVwL/OH1nWeiAl+Wu
GCxyTVr9pDnw0dxPpNVWBkxWxA3AzbI6UziCLMuMIUVhwJQ1EbhY/d8jPCKNCbH8
rUnNeBFH4rp3oljLPBvlbKc/qVkPc7Mj7y4pi8VqUBScuCXMwAdfNaJnBPTJkecE
jqk3QiLMTkZZFwjKxU94WHwGk0IIXJ9hiX2tx7XZrZU4U2Qbsz+czIPi6IRPm0jK
6Sqx/f5Qxly3VaEH4cWDHPGvpUoKUIZ4WPK429u4yT7PzM9OoIUHWgISeAAkMF2Q
GRx3NWHJpyjdP786Zkewgz/xhgM6bvjebCJG5yn5dq87BL63jtfVU7Ud2KzlXMGK
0gxY3bFvlWpdIK/XSwnGGkMQOwqdA8Uig8M02iJaY0wo5OlZpcBUO3IVDkQbdvwZ
LPWxlaoB4r6IeqbQEzAdfdK98KvDzIV6dI3taOrcg4MDtjVefQQxu9pXYZ7YU91J
y0KPcPfizurorKf5HR03kFbhIC6c4kLzmkwODnz62ii7H1/ol/MHiLvOHZuTnGuC
347FvCoDenBT2/5yWsHIYqkS6zE9Zl4wD5ePdFG1mH2D9ldOCDRlhsONRObiLC9p
it96MeBzjXChtSHFwV4TMDWLxbYZ20pZJq3MPC4wW2p7MVW4B/BBRWoG2IlXTxEc
kGoE7KYEm+FQy/cxifetqpCrgLrO/sirK+0+6CogrO650QUnZmpevDIl0xT7lVif
R0of6EAs/iHhCwWhcVutnwKSqrubeRRP8cTJGDgLZVuOsbzBhvLNO8vAiHaViBhA
X/qzw7t1hl/y1EjSZozrVBrHIoaIjzfb94NMVe/MV/dexYIlepNsyRnI7A0A3DTd
RwBOjOid56ixJIn0yph8xwNnT67MXtANGtiDRW/wXRt2n2fWWpBjX7MNxyQuEOXj
ISqNErfQaFZZbnNS83p/qg6pJkG+YcPnCTiBn3riMSkXHQLGlDt6KCAvkuhDbLxa
ShqwE6fiiApr1VEgaAnlPsV/rS3pey5gsnb5VLUdRFCvCCnTKZBErTB6li97jW9Z
RcWEND5YmXAYyZntCIYHxP448Ur3OZtuQzkzuiatsEq+Suym3TQmNCqSMxdYjQgM
SAsqTn+q/IwM+TQ1kpMXCQ/xTmFiSwe5a3DDx342xHNMib9/HRzR9/fd3x0V3cz8
Ssa8ITSfizse2tXCc5RpgNTMHyRWCmqHgDKqoHkZhSFFVU5eZz3yuOLiPpBJ1ap/
Wc3lYDCC7Yc7OxKtiu7oh4i3GtyCAujvWR9H45lTAr2P119mxkOWh/K8Y46Pm26b
+eTYFJ9jZxNVQu2RF8SIBX5Xi5S3vm34K/a0scHp1HhzFSlUJ2UnMZ2Jqs/wa2ge
bhJAaNcOkiYDzQwW7X6y55RQO5txZZ9hTNQgD5Cio2AYDAE3CFhdLbFxE1J3DIWp
O8u7Ric2vTn0JWfl8JGOr/OA0os9rQwe2cMSivKhi2bCfIkvmepwgB7JgEz4fG+B
yJtWpvAjY9nCnxjNBDyIEgq8fLNa9Vm91gkDmggPyFVS9f8egLrtg+3yh0Wz2TKK
eby3iFN6P8uCL/7Ba9oESnKOuvE72a60G0ihOeoCgBr7AWOlksWvrNShO9VS54nq
s6tsZvWkwTvnAgz/u575Uhaa1tNq2kJHSQb9j9aq7YEnrqv4oRgOysLddk8Ic0SR
/x3NcDD4LlhLxa0/47X8AzaO/g7X+Pt66SDzlMhGI6XsbWPw94v4aN0dJWNp3T1F
ONFnOlfr721iViGUvhwwuOtNuAr6ATqnIxb9rlgw1/SVKm4Jd4dsHq8dOI1bPV9A
jf8olaCVGai73IIDOUeCybhY+k3cdz9TNfU2j7Hv6ygahlOd00iAMy1jGP2Uycnl
/xnYA13dPWPzL49r2lg6MCgMDCBf+9g8T9EcGQpHXZ/UDLouj3Of6LlFQ9UCFVRD
Csi7TVEyiJ8Lw6dqphyT2r6axtaCByYqLdAEsGeUGWPbpsAflrA9dgSypuTZkPl4
0+Ep8t04BH5B4uGad/r6JVNZ5tDWZURkExDExme+q9m3oyDU4ujJQgv1Gy2nhxIB
dNHyxInSNIumPBUcoba2JrLYc6Feiwdh67P4Dfs2EL+XXfEXkAciPq8XMhqvD2N/
sdrj8pBlcu5NExSqBUMQqch9BhpbWBVxENKGulPUsId/jvO1syTiqfGZAmXtwWYg
r/OZyU6r7U7zlOgCf9a11YSUJtI59dl/nbxUoMDL8TO24XZP75rjcRJ2/4+vXs/v
3w0h1+AVbaYCzEbjP9I5lfHSKZpKsJbBA7+wL2BOjBSrRyvlfxifG7hNIhTXkg6c
WK29XnlmJSroG4k7EhB8ApSGCDMV5odxplezJ6jIlzaNkxy1VI7S3F65heJ68aQ4
atNwtKVD0nKCQYjIkvn+fJLdLjvMDCfhlxdH+jqCtTEH3+7Ndxrc/ZjZhDLv+bCu
AQQw8C9YC+pqj7dRPvxCmja/V6h2ha5HVMwtfeOGt/Hb8h7fKAn+qjS3mE84oNyh
5Doh4Rbq6gM4lbRNRR29NwljKda+61lDdMU2CFUH4KPDgfcOu2nocsmyO8axNL7l
15oXg1VlOYCpMAZBJ+xrv59Nytg/B9JpaK81OaTtAS1AJXHI07CVTQ0JM3rCJGGI
9/H/uZkrN9P8cCpg8F+j/Q8UanucHz2vgY6H1MZT+1X7yOlznyILGQLpdr+OMOlj
Sfh6JbQM0pXOfErKs35EMZDcuTk+QweCnSmjuT3SC2ZQUhJvIGpg6Dsg9sUzCIQw
8pqf6h+UDfwt1t5IGGS2JI1XPfFB+FKwPUWowmWAREgj+As6ID+lSTXcrn7pHV0G
e1psZXUyvmf3YghwgtKL7YzlmAl0JWJp5BQ3Gaeaa1eWPPPVVBFoXqXRyhd4AKZ8
C/9vWRUjJiOieXsBZ51s6uMZ9/VZTnOZ41ruoLrqY2iAyFLbGrFXoTXYOEfxPZvg
64m14+XICkwxsGlLPq8rBrlxBjxO1bLJDxj1WGa9L0wUmfJUxURt7pB0haB85Hjq
Sx9sre+zEfYf1lKfDneGDo3yRByTPpWoK7zYWaU/3gyWwqLnX5aBBrVNCMD21Kbv
p/zd22yfynRI/s3pe/igIuo4f/tJLSTsUu+bqQKJ+ZhIWGlbgJOwY8n1iU73eQvX
a7ZQtHsjQ15rQG+w1CIFZUnBD+Eoadh06gJzvXn48lPty3c6yTNrR+cItdTT0n85
dhkhsbfU2lRMJ74C9kbiyxWedtoAtEUrtferpz69fNqtkpl+crc/wvmvIwZ0fKeA
VXlL8kqqOmss9Zih7+yAmwznHzNwijgmxB+9vggofrI3gG1PjZwmIBmfYopPFEgc
2uXVyYmKeS3jelq9n9SqM+gDLX7pjOOZ9Gj3KfBMYvCWv6Q5F9ARFdA6/KeDFPkr
2g7Ko2Yee6PF4abbAEBNmHqMSDOHlpgwGUog6PMBkAlQp89BSMi0O9Z0FbvcD10q
NFXvuinXJZr2Fn5Y/ky7fH7H2G8pog0WCC/DsmK4pBs2hkGXCTLV4NXt3a1rRldq
/4KNqoiORKq9NSl6gCR/Rl7SObF4reMDHD5x4sq8wagqAAVlp2kfzf3gZmOKw5yj
bKXNsqoeilvcv6M8k3CQZ1kG/a9xYdO9007oCARXHLdZ81iu3pIT79EsigmUTvAQ
FdFMQ4dpBk3rpUmeCH+ZLq+ZeDRYsSnRoH/6AYkdYM++zmZ+2JeL4XhutaW1QwiH
E/e1Qd6roeoo/m/NJElRB1X/98SwLyHqMzQK6328SdOfBEtGxjLJoFTC3w9wnuw5
cMojmKTrLz8tMkA+G63RvYDbA0J27ILuhmxvOSyV2mDE7ngQdkYIu1WIJU+ndR5j
Stb5Mz3UZuRS+AhVzO1XM1Yy91qaNu2WoiNQILM/GbIzIM2BKBHkGPwQ6SYgHJay
zMPMqtbgJYSoQDN4Q5JCxSjQF//bKl5IS0zubCwIVs5PWcs09/Lk5DO9P2FbL1ZR
10PjMvRHsNm4pB1N1/NRazs64M84F+8KxcBIl4j5NiBGaSpl6AxqseYziTpG0H5p
AyCBwV89rOUgmbF2y/Rguo/4B7Rc8pdpchdnQ2Z4C2dda5L2iUNHqd+AP7m1l8yM
wNXxl5PKBHVykcPfh9QG3EQVC4GdDA26r7Mvz2ZRaAgvmIk3tEPiYy1zQcZqH3v9
tQyVHoxCWmoMS1AV308B85ems+LBl/0MMn/p30H+wr56BCMim2dFrmSaEFl+19Qy
IDI2ceeuaB+HoL4lpcrjPWuLo/ZdCKOcM3MMvz6oSipkkXBFB6RilUhd12Dk2gMQ
wpL36SK7AYywt4KtFs3MIdwcFwiHWnms/0Yc6Cvb5Y1RrAH93jJmoxawnfRA6K2W
kp/mZxh7FVVrIzb1/0oP+A1EJkZL2+8FnTKPJY1hKry8OvUChw5BLTZ06u9aGOSt
d/kZ772yJFR+AE3obQit9Cjy8W3UPW9/yuJYfVkQ2t6LolyCWCDILFP4nDQK2QxJ
RXf8HHZdCZhvo1pHQSFxPibBdwu9r5hr3KkufkhmpC1OW095s3ZC3zk7zQ9IcLCI
gQDjNOKrD1eqmxyz2lwVqxCeEdrONTWs0inime30ed+9w5vYni7J1fFAoT4fCqQm
Lu+WvPLVT/4NTSG47DIWkhRtYfCQHwy/MaoHjiwr4Opm6hqBnKwdWFaxQBdy7tZZ
s0907spQv2vUv3UKiWM7wMegCjn3o8bpeTIqWvVCzG9Jgc9EioUUgltyJww8K3WH
S4B1MVzg1b+U3pvmpQ3Nzz0qQbOkP/gilvR6JUZzg5LsniiGHaK5+LvWm2auuKpT
/lr8vnLOwSDbEG0CrPjRQTfntK/tybY19ua2/p8e6rx55Lpe9LB5AyT/NlP5vC8z
V+/d23apyRKmHOa8Acc7DPo2WuC424wv0h3FA5hImiS3h9egNyLrpBIZQR5m1nQQ
gsovnNesXEA1szO2vZZ4Ya6WTSK/h3hGr8xlIbHgluQPwfHDQJ8FBE4z/FUDN5tb
WcAOABEYBhHTSyrAUD/TnXGmEmeTDnkl78aMG181HD83VmLtcv+k1klwZNa69S1f
GgEaSMigc5Si9lsKBk7rme0I4cNe+9DsPYKaKHU3dVSLx4DerlEEqXE6sR7r7F9c
bCNSA8MiSdycWd6wr6eJMvFA0FXDgxWIgRYcZceG6/25STL3jt13Tnl5PnUUD8xH
vjtK/iSGUNgWsk9BXGbjBuutVR2rIIBU57dCiPILZCz/5GD2fvxcM0k+ffuNkagm
WxcJNfvolkcz4hsIwMCjaKKKokOsWbvwVMYaLKH9GNMZ+VmG2EXhh5rn0eREemFw
tFrhS646Ha7BJZoxG0LpSaTybvznFQPAVRa/1MFGBVDEUd4JnrWOqRrk3O8Mdwt7
V1TlXolosoL8wCtsiDwRE2UtsdAeIdW0X5RsH/chPvkOtYpBnPWoZgaeLEwMd6pv
nZKPkNR7qru1IuRP+IlYdnPW+1hivJJy9J+LFuJYUox6Bfe2Y+apU8iyL+bp0NPV
5QrePGbLLt1stOZkmMl0ML7hLCWfhXUQ51XBHn7qFV9zvUn7vemcoJ9GEH6k2UVR
4HFYxqCOEJsQv7VIKaah4omyk81qZ23AYJTUIwEMKoXNMBPKzJtRjdtOvxgDxMCG
R75tySag4Y1+hPpIpnV+JerJah8W7mQ1iHPLmbfnrJn0MjY3OYSCDuzlo43Buytv
3FZB8pXMfKHvOwZK1DB69nl/94X6GQeUXodAlrb0qXf4C6iNLTPUdyABem3hObBn
Aqv6TsTZZrIpYHVhtAcUCtW6hZoTpj786sxZRwOU/TAZlvhrsWm2jivyM5nQjW4H
EOngdsUTP6uXZ2xeJY0XUpPVK5NetZEjovBHz0NkpDRCsc/NkJpo9fR09EhndVSn
YhuhZvi2rGY/+zU8VQIdn0F7MW1nTPosIlYJGIWBvyuYLj6DmQ1gQyN1SgsU4FOc
vDqVB1/JaWxmD6Y6kMbsVwW6Su6RrqO3zH7SXqPdD0aJDtcYQnVSBsFSFt4G+uol
68bBLC6wOmE9f6V46r/gmVQPx0X+xlqlac5XlO4m29Z0igPH2+hCKmrRCsnySNtE
EiLTccnlpakmRlr3IpgN7lnTFnGYxs0FbUoT/sdNSwLuZRsMcEAN3i3DenVJMJbn
jY2au1A3LLAu244fZcZ2BgFkUMv13jda0+KgTUqCEWxt6Z/Dan9cwbRezSiqDh6k
Ug4tlbPSaVKUmzl0Ool+694Gxml8EhVrc4fk099RsEyBPQZ+I0t1GaghaEPwlbuZ
/XEo8mmWVO6hxHQXubAUuq3SOMs5xhonfs0CZzQKE7xv8YY8YwedMqaW7WyKs4yU
uCaQsanxol8lB3iNH0zGMoBjg5prYlbo33QbRJ4jNTckKRVjSsTVDM9OexOMOLVZ
99bVxeVQbFd6CAZ/QMj9s9NsxBJDoNy4+kXpau8AbBrynxZhdDcZREzi7aEKRecJ
1WZA5yWKucfThOirqOyns3lGVIe3OBqOUwsXgQPMkp9Fiupj+VmUZ/hWEwAxWG2U
f+KupFnaTZz/YwLRHVdnLdVFwBSH8XUbf/t7ZV2CeA4yy4ELZBbBf78+9Tadl9pa
5dvENGajjlYPYtPZlo//0wqdkV1sSGSIdSB1zK1RREIPBXs/YxXTj28P6u8LSKRo
udLxigVXb0D/DrLfTQ9DqWpxJKnYL+fugTE+7RGfiWqRs7RyNF7oKtf7OpVsFIQp
WwcLQVHLd/9bJACaJS+ZiAc0FRmhUHrFawBnr6a9D/i1ui+9ubdwrcEfpk58p7Bq
VuBDz/eRMlEskt2VCJlDTITPp5pJ/bu+e/l0dVMCjSn+joOFg4QIMj/Qj76Nn0mN
bQfeEuQ29Uur2F+SzAfuh3LbmxoXk73jp1tMpUK0ymrrvxPC52vF0uF4JUM+JIFI
ahZnQDLXqe3DuiacQT/2iXfYvW8lzS6nsJzc99/Zn4LXp1HFEUnen0jf7S3jZ12d
si/qNQba43N4e1sW0er4SI0O6DgeosG0sDgy2fq9VOZtK6iznaj+SLECAf3nuGxx
G8s/ChaqCYZH1x6YDVmbml0kTeUZXWg9Dv+acSZBL5CPfwer2PuTS+NM+cNUWDo8
jzq0Xucd2jXJzysdkg+Q5Gzb5ZzbSPTYsWnmqrgjY3fUyCUt26gUcryuzSum0RB7
ZAqYTOTIRiQwUeRM//N1GroT4eYFrZ1yBy4zJcl0ExA8PbFF1cE6A1bDimGnQVbV
590Ylzn5nL4msqrqoKRYHxRpirPnXVEWsza9qpVTjcJPAyqH6ROyM1VLG1Bt+IAp
NGWBm3H45X6yP9mZalq2THMClI4ocxtdbTCai9FQrtcZOktdzDvvfv3zYEbajsPX
snVC6MlQ2sEaBfgwHLjFjDFFEEyI0NtDN7hE45yBv/gIlISYsR8HZvvY6B4WQF2w
7t4EVAYR5xeO6NGPF4HgjZ9lD+xHvdC/VfkWW+wJ3+uF2SHQ1r/7tOisRJbfFuo1
OiLtyg87v26hKqUQ7UCPt7OmdBPeHBIOePXbHoggIULuF6VSqCOCjyul2HK7rAgc
OrtpPlc2pv5abxSRK7+QsiNUztFrRefYUcmMt5aVRayI5zAOvLggwrVTnwit9Xg4
ayi06ppuj0a7N8O4ABaQYlah2Uu4utdYZCh++13DxAsEQfcjvpEtWfVZVKBElzvc
LJcfpY9yci0KAdFMxmBdoiG2IkGHCD2Q/mdoGTUIn9xr1rQQC+p/4wWdexokp2rV
7NbTOEWqXGLIFbKCE8n+bdnJwtfJDuIVVFrRqpZDpPeNoCERIu3gwFX7jtDeNj6i
sCgbWZqR5bznlYChrMHMUhU5i+ong2yf2/m6DfY+LwseOS0BexDRZfyh9XGxi8iM
yhdNYWbYdjNNtEyXY5I4D+gPH7TjHh0Wo8pBbZupTpvZ+1tb5N7zQqeCxP1jbQ93
2iBB7dUVn3oSrK6yPdnUOh1jZbfPZrg8gPCxUNf64GEcBX8esLNQBLp2va6sKdOC
3789dYh8DTPZGwK0v5hCQ8kuPCE12Dt4Cyis78nYPi+HmA3n+lKwrX9ay9HRbuP7
hNd1T9e9ZVMp0fIDjMkNKrLFgFMKEbc3ayqnXgaTEe1O5P6WfYegCA54STKO8iEn
oMRL2x8j1RIOI7wbsEikY8V35g31o91vagrfl6xzkAiIQiUAIaE3CEGqN9Cton+k
1pIcwjvYj+EwG+6MI5hy/uWgUcGteAlKbm+PQNngxNb3+wkeMu5Q367bzylTWaxs
8wiwQZzJ23JqFgMnA20flwFrBedFnCoTbrRB4VMJguT74GL4GmUlE0iFvbU7wc0q
0zz7IEhvP0GugR3dIBK1iuaspK5nLVJfF9gLvVDXpb+JMwovHGCxqfGyXDp1g6va
N1rZdCv/fVh9NC9wdLluJ9qs1i+2zcD4DMmMwdeUpBieU9ZknaJx4KOavYPybARr
kgTjWqdQs9vQwtrIPW4Wj7MqnFamjDKZbQ1DaAd+HrSXMhxr5OHKy8dlghMHCQJK
bJ05ZVxwi2gCTWqFY90S1RNX/vUU99BPQF9jVCrVpDtt/eHp2IsnOJKZR5WKeS8Q
a1iLnII192gMj5Q62nvL+gzp2d6hhChM9ZSl7joEbE4NOMOh6OCcL+TmgSya4rXG
PedeY4WynnE2NG/LTcEUIlLW/6OVE8ueAisj2LbpOGCBOviXbtSucRw09VHFrI4e
f5tO/Ktwvg97G3savEId2lfxh61WI0yydp97SVE7oLk+j/iLTSEgu+TBzdeB+J5H
0xDS3nGu6AVB1m+ivD0TiYTGtJPfElX+WpyJOo/ZNNDg6ZMU5XfQnkszEhk+7TBB
7V6KUkKQrWuG/THKb+m1Y0CgGj7NOQMMgHwm2xA+JXjye5CfTa2R+2ThTHvzuD8I
iblL7Mv9Io/8NTZEvpsYc7HO/fyI3MGzjKbK/LUikfVDTcS/0DNHqyEsubDMujTE
hwZbN7Sl4MVaLkpomroJVWA58Dy0qENPG3DgYOpJ7xYDPkIaQabc0ZtYyC5U8NJy
dQYmKVds/oqWN+rEVURcK6M2ZtuNA3M3kNP0SrNzkjWxQxHtiQjxAdyLJGmYuu89
y/PUY74lhZWAmesmUCqUdl5ag2Kuf2x8qnr1Vvt6bes0J/TF90zlHhIU9Kd1d+xP
nD+ovyBnFlFIoEyiWgqN/AknYh2ghRxYwC4JFR0sXMdqmkNt6n5Dfop47X7lqrqP
Qzcb7c7PKEHAqxdmZ207wZOApzkw/y7PjK+Gts80p3OMTbTJYr9Y7Q5puPFQBAM2
E7W78mVn+M/SCtRnExS1sDA1WnYXVKUOe7RHqqkzgGmTrb94UH4tko1J7tipiQou
qMSnWzO63uC1DJ1Qq82GuCL0q3tluoRT6JmKw9WbZTVMtQOanH+sJb076Uqh/ehV
XWRFR64/TXbF41DaI41LcLt+eABrjCnPTCAsPLRLj1b7O+6AM8WqejoRJSmZENIB
EgVG1HqTNE/u6L0qq8hHVAoxUDTSPp3Vcf0yGTtrTBlr3HcukZDr/1GvDdf4R6gz
2KPPppiw3/DFWbjHCHES0pEoRZnKtTWRx/4hU5RcLqYnSFxBBpCTMCu5n9diFPFq
jYz5jU9Nwc7AFlHlIBI8x/HXt6qFwMt6rQJNghe7O1580xGph6duUex9JIXHuL6h
16ykXnRJ5BFHxpeGGzIuIm/JhXQ/VrSmf0nXvIW6bDZq2ImYGmiuagUSpVoMww1p
xaGUzjWv7x1sKOuekoO5KTwXMX4qDOfhvP4jK4XbqNrxvaSANriXX8GB13y51MFl
0oh7SSnmxBNkkxqTXGIhuBrH/md4K6kRDEWRzCAo7VXoBTpLFi5ZQd4lllbcagUO
1uI4BurOTckQlPvFLcQPtYDBiRpbACdyrTTX0C2NIda+mibnKJyObUUqpnfJ3h4c
n9CKts8ZvXYt1B1AsQQCAjGf9Q6ZTNjFxS65oFu/YbBFcmhPb90KmKVxOXkBP2uo
ip2zZZaMaBBz3nAPhq1VO/XmkeVDnqE9ZB2bNz9DfFYrvHvyIIJwfLUlTCzqw0Gu
O1Ght5SNCr19+NvGhCXOE0T9Iy+ygNw9FMfssJvLu+iKKdWp5NYvZ80wsqp022fL
1ZamgfC5EGemldWxv8+Qt1U+9OfwJNpqUqnjq6QS7aNdQujmwczTheyByX/P/1og
ORJLhWXR6XAlS0+mmD0BvpT0FrzBrvkTKqQ6wqqJ9mf8vCVHEP/UngQQJOiDjHM6
+INsl46oJ2KUym3BOkEfYBBv/mGMX0w/UXisg2zyOYBE7QxuSvrsOs2ZgEyQPQoG
MeDFjP9hsACxU2OwUSDhxZNG1C40XMCmZ772/nHZyYhoV3JWpmgizeX3AIT3aE72
GamPIxfeR1lY9G9tUq0wmrWaaIOf5KAWNQg6xvUPwVJ50gVeE/gdV63kyhh7YhUN
Cn3XAuhAvuoQBZlrT6p5yiaijRsBQyuViIDXqPnqFUvjT5Pvp6qX0Gu+kRGPtbkE
cW+kib4beuiwlpReywGwqeEkvuJNm31/qnaq7vUOYG6++C2vF9lLKTwW6vm1Upk6
37gADx4/IX/8OCk/6NNKrfdZYpOCLyQUeTwTSIvkQeBgnIRd1xh4vybHV1tNWZ1K
owcJwYmAVkZH0g+S2RhsfLFJxaWfZRdT6X5o/2hL5yL3COL9BTAIK46ZWZICfvAi
KlnuZMnZscqqaUCiEnKiPMlfobARdfpVlZD6w9fkIGN/y5iyxZohUIkVR1PbVyUh
a5KX0/JEmxRCT7Bf5MfnLm9ToNjU/YIiN02IeYeDIzJYSz0GnqaCr0ZRNX6F/5TD
mkd55GIStiMYlLWbgFO9bPQTyvIJC8LqdlK8WviCb6Dp/w0wNPIh7SN51YO7CoKi
stfZSrrrkoAJ+i6FkR4gHcG9EeWmSxNdbC0S2I43fmUejb8aGA4igQwF/aIFRxi6
bSm8I0DM/DSd8OLCR+z25Ia9vGYAnvot39bdS4IX3yWS4aBi7kXx5vVAfkWiT9N/
qCmvQgnSM/Hk6QNR4LBx9zMTzQ46CjUNwD0vA9kwNvr4toyYyTIC37bbJkGgICaV
0FFIn9u9L/1Wi76QcNjcG26O2KcHN9uKw8NlW11/X/oGRIaPnIgOI1xWVEVQL7xJ
7oQ/Hq30edQDakmkxf966S1wUBANtIcCbsgAbr/bps3WZ7b5aR92kGJGBNAtKm1j
CyFvTIGl8/2Ti14e5KG9b60gYsvCYa5FX40u+Ai2VyxPugkmcJUF8TZAfvZyY2K+
qE3XQTXlzMUfhu4GQQPZ699LrP1hwpqGqlO6Z4FaFu82Su9DeSIL4Rlv1m+hXuU6
hXDiAMKrdJ5GQExVhKg+itPy+Pe2bsQiI8PR4Ynv/Tsr4S9UlTRbj79OtTl+cgyD
aLMJq466EiOvKYeZAn+GOp8CZtv5sEXvY0nvhHF3z/hJ0LaKhoCHFmPuh3XMq9j4
+HXr84p5XoS0w/x3/Fwl7FLRj5uSZuVrRGy138jxNrdtiD8trmf+EtznblaBT805
fywEdTv3MhPI9/HScdux9xNs5hUM7Xs/VCXtFstmCD++yLWbQXatAoplZUPyJLXC
WGlioHwPqAm+Gy0ezJI9jTyaCfZYVMRJ4kfq1AUXEqDV2peHYhSjgA9PvKNqNKrz
vPcAlvLay7FCnr5cE3Tbz7Z7V2QzIm9WXrWl4W0BIDNUQUZcvFV25B/4h2rUxZZQ
LUq2E6l+h2K7D15AZTyZhzxPmdNdFc21510+uSEw6grwKv/uX7tesfmgzyl0i7M6
We/1qjIvnh53qLw8Aid+udL7ZQsPp/Bgd8eyCY9u1A7te6uSXQH5BERl6xBl5w4B
SfpuMll9j11U0hwmuyvXAZ/AYsZCvPILNG2z0eSOmsuzm039AwY3Bce95VHPW098
3fQoGDyELTkrSGs6HWTZc5jbN/8zqkmkX9s5Y/nq9NI91xs3xI3iC+CCpbhu/wLh
tm4nH0A49b9TijMSEUupbB9/sXXZQwiz65oCJ40cQOVmLtSlbdX32JGzsRLHRkp0
ssRigqDrYG9IBAppj2IFHZep8hxZoOFkYNDosMgmbD4/KvhQWDq7reZzU28LxMMD
HJKcuztnXWlFje4sXrl8J/VwZI+/6it/yGDHj7uB/dzkoPX2BXot/W/6K8EVAi+h
COZTGq1ko3t8odEKjDShLzAJDBVP1iqy+rtTshY8S8j93SulEFcfoEJn8giaTqz7
fcBXvOf4fmYAdLMcVnW5RANQPm0SJ5SlX1rKmIoZXTn0C66oMNpi9+3vAnChzNt4
G9o6Ez7TsCCEljAs/232VIeygMPnlKmYdpF+jlUxtOXbn/sKJjAmQhFwUn4KlDnS
OUh+PhyJwZvOcTO+3n3UnlLBLcSCOaSnSiBU9ZqaujAuzp7gq0hXggZt+unm+MFC
01tVb6JYetCiwI36ThsnyDmcXVgn5qjUnUjVMsvKhrtY8iz6pP69EI0APg0LqGAU
aLiBuUmq8B7rAQ4ru4hN69XoEiM9N08Wt0miLo7dQ2aXbc+hyw+P1YaUMouyzr9b
Fj2wWuLjtIGgNF9ecR0Db5vTwJ9CN+eYjeA/de18g0b+LoQLuxz61DQe1DyGz++N
zUVC68cGnGrrF1PgtQSh5FUinVjQ336EfvOJmqZpcsevItafSxXjiVXATn/WjSz8
E7wzLeJNwg0Z0t4ODGXV81yqIHb4/CxfAiiPYCzsHOjiLI1Qfv3t2FJtrIQFNRkZ
1zUV3t8+xJ+07DNKmLzYCUmxhzNT6gpNC7r53VfL/r57R/MSPxGBUdjKg4Br8leR
3bnkNuNNTYqukrNIAIv4DYp/pu3R2btMbHnfPBQQt2CEn27fzvq/JaLNvH+orrch
9G8+wPDZH/d62lkkEWnEaulgTILej8A4YPvwl9ROqsGLuCLLbK5TM1vyJB5g/5lr
SXnSTa3FNvnd6BfSwjXJAKGdMj5JV/eHVdDDQ8QqKbBOx4eBzYIvT1wFw/7kXCtO
rQiLo9uqt3LwmK1S7XRuzwH9Lka63glTcfOOEvOCg2xTQtiwTtLZi4x0Z5gDp/gz
AeHTYhb5KGZxNhWpIT1oAfMADSL5MnPcV8zpXwifUC4GX1CzUuiKBALKzi57ail2
VQ0aLFPYvVIz61OBdRmf23b4+hJsYH8BhrbkKEcUrxiuMYQmVJRT+YO/Pdxe66Ly
3KXcAPGqovjhmuPAjVWpx3leb4ofAGckQAxzwr/UYR7DfM63E31U/0ksxaETX5a9
q/nb1OzhDW0hb8QyXC7JSf++kUU0MK5iKrCeeHfUsGIsXdNmGrlHt9stP0tI/aJW
VaflTC7IEgHrgwzgxkwcJ/Dx8bGmUXzQf3frPK+49AjLvBepfvqFkoFXJAoXl5oo
osxSDUEW+oKqyAhTTAnwVwvei634mI/OfXAi6Yb8UkG6WWfeAF4OIqn/ffcxmnCh
VqRPaqEHoJ4f5GQHd8W2u0w9vP8ERb94cUbvYTgO9szlbuKmC4pHF00ayBDwdl9D
9DlQgbT21qP5UeFgOpxecVEZm9Hh4i1I8zVeWCZuhjtkFtgRJBXq28B35eV4RRNJ
UdsumReZsHAFeOb/HttfnQ/mPAQdLDEeOdUGAXKeO5FKfyR4SVIlWnkYSlsHowxH
BrX9n9U8iOw6pNajCP1i6qNIuUNaGQklL8QMyjTRKby/Kp3D2ijWf5MJMClxVM5N
6J6c//5pX2HeDrHFrAMboivpvmwwQ9/mbJQjOYrUkAmd6SzsGQThmbK2akPVa+ze
8RIW6YqvLtaVzu/NiFzhgBBGpBWH5lZObFKPhKO2J7w4CinToS6f/Mwc3RmDZy4b
2gJzzXd6GMrox2fFsPSmf/gnGqSTfpkJo9bolMY82uSoi72nHY256DrbB60ub9xK
Dc/DFK+cPJSNQUj84DWZknNgDLLVU2ueT+iFLZ7+1BBZzDdhy13FqORTT15KdxT8
caJsZKgEQ6fYCofbdNoRIg1TJ2y1VnQQkuEpHoPnTfyodIUYK6oJYfKLCpqt5PP6
SeKGC9jBHuUy/8OnBBcDObx8k4ilhLVY6lpiL5JhKieN6nwyJwq93AMLVFQ8PMdy
vsXq9NT7tKW4QqBezKbJqtmzl7VPAbQzIYGGnfRAFwsyqdZ/hZ0qw/TXCyOvaCQW
n4CeS+VkBVZLUMY871YjbIfXO0l0aHNowVzVFlVrQX/oJj2M1alIRv5J/eBdCNxE
8UKERVT0yP5WZTVQ3ecRilAK3OkcHfWWGRTbFV0tggTZhBRbdyKQvrXpN3voxGxy
z2kU2zqPl+tmWN0M619Hw4v/ixHnzM/hDcL1NEHZfEXKwATZ0vEkD0Va4n7JA3nS
QN/ceoQHUhL2Ggi+istFs8UBlHNLiP3x2hDfFgfNkgNhUYRRVC7KIX8NcfHm6hqD
9XyjpZBj3msx0mwodVGWAe8kk0ldyf/WVfD6XYTpSZ4Bzclaa7ppLssuHFkMIscK
L8Fz4AgZKeP6WIDY5DK6PhrleyMVzqlpz1KRKYFFl/KKmorod8sdAYORVOrvBpab
4PUk818NE7tUKJ13MH3jx1noyBqn0F86bVEM6/mZCmZ5x1wmfY5RTrzEikvr/S7a
tSznmaFcOmZU94p3NjjmGGEC1xYXJUOSoyYRpar8oYbbHKINcEzUxOsJtQ+sVAiS
bcMbNJp2cNNMix20WLOlQ3AUr6lUhaI4GAqA9q7csPINbCk+/5ug8xUQVPUBXaCc
E2QWBscuWBtkiOKJCHZhcmMu8ijzpO70ssUkBTVNF7q4TnnysClEGx8Cnr0dYDNw
98dCNFjBQbr5XcQq71h1393tRp6piEkPWK2sJ2LHh5qLQQk60rtU2pvTgipiyhFR
XRaBIdWhCLVQimB+g2BgYFig6K1FfVI/Rvp9k0bP5tRR3dYncKyFXO6lDGs0NcSA
vn3zTehHGfZJisix326/pzdA58DLI3MZUpw5LgliqJ8SolS1OmJ3GxJraqoRm/pq
JLe9oQDFlxfbPYuB4V5tV1ZCe9KwF4tB9ctr+tQekMAQkU8BxymVAXUXVor0jfws
urcoGKlYrFiySOlMLgIs9uubUAO7qomMGHodmzfXa5dpxSj+RekVRwW+5/1VsC13
Z6NE5HQb0MDkca5VMXfiKOMnYzAEbmuKVfMKrlMPsU+HkjEcp4lvHR3aEV/d0IR0
wOAuUXWoevnIZscur3PkvLcmzOV4FwuWBkvNKbSuFD719JlXJDUpiIQJcxXED5I0
Oqpl8QKo3cqTml22b4sdn9AZIFKmwJDX1CjU6uxjiCtSAf2MH6f7k4enRJadapw4
oYstIj2ImqoZ98M3j09O+J1yPbhT1LKcWYNw2jrGO6t7JbHCytszSBR6JEEEr2bC
M9/TrhR4LPwI3ZI41Ax5Gqi5GkajdrpKKXnbyIfnATtc5wBHXB434AA6R7LMo3lx
UJ23YCrzTIdZWQF72s20Mcd8VE72T35gQzJZsl3hOwPm4irymavQdYmBmtX5G1zN
v2M2Tl1MWQ8jy6Id637uXxJXMOo9VDYaAp07CbGP/ImcL1/58+CmhvK4C1enaZmu
IJPnexpHtNsIL7czTpwEiAHJ58ZJOD7KelNz9pbjJHl7PAwPHVdqdcWtUBqgirQn
jtoGhR27xFs0KcxyrG7114YDn53UrMTInO2lO6d54lHEVF66g1lX+tlPSAF2hVS1
+ioka/ge1sANojS3T61pQ191upxXQyV3Ot3+AgfuAmwvrdjQ6FczPLIp0Ytj3nsX
FSeIasNDSVs6K7HDYK+vw3P5qBOdygL3z3+sXrCgbmSSUjS+lEaI3Cm3G4QSPcqm
S1RjiWDR5GoGfMIktO5udC/7saK7jRFO5/lioYELVZBcthdQJgcDByXW4CaVshiQ
QSctdB7jHP7pzHX6hVGh5bjP1+V7cJTlzxaME6U7qVt5Ssg24higqXC5hezdbzd+
yuEvUPOR8W8+121JLKQ8svUQwizimE1wVlpJVPlYKzEYGGB5ShmUFKUui8TMtRmg
uZIXlsw1G0OHt3wkjG/FnPTbferSHsu3nQZNg1zLjrMm5xAk+LywSx4wWM6nN2wz
b6hLuEtD7CPSb0ANwCEkbgfL/RX9eWw5mJno1y5EphlRXu0FrECtkL8u3W2tUMy/
1y5C5Nj3qW498dpUzD3YgADTeNvYMaUb6hb/nuay72Lv8T+BoqvQA3wa8mGg818a
uibND7TpNCDYE/NnF6VQ1q3aZlX80aXNLVm14VzpZCuSbBwffEq9Anrs0RtN4v5N
cKJC0VKwp10ieggPvAa0npaek7Guo6ujVFxEznDHI7BHviBihTAY365Eoqf6HszU
MMg9JNdlLIrlC0I6CS8Imw8fF2F/rM+wNpgGM/+QMs+cFb/mkSC0AEEaipzQDdIX
9k0XNvyW4aTvp9ldXvMUv9mQD5GmX15EhjTrZNHKX2J9r+f+e+VsCOBsIG3am6hw
CJKQHrVcDw2TKxWIaTOe+Ex4IFg57pHH8V85+ZeBtxjoAlVAIWG0fF+6AIUVEyRJ
9wAmZuPW9FxacV8Y/CgmH/tgX6n+RfRuhJB3OKStXfDOqzFVDJXwCEIpJHrvMFtn
dfLS5oUs5UFs/ipTLYDEBP031BNEOrOYFMThOdmutAGFjbOk2dPa/kEHkFn8U+Pp
1UakQK2Ick/39iANhJ3Uz8eWK8Q0c9toR3b1XvK9Cq0CSp7T7a4yrjRLq8PzzMGG
1Asq07XP5kxoo6J2TyzDdvW2taQEPc6rgo8CF0bL3UuE3zQP4+QEKcaMi3Ide2q6
nwqsxFku/qHutBWY89fG5lFI0H0d14L5YqDL+ioFJINq9SWJh1XieNPxW3zMp12w
Etg7YHFqmbTqfpoYPwOMl6xWDxm94TGYST8pI7yq0P3Wp4MuN8U1eHr6h6sXyMkn
Kle3mEavXRy7OdlKj4A8KPAbmttGTPzxJGrgrWDby2ExLvpyjNO1mgYio2vM0RRC
tGwUeaYa/c8AhSm4vX9l8Sjy4Ae/WI+I6+KUtH7jdDiSb5P7UgjvP8Fr7s9I/Vj/
aVOLKyeQISx+jFsQ3o1tjtt/pWZygxK7IvPLWUZ+xs0j4pxMRNCTIm7Og0honKne
siLvA/63kyyAUVGDFg3nVMoD5N+AcVjLyTEvNf3YeR4W+Jkcq3kyGgGjcJhm2s8r
2gVko+ISDn/NjOo0UXnBM8UIIdFsc859cFWcyWWOszeipQXJIfb1IBXTCK1AnPa2
HZbgiW/Vd6PQGN18bXXA1l0uFNNfhhokhMVy6kuNDhPKrjH9fMv9VgBzQWPCqvIx
1aV1X/pIGVa+7Mj0fBS+yMmbCp8g1g9Xs4Bc3ZNHmJZcGYV4R+JdECjQP30toY5U
IHAMpdPUPElGw2ZjVWaFG1mOHUvX17a1JKrM72AjZB35Z4oSRi/LNXksY27mGxfc
Au9RbQ8U3XWzlh6JZWcjUafoTWgiEwwJk+xPEKcC9ThshfETpFtYBFyRQqWaOCgw
vwNVdSPE0Jyqm5gD5YIsDS6qLjdgIc1ZDcR1W+iZmrv/StPWq7o+dHlW+8ZEruIl
8zhWwyIpndi4dfqsT1UAgVaL4p89LW1sWCCO2PWUogZ58yCZ5aippsIEQA0ehOvM
v0Id5LGX2RxPJ1wv5MB1B4WYyI0D2jWiQsZbksiL+DYVSc6NemVKDGNP8w5TjtQi
nASwgKHzsRqXZ9Sa5eID3OWI2/LhzYh9ZRpaWsq33meLzVF7pE8p79fCs4a26+KD
bUhu/0RVtLM/wvORhOEmxxkZbXQb+dppUXT6sGkkb+Z/u2jQZNmlhl6uZNW1BMOW
NFU3bNFhFhfd4Y8iZqIMmJZtq+9gAGIOqaeIsP/Cy9SgTGvP/4v4QsNODAtXLZKE
U7mSm6i8DoZDmkSuOOS7J11n2NtZgL1iKbh44tLwCAL2BXjjU/fAuFoBsac3hJdA
zqS8JhD4CToIZLHDixVW1axsC1pxXF3fQPhADLmCTE6zBNjRdUm+WgWrevR0RScb
RQpo+vUqCevL6vXzbmtYuyPaxqokBrFrS8LgUIfn+YXka5WOPUvm7BOTw8PABK0i
amZXOecVk/6xHn+sF9Jx46Bjozt1Rq07HBL9k/S8kwsc0eCD6Z0Kh/KmNZgh+1Zi
MjO72vFPTarsHDT/n01t89fGQjZNwTDGFepnYQS7V5AzVCHGGHEvP/uC/iyn5JJ3
fqSOw3bj2gpN/kA3fznS7vd+lEaWmahDiTSV/QtPCT0Bdg68bIhfA5VDAq8RptLo
xFGMe/lh76RB3aKAfN8kXcI4p7dW0HxDPLNn/4zjEB6xfqJVry8GW8E/OpVkRaEi
GrZ4Ecox+WQOscv7q//3lOJ70TXfnXpBs5wexgxI+6OIiWyibSDKhvni1ks5+gel
6btDSUnUlEmmfcceKfjW7NCskhRekjn2JWiB+eFMUnNakj7ke3oeXld/g8htXipz
pNruPz4vp6fuXHs3ymvZWRHEd2Ya/gcHF0lW55gW3vttb5Hnh5n7kL7b71H4nf2E
RMIPvbf0QGqNTK/vGu8yRo/Jp07RX2xmB9qsfpFvVtcCt4ZwUu0WdIjQXdYb25vX
z+3vhXhUbi+GjMOvm3BOc7stLhE05heCMuahDtM8yDgAMxt/rNz3dlsFGd3jKpp8
whc1TccUq6TdNcsx1jINKEhQQPGQEYDxmYMqmz01UJGueNzu1mgW/Va+SEhZ6f4Y
pesM1jz5QUTjpxz+khOmbjO4C5xWg5DAo6kvYSphy79Fyd+aYVuDX2Aburs0AU0V
aU8cZwp8GyeW6yG8KnuaVed5svrHMJ/JSrsXFjcvD165Olq9m2YR81eIB6cFYFxf
6CVvqYi3bF+InMe4W3xGuOeSTVARNtWCNGKdR4yEJgB9pprPSVmzFDipuCeJLOgo
bY8JTiJ3PVX2NtKivODDF6iwpwnGdR91PgMb3V8uX0Z6q8X6IEbiMI0aWc7hFrcs
7xZd4lZiVO+ctAa/DPxu3GCgnat1AJqahPFOXk5q1HMlTz5KIaPPQqWzPKtTfnFB
qxtaetqJj8PQww6CsnyjlK59JPsxb7RQp/j1MkJ/QQpcddwYIZI1uwymb5bp6+Ke
ofw7XSI7eeVr0rQ6fYr9weX1adRDVNbAUOtf5G4T19RZYBc8HY/I13/yZnoEZdD/
4vgdxTeJQyysT3Ss66WzALiNL/5HS6hLPvR15XASnbC4X9eyUTx4TvLBvTXWd7UU
R9Xtqp0PITQ+UPQQI4qkwdmeoRy3s2wlXS9justS0g805V71+1y0v0AtQd6F7Nph
jRSxZK/fFlGkKo6fg/Dt99Egt4GHEB0X4HoOIkH1pp/BgfcnAKz/McIbQruC/4f9
zwCzqtyu6VmWMREhujMDjnpH8qW0uRemRRtxmvFDYFcwt+IUe4cBD2EvgDt/tW6h
x942sc+5semaFoB6e6oHwS7HbhviqWPtTyJWCcR2rJBhOq5QiWs6Sb7PF0MrgmUI
XbnK1h/4MFnTC/usBRE0y2QWgx6VuETeQrhIKUWEP9cIqG/5DBPIumc4AhefbZe8
7qJhx+TuqY6CVRKN88TlIbG8Ul7pH07ic/ns9p6pzYGGb0NnitdAH1OOIc+uJJ5y
e8E0+RxdXV1UkVQ9BNNSl/MFvMoTg91yoeYxJgF5lawCbHpZj677uMppBtbyZBVU
nWVwp8JUuwf22lDvPTVQhwaQwb8W/f+MOaLHAiuVZxFWP5kJJQtatZ5RkCY9EjeX
C7swkB7BxCSLSue0QlsArP8Vr7r4wWNQfbV19y1KVFTODw9Y0Gyq4jff33lyT1v9
zV5WEa9d7ckLn5jiByN6cZ/3RtN/viE5rNpdGd8O4iSvs+qHHT3pPgCRL3LPJRmV
iN6Zi+HsfUITqcrJvjv7PPNj+rgSKh2k8UHGIecmk46y+vPLDobCcF91PbBiZWFH
+7aaztti0ooB7hMbVefPA7GkOjmXAXeqbRqszaIqoY//W1mRQT28MTFCHiz+ilwY
PfpmWoO54cikEz0CdWD+a1dnauwYc+dZCgy2tmpRKtL+2NmW8mDIBv/pd6NMSXQU
Ul+c4yJiv8Xr9l0XTtB3xs53g6JgkYByGbIipvbxXNEm4rU+Bh9KLoutdfFlqD0j
F2NvX5ejCOls0pJKTfR8AKiljcQH9CZoMQpuVw5ZlGUNsrVr63noC1xGHNo7YciP
QIoldBuL1S2gFt6o83J72E9N6xjhhW0Vehxa7gIM2QHvhCww5FSMwGZ42YupVGLF
zgsLNiXUvh/JLbPUwmYHSFfzp8dZKpBIxIdU3/1QiZSJk7gf1LLXxyLCTWbWU+9k
3xbSJyQTQ0rkpzkxMZM2HB8SLNkBZB3ZYx6s5DsnFY4Q0qaNixDGzOdSOSL3ca2s
DmCwKo7FZrCu54J7sbmJWPI7xNKxhzg+i8ps/1eGJ8DrIgYB2qID1tsXNieMg4Bi
nTLQ/nwrb90Szw7x7X+n4A+9kItu/z0IIKcQIGqwH6lKX7u1Rsyjm4O1bgb/8VnO
Ut7IUtZutcv1hY2MENUgXAXuqK3OPglxtzaP+633HhBNRuGwwvIxsP36C0RghgTt
rI5fVTnEjOB214rcyyEl/TqoJFmI29tki0cSVeFZ1iQhoUphcZD2bmo+g2CfEAMf
qc+fcOd/JHYYzTg9CXrPXDkiZ20+2JK6CcclXN2TYG4k4ZtDZkKgnDyZqd9D8RwM
W5Cx6zdZcps/pomZjepTtz5fYYupOYvdosLV7uon78rRjEFlCURhVqLY3dodJYF0
ZndmWAjfwWtPBB0BO0f/voexAkZtpZ3ukq3R01wtP/NGixJOuF6KbjNqHg9Ttt+n
6uj+AflFuSeqGSQXmIGwcP5CgWAgwkz0BlhfoZJ8rR5KFp53Uf4Q/hNPxaAwh+J7
H1WVIJYhu/14E58l+Jr1jk9ucHLU1qXILUP0TjeGZr2/8k6W6ihs93N0C4D6lPK4
zw1eYs+Yyv6qBtOAwHGBHoFexvabwqemhKcH7dGbmZQlTsv2miEgVSP8iZoTWPdt
sQTUid1ueL6ZX3mY164E/LW4mP4cO8hsxsRXD8DIBv13Ss+XcWoOerCNmLpiVX8j
0Z29ULCwTdC88E3rTnv0UL4f4rinM2Jt/K7kApOUryYocsA+hELD6ihuFf4fs8QX
n6lGZE9c9WlVcSY7+tt/tPAFHx/4kXEABBEQDxOedAroso2Bm1vTZcqxKcw83eht
ZE7EJVRQ+8pUCs8zKG9mNCJeRRrDXlZzNSRwJBosOOTCHq49Efd6lKdomC8v7vzm
nEuWQ2B5D6b4FMbyRNV3RIvuXem5oka1vKJCiCEipJk8jRNwQQwNW1cY+J9OxtGd
AlGsoir4LO3S/XXKC6Efqn+ZKec+ceaGVpYPk7czx1c4UXr0z8619ZdSIDRCYpxM
DrbNZiC6drn566Z8/L6P78ZV+tJgzYqu1ndJWixW4+kOZ8gW0DReTvJ4n1CUQVjT
leZxNxPWKAOj3cs0OLAvh/jtjwllpAg+DSAhgcvqFoJzttGLNnUE4x0VtK0X4kUt
XhqupDX2pYeU0UECkXsEBdBF5luCJA9oeQFYbLwJTg129ihfUssCbVCycbk6P9uR
3Zh33iuD1ci3ynbuV8k/M6sTxhKmhpGLd+K0ICXI7BReeeFdEtHljSk7RYaY0v4b
FsPfUgJkhOI8l89ipiONL7WgSGb6Wqlci/So5VYTC3skEscxHPEaMFhl6URQRObx
+Mwbc+nCAyHnoi4EGnjZNy7rVALhHE3ZmwqxjAehEoC+lqCXbNMGS6Jz/UHITHm+
NU0tVjzWbJXdN2ewwbFjpwQb5eC7IqHJJB0W9pYp4UvSzXGaqI0rR3L7tbsAy83Q
bZ1KF/WJoP9tG3hs6RXogOFQcj11TAJyBsDWk8+sCllCOFxgryv4bPi/nMxC6Jz/
CNNYOpscSpPO7Z/IhT7tzmKveJ2aKwpLUOkHFpETLhipDg9/gedO93ecjAkfP0Ya
eW2m6oVZoh01EJCDG83bhDOZcMG2MHtxG3arK7rUWQKOXhWJW3Gi3GQS5VpGvCTq
nKHJqowVCfkaFjqAYgwpKK4o6Z3ijUo/UrcdJWFLqSx6uZb/+1LWJGF+FgGYfyug
uA2MQAFO66u4sUbOvrz7ZuXlKfy9P87WbXuYIs8CIkwODruoWte6QImyxeBJ0jnF
8FZvB+TbhomA7EGwDN/rBd5eu3fTesrDb9betljGNKKr6/toU7hjUoqobEDLtBJi
Yitkf0AqAzsqoNxXwP15x8mH5pbr+5GqNpd51f4yVN8oBma+qdO08sOVm+0QO7Ox
A2y2T/nJHSlt5mei30tmkwjceR4v39HxI2XSt5joU0BEwUWh5i3D2PkU3/bkPuw4
r4nNlqHBPR4pUQB/2sQrZXRA9hA/jEv4LdBaT7s+VL5mBJwnVhnqQW57ZqOrc2yj
QbDT9cJ4HmIQH3VWNZwvkf9EcDktzaUJ1d07vcN2RMP3ctqxpD7qXECusA242iEt
ISQP1TQatENPrOQv0DWoHFSGWonfuBh6QhdUU5g0Ys9nFSIbF8d8lMYT5alB3dQV
POyf2OsNnfv3sMh8fDFbh+UbMA0OGA0XJ0o/4QhJF4eEQ+tB5PXuXe2lVl2JrklN
f5NfpJc+sz/5f38A+73P5ZhLx/ZGCzo1bRTb2bhJLaqG48V5bPrakc4HQDM8glIC
jALjkV78vUa4VLts4CriI1LCxJrmmTFfAd3aZIOCIREW1zm9mnA0odfWE8NjE1dW
z6Lpnve74llC1j7HuWlCUDCbCK659PuC4ktMLN24IckUy0exLi/LhuPTzhkixHQ/
1/RZYJGnF7QWduWGN49IdVx95LgYMHCjU1P8ZfsEoxbKtabGu7zgcObxUJKBEF1H
6Gv1ERtjZxrAf2svDOlAoLxSuOCMMOAZi7pAF9Mx2kuPAvDh9tnS7bKWVy/MNZL6
YTx8i0kO3m0LxqB5ikRTH2na3I7u0bZwrcezx3meQQXBjnjkqTHGArJhdrqLcfrX
tSimYeoSIaXl1lN0wnqgGJEYDmSwpxvGy7G3wZ7k/+52jguZZdD0zUWNaRvmCq8O
iUZajeFtirCX+UWC8XcCUVS0rgf5Hcb/z4XkPCyqbJx0CpDsC3mSfBud/AZ54jW0
46eBlPFjGHC+tF5ndeceldwJNMrIPJjBRmNHq1CUzRhrbFsSv0ODsTo7/AHZIzsr
TALt9T4PBT6xKeEfgjPRWBTGu+i5k9fz10+NvTWcATvDWPevtdh5N03In5n+wsxr
Xnz1QsrH8XFxCA+YyU+Sun3xvbRVNbQeD2l2l5Gc3axJ8QZPep2rUwJCJggs34Cu
8AlKyp/2mHSS9rh4D08prP+8njgD3NGTRjiuc+lKZNpa+gJvELKyYf70fWdjwOab
zSfYJVJIOiRwl8aJi0uUtnRmwrIwd+AmcpZW+U0KzuKSWsay3lQmPNnq/seHn5Cj
BpYe4wHcuMMTD/cRExd5+VgyyGUm6tw+P4unTzcNLsICXUzzYSUCxr3Y6KYwukMI
wd7OC7j0z3GNG7zbCNwoW/7GzTbgu316y4P8KdplnsrZYUOL6wdvpE6ATKIqiy4+
wV1TxF7i5Be4MtPpVQOgC/fIfnu3MSqpMB9HjE/N0m1msaFS98vMMBWtwPoEQZq7
d15eabpTaxjo6FeIBIYqsO21ui3nlDP5y1c+KyCXWdZFK09OVxgCu4c0tFENEDfW
Xie+CfzqAGIqWR/5h2Umac98A/eXvKTKj40qkDdbazQmVi6Ygn4S3xEs4cNhLkrN
UobM+rhTRnRmaygKlutju/CDvfEtnEJKSZucFn26qvUgomDM4HeyOK8r071jiqfH
SfBPSL8VTwTpYX6J6NnGre9yBO4+oo8MkN5wmkZH9SqXgyrehz6h2hs9EmYj8dBW
CgJWTYokW+ye2U+dEZMGxjt9/ISDt4kBMF0sUDMLkSo+OkMQvqV2mVwhDgWsiBBj
XlUWB/QU6CecuNWbaK9do5zQCkIU++M/vfELm3QgdTEXDo9R4HbeRjcIGya/69uT
PsHvyfrKzIADGzKQoxFmfkPSDv7jtCl97ESCuQulTOqMSCQy4+c7Z8UW5WvOyPWJ
aRvqrMEWfGz2tuNZD5ANCQtU2qiumFn5AThe6kaK5HXB07z+efGvqA2YSRd0IGC/
crrH+5Q7K1KZcqGNipdH9UOY/KkBznbvoSkQSX+G5rVlzfeLFYbkOCfIw1I4QfKi
s7l/VUYLhl4pEXu1T+K9heJt7v+aiQ4bqxX42YLLulpCUOoD98pv8kjr3hgTGvIm
I1sdnrltdCt8r2PejNAiK4JDkAPucryjcy9dBPU7pHMDLd+jbpmf9i2zq7IDY9oP
KuzLmWZnZhvbw8se/rxzFvQyCoY6aBv9WfxfelA4zQHPWmjVc9iIIGAbLjtATDnf
ZRXlxqu//DMh0eStfovS8d0qPszrG3/XGVsYedyVaC6g1Z6a3Hvx5dgLWz8TiNNU
2/IuKHtJwjAR5VqZEXb2I6OIo/4WIQEpcmCRYvPOaxkKN48N0QU/him9qny5fMJ/
Lyr0zE1zwo1i7xqlV6JdihhiXxjsfO6GdtpL8FETDXewZH+hfRsiCrDwheGx0ftz
kV+vmSgITO6pUGj0o7QOhqlwDV2BzjQvu4z+XXnw5V+M/qZQev7TUV7lrAxeDaOT
Z7DDRvP5F5Ay2KwJL7mWHu+Nultwo9uKTwz2Tx070iHxVVssLsVBIXqkz3t88x4w
ZEWTAgAP6atPzY9Mo5bpTZtrmchfetk3VlbkH6uxLcH0MOXw6Fnf53X6YePd2TeU
n+X71W6I38ROMFAcu4CcFHiDYPNCUvrKNMvFPgd1gp+uDhS5KzwSvdjUAj2+riut
0FdqI0yiELebxxF6oqRcl+X2n1YACaSJOz2l9GeUF8RSBzSLkWbo3k18MlerCHv3
GkpwBwBt5V4G7mYicvaGrbjU9FnRDK/kW2fvOSv3ssfHxA+AGddYF62JFsd8bhnx
H5t77fSs51YFZ6nlE3klSVeNeSiMOKQxQdcAqhew4/L6h0UGdnDgKhy3dVLr/Qv2
7+sZlfBup08tJvW3VsmMUOzp3kF0Hjn6YUR1QfnhyUfdtfGN8Lc9cHPLIZCf5AAS
1KxYu/pMwDYnU8aE4juWP2Z0e0HTz+1hYGTjh4lVRuS1aZ8aThovFy8KvF8da9lR
je/gvJsBR8b4CKaOP6qHwUMirLcDBbs2zIRT7MHT9SXJ9XZHwDNwPWIFdXHIXbmk
jbgwX1WC8gdsvaRsxaO/TCEUOR647k1sFHkZJq3aFINPi56O9buyaBa+HaxaFuYV
GyY8XsO9mADnNNlmuQRoncy/NjHQNwXL89kNXaIR3Iqa8sMJMGoZsiwJ0N+wCGbz
gs58T1Nup6nOJALlsaiR75EdAdKyM5Z76ZPiLY/G43+Z97xzZY/yyWsdemPyye6i
2AUWXKw4tNpfCeguFZ5A2lo9/CKuPA6n+flG9q4U5SY9+hWmLGqtbNCB9lmAY7Qm
sB+wXROxnz/L3mEJmSxH9pSXcraXQ64aUWb4l52qftR3etqOatc5QxwpyscrNjfN
J3ISJNw35IDSFlYF8ZKjNAaZRciRPOQzwoByqWftwilfVZ/W3KxdWUJ4tK94H0h0
R5m/GTyD3myTowjF3ZwdbIeiWpW8m8p0KfleqFwN277WSyVy4jUMztXbuxIlTsEg
Y2jLvLRy1ZJzat9+CydJ3+H3dkGW8hiji5tUrtWkZr4TaaM6QK4BT6OCKwcPalln
IdT9HsrNC6qlEz4FwJbW+jqcqzFYtG1KI3VoEd5s7+34PEzwLcxt75k7yiswZoW6
PFMGzXf1NaT33rTyzgaZ6k8xn2HWLP26EqcXap/TFw0myxLZwcxsYTKPwCEyIaND
xCVCetCyCJGGy3oD1ZxO6AhvHtmuGckaeXsUKQ1IigYdObtr3XLDPRgKY+vPawce
cs+SL4qlPWS2+nzFWl8pT3UwE1YfPwlLFiVIGS5LYRDwZH1J5A24cMVmte+aLWXH
EK9xVpHQysbKunE8Rq/tOyqUbiFqSCnYqbUJw8tVmXpc1ZJXtSVafeO/BtaJL3WO
CXGVIhA5X2jt/U7kzZxLwiOZ4/OOv1kapOCVoRfvQsTG0TyuHRVjJW7t8I1GuRO+
/86Rll6HFJ5NrzYelieSXPib7/KQl6cZ1ldtDvjbWkqE7xTOqOUdOfjeGat7kzNT
gWvExDTFtjKyAgrWOXzvoyVzN0kUbLAFPb9jn0vP6qPAG5NFPM10jL/DJFlcAIY1
izBl7skmpWhmsu0rAUoJLGJ3tQGLnp1Pic6dTS1mDds4ueM8udqZOvuS5W40Jw29
nNC26NnPiPE1NjDfy3Hglj82KX7HmKN+fbIDF4J+iiTKYHeUYJG55D/RMOTO/Syi
nMcpb0o7o1eFTUHuQu/q25ReaaYcZhjDhkqI027Ox1ez2VwE36/RxumyhPTidTn7
Ki/2e+QUb0cvYNq/Ujr8tjb7lSydatdU4tEBd0zcMWKsVgXFpAhFNf0KIXI02Tq8
vsyUU5OXqlnKJyLsRRUeloqheRQa5MXueXjg2oMSNlIUOJr19Nt7wFvGi1L5ba1G
nPXFXsGjkKlRYfbGP+l3+X5KzvppdrX2pITvh9RtfywMm82UbmFsLV9l+yICaNXP
JNnj4VrsPEiiJ/Iqzi1VpYk3OzFwtpI20gJ1wTvX7S+k2/Uf79Amf2TqLoenf32D
X3LeqxnNB57ZvQUHLcbF8Vbab0kHm3BC+XFesxnZYHW6i1saghVWoWn48mq+DlXp
vBBEFpJ7kjgRl4Uo43Wd4w4OiaD0ls3Mu6bFIoNOe7lTkB3hLEB4Tq8OIctgTiHM
REU3EQ51DHdeIVhmTnOXVExtJnHih49Q/1YX+B6KAmP2n9azZAsxUdEUSi0gUAMt
svhGiydIiMjq1Cg1/2SXpGnQEAM063NjFWhrh6aWZlmdSReBEO6CFGjO/qmDpgkb
G9WkIQj12QoR2byG1+aSYwjgkJyi8Q+42Gjk3LJW7rZbX74rf4LsOiKAgGpSYaFN
YZaBKlJgGlRK51oIMWYU3i6frTEc/3TTtgfGS0j5N5ggAw9L4tQ+fPJMGVQfx9Oe
maLdOQx3bQrFoTyAOnikZ540UTV1tZO/bPzlp8Hqs9fv0sWBaAeQhrYvtHqBPjdt
GjeueUiKubKKcv4bKeuFYbLj/PxxJvCHtP1bfJF8kXAsG3LYHQThhYJ711fN+0YM
Ei5GLpRmyotEnPrSDQh0CD+6IVNk1hAjiquPF6ny3Pxc4bnF331jtaBaRyIfi8Lc
526wuo/DfVFtKIVoXpXl5gxsJo1/aXmEnv/p9Txl4uIMjqWnXFA9uoWy+7JlopMd
VPvkeRmviSCNX9yZH6j0u0pYcczX8wwpNv4DvnJu4SX2gm6Wdi6TnOSHZif0lSA8
czHHzTxkMRCEwyxL0QdFx5OZI+kyPEnay64sZD4qbX1PmSjS/BM74o/RnfjY+L8P
8vySYRl8zkDsTb+IjPKlp0lLfUUW0QN+K47k3WSvMElaZ3kNFeQGZb8edR1DQA86
smldnvx/O4uEOTt5Rx0Nnsya+WL3u4aEGY3jhJ2KuzjJZJWvpjw1aZWnTHZ67wBI
SYAUo8sYiUA7CX6UsHUlwoE+dH10xsVynUCjJpW2YD5M0kUBz9umQnvvzpBd60UJ
Mshtu0sB30VvVDslObFEROculhyNMOQGdSujEjRn+A5hxRQzBY+VYZCWc08O6D+h
KxH5vqLIg8QEfYwqfwfYdUeqyy6Py7DSftp8oGo8mpwh3HPXTqklxmxWpxhWk8yd
d2uBUIEl5690A6NTQ4pmgvVKcP9Xvc3t52uJ6kTd/i+E1lYiu0BvFxwh9byAXyFH
EjVoxgARjHnctggY+zEk3G13WvBpofCX9b5XWYn+p/KO4cDyxwiYTK5Lj7Ytk7Yc
l6uLIVk+x12NYdDuuM0UFOlVI53P6u7OAhRh/Asf0axS5ol+eX6aCiBsH6fF1IHK
/Cn+1jIQoEF3kO1HFnXl3rD5tuCXXX0gdl4pCvaa47xTYb9Ocq/bYXgKfLMX2I58
4FEtObn+1FZsFUDnzonj9GI22qiRZluWWiH/yqyD1L6gXH39tu3uCgn7BwsIcebl
lJqyJbcZSVlQQNWfw6+8QKIGvW4InRPx4kDD0uIEY67nPnUGvziLLbrNK4IL0zSo
xdz7kmylJakzfBp8qx+QoNN73nBwp1rXQIfy2Bm/mySyLUXH+drs7oKX7nfIH3W2
zZqVQc7Y6TZAGcZ2+gJTvX9Bd+c2Z4NfAu5lgn9LYrNoSfzUYDpxohO3kooWnqjN
CV/Qq64Vai5BZj3rc8cuN7t8o/MF+HMSTVlD8Olc7HfsTRb0HDCD4pW8vdz+ld2B
3keFngZA7suuRISA9brW/luBtpJTg86oEvKML8UYQ0CvE+vFx19U2Yv9tEH++DNC
UEtuR1gtqIBsX3jitbMZ/ol9PdVs05mewqZjFe+97IDshKr0g9HOxfBUGOP+PEju
Z4wuHz+nVFYE1koJv7hKcu5utkJ8dtxe3wxYmOhPifUS4YJZHL4VdTahp1qKWlUA
qwANaLK2CAHSf6Wto+QjXz70ay89rvOtxzBqnsJ6O4qlKoTIpfvmOR8Q81F9xygn
pFXi7s86F0nBMO4GZwRx6RC/ErmotZ4B3CLJ9Lj6c1QgbBipUmJJ8AE5UMUdg+/G
Nq/PX+PCPMHbIJ/rAzYZ9dD03t1Sml/SRz8/sZridN87WEHAkwQQy0+jzfkhSQIg
pB6zwCESIxgsSBEO1wovMrFgo5V0/Sq/YgjviXTFI2KzDdHKepmaZHtSgcg5lNDv
47rvY1jQnbN0sGh+WyW14ckIzGJt4zCtKffUV7vaZRMMFLQL6WI8qebdELxTu32R
FTy/GeeEZj+PvBICP8suybIoitHQ0rpFNj26npOv39/nDc1qbC0LKcE8balHCYh2
csqXu6R2SPls9dls0oJ8e/G5TmFFz4oePup+3zepVUHsvyYiOrPtXvxgcbHdTaJF
1EMsff1x6c82k9SAvAQsY2t7DCwHmCioB4FidrRwHqCfD59ASymJGuxghdCI91b1
rM/l4xGhinOQp4SpNxylbWnvAsdWa99gLGdcqLnwLCbNjlJZoPq8sBVMVeZSw3z0
oNxfE+klQaXuiv9hC0RXKx/gQLT8OQNcIZoqe+uejBoLo/y2cTz6GZNHPzxYQw6l
XAbjeDioC28mTUbZrIDJEBSVPgFbw5pDWG8iik21Bq4UZL94ZwESV7JONTw99hlj
d/nZ1qCJaVJeI5kudkkfZQGLZ+KRVIOxQnWxNCOHJgLEVpLBDH2Lua6GvH5FVZ+4
AiCL1bZhTl2kAj6FUxBb7nunLpsOihNKo2ewL2KuSkwbO9GuzSSpYvU7VGEioHNO
EG5v1uJl86+MVrLaGTNtzPYwBPdq37XLG5x2SAQeU52XNzhmnj9xHUc2F0OaOetu
8qThIL+gSDnBkk8WCwPEKALtDvWSa0BJuRwvYLTfvyyfJfms2fYJEZOldhin/pwB
OQ60fAW4LM2geLhr1kPAJ6l7x38L3HQAi00ngP3npGTvBEVXnVX2DHh4YecPdGS8
aIgwgkxFnyRtn/jLSAex54QfR8KUhr7DaUPUgfj6oUkNEvCwRegs5T+jpaQX3R0V
1jgpVd+jcglRiAnbPoR5KwLd4jzM07DIILgsWK8AJQTIYP/4w9rn4t2rkoRMrEZj
2PE/gvUSEcZjb2pLLBvba293z0dz2iDVQILVZ4RTnqcicLkoV20RgeqvP5/hq4DX
+pVt1EbyQXjm5ZtKBbfKny7o7YKFYbFqn/O7kyamHArBO5bWPoMGT0oiFMd9jRRV
T42ybRoBrFyNya/JE3jrIcfcpD+5JmHuf8ZC/CdGog69bf0YgjRB3+z2mSAmemE9
nURZ0vKdd7zEWGl4Ohos8VdHPQqPVoI20YGg1umpA+7rLd7MlxD7ebh0qXTQXsyd
D4lw25ez7MRiV9ncIAWqay5u/ETajmybkt88c9x04KPHxtlFCqwoKEeQCjaCTsmf
lPLtdrEeHUM16y1+5oFsVC+uev3XJbznCJTX8MUHP/QXkw2GE617rDwfoiU7w/iI
HDBnA39VzoC6ZvEarZSJtPpRgUagAiH3xejhu/V7Lci+Pn1JjrWLWjFl688yQN7F
tYntwH1tDju04MyeuY7XBOhidc9ae/OvialgzCjudXQuWJMbPLalVr/h5VeH/U9U
8+iemPU72vIFtUt/X1S2p9+gC/DGs2IYC/k00JSxUNY+Ve/so+7L3scO5aeFZcBX
pprSskt67t854xaQheZ14FBmDZOvSpuCTdZkBEtPnxadVJ0JLtyK0WLjWB7xUgIE
bcHaiDwvz9J0TsUE2vj38hFUqwtba6vcPpHvxXiG2MjYwBIHi7YUJwWF4GuFv0m+
FNVpEwxygF7DquiyB6OHOxHSWvK9QxWXn1heNiDcGw9pQDeVdqE5IFxNQassXdBX
o9u054qr6jCMD9TPjHNjAD/QtqohJFfCBkctIfCpo+kRP8EB+Vcej9Wnnz8chcdp
NP8GWt+mLF9KsLi15cmoo3bSyoF9+PhLYSkThrxH//lLhAwITJBfPpaZcxd1Vux6
KtnED5dU8PyeH0v64wNvmNAvmsA7nlKgHEIhc3QArQ6Nsr1KpAcJ8vBm/gJOEWTe
Nje5hskKU+Fx4fklGHS6hYxzMG4QV73I8ZiNtaGWHStfPcM+OYQUMQOGwh05uYDx
xxpnVn1h2dGsM/JNeusezjqMwIjpxO3TPcLApdOZCI8xdOpeXDg2LNEFosVeIRLC
9luMkHKYLlfCu+jqmHwMrcCoHT/jpyjBzUx2NS5OrDDY/dvEvuS53BrF+9TIs2lO
Xzbp+0cKPHrmep3sIFHBRXM5aqA6St84g0TFSLJebnpkDHLPZTlrGUpMja8fHWHq
LrqX/ZMMKjopCOEsIZDEi7+TCgrEPJdyrtD7DdxLI45Vf+uSZEczgdsooTDaY80x
PKewnGMij6qV43GkbtJU9Dmg+SJeUrTKMd/n8m/f5fjEtYeqKwb7xY7MiW0hSGvA
rPJUwXEhsfdneynlwLm056V+xVOJzKZB8mHOb1IQgcZqdgUMLUFJNA8/Xvnsylvo
6H3ANAG2Kt1J0veZTwIFhAYd6cAir39mfOjMk1WMChNuHak1YLpHItSqx2gQdSJ+
DoFSVKBwji3nUduHK4q9yoyFJY6Q6/nhbf7Ce4Yx8W3IGMyUiTvAIVqN3aKnUDBp
aeIWGQHAuz7Kvymj8hgeQRVd4tzKLZdJbMLEUMk4cHUYHk/ZFwIONbH635Y1iY/J
LpjafigDid1Udnz48L7EJh3ST+J0Qoq/97yHGmzotrZuCAi32y5djNpO0PnNuoAr
sqW28kCrDcYYOzMsxTnIb5PvcMlg9b47JbF+xPtoXw7CdbEJNdtHNrD/fcbOgmZb
Df7NiytRpWX6f4MOv7zcsUkcwYEdHTL0WmTC+41h4jn61r9el2I7I2WvSrGdfe3i
IfraIv/DdS/2MtgjRvMDXd5yCKuPYD0B/ruEC3pvSWab4k9GOEzOffx8RDP9eimQ
U8rn9W6EWSiSLO5frUUe7B/MrUk58oDlfLod8nUTbW3A5jzCbmRrPPTZi/SJkhNk
WPfA51cQcuye1GGcugp6LFmpFG7RkArR4e/4E4UUJiLm8ztSOaVh4pIteGCeOovO
QoXkBiisvRbXM/YmDkRGonJRQ+fv9CuGXlsMwD8hTbVMTxHRHvW+ZsCGHJ/HhLDh
3Yt2YvnnrUZJVT5eyrWP0VRULTEHz5TG/PH/XuNQZBsRWNtsAQH/q7543tXpWmjA
WjCeht9vCM8t4tisNAN8LIELyZG12VR92LfZIKKNfExPpOyzmqrsZ2T2HjoEJvXj
ER+HLPHLhW68Wt6gOACk5crLZVMyCn83MFmYR3Zur0UMHgizVvOUhlui2A0eRmwI
9e11bFtuNb0dUXzbtqa7bguxcjAlPrRzOjnDhO75LO7gkAMG1uNmdY1dttiGnWfr
G9QH8C9I+hHpygxVm+BIgP7szeyCLIquZAtrp7SCVL2+E7wTCjGPkl5xjaXnXgDs
o4XY8HNMgTUmlm7rWiycI0KLz1rO+Czg5KD149b4Yd/km2ind4LoVI3xVs1b8xsN
AOpmpv2S95WzrdJDJavA0h8BYlW8Jthz2nRJv91YRe1CEzwgC1bk9nrsRoiuOr5n
2NAkadwb0zAVdsA0KFWdPA3WKTQVD3hTm1mK7x+MjQXfWuQVulqeL5+z0lcqYfAl
acv2uely/ef4PHF/eWbPjeDFVrmZNyEenRwI4VAYcgZt6twPjWKoSKcjQFNuEwTd
bXAmDiIn2zRnEAxXhZicxP+mawolIYg9r5PYe6w153mk8DrQicFKrpK3URQn5Z0t
ikdGQqd8RC4EIre6vfq8vzVIiebS/ZEL8Oas7KjzAnESxyVi8MYATVzUzVQiuUPm
kaq2FO1TiDlx/3LxaI8THle6v/jIwygwBl/a877xhKTpMNX3bojBLEbfF+QdV1Et
QERh7p/Ciq/3daiAJ/cDTCZ7aoj0GNdUIEQQ+1Mwbw5gp67GVA/kgtC9TgLQmsC/
loE3QWr42WbyJCBnpm8VAc3q/ZA0AnAMPAi5pmbuJGQ60HD63E+IciJfR2oR3i0p
0XxHStBoj5xaTEx4ErUyKjTONPoXvmDdJwe3rH0Qgvb+jdSfZxZ1KiqoU6swPHJx
sN2CIojNUjQ5zWWz6M+3ohmubZd1WZRdJGSI2h0HwpuDa9SQDDEq09G/1anbYTCT
RZ/RviuS1Z0wMF7jY1GNoeKzvwy3s3OLfNRnypv68ROqv0UYbKxll90t4hN49XUT
KpyM6iB01i1v7fdyLL+/PRqpgXQJvKC7E17HIMQOR/aFfrA9juw68069nKmRahcS
5fR2ZwItwJaRV3QuJQyLyWTobA7hU4Wwz8YrdFIBRiCFCJkZ/2Dqte8IbW0Bv3xU
cy79NR49JH58SKUcbKNDbaZhx3TTqIsIG6+CtCd29oL7AJbXDOJHzVkZCv5Z4xuc
FmDP6PWvLje4sLdlVrUygoGNDXIhCzJVjUVOblTH0vpz79gUviYb/kkp9hbzQZ32
O39Tl6H/YU7z23XLtAGAgUdqLHoaE5sYz6hdUMETMN/NmIh7Y/11De/5pernFEuI
YRNLbhe93AOA4UHPsXY1Ii/GyI3fByt19yFmV6THcP5swW+60+IHKdXmfPg6JhoU
0MJGp3/C5R9lg/7q/IVaNWcccE6chw7LeZ8/g3pCyacT2W0TNCtmXsJBZe34jwJo
9NJqykYfQ83PolvZkUB5qtRTmvE/cYiGEZjqvBpLEVc0dPGxOrZfNRWFCiD1r7GA
oWlEqM85WReuy6fVlbSr3bNcFqeOKtv1P5ZS2oMRTKcQ3ZnqCjxn0CG25Ol28Lyb
CIkym4IZm+qQmaoNITYu3pJOS93H8Aq4zIRqnvN0sVwCyNK6IFcVSDcewEvrPKeX
IkcxgEsykSti4MzgvWCIz8Jk5hi+c6u+lSv62rRdH7it5iEf1H1SLGu0yitD8rPC
MpbHIpa+9BhrIOBdTsaBVYF65fm4aTnZR5D6+ZdqKaKhbc0VzKafh45qd105aw3s
oyYQHFLU5B0xnlLpOlVFR6oBa2QjzbwEwFw+DkwAyvlIPqIc164WCodDba4c7yJ8
u2HplpuhYPv4NYGgokkXXI5KYD4KW8JAcsXhSS8OShI1zJLKChilCW77t8ZrSIzF
lidg1yPc7tUX+QODcCBYvxJToYyST6dhK0U4mL5pzO27HGWH+Hn/aBZcZwzlXB/D
v667J6hBEmueQAx767G71lyQaDBKa9MyEGn7vyU1OCm79l3GiUPws9dDDMPe+fbP
lyqDedQNcg/ox/uMuJ8PVrvNekTcI6ZDlkyW8XkFoW431CUgGohVz/KHlJ5Q4mPV
v8rUBJytEMdQuKTFCLW6dwtTJ3g9SNfcHemi5Phj/Wnt9DqbM/RomUu5wwoMWhu+
YI7/X5anPZLUBc9fToPvH46b7W4+uQHJD7VUHY2VyKxdKu+VC9Sr/e5EEZsTLkqM
KE55Hxoh7NLLvYIzHiBb2upboBl/bORBm0GRU0lNb5FxPJ+DgOD8UsbZWs03Jgvk
AA82NRpIPFFztu1JrP9X1cYWkniPQOnaFUAGDOo3ZbUkECYA0NSt+6IkstDvl1MQ
+h4Bh3iZs2yLWkdGR+V64ZFzdHc0at947qEgTqgsrzfspOE5pU5Acbhb5H428JcQ
i2KN4yLBo4ulP0ALMb5+VLX6iERgIpvBpzdYtTfA/zLG8aUSFkmk2GwWiGX3+8U6
Kk/DQ0zl7OUFre96pwvaOhhFzlCqj+gGxNQ1arMSXhcar7dEQV5bUUIEaasRcjdX
dcrKIEt0X5+XQ/8f/PR9q1kSXZEcrdbgBaCQHvoKfYCDtdg6173FSiAmOFJFd3eo
juM4GzVdbXaWFQ7/1HUe6VdrNjMv7ws+CMpL6o1jEAolMPL8C8L259SnRK7Z+yZm
yIjFPMjoy08gNWpNJB59MPUUATQFyTYJJQVIHQiNkjx6Quuh05jSdsrd5N0QEkqh
EGmvH/lJlH7cI5aMEUIUCBfRydlgkj3PfKn0MK2706j1wPGNUkQ/LZDQt3ZW80G3
IKEdqPM0z90j/zyoqOT2XyXPuMHmJuHLvOhuSf8+9Q0AnFmUbxQ6j+H9dDYHC9xc
oOc4TrbW9GULJf2s4mLmAgHfs6bwY6ggInWRMBRH5i9BKc/EfnBkEaNxY3zu29Pf
hDEsvOxC3mEhkVILXKaM9KyjqvzWQYsN6U/Va9HkmnTzB3MJAr0Ae1xvDepokg0D
53JrEeIdGldBuC3JZwySRVmqeAdcRKboGMi+hBbPZjEevQ9arQslqhX1qwgKo0f7
2BXfKLqhb7nNOxxJrZkn3oGqZoyNiIPbL4pscu1YoeMKCQcuaqeyCgk4Gu3dQLiZ
bvm0R6mhFb1/oP7JOGYscURZBzr+UuHMbNNISDS1tjD3ZvSXIRaVx94Z0DICU2zn
86bXqDLuzF0SX/vXYC/qQp9TGvFhSLiXDcqOot2wqxE9jBF/Y/oWJM3jPsWclc2u
5AJFMIX+YGy1R0cE+6589e1Wd4olLfSUPxJTVIr3G82GgX8P2wU2qfIbGgb8eBAk
SqsF5ejtRKOWq8/WrqV9/N2o4mrTNTNsReqHe95i+Wg5/BFRAp0CCfdug3O00FYx
AseCxjmdnmQhJxjhuWPFD1WlAi542Z3RWo4R172MDtpHpZaFloq4Gb6U+mh7N4Zm
TngFHd7q/g5eggDUY2rEfX+p5ogqm85Zjxkmb1exs+e9eBTAfF7V/r2vO1Av+5iT
B0BsANUW5o1nSLJHD1K6bOAVYlKNVsUK/3r0CtHLrtx1aRfDntXZbp3vivP3uzOe
0JvgsExgrbi19djdbXUqK+qh2J301t1/2okDMzOOVHI6Y4MGW6aJR1GIROYundAz
tV8ukkNR/oj4N7VsyZuuqWdr5DIOg49xkx5tVKOINzBzgtDwJmciZUV/WjnVRG47
hYq+J/rtJurNi19+rtlbC8/yPdugkkvaKxSUlVz/z41/XfgEYbiFpW0nm73JqC3L
6DpAn1D/DC2wnN5tW3Ti6tO5amxVWpZUjRr/rU0a1mGeyXFC97LQGSKf3QwSfZet
C8aSUpm0HDLdVtczYlFb+jxJE/tSmDYmVM9ZPMiBKf/HJY3+aqy/VnCO9b7ZJ8l+
Tl/zyz579dirzr2iYWYkSjT2xOXoMujtf7XD3N2DlTXwhx1aX9iAM5kpMk7a3YFU
8hs+oITo03sBWOxh4tO2VYZFzkrbd3BLimvm8/KBCpp2DCo62L7/RgCge1zWRlEC
wEf8P0ux9bAdTD8KbR1CJb29HbijVvHQUgjJr8sfDAol4fW9DuhZkTnUTz8/GoY9
vXeA+fblyzb5DHkOfpr4QtDf/6bDEr7/lgi5Zi11Mj8QEWb99MmDHfkIKTqJUY8e
MpJv+hKX/u3h5hZn2SPo6dQXlHBF9ojyyn2hTKUyQY11SYmofhVj13hPNMunxq8O
17A7i/tmAGD9WdoHxR6bSUZBtimmoYJytHKg0Gw/NP6GGoyN3O75IXEmHthYJcHd
Gf6L92J0aStuZOTM6iIHmUFcuuzYG3aLpUwRa3TReR1/YR8f2wKfR3D7e8qS+xFM
P9s2AivxRe9gtPxeXCZEpp6KXoSBcI6e54sqQ2hmOu1cvnMc16eUoVql1yPYoaXK
L2i2nPYWbV5GoFANRx2Syed6fQptIiGG5CFCpWyH9RWCmYNW6+oRcKASVJbOWAmi
8kv7SiyduOFko9iVvy+5YcKfED22Ur5pdphxX0qa6+R9xJpnvZBPGxed+avUjkhM
i3QfuA8PgYxNKWZGy/PzSc3sZG3jx07ZcBsboEEHejREbHwiZ7I2J383of+qO1vT
dorcVPzgl4g/ygTq6oLRSSd6X7wZEScsrM1kF4jIINB/gFfgREZBPnKs2KYAYVij
IJzSHn5utSnyzq63BwEK1MZofH5dwFCrZkI3u0fnPoOQZisNMCdMSKl5QS0lTwoO
xZYyen9SDQ3NFyXW5Byqmm4aDXkd5sWMz1nXWsNbFNUf8BRYsBAgfT2IpOgLtZnt
YsLfgjDdalJQBVRSKqqr3Wsb8fm4xdHKgKeuVUzz7hrnfE3bdK6lZvLiNOV9yOB7
FhtnfrQCrtbXzLpF3QbReTp1ODZMWO5nNJ8g+pn95m8qGsxbqfOB0CcD7cAXgawW
uWHvQ71O0ZS4P1TQutzF/DOmLcO5nZVIzwoe5pJgC7WzLZN7dBbA5q3Aq55R92KE
sqB+ScQ36naSe2uH7SFAeK5HtrwT9HNVJVTifzL8pOmFQ2dppzFTTaYyv7w35SOt
cVM5htdretHftN+rpWxx63IjXM+yTzb0903tGCDQJ8n3fJviYJdkSkNcp+xBKu7y
yFiUvQIediFcBqJbRAlWiMVNXr2rd8YSDXLiBxnJS/dHua1rQ51EhDpifCmJ57sa
nMxWz4fMd+OYI+oVnsCqSHreZ6dA7tUCVP51D0iSniG9lJLZ26dR8ebVkCjh16pu
GHHFqJbsDfmT1xP8o1tvi5hcam0slGzeEjEesip8BzRD8Hx9SweekUpZbaotj+mz
XqpvEd5boF77M4l8O3C6UwyD4MUPt596ddWAqn1GOWNPuTBvA4IaLq3A2Y2orwND
YFoRpOakBTMt+SWIotp725hMaDa7AnDUXT7nxgfeDNsWFmpq25zb9G3NbHIztj9s
bq5awSiMv30e/pBQTyypWolrL1WYMkLyeh+x909mpg+L6ldpUh4oqsQbQ8uTB3xw
/RrbEauM7KTmpSgr2FnYnMGUjsaO0OXRleIRF0GHDmPNSKDjXhWMA5bzs2BxAuLI
FdGUCvn4ioWjNJlfpJhNHfAy8iBbStCB8Yt9300ALr+tONg+bCR1qYgK8Gzf1iBf
xzBCoYCFCTkEr+znRSV7K2nLXH2OjqExy37HErrdZgbRpTCN7WWHZTDKxj2yj+5B
EL3XspL2QWHPGgZ1NvuVTej8JIXMAYzjV81YEficy/r1EOkxVw6aZ1GRMxVguoRQ
T9HsMB3YXkidPZKEh0ld2VfMCkTvakgg+/mQj5vCwuVBAhJhWqtFT9HQxYOzUYwa
aM1FkXylBbQDvQa6mTyxI1sS1Fldsr0KFtMX7VIMEqvPSDKqazSUMZ1NxMhWPlxc
/gCeb4clJsRA2Qfz728MnUuIRADDcQeystF74hBJVUrSnqe0ht9OZN19ghM2kHBo
/3EqvNA6PQ/V8QVYxtF1g3zswxXC4E6m4ABy0xKXguApded5YGEZdRmpn2gUVCa1
mzmzRu/h18421ZvucDjtsLONePkJY2CFgr1WSLolvdU4guvSqdOmF5mxVdUl6KMw
STl0Ua5LkSw8HWuQE8fyIX5TNqhToebSBzrz4IBq5gXnwkvorgOU36Du9syJQooT
FxWjPCaz46VjYDl5CAskHZPGPmfzxRg2wkgXumrraKV4ws1HTZCOxaY2OPtKEl3f
m/0g/tcXjCfLeOWrHen1DJmU13+Fdwo0zXQ4wklS8mHfVr4LMrgAwGLivHTSmWLk
Z3NS8zYc0fP2eIi+Ubrnt5VD/CbjDoqTkIkos1Fj4GdCqs2nETjW3Kdaf9YFUzK3
oWx5RR6et1RfY0YQcPTm6JZCRoIhrAwMA1wUeLCxkKkFSxfav6/Lh4AAIqGwRZjr
+NbChw0ct45jv5aEsnrD+cUrw4glX3P/PvJJkTGTGQ+z+inKG31EpxnMABYpDrpS
ZAUjTYhqRFo8/5pLo3c2VcWtkKSeHC3zuI2GqRtjItdtpFJH9YHoq5qpI/ao4+yX
wL+63mTBF9JpuqDe9+HrFn797+KH8yK3PF/+KhcRl+fzmxpTv86df9RVViPPzX6I
UxmVeAxHqON0sIdYKtrCNKVPJl/MDIvdYiPpv1AZIpNVkkKwOrGaPkdjZXqPcYmR
KDg0nF0reSspAXEig7wD8NLj/UwqXh13ErgnQ5FQruyMiXYphyog/jS3lMBRWhxf
CIL6hO/WVk2uXxriIaHkKaMdOSZ4ZhIUY/Mx/ZWer9nwLxpblCEcC6yvhLvlqR+x
egKbc7dht6VKMM0lJSJ0fo8Arg5C9TDwp6BYSEWo+YLXgiPRai6STDxwi+5OmHnb
XhdNLf9vOeidBwx9wQAJRSqkpMB4Jv+q8muyBDfHPcXkpiJz/uDoGdvmo0K8Qo6b
eM91grGNhsBao9XrOYwVQVUZTpVvBQZLFQ74i6KllcabgmBczDoM0kTgP7hNGq6L
MpMyDBwJMz9Qq5Y+OFrh07jrUM1mFWOXR45ONnYZ8DX6933QUBO8ycvjxI791xm0
0aShsQaj0mmqlZ3CXKkUC6Zrn3jebFOOP0/pnmBRGm6UWGaSazxrZTiHEDaYHIUp
K/BTl2P+d61fHbU9JxesBzxI36SugV2j9Veq0lxqDBTKB2cW1zsWEYsr866dtocz
aMr0aStikcUnocDTxQWTH8dNLGsPeamyGSHjlFZc3lN8xLLDQCt5PDfM7qS524bx
yquJTCS8x/QFJrgwZ3unVVuFDOt5kmn4cju5WZ9O9szZMshOG4aRClHHVpqRnygL
EgOL8VFY2tMhdkNpsFjWta17QdY9tn0f36R5ChjQg55bBuhDqjKt0c9jGhK1rnoC
f7ADPvNFMHwsuPN7PAdEFFt9Ek0ehO8/iNKD3Te6kz0hnrKjAIjqfGOL+Kh1Xjvo
MWV/kIPg/QmGppKUMk2x3lZUe38SeyFVW/AuzYMzpm/X2KL/5ZHYUP6W3avXLtKj
hMwb4XnZMiCOp95+9DcXKwnB+2tCdxE+kDCPEKKRdLlTZpn4+2xxWIoTkCkMxgMC
qs7SPbf59Mz3j7QU8N962s6W8Tocc73TFOtHedVdm1WI1zTNS1rbbP1oDJ8GOSYM
mjxf57G/MsZIckCCUhmdYsz+Y0He0TYQpeOuDKZ66ItROWojWkc+WGKQTsTr8vFM
1mEhHhHI+7ZDUMLPKKSDfqCP1ZIKh/IwUCVykPwJNnig2FW+voaCHyGWce7Xqz4n
1a3mK7g8jNyj6xFJz8Um5DSY/T4tNDrMQsMhHK7fAgbr22Ts/7gFSQjog4P/gkdm
YimugqUpR7iSh7FysIzpL9Xt0y4UaluYW7KvRy64iOOlnzgN41ZHYkq78c1wL2B+
PpDvnOzYw6EDLFYVeQSh98tKSl0Av3txgbtG00/ODUh4gATq4GzIePINzWS6Pl3I
DIKc0Uk5uhjg6/y973JSDpoeELXlH2d/s22OeDi1aaojyo7H6rCfH0oS1fmgUy7p
XhSOVfX/MyJnH2R+VamkgV6/tJ3NOnh8pmZZaXtlUcMRrmfEHs5kQ91kIaywzHTC
rjYLb//v9TZMuoOYQ82HRJXpxbcRxOIpk7kh+00fhrUhcvJmIJVJSoGYlSeUTJMg
jS37qoeKxkWvYh/5tN1fAblKwx8VTetcpJ0akFvArbma0sxYnR7SAn9fO2FSYULq
GMvaapc23w/Gwxu54aRdXUdsrghQAbYPOp8p21iVycaY6ZnY36uRKfAQEG82FfVY
MTGNwJbQYB6evY2/jtp5ZO9xIUNZZ7czbqpizecPaRa8ob9Wgs7vXZakrRHwOUDd
sZfncK5GDCMSu+GUjffvm7AjYMnqaVVu1O4MPU1ntYKtq/pyYZ+zi7CPuWotVAT7
EKFIK4j515BqPVVFR2SDbEc8Uwb+faQ8yhMMDjCguqYWfJfwf6yFBzQdnkwi3ujR
W2S34Nk+PwINvKI2xGLNAuHS4/jlwGpbJD9HujxX+VvPSyySL2a73C/eWfNdI26a
KvcmV6pog0IMeqhHx21X7hlq7uy43owNlaAnj71H3aVobubZCfqr+tPJ/7MYCrKe
0ac+bWbR/UlFu6OIIPFx5RTmctRNbVD5c32Z7/E/mJZxBMCRnLNOUSPbFqAZ8zE5
YUBeflarpCg1tBAEeyJNnnwxw2x1TQuJzlhIq4TgbwZkh5MIZCQ8mX31anj9uM0t
skG3FJnF4tIN0YwQcZ65TXhF9FBR8osQ5brRQOicntxzZ/7TKzFNWYudLruVDe1L
rFfewKWTiuaRgp8W+UQhR/TkuBtCR1q4qABcyh2bXuH7oTxAKhRs6NUxdgqD70mi
/9qYn3VYNblhj7cTt2k21613N+aSw0WVHeBT4333d7PKXAZolb+PXk2+cJiD6BN9
Jgz6yVq/2qWqIwurbtEfECXSpSxkZsp8+D4W8JRATZfzT10QHAqRrQBtS5qpKjfF
kNR6N5cjS9wZx1KEm47+lho96P10nLIA1EEWjlrb/+LUvVaBBl4gLMP+jhRwgmFJ
vnDnB/Opu8BTcotR2SFnHt1+avjY3ZV7ruChKU27SDgx+OV3bIRvLQL8Q2i4Lz7z
mLzbePeANZPhlBZWJsYDiiQwfMUTxKhnKVKyCx1yEd1A3FmzhO4WdTPHQrmzlrX4
SWGEBysjhhbY4MQDejn5rfGizsLbmF2E7GnNgQiaKAEv2OQrgENvyIoWZmJ58BgT
rFnaTPSnKSrdcLN4eSX9/Ta996m9lcxW3dvH+gJBLyhNCinYhEyua1R6XhO2fqVN
RUBvLNK4jQ3xBDsEBIYM2ZViVyodeUNPp+DjV/YeiOE9VQVzTV6Urwaji1BJtzsr
MELYN4+oa3m6uLQlyxrQh+pqTTY1Z9MvjrPmbGPcrzgcK377KM+QSkGaFzAT8ES2
akvkJSF4APD3yyeFnn/2ZL/tYo/kjhsmVsRoZi57jA5YWnKqKxDzQMzaqWuKsflW
0DLikxIUEpwBCgk2pG1cV1hUPeIXE6wMQHvz4TcmGez4j1u0vc0DP8cMKka+3H9g
gP3VsvaWedFSDjS8csxpsawtVOfLor01h9cuwq0ba0O4wjZz9KmmztftsRLmZlS6
sTn6rsWHP4fDHgpX8PC8r8BnHCia98NNnGnP53LvkyOgFbd5/gfb9oqPSLbnZW52
K4niCR8+dGRSsqa9TXoihZALBpsd6+s00goQgU0Kb90CAZPA0obqU3xEzp92flwK
ZXlNZUDmQ+xD3aDVxq0b+RXkPws2i8edUFZRmIR0fo0sraMEoLcfjbL7dPtf/EtJ
evypQmp8oCfINFUmdDTx0Z14r9aNcVbi5ekCCN3Kr/Ql58DaDcz63L+NqXq91nlA
N0kV5xBpmuk3qW3xc3gLLZSQXGxup8WWVgJ9gWMjQME3+3G6l1w2bFGVGQR3JWxm
nb2XZth9nQ9S9Ir3jPOkEN6gR/pLWXID43iKBQJXpqCg7dlVafmqiG+GZXhY4sD5
Zua8EjOzbwscy9Cjn7OZxDv7nglT3jv107XrTKycp0Acs5H/5ZEArk8eVsfUBlXv
Rs2zTYjETkvwVIcZynXWJ9mCWANapYWVUwhdt0b1Apo8spiDbbLOzLVGvDDEqlAK
JeZ5MftnsRT2whVS9C/53UQafk7HxWsZDtvUX+farKugswu162Va4y+FxrofTqts
jN3Xno4equHHUj7AgMETBn9sLLjRGBNpDxjjj5vb5olmYGiDagLwhpEuhLrFQle0
tju6Aem6aJv845mAOT/Mjx0VWmH+t3lE3SwoV1Uny0V5Ougms63NUqntxLkwoAWv
rpgAd7wcnARprpH3qUslI01R2fbLbZCj+BDEFtzZL9jTYhwguU/GGncHGhx2jkZx
TRAwx2MKUgjBKHJCgjtJq/9yjdsBRe2tXx1uPN3tVMtwoGiRClAjT8fRh+xIeTUj
gpJELrokQv84qZd3ybdJK2LIEfVuggYvgljQTy8DQrESXIakYi0fONFMCDQU6Glb
UvxrUU2klbBsw+jxN8AgRVh+8b4MA3vGMcT0exlpFa2Ix10WmJrS8hOCPjdD8wpV
YbUYNyOb5WemvACSbA55gTQzT8ah7VE100nD6CIRT6esNBHfyvjZ4i0SdERtMC6X
SIzLXlQ+tISf5we1rYmxoD3MGNkNOeRz+PB6skd5b0oyLRa2E+rHxj7/dZiRTN+Z
IgUt0zr3NdUkSl2MfCgckFUcHqj1bXIIvpsyNO5Rd4I+/cNzBAENdsvi4uyqf0lL
nioqo0IKxPyxuMpmM0OT050timkAwVNnFjynt+YNyVFbEt7BrPB27uoKAybtXYCl
zpp8knOh04ZPvNroEJYPYHvtMPmx/D3fNJT0L3c6l7V75XZmdbO2xdwJUr5cme5t
et3pIIKEjgVDtxkR4/OzxnAGfSpq+U+yy9ML++p+ZHSs7/aXgaOXUn5FqN7CMbCL
d3NQaKjvXuBga9zSclTJ4Qzgo/LFwsPyiBRUG+4RwV9OfNckNVWuCwkbl8fPVkK2
BdlaTCkO8q0CLKsopKIuPdr6wkpJa7RuJnQ9vW/VeuyzdwuNSiZMJyhQTK4yjO//
o/xMGopfMf4sHdKUXJ3axngDh0Ks4lktzTbjjhTwGIJeqa/Lp2If2R9pG7clPzj5
gIuRTqMKcsR8Wtv7cldj2CIaKDuIMiRLcolZgrBtGCa4RiYDk8ynvcbg2+HOAVad
TQTal5fIBK2Spkz03SFZSKCBTH22RU7JbAdQm2fKpjP0ICX0GhwRtJ076RyV892A
S23yEark7x72gzmsqb0vJ407F63kfJVA4CXSsitYg8gGV2MT8V88p35CGeZg41SN
uFLykLO9hFyv0NPldrX/OA6m6FSGCJ1siALbF+59Z9u2TrAeKvfiQdktPALestMB
FG3QCgdizbPfTf3TuNp1AQcyZ4NO9KwdCgIb6aoUXLoQyRQI2YGY2jFESQycUwaE
TbcY9QBWQESkitGx0p2RnlpsGEM+HzsT/yU080Xc9BBJuYRTDWdaVLn7AzyblKla
FlhjUOhiJtCG7jLiF7KVhJjpmYkrvuNCXD/xroOdHVqLOtffalTL27qm3XsfLetL
82R+tNKJxXiCDJp/jiQvkxeEzXi3qaeiD4YXwvHXARhiZ8AQrQzpTZ6C38FeytKn
2v+sIkuKiNC3UCEhND+t8tUvveeyUzC2NsLjWEgIHSrtRWT3+tIF9AWH8MGIEzbA
X7CVMB3aqIoPyZiJ83mGgLyCNwGGI0Mp5TfTg5q2gTssVzdfvTtBXA/TYhAZlBuU
CN6ppM1J2eTXfkLk1uyLRO0PDnihfHvs1awgHzvq+gA2Bt7vusihlyC+4/LczLoW
1H2Qfcdkmjua5qgboJyJi3OXI4ZLZAb5HBRlma+RDNdVkL/jJJa3udW3ZIfkEBTz
2VzBuAiemvLFSoYILCC/Ki2L6/R7ppFLHOMkYmbyis61oAaWMw3ThX2Zc5HkAjwG
X5YHjis9M4wCpG0qdTRW4guMuZN2hIf/3uC8HfjU6+ZdSlv53DE4RR7J9tSUZPQF
/KP+g9IHxWjJ3JqWUaHl4ZjZ78i4nQq3qA5gjSZmsLTqHs7ARYd4216xdHUXjTzU
rmjtxx4UyCKT4vj7MHHaYuPYAn/qwtUKI9IzgyqcYRWmUsdiZnzYCXWu4Lw0jnWp
JnBsI+pUDPuhz3pq5baRQSHzugqOiI3AjggGidk/vUAiNmHUs1oMeh734H31dZiS
cJrbmauXvZvhmScRnMd52hnALI0TBAVR6SwTdEAmjatLStbJCV3qfCsGyWpcrJMu
vNYBaicSVeqABbEDmBNE3sU13r92Wd7QZjPxZ7/QcGDQDJbfZddUY7z2IwLbrMCI
FsmwERAcuUjD0Ek0OlpMueNQCIPNaKJGq9E8GzWNBgfr7x/2/QJ6w4aDOpZldAru
xszxzxYGymKNWcJLyP6A9puDFYMsxALm0cPTWiV/jNcrDXLrGz4Jo+rBVvmcIW/1
N7rwRzi/8E6iIpGWuMZc6fEpGFpi59ZWJiGvJa/EKDgksDFeQD42A+zCdDsvTykB
vE7VtSiNKUhP9lcQQnxfM6a/utOsLyXEo1D0dCr2XHa/sRQ3Z5uJGvozUo20r9LA
Gj4qNxE1DF6RPSeoIWNUix23LjL5Li9eAOcJQ6mWPRY4GMAWvCzmBfpaZ/ANQ95M
Z3J/pi+YulAXFrP9v+pWEAsfhE+HuTVz7621LGfvPiCoYdZHL6Ys76suMSkd3XpH
PA8O2Q+ME8qTtZQmf+3Mxsd71C6yIUN0LI3Z3psZZ5SQ+9a6YodQnHy3Xahnwxab
ipkqxgPkf6h28kfszMmV40UhJJvXyqzjdeDZ3lWT7StSuui5b9mJfoppSbj2McKK
DqKCsNt0Bq15l2RoPyU3dS27yB6FsndUGFALfe6BicA4ckUjWha1QoNW2smoEuTY
5rXLFtcVhanv41w/fX99+qewaXAXEXHiiZn3OQFLOYbUxCPTpcQtqeoZKJ2oYF/j
RbBJvhP3QWWOrUOm793zdXISj6NdaL92cI8fGau6cJ3wpYje7fG/DTCoP1z4nxLz
0vMUvVlrSNQv64pmpgRaLD6yhuy76g7/LcdTxOEWhPxLlkEBDL/G3iUX5jzXIf2X
vPqLy/V3eyir+yR93NB6+zO/LHY3fFettxYtx6Bm4GMGSXjQPGXwmiw1kNzMU+Jn
z4ewmfZfz/C+Fj7bKrcutbbHqbWf5PY2XWnyMw/l5zQkiCq8c1Wq/fXH9xlJsJKE
UqvbKkTLD54w7Cti0GtRjT2fxx8BSUfUtGKHbPdWIyAbDUMIJMF103jjyfVv/i/P
0FX6RqiDJ6+Zhcdjsd2kSIjKP8dDAhyH1Vt4w5p8t8hQULbvOkCgrwYKBjVY2drr
IGz37X5L8ElFmRtYxqjmo/2xXuIXlJ51aU1q9k9Pxzb8Lr/hzZ1VV3HqYT2l7+Hp
aaD97qaZ6DeQL59m8G/I6z7RkEDo87kl0whNafOcwA5kXXHHOIgPQcraxLY7VqeQ
Ch2NQtxz0kzMgEnH0Gm8piGCYGnKHYvJ5Ke3wd0u3O8L62QLPytQdfcuW35G4Yfp
quQLpVnfbz9gPdvrp0aeTG0wYPCZZ3rfVIAKGUJkTJql0fCk1ab+Zdod6EzxTc3R
VHnqcHTK449IReDFPK/ZWPUGK29ytgvkhCw3y0RZKi1dT9TWzWCoyYudAJub6tht
wPe+/faZ63VxiiEJDJVkFMwXUTmWiHuiosfI71Gp5r2er2KZoqnXMmdKAu0cVSmZ
5njG30aRCr42Ynul/lNWZEZrV0cdc7EPdz6TsEu3PmzQ850HtVz2W1amMauiCr9+
DBcyTj/xldXxDbiMnWpjlHNR0HanZq98tzkadw4Hg8uiCGaFKrddXMzTv5/ujJ6h
B+qALa6ONM0zj7ZgRu7xISjL9qoFhgiVdtZP5p6DgoFInXEcdZRzUQ28ERHIdJqz
c/5xv3z5bZOq9+O7WbZh89hO6Gro2D6XaN7usM9/J+8GzK9GnjSMb1X98mg/oSdD
EpgvpLTs8oEh7QF4BJJ6ZNTC+OgTnfjnLNWaukcjp/7XYP45/fgKwD+pO/zsmHOo
sX8+3EegcikoW7M9P30jywh/0p94pP2niYmB5uyVHBSQvJ0xgW+gX296B+xmnaF6
rY0a7D5gI+H1MGFGVeSc/ophtrOUWuWg1HzjLsFVDY6xceI7glNkk2Fcm+7Cr2Ey
piAoSW4vAIKYiJWUowCoB1rG4vRq0XfLzPRLghh6mhTEKkBw1EpdHdkcaxe0rQy5
mxuVYDGPUa7qqJA0or/jteJaX0lr2J3BFIuwzhS4w9qgxvqb6MAV+vvjWFycma0M
biXfFbaL877gDBgvdV+/VPPYIxQiUbzyEn2kB+ZsWry2hu2xGo+Y26w44H3gFBAQ
3cFtmF7mRkyYqUv8Z+wLfLKWsxvBKvLbuui4qq5JEab34a55jyaTZjMBjoRLMd1S
2C5ow5XQUKRQ9i1poYtI31+XJrV0DsSZ4zmO1+F6uRjloVdFYJ/dH5+gqhBFIb/A
gtM1OWOAcMzboqo8nzn0EUYKMrAG58ZriQLUvcnOuljnKp3iYbWLaf7YUmmQkmiB
0DnsK+blv2Y86x0zzQISYXEWMkgZ0Do1cgD69FXJdw1GsWydUFns6Nwp3UHP/BjS
9v/IOGHKPpzIPZaq/s0WkhsbZZFSaE19bcZGlwTtzXg5RJKDVKjT07AKL7mnYiOA
JN2sTjAaXrfOf4mnkrb7alDgsNBtTkd1O1D/d+ix2nx924N9vT8qyCEmDbrZ6uKy
LvN6cfF2YHCu/f6WeuKy9Q/ZvWP1HZ22MP2w0VgM2rIgHhkeHrgeJyrXghC38Bgr
fiWmzSTNhgpnqEzcf2uxRYm/DOPzCHUb0EbOWdvOdXVDwDPfGbH5dqmZ+Y+OkI2/
sGTNBYxTaLwr00Kr5kctE2H028wSIj2VrRV/JjuxrO9w7hFg41pKvopTvvpy5uJb
VmR0Br8Qyelx3eJxr7kusNpEgZQMTLcrI6TeIHkK2sthhmiA0tGabbSSknTqbtXb
T/R4IU/tAKdsDGDPZoiTV0/q2Vd6AugNe0g2G/tmSf3FltWfU/H1/oeh4dMHG0m7
xkYjmmOm1Jh/MQdTRHE5Nd/BJklTrFizNwdY/upY9IyE99WIHRpBTEBg5O+QvIch
IG6pIOm6Pn5xpSFmz20TmH7wotnTTsL4f0FG7yemSHLSuCERJMZq0Cnzq4Gwafa5
rqR7NWm4Dw6qaOYktKzeZBcu6YKtjBhLw7pVqycisM3vf6fjmOoOl4gNElLGLcEt
37iPVqa9eXrQ4WpG/ru3D97DqJBbzFYgUW1EesyVA46h7KHgqiSs+2PkInF8DMTL
sDWVEmeBJ2Xl003mrsAV7jy/b/uzf2Lk9sV6VKmNre/n4fMjH0QDgSITx0w7B+wg
yF0QUoM5jGK0f7RrShRzUSY/oDmUX3govCoVRr1g9fX1ut3gHmOUMyDWwE1po/JK
BROOEPfUNYIsdBAwG5RhDxR5zaoOVjwK6Jo6c44Key3SZmZMIB2C9J3QKLNVOGCO
qWWgQwki5Hy2+78sMjjaIQsYXi0Khkk+GrqsfEAJgjgFCRxQYwcl/g3g43Kchn92
3udS1LKStRoPVe81WIF4tSN0VzsI1LVquFcRizWzvbSR28HMZWo1lBwjYB1tp56I
LaKnX92AFISLyT5vyCQSBz3vlPR6Jw5I+6XYekM3svjLkyJA0sun2jX96iLioYLs
Au0JPYLXjjdklFdAxCopP0sPr0cJj/RIMcfAuBFu3/x7nm8v88AIDfcAc5JzK+cN
z7kSWcjBM0A66L/k1tCqCY/pgLwU1997Gp5hvL1RVJaX6HvxQd1EYk6Un2Ulqk8T
Qzskv8MEkNIAlRWf5GkAsx7/zSWEVSSwGbJk7QofJ5X/Se+LO1SdeE6o4dMh0EE/
lrcW0JPPqpj1xa0BU2KfqfCIMfEmqZHelkoOWBtZFovYmQCmbAji75VxnR2R4mQq
lSJiI1KPbYa+J6YRfBl2MiPXd/3eatark5SvuEHXdMFoX7YI1DPi3RF7IGtRED8h
5AFZr3HWtOIpgwI8nf1iJ2DZE7QXvhkR4jc9R+XMrRfv7hyxEgZ7klinlIs9CN/C
z5CFT4VXJ2U+WWW32fvpK+x85rLUYaAHneBt234+uMEzIlqj/zzQFgf70JVT1bsu
ZqC/CErFe6Mw1BaxqtIwT4TqZ/ow5vUHbgz54Y2IxfIKonI4JxKDD0WsGHhSlHV1
hdR78AqofZWX0U3Shc4XMfjoYeD9EmDYzLsuSRqGyhQunnKF5j2x182/pPjc+DfV
76H9ZsK12U7eIGi4obE9SJLPaKCOrwftD+xS04sURfER0zyCU4++VriknnVfhwBB
/jKfY72Srh7by54cUAxSsX708ThBM5weit1uKb48CEDtMwVRbtlVhAwHl9NW/f6B
A2lLnAvF+qlnDpIJodrLO9MU5CLCb85f/bCbYSC0gkuCEqpiUG6YRhTyfiqt4S+J
kxq+Lw2lW0wtQ9Uo1h6ug7I21APnPjSvQHvtm7uwYmRpt+gQJ6KXHSHuivguINqj
pSuOSUoC8QLzFKk0HbwVkDxcH8jDTYOS5BtVRNO5Zxzy1uZWtE/2B5JXfg7l83Wo
5TIF89kLnitfIlsjWYlD+tn/u0AmWq25Hjp3oGyHC3Q6q+vDxNSFxDzUqNkYiqri
fBx0X0XnuYX+ZO5whJ5X2Hp2IGPRtyvuWtbltEO+78yUNuvKHuoujKYytgAl5awg
E4uezfCyEgqLsjtX1NNn67cTXH5enhLeDivEDW9BBcBKfQ1+W+FR2aXoxZ5fOgrH
BM15PkuJMHOWbODqOs+BKAMZsLWBnBYNWf2T8xWk4G4Vv1eXOquhT2j3YhImmIZM
3GRfo8yDUXijc9/E0GlWeUULBzajz4NN9k8wabrCAGVKI4BL6qH+i8rylrKP7Kbg
8tscYO4KTFgQgSQFD3q8wtsay68mqX6h6aj05f8IGfwg///qMuaqEdEGdbHq54Bi
VJaNn+H20nm+Gj7GvioOHawQjG+mmBlpOM7by427pRg6e3BgtgLpQ7oGocwTQY27
F08mT6R8mEVl2uw+kwYBztyh2PISaKRwv94YvpqTZQSRthfZH7E3lSXDGgCoaWLA
2NE7+frPOF6Y9lwDc5DUC5qjdTrrbepriNbeIgG+VFAk3El0cWFeMP9NTsGKONym
mZXCAyyQErJMLDjmyBA/c13vgQitgMQGh8wPTZsHCnX6PCnUtELTteZSquuetR+K
XO94FFJb3Bcfrrkhw+Ecdw63pMsqkA22ooX3XJKilOl7ZzhlSmuuvLwAyNubPeyQ
4UDpDu7vQ1zPs1J2VSWRYZnGgCiLP5kCeTklLBbY12/WwyySwIF45qszBZMn0FVr
I1Gx8Gn92nCO+5GUAE2Fcv9APkax/Yca4FKmCxvOUiHVkVxZ2wZz0tGSgbimly4P
bSPJnUVbXxyIdVl+k+itYfhk9w6kHU0iD9w7QYPkvGtENsI0BijaNoshIE6ieP/9
QHVdWzX6us7n5GDpibAjf5BlN9xL0l0Ndx7KAHv61DHeHYdkYk7in0GjBXw6ZhfT
rH4cTHo1JTsjaBtBFXlTrJ21EzFfLGVp/tjHQo0k3Nwi1hnSpI6+FpIM/5gzEEIx
+cwqSaJWJJ8p4vAMvCOOnFqktew4ehdS2zb/Dg6aG0X40QUJ5yimxqAkbBI9HdVJ
haB+ETU+Q2k2ubTpjwWZLFctaH30KGBk3SJJ3wJylNnJRZAK/ZLFJmxRwVcJqz1y
UnPsU7vIw2bgRJXR44wxQ6VxXh36YlqXMiORKGvFETXlM434BusqoWzhnuURtz6J
YJVSN45CXVYKLDSrRVBhxhS9WD6SZZGQD/rYsaADMR1uJUOv44NLqqofSUQKmnV1
JNfmQLegPft9856tVmt6e3JadMrGSBkFf8vOapGuzK9//aBBpWcHFGJEwomVnsVp
8a8zuOMpHi7wr3FdnEzBVvuj4JJSuY3A+aEFp9RmpFDfJY+xDdTq+JmDbC9PNuX9
+KcepKIY6NeFeHOYaxjsXnpg9SUYkFgaYDzDwlCtYOK5TT8+u/Xp9VH9Jjy0kRQY
wVS59351YRqkeizzYCuBnsaJ/A3fnRDkg8PO9ehmUEtFUieyq6jHYCRnVB1Ugf8A
SyavXAK8xjHRrNoEoX2h/GBYBb0gZR6i+O4/93+tCZ1J0kaVbqUT8YIJu521zBpr
MiMWVmHI7wU+CmEf83XgGB+CaDgN9C8fpXgw2m8KNCSuY2Bq5J2aDQHTLygtUzsN
tdP35bonrMPFSabDwnkTC3vxMByB55n0d7/FNKyYfOOHeQaHFIoy/ikVmnGN80Yc
5ACn8NzuzwSQ0ENSBFaXjendr/FHDShEKo1Ro4LBvP/bZp+Igwbr9bbmNAB2MTS+
MMrflRCWYcePcPtFwB8dkxMrbTeEKn1FbqJ2ZUYsuC4pohoddwsQ75aCXzNi9SUl
Bz+GC+Wn7xX7RuA2hvZY9f6Bt4hjo0eMwcuUD7H/OkLJcXCaXSWld/GWrAB46fto
lVLzxo2HahjzkShxjULNEmVyObzZ07nzGCBlk/oz87jlp0MVMKg06QCUG7augv4P
q52RwJkDPX3S6nBEzOUcOcN//8WeTezf4QTxn5sZIJRtCCGDZmZQwHCl0nADFiAP
JD/xJwxNrfB8oenv26+p55HRIVOEoEQHn/sy9Xrb7AAzMUJELTAsFUAiXeZF/1VR
3YgQthheDoJE/Tv6VCk0twPBO0lSol7ASvbSTgWcJsLObPoAmjPnUkHQEYd/KFbj
U8+EJNoORgRJXHN329SyZt9VHQvNBRfhgu6ubWHi4gn7xUJZ00nxutySmMQS60/v
RIzER7o+G8VJC7JiLlka26rSH5BMjfR/S7OyFmxYGe0tyxBVu8fenOm3b1ui+P5U
Y1fk3CZf85uWu+Pe71JhRRyOBKjo6Hi3VeWvXa/DrwuM2sY2g0QbgICAuexV8zhP
1sjo26rfDDAyPQ1RahjdGWfK6Ois7zo3LWmXwrQs3TfVuwUXSm38FUAsRiz250Bb
snji7VgmyDuGJgq1535lE75fJST0zG4gDulVycFermjFSBI63+hhjpWQCW47jA+a
e3yHZJ9uQdeKnv/NHm+zJJC01PaEc7NbRT1kWZMxd6btA3IP1TrdTcQfy2+unKj8
o5jdrCGe+vP63jVK/7sZEHnmJ3jrjXEHOKsmjH97lKVkGK0svoHA9R6ggXqVEIv2
IO0bpPRvbM3jKMBrEzZ8TwP846sMv1fsYumkVgrvwPeqUlhS/L5bKiQlbsa+7LiQ
L5wCYOpgJlaJBQehA1WLClxDPM9ejHV0RPplpqwzJEkdnMSENvqgwlbEdjLMlmlg
/4FV9WAUpTOo0Ph2v5F0bqL0sU05OzhTbTS8VrErn4o0lJ49aa+hITLCzjsGx31G
t7vSoBvwvKrxm7afh6k84U3R0sT9pdl7m+Wob9Z742KqfHkT8Xe4beH8dvY+a940
E4REs290VVHXa+7QVSCI5R3ZFjG+nh4S9kAYnHXHaPp+Ye0/Qv2TttpVLbjzr2MB
QVwsoZznpYp+dBoD9qZoEdYcuYGALG9/cR2+VdxWGuvG3sroD3Dm653J9+AqxLJk
mJtiudBabASCpPGsWh/Dr3raepds2xVSzxKGQWTbE5vj8uVJSKYC53JnttFergTu
hQjxHL1AYXvWLBDCZURruTv3npVChVo5bHjujcHBy1lhBEBa8BLzH6i8MQbZsI6k
feCSbRFzhLXTohp0dbgxh3X0Kz4XIHDXKXPJa1inzxuGP++lVioXUdFNAYjn51Rz
d+JZdDLqVqsbVVXltmTbWPxgV4pFxexvZGpAlgDtH/cjYePIGlw1dQlE0cErFjzK
Zdcrx1lKNUDPQjr1oUWwRotzrVl5wD5GYG4O0vn3xAyEU9m1rruMklt3CiXred4B
P196a8bkLeD6xaGEhrhNhxhaRWAi+pYeHjktQ4Bzl2yw7n6NeMZb0ldw73jv8lbt
9Obzb7Pv/my2VeLqAtILI9gyVbjSRkLpmYMO+Jdzres1Y3UkkqCLRMmSAkGQPD2S
jd3ahkb9d+nGVlHJr32YN71ulzIbCoWBQ7S5arBnqmlyps7ybZNVsSOOiDA/Ed8t
gFi9rmKzv0bEjbm0kIyiaL6tFOmfzIyNzI4HmpyG3O6adhNUUpit6QBvDZzx1h/k
ldmhfgSa3oT7nOlUTMtKmtaBgu9l2efrpiJ4zGWfgLlsLAED+QygoTpoFik/2WGQ
ttLb2etnLb2T764ofvjxJIUDFQ5wkPholh1yWuHbF1Kmvi6+2a1F1a4XRk4m/ZAy
YrIROZDNptM3takgi5I0dWQXpLHvAma7dJs6LDyNfoea+zJo+emFbvQIBXF9RK4y
BApIbZ4YTJuIGSdIz5nnjrmrgJqQxOsBE1LGpUxG0XLKsdZy1oYdiYQCQkCwbdkj
zBflFDLN6h0h5FAJmEgo0f4lV49uAUjl7+zQ/1HdOuG3biXZ7v0gC7eZ7EPK5vZr
+fIEbKlb3N9w80fLKoopFhnTuqYQ90OvzK0lPaKJ1s8k/EGfx9Na0LXz9RT/2uth
L8CMle8d6wfIGOz32KdAmbmp+QjvousxMl2Kjz8ZceTZ5I2DTRDa3LaPg/sQDsAJ
oNy8IkKlm0ZOv4sAFvgzrQiIxSIQ40TxzEBuLGGibpXjS1ogiG60WsI0ZY/wYDoM
243OvQizcMK72zvU2b70xxt189dyEDUqbJcFxLeXlsMfJTrllP6i3KPNkHrC5Ciw
tSxPO2NagaQzjJ3T3URX/L4sQyLzL3cx9AD4yguqUY8zOKERq0JnR3DdoXjWNlQk
MvudcsqtRBSDJ9b/O+HdZYB49u0ChLeqYm0HkcCNoUrwlJTAYyDQ13oBBgQykeSC
Zgj+LXU5wlW+mIqwTxxvvh7TpUEiyGxuO3H0+ySVe54BPxJSixiF3jQ5zhZJXGao
8hN60PK9+9gCsKq17BToIZorGy2+V4+B7W2HPcEqBg0Tf+VBonQYbmlM2Nmoim5R
9kk7Rn1JjGw1VJNghXRbBz7k3Q6JV0+zt88qIfeWag6KSN4cyDuV5IaaLzCQczbx
hWgvw4cwhk8Rp8pjAsFw9JC4bouKy24xiVy9spI05OO6GESf8WpL5jy7eApaelsl
7+Sn6E0F11qduUz4nXDpBue3Obzxj2Rp++kWxDPgTF77GQjmvzKLtRUb0Whozkp0
gCTIVEb+v3nKW9bICZruprJO7OATvTYpM+tO48SyYghsvYRQMX2LQsleHbJmheUP
ztOiZPyClNGabLAwWewMoX++d5ehGnUlTKPIJsoE7PCuO49LnJeJBXGgKeTu6xNx
mmA9rE+5mghWyW3mciGSXkBAaxn9z4qqKECyCZwxser5unjTY7Ehp+A4GS+2z+vH
0WeuwWwMydTEvq+zPKtGB7qHWDRSBNNHoG1ClQOVOYreyLWSpeMP6SyL423IMOH/
+C9UIy0lzsxFg87Q+FwHgdaMJsXeenp1OGILqmnFul2ORFqbpnL+DIbWod60y9pn
exI8hmRtMb7xVQ03cULuobz6yXmQ44jhu1TZeMdvLWNW5zG+9/zW4YIzTQ7j58R6
Ps1s2ECuN6p3oQn/1+a7/4NNKTnzjdrG6JC7uowWJVFY09CSnMvqXpLG162MVGuc
1didJura7AyI1rnelNtQSymDUYO9Ip9JDCyKyPa1vNPP6FlgmkOI3u+XrXX1JqIw
/dvFCuX4LhW97iCn5HdkFQII3NbSBCauQt1ysjO7iS1Fpsn1Evislf01ckK9qjlj
ZBBVTRisruYPrajYjk7v2hXFAuJcQSNv3ReCcsGmQ5sfYYUCkYXV7B6FlT2RoiC9
n10pWx91zWCRbu64u0xxqwvjuvrn/4raFqHFsPjmx6ykgBEnPDhdJyeTBTAxZB38
MbCa92uZVTqQL6JtnQArnNktf9xGroywQlIwxqIkerY2FAflyShPDC8i46g8g13D
cRwtBFiCMWhC6yKakmRMqcZ8er78VUdmcWdV7EJvdoiqNmmgrvTqcdms0wDYFjI8
riwdZ5xjQoZ5J8L4rxxlKD3uBHTEAYm9wEj7GSNB2Q7hPF072z7OOGa3TlN/fhUs
HJMHRP1g1h+/V2tjHyrpQZj7x2/sSJAcC7n1jQeAe0AYflrCO45gvk2GJaPYKHSz
GH7YTjB6JlHIz2XAj2vmXr2LEODQJ5wfSugRWN9wufP6JWAIuhk2CLSlqSm2mnD9
UsYUScxjxRtEFOBjuGugsNPqa508duO8mXfpoCjIo7REEEUHnM6drxYODZfgLHFp
52JDwE0hF5jGUuDoPiEhnKpEeKxZx2t8Ieimwve7NbbKTaoiJDz75GdNoVUVdkPS
jqd0TbzOq2vrc/OL5yjsNc3XVHTr3chmv+V/tvkm/bWspmx5O1owp7GcR0eqPwoy
/za5TKVG0yCSTZuwkJp1wW3gmz2scguCCulCftGaTTy8bPsD0voRyHW51FDUlQIL
2vPwz1UoPjDT8WdXlEtiXGGq5/5JvCV3uk0cs7uie+UCYeDmINhutPW4ijZyhrHs
Ba8fK1IpBhZIkcfvvlQv573FDPtOk2GwYhmZgL3NTb+XyZQh4qfiqGS1LBgpALdn
a5p4jnx+dOLgDWwysWWir5qotOZrSfDNTzmd/jPkUJhHI2RcNlpdqAJn7HFf/aok
bPTcyJiMlohfnv0GByIU8Q7uO7VDYRI5DIg7U5KI9EEfosz/2GTN8swaotG57pS8
3EpqmEFF3/233/YEtk3JD1X/oL3I41s6fIQZMbsCd8WEAIo2kdjNLzqVTUz3cIu8
U5poN8HQcxx7UBbLVBdCHpabwKgw3zZ1dLLw1Y25HypwDeIYe9fNdkyUEggpsLTo
t016KtMrebxD3cZyB8NU5SWWwnZoqVmlkrBooNWC38pNXj3DKxlZ34U2XBJVu2xB
zDnxdbPe2/qUv7QhhfyksoBZhJfM57aVR48CgjtbU8UGYW0DSAhZMDWPPdtlCJJg
cT2B1zGYxIe+hxk9AqzqNQmdeu+o1y9lVMci9a/7o8gl78VPkQiLw1b3tXLNu/xT
aCclLnN9AhrLiDGMt5qgT5ADVlQpyS0bx5CRZ8dcbTlWIzP33iwiSbAnzKZ0QlUS
0VSm9imuCE+zoBs0Zx95I483OwGRlOg7dYvON3jF2SqsIxy6rBS3TAx02Hf9sYt6
xXwLTqbDkOQF1Z3lcbws6jgxXjcErDnONdNC7ARHSH654PNC6X1RvmHfSyxbMMoK
hBE1zH9RKd1s5NGD13klNt8Ew2wEZ/pQaR1r6F+NwhQ5FQofYJ09vrlsddvxWQRU
WUkyNNeP0N35Zmn8Bhy++96VnlFXDAim9x2M4VfAfFBSxtj5y5S85EqAr+malECS
hWf+9w7JUZsjP0LHFmL43+miezR453n4XCIZwDmiXKKe9ZOITFD9FQmFV4d4dnC6
wzFKSKmU56bFBiRtL3+2bvG6qywDmtliLQoeva632n70QcH+24qft2JHeMBZFyI4
lQmdz38FAgcvRZO7vPnZpdnoC3uGkyVYeNoqC/HDXeBAovQsdQnh19S/PuQAgqQ9
hhUqLsL/TkwgZmWodFvl3IZkx+fPELJUp8vBtXu/etbDkP3Nn9pFx7HTbmA5H3xq
RXOJgne3DjQWGprFD5R5SqcWujbahW4RXk7guyj3xMistgOJgT2ls7zodewL9x08
b3GaopbCP4ThaNkJgw+96mE036DX2NL+wZ/Gwi4yKlMS+tCMV8ZiDhVPGzJEC8YR
fonmD7r5wa+HVQ9apBq8C/po6yijPnWdaFjV8yfRSYntZ0gTw8xolqxmeJmy8SV8
OB0D9eQ+sZPNyYTphNFvYm1yA7/7eNEV5pm9MdDETu1a1TtNacY6dW8etEh13Nwe
G9883BPbiMeLrQ/SMXJWCz3c60lb83zoIMaa2HBoL0kxrw57t+e+FLsjLBmMsL1s
dHkQbn6A/YzpI1SL2H82SfZjQ/xM5Pw1XR8t947kWI1RwTsKZ81THWsH7b+OUD8y
TpgP5iNsn+RoFc/3J1T/esbOdqZ9lKS14yWqiKlDJPBkLgt27PaY79ddR1N5luPb
4W61Y/2CvQBV+D4/KckAIWR2QMY+jme1qyCVfSkNeZfD1uaKj8Ayn4bnpV3bTXlV
WK0RvyVovZSfH1JRGuaseg7yRZ1cerF5ElqThBo/GW46gDdwSRZlGpysrwosiTd8
t3Q7iyAwsH7OkTNB8Gj1nMoEUSliMDSf6+YwQzzUsxQiuGzpSjTGdH+Lz6+ep2q2
s384j2R1D97TyUuvsoeQqMrPUdE+vyceeeXVD+bhci242p2DrgotoHSw9W2tQDY+
eU2+eujIy8KxrRjbtLUiI9scxUqcnfq/HUzLRm8I6QkLc4/VIdkgU0Fst9DUa3wD
cwIlt3MpUoUXl5hrPswGnXc/qXhC1bHQ9rn1Dt/g27MprFAju5fKvpPCVBkBXx8i
8AGzCUH83Z0qjfkO/EkhG+nQq82ueiTY09zyIUlkq/QewmlgkdmvaHfbMy6tKA1w
AgNz3hIVk8M/mUZEIiDBYMDmiRKi5CgogbivI0Zly0f9lHnVck+fwAWFAOd4MVU9
rddBol/C/Ja9+YtkyO1EWJZNBN/D3mS81pl7egWdq5c/DG3T8c+D1Fh74KYfhIlU
IzlIAz06F2Z0MI7DvJnHJs+RP9iZ+Pz9Xdl1HwBKDPFPVM7vPgWtKrP06a1/r63d
4lcsTURHGshKNM/M3pNAsQqPf857Pb0ZtVccLx1mo7pmxlU5YXDLjR1F4HEAaEv0
hMNGG9DhJzVIp5B8XRjv0ppxQy+NOqwbh0Ykpa3Dz7+f7TopE5CEA9xCd3LrKlUc
hFHJGgl4t9Zr02S8bhLDKe6b0IKFCU4+/2+fkIMPwpIBpVXh9LeREkQlfR+CuBl6
aW02d/NOcBL7SoiYv70PnhKEfmLbw4rpGiq67QpzclDP8Sb58Q/a01SQ3lps0VHI
Ut9Vfugbo7GTPvp3L2B2jeyOmO3FyvOKomUOHk9fw6L7TDm+ku0o11nCG3vgSpu0
wuhREP2NUKE9SMUAt6JZzlwxMb8h0gSxZRrFovQ8cSnXtXUXifOctCVMcQt7SDvC
KhP6GYmFhcG6vcqpJDNp+42cq0J7CgOAARey+3KM/8vxWyL4FB4JGClumdj62hHr
c+tEXGhUhwQdReND2uJV92O4xgG+kIWWfFZL2WBnxkETMYLz39K3JNY2R8EERyWD
+u4NYgeXKUutusGe21698yIik5IXhgk2RvNhzva5jbRp4xoRGP9E0eyuZW2fS/86
+SPnySWqZyQXh2TfrEOLwBAQilOChhZZPoOxKnMnt0YN+Z8gQiD+gVFssHwUgV/A
a+bink2dubacaaME99glckjYjdUhYdoMhm0B6pM6IQiuj1bXeRi04v1ozgWfj2PF
R8lugohiQgZxXc+S+rRI3SxLYv6VWPRns42hqD4dyqUd1c3MoF5wJppSzfzT9oki
xBSU3nn+tFPfSI1/xFgbgrSimqNC8ZVUNBJ598BSv6fYsVDJsSRl3Xe8ZpIrNaTl
yxMuNKHWevcKKi8QXv6ZNK4hDOxB9aBmQHbjoGGEWwL7buURXCIkiF9jH6gk5LRW
WClK4eIoVoZuig/MY0e7IPsJY87Xu4np8OuABLyVu9vSzQjyu8RUkeSEzFhOH+0r
SqW+OQTbKht3e/x9l/O7lyW+3O0A1BoHWJITOKXwUnwLPIkM6Mj1xSQ+vKnUYylD
EKQUeUMyiOOC0Y4sc+M9XkBixp3h9HpTRfBrgktyuDCgr06mg/QbANNs/7zBpXSb
hWf14n1kfRogdi+6wc2YFZAeaypi/j9jwRNHdjrkaPehT71zHmntDqI0LT3IINYE
XpfmNmNrOQRGDIaR5LIe/H5brSol1vSt0r0oZY3OHW7DkbWV+7z2OqMSNRNAtcKn
cQlzhZv6Q7FPMRktljs5Bbdgsxyoui1jhrbPFQGSsfjXTZ40BubQ3g+V3oEFbLS3
HOIhTHoqTfVq/6XDZRnD1aZnMqFLH1k7pOtgu0JRhZPftaGYBEqjuw9/fvrhRco4
eIO9+lH1tmpPlfb7jAhtLfinUMhhLwNIv8Wg+IuuSDrmHFYcyOnqmNaflXXJ9DkL
JU+Kr70OM2PiYwfmRplcnaAF4ip3eGWRmLzLkhF2HXNYmlDRr7N8FIzQwXkbKvj/
t4xuNzhBw0Bwwg4lY7e3lf3xSKYzDfZbo0XVEMh8RXEBoFnsSK88COJflcz9S0qm
YydNxsckNHSSvjD/i2oLx8MbccwKzAwMgJ5oP8c2rUh8/69L6rYhRwCI/vdkq+AM
4394nP3pfGm9pXrSqH35NUYPsMc/WYIVkp/EKsCMf7CDOGpjnl64y9OoF1b6P72d
SgyWDiyPudItkG8eVfI8IiADH/XKDafTU/MJZC4eV1fh5l6T2Kh6zywN5W9tIQ3i
G0xCA4Ljr5L//8uyTEyr1m3Ybo7aw8jkDEP2DfhFKAtLhDNan3Gb7WI082TXGHpb
3xGtxsteEapwOBrYYTi1lFn8/W8YHedjUvq25xGvSVxMkqrA0XadHfIgfZkQzcp+
WR1CEF9ZQqxVvtBOXmWCAW6BvOo5m3jl+WcmFJ12/sex3i8A+pDPHhqpu7YngFL+
jpD42+/+/L+6IltuZODFBsqcRXH5bIAvet3Xi7ZTxZ9m0Ot63SK8jq+t2iKZR4m8
MMd/gal/ADhsyakNn8GvVauHWhRVCN5cMyXdUVdj4Ox//R11iHWsQcMqQAfw7Oq8
0btgvTPJJIEjO8x+W+Q8PCAWKFnjhc5HqqN3yhADtrUQ2XPvNBsm4xMjgyvp3S2q
AywpmSdUAHDsAbA+8xAhd4LQgMdVL4GFhRVtwLdhpegqtjktci0MiH/Xyg2j5wkV
DYKnag3R7Yn3/gK/QQo0uTO5bT9qwtJOxgnRsd1bYEypnXoFfADRmpvNP+r6UHOs
s4/uhGTHaltYZuXIBxdUvY8AWjuyIwc57yX2/QEDdkQI5fGZ1IsMR0UR7JlfrC20
a/ew8A8ooQUTlJH+NXRAKwZlGdT5gSDJcCCwYxOv0H490mESjQjfuzSteThKz1HN
prtQFaILg6k1+N4cl6pBt7i2PxDPS+o1ygMb9/K/TP1TJWw3lgX/3THfMt/Bp/0S
7AfxLSe2IwLSk1nsvSET5TOcs8BDBpHmHPJaEeTTXqoDGr62wOS49q8p8FDHTGjZ
miYe6Nk9l4/qTqfQeL2A0P7mtkLaHl6HysXnb2108kw310bIlx/Ol3RmWJvLfSnA
ahbeqZNkXSIkN1+hzyELMxrv1kGDlJxwihLNgzlo6MvIwcCe3ePNfkbISHxIcdY+
hxJaL0J+tP5uyVJP3cDDI3zAkc6nCvR2rOWvjjvgeckuQelewfNNbBtl6l7+ewBZ
Y8ceis1DEqpg0dpPVu2o0NZj4Ioo7m1U6a2Bhx3uEPH9knzkcdpRUNYECkpSJDJu
UYXywye5uWc24iIC5ZdWnBtS1BjnfqRspRd0lwpOF/N5HhSYSqFls9hD039F8zEt
d663aM8sOr3YYSP+pKsQ3bePk+AJ6qfkmvOlEo2rxUQ+CSuyKEC/z+LK4eQkAfO+
fKQ5Uc3XvPvcIV3Gx+BI/10MoSUMyxkDp4rm1wtF/P163vZfLBdBTuMrSnFLXeic
srq5Aj6S6KoRZzBtX+ueYQ4WNDMxm/uHAOoF8C2TpH5jWjFr0PIP6afApfIzKXFP
I6M+DR2KhR8rVxwjXmeWADVHzV0f6o0/ce/DpDVIK07srAJPdteT5ZHIrSDsmV08
//iWJhL47GoIaUmcZOlOvXqrZiBMGRYX03DkdJHNYG5Ng1m4ZnsBjJw59F+oxY5s
y6Wgc7eKGzqcc+HqXnoO6w5Ku20fcGHl7rivpDSqi4YHF15cXOdHhhzP7MTgieu/
x77UM3aSx/WN2aMpOPArEAvtvDeykOKMqifDgQl08zmfIuPSeRoJmVmOIrzFutgc
bK2ANzmM3TDSd2yX8u8E6kh0XQQumRdeeabiJINYbEdOj7NxqwMlv1KD2/MSQCDz
I2euSyVShPCosE4Tn5hPeN5ZlLUUFaFf+BiEwfPeTpc+uRw7ep6k9rnjItlqEZcA
18Q+pB+AxCd0VGIQBT/FHZuoiGQClzfP6DzQTTK3BCZF+T5hWFcFwCYS5KfPYbZW
qjk+bulAm/lleIJI9GM0zbPpfnUC8kq3BOWKSDlm25uLaLidk0lo+xBDmpo+pvhO
DHAkLBu0USZb9AlNGAL0ScOCL2CtHgrViOSjdXncAS8WZeiqwjbyZ7hZxUp9KYdr
WpVyr12lFbnv2LJBaEJMeCOyeR1NZpiidQLPZgmsZC1urAN7p579hLZErcPr+m5C
K+4vK1oybhVuXzsbw62MKtO1tY+mDO+H+h8KxsFzixw6IikrTQ5oTBwN22Shs4Ty
virxhhnsGGGOISk84FchTdqSYdRnmTGAXQ0376WQHZ+eRjlApfoCYoqT+r8U6JOc
j6zQZqIFvtAi1rkokZIbrKj4aH/VmiZSnmBbVek0+3Ax3KtIaMI83DhQIXsXMi/L
AHASMrmyHKW3gu4Ovi1XLLFmk1Q+3NiHMbRG03TlpuxRjP2IZwRY3Fsh0rLppEIj
ftOLsS5XveN7CcVbWcWzHfoiNTsJB6HdSA3yjs2B5wN6nMDfDBPGm3f5h0iwUFFf
MxGeBss8uVUU02SCerdzcPS1/3S9Xrg+hnRVDTLWZoJGEyIB561JdunSxuHCtYZw
m5cmj1/iR2fx0AuGwA11P7Vf0zxU+7zPTzb9BGBspTutFkt1rma46Ios0LysRLML
2t9PEY/hhiXy6vf8AGrpdmO/2ISz11BV8L3INNUCYbhkXCg0Ex06CFtNyxU5CbX8
TUNks4q4EdBsjuVSnIwSze+qJMHo9MqhUCM06aT38AFEf6Ydgygc1JYLytMTRxQE
RvX2LA6bRrFXWdrcL+yPa71C4708RmS2L6riuKWvLnS9ONBY76f0USW0dfUhOzNx
5buI1sSlSsyubx469Y5meOycMIjYlnl5xk3KT7AdqN/y3JZQBR4cIyth6k9NvcTq
PYQRd7yAgdg2uI6RtEzOhANy65rxJE0Pz3SlGEN/BXbx+SGyg1J9UodBCU47rTNR
rfNlJ6My5457WMz4ASzlRpR1DGawITS7DtxMoMJj4eav517IOKGwsXnBIgdu18QK
nWndrV+2YJ+O/SjFhAUT0i+VEMie9p35KjdT0F6OXlrbZJgdj4Jd7baIb+02korc
0gLjef0EvG7TYDG130RLcreT4PhVbcu8uY3WXH3o26sLzQPadbahIy3GAlH20IrW
Y6YmldaisxGvJ8H4h2PTVTbHsQpX4eHKl0zTS3SZWOeBEwTeCU0+djJ1b+Nz7cvA
P2zo2E5JtUp3fEJTMYAdHxrAIlgO94OSwGkpQk24TDfIqA5MTXt7fxnodpQfH7Pj
hZ8XvMARVX2FRThLtqBuayxwnROfyqxE+gNLrp6OKNnaJuITn/clCswdlK9UyBYC
5n7xEkqUAQJxzkzHspKmcdFvy/PPDYq6TgO2q6VVHdkLDL+DOxF0h5Bh/9SVf9aB
4NLj7VDxo9MGSAl/F4f3iOHOPi5/n/lefnUkICrf78F68Ek8S5McwwdovgrVmVlZ
NaZIgWOSBfuMzIvjr7phno+HCG0SP0KkyoaNxe0qAXeNvj1oSH3oQvg0iOhIqDnc
qYAK85WYbdsA4feQXl6Ss/nDit+MnlmBeA/67hGCcdexHTdiCA8zV7krroWgNOba
X2oNJMvkPyL4UCSFCX4oRAhWRQbGs4xedQkKpx2baOV6i3Gsps80MV2k/Jxtzici
H2btqe0DcG9is1KmiIEDd+LgLHODaTjJRgWJ0Zi/5WmwdCK9zcf77TP7wWGnPGGZ
QfQ8jOqC9ANbLNUfoHtoXMwW2i+CCo02lFxAB4II43E9rVn4w1xxCDK/XVurdmSJ
77xSOx9n0fQzOCfskRWs22CHCZsufDsLSJVjlH7HG6paJ7bKlaXvdBCSlg5hy+wS
hVRG2CggDq8Zvu0G2joY398s8aPB72BoCmHXLN1s9XZd4TMmoi8t0gVKK5r6j32c
MHCgsx+J18sASl/UD1Ztqt/Rnq/vN8n89NqiU80Qps1rUfp4hi5bU+AihJ2Ll+p+
BwFq1mo73JG3iM/HdS2c2Fqhb7iafdcimBqE93DZrEAUVaqAptb2JqPAagpjT78C
mFOSKYom5UzLP5giC/UbqUUnc3+lUD+OrtLjLU02NuU8uA/WESSApSwPnQaSGpDf
YtoHgMdZjzsGLpX8qqXrnVLMAxaOsBAJstzaoTLAT01heM/E9+REv3aHHNX3wrtz
9CIjChVgZAassDPo+cM4jMOrf7E+v2JILWCOd5h/HGztanZLWCRcQJFTjxilLJZH
8Hr1eYNJOx1j7dKRGLe6La/xTsgB6V5Yg8MpZmJChIqX5PGtidr6RLKRkXjUGj36
Qlpx225TBkoCiVkZWs2RJZNwSzlsWnoh155ZU9aH9PcaFUzKoR9qwizmf5tGja9w
ofPmkOsI/jQBtcD49eW6T+2XncxDhTJUULhbm3K7NQI4aKjUuOD8qGtQIbD7sLkW
BU3IN95SpF+muLBGkzkrRIVMSYJcDE8ZsnBygYlHvbjWUCtS1eIBkrB5+buLD9wn
Z4FVqol5B4W/Vj9gmaUL2HpVGiRRDqEQ0mtVu/Q5144P1xqYNwjwUtgjq3YNkfCZ
D8/QBC7Cf0MKW9XM+M9rb6V7sDM/c7eSs+YpKjbH2SjVfY2JdbbeOUceWCimnHtZ
3QCyEZvZy0LiBUTmOyfywwDiJeWHXs6tmNke/4q9rL1XgRjcIv4ZMU9KnGZrJMyr
O/gVrq/YeRAo33b0i0Wd2QkfViIHCpeSYL1hedfEoPH+lvB8H35Q2O6JvSYN9Z8X
tCr+QxCyC6Q1C/8u4RDzJ+XyRBlDrrqWtG7vOo2BI/vPsZGl6XGiVOGgfunB/iAL
xu8LY0PpWO7Ix2+j9ZkP5u3hOPQqN7IeKCJW7hT0DUYq7paFG0biX7ciAU/zN1JA
LNvyUVFwLHxQP2wjsQ4JKqfqIc+7t2R1A7YO9jC/uHCYtcxmVQonFHIDETBkSCoA
UmrGlfyjix9IAvWCQlz6d+Bq5/pz61F6S2B4NiVcExyE8XKvDl3acQLVK4OCTBwf
RJ/Ccw2HlgpgFZVSGZCMMuzk5x1f/IgotJQ9OzQwa9qvGFgAfsReUojCSRXhio+h
BDDt8tfLcP35Uc23AuOJMSebYZEluf9AbkCLYXYhYZqu/CCBZlzrlQonAQhUYZsm
WPPbcnyfMox3pKjEbWhZOUscnHOk49KpHTyfsXjt0KgfJOWmtOcn5ytDyKy45ffP
q1jVCehvc9d7OAIefzKWx9GTbN+PnHt4pBEgilpToFvxYr0n3zdyXlXMiVn9IZ75
AJlI7ETiN7d7jFytAW4BV1P1i9NgDM/smf93ZUrEKalad7sSgpptLBOmBopaYtj0
u3ZcKbFfxuhHO6mg9BzVliBPRWcPRTI2m3NZezOzN1sfaWKbx916RVpZe7DYmdP0
iTDX7vNvkksg7MzveKEnLQVlU9tQ6oHnmvKp8GJxNOfnFOiBq37O2C4tvk7OXIe8
lmyDs9+H1xLeTIFuigpWsZjOFwEVeZXJQJT7f6ESSZS1YPCfC2V4wCu4wwfctLrb
XFsXJMxJEX8pGOXObCczCbPWTvweRqlMQoiOd4N6QkrnvoOvg5avWzvob5sjKZ+x
GrR6dAbLpwZgzE+LahZOs3/hWJjcUTRiWhomuTTSgOJWp8vLL+YafxMEq2Jp3uLO
JY4DW9xLE/f4aQuSeCLqGvNxNfx8m+a14Kd0yrXhfWKtOn+NyyFrPpxFo38S26gn
vrjdMtUPxYnwak8fniWhSzry8cEm/k0bMt2aIOmN/xHYovUGRxSWLloQPxH61GSG
CG44vCH48YPhvd7JgAAOg/1izvypgLJ64DWLsrB/ub3fq8uHa5gky0OSf1z7vSMg
S+d6/1UcCmSn9tpsawDC5so6ZVN6xjA57Ed2WL/FLtWMoARsMOZn8ZBo+2wvhxyw
D40LVW0oIZvy3UgeN2sIYeB3Zpo1hn1ecR81oyy7Bq1KG1yGhS3Tok1j2gMorp4h
E8Gz4UJXu4HQUpwTxivl6CSHL/Le0e4q7FukELu7D1Am6X6RY7Z2TyvZMJY7ZfW0
JrBWJdYz93vKUYFDi3KIdnlLG6Jfbs9A0j82Vmtq18wNmiMYVfXDF+pkaAI9duCF
oXpsKjcu5PoaIlQ0L7RABYDLh4PbiaHgM8cicdvQZZ1W6Y2wp9kIthMv301QZmKE
/ufQ4MD/htlvSlyfzEvkiQKh0y2vEqDCra2WM19b5L5wK9nEAHrCrXIMuOHLyBHv
z1MLg0ZtPdQ1AElHOfwO1dmsHrs00vlbnJja3ols3Bkn6DdfEaYgc2xdF9/XfqX+
OHOBICuJrJGFxM1KLbGSDLqzL4XfZF8dL8jYjZtZpagdeCWRAl1eE0ZbOhJ38aB2
AhwWNcq/zwhlUzFNd/nSwuQJlgVfMdToLR99NF2ZeqE9WS/OoLHKy/bv+vSk5cTa
CGa6Y5L1Q3q3WzKAZdpabmuBfGGjKsjWh+XgvD9T9WiA1xK5FZr+dhP938N5TCPD
t+Jk9rJHHQIY9tAdzBcS3HMfU7jHjqfNchJ+AYEYF4UldedL0dBCcQC3neHc21oA
z3WyPQ3rL8PAypXd21nl7KluijVXspAfziMzjtl5W9tbfkMqbcSa8nJRvVZxQ7hF
2MFMusZllnfqopL8Y91SjZS3MQzehR3HZbwcVtxeFKIuR9bfYf2TiMMa3gGkD2ou
fPBiN0Zlo40Il3zkIkvcckWSar6zpmymWvJ0b63fuhodlV2K+jtSfoviIhEgf4T1
ZJRtpnNpDKpUUYwxCIkQgAHyTUVyA+Urj2RhOPWM+odlMUsU+7g1VORi7hmkf3hx
n+fYjGvYinktTeZVkF+VFpOJq9/X5JSEyaRyIIXtoAIgBcLTUV80sBiV8CnU07Yg
a2KHux4XXgXxuaAsh4fYo/g807zdc2yNyowz4HfKZnP1E20A9eW6ySxmSqNAyT2Y
N4wxSOEC2Y9WLk4+yvJlTIT0UmNRlWqZDFt0PfFhzIbTGADR45FNh+U6l3L0X7eH
MQAo54wJCglWyBteCn0/bpIOMZDFaGS2WQsSv8k63ycaXKcgt2E9yn7A/2ZyKUu9
DWX8FiUZdwUnDQeaDXzlR4Bl61rUuLd35168u3YrIEdkuPKBn81BQVVNh0YZj5y8
XEU7RZHcDHGpTue5hj6yPr1h/kkWVtd25AEUbimvd5cPhEdbQx1stiA7SR8BPu1Z
YbsIZTWo8NPV/ch5i90usaPjI79xaCVpXGD1r/Ijj7/ek2dZtJH2mBR0hX5c0nXk
JVvOgAnfdnV1dPXP7bHASQrskmtTkQx+Pq4z0gGWsghVTIJUcRNF4+9HcyusYmyG
q5L54kVag/rGcveVbJ8N0FPydwmYY9egTm6u6t2h0KrmCFwzT+MH1+D/fQZXaY81
hhi1Zf5nK4/7KxbhkEbBKRE8/zLOqZrWJlDjhOD41ZSBOR1V3qASbGtLF6W0dmwn
7X8BftJXvin25c9TU8zmFCSlHZiSYJa/1Zp+T8ZByjRj9w+mPdzZ3ed2KYJwPKBg
nf25mwGdg8MaRTgQX8bcC8NQZoyUPkfKo/ZfH66Cfyr/zYb/8lxZ6DMpZ0kOkjxc
fJ5s22mibFuMSmxhT05RN1dYilany56luefAYYpChRbfBWgYmM+bmSF9v8pRfJjJ
V0QqQXm6S4z2ZKI/6HkBoXI8oVM0AbyidGp68EA/lvstmMUy9xgdmsJBNSneaTf9
1UPYunciFHkL8V2w7tIbQUZeRyMWN0hvZfg78ahfY2Fp57/3aWrvUM5g7dNostw6
7ihIMhnbkVcs9bWBOxhk848sLQYqZGTTMZcVOoI/oFCMXtcH0dK4kunPyQbbwSqj
G46a+MDjN1bdmUYk6rds56F0e4hn4kV7apZHc/j2c0Zp48mqkIiFS2f92nmhv0sN
4BH6fSJm5ZIPuwLeznKu0E1ew0vTQ2RkgfU3X0Oyd5c2gOYXcYHXs1CKwpi95GQA
xAfCrxuRje9202d9ZXNYzFnF4KWQSvkvdX8aKdntiaFo5eYeMaDRHty5VRDoAOCa
pa4fnPKTnpql1T0mUGi8JaqqR0GVeoa1Y81npWUvqyRA6sN7gc0nlIwJu1y6x3NA
m/essb2BoOEC2eBEczZD56QLjQAvAen2xCcsrsj9jP4tBPxWDaR9eQ1qE29mXX+G
4SaIfyk1SrmVTOAV4c6h7+K8xbtgoAdSfSxTUdBreOFi3CGX7RXDBFcQ1QTG5Ic6
vwt3ZFAUJBZyDB3tET6K5swiLw+8xWr5L8eLdwnPzdJKEPFa2KTy5fH+Gu93jVtl
6Rit/Bs9e1Lj7lIta0Jdsix+rUebErFq1As/WGIw9lrtufaRZw360RKmxDQhtUoA
MSCjcK67uGzXyesIXRdFWpaGVXuKgaO3jM6OfCKcp5kXEbFziUByUmkMYKqItxgQ
dAYnf4JORY07+UquQ4QEC/C3EshAQ11rMiu/VyOIuw1SFrk7CdnLWlVM6h2+EOnk
dF+qgDdmPHFH+TNYPrdhuPjKsv+1eZk0rZXgPqUl2ARKztPR34SbRbe9HKLrdenC
/22P0nz0mimswXz4d0rBiIXWGYGq+B13S2Su7O5mgnM7EnUIOvJdEDZLwcNxxeWP
ws2kENn2hmTe0USLaaLfa/C10ViiyZKtrJwKkC8Sdv+FI6TnJ+N0V6ILU40eKChC
Yu+BHrf8igzvtnIli/XjbJvnZ6W4NKgCEr9UMjJR5TVcm8YaDRkrRYpgOxFpA4Lj
CQvvbhz3FaIFHmm7QD50dcPBKEz5nW9SZllSZFrZN/36Qbaoi1TCIw6tPFjMR4wZ
Vtvbuj2EzjR+NZFWnVQH/lWJX1gIpAhVCGKfDS4elOU1x7pd4CjaETYUpjM/lNqq
+yek0VzFkUme2fgkTe1LudV+KE+TmZJ5chPZlmgKgtBZXuvxKhvfdPUvxJp3cjdl
PGgjBNnpgVhe0x9oBMd35O43qpNm7yWJlaJKMo9ZJN3DEzuCKb93/W4fFxYRUrGd
vneXRmv79GM3+5OetH5iiFhIBeovPZcxdWf7uZe8m33VmQGF6JF8lQuW526HhkWC
ffxgVWjZ/CdcjgY9B6NVgJ4EwEraxgBAt4BY3oxgeursnJlKoK3YQurzVk/5Yiu2
GqE5pYJ0SKj46I/sYtD0gTYiTWry3WhnQi8SdhIxN+0jJIdLikJqIJoeOqdQEfeN
Kdj5c5SVtu81rTNfFcn+3ouMCQq4uSFzaZO2os529NdFQWmO/XBYFbG69KOT2JcF
88F3H0oiog7BH8HTlVXOOXzs8RZbnyJAsHj/DdMAsq9hbiqcOTmcuiHiSAb8nWSK
iAwY9/XYQKPbSz1cJ1IftXkJtLrC/pmV3DeHYTl0S2wx9gduZxQXIBL9ztyTOuA+
Mc5zofPQprxaK3jqG2U2gxe1Bt5/xtriTiRGM7cXDzimdfcUbuUXE2qE7jWvRm01
AcuCGBTjZCat/wp+k6RqCForgZTehenj8lYfEq7ICxdH8aqyO8nmc0b6FxBjvsjv
W5dbU25ChtzV0glbL7dnsJfvdJAhUcB3yELWqqUhth6RXtqXW8vh/2wZmfo/d8LK
GyK2vZ7y9blh7JAXkGITgipVX3HwVzIO2mT+oZEMcTz4B7O9ht5h43fph61b2KZT
Q/FGhGyXY40ZLSQvaXwcGCKVkC4tMWbsTgfwBTQ8r0Jk845nBz31/8RQcP+RHGTk
3PQTnZ/A49TOFwBLsM/erXRoPxxa+Fx7vUFUPqe65TpRfHEHVvpd4ou0jy/FgBkG
Z2Fj1un6Mn/3AWNEbtJ/vELuBMtxJ/SbEso+uCiVEZu2L9q5YImXq7JziQ18Q/Om
ECh0e5lJJtl0DOMiI0ClfcCbNEaCvlwcUeeBZdy1TKzgkktnwYFujOn4YVcOFQWb
y3pasbctjigciv4PyRFSEGXlNJf3xCW4ymHoEibY7FpSUohBLs7SvMeGfcUxoSfr
R83TBuHB7ibk+4ta2Hsiu5Vq3Qk6ijgkGeV+jFrnn6wU2ULqElRb9E7iO+VutcZE
dCMaf4z2mFt42GxJMmXxkNoSc0Z9vFqMPjDWaCqBEx6AE6ahBhHx3/beJ+onJewy
VBJnHNDMTL0QBGOvy+sgthd3TeaSPf8X7nfwVsg1EdUvfSBfiQX7ZaU4Hw4PLnpG
9KfwsP80FdYkdo/0P7zuMcYd9TgceiwzPyNAhGb8MfSlUxxlhthipCiOTYiopumA
K7eWaSTJL67YqN3LqjYABwpGJ4tHwWWYPLuDSZAivWJp8y5tjyonrGhf8JqBjySo
Yd4ymKz3DtKStAPKiSFW2o0caq9yZiaMhiqI56FaPS9XgSW3Ky01u+e1Z2R4QEgV
W0dZkNY/92Xnm+GJhyOOmbE2WOhf9oXe4YrrImGwICMloeujHC/yhppegFoXj6C/
JVFVadi+iHfZqZX7kQArFugxQHTfWmvtJrPUrcIWCisPeG9AyVZvXbMgVK71UTaf
9lJfa+a/QuUa2H0uQGnA4Ds+qNhKyYNFeayjkc19H2yQbkjfbLZmgZL6aR9NF8a9
4gTLufmuMGRnJ42cwvZpZbxGU87GGzVUgDcWf+DuXYP6VkBzKPERZII+uO2mjGWC
0gwXanthny34RlrBTpJvnsUMaasLMMlcpXb3B5ktQMB3M+vzrQXuYAYNVWoy8aH+
yLEwxoCRLt+IkkcUcQsKekn4Frn7XPMjG/nXB3dD7AFfCq8JN6lKguU7tw3ODZ6u
AuYS8eTrKo0k11NjBS+F2cCKSkcHn3E00NAK8zIgHBN7DUhn1J54xG9ULycp7KZd
QG60o6vYqw3vQJGHaMy9RslBEItsEyx80Kb4MXOqFnVUu8XTkcSyttyXXmA2xKp3
gydmxWPzIExFK1D/6MLIUqIGDZBH38hdv1heZOoVcZ9GgAX+joNiZc7s9dXhIYKZ
hS4kFKtRXGGnwoaroVALbFsARYhdqJz8J6ehKcQ2fKUc1zvQaBnNTSnO7IodoeFR
iA2eA8uVXFTyM3Oj9+U9TiI+3ghlDobaNBInt6044blBsuI5sWVkT08SZxh/db1B
dccPnb8hFVI2s+Ox+OzzX8HtydMb3iRr4Wdc8Lq9bxtmdgezuhW6OMbsOQbjzPBl
XB/aIshGn2eQBZSl/zUZqOV4Rwu5YjFOTUXzu8vOXzVglDUWu3olCM6ouWmi0Xkc
YE96zZqZs0QN6FCRdR6HAiE5sWMQ//dPCOkrBpQwNeF/zled0D0UCuF3597dfMc0
mzcwuhAax0v23pEVM4IiwgJs+sLA5fjdHi6vRCtrbhG5+3yV4iWI+gGlEVGrvu1Z
uDiJNBLLkFdKVTkMpbHLMd3uZAUGUTZfxpX1tPENn25qWO1n6FgkqIONd+n0ymDz
/WJ1loQIPrVJJcfMdB9ae4oqfBs5KWmRJvRWEWqokr3Bdv1PsJFxBMO9QusQFvDw
esR3jcDtDAlcUw1+vlTMUt6At475PjWqEFImyf48bVwiKoriCd7QqvMV/7yVUBmw
oI42bp00zWE8qrZf/tjS0r/lJZbMdL2H99aW2cLyfvLVnc2iD1CBTQh6mVADkTIB
mDxY/yQH1hl+Qmo28eK9CkFs0CouKccIwTiKE9qUiNrhXnP8n1N75bjaJejZTQRn
vqa8T9dS5LbJXs47bRcuPCfdP061U5lZtUJrtDr7QWwPEMxupyuLxoqnvt14k/P1
KxcfJSDMaZ+IwklkQhb2lqXne65uvugVJmfdzbx8aryOwL3KGrA6YmjznLs+A1ZH
xrplqJVQd8rBLaIH0aGK4x3y4byi9IkVJE7cb5sq3bI7BdIzEpgTED3eDMogRlW6
AKEG+HEI0Q7zrBHViz9ynQePfigNnE2Lu2gowr6BCtM5efIJigii43CSo7lmwgDO
TJ3DUA1B1IPSs94JFBbHd2hJRvRsAdKDD0H5ny9mQnGs3z1G1vM6JfWdI/nv+AKk
2+XmmZQJ7l4YWwsOVO9R5dkADnP/dB5rYaAZobC8ktDmvmA4zm2C9iSqQ1v8EIX6
EKGQw0CKTUAx/mkVjyslU1afQGgVNaamIzCxz67NfXr//L/mCnfcs1FSVlYisjR0
rMAkHG1+ZCoiJhwdjTbsGJ0S1RsqgJu0Fgldf/lo2L6xgLO46UxrAh2LkX22wxUC
Vf7PNbbyOwXvvzfcOJW1gBQv58SSDqntlkAgJgfjx2mrETV+/G/hlqhx5xMFuG/V
qEiR0cKimxkEzvpUV17IvnqhmwFo+x49Wrgu44SfYxPegSDhbrIcS+VzKciuYT7Q
/6eBXDRmxVHa28ekl6o4nxXduCWRwBleBLl7BiWR3og0iESNuDPXFUd56XphQfsE
jNordQf303cjQmAME0u+PwBlor8hjEgBU0n20+EJkt9bm6GYc+NONxBE7SQHL1+J
oZAunNNLR0mqyE2OwWY4T2qr5eiEPeLI7TTb+mxllhoJ4aFK6N836FPnMrDpizHJ
KtdDJeGEvSY27R/+SNMGCbfX19z102cdNAfkcJWBQlN6ZdymlfaNke/5ckGag8a8
+PtYHgR0WzWh54Mbs1rvjwmsFTrFDIr89U9QcJZgYhxutB+42tQsHoPhS/RjqCnG
x0euFmwc7rOEQVBPJRnrvx6NJy6ISINXIJAk611wAPlz9urx7TnYxZBrYY6T6M00
NTgArP2H3t2vXp7Uov5zDCv+3vgxQw71g6ThEx4QiaRDGbgYyPjJ1FvBLGH5Tpr+
Nx3FNR/aXOZ5MNIuFn3+EaV9nJaCfuqX1JhJmBZG5AkgEKMe/zGWyvG11mlga3O8
Yks1gqpiKI/Yxf77KYdAswN5jBY/YY5X/OPG3/z3lvisucsOwjFMLVY1boYHDETW
3PNOnJUXEy3ZOyZ18zpb6JE+VhPfkEjVco22j7zDBMXt9WpTh243sXN+HPiOoG/t
6xc0e8rByjSLRD1oWFGnoYFu/eNH6TAnQGMC4sc4wn4K1f37KoV9DQ3FscPEjfpf
jab28EwQikGdrhBg1Bq8bt9IipQwnoZkhYt5DDBmTf3MpYfpa/aVoIi60pfnKLh6
xCM7QkrPEwP/I+7pFYt2EbMkfK39r4L5I5U2aVjlXeOXt3o1eYViZ5q5Bxyc15Fl
PZGDwrUFH7J01DzjVIj7BPiwtuIq6do7ArcxAY4rF0BxLtNogM5yTQhauX/GRLxH
m0HQtOQgSv8gzUKNCsfhEZvVmF5VMxCeiGjkdTSj2KPiEIjgQCmSx+vGdjhegaDQ
wgTLBFWimAwUwhuMQ0WFEOrMIJHctpKW0ZRABqtR70XR6gfiVd8j6qeYgCkulP5Q
OBreEMe/51TYhSev3RLLyEI8HT3Hu5rP+srQshHG53fkutgCNkbWB7Wv65KGF1Fa
GphJGWt+fA7ugGEkzpefFSHDkxxyhGCyH8pg0d+yZH1VEAHO+c1aFWR69CLe+U1/
8Fr1T9FWhi91lwVYrvDrSF2AYLjeDxZNgtIiHB370VZc0wX6i/csKU2Quqri77lv
DRNq/uhljbk53BMH4nlByImJ90G8Soks82x1Wt52CTWEVRWedUzzWzCPmZhkBIcv
33LGJB4de9my88Pyll2mSXGupF5Mcl8R6MVhCsR7wPrxbu1RstAIAXYIIYXOkOML
lqkiLW+DUPG219XEb9t4JPuhxlefUYuZJBGZtbnELTrMxUylk0yBgnm/FCmB/55T
uzlWoG60fxQhbSN7KWPslv5e4UHGBHqPWcALTwgOsm5LhWR95wX47pi+hXzuEI+f
AjZ85q9ro4iDAnVu/94opNigKKcmZk/480JMOO2vCrxpqZn5wxRxZSBMbl6f7afZ
plzYNKP9jV42T2ySmKJwkn6XImFyznuQDPvHLc6fJcXZF4/iQrl9tasMsK+RnzVM
ggUWBUoV7wgvyyM3VLgJSqLYqD0sRVBOXEzYGqCJtoR1vSEeVSI2goSakgysrMBA
9TI063pfpYze5uw6mWxaE2Vw4yBaJxrvTDdkKz+cPYzWlIKsRDTYiRWzFrXelHLN
ARf3hnmu8qRE7H9krr4MgGFeaS89fVEsqHYa6fFMnl3Fr9SsTMNJSaQ/o2DlvAF2
nW47tuhMknkr9MA6ky6Kmx00492lL/yKIqv1gztbH9W3kJpNxctVRhuGOPlpYwxh
UzwpRNIj+2S5DsHAXok/yNVPAxCxH1umVLcjetw6P2gyiFfdsW7I6VSlu9g/MBQR
jmPW71Vv6R5SNG5mA9pN+z2MWOtGTDyYEqmrwiOYszU3cl6gRDe5asrN7rm6h2Ib
REB1lD3DDEvWCJAmLa3+EqI6Pd/Xg202Js6J/t3JZtiTb9w3AttevmEM8t88N0y8
pl7WSi+YrPKcT8aufdsQQjRooE5+fJ17px5K5By7PVgMQFApo9b+6kQk1K5r485c
POkXS0i38CT3XbwSCEK08tG6xSNgZr2caEsX1L3h5ypKTyXXX8Ool5PhZv0ImHpL
jDo5hVvYKccNE8YPxX80zJUrpwt6pDptjw2oJvrMgvpsaQ2kPa/YngRF2n0qf8fe
IcVgJ8n74paMB/FiWMAALLCfYvLlGKPF6Ael3Qi6M2HnQzntQ46Vc76UPPOivgT6
nclzGUmY08PGXgtN4tItDbLPDrXCBk84EJWmmCoibgiEy3mB6vmr1P7lHu3WMrDO
f6zIa7B1W4uXrYyRKUE49gxzIq5Q2m7oypzBDdTrm2j+ZUglxTt/vyC3VlG6k5+P
LFr6tHgNnwKyzaDkbB7vHoCqojUaddFkC/WT6zpaWFr5f3SG/xzjTScFNt3ejNqN
auUGq1U4yejl+orn7xwPhSO/9ixZc0rc1IaRbKEbNUx5QQjVSEjdHfpuRmJSdhVb
rMlqeXdRxdsdWLkHhFEF15/rNBTavNeFQ2xnmd2ZnSQ6zJlSLiuKW/ZFpL++eqWS
dSYzqiQ2u88GvU6EUKezvK1NBhz6xWyMKUXo84+xoclt/hGYjCTsTnzls+muFCA1
zTh/4ZklaPbsWci5hLMc1Be/p3rLDsqcYOMTvH/c8S/ivdZUTsLSrlYm5rnURTgn
8KKuCsZRyt1UjAYcaDj/3GlCIHjD58huYMYcPzKk0V6kEFyImEj+36lj7I3i2uRT
hul4yPs3iCqPWcHG4lqo++YjYoqYuLQsY/YUBCdzPxR9N9DbEJ4i0nuIV7W293tZ
0+IEqnHBYmkWOycOxQ0sDf/+ZyP9NVaficROunDaGzz6JCuqZ2ekjKPz2iPVyWQ6
qr6rddiohhf+pCGVlivzqVkGkcSWxaW52zwF6AxN3/SixoO4vzUtrFiMIU81hz3O
9/JyKlKv80KJfEqZEqrrBWDGMCg8YzfdhbHgB6oeGeiaJ3BUYv88Z++ympsHxF//
LwoypH3gJ0vP+MD12EhYbyHKxyaX8/bV43BPauR1Sdf1r2M7rsiXFa3nhpOr5GNi
z/Z/5bcW326hhZBTGCmCUaYbH/HPt4UtVpZRljfFF46E4WikmIdEdIwT1j5RpY9V
aQ3ZgcWgs8N/wEEeRQ1cW8u/5aMoEojYNgQgOyfYO/O/QddiW8B8aBvgl5jYMom7
uun1HimABpFqRVaPaIZNYBAOuGQntWvlq4RlTTnqX2v1ZhWzsTCWeeH5vJLUADBU
fAdbUMI4gvZQyGtg4Qx+pVEcaNFHZ4fsItPMEucE10Du7/fzLLsbLksEsEa0dfLr
Br/BVqxAuVVrP+k2oWRdEveyJBA+lIte1OiC1y6ap3HlWIUt04i2J8IZCD8aBSDp
5xG5M+mqT621zLEGhxb9MQN7JXGpwy89K5lm6f7H6McSM2Ft66Q8LKGavqKb5J5l
Yp7Qf1GEJEDy+/GaCMDJ6zKd0Y8Goqk+Fld8N8cQwgVylEG9feu85238prjfnNgt
5WqwfLKChB2RHDzkZcChqYu9Y5M7PfwDmhbN2+p7lA+Y58E4EMNAItAN5oeiQ4SZ
TZCSIVR6Ko4FVwWPa7+zDFdUx5UwtTdCV04sn1pWkj/H/vClen9h0869deYV/1O3
jIWHL0Fqekn3t6xYHcYPTm3nbkms1mTnD/DoA4xS/N5sRsVqtNap4e30Z2y6qWMP
n8Yxol2GH5xYhrFurwzAVE1FOpVG61COhl6kn1qg3Oq5kPzqzbUZ5MQEg6syD1v5
UeQObxVXicAwoUM1NHbYXDx/6/gvKXfGKCNqZoTGUSxKKa1pjKFFZG3IlfAuXHgr
/nSYaK5Lk3X9jvjbIy+RkCgSifGScw91LyxZNqz5mUpzwaSskgIpZoHadvbb722t
LewZQ7niwctxrA1VKeQpu5FvLRz33sxDS1tIP05fn3zNk62rEXhp7ZTwyyjb3yGT
N/+LF2QPtlKik8aiHbvSXCm6/EEdiiDZLPeYExT50B6m3KONODsGpbcGSo55koH8
yutQFEoHhiL1JJ8l5Dd4NcorlJcY6I3oXGViDBtKEhzFVMPUVoPbpgv+wqrkghip
kqx8mPQiVFYiOo7QQ+OrPusHdQk/m8q+VmV4TIq7b7zWpKJzA170YY40zoh9WB/m
FlOgNO+PO/LvmJg9Aci8CfAPzWKyjXQh8C6vJzeSvuWuCJ6mifQ5i/4CGJVTwQWI
Txx8LOytJ3bwSvi4/9IJO+4yJWuZSuNnVj/tvDoIUwhXAzMPqmIKW9TfiCObkcEb
k2felDe0j/CjkbfX/7zzPRNEKW3//XD4TCci7VRqgptO6aMVNYPBCwGVXRjGJZXS
8bVcK1AmIWe8FZS+k5daoFokaquQRXQq62Pe/41WUrWEChz3vgrU2vPdQIaFzcVC
Ii/YtCpeRnl5vFvwvLRBHwe2TmqY1LSl1YyCU7EVBJx+q88fzWVY8zxA9/l9Lmw+
SgAl0noRGGhA/wLWFDjCMvv3G0cRJ62qia6NFcUV9GZN1Y9c9h9pD7hG+2W3W5bh
XBolOOVoYT5w+i/MQ7Ey5xXwAConHXSEo+N2dBylfquO/G9Jwdmszufde54qHUq9
lxe+rwUkdX+3hJ1N265qhFIJ2CZtYetmEyBoBvGxZf71u4XOi9bjdgbMbrIAz1LW
P1WWAjbUjU66NirugR3XzxbuA8sMFLtS1YzXbqFvmD8zNghyu7DU9UzTlNG2RTYF
2gx9QP24REMgYCS9DoMfQNh+3k7EJvPYpypkcqynZDt5dEuUxzVTf3ndfUhr85zu
4WHxxxLhy77nywLo3zTM10ApMDBBotiHHBivb8oreZMEHhb2QZwyzMkQxf1aZ/3W
OyFvRaPhF0BE78UnLlv/I+ZhoSdcPQvE+p/OvfqWsp3COh0Mybfnc+2GkkjBLuJE
gXLLC6XBsBSAuLhgeeH0QVztOA13iIxlGvH8a008imeGNePiCDs82kHUGEOgfsW3
nJOwBCNCJCWdtV5R9Dp/gqs2Ag0xbsZk6gY4t5Pzpa0Iw//A1HqG9W/AJ6GBo63j
797/bgApvUJ8LfiVe7nM0w0MB1C0Q11J7mV6n8HG+60x1JiO+rT+6pJfkSDROgm3
eZFMda4SCdf5WZaDXJACSCTEfbKhzEzP81wW6v/dasLBr355vWYrs3qkQdOfyHl0
w+GvOUM2loMq+feuUJN4TstsRbuB/xVcfHkJ07KObIxZmgXPXROWwy78Oyf36stq
dLYz1EL4vqCqHLUT6lCMJkz1i9XaboDWsCZ3Z1Lswj+dtz6zxWkUOZ7RnzyTKNFr
krEypLd4gx9AeOp6DpdagxA2W3UpPYDY87DOXaU3x81nNmCXbOe7X7zUK7ILZzLb
vmnXB0CX8PbnR6J0Pv8l5zFm/2Nh6cCD+ZvXZffNt0WnglGqb79yrz9JBgEi5Q0+
1AS6XssVv29BYfHkE44U9oy8x7cdA3tFVmSm2IoMkefjr44KlLi4ywjHNodwwBt1
ceAhCabW0WMQxXcMpLIi+mdAh8M2W9Q5YJ4CvwwLbv/EyPTg813NMbVb2EqnfRLk
thf3DjEcbvLxgkCVGZRj2KCstxVc4aSBy+mnNXdUEydFqFO3elUI8tSAxP+QDzXk
W+Bp+MXdi022TbUPQsgN55v1eBOV7PdACLzjLyvQ+beyd5nC4JIuwF7XF1OaDLGN
RbYJIlEQU4w3ioVQgxv8JOxW6m9Ero3ktT0Tcz1zxPU/6Nrf5sndR/rxm+mjMdXz
8BKgVbe7yPmauzSLY9/AhujamasZl41351glXuS+qyv72ao4+MjSACVySOoN9WXO
D2SOPsjxQx1JhHgov6sxgNE2XgpyV4XYEJd9R+XingjNExawqVAq0pjh5v9g2Sh9
qVvzSE45zlGY2h4vERwcGV5IzLVowGfcvFfiDpHTqGx0uCqICMH317aV0Pzc5iNl
tMVBoG6rikjZB10SrwXDx1nF/KTldIQuaMSENYAeDqhMahgtKghzVJsu0x/8PN7X
6xnJkx4/yTazCO6mOs7STZkdTfHYOltG9ZeZTSRJ9KvN8sG27OAzkJtpO/y96SVD
WxQ2OZb3uFVfO7+YTNp9ZjZBdwOcEv/tzpM0tVPf5kgR/5Sk0b0swm3yJXgFoIRn
55uDoIg/2m1xVBwqgsKvUhpiyxsWMl1dETfhico7QjnS+EuHJ7gEyRcVxXeagOEv
2hGjHJorxpZvVNp9lAi/zrZPGI3DJmBQ5SAOXjGbMQR0HGvwWEDgMsfL478sv3sP
92r1svEKVFCVzO5DJdGI0MwlKavV6ogJKN1kZlcGnFgBOScJ7PLfa3u2cKBedE7z
D4sSMzReMAMOWKoqJp90u8o0xeYlzYKg0rEabSMMfB0+5Z5whxUuuQlMpEsHpGc0
ck9t6XIEnoGpaL7YbksRKjcqlmsn+Ts4P4uonTbmNF0KmQWr5cFwCRUfTqo1WGvS
Lvq7HiafGzkTXC4XaF72GdWDIzp9ovosoQpgulFrmBRvNXH2KXa2QuJq4lHsOium
34uQWwspricL0QA28P9+5EnatA2N80OInWpOSkNcTuwQbFqaD4vH2aX3R90peF7e
gICJQ6jZE/k0TLHUy0agHgQq0RyL+KyLcPU9QcwFIm0ls7RPaScEyGYAnLe0P2rH
ITGV4BvZzASPlGbggqqqf3b4fkmd8LCEwAnTXDo4q4HZ361m+3/cYjYBMOwfMMF3
EVGq7vq/gnvDRk5p/d5p6h0L/1mGu63wzRFSOkTDIzm0ngy9pBQEm6rPFQlu2FYb
AgR7S8wfsQQaOhoKBVEFiBn2qAEADeKWST+kV3CBNb+R2DJeUsVQ7xSVecmfMN3X
/fYcxj8yGdzoWJsC8WQXHKzk5mG7KcnsiiUaXmOCtO2wCeZLcTxMfzkn6d5gPLqB
slXQGgz07r1ax0UazwAIzjBfO7ty8iXP4R7jgcyUYjaXaEWy+IDMtSKZ/IB56ZRG
5XHVOu0YWr5s/bl2+xK2YLZUwCmVNgcoWVZaMkySlXIJMaSuS9XYYGblMRe8DIE5
Oz0ytYP/8zQOtmMBICi0U5RMpLEVje9dnqbimffM/DVQqlzSAwGEga/Knj3oXbE1
ffPuUELG8uyOULYuLp9b91bTM4GcF8qxUqxpGARgPQR57FolM+0VPuJxyYevspZl
mNzLjk0qFFU+iy3j/fjL2j2Sxl/CBG3DZH1UxHUdTcnfJzTptiZ7m7jvE3OtHnt1
fuTr7tguNX2qj89X29AfSq1cgGIRJXSmiLOr2MuDKcJiTMFlZrQrDVPTjsn885tV
uy6ZX8CascoURe4IeCpqoSEauRygp+50rF4CUXdMR6eeVvanA2UAxVDBJdWRT5m/
WMUkT7lv+FLnXp1xtesv0a/bGiQnWPpNgs/613eJcoblt5K35TGx8Lr9C9GEBl/+
LYoap2bWQP6nEAm0sSUQ+LPuMLL8Py+cz87FEWGjuTquDj4PAU/9IFsp48kpAPZk
aG20Z2vxiPoNWG3nmz1Azk5ffJXkt/RMFJWfKwEzAUQnU/2ZnguJiM20SNUmpM9d
nzdvWaTfu8koVeIATabmQ6uyZNlqmfClR8kQtDx+jF/WFEYprXCICOIAov0Z5AJS
L+MwtKSXCJoLG4EhpcMdBe/uH/RqnEg7yN0Do5VwSssUGJpL6rpGDLuONPd2GugP
YLQGpCdTcKCzgyO9CtFWyrYvXRpbhy+npCepDSsLxNOHH2v1N3lokTYOoa08MKUl
g35ttikfmb4KdQk3s3vTjfokxsKdn1SoYPY4Kts+wKZkw9x+5s65H5aubh+usFHH
2/NX0jNwyrp67n7ZGU5HnNuddc5W8KN2AmNj7V6F/XCN+m9l0F9GjhWCDaGY3Sp8
hyWIPF+LF4102XsWqf9JI1afTChkc+/lBUK8BbvladhBA7Kfc/hWd3LqFV+DtBUt
lNSq+omI/myN32ctk/QUzmL9a+k2YRz9giejuYtJYIOYjmGbuDoYicPMIxu9vgPM
SmzFuqMVa9gaN46VAezRCU7VZV30IgPXvW3yMMp4IVROQNMaJkLYpz3yjBog1rSf
ln7tpYPVbum5Stw6VX83ls6SVwfhLkFCmvL+5M1UR7ipCc7PnEj7RswVPbTCgQg9
+yqh40k9Mp6MhXePuCvfgjtDGkBF2MMfADk19dAcXprUSIjxKbq869R8Uc6MXizX
QkrRg8bwa+KO4BFZuMzKPr8vJvUZ229xTOBKVNjP1lLOf+SqPuVJ8Pu6dKjvuIF1
pezqGov2doZIakdLIg4iHabRPfeLUD6dCB5gdc1snwqDi7JGxWHHJGUTy3J2eo3w
YhJL7H8oRkYPhH3gTNZbh/Z4ap1f+NnyKcKH4hiV2UlqRxKt4sGI76ILISXmIsVu
TwDpMvh9paFb9/bSLK5bi7gmRcNXw6fUdDo3hvi8v+edKrWv5OGCKBec3Ii+Tifx
HPeBivwU+bLqgthKS4psNIuyZjIdgTJP4eIdbvBeQAA2PjRwXS4ZLl4WbWVM67zm
qJUjCSReBcXUjk/urz9UyeUEnXeDOzKVEhZbyUJtKNQIEKD08rxpQHMCIAq+kn5B
UB1ZJfxR8gELbSAilBOJ+nVSL0vc2lF8K7HT56XQ+0WglePJz9s4KLJRLlhYeque
31+3RBgXFP/veMDZcMzR02xwEddQPlUOaBGgpEgf9gsD0qIQes001VboGRSawHEt
6RY8L5bqps+WGgf3Q1KXvL0YIIym13PG0pINlbD1hgqO4XtmByLScwRNY5HWNUXg
fRV0gwV7pxs5G45OjGqvnDTIPzrZYaAlWys7/HPkJq3VbWhd0ldpVVqcmFhPuaFh
+d90B3EcexN9cJ+UGzZ3JRbaqGin7QEm2StAZOmyG5+hIvkfcB/cEiS+fd0e1vuZ
qRB0ca6rQXdN0G8AY32938lfZAzcYC3NN/r1FkdgBuyOrHc99A6tk2Bv5HXwKApI
/BFm0lM0K6PqH9C4NLUZdZPZ09VykM18GMEt95UzKXefT0yVZATcrfyX4cVFWXt+
qbHKAVbD5OT5IowcYw8OSblkXPQhVenAMqevLZLa4Djsw0uvRCkB4Eh4U/gt8c1y
fAjCwtzh1AJcWOYJDGzlUUx9Kra5jf0uTzoksWkkgv664Lqx7P2W8FQoKm0EGB5N
2P1ZhojlJETRaBPzT146LlWJfk4HL+S/Z3MIKnInOsPFggRkHrRlJ59+5wH/q+dz
fg/2tIKM7HRNsyJlTAcEdE6WsKQ0tMhY2Ou7gSX1U5SVok4wVH4dg8M3Q+JAqVCD
alYUddsMZZGJd4NyoqMk8/0gcK/4YrDTnkZXMzCHLnLZovtQH07WpUUuKRg57wp6
c3pMn2n1t/cB5XvCwlbTSxuGmEUO2YSx1jG4BNgQOicKGYcnAMiGPeO3i/RyTQhq
t+x3MLzrcDMzA0iyjdMsb/jEBB1RM/X8ua37Nna25ILw6rt3OJq2eWe6fJzxBnck
3K75ZOke9P5rDcBKNlcMQ75QkLu7o2xm7QrdZd/4lQa2ZuAv5A67iDaj/I9laYA1
QLgVy/RbCGFFxeZlAJBJP8ygpM+5QQSC5d889pUdx+EXVaSBV0U9+FKDpS52Ahim
r4ObTvVkuDvzhA7PC8QOfLrq1y6X4u09qzDTCQ4zDJYjXjC7adjIo5LR0iSAirlA
Qo8xQb9nOhrQueUuFGsqE/r9M4XEku0T9gFenCXUXfmLCLZadJy4go2SGOSlH4/8
cissNL8ouiln6hJh29qF3NT0scaQ6lcvcXelasX064FKDpUKLfyGUsfUn+keBaxR
gOFWYmnajAtQIbpTimtb+wdzBpHi3lqVAazej5emQkujAM4yKQEMqKsqOrWwtZ5x
cyrLB4fuVJKvNH/DnnqHQgpoVU90MgD9piphI6sBt7pzpqDDWqBAovIztgciuti1
qFbV30xcLsn744YDe5CQUxIS4yljrfx0Mx+8dwqRNSlIuYALGcU7QFpj7qzsjquL
yhW8chogsrF4uXCSNI4UIAFTFvBPx95b8lFA6uOqxper1t2hhkNnfgWcqEubfSgl
V3Aa8iR039jTpEXN3gA5J79aLqnS4Eutty07xD+38/HSej/P1uFbU5bsMbey/Uro
VPNrIsvGGbHmkrc9nc664W5q671qCUjLsI2TMQPUO6Bairem2ahAhgUczDmK8SFX
lj0ORe4/4bdz3v1Urj6waKaaKyJ6zMobL7rWyg8FHG/HNubuGUMCJHIZ3Xvq02hh
LlScDLo+JcHPTKY4zNfyGcSaaKX9cKjmX02K4aC58K3CnvaoSU/Q6ElxRsIVuzPa
+6sBO532J5x0283+W6sXew0AAXZQFzLbhfa9raxAvKuYNmm1rXLdq982t3/btfug
nVzoci3R4/1bicyxQdV1OUihy1np6PbA6H2NCiMZEgL8Dm/p5+ge+RqaCE+Jm3su
QsA+Mg4jdRaVxNLfm+1HNAY0nfqaPXlUUoooZ+hbqHWf1SujDN1idfJ0/TDkUUfC
BsCck7cpA0mD5/8sF4AjqMAB/++Lq2eKsu0MxuAdtCGoNBdoBFUgm5HemDnLjL8u
QrHiVsPa3WwG1Poxde4qrALegxwBkRmsGn2r5jiamsAd3bQTEEJSW+yyLaWDHRTz
3UgZnFrb01IEOOPQhccWJWfsz5b5Drhou4WzBUAfN+1fabEBYxccHPH77bVNwrQv
FKCksu/YSyBidd1LehrXHbhPGENZs7v9yJda8skXW8bMbcrc/E5RambS+W0z/DU9
NO0IwdkMgUSe44Zq4Ql7r2SMBt4Y1QsYgeQMOvLHnBWsIj2GLg+TROD13L3twojH
cZsLnEWYaSrWdxb/SwY3QUIWWm1rpV7cLvCZ1OBJaFTOzWyIB8ZPI+BlIWzTDt8e
ShYFVfYlvjPjrn42tzKSImqPxaR51+Tp5CRBQpNDG6hAM74uXI3hbamBU3DqmL1L
Fbu9pNCmbIKXrzexLIZMMb4CZ4UeNsa1L+xQ0p3dpVe09+UZR3bLbpXOm2ZwDD7i
J+xpUTwSZh+ksv0B+fATkBcGy8XSafPiWth0Q+pSONgbddj5YcuqThyqI8AzELiS
Y82fEhplyd4lgIz/i5aketZreFL7TPedgiYNLhDnysIS0TDjtKsuEqRdOTltgrZV
BQouPAaP4r/3IWUE+ix5kSg5TajAIhcD01cApRlo9+nxnc6PId1c1owvjSTXkgnU
SMaVajhWVzBXf8V7XA9y06eLoyclzQzz+hWNPNAQiNmuaxH1KIK3Dz0D/cgpWAJA
h877OWhnGryvHMFcEwTZBILt89lhiVTuZilPcZL9/qXMx2PDmNp8BtuWqKPITf0e
JCtpa2jBsz5jTMUZ6xCRNx0qHHIq+jSTsHj/uu5RJW04Ho+ttzTupkrIKelHCDCk
1+sX4ZrzeVrKI6OMSl2eM4K6W+/xADVuOb4w7pRWla2Wx90T/a20i5dJhmaGEpvB
noNF9J+mRv8Q6NhbWEOH2Yl6QN99Pi0azN8bIEY3MZHVbv3BSfjU2FVPdeAhOqBC
Pbn5K6PV6Mf9S2clTVJEydRpR/VHt00NUMxamVnNVoYJ1D1ykfskZnJT2ourJVip
6zXgUAvxWQ9eWJICEiaNvmYiLNHQNCsVlNp4b9bsopl+2hz4l/8DMsEU6etvDkCl
ser1d03WCDxfDfzuoYAdSJbP9b/K3ao2bVuYigEOsmxh8ldKSOQsNtvQRYNCYofR
jlU6ygO9Zo6vfZwJdSG2wfWxC3awT9aBSuvOQLDD6gp/MNVmzYTAW5UjduqZRtwo
84kUi07gQnA4nZ+XvK3TPr0Y8lb/WXZGJloxvmx933IJ9SexNOjaO9BrPyWUUkRm
0O87R4WUUVPI8r4SK8ZCj8yU1L5aJzK4XvkB0PzbFJTKDu4zlPUJLkndJXMCfNfU
/eeIjfaltBYMa3WhRGEH8Wwq6iIpZBsxe4cK0q32ghLrA7M+jXMj9zlYLIuXjc7Y
ueApo3uJ/cevBqoWbScrPIFxIKQin9SgKN97ZJ1qrRnfOn68S2JHXLVMmtn5BQRV
h5w8cDmbcijwROcyIOrG4O/cJAEQu/FwPZohswe1Z0ycvbrh+jmWs0daQuHAltyo
1CcePwyM7S/2Q2AMiUXmBw6eRB+CoE+dS7B/ScWUopp7FI+0lDKFMQTZoYzPesHa
zHbrcxPdi4VK8B0Rk6EIP/ZMZIbWYd469lDiDezqqk9SZAKdaJzGvlxf23+8/eFg
+9q3i02h1s8UVitcbv/v5q/G9ArgilTuvtcssh/4EDqgV+CNzAJuv/RW7JvrdKL2
Js1cWwma6X5uvXLiRkCqBXeYmLu6Tc2Xh8nBjRD5Ck4qFGcJsvq4N8xnKT7wWuNI
LLK0ChmPvgblz4H7Tzbs0sS5meFj24aFxWj5lbtWhA0dXPsRV8t0C1WGoVUK4dqr
Eqc2YNMI+HNdjuLOP0HaX+FSzO+uBjLHgv9eZxJi3SL1TxbuGLCjmm6mRFZKZ1or
rTgYeGKonjbLbL+vIQrmoCSrr7g1HUCZf4+vsvi/hpbM3KNbarAdjEF07tDZpbDf
NwFOIIl8DqN3Td2CcMbVDCN6McQ7vcKWKs2GuX1wJjzjf8RkRd1tzVj9WjT8Kg2g
wKlaP88Mshn7O6VinDrhQM+R26k8PlU5RyreaF8oY6JIY9xTpK5Rt7rkp9ZuvQzb
5cC+YyeDY2EZDYfcKcAA/TuJav9ZNky7Un92HJnNwdveHAIAIu42xt3rGYkUab/M
xAB7poRrBSnvvVHbT1f1+WUGoA/RS1Oc4hhb9THOvbj1321n7gFuplMlFcXMz3at
eMip4+PmfAvbgmi/2wEiiY3JepWcjIvAvVktb2oVhpqpFWYaney/kGHfq3vGkFP/
+blbtPQMVdDpKW5KJPZQrm2ppwAXmqzj62q0o0cVHVOuKJ7aG4+wJh4a3vyaWmBw
sLKE/eoB6PBLSFAkHyCcBPojQktrgZzi0NsPLTjM2MYvxiDSbCDXhsdmLo5qf2jl
u37C7LQ9qUe1Uu06QGItpS8J5o2N+n4RxLNmNjQwnXd2KOmMCW2oTjPtyhNHm0ek
W1v4E3PAZBblnzN5NDrXwfRREAFxn3glInYIcRIPMpmGVFy8+Lkl8pyPYNiWgKBx
ZsjDOcP5WMp7RvYVYLoLo3642/zIUf0NjbDHeoJlEWukwpFF3IP7Ai8m7FDE0G+W
I/xK7DQM4M822yGyt+DjVUaKH1hSW7FoMqIWz2ADVjSLXNSHPIwJEn3c97TQJSbr
MYev0mpIqwAalEVoHcAL4spDCzukpZl+isR4jxW9Ide54/Bl/g0rLR5k2m/CpBjX
9xSk9aCJDlNLcFapGPPBvVpr9eMnY26FQVu8IABzEUGBXpU6bPZiLBAPckDWQrpS
xzsfzML+lsDMMfWX17MRQcrya1PMK+l+Mi3CEYQgW266yVMY65UACN6xPXJ6jG+R
JuXhK+oeTcrzYcpC6qjrkn67583nIgBQ4LKaES70DbipiVbSeI6ZSwCfeGxZXQMr
PYoFir1xHleez6Ul3vWVfBchJ0Fdgai65vrq1wCNNqh68wy4bilVMAK/t8Qvmu2x
PDa4k/WvQYFbdrTXClguhJymIgQetN5Vnwt9g6Eg6RsUJMo3DtKUd4M/gbQmXVH0
l6ba8gBqUtSjFtw3uir3dIJxauRXStwgIRTxhV4M25lXbqA5kRnUuOT4woUXzqZe
CagGrynlkXwSfiWBh0qcrcx6mA+dvlUgYSkMDagtWwCIpx+R8Fx3tPm6L9RDexZB
hIXRSrloNe7UOqRc0Q9TSgbGNjRb6jJL+a0MGsbANYPO0TPQi0rh6m0yDE3wyfdH
pL302L4lFKbeTJ6ObwGVcEFoGv3ZBkk/jKVakko5F6SLOSD5vUOJq3pfVDjI1poY
s5GgF1CEfMMKztCCf7uggRqO4i+PNY0OLX39h9QG8l8H4UNIk5K+t6Su1S9l5awV
WAyx7Z8347mbqlhofBLmtr9m4zFsakc1pstHcMM8FL49EpfD+Jv4VadFVjNRDq64
7c+EGpbmvCkpBbjHRZXznSKnIiceKQQUNL66tLybeVr0WmYFmiakS/gCjKiRP4jb
ljuQV3ebx/x+VweI37P3NHEgSC39wbGo5w++Dc+hnsdqRHY74+1mj7ieLFskMl1s
ZDay4CDh5jbDqnxTfWAzxnBMOAdUlTfZK6f5SjR9+gUFSVVFwOq7oVMo3bhQQ5uQ
wo34AfBmwYIcW5lmKHlLGuM9YzcoqeTDxT4uEahpmXHl63MFauZT95jAF6YttVHx
V3jFXCDt90DsmxICI+3QCKN9SG2JnBFNSrEcQaPyVyVyX09Q+T5+HF0Bh9CnBgTX
sQjmx69229DVWJTQ9/dRymc89EjJ+xWxsJFeRQZz2CQkU3bZYCXhHnUiWm7k6k5u
SLgpvdtJD0jLHsCcPXX/MYixOBImbV7BD0ttoCyTRGkfsZ/0y4SxFEyZm5S7QfVy
3vNmkJNZjN5AfYbNYHxqemyJeL+p3nWlgQGJs3upfzKOP+/b17o5Sqsq1g9rt5Jx
MV2pOUI9CJG7qVwFHtk98OrLM6/UuHQ8M9uqu9iQawewCMjT5l4CXcbcHcu8zqKM
i/Xjsl+DPBbcs5sUCkLoh78h8HofhEtuzLODYeqRVcZKOWmlQYBroIPLymMIPcpo
1wr+7KXjfzTpFVq+cdZDmH1sJdJCFZwi/S0trz2bDq4Bv1EHYLvo5TTHe3K2STax
VI8WmDT1E5eIZySmMcRAZaRSQs0O4YbTN7O/ViLg+81nZpT2ahQqoWJJKwE0nE6r
jW/GhL4e1USEif1ipFVPz9TEf8umPf5h/f6q7iRbLS3GRRXf3Y/BJQBfr93xqZ3r
CD0upgdWJfbiHJsZ0dK5kXtkAhNfB2uwWLNqCGeQ5LxJXT056ClM/HX5QCJeC799
SjZXGtMQbOMFcjhGdgF38YyLC8Z6Keaw7eFunZOB/YUaiaReM172Cm8DDKz/wj7C
iIF4LB8OK+M5WpTAu+s90lshZthDLDcOUQKEDZQk7ELy3nuJH6Fd6GaTB5RLyAR8
LjF5BHQnl6syRGSF87fx/2ZCXrQmvmkFLm3GqmT4Ug68qpvhQktDUR+vAtE1uf4u
/H7HmNL57sPQn6EwW8u4OB2lJOt1uIWAccMaWjD1qCcX/5GO+tdtmijTnqX2iPEA
rYMog0j8XYdUEVQ8hLs/UjNnOtVGt5VTKTft2mkDbxo3QI5lSR+aywzB+w/t08T1
8ncN1pHkmYH8eiFitz71schxLFTjZAqo/XpKL42k3woimjsvKsZDTWmxTaNDcJXO
D29sY6mF+GUq9eqBM/q6uUgozN3ZRK73M+PiKDTZilGPjE/6pvgcyqnTQR7UGhuP
LO6bZttiVaXi6ZxyB0qwaGe18nN+2yOgi5LlDm9mBdzUpIieL/r48bW6ebK4lO+R
061CcpCkBLGHJYGYZaPkMo2Kb4x2bbLvMrmgs71nO8lyFK6S1LNPXrnW9HhDaxP9
hfiK8lt3peYc3OkM7rL6S/LaZjzhHHhUkbjEOaeCftPCTDsrkHHCdFiInKYHb3oo
ELK3EC7eDl+IcGribnzUzfH+4GMRYj2KJH0gToCUZ3HDKWbt3XAjMGCCPfAHdmUZ
zyf+y9HZ0hHIxtbpY0hZ3pCD88832r6lv4YwBwQiXNoFKu+Q6vLvtYWcTamXb0JU
TdIRMXuDRrpvz+McPJ8kQk6Z3V7LwjlelTd3HeRZp52bCckMq6aC43dmob/n2wHL
V7EYDUo3Z3qWXYI/SiXsWNNshBdkGabIxJomY6NHkyhJqpfyzTlE33Spl9GHpYcd
OgdVmqxqSH2qtHIdaWCUTsRcchajwDsU9YxQ89KvjhOqSkK5S3dWRvqpfA2G32o8
XvcYXA2lMrCP/Sqi9qxunHRoUaxmXXJOm0P4503LlPtQAnvLiMtTbPcakcCp5vjc
ODai5MPbF+oZge78EJYnZZ9/89mpoRc7CI10gRxGZHPDQB3diboBvCdk3j/1CH7H
15fiWuofbT+1latAsVWTF2AHbDRY6jMAUI3uBP5JtOGO7QAYUhDm3MHvpz34DsCM
In01/GEV8uJ6hdx8ZdfY4KedWXddKm9PxwttIfVjjOFUcVb0t6RW48p63b5oshE8
oyvpYiYiksS2iNylU1YZvky4h6Mxk2onFs396a2GL/PgasAOwYJXsnexw19liVB7
Asxa+3AaMZ1fpjstPZpGlYzaSDCoPGUN5rlqwuH97XiR/BB4AMtSWvK/OdOlURIr
F9JcXFTTvvuCY78MmbG9YArKQdHMcf8H0ZRzk9VoYx1EEHzPTGpAqvLflScy7nM9
ooqf0q9aVE8LXwNMA+QLTtwswwSrVRinz6lBPkHBMBFRUaj80c1tz+tFn5tv4SHv
RE5IGs5Ip8JvELtvEnJQ62I0IlEL+SwR6M4SkBpuFr7gc7RRCyON57FvOudN9pnm
IUUqD9ZEJPVoXalvcsDzuBvCcMe7AN7fBoyfGQWRNDQH3UhwinkSE77+znnkWU94
Q8AKs2ecSb1bThE7qitY9raMoiz+CHvyEfSd9bzvbdgh3N3/lj19FXItN8vmjZEL
f960VzXFkDeB59RNxmarvuu4DGUARtlGkzbnAqlYZDPJ2arMlQAi0f3ytA/II4/+
s2DlHaCBpJ4xJBMpmaVshv4LAQ/4iMiI0KZQ0XhgDWAp5N+cQoRLSj29nvaoEwG1
dc7ZEOxHtzf29PKp2Imz16CSpB1cMZ9vbncqEmJJlPjCpdrXXIHC1wbyakjnNuz4
XU4tFdjOtcBfBft0sI7xK8ybFMVwZ784nvApBSnOg2r/Zl7PvCWYV49p13S1zjJd
pwHbjO7hGBTob8e/nzxWfwEh0P37Ag8RN0eQZQX56vfWpnZXDK2/LFVKOZ0RhH9P
+Te7Xarbcc5u9XeB/F88h4AeS3V4+jx/zcfeR1LEgfACQIlklJY+WOSPRzdO71hh
blalemjn0AFFVmWqxnxKFOB2I/sL+maRNrcxbHxHchxYUdB4bi3FkXAa1zH+wbzC
qReT4e1Z+JOw8WOxHeb1PYzTHXV6vqVAgsYR+U95JA8PYqWkPVr0UdrUkTV7i+WM
yiLHpY/9rJjacO/SdGyGnEyRaN/fSOZDvdDTOrI90UXV9ojPELJxpVHJ2zoA94Ff
iN9VwmherayH54jL+hra4X//5kwyoyHKka+Xq7wfQhnW/O19YXdqJJ7PYZtf2Y7g
nMGZPOpcMdzCkbVVQhaoy8KyUDhWKiyC3FaHlbog6lOSHfDvcsdOXX8pSiK1rhcb
79kUc6GGjxpnie7RUgHUw3hrrqDOgXgT2eyWVL8OZ9F+hbnb9Z4ysy9IBE4b4fKQ
O9TSD6L2SxChu5Wx1M0+R/aVeUOUJ/bqVJgJe9bX10As14FlNnqVwpANRAsibtqL
TxbhXbqIWBi/RSw4F/5NT5d8LOVtpismeJaD4Wtl4tOTGFN0YN+R+JnXfmHaRH+3
Dco9BZs3no8PgZOX6P0sNK3uAF9yIWexbcHe4AoEyczLUBxufbJYKQHxgILw3uHB
cvY96TJQzSBOX6ki5eFL6vAi7x0jzAG809JkU3PJajau84H2Kfx9SJRQdksxHMR9
yKrbbNKCOrV41xWmAX1HuFhiuuXRJ3vsrX/xdKn0q7w8aEVOgvM68390Diod0oeB
4j9n0jc4xJoicvEnNzu0fXTaZGUl+KAR5HnXAxGM98fWt4aTQF9djd0bNjBOBbow
lnH88cC4Wexg93HGBKj1DL/vj8xdhyQbbG0DiPEiSkaDKGdQMDKuWS86m0k/bfyC
nOvinODs4bATp3rLF/hTI5oi2YuMg2ms66xn2RyFPeJtQTaGEFJ5Q8tLv5gALBJe
LdT/K+C4+iygaDIVgCyfAk/cUMhfUIVWjx3xr/wU+f3PBprKNCEutTEkvSjRclUl
g0xM87QL8z35iPm6ZXna8oOFIUUiTeQD/hB606L8nYwbIgrPeScUr5TZ0I/b5gxm
i0vrSV/UKd3UuE0XWEZS9nDUMi9Bi7Y+f+V2CsaExndyXtr+Rz4n34wBtnI9cyt8
zJOCv1hu1pHRAtuDlefykKK8uWMpUwxlN7loAdZi/FX/803LpTlWQ8yw1qmyAzAm
5sq0CGlqPNvuJlrvhNcY3DUk5sRBRZBVr9NJjVdMYYs+RvWKnUEqJDqTmWkLSQ8S
p6L6SZMmPE2fiakViBv8jMehGYGvmSWpAF5egUuG/xORPmFtliJvrPya0G/Tk7Sx
eRPb6zAD5+09n4rH8UlxEQhw8Z0P/qFrp0KRgN2vycT2JajTPTcREOb31jXXoMx+
39cvsRSGrb9TItFs2LTWZZFeSbPbPrGm9BpLM4UFF1kS1OxZ8enBAzC3SoEw9y+r
0V1i13Rq+hdnzMaSfnajmnXco10ZUM5b3zeYKwvsqjfvsumCS/VLxOonEWYTqqF6
DaYWBqwwz5cWSmRwO2ARB/J9RnEN0GwY0Qlb0ovPOHIvpCsZF/LHZWzMA+oJwJKx
limCWq6DcoDWzL/bc0zgwikClUeKKy7txwzZ1fV3FlDj12O4jfYQADSS+oVuZxvV
642xzHbkzVrOEdhOttNHlybkMA3F3RuxwCtGk4RmwK0x2XOIlCyfJZ/4/VRLc4xA
widOiBv5KhSOtMpIQkURrJUnDSgSVyx+iUtVNFtPm01VS4gASUkwuKdXwwt3Oh+z
oeb+IWQlxFQN9W/fuS4m4xjg8vCjDNZg7Wmj3fmlcovi5SiR3Baw+YgsvwxhoH2s
rn6FRSjiGhlpf/PGBAz+l12vhekOsQ9FJQH8KpxBPMSJJTx2Oc2VlrbDhdaeHHGX
MBG/VALRwHIBFgUcOq14KVvbdElfN2BUni8OcWs8x4iLV81NS8Z1h8yGip1KYcTy
Y8Nb/EgPP1qAm+jALRSecYfX+NCbvOU/VfIme+okU6zMXwkrBCMQNqNxoyLr5r0z
POO+sZZpo7rFFvNJYuAd24Eu0VlV+bdIptjRMR0xgs8esGle2+OrfomqCRX10uMX
jY9R1uYRbZDyrbYlPCoHA7VkvQFiKofVCim00rJWPgzxbzK/c9zeo3JDBKfcy3yu
ZYdvWHlbRX+kK2b0MTpUvdx5wWZ/8AffAqVRtUJ1N+ezZclqmZVtY63q9lW42Nsy
Uv+S73mEpT2hRBsvaUw+PNkWCf6+n4wkiiZ1Ryfue6GVVjaAzIBd1d2nFWECYCwg
yTWuRU33z/owFVDwxvAOY+KKBTZMqjDAdzC8vdGNLEX6Da40QYQQnTShV0qR7Mnr
iryGiM/s/IIRDBRsp1z6942SZYWsUZxg+QopHM+jndVTUzsD2GUQrUr17ypyvca2
A0dymOjTGRlcbU3kHUHZBIzTkqHwnS/SDcz/x6kU6wVbJ5w+CyM01HPvTCmJatJc
odLlzWuSoGG19hFzMWYM9ThOML/OATHzK0SK5O/HI7SoHpyQ63EcCpWZ/h2Hc71X
KT2ZQ+gqUK1KmBN7YxNEGsWuRLFX+ZofJZJh1V/e/RB8QSRj/dEo+9lDc+aEbxrl
YJJ997FO2e4yK/NO0B5NJkVY5yO0tsrlcKcdRJXX3G81MH+SKNGy02khznGCfeEJ
56CfPxDkqXZeF05OhYMhne5a1FbHcmUetQlEGQCqrzf1v5rEJWA0PEdRUHDcr/JS
5SRHabbJ+MHurmxVKaYGxojm6piSSmeNuJVj1PyCYGu34Y/7Ikueqx9GV2emfu2/
rWK7Zse7xK9Zv2UQwfBP0terceG3gHjtMb9no5aOvHOXe5GvwnD8hZwjJWrTQOvp
xKHh+rikZeYHslCMp3LIRQaP7jgn7eVfPeYOmRSg5nzH8l1hqpBWsOHarlHZDVay
PFG2xV2Hu2xX4j1vFZ8mXzSDKdANdXYnuKKs5SQPlfYfMHB7x2e/F/vJXVTFuknA
yB6LKyDtZs9HIh5fgbzDUQCPSGdAX+BwPNPOmV/Jo1Zj1G2yn1lBZCrcG9qc8PTw
Q19U6d0inBWCAEUcoaQZLn7rYLZjoOZiKzjElQuPihXtXSDuMpVSsx/buihpEoX9
+FMAht18iYLnxwusTbWKwER4gq+Z14n4UKTYmDmIekmOzGD+x/PB5rxdCN1Uy9DE
hYU+PzWHeCqnXKbCmqAeKCS87/bk6mYi8AbWPQz0hrrrYZejnw4FdIcr9xl7t642
po2VLnqSTdXJNi2oQHjlAOkHfcwSX4AgzuYLcVyX6E2VS1PJ7OIGJFq8agI9vkws
UfUxye97GpMkW/NvZFaNpGkTvM8GL2PqwT+c6MoMoHi/sbcMRZ2vrPKEQg6yFpLc
iPbRysQJSiagBpnewuiI4Mlqiz/HMzq1BAweJTgsjOquhCzyxlbYuQAcOEOt19X3
Ix3pU6bNwh2xMlWQ4lfGykAE7pt44E4O2H61A/lLxQ2XysMqjndJxSeOfTi+Mv3Z
bUcR6AMSWjbux10lR8djB/Y/insvRBwXBap/yLDeEpjmMl+y6G84H+eijiOPPsvk
/OuJhirfPf8dhgiR6Aln0igFQjzMnCh/jdPFrkJqlKH4pqQcgR4wpuK6/O87DSeD
eIpvNuBeNFTRTrBdj5fCEBH8p5lo4UPKQHKAg9S67xawKUEOZr2Bh0LHkaV9E+gq
L4p1JxSDHW2LvfTgEb18KnJ1l7vNmxAG8mgfPRYK7CJ49NZheg6VMS6ssvmfC2Ir
5iww1xL8Wt+FLE47TDZOAc99p29L7YEyt/Ifa7hmMNh6KwLfRsh/969owHOl0iKd
6G3WJtmpnhTTyEbiZRdCvjs7rTCtAU2/Ix1Fbt4J0aKXDAHgvTO87TvqXZE1mOBg
HFT4V9tOa5tydbGWKdRWcN3R69eJxLWPkFDK3aGFQEOSkfaI/RJoMalSfthZ/tDy
ZOtr8xm2v4FPyD4FrTomRZahp6egCnzRTkS9p3i+P949nLEd8jA2lnmc3KbepAe+
BrTQjuLjXVSHrZ/6K6eTEeQGvQ2fHip2vNDHaHUovvOtAuWHHUGdTBLkAYOsT2+u
lXy4gn61ymLELCS5xiwAgDtzWr915wbCDt1NlHjHO1hxHMGL1/kc6d4moSBVcka7
C269hTXezH5yWb8roE14jONEKoGjf9YyBl0zhqwR3MG1JXJY3gRzQuKN+/FbYIoY
8l0CjgrdBxuRQIoJGYikczNHZJkyduabRSGeFC2UqD1JeJp+1RnD+J+UHPnbq7St
3M4eDHlkguaSMMFZYEkoCSIyWTCgnNWjye5wcYNtQKGmoVF5cM/cdvrc7iXXFC7q
hx2uF9lheAC8CQIDTFrRuBVrLxFma/FCs2q/TiflhlUH8YBzxtqvn4WKKmsNbZHL
Nge10E76rbmVLHEZGTI0B51ZEztGUeHD5rHliGehMRY73UidVXEwEkksn7LCqPNd
ucjZb2RUAh9vciTmi0oRcIAz/NWy4W9N3siHOoMrjrG41SYG+pKRo0tVc1Grdh5Y
99vNTZ4nwuifIJP+2BWKt0P/wj0U3bbo0furOxxggrdmnltXQ7yz8dXtKZ6TKe6O
dKBGUpmWUfQVtlS7N3HunWtDugFB4tdvm+vu3iJhOTssKL5UNgoPGqEWUCNvZwvE
Y+VxO3uVMbn9E+60jtZiFybxpaCPEgSDKgzM1bXZ/EEV2QBoOciYM068Go9O8Lfn
V8P5+OokNzyPb18itEFamww3vV5nfeR28+yv0FuEiRxoO12OyksxqRmUldIcC4mw
j06IEJO/otYWaI/jqUzp28zfjxj1lyG7FgCesOhh7fqsYEsYr1Jg8NF/KDahNvUi
xll87r7jjAFNP9GOjVwmbEBs0TdlCyIituQ+ZExZLikR9GFaw8knRTraqiANrUYY
9So+BjyHr67uWW3NwNNiDSK3SjOuFMdh1HPvnE4l6NHw1bPmUcXyNqLtgZrby0DB
klo3dF49UsUd2NMBlcVZErx3SDcLK3jrDl+vH2x8/sC1npw/kixs7XsDS7EaPGg0
or68bLWN4lRjKDeH1NkfVlBkRlpUhU7CSCcGsYNB76MHoecL4jUSRUr2eD/hGG0S
S888xC08i9k4cqEtg4tpUBjABCHyg0CPF+CCj5ayKaahl3aJ63vLAy68d57NEE0S
p3TYZNrF+DatGR0+yPqO8ECU/O879Y7TYWujQIsoaZZ9A8bLjdN3+y0L1F/Jhs2e
agpdkD2MnDegX8ZAa04iaT2ytFq2MmYErUPJzJwVe7RUhYtG0EVSebn3hGkiNUUe
4FoHDIVHCjh5YNAEYXdmMeSlyvVDfzIHNK5Y5t4ijGfUGd2mlnLNyd58GmEpxXev
OsbF8bFJQhoR4Q47c00O0ZZh5w2NvJyg878ERcQp8toHBFfQU7C0+lcW4arMJkAG
pXy39n8+guJ2K5taUj/ph41nlRxIhHl9akb+3ZZUVQXaJHi+DQUi6YQbwWCvNx3u
wObTQ6+CweM2cNJnu/7gwblqrlKyBVEPrOp7zf8J4o1TQxdnlCRXwALHaeXumPIr
V+5dopkxcrcUhBU9ZtNQYGtZY0teJsOvBlq+44fm3jfZRWofFCFZZ8dp8djlkqjf
Ox1VQGKLUbn5KO1IqisjBeRIiMPnFqgvJHnwieITXY8cidx8AzwzIoiM6dMeHRGY
tlK+itwzKk/b3Z5uOLUV3VVrPCOkaLfD6Qv4yS1LdbYYBBIx9E2w2Xyd8lYfAOEo
XbBt4ByzPQyX///S45Ew++tvA7WQpf5Mw2dwTU7WH4o+gDurEnREzvXQUn4m96wD
7tdrQLs/R8qlbx99tZLBJB7YHySplhbzQTrHaIZRMiujiLA3oFRKZfjpF3/Dxk7D
9J7nECFpX6PRBhu7g3zNLiYGzCYuQC3JVS0bmRWv8tgSrPksFDZ+BFy8D8KjvsRP
fgbShzDr1QPfWg/uyDEMSvKw+7U8cdN6Dk4maGzaH6VcKKxWtm9RDbQKtCuX+L3y
jRMiXzGs7QLvmiZj8Vnasx2FcuKjhInqyE+CkErJkRxAzIMdSutLlaozTWnq8neO
5s3ULliA2ALIyMUu3Nwtvf5fs4uUvWMEyrXB9ZSAghYTm+SNAzBWqWC2OfZ1hB2M
YYISYwns469I4FZTgxn8h5HQFwBkG3ZGDiEJX+hLfLZdn/h7mBbqao0jNqcDrgiN
QN/VbOON/wqW6tk7SFlx+dm1ZO/GIt9dJj01io+OXwjuAGWbX0TZ2kVvCO/ITXFf
Jw+tjTbQT6+tu/RgI0QRcT9Xv/Fb5cMHlUNYl7aYtpBZbTXVQV1E9ELbBPlqrKu4
E7k60AJNcI/zQpKVGG+d9FJIEuWBFlF7S7KQZZwAK6O0bfpC0z2aEBXJWSyQgKXW
0prnMklelvA6Sl1NycWaAEZIsNyObSq5fbX/qB/kb4KkImBHrH92eodRkGRFnNKU
mG3zl6aLcQxDQSeuEuaG/rfg9SFBfmv86Om9RCenLjBLWebl7U1hSeqkrts6uidG
3daauy3dljBJfdohRBv6FgebGJLGe33kLlfPZZ6hcIqfiZdyEWunP9U7+ocMU577
6sQNbWc4UgC0HUaYBFkMeoMszRoXbEK9x8OtuiC4u+6RO+/L7FQHPhEoLLDGN02U
P159p7IdOnLHRe1tVo7Te957b9+GxhvcTopjfj8J0Oq5QpH3cu8XSncblEBUAtKQ
WbQF0rJPFVU2YwozeaEAyQHDVfWXs/vtQJaLHtcmuBGKWntfT07nsaxHQODMoFep
biveubfGwM/jZ98FJ8TKha2aqzDpkeUBjhhr2VcAokFh4adiigU+ZgTZmvB5gdxa
BewTgf1uuJX8PwsXwflUYWGBDD09Y7wCXZ81nblqDORLMlHg3ywuu0Co486jZLjw
xoTtk6h41l1E0gkBBCvUOvdqltZRjQB7RC2Uvr7Kl1mf6svvy1RJkXLTQoGloLAc
qJ0TiUIMl7yhsHPdVEm9BeJ7+5Vhp183UkCM+why2L6fKuPLkjc1/23Ue5bcsX89
PteOkKWds/ZdkyOTijJBXyX9mdczLY6LzIhhtjqE9wbeJ59PcpwWCnDBn42jEzOx
GVGzgp4UT7DYCYqWWVZJE1uHcop9unUNDqU0uX6AV439D+9iQzlbpTnzmakrWVks
aUeXhxjwe/XZ06l9/Kv0M+W3AvN31xue8kDhEoDid2zBgIqiTIqFkTVFBk8g9JjY
NVoSxcOAdYJOV+JA2aivdUTuBi9b8u6Ivgk+ogaA9RtJoQQAMohf/d7/RIqDwcpR
40Y5g4UpyO7H/z1N8llyDP1QKwJoxMwOZ6NQFStm/pmABCpHMLsMz8P0N2C0f3H+
kCc3TZ2T5O3BFYHAW9A7b3OHZis4h+Ps6DGX5uE6tJ3V+JsVQ22q7CpLXTwg4gUz
25VqtwrW3/nbB7IOT7cJT22I6LiGcVOEzQi+Qe8NQry1SbYKmHbg59fD3odfurDo
B4HVFOBHpPrXpYM0BF3DEo5xNYPF21NyJ7gof99K3mtz3/ivnDV4HSwbokVaPoWc
nBL6w6VSfL1NJAxSxJVo1sgYw4MoWNUKBhxFrAXdXPuKk/fiX2WL8aveQCUp+o7x
XusVisj6QH50xmj9+V0FukVug36asB16gfD5nFSMKsqd0848hcoz33R0nCM5kh0X
sbfqImceevEfvaIs7jzKa42ve1MSCh4K0Mylj95bUwTawS95pxCMscKUXQW+jq/r
+CQiLFxXbzdzVzxDWFVBwaUny1kHXtzLF3kDriFVzNXa3x8ZTitKZChI3nTaOciN
b3aNfG1hosuhDbSM4UJ8drrIl7CPEv/MY/T2JSZjbpHffh5tfNHRxSTjPOh0bx7Y
MHNtg375MurumwrIGRtYMGs+Pd/MInZHgHl7ZnTVeoB7EPB8/abJ8o0b8bkv4DHY
TKd91imlaLT6TDh/pm+exnt2aX22QsicyaXD6dk/nh4VlwhLGT3Fi44MYex1h00H
vgk7mIehpm1HsOhv4Ew7/HGzlyk3H+FerWqiMOURAIjG64MwhEU+1s8YNK68ectL
oT9K8R+8wQB/gliqGP9ecVHfa3r18vXYbm1q3VzBoB0Z6VWgy1EXm8uFM2j3M/Q7
gLXCaICALJDApQxWBux3ma3mck1E5u196xJNflb6g5ovCJbU5CcVZrSTTVgKz3gs
dUzcUJ+ntBEUbwJxr5Au1QrMsPPv/9DSQufLXsa+zOjoOpYUEWVRzmX6HFhFWqUh
u/hrcjutjMF78/h0Z2J+MrcHARbjNlnlKjVOF7BfeB4VG808uJhV8yIjOmueM/7e
jDKpXnX4s4zqBCy5ZBSQa+KoXEx48WZ8lLrECjP7fihOKjhgIS+BY692T8tu4OC8
0bTmo/UiNbSTWUimaP6gkofzy8rIoC+kDVuOlQ/2cTHBTCsEzeWmTTwwLK5tEoLj
tCi+KIw+/deYkinCxuH9MeUFFucxqdzLqzR8W0YAHAcxwbkNlBLRz3V/MbLu/n5n
vh9X1KmV6w0cRj93r6z/nuqkq0QHRJx7AjP0gnzpEN2XBOoz9cM8/etyXRxNQnPU
iTcBwW2UuCBthshUKBJh5HNJ3kcu2M8W6dQc9k/FeKAPx/VBFKf3kz+zEiN94S9/
9jlTLfLViG9XjVLdvJZ2fqzNFaKAXj7R/C2+GP2ORDMiJbYmQ468Qyw2fxDRDRdo
pw05jsJVl1bm//ABwouVaYoJ3lvf+Ppd0pLD6WxRyABs5npR0INFilcIsozhSBvI
WnO8M1iEaI0afHW7NNSTwqZorMY9kmQGQCTJNAkhxEFB2+P0eykcIDG6c5Y4qMtS
PFPDdGkTMN0/HcHEhhlKJLg7+ked29DpnWCDxOGAlxyAfOYnMDYqO6VgAiyMPaNt
hzBlsaisjZ+FvaxcCiyqPHlrgmhUDN148HY1SbkM5kmSYkedBLcHmgul5lL0/ODY
1zSCHS1TYF9QqaB2aPai5qNLf5Jk5vwVq7A9WTQw2EuLHPQ+XJW/tWw4afUTxDZT
bAjjFI4zZWOAbdtZdVXPDhA2XqwnZm8VFNhLUDR+mKUTnPkW+2GCJurWwnRvT49K
ZG7UfAUsYIDRbLlg/eiF0suyPZK3Nven2a/rvPWxuffziF7B9WxhFeudar2jpjlw
RphCVdPfJSUC2JCzZGy93UlwrgA6cfQxMwvDeqyUNQO4CzlHf9AGY8QeDrbo8+b7
BitNiAWZeS8zO166Lt/reQ+rPS0U7BurT+3JBjqbFs/cF10EMGlXNK3BJ7mV0Mez
QqrJW9AWdv0acmiqEcx2jwBujFEubFDY/YSnUIJXSszMsTyNnfVfUfpiRUe6gk7v
tHuc0b58zj8z+bZKo1/BkjALxdkDx6W8NaWEsa7JsH5GmL3wRnjCkLm2L04biWxH
qSvmunsHwuHL7+X3rRn+hQqBI1/XPBRUCGKp1UkZk9plpK25aQ4aJwCFNvh7lmVv
ussOfURVuC4xOsZ8HNcPIFTqx8VOwMYJ8TBavRLRElsI36agjZQHkVjFGoTou0mD
H49SP4r9P088kBaRrhpjJIY38Jmbf4I+FT8fKLILadf8d22RI7GOQogVXv+PxyyD
Ru6hR1O2YOZJPNwPCTmU/imU+qHZUxjaIGDQP/C3eKyCU/6ezZLKFrXCyM1Hqrg8
nLirmefMJfFQLuC+2eEVRJjiFGgbdvvcQRQRChlaMDVeD7fx3jx1FcA3I5Fva68l
kQIUkdRExc4HDU6qhEz9NN1C+S85MMt+ofMWKqnBqjlGYjmZp9VE68QmpHnBzcz6
OOFHfOgQ26xcbm19TK7G2wclY31JFF8Qw2g+iOCIXXZhF5v35wGxiSd0gkX/u1v/
ksPbQYNEy4hfgMJgi+SOCum9hMDknUhX6frGsAVxtYRIz7rynw6JzFfXBAiB+8mD
W3N+WUIrNF5e4fXr8DqKMHZnL+x3CNx39PuYJ3NhdS0hfJH/h0L2Ctnz9i6s3nwY
+/yQg/Lvdj1qf4Kqce37sx4T/wC7Kvgxo96H42nOQXpW924tbigqnmxFS5Vxid3+
CxY7AWbzLiaCnQc/wBHq5k6wB0rj8m1XlbOKPiPz+TMybnHPiPHmmj2cZ9ThL5BY
u0ie1tY4LyaO8qRWbxmgZcyK1uE3rMHAxXp17FjDLzGO//3rhHgeKQde663/rtdf
t1IkonWLUVs3duR1sS4gagRtb7HL3WuGOyQipOiM1ZYqgEYlTlHFIIPtYN0W3rFy
5H1Kk/hAfDhXogCNqk6nSqu78mX/yNM5pw+LDPWMJ6Mhssk0RPK0/UPObjz13vL0
9haJzdKeEzc+nPXER4xHV19LVarYHUwkmMJDSP1+vhbKOJMuwfakVz8n41jStLJ5
3ePKo34eM9YmFHiqveeVuafL7TDS9O+2xNjUGBoHx3JyHgcL4WF16A+nBqYKeDzj
22a7GOhVZJj4OFdLdGk9idk437RzXoAe93/ZZV0DrhyiIPba1MK2hCqsRCwP4Tay
6qJXISp3GdsVRvY/z2e8bDCxS04AwHrlKgibb5plBi8pYnaTwxhC9FtAguaFW2EC
kNUyX+Aa3OFYPBXw1cXDbX3WRaxialk11wK21VtpadvXR8qISsYh4tx5w/WCypIr
AHYoadtYXNBedbBcKCLJ9TpRIc7SwX8+JQPX0EYgkm6jqaJWkTBJ6Qprq4QfO7YK
qt6bCFoEY9vYZg9QK6KUPU3eWKEjsrYCj7taVG5l9aQ1cMGlTDt7NwZKAgME/NQ2
gvrJOhgfmPp3GrV7AGwTKWgFAtkLGiIdBxrxCvSdofcZntgQXizMEWMCxSEk6IKw
BBlNtSpj4Mke9cnYkUTI/CxG/6MFLYG7wRmquV5xMxita0C/akOAQyB8RL5bFOnx
EzDHw/p3wr56ALKsKNJB96FJ03h9bVbSlsyaV5WNhveNL8TdNA/Akc4dxzu9Nr/X
ljJA1tTRwPS9+Kj35/S7T/DYxOBW4eNwVqm+PejWZe0XC2VcfSuYUs6wDZixLTps
c2dlWLgwC5f8I39hN58QhjBjnIHKU5vO6EezpgyPi9IhUvQB7IX6xd5VS9Ccp0wj
ITDe68svHeSYOXb/7lkPDT6T4XEgLwm49fgPlwzQUKdrYAX4EBX6obBYVoso4tVG
WvupfnneQ2N6xsSVmke1HDw2BUCMLkA0uLpPo4K6ARAwVGUIV9WLDHoV0xyFMcur
OtHYAlsOflGx1xxfcV7Xmvp999ArJO1Bn4mYOQruLHA4HqrwdxTi0XDuxCHCBIrX
t5+tizrh7wACBBwoYw66P3sIJT6ooTMGg+G0OjH11g7wZlqxBW7vBL/PlseL9Mfa
ecqBRB25qab+GlOqjmgMjT+DAxiUjQe6hu0z3xwo1PIVQQuIHp7Cocq/LHOjMvgJ
YXY0GJXuYp5vIx4fLUv9738Tcf6y1Vx5Mx1NWEwwIMQWvql4kLgewiD8TdBxm8jk
kHK4WxFPw6IwOIIy2mQaYyghUurWKzIrJWguykGgBRTDIfKk7r5+maJzjSODN35N
sX3BxrdDEty0lBHba06D7AE5APCfXa5LxhZ46g0QxbFv/zKqUlHp3NBjTTJhf0m5
kVo4It4znklpLkuDhbq+aAINkEL/Zl/j7L3Fx9nXmynrPX+YMmIRxtalWMNguxeb
mg2eTvYOtTpkF9da10lh6XZkU4JmdmWioWHCLocTrh8u0SRTgZNw/ARd/A4LbOTu
Dhrg/HrO5bDjNzC6FoKNP3E1Ot7jUUn/Zh8dSEYZ3ODPvFq0eG9mOH8TMqskC4o/
swAToveHPMWN5Mj0NdLX/xNEG6mLaKzHecdbqouFfZxTpXx4N6cHec/Khsq9g60h
IQh1u8vtYUlMjnKlKhEaOdNQ3rixu0sewu9mSlxuqKS92MWYGosyKQkFzIb2qD3V
RkbwgazQUkZ6iAtUvcmTbxW1rjsdX6BqnzSxyp2By3OP9baEvEDFQjn9dqjVPfFo
znTqe5uXlE9O29NNKpMHgXfWm+cEkm2lp3DWk9mR1/XmWpGAvmIzLQXbb/hv+L1R
QepA9HCLVnn4T6NqMoOxACMq8w7Nb18DQAYtJMVVwYIdnefm+sU56uKzT40U+z2h
8yVAMSX4T6ayqfXA1p78b1S2pFHE9NVghefxp7SQpeQssB++3oLdV7YkiXtL56Xb
+IWWl1ua+pbtDewW764xWHmOCflA4bVngDiZoqR0Rn85yy21AHYwgiyvhxYXwmiQ
lN5dINjQOGjCyEJMeHzAN1rTIVv3Khgwg9UBnd7I+MB6BNWWpa201OPtSy5N1gkL
iTP1U1kn9JMRKWspN57HGZTumKS9G7WXbjYT9C2OU4mSEropdNyWBL+MuxmgqLpW
RNGSNj3vVfSgEWmOTYEYPb1q9FyOl87Lr4wJvx/InujfquSUtRSOKjesdaG0rhfJ
0yg+XkF4G2dS0EnSIw3kTHmZhdjOpjeikPsbTis4R2fWOEU/rljOuEnvrQ9RCcAQ
tX0XthMRWTl4BIWeDOoyqWggAW+55AZyStpl+ndpWzIr5+dFmBADc9AYL0z3iZF/
4WEouiAhn8iT6ZX1Th4322UFXCY9Psc9dn8+SoubeAkinQ3PH4iAQVMf1hCai0ar
vbCnrzhcBVsmt9cJCn8pRunllfl3gHQz2kWzoSE4l3gHuwdmQUZN4t2P6BP9FhT7
aV3dxft5AXC9E6YzyxJSmfloLmHNmfZyBS4QCYRCiuxe1ylXEXL7V2sS5TvVr6+i
NzGaFhis9we+9Wfe5tPlbH6Hk7F+G1/T3348BmtAAxoQUgGiY81JYr2748Ht1I7M
hYTqwjvOIULqWDZmKQQdV/A/1O6S5J7A64A+xFpbbjvIojXBdYFx2WtuWY8O3wZh
vKcbeju+Lw8XuR/ZBbcFM3O4n8oR6X1d3JbEoFh5PYwLyL4f0e6HrwQCMoZ1N4TZ
GlgWv8xSPzCNKigCvjuEqAVi215/1iTikspeoi35H5SHDVe3EenLZ9kj0PFC4WI0
mYQ0Dh+kNEDTEx4/Jvi52t8l2836t0hvhrinalAu7cJF6Xwi/scczuuKv4HnIYOt
+IYulG49erV8zAuKyp2rrL8fFz7dtFuDPvzOj/aD++qwmO/ILCfUGHrqRRfB7+HD
R60b8hMLsaJIlnN31e9yJlA3T2vJvHvn/msfstmch+JvhfdHvk7AOfj9NCjucvJJ
jke7qswrs/M5fdZBPtTyTYP4E3bNukCNUC7pu90chr/JSNqA3SW+05tcsSQb335F
GJEMltVMoSJjumhJ8uojKgoNvuUKFc4bZifSkFSoMKEFeqGRHmsSJ4P6yQzZMyZj
9GvLqi1WpBEY1TaZnwzQ8hrnNBJUSsTt4bKXpKqS317BLL8XUCBrfHxxlJUT4u/R
X6k4EKKd3tSuKvmkOnPKp8KlS5ceSEbABlsSUOQN7gEpbcnMQx0C7xXEGrnhL16x
PH17lE1UihSmQwvFS4bh4JfR6cWIaj+7RNnfTs7k+0zZ341VqjJEf2KNjPsBfF2j
FBWdJr+CwWFrrg8U8U5YY5gab/cCzLbgR5N5+4vJsMPSOVBta/1IgW7flxB8bTLm
kFZxE0bBq0i/ZJNX6k2XdJqsL0K6e+SewSJfI2kWjwZhwEP2bM4nR9y5nqDZKS3C
3HGwg5jFzrVBnl0DgOkh7f4tGG+qu/SejDJQXiRz8ZZjilAL7sBODDkx9mDtGDUB
B811f4DC9nSp5aEolzBFFI4CmVjLLkJH5loC45jYTkL7TAApb291XeZjR6KAV/Go
5aD8iqF8br+BLQNXNLCMWjAeFqX8lsynXxVToAziaAhQDgECaqYoKCzylGUdSPmo
kxvgXrinUwblLbcKOxtYm94ZcnbM+oHqbowfBFHItCjao4fuSALe0k5ootLofTeD
qNhKtquTPWHqdYNxEnsOnlDGs3DeypsrVVESBR6cOql1o6wWvtCzR9Bgae/2WeEj
FkjZztGsfo6ET+XXI7ORWykb9dadiolejfa+2A01pXYIM7z4I84WdaWLu6POKABy
aYFK7HM8+FqHheqw2SeiZcn6V/HpjlIJfJleZbD8lYeuZSwC+yu40AiKBAmq6jIc
xJvnDQNramVRPh0FUYcoPwNI2o21riFUfsmAM59HGY8xIzqVa6GwLkKZhGntBGgV
Tu/phNcAQUolrqaZZPAryZShAeHuq6etRR+7qCVUFPENfwtX/1kvGWmMVXePUvJU
woVN476S6ZXsqhu2DhTSZyF74s7tsdYq91Qgw9UHILBotOeG4FivOjM7R2ptWBiB
RE3pEEjPXv4rYbC95CA1MOXba04F9EdD0UNsCMar6ReK6C2smkShlk7iENpe1Mld
6U0HvyF5NXDAahWyjoPmrZ+d5ZCUlgTXJmkB/ffkZUV4+uuDsvtP1mQoTADVA34K
04Awn5p6FBR+QKJC5YGee0StM0wvSj/mBBjnvpr6mKpqmabakZxjIV6SYP36Ua+F
wl3nE4o400v76OCZscZfGzVuByotbndS2BMEuhJwmfs8rcSV7smuiEMH/FeV1uOH
tQkdDxTXVwyrg9bOIGnMy2JIYM5bn6FNtVkvXdIJRXmDFgNgoroq/FrSykOQRNel
J9wZ1Cz9nnkRaLMWBVwra7UaYWuXyEF8fFosnpogmKTOzh/rrlLxWOpmuz859D74
ZDG7WFDEBfpQ3slKgoFZgNw05y3phq3EFYokiOjQzRr0m4YHM4bAz1X7vT4SVEwC
yTs9ZSoT9iStujzJHjZ4I2XwNpO4+/M81tcql7vQwjnwbf5vhw3q7byaOvRkQqYG
GfrSS7aiVFFrrd5cCUHMP0LYB+YJtvuTULcVjns0ebIrH2pyUIgLTo3yP82gEsr6
ezLjh5SJDlNB9MDpvF9IAOZAtd55O98+9ZsNDfeIIeuypFbVG+UXAY0USnJU7DM7
LtMgw0sIBiwGhtq2Br7LtGp4K0p5zl3WnibrxHoCRHA4Mfzir2zHpBJbH+HrJhSl
MRuxF6b6Hd7Y61OHLUPYmwHyuYO/Mn1HjZV5Qle0pyMcBoSpDm6PEc49zVJ6YgWR
bbLyHDLNUnnWauDRlhUglJB4AEjRfPjmAkChD2zuy0BGbCvYZ9H6cK5+IlAh6NWn
6LlcJP9ER2TLJszI7zQhywJuusyt8WacnR9sVRy+G0LmPE8cBaN+LMzJab92VBN6
FBeo1TA9Q20+r9EG5waiDuh2Z1MQeeeaQZvPZomdxFeWlPex0VMzPdR/IJeoME3o
3q6t7LrdNKy+y2SvYYp4Hf1eCNw3e/PzuFf/gJAzywdraQaiqJbv5tGtlubCOGnC
ii2FA2cO/+KM7k11mTnF+pfwiteCWDNl3sIw8jeYwv7nqIPqEkBcSDskUKVrmays
jCgrQgw5aJL/B8PZzqV5MiB0OEVfL7Yd1Dw5LXfE2IChc3SOzoHwLNayznmmGM1T
2tdkJ6YKhfJ/4Y/q/3ZDoTba9PWf0edbAzCdm8x2/1I+7j3Qj861WyWfhPgCP8Fw
DiXjewi+0N0KFXv4xHHXFW7bXJkc/AiR1ozrvDw+i12recjAo9k9Emjfi2WkMIqB
rwft6HDFQzOvE+/cdrXOfKDGFsZ2LcwVyND4kbP7QZiOQaDuu12U8rP+SdjqOOlP
ASVl0DgWXcVR+R2ByUcuCinLh9Uin/nrUwe4fXoeNk1YQIYj/jDDHFCBLEnQ2r5b
gExmoOYTEvYaUuPG5darTRQDRALAKK9ZMz4I76UgqvQ+/kH3SOFWlWyup2KCCgOL
axQsTpcVi7nsLwBbiNh2Hn5S9XiS8qQ/OMK5/s+ryJLy3P4yzX1hldpZ88B4KbPN
5WQaWQX+5FLTobOP2kpF4n0oVR4zsMOdWd14O63fDb1AMQXg7upcPxxnIdfqDS+4
ponUDa60H46igHAMIvJlffWM4AV2nS3tKDKLCDwKeboGSNVsvk8Mxc/B16nSJfKp
f2MHlo7agrxFMyQvaVpO+S/zpvZA4fcBeFFyy4Rxae4KkOATHNazK2TS1oRxV0Ts
Is9c2pt4SCxvMqsdLjcI9A5USUFNhGnVmN9Y8jTtJ/3rWVEc7gHpuwgKylgrqiGL
xxAliZKI9ZNXxcbARX2l5IJvvJ/eFXncWK+Tma5wu03dMZPJNClGUSbs12eE7qJJ
dbUiQH5E+jjubTkhw5+ORBTo+cw6HyT0JMlhl2RNY70TrKslb2S1ffsef09iYGib
YoF6zMG5X9H9Sedcfg7rR7A9mpd8l+OP913FJDwKNcg6xjD1o5p5K6Wq3RXWJSuP
YTRpwAX++rEBQCQBaoIim7I2lUTnKVuSlf3ifjs/axB10La5tLLUSDAkjvo/qPVy
Lm1c7VJpzfkoCkflbyMVL8ajiT8LDvzwhLw6TaXyDys6O9mmmvo2eM9UtGKCqtBA
1djfMb/U7t2wNBh1R90rUnMupnnWxESK7LwU8LzV3dzyLyUkVHOIBC6gn7tehbCl
FjvJkoDThTLKhhRMI5w8fvQo2nz/+sH0cN5Hlrbvcy01x6hWzSeRoW+TcqRoIqpy
CiEeyrF/EZGhAElKhHHmx0fKpZpCJXM1/WwqKtm4cg4VCCGN0IgNZ/cVVdfPX5WV
HdupsWZABI74ma9jpi9OzuuMiF66XNA8PLf1aShMdtIyP9SvHJSNXyBzhpW+zMSJ
g744O95/SblMirWg+taPzBrHRIam/KH9lLUyVXo1r2y9k73Hhd54D0Je+kgd2qF9
Tgc+gn3Wy7IJhkOR5jrybO+zatuTRX3KbkNVYCRw+71QP8gb1I3iTOOjoujXVxrI
+bbPArD4EL9yzKZJi2cFyj2x7cTwEfEUA/3qLMul8wPCWEI6h7LGLiXnKtJClLlI
CetF0P7hDeJize4TcNFVS5pCeeqxNNpZNJH0D/x5M6HL+OPqQ1ktG+MdeJLo06EZ
247ES4J8kLq89pDu88UGo/at8GMuiNju5W7mEAT6x6yfRiLWPghQmaUxgfUGVcPU
32CZIUpPif0YrgCkFNJavk2hBr/grMMRhbLBrwDR+ykxxX7SSZqV39rvWbxAz7XF
g6QZexSBMaCBfileIQQP+70zEqILhJzPhOcyxgv59C6R4KSYZmOCLFk9R0Y9r60p
w/ZMGekS9+cnH68gm0Cz/Jkdylz3n5fm6skMjBaR/a3aD7NslYDG3UrbPOtdSnS1
oSaq3HU6Y61zbeePOL4itB0FYYE6DX6GlXxyAYZjmg31e5IrCqsn/muBe737nCjl
pUdOYJ06ZFkqc7qNpQ7g8JzmccniYmMfn4hAz7Ka4TX7SpGh7D4vE9KBMbgh5Jgw
Fdte/gNTgHVZNMvUOA7/FZNahS7/PyyWbZIh7hTBCbvKGcVg6E1olTo8XPEvzj/p
r000S/LlmLEqlHb2E2bcbS+Y8fHlzvilqiJO5cfUyPxUqpjI4rQwQwu3GWH1tri/
jKaYmwazXxtTxhTT5FSGl6xgofxQzKP418y3PJem7JyE/4nB7BdxA7LmYXqWgw9P
5Ao9+uQ2FrplKWB7oiHUkjb+37TnOZ14aGYqWbK7zvFbHhxyn0LugRiFIkMLByno
18czpGvQcJwBzQLs7v6X4LYlInnm2AFCmB1wX5ou8jxyuD5KGnH1zOstf9RZZO+8
S+ZMPM3lG1N6dtSI6pPxxJycqn5tb91pBADdqdJG8BAyiFGKwSBi4My5YjT25/7X
bDnUjlYL0q4LDbbtb8E2qOQzzpUB+Ui29Wi/Nmo5BqSjRpntsDE4LCvTGc6kcLeB
2Zhkh4o6jrv5AKQpycjrvLuq17e6jIDRCnfM9PwLROdfGmadEezSYag9M9AxIihv
i30Q5BNb4XsGgMjSgmFgQh2sesfNE+VBBHF0oW7e2fg6c+e/XJu3fqN96FNwKnSS
YsLwZy1yv/cFT2uYt+uOEHMjlMda+fmKwUKdCBMbU9Y1Wmb4HkiPrzePjeYRUTuQ
qBphAV8hOZIm13LND0wl7Tg4VKi7UqcRJlr3NvkM5aua+S+w5JGnKwRLCTikKR9H
4frVpxXg/hf8B15w51CkD/YlHLIXzdLMJQe2S/rU2qLPtPtCiTwoi3IJzIuOOr1P
vnHQl9AnMoQTg0iIPF8VgzGlHjQ+WI9urbU8bxsL3xvTfqBQ3Hl+bV5eYUIgQHGU
bgn2jGNtMLqgqr8vZMwa0KG+AAe+/+SrQwrpFKk3FuYWEOqAll71eeARoBAiXAsc
PldsQ3QvS+VAenHGkU+QPhBSmOy5psmHGRGcRzaQlp4j6rYhslwFYPVB2D6bKqvm
7yKVANhcVOrH+jNu0s3fZt1wQimInKROsIrrezGSeCdRhX4jdmdbQVe8SyJWt96J
+7Kt+RcFGZ60vhj0L4QeyyvD3Ax8TFik8B+jomZmcMXESjLKJm13sy/Zn+zUvS9/
U/NhfBAlwuF/AreUnWkMeJJSX20BmgFsSh4x7D27kdH3w4YemmS4Rbn15aDYNkJQ
eDEIn9xdrZh5ukrX2eZbUJNJ4l7VWab9g7IdJZkpb6z+FRBUL3gIwSdbl2qYROVq
/pcEf/UIH+bhPtGKIstEkP5oGF6A9pOla2InJjX/21gO4KMI7vgk0sCPjlEhKRXo
0qa33ypNw6eRWovzjJu0+P9uExWmwhC3RJb1p0vQfWQDzWbdM3Nm+rjqVv2YImwW
4r0oZOqoFZTAfqlvnSPytMeVML7oXpMqtGJZ4ifr6Lm0X5E2GoKI8ZN9Yuc8IbEs
pPZUWTDh/D9LYmWqAYlkfIrUgzWp87/U4ZkZF39jEa0PAhbtRYY4WT31M2KqXtpq
TUwap1EEVyRw8G2O3c4zMr2hDYDq7xS4ZQBXEwuRgcAcfGIKrpNrn3cSHHJhPd+4
VdlvPN2eB6R5YTwThgk/4fKxrvrZFz3PbBcAg8ocx9L7M6SzZgZdz3K39xb9dm3Q
yP62IOBw2cvcdz/R9q9+TZljkmb5E9BWXPhFg9ViuWTHcTOTiCDmwPhGUpyv7Wa8
BtYip0hQb0SXFr4H4UPK9DMRFm/0hzHKb1zrJ10HxuZ2+4c4LRA3eW9narwntSN3
fjwtPjai9M3iyuSPIa3KzrgKKR/xFOBSikae9xTlkyDFB0EkEIpZtX4wzHcvJaOF
H9Jh1E5Vd3DGfUnFHGiXpuARMLR5R6uPM9M42cHweE1/J1bcjc+/AXj7xbo51d7E
IvYkLCMe1PGL7q8B6G1gma/HZadA/BOiOcKudazG6tZEg8AYDuJ/awTdleOh/2IB
MDe3hvmiUEWhwrnzsBWXH5OndA4wnOKh2Fx7BGRiwt4MFfF3J1WcKWO3qLQO/P6W
2T9KTD3dO4a+gesj4ecCYHrg+jZRWtHzAsI38zt7iRBEUdNVQqYTaPYKYKI7/35K
AUjLTzexHHA/7ifyWatQnsb7zC9kmJdxv0KSkCpdqOwvjjajKh9skD/Q49UMsJba
iUBqQU4PECVdpE9XWXGWid0hgl71V4xvj2d9A9yn8KmT95HN/xnA63NX6W0jC1cn
+sninqS4F9eAVWcBDhVEwN88QAUE6zrd1qE4IidyejKwsW2cB3Qdjwj185kuzuBO
EGXXIxGB0wSBAAf6d/pvoGxRWxWnnvicb/Sz1BChGh1RWYC6WjBdEbIxiEq/kEzU
aRe9VkCV2k9qLchWRe5nDiKgS+zM/UGofVj642Mw1HkV1FG3i0vU//XeqD0FCOlm
6c2ODD79fzshOckhfesIwtrXiJyk5jq0ZXHp63bKClBYIAqfXQ/4LT4gWgTpEIur
/UEvFWk9tleij5pGlbDpZRGgjqD6eiXn+m/9RR4LPmhZRG77OQjPiraCIkLslQPZ
pQvBjcyzPJXiyCrBovFG5dJyENyYS0QL6RYkeGaMT78RbliM1ItKFpO6/ab+QVw9
R24VPBTgGaSjyVDGMf7+IjZ+8FlPZVwyD5/TdI49SUC7K8TEh0rRv7wkTTkALo9z
47LLYI6S9cbsKAR2E7LepRrXnwurBhe2+1JmVYhAkDElVW8RdimAlXNHu9PGzjx1
OB2ZEGFwFQ3kEqQuPRAB5haPMbOgAqx3RmFfmzGSuovL7gJObqHJnQtiFZq5lfM+
SmWrBlBNas3iAOeHPG8eD0rRv24dLKoIBCN+i5cHDYRP1IO66/vfXaxI2cBiml0P
krUNNvIId/WjbJHgxxF7poJm3JFuDa4/ioTXLxO6r41VnnHuTnHQZe3m1w50/XBX
ERwEr/6FkoDV+hzaIYy4rZ8feIH0g9OnZLn3WtMdprZBZvmyg7ShE8oZAEurejsk
JO6kMbNu99VcE72enMfiv1u70igodKXjvW2LIGusId7vSGnvMl0v+TDR+drvWR7Z
dSujXYuxca8qHjcujAMNaXuunvWmuh6sYVxMaCxaGTAvZiukrx7g0vIUCJVjsxcV
3Q1JBYmDDfOe2C2yA/IhPfE+0p58JyZDTBdOL1q3e40DU6CLCITZ4VywrbRucdXw
aBd5KfiX0OFP3tHQmefmSdl8H+CFnO30HvgCW39YJF+0+wKE62azOhiBNdBPBXLa
yz5gW5qsi5VNR9mNSDsF7IOjICiZAYLQU5JVCU30ZLFXAVleCNNx4qZssxYP/C0i
mnbB6vgyPdN4i4uY2wzyRtpaSSChp2WIo8XVjFwg1tglcH+iWmIAJljR6g5WHSiS
X5F13ndHjK1t3J+0AvfmObAMQtgYHCdqwbN5XwUiVNtmoH1OWaI/YhEm/kajEcHi
wF4wivjRHXKYcEBWVRzJWj/JYqMl3usPLtSMg6mHex+/Pqe40gOvLCxl/bnni+aA
XawUqkrn2ROIu0YRTjR6pzJ8/wbJ0BvUKzmCTr+MLgXVzjB1u8r0AEdJ720f1ecz
6EMiJ5slW76SlU1iW4gLGhYyVJhKOP6wF+D4OZgvHTtL1l3eOpLB+iLkychuZcVw
hjK8nuoHX4ZSHUEiHZ1SSUpMA2gElRGgRWrwSLEaA5PwJPI4N6yZpuKhkuQjI3DP
3n2DI+iGeOgXRSHFab/j8aEuQxVBwW+W3Wycy8wuRmZFSR+PA1YDkGrY5lP5aWo3
6SHRLdTDd+8UsRncp/S+Yn8U9cAfeq5oW7MynOqtuBdhzcF79MK6JBaXXCj8ccBu
6ZtS4QBmfW38+Zzfk8XK9zt3wvsk9olQ3A8VzFZx4nYTKgywVzdy3t09GDqmsCd2
HyZhdnCCVtqpcSH/LUaUggxm6UNuZj4yflwQ9mx4AoYgmb7LrN73a/VUMslOy4o+
1xNDnnaQ7n9vjNYhKmt7+ZPmjKxNP/1ln7ZWljWB3ckBIvtDkuI0MHkFbUsLu1n/
xTa0f5xDS7rrOhhGaMsMrGnvi6WOFNKyDSO42yW9BWqA+r9KOMv4KVnSkt81RHrl
KQaG+H9M/u4ystDa57y0kt6fxMelg9EdDw1Vk8Sqv21DAE6U7r8zDxfBn4/6hrxp
Q9PbwB6q1ffp9bj0gcXFhd8frM+jA8KGpdEKs6/oa06dJLBj8qsGTV5sFMQyQBeQ
oad0TU0DekanWlPsTYLNLba82lHV7B0rHqJIJL2dbfaF+nc7bRhZL5K0zOn6HAS4
nMX9jexeqaF4KUXIZFwkUY5UbzmINkjeU2xqKD4oxbyieYo05HwxgOEBn6y4tK7T
UIkr3Dk2iBylRrlKhL29bYlU2XlDcH+79YN+cYPFxJoYTCq2/scVCHhIi4hyrCVl
xHhp0zbExbAQcLILQrfcX6j093fUJkejWrZsLR8hb9psUBJNV3pFHPSNJ1c0TBN/
tfqlRAViMLifQBNXKm3QSTcAizm9h/aSHezwCupyuDD60izg8qDsqeGxCu4uB0DF
WHQ9NDF0aOrGH+KMsBAxroRrTSESSRG8B5fTV12qZ0FhOQERG+h0GpsHhOtXsauK
wRRyRsBIEVbjAEIYDM111Mxs23h8srSKA654DXFpBIySxG/9OY7bSiACOeDMdACy
5FhuXiIZza+9zOHfKM06L2INc5P0FFNSMvvpzXdWwGWRxXqSM8GhThCAlz7ozM/r
NUPGPYIdNJwv3NYktM5wUxG/vW7rEcDrp9APIlxkPCPvnKx3bsUDYKq8T9pbu72Q
p5nccd2B9AsaGX7hOltlkg0vankgQEGDJR93zHlvavJSGQS5F21X4FkEHe7puoNq
cfzFvw4n7uFWwMrZOkUIbGIYGwzai6LhoSt481RFLMLzdcAFZH0H2xmH+9Mxj0gU
BsRjI/9bmclqOSJP+0kYTXKKCHNHH98hSZLuQ/OTDIu0t1Oh3gQ8om+eAKgXqJLX
hafs9ddA7saWaY+bC4OPB19kqFlceHyFlThOF4kTFsUkwjXtVOiXAvsFEmX2A6qh
EfFv5kcTsXxG0eAJ5ooBHKQ016JyuVVcgWA8JD4AdfiUk7pMA/N/yIDfH2A4j1W+
xHuLLfcFnatlLz/qMIk+3iXVA0Jc4vfiYwwX/SvIe9ygNAYT8zqtCWBQDRrCyp/y
WhZUZvDXulo1h0JT9e6hv+hWdymo0eD9+DIE+K2tUjUykoVvt+HFysH1bXApld0H
0BHvWDn9gbsgEh2E1wTzkcQJQBkxbJcyIc59YMLbieEXVflVfMI04ZTDA30IMIB9
HbN38ayw9oZCDfJYfZukB20vNB6bTLOp7WySkTCSaEcQxqMqP25EpLAYGZuyFvn9
XAxMWFKprqyReid2rYUV1h+mI1BNP+uPK/gNtSJbradJm5oqzRUB//q3Rg5Ifu94
YhO1EZfFg+2FKXActW5K4kGM+Xef3PQPPIUL4Vj798L/60VMWahayM2rtiIoWJLF
ck2cR5YS8hXDklvu6XdZ+hXqPEVfYWGmqPZiQWD5TSgfnjR2TnOz7eUEuPFAZ/Tv
2pIiSayifmm74qkCO/i4lVuLJVNXVCX/DOLs00h5xheoaGZgO2NazVnzJlab9SUF
8Ra0gYdau9NadpJcZBE0Y14S/Dz4XK5m8d1DVFCxz1bKUay/2ZDFA+DaqYf457mp
htEszbU9lsTWV67M553Dfh+bGrS/pCSozOaE8sRFqP6+UE4RgwtOW+Ku5RN8C7gJ
HTiz0+ULvp7VNqzRYPe6U8vI1gxo8DIybLoK1ca/r7TOogT0r3ScMlr+vdz0LEm3
Kxv0HUHK+bxFXR7UqJOYN6U2Fu5loaUqtLRVrLpoBTL0GDkheE25Ehuq87bS+Xzg
KienNsBmVMEmDM+i3UhuBmvnK5AMMuCQpiEOViwDMzoogieW1K671olYup3JQBmS
sbPUryrbXH0uSIg7++YPdwxEq4iQ3Cs+FGQmEOWDU3pL+iH4RZVD1boQHY1nAInS
YJXav/2HVRSeh8nsYgPRtmiXcUpdUsO2tCB1N49rd8/eG1Y2jlQ1AarAizBs7gjB
p1dWNiXHh7qE0Ks5Ox9iW5SCADGpFd+icQ1JH3lxW72FEZBhEyU6iar41kXIDai0
lIgsklkZPiaNI1klS6YjrNGFJq93kTskjlPScKi3xnyXl39eBhEAPhKtIximhnfw
dcLLKaq5NV1dzdnMRlRw5DgBEm+T1om+nug8UrgDfTWpNzIrDS813DMKsnrzTc1m
cWMWDmpsEbBmHFV6oZZQK+WIqE6jxiIUxxNTC8eKE0TN7IAVLkNx0xjKtarlm7xv
PqlCalQC02yh9QP698SfOChy1LKPDLzuprffLHeZxD6rJjFKgkhkzPPyEwUckxps
V90lQ95YRdTKSCKNhE7CbbnRVpXRApcLwLAIRJeGEluZVGMonGQLUQJtNnTGnDpF
g5pMkHwENj0BDBNEaFMOTFiDsYrUs0uiMv27sftXDT3BcRpAaUElEsETc8P8TM70
vAfhiN5aT+n8cWxmZTdsjctRe0ojjb4W8bMrqLGiGlfIcZETqdVpu13SmDNhg/Vi
h4b2dHIg/z23mGYDgLpsVy1IAS1r8qqlPDRb6+zGeY8ylarvZgbZSRPYbrSq15U7
5dz8HSKKq4qO23QDBDVgljPBum0eFv89gm6olJmEnmbMoWvP+n3/8NqP24f5CLXf
T288lga85F1Kagi50OwjTaCjeNRtUiOMUS5sxoE+98csrGMgjujz4GDSJ7GgT9/f
uisgHpdWyAoc0Q2TNf6R6IWZxPIU5Wte6F7bN+Lnrg3MgJsgP2WU/HUO+phTo6Mp
oNm44Vm6YI8y+fIYyQjioWCus5WAWYygyke9Gnn8EBW17E0ItIl6TG8YoRpCMptt
yfVqPE7uRYpzY1EVJqqrf9SzZ7DkXEGoBCUKW+8eEryi/vX6xTRomr/QPh8cUfS2
m4SSTol2wq5yOOF1qYTBlYzpi3EWg/F6kA3sj2VXXDJGIJXC/cDH8hjzzGjs03zy
8ab7i9hXHQqyypteGyMMZQHC/buFWpUZQhqBNaBRav3K/Ui7jfQy2JisbM3ceAec
IB3e31l6i+c4zlKM4ZGFo5gMXFE2773o9hpTmIfG6h2YHfCC+YJw6qk2CKgM0UQN
+jW+O3e+zlE1/MXdwxLw46jhlRR0Jqmbd5G04HdS8v+mM+kqcebBCYF93xL8LECj
UAqmBMoZidYzOAzcZnMjN96XH4JMjMD3DSSVw0JOOKnD01GZT89gtOos1LnKHKSU
5na3dsbfCyRpyDeAegxcqU0XKWyFcZeISQOQ4l0f3vRHDH0hfZ1Z6SucErBEawb+
e1YZ+KlXq0Af49zMi6H7hS35QLYNS04N6XMbUQVioUpefpOLiON2jvw0BDnxfJ7T
aRWqRWfwBXuW9qp1ib9wV3XU9d5jZ6v8ioe1lAYZt57cWJtEkpm4N4fKVZrStMhg
4KVTfNDY5uXXDRhFi+5QLLZV/djd3M/xamx/GFUCfQ6H5Y4ACN8nS32iqB/HamtG
EOl4GY+HN0CabU04FoyKnttn+7OczlHzLX5nAvzG8aWYjJWM9oAbFC1NHbO9DpoG
NSQoj05UcOpmL7Rb6FH4xs1Qq0/stLavbBlO29q/LE1Bo8WFXOrrOGeOh3LNKSFr
km9q+wEEtLAxrm5mkeIqPiDwChHrEpVhv9ql6ltM75cHk2GANYui3IA5r8zWwlUY
acRg8aHIc/9MXL+DrED4Pv7Wa14SgdZWRU6MAFUYaSco4BOZlhCpBhJCsgo+aQdk
DcjdMcUHEbG1gQ0Um+WCiGUzFBbKpQxvesLcvp9Ki6HfPdPE1FznBVTxQxF55Ttp
9tIO9imcuAUAhS2FOqjyL074TBcHFZy+pHZx51l8xAxva0zwdj6Qp8/4UGsVsxOw
2q6V85wMjPPfL/KvaOX1Io/ctEqUHdvxNweUSzuWECl9knb6tngMTMfezcSFKoKQ
sVodJIMvtWauCj0Tzzay01E25X+Kbh4D/J2tn/Aaq5rVFdTcAPDyVs5luCmrk+yR
E+mpvIl90FLKkVUA8WruFVgkoSWI9bkLylzSe4d7EN91HZipg4/DKrgAOPsoo9OK
HfJRpjL1j2jIAhhnbt+ch+Yn5kuikA+qqVMDOfhNCFMVXFVfMtuS/G/68kC65wp5
UgqyA2+R3pRt/BlAykuZwbp9CUAmmbTfD7H82oMutOIE8BVqtCEz/f3RCpMSnA0b
4rgM+F9EedW1aHlORO4H7vs6YjCoBMNwFrXfynVPU77zCAJEbGdC89h2mf7zUAMf
Idce7vbO2gChTKFXr1D+nyXrQkR1Jk3mHlVbT6Q0BtkHyYkAlrGxGB3aiJ6xFU13
j/tz9zGB4t8Y/F/ejZdJaB+yxAHkDD7buBL7hDdd5XasO7Z81CQzvvuGWzg0EHW6
yTEeQ0t+XMr4OlcIJY+Nbbx+pWAmo6hHXwAIVqPpQsbW3EWrlmZeD+x1BkgDsvjS
8WsoZlY4hVtzyqcITo3zk7IOeb5mfGzMX4rCxqxP+h1RZdrQ3RzGYVggnMBBDnBT
btrJvftt68rHckEwPRC6Ymf7SfFv9/4ghlKpVVTqoLTdvz3a84EQVXE3aSdcy+Zc
nw/ESL8VRzCHQQD2ShWb78X2JL6TOIb9eMyU/nhh0tuFkIPItgvWtg/JbjQTLaVd
ztATcPazgCLFDeZBgDtnYyBw/DMFX2JMe+L1WFMTvi4pEMD+nuyH1L3T48AA1CzI
tLPDiyoSkQEzHGkV7NcrRLM0nBSWelEU9f9HULSzbI/inzAfQGhCQ4OwDhco90X2
EMG4A7a6ZZpxxZVaiV++zNCqqmWu++YY8gb4vrYrQTPWf5yovd/gJWoJLAMOD0/p
s6+GsKxUP0msu1qRmI/03/mgxMg8lNN/qOkgD9FYQCdK974dVgiXdKzLhKSu7OE9
Gw67CCILplL8qNGpBzoA/lT96PqyMuXMATqj4A1bhurysQdymk+Cd1QO94hZKSRV
93Ahwuussi5MSh17+jKOCWXzD4fgcfyiIPL829/Q7KEawZh4RIHTsGNaigZ/PwlQ
8QjG0XV7Ts14MyJcgYvL2b9y3cnCZnb9hp4yRsH2gAJQtAxaJeQbv6iN8AFsoD4F
R3mS3p5suNxXthwYULX5kDo5ee8W2JrseHWXI72JOaGhUSYHtyFZ+s3IlAj4209c
AHoGcxv4F3ks0jeRX9AUhZGwTCadO/u28zuRzaj8pQUN2KGdiekuitJoqAS3Ljmf
Tkl87e1Aj6dZ6iEmdNr9oot8sfVI4DoPy5NmmDiz0CVu5wyjcskQ43p5sCknDrmT
rM05qEhcTw+3GNqHLMhpnGaPN3v932dxDCJ+V8zB6NCFuGMoC5soHys6vRGS707W
rqUMeCdjJT/SJlxbkT7Fw1kn++l+G3atR7HYT0W0p/cxSuxaL5tRM+ydZkilORH5
xFKb36+TAYEyQVIYZnVNmJGFjsfOAskRBWlv+pteuZ/TBF4HLrNk5NFD9aSEzQfh
EvJ4dMh0hYGItLlmZ0grDZmkfHIp5vTPqR4Y05FyYyJVFkElMUgeo7QRPZzoEZm4
PpJeNUrJouIo6nfcKX/PvdfAEK3RyJu/7LrWlPna+nCvuo9hWAdSTHr+uQOUfcpS
c4m9s4jhBtf/rNHWnOVxZvT2js+FgZ5n8S9EMaOL6QcZD5pQdiCfNmee7Ot6TqNO
YBF7GLn6SgCu1fAFkffLAyzZ7jiS7sogxd7biHFf3vx4twHBTM5TcUGvCKIa3gGE
68lsX5syNiFsbXbbbGfAj5Yc7FHCcbmZDHN3nIOkZaxIwWQXgu4rO4MjgPkCYAeJ
iAqRx9FIVLr/KMjpKSZkOK4WXxVwBrfk4Qa+YA8Pjb49f+MZIPa8z4llVxM9gYA8
rI2rzd5ku/xBmOjSdJpPqM6mudRiAD0s+Ge7kgYPyojzegkl0o4eP3JOWZjD0iJa
jep+0na1JwifE6ObnxiJ6rtXzj8MRNqoZ3aJMTglvsMN5Ih4q/ANbBYNN2qsNPHS
8fiKXFVPubnPZfURHfVEDSSJfSzE6qiXE4USOn4UKLRILNx5oPFHtNdUEyUMSFXt
3TN45IRo+UiqvQV1WVM2BEymqXZwu06XmsqTGE8s4ABKf+X1Jwj7Xf4qxXW1Pgoe
S0YSTDVCtuFRTVxwu1w6wKsZAYVH+8r3tugq66IUDCVf56fQjkM7nZ3pWkmtYzYm
fCQTBCYhUF4SGejnpgE0GDtU6zqnpvy0YzudcA90T3VpZS+dyeoS+YMf8DinQW6G
OFsNQQxcRLdTwhZX9oyr+lzwPHGzL1dlW57WCWGSFheyiTjaSebxMw3h/RPsSmHp
m9rzePUBQkbADY/Pl0W3uD85pFuDiihvju5m+SRhOXIEnt3LhC3OxWJWS/5kP7KV
PS3UX2wm0M7LUgTJz0YVWGQC0C3/FL5mi3YKRgTlcZ/2bwxXEvEGMO2gi8hz/NF7
NdHLvAHbHwSrvvX8KAaLjMaz0WyoUyDBU0DI9pl84EVDcH5oExoJg0QXTrAJwH7d
lqUdt9Ccvnxdgr2N3uFOe0931nl+6BDInWhoS1Qpq2BX4VIbqNYm4uQfNCbjrxEq
g2HJX/58ynyQy+O8hD5n26Y0RdGs9Pru4rHW1zky0n68wILlI+EAr9YHexkhyopX
Tqr6WQSF/EJpurLLTJtDxrrhk+nMbEPPS2SWIrWxW4Wsz5IAd0ExMFYYVbdy/QEj
0Sdei28WYPLeowf2ctDR0u5kqXweuX1i0CaeWT815kiJuMvG5N2AlQ8JLbuxZrYJ
gwUORrUZ833LX2GXifosJxwE8FxCbemfAC0Us8j+Buvrp15bVTmWZOjBzoSw23WS
i5hBvfx6Jhd7Bm1F+1GcR/whwiRRuHHcmwGd9MZCSZeFd3t7b8XmoKMLYfgUe+UW
USYNOIXHpBcLiXNUh/ck09mM7J4KDRHzf/ZMuytG9uzHAxY3y5VXZb/FDszIBbgy
SsUZtKQWZY0ijlBLBLLoZeYrPcK+mDE5V7reYy+FGzAxVXLxcF8zqgi/WKXrIZHi
CWkJWcmUlSEuOZNQIVQDZCMGI1ZYNfNWTxGqOd7LLI4pdjuVXrCLd5br7F7T/ePz
qL8T+nERUMTIyimbbb8QF/QhSLULXxVUGB6XHX9rKhiRykaUUEuWXWHJw8xdZ9Z0
w5Uy7Kj+PALdQiCnrhHXUL+DyjFJb4gR0M6ucERmHGEwQs7PhI+Td+s91l3ukQtZ
uxVFqkWSWX3nDEkIdAosvGcAcNuVoVTgnhNAMu5QV8KekbU+ghZYruDoLyFHc/NM
sK8t8w5+hTNDBjIyrveEvLBg3YtPUocDwmKD0RJ7ZkksBI3aCkH3Bu0oYdRdFZbl
3iEuLUGou99rLJIf6Z82B+MLK5k4t0HCW7qevNOHQ86f3J6OEFAlz+H3T6oaFgbk
23zcHIRRIQ0AwwUWXwc+s69jwIeLXnwE3SSIRVl22Vu+bFi0RAe1SLR6NsaXgDI5
kgs4mkU0/AIav0LAm1Yj/R3CaBFo+Xp1nESyICts93PDWvKtw7/f3pzkSSgMB7kB
RvmP3DOMqF13JJtbh1kmfWnRa/iisKI/yDtxGXdKCMkaRYmoto/2pzkeLNSIzofq
ZNJHcqmggc1fRzP3OQ+vW76fIExrKu9t9BL6zSzR+TGh52+kR7Kh4QVqWkNkgysV
MTUEKoEar6yPjh9cGWo90BxkdGELDtrcs3veoFh1q95p/jriPo7LLjgdGlZNOe5c
6L97sUCtodllDqtln+BgeSPh430hOzmxDFvRclXvb2snaERkAnS4VyMQpY5Bzpy9
3A4JKELUUdenbDWOAptoC9cQj3BGF+ts6GutmdIL8zQOQUWSWj2HVvkKcvo65P76
n3toBTLcGBV39sgrC8g5UDDPTVIgT6MdjqCCqpPgQneaVdM12X/ZTUjCGTCJDB/9
gfiAZqMMzthb//rir5lGmrD+DWQw0HW7dstQ36mLtJFYadSWm7PqyPn92KCcEiyA
JvnTK5CXYH3uNudT4qaPFwknpvHZPQRAseAED06m/ZjTxoYO65tZ7/Ks/CaM2QEJ
AKBrzlHJhroYI6JVEGF2U2eS5A2gbHlCP1YZm/VSEF6qIpoPVQhGf3PiLTh1e2eB
aJpo50Sg4y4qNEypKBlZ8sMQMBTfKwr0NaOS4TB7jwDOHmFb/thrfxqtAnrUuFx6
oFIYV3EGS7XR+9D1lCTaotmnW3i9THqoovlk2cL6h93OUI8mBXxXsQMFOMKlvQ4c
aK0CJ3r7IVpMCE2UG+Dvhub3XdhK1DcdVfY6F/xTBgaBE2Y0WZ34NEckCiPwLXCB
stJzTlxESiPtkeN/00+MT4pIpibGBq1v9R7O+e3HIKAd8EaLR3CKYXq6oVIaUVHg
8Ej9JU6GasrEt2p7Yv8LZtHjQqBPZvJU68fa/UOCTFITYA+z5PMtyOcoGkmfhBM0
PSSCRAqXewej2zNV4H2I/H9ycpwEtZO4ZssKcqIMK+IRfjLKmfCRL11sGnNVRX5I
8yBqDLwKyNNysTseEWQnuKsrEDAUebgVISDdiR9PMgn6nf7oJDZjFI5VUFkp47PP
vzocx5cfORY+td0v/jIqcomrMYVMmruyVeeB1C0/hvB+vtfVO1H7oqgYBQLO9y6q
QX4qDkN8MKgqrifmEyQ1jhXFO5FvYcMfBJfzIGJrk0O2Y7eRpMnULR3yqvodpIDs
+5P3cqkiPzNarWyoEkoX1o21b7qU/mINBNPhHd6fF+TK3HgiN+tkTAjvf8Nq1Gcw
pN6PEWsFU/e+NLO3cKVJE9DZG1SLaw7Mn9LZBWTcyJgG78B638z9GHK048YQjnuK
adRHbDDIU9lUCVM/7ch0OpBsykN+gVlLm34aprxyMzlsoJVlq+btnlcAf5ftrCda
+NekbOPX7DuB4KJD3bpyknzYn8r265/xjJBV9ro+GbLGxrrY/PVbptpfZsJ0VNCv
FY7Sp0+CPZW9obT0hKfJIOuIQCC/qRc4bjQFKtRK0iTf2oV9pgA/GoHrLwze3x8U
YrPh5KodsDHUVq8e8NTT8oCbNrKFbqdmE0qThX5FGQrmFru8Ea1l14K+qEt8WJ6S
o2p2ewpnfDDlX8wIJEPvO2NGzZRuQPMsmfy/tOcnmqys4GffkDqffGbEmSuIpioJ
EkAMrd5bDgVQ7ty9cww9aheihKZNWTtfgVEmL87sVi3eYZgOvN8BaYMD+c/LqLZj
qahtClQHQ47DgVzdBSNtelnvI93tjBchPDDyO0WtjsPSdoHgP5X2at+PVmkmuPRT
Q39Ik4/slWo2D8jvDl4y3G2MjVRP54L/Nu8AKa4doddv0q9e4piPiZsUeUnAMn2M
txckTBGGKPpXyTeZjyR1/Wi95RTikw2ecRtM38Di50FG33i7V4FTF/1R8Z1BY75O
QdZke35KMbQEafakkjjtYGe5hCAowZ8DZJuYrykrbgPEe1YaWQITYTdmFVsAm2RJ
aciKnbeOjO5YxzkT1eofxY7Y99PPCsihsCyOVivZ0+Jpvwo3n9iDsP5CbSLB8E6G
WEvplY8XrJ2kZVyV7+fbYpgMxg1UVvdpwoyLYUJZ3q/4pMqn6DYSALt7KqCrgav5
kkh8bmMzknkFbfOhuSaiw7smFyE1bQ4Qq0CL3y3r2QGpNA8fR7iYxWMdKsO/H63y
79qlw19uramHYYQumYKURc7eexb0iOjP47gIYjrcqGlzoco2sZfEB03mWn6iu6rw
ZdlfH6NgdbxLQECOJX6REoSG8wG48o5wa1sqE5WJlI/deTwzSCUXYIkG2JCBMYPk
bwbYy6p7L9BvV2qvVjysmkMfXkwHRmVQZvtYV9eQZJL4llmalTCdWKOKTEav5BdS
diVo6C8ykO+bNpXkJi38K8NPYzY7RGf9pekSLaGIQ7pR7jbbxfdq4WEXA4jtNK+x
ZtiCCLBIMGdRLQE/50+OjAjoVLnlS1O1NzOOODzLlCOkb7N+96dy9a6C4RPFdH0r
mlTZ5FM/BnVz0QVNhLD3qPmzTTu4aug/0QEZm59EHqt0iNs5RLLkis4Mslz20AoB
glx++Kh3f12ZaGMvFuABBc7ml0jyHP4EkFdPmC6yFWmCOFmdQMfL6G74c7TYo9bf
LHeH8CqGHmL/10RtApFCzOH8h8XSxr6qy/8RvFyAVOiYK60W9kL1/WbMcP2M2iF3
2ZSvlMw2d6m2etIsTp1Gk9aQA0GLhI3oekC0jv44HhbEiBXx6x5K7eA8wRtXAg38
LwWs+lIuoAS713fcWDl01UIl2vjJl72wWDnRay2sLpZv3WE3Zby5LQ+DpbQMBz7x
DrmdHreynrqhQ2itDn2UfhmQ0sX6D6vM6UYKHLxY3b7CDncL7k4IV2Az5V+75I53
Gk63BFASmWYniV/FhcYOrTvnelSlMnt/k3x13KFPnp3HD05ia8Itgp5i9JmteN3j
uWcIDCz60hUPuRArPuT8dupIzu6w4EoFHUyi11JApkKVrOm1OlR22pTWToa54ZyY
uUfDXDhjgLW75KTgT2YGnRz7+YTqk3CMvbhXKmxOllxspLexcvNnWyov5t5syQNJ
HftnWO+sF/Lkq1BvE+H/s/qIxedu9YaBzXiYiP/w+XxmT6u4exDJ5ytEi2KySIqG
ERPX15vyW5O9IWFZzchpvMJ9uzbMgfu+CXYc0wmpvgn5IQPvBWCjbZkr27+O1um1
mcIfvGzJNebrwd7i1F0tJqrMAg3Rsps27qO6WOQVaNmw/vP6WEpMGXXQr4ibdW2s
tNJS3bwnrncLh5KthJ0XOrw5pgiF0PO1i0vbkHgnwia5RNn1YpDXq2IqJgQaunU+
IKhpzWNETtul7iDr4yTzvPYz9OUxMYNKF0vcztLJAUusdmFP2qWnKricBItE43On
VbT/b0SiRKLHJ0AJkV2zvOYr2vHrbVlx4JD0vonYCXiO/KOfNhL/Zla1ixe6A4XD
VKzKrSXMQPQZmXRDvqRCZeahkcX5IU2PJV66kH34lv5eEvRthzcdwQR76s6vHw5J
Z28MwzLJgs6mKz8Acj6CigPegNeoxy24ECMsJ1/A3Fe1dOFm+XEZwofZoKEXzMgh
nc5qFot8PsrLnqjCBV43MMmBmVh6HzLZN2zH1d1FGTDuwKCx4pleoQFsjf9QLrLe
TtPp3pKbxjjNp4Iyu539SsFZdaNHTxZyLKtoclZo4EFW1HW3LpZdppAgBZ96s/oY
Zw574LNHmzrqtGtvudiHtNlC8FffWaNEE+HReYF+aP1u7KozxHa4N/LpFUkoyrAY
809oFjEL6YbsO/w+cstQkJsAEbnQ8j/tf5k4BWhQAqKP1BDrr1JA14NfPY61c7EE
xW3cTiGyXqBvj0rK8dqFDmnUNAvSn3YghdSLq1kXAlkhLLAOOwq5WfVDV/PGaHrQ
8a4LRJhnLHrQdtwsY5VRppnadmzvHvpNk06sOLfwu4doX9yN/d5Kxk+GVAUbnZyJ
41/wQXRvr61ORKCayExa3OOGn5zntpyXKGXzgqwIjZgZHR1FE5ufGIBFg926SZ+t
GmvSVeDVk4YvItCcR5iJsuAlMheIq3TS7Wwmm4ywaS1phtnivLMn0Asx+/sdqFaS
AbgizaZOTuBsGk0UCJgOJYC+770ON1FIymUNkVlfhp1Uf5fSIBY6Vz3z4MQlnX3+
mjIW5VnA4t3I2nx/hEF1C09jKeYa2Ydzr2JZUiPb3NMZioiVbO1WYAMArtrszSt8
LhyHePyuWIrKqgDVo9R1lerXK+mo2XGAoqQcPvbLGByj+PV91/SKHM35El0ZsSMY
IuBbEaaDxS38f5TW8eysld7QYJY53gHiBlhxcctNk40BZoKwA0eqpa0t3Ofj74bi
zP11zJCLzOHXc3KHPufNcRSichGyNKMpa3bCv2McC274vSo1ZsYFiCw5yGYs4BLP
fcNBBrsll++EB66S8HggkNe71I5MS0t6OwM9rh+vuGg+hEg1LmfOD6fW+kW6i+Hw
VS+4iU4aP9NdMYIh4v9wjkaEOTsgQzzofvcVj5mUo1RaFF8oFo9e4wZMTzKrvRpw
wfkg6AoGcY7q01pqlFK2MGUopcfxyMJ44xiahiksZKNafIYH2qUdp7ZTNF25zw7g
q+cx1ECRPeV9ZUWUWkKUKUlj5c+MXHhL8r3QC9HMUtVa48/turwTJybTdki/2d6o
CHgAkvxmo+PLM6koQeOiOMXDJuBCrphjXcrYA3GgKIK8UlN3VCGzUcS7zEjJdFID
kLHvAu1auRY0O19AXvcky4iLI2041wuUUdLeasESrA6VFe3VvhDhVl5S+gjDnvK7
KkezvdlPT+3MZDdMYnJh458gagiMu8vhvzaixeVMO7Ii4kGVMtcV9OBb5mIGrAqG
wNabmclVqL5kuA1+N2lOWgSQYg7BCvXALkPdvrczTJusqoNG6wlKXl89NjfyUXnp
ePrq4iqtzfL0RLhC6nu24I3qq96JfXaVAJgXV5kvX3kKpx2NixEcZarxY+coNj0c
mjX7So1iNKDdD4X1SK5FVoe9vjVw7gvW9TMh1pnY8VFFZsy+SMbJSSziFfLnP9nS
T+dKMcwV9ZXQXxZDKRdpj24lErldXwJDn1AOR9KXRN86JalDz29heOJauXXhW14v
3eflSG0g2en+nNqIzhHoDzhrZAIoemEh4Ihm+/fM9ki0ohnOohe0TAo6fdRz/ENL
V9jvsmiXAz6xXJ9POUvrVnGQs6BWPEByB0cpm+KCs2oMCBGoefGMOrOliMIv0FyF
cxgoLxZMgmzcAGi88f2LJFELGdKUynebCoyybw0h0QEhXF0hFztXzFYxWiL7nvry
8c6trVta29snbSSFdcFcQaDPi+ko0PztV5+xCnH0BstjUVGp3saJR0KiyWtk/5/W
bXHj4hIh/G39yF1dCd3lP+S5euwwcdw64BVAiA8RRGbJyz0edJbH9igYE7UMmCpK
e5r+BNpyHUji+bCN2xsuFlHiQA0exCRFiFgjh/bMOoCEFODrboRv9qkDoggcCoue
+bhae1oMzU3nWP+392D75aWrgKx08bkvHEFbsaPCvBygREJDKKrbmuvcNed1u7TG
xsDyi0A3zTJzCCYowdX/+iH7AXKcq5IfPvwCZ6iLvGJmx5ygOf/TNYh7GYjjTl2c
gZFSLZhOygs4fU9iDoAa11jsld2RUFZsB6GDPCXVl7xMJDYqcyxZ0rYbR4jfZG6N
QhRAX7E5LkspnA1Bq6OQHm/WD0qzHimQLHT3Mfg+XXQ/WxwtFl9n1oeseRUK4vnD
BPekGkQkoaAsTqKpRcbLSK9mYa7jwbROW5n1moR3w/n7seb1Qdq2YhLR521N2RBq
Rzp2q16CGgCIOn2+ugwBzRqwFUX1HT0hbzPmfeeqadVrvWzflIbtAEPg/4PvXA4i
fc+DCjvmlQZppd7+lU4XQbJ/wZxtO971bmp97feO3nAMpmDtH+CLkwhwR1Wn/YfK
YIF9fyTrSM3+0n7VFX5xgUAGNIrySCuUzFsfTeVHvp4P4coB7FnGFEGvsmI6/dO5
mGvbHfmG+vjuzqvBg2Ifn2ZrejcRzaUS3ILokvGXpQV7cdjg+l2RrfM6+XMH36TV
/WccI/4sFon/wMtZFh7Eay6X1jXOXbZg8V+TLwVzUKhdRebUDtKz/w+ZwIom4Dr2
zN9g5aup6dMxB3XhPOKNQpd/tcayXWasuY0hkjotsE9whFn0EFfewotnu6YaKDY2
ak3CCPsDivRwq4Xcy7GyuZQz+SSYNGzArvvTF2yZ8HSLzlJRZg6tQb6RUwXx7uAx
v1onmX9Uhurh47AiLiqJb/AGCxiq3BLky0gK90gaATCrxkTXg4TLNsHvR1MvpohK
7dLf+4PD3J0Ue1zNA3KJtUaUXKJqgqVJMhkMCVvY3Gp+XAsaVE+n4PnNVFwmCuNt
UOkZo3TrDJkuJvhnRs62qVIndn0h9puVUQARlpbKEUEt0d9mBvJYsRlLJjxsBAvb
QHsoVdqI+5xcMdyn27sLGnRvXZx80ZH8ETJI7TJOJ51RKr7KDPTwXOfxdjAZBJx1
WzK+IICeGmzbAFhBJ2HguVCBRAg5vCHnZFSh92yfOUz11LYdmTCVfTAZXp0/nIQH
77ZdIodVsxU6EkuFmAna0PrlUT2mIE+mET6ASqmC211pkQh74W1bEAYbqRYvS2ir
CGpJ5pW6j5FoO5lBCWU+gi+gal+AomafDkpLK8QCxW0NsXQd7096aCf/MiqaaqNh
0fjxZi5erQrmIL4t4uDn/AGxrXg6b83McUtmOmSSZlempCGNYJ9zyqxR7KndgL4b
yV/WVu+lpHI57Lt+z6uQKb0Lt6P0lUPFCebiKKKG/OID84PCYJB0g+KRhW2aIzxI
Sqh4WzN+uir16F6t+PfF45xQUqcXzZ4xOXJqtjieeU8R2OjSzptMQCXVqeMw0FK4
244kgxWdvl4PfWyPrG3OaXmJmCbaqWCLdatBCGnexQkxMESjKy+WQz6QU8bqTmfh
d7bb+iJ4S7QVhVjSaf8tKBHvDW6DcUwCPA2ADu9eD/iNrvVPuW6B45TaJfO4A9nt
Q0TKHkUI8Mj68xsjhs4GvAMBAFc1R59EUk7ydA3kOURjqSI0OZOrGB5ytrX53rz+
hoRJDxjeSMQlVEJlD1AdSkBEMX87dF9J0wPAE/kxOHx+4BYtn4wfSFf5dMrOkVhi
uFFIMrUKqm9vsJ0IpweZNSJEd0vdalyRWPgs54qHXmKI8oGoEuMoNUKmFNr7v7O+
Lbpw77otrXiWc7Le5EkSiBzstcGIr3luC8DqvgizENEIVDkDXlhasDrzPcxOflCx
BcKmcGn7l6/iY7kJhWV6JiYVzzoRquyfQ8HVAOUbB66ge+n7s4z6PAFrUMdx6OSI
wTYlIEe6Abkmd1bHfNcsB3RfephersH6EX5RbrD7FT6n+McH7yWvPeUPxSaSSX8R
exv15NbiDCsPeXpw5vv4hdBOYlhbInuM85dJhmx4EWi0z2y+MY9kIq6NvTneko9J
wKqyG5oFeL6HrnjTESwovguhmAIuV/qtAXSvNLVkyB357aUE1mVOYHSCeqHOhGcH
SO+1kj2Cwv9VRw6ASLWPFuZZYFcYUHOMVgxJst6+niY3RPEqW7e72hiYkZQcsZwn
yE1vqN56+OWQVx3zc6mvgiDNeVfDU8sf2pnctq62TxE3QqWMTE/QWqKlRwpk+pgn
SxDTVU7NtrctE7r1TveGFk1XhmmIsGc5oTgi04p6z4q8BtRzBendl6nT0DhxJ2ky
9Jd2Co50rA/JMqy8BZ+gH3Ith6/WsZuPq/shPm1ra0qNr5X+n+vwwCr2//4EEYet
a1WyQ7scNCgDblNzdVWGaINPG47aTo3HEl8m8s2HH0RGM+xO9/5FZgHhLo7SZD0f
EGtxA+JANSKoe5s3gSgdQm2Co8xDelLhX+8Rx2W2P0RCJqlwdWLH9HJl9RlQjLfV
PFrNbKRonMIc2KzHaoPblnYaWrOYYX+StnG4Vyq5OkL47vLN+oiqRv2URO2OILRn
6hhc1OaGZT2/qLVG61qQe3X5ezeF8QIbHWmJjXCJ8NXzbxW35/hfdvo+kYoq6lr8
ZUJjI2K8yR9EuDsqImdepQFd14IwvWi2oOK/OeWABWmTdOT09u1HNSKou7wq3jsG
EoHt4X0mjsxdOsl+9Ha3L3swmfflDrnmG3PDjwhN5Oor0HN+a98qy7cIv1ghRtQP
CW/gedrgd1YLvHFrNkKlHmFFnaOnNzZtg2ln2yojVZfi9dYIaamPhSvV3kv3xStQ
QZA80A8JkkjVh50VQN9WYvj7079FpKSJYOf+eIB0IB2yD9uvojaZWazTEnBTZ2Jo
Dh13lS2PNCNyrmBo0P/DyuhdmPG07YO1oUY79EOnqG2LtRlscYoFAx/R1m3m8zBo
cIJ90R1ydIHOJAFxUaHxkzN4xkE5gemLz/hk7p0R0a3LkL1y9gSbr4p7EYRRQIgE
hOsOkY0kDCarsWmQx4KaWcm+Kszs3Vf3Q4gqQ11ckYoZ6GuqqZ7NUiA1kuwk3Cyv
q0vC+yYs3eH29zo6O6IBJwCLLSpMUttgRbfnqGyrvIEb6aE490v6Cd3R22P7RztU
QHih2KJ7RV1JPrv7xPkekLblIBjjCBOO5m4Dl6itOGrt1PCQj7Ov0rHt8ImUCXwB
UICMhpbZzR0w4WnGwsWSMMKxsXoqzZ7T+BY9XjVpAYQaoS3j5IN31RR+bZTpKTOT
Lo8yNICIQejK4GsOm6lWjLPZUYY0Ua/oiUt93Gh9YYPUvmtcuh1i0i5ipiwfBSlX
QU/l9Qqlt3tSg1Tep7gAQTdeZ4nyvFXw6CJn1L0Q6krV0J98YjssD/9yEHVQz49z
hLqpb2TqTrKk59pbR5CIxzAg60lLZsliQMhVLdjNsYfnBNsiqoRcmBlS7LgCjRzW
oSkgw6NHhoWsHKr72qj3KiwUd2YNgmBIXWIZVGwb3GQYragfcsct71bACKAK3PRU
vV4j/jvk1p5OiNiP7sbKSOX8xp8thc80MqnCG3HwvqaQP9MWFFNRPul0c+zkA/co
2A7O0NZxM+3RmA0MKvGQyqyi0u2skU3UN4Esmwzdnf2zs8jsB4i26UHvGyiSZj3f
SGii9TN5/KchHTDbU697x8DC+F+/lHTdtJiPtswgxgyCY8VyUhJoeCWP4f1NtSA2
sKRgWazM519QhJgOs98cE1bKQNrOlGRchcW89EAM7m2bTC6eLeL8l5z1yUqHsbl6
oWRERk4CRuzySo4wtJjRJO+mukxzO8Rhp+iroEHyW8nu2EolhHmOn5PSrF+9V/cS
Al7MHEDFBTRwqcFwHx/gLm3kCcpl6utEyXYYP0PVsN6pmivh+H0TqwlU2KuPNtbB
0WHDnp81MiV1xSpJcLKchWYtfpE4d7NL18CqNVMBXZKoODGU9GM+ZeZo3AtQbQ+x
oGrburJHKiTVadcyJ7qcGn0vrtEnq24e/QKBLzymJRJCtBm8VTy+XuYwSELLuuxk
WoofpksU1iaSSYCSHDuqXAsTAokLFX+tzSn4jErj6/2vbWiH+6JQLgLn0vpD9kR6
ksv3EhyIAFRvUNduKig+AH4eTVjkWnwObfSRFRpbQuLUZxKEtgoeyb6xE3qSYnwn
5h+Oc3YjX3Gm0C6v0x3kqykVwBLAOgCNUv6tbn3GhIsRTGRiMJV06UplNR7QyTxC
wMkKLK1x12OWHWBXbUKsofqljCrOjm6vBn2Obzx8iAogtM9lOEWHWrEZuIV0XDJ7
FvWwXs9gU6ZEw5NwCsk6V2yZyFUlYKiD+e+i69Eph4A1oOhmMNfri1bngdEcoiNw
NBQLEVqLK6SAQ1ajX7e3VrUuiRCP44QhY/gcTFxwQidzpXP9G4/ddgEye9m3lsRN
EETtNlImglOCXstRoobUbcHQbXoCqFgjTyI/hSdsKCEalnmyKr2Z02s7Z840wv5I
zwUaHmj8Q76P0iwWum5W3IhOXQoRCa+N8jgVVlm+FWt/+5jGM7Nl3/gd+5qYLgrj
kydX7j+8S8/8yryV8sgFqXZ8bAyN82Yz21UQnjsDO2MO2SCzGLTCH+YZk5c8Ps/A
zmULTvfnt+z4e1BE5Z79BJqnl1wxYta715N1vGqAujr9SGi1JOvtDMGLucpuU6wZ
iwgU5ccAquEDsHOShQF/hIuVwMQngTRKEgEWusj9d+QrybNRrNZCc9uF0TEBsbwl
y0uWDXWH/S9im+g3nSRXhA0/UdNDKZY52NwJb8ANTFBhn8BF/w8zzreQrafu6gds
ipI/WIgDnN2IuEVc1sdicR6ZCSav9+bLmoNBf6W7a7it0kQO+ydLCvMuSenqfdaf
GdFcXziCmoOSzVCqZ+YMHY6nV7ypAj6X+TkiF5B4Z1I7tb2k/1P1kULUGGcoS9aX
cGw2SBTJ3dY5VPuM+XsTQHmDJt+JDAQXJeWt0VbnWybTYWu8KZR1opfGZlfx2QBb
+IQElADfFWKX9HDmp620Cf01qXyZ/9vOb79K1UvC23L3x6DNvboFbIZBNAKGD2BM
dCbVNBYGh22QXAE5p/5VFq3gqoiW4JI/IYmElZdoTPprcLn6DEAEIi2MHp9frwAg
1c289OBNipXpT9EfJhNrxK9/l0HDAxx2cXISKmAwWquDm9xZzfcnnt39J/paoLrN
EiwKFm6BwfjtQDwTNXiAZuw3u4zxeMRcuYbadKbLn6eMSzmNIEpJ7Kkmo9lw09uY
lH7cm8Psr4cq2hLa2YjrVcmOGFpruAdT3icpxL6AcITBabfr8BzqKWCkNuywWTIu
HgEO/ZbkzsDgC0pm9ceycgoosymsqMfTySa2TMBLBOkHuAsf7V501TuAMaIwKR8j
Qx5saTbLNECb+UlFlvcMMPHTUNObNmPuX9FuvevYqzK3i5Ia5gkiqOZ14k46kuNF
x0M1wMULRm8IxHPX9Nv51P51pSt9MG2VDz2aqgvb6sphXTeRIG0UX9ApIIivn6sw
Ik6W8JheOONYBdvzt3VvB6jPWtuElO66Db8jNk403/62g+txboGOkG5YIyvTvvqK
yGEBaiY+iBnzOcZZ2lZGkPAeQq0Pw7ofewiwNlu4+CQf/TH+9v2JXGAyUDYd9KT6
l/PCq8nPFLYdAVOd50G4nuI1FhvTLn+lr0hY/HBOp7wsH+dGU8eyVETh189/Ox+j
mL32dcBaDzZ0yxcVFuBAGpqS1i51b0TTfdF/Jd/l7e65uUe46tpElGVauimTNCHF
xe3SR8U05F6PNYTUx85Ed8rtpsAyzw8W2wDY3l+lBrhTfcqRevGtA1H+Le3Q421g
GwiNKjQDglbrMMxCLDS83DnxFo2brt2qzlMQ7hqZRKO5qpv3cmm5OS+HjjoMPoVw
LI0C71kkJZMtjKrw/KCxQM5KB/4Cp0HFNjyZLjKCaHWtNwhebEH3wOBje07SeRxG
lzVuM404+tDM1fue5VaA3L8qHZm2lBgaZ+/+ZdEfJnMFdy7ER37xr/unn6a5hWEi
llx2wsYpGaJ+eXz6Btf8lTK2zp7beduYNQ8LKdj2GKCGhSKGyGJ5QKLIy0fRw/Pn
oueKHJsOSEWmNCBTwIML8pQPxeMoplWIQUz0uMFwcAXQkTIF+iPBA2SEITyhb9vz
eQrtxTHcYhtK4xIEPB8DLjTkrSBn0H+IqO/iHs4mnSQH9c9ZNQQ8l2bu8JNSZrvB
rY56naz7PS9uNtpJt3l+D1ybbz6gLo9Cm/sWG/wRpesfeJXKflZQlRzl+Kgcg8zk
XzgqRr0almBnzgyeo8LhxZopKln8HBZlqGfsqECgtgrqBPBaMrnmD7qWMogx7a7l
0SBpJzSn5C4ugYwHDWlnAuoa9hBYI2KyOjyCmkT3pLylOYkuG4r8tiJ/ePDxT6A9
9TsCSaa4WT5ueKrA4hu/rf5Hpt3yE8YuFq+ZiAVeocXLjQI/q72083I6IZfxrcgv
W2PtO+wlC8ApcJuDBLc2Y1ryBvKeSY04J6sVpuL6KQAvQoHBaSYB6VVd0v86COZ+
8b4Uz4C+zH89XvtIO2Z8Z/zenpW0525pETRmn/MzM/EmQYEbmEQmVYK33RlgGkkh
95dSrMJp7IsPMBoXtad/YVlO0Z0+UbJpROQz6ffz886XD/0MjBD4FyClqalNp4x+
T3dwR6isFeS04RxKSHr0P6ctuS1pQc9C0P7vooJU0Wic7z/vlL3mMt65Crle4noh
jU9AODjlzr2XbuwpHFOBdicSbS3c4URSARxJozRoVM1wrzDz49JpWe6UCwH1Lh3/
aG3QPXzlTa8/DaEVz5pXCCP6b0Pr0/XJRYjUNPzBl+4L1y7b9f7GJTNCNweZBNsm
JyASHFxFOEdfNEwnE/3GZlLWEu2k5HzbExCqnfor6eTAkr9i39ji9ziapKHgCz8o
bHoHshE+OQr+jABJt4HEjDR5EWeCRerrJgpfaD5bwfMeg2Q66iA2zVAFzSnHyehV
kIF49iya/Th7vuALVE0OpJWZZD4JUZNZDetTx5Zk24bHDDA+ekhxpXDzpz5mhByc
K2edQp9+RfNW12KshJ4olRQExWIg7hr5t1z0oYwEjNODmdRR0ZEdClQYkZEYupEb
VxEgYBUlNDqn9T6KEkxRyveyFzTC/JyLk1cOhD5TVETAgZbRJzeoX7mBkqBdXkU4
ozm4bIbVybttuI94ROWk/dNDSFOP+k8rOJ1qTrNocFKPkVuUGR2IhS5ZSibZO9Hu
STNO8a6ib9fuWieh/3hj9bN4hAhvbxp751cLfzpZKNGTBToDH6QvwLDzzp1NgTpK
RVdeIq26F3yaU5gihPo09j3S7diWH/Y+lW1kunVU9EHSwxgEdIkCiH/KljmqyRVW
oqLv/bPzaPl2Di20aCJGKvEsEBA4H5FYTML9/41yonrIIUmOlUgbTRd5BQGGXcqC
HVz/4ccratRAk9MH6vI9lylswZYjzjFb4Gbg4T2JGzugog9zHqBKUalmQgh8hicc
5LfDVyvFV6k/+ypW0DBqZKttIeu1o2nDbgC+HfGkVD5KzW2rpvrqM/dyuXKNn5lT
FaqX23dK3p3366PYDty03rZjgIfSbqECYxhklHc2QyDpGqN0nzZzTzGfv22zmMjB
XBwWq9bt9LR2xfnbV6AZUh5AiV35ydsNC8cx6JgfcrwAm+xsLOsGvOj3AHug+pPf
FLdEh1sQ6QiWQ25HkTbYyy6UhFxy+HSnN7WSIIoPXgxSzSfAwYjgNwvO+3I1gUMq
EFCsKlpHhli0cgqlOmMxTjeVzXMu4E4W23Ygg9Y5rvIEGRAU3KJdvo6aE0hfTuLS
rOhPaBDNu1U0kxqRwpgUZ6PGG0Vl4jHyLSXLI1o+4E4U8aXBzMDGvvAP1Gufc3GD
FYTiSxDXpCA1Jl3gS1x1YpnFJtU/i6kKCX7F9N5bwox3cWvnlLdrVr2SnTy/f9ea
FUlCnGef1iJvFapsIRmm+3olMnr+yZbKkkDXfW6xB1s585ayAnWU2PwnS1cwYWLI
4if2eGz7l2kYVuyoyDSoorIlKw+bYoHYHWYrX2mhKuuKfDc2I6BiEke0kcy0GDhV
Gz3bIP7IroNhfXq9xiSc8HUJ910kvLWQ4lI7wk5XCZ5Y8n7GO3NWaOaD+JvsxqIS
j7tpwJYV4CmpcYOKeXsOzk3ksqaZQJrN22x3ODtqQU/q+Y0pKhieNrk6SIPvgD6Y
UqNNW0Z9tbPpovEWDWsg71onu4hpsAwbIGmTMOmt8V8W8jKols21JvdCfy6VbodQ
7iy9Hs/mitnU2Q7+jqHUN5zElchRQanl7VrDeB8CcPSWCc2R9re7+tEhOm9qyQD2
fkJ01YJg+6qZ8DqgyFkPBolWn8MTkJi19U/zlvtXrygARlLMdg1dyW9R3IT5qZDH
tYjrWCjiB6EkC+NGqQzGkxpbQs+OmjKjxhRGNt3pS+QV5vUya2222JBsvLWB2y3e
y7eUCOTkQ9TdMFOfEXBTl7V4+zwSQw/cOeB4AWJarCx41P9Ap4puUmKxD9fhYLuH
63ZUQisTHguU6IBUqnYAalfhH6GNVshZYPFUbGvXD6e7ylk+UaP5hUiB7HRrJQwh
/asDoNphhM34YLjn5roL68GglAmbnaT4QzGNSaV60tALC/0pHUAKOHxye4iC265r
OPhSCa3x932yjkIlpFKNJ67+B0SGGqhQ+jHPTz/0h/qFIhesAT6OZr4m7d2lGPZZ
DyYusNQ4FgWeuhDXiYDdtO503Z5KXFdInWYk/Wc/j2rt5GcGhMLfkT/Y+wa6yhQt
j0C2/HB2UqzUUlZSOx/7+wua4jBrIEflal4O01+nTcqm2LV15E0dbve+qeKWgyC2
y7HBdjlkS69CKVzAp+kc41hXNcmZTaMCVwBzUgjfnhXnrqYhwvjXo05FgaJoJjx2
WSNB7gaFeoGNiORS6Opor7ejZY3iQp5YXXrxvZBvRbahWJ1xnn4k00Oix2CnQ02k
W+4C8DrIXj2+EVa8YdsrIJec96JSJyBhPQK3JXeqG1ejoEuABEgUK+A7a5Rafjr7
nqsyOfJPNNRrXfddYY5cK9MJFpMHVO5lvNySyUqtwslqq440AfvM971KBPV5wy+q
CPtq4zfXKiMbAQRYSwTyRtwKcGul2/bchuId1SHygG3vbS0zYZi6hIEU6rwTbpjH
B4q2/7/ckFRfiDVW7LJRWVdxJ1XIFzUyYbsj1yH3ptifOQcWiuxwEOKmCiSONUlg
VfBUaRcaDc9SYrN3u6WSbmVUGHWVpTnmPOfh06ciiz3qTTY16iNpOhVxTJNllupP
gRlMrk2Di0uUW8Io4MhJMRraTcFODuPGLqBVVWjGK3btJ8BVo2fv45hhikyCQxCu
RgAOgm8C6L272iZdGyGXgaS5/GHxhBKh4B325rhhyYvs7F5OLoq476N90m9d1NQq
9ZHD0HhQDyGbAPytemHauRBuaRA0I0Kh4wIDxEClxnogrGKHn20LS87ilEkDI1q4
eZ2wvC1kjXLU4aVmO8MN02V1Uw0T49ah/3+oQFyRumRjLN3ihhRzPT5haE7a8j2s
ii2BB0e+NfKPZHI/V3SKEXK748o6YKCvdBPfeX61OvaBbj3//jUEHl3iqKaID4wd
RLTD6vZw+MxPGVghJiJky0oZcwgDnF68mpjtBPOnaM9iMhVav/Z8e9E1FSg9Cr3U
316pxPvPy/NcH/DdLcsnw5CbLW4IEBcOtwaCb+pjb5k+C9y8q+VHJ/x1H+Dtq676
cep3no868gu1odmcZnb+x2VPXG464c12wjysdHcJvZmxbg6nPu2qOXxQoI0/8LOf
iwal1hudcj9mb7VDOjEIirk7z393YouYjkCvOzY5GROk87stIHFsuOj18c7lnqbR
XASiWe93dMszUk4JdFIpOM6MNOVBWyXQUi+9neFNOz32C74eX6kvbrid0uNzs0dW
x/mDafzaAmzDOLoeHg4Ho2Up8YZ2e7RJusp8m+/PpCFnU0L+PUrUBPuGxjtldrZ1
XfYIUtpegMsI5Af6YyPN3WRKuVnADv2EccZpvQidb6wi7WAxwuuDkPFwvAMovLAH
JQBWkbMtB04dGNqzipPzPlw6LGCHOW0GwFC77pK6dgngYZ/z+HQ0wUrixF5tSS+K
x54zrwJKIEx79DZbeZH0ioxXK06FzgO7WiF43/SkRr7jkb7uELwLGpvyjK2HNhiC
kXUo8GnxBzKWa4LEnN31OjlCCbugEEd2Q1VkiUbDnD9adBkkM5QbM5Ds7/JDfS0a
Y4zF+7H959Z/Y68zkoJoxlrfKBrFpMxEm0A/Putvp73cEVq11xUUap2irHY79Pl0
do22yo9ih4gwVc1aOtBBMoj1XjuNTYKtyFB+GS+3Wr6xorby8kFzzJTN1PMDM3YG
xDWrWziRUzoJFbewE3UeuqqCZABUAKfZfkKv3RlS+Qc1DjHQ8P2tQkUF/d0MwK8n
qXlPVkwg0AvdWMzeDykJQYex+JbuCjBywgiQkUyfFT52hmcNniLEn9cjw4mbFKKd
oWESlnGZDhAg0hReM8vpdZkKoscWkbrt5BkUvSJvbuHi/V8BR/TmtTqdtj8i2IH/
M0V1JxFc05rQAVpx8ULRGD+9odeESksooJGMY+iyekXpEnzNhJg0jul2UW+LwLoI
OJ5Ts1VkINIe3HL1lhl+xVh+6M0HM+oGO0Op7nZCmO5it/qYXnK+qG1LW1vUYGeI
5lcZhfvkoyRHSc0ITUcsEjfsO0j1uwGVPMus0gU73/JRoyBDepMppSXD+hESVCeb
a2J1voLW12N/+Nk0HxdB7oPtm4sYkgwM53sciKT+Z0+AtNI1Uz1PggGil666W1Xh
xVyFnE5bq4ZlAXGuc1mJ02MZCrAf/D/MNWBFNi5D3Ksgmv4h6fzIRUo+rGx5MJbH
UGxgVvtDG82fwYIbLy/Ru5IrQV2sLmoPQevBN5GFT3bDob3JNzbFrPQp3FBIMwvP
BEvpYoA5yjjc5345es0Vv4ueteriUMnptwrWzo+0yTMlEy1JVyMAz/jD/4Pa8VCP
BhcRCfp27Ek3M7n+cDkDFqzy/unAZ2Mxzjv5NXkmsvwRrYT7eIMbXG9lWHmUOtNm
qwM+2UbIARamgdrzcSXlTswqxgTui9TcsoIw528Gv8zoRU+zIGP454V/qH++gyF8
sujGn37EipZbZ/htWt+m/niL3sM+o+ZUnQHezP6JcfKxV8mK5Lx/+Rbd1njHkJoZ
F8vZpnT6I/ZHCkjRdUJiZYwXPzD1T9HvjLiMPj5hyXbKXbl4S+pmCEYiuwHiweId
RBr3DfWY9wKQLCpTcpNvRLAOfNb3P7lMPviHiolww3JQEzGw4dMJ7orSYkQWMv9f
e9Kzv4EdH/GgGlZ72kUjQVS3RVBmiiNsEt2yj1CoJzJSxh+accH2FEMpOrJMnWcq
LzT/YwNUP+XDHx1ilIhY5v7sMTEB/fRzyhVaDUGbqlnXXcGlS15IB82sv18H6dyz
ZKuyzgL7LKSnScuujf5o4Cd4eE/oGWKNdP8sP+QpfYSCWlsTKdWdOVDFXSDxs/o0
nAsB+B1cruug5diKX3CpnVUeOky62Xr6xPzParwkps5RZ96CSBPeAM8Ds8UitJag
2nykjFWqqNDeYI/ZylY+tRBm+Ujaod50ONV1L+hA6eFAHhA5SvYFe2Lz82ittzPv
Z4AoARrTm8xdyryMcGrM7Ht8tlHRJyG4IxS02xd0B6F4zOMYbl0CNb7kVgX/LphR
iEWYt6SDZzwUbOWXv3Y3OXG43IZ5kqNVohLdWMfPG/iOVqNpEBMUNeFf5jZNxBZk
izMzVS7TGs1KFlYMnnct5n3w8TrDgdpejmtqf65cci4T6011Ac0J4CWkwl6PT4MP
W1Jt4nETnTkLi+WZlnRu+ONy7mW29XKZGXO4esmTzqsiv5gKbeLTR3sda4IhCxiK
jTy3eLsDvOMcHY8UGICe71x5iFIAPYgTSXUPDSHGDiDqmTQ+AFIFWCVTMd5eiGdU
3cx2QONkFGZFbCbuRBUJwcO6wGl52Afcqg1k/MkiZCM8iGbnSkqwEJltkPOaFNQc
APOMgsZo6Y34YsX//t7Nak5u9m3qF4DT6K9Miw6tonwmaq9NHzZKQXMrepEQRzGK
x/oB+th6ncHQMsY0EedM9cbRaJlpQJQzTsCFH75X2d40cXFCw0TtYXC/Uyn9+fCh
bh9Ye0+k9ng4dJhvx0ckCXjNC5kdqx9lLxqYMdjjoWerPWL++NGYqoetivFEufdk
ESO0HcEIKA7D3aGiktZita4KTGkJrUEAXUZs6nPRNlcFXQBhYspVXL13fpDBLbQK
9YTnmfdwXZtUfhYvXyv3KHBpBVCYHfgNVyKf1bdVp9jLPlpJFm9kSg9b4vpJhP1C
aOQ2TNd1GjOHeuL+Gk7SAKRN4NQDfwRRjX45BP8mM3fd1iOosRbh82dEIHdneINP
KUkos1BLTxK1NyjIW9JGl+o4CeZ/qctwHkakbxJRHl5GI2x6HzFXmQ+GnAgPcUdg
XPpoTIqtQr6tE656rlWsaBk/fraSX5FCPmVYaABFTpVliiribKbOPCUKaRpUCQB1
9Ns1jyeovmmjFsP3fyLJpDpNBjIcLFeWOadZaP/TFLbnJFaWAlJ91ID26DFdX65I
HS8M2AvKzHEJFMUm2pzrsF93+0hJBz5Z4xct0+Q9qx0xxXh7u7Il2Fd33zQM5iLB
CoKL0tuCEJQRZ17BbdPRD4QEiPL6/qjXr9u61dLPH0PcqsH4ehRkj+X0kfDF8EGd
xd1h4S1lHa37SFKeGRQDiLpv8Osc6Bh5M5QJT1nWThxQFJXqdyvLWTPbxHX/J/TJ
jPcT2FEq8to6W67A1LYftAtIV/T1E4Y0Q5zHbKKa6pVnkomUtQrDhU7+tz0B0W5f
CAa8c3/wdt3Y9YrBBn30JIN9Eng2x5xOsrH+zpT5xv8i16cDz4O97KZd8Zi9oGkd
gazXifeVpsldCTwyAKZTxoKEURL+gA3JTZ+Ribv6NpMhAfI155kHaPN129UqFBhq
Cfd6guWSiMSX3XMAA+oYeRfMfyaEosjHrs2exC9ItBEQpIgeWvqc9v0KJenrK60C
lrJMfBQ3PiUXB3gAbnO7pIsQm2qFQfn1FD1c1fz2wOTGS6P4iHw7OY61kb2K0SLs
V/p+5jX+Cm1VaccwRAfBCC/txWMWYKiJFS4xKOVga0RV3q5kD3Zwlq67vUtf/e3j
Cx/oW8ankKWpk+Vn+8OlAgXQzFVumzy2zjtKxmR6/hCOrh/PJcYjlr46Ld5G6sHD
6mVuEluC/Jyzvs/6NENAB6grLUWGcjbmHTX+EawsDZbIPPX3ovoCnf/aD29061W1
lLky+IvfgbAONcVgLTExece/HfuShz/j2HAwzjxlJrDmUJuJDT79o+9T3Wo2NOwc
h+TjxRi2prSpVYZfctIbppmlsssl+PxocFyDyoG952DpofcXyGjLeIpOjOxiPMoY
OArMWfAIEUmcCr9TRIlTCGeVdWaqZvY6XuNDJZNPoe0LnJmFNpLS2uMB/QZIONwt
GcSiA1gUcCfVOY8cqJ31QMpyf+VJhslbcEYBcq3jShG5SK9K6taPWy+fm5wUSZlU
kahqc8mkDEWL+AcfAD9k3tfn2+lFoYIeZ6SXcboVyll2R9Ap4+9G8S2kPIU8X8t9
hPXnO1bxeH8ipFi9Gzsh2O0KsYB9ZDxwUAAkBthryaz2TSD73lo6Q4PpludfH4ix
CjGhfAl1cPOoWauPoE4/vPwjiiCyqnFvXJsOYPE38JvEFB7grQFTrRsCVHf0x9u/
H15fkBQlXAH6fDRP5P19oxsKQ5Jj6D4c4MOlJil6qTTUNrZFYfoKNOfR99gzwAOm
af3tLtRkUIi+UOSqlLiiBObg/4ZVh2WNyiPw7EFswuDMgIIHclHGkEzDTS8MfbxH
2DkaDRy0VpL0Lyg8MWIxyQRSyVttpv3mPQoZRajQlFLnLSTxvjOutBJUfFi3j1pb
ohLtMizyZ2Ec61bTnjTlzZUSi3oISf5L3P1Esnc7VLamMpgybTP49ScD3Z0UzEMs
rXfs6d2/JGj0wH03WUwAyuC+lliT+3MgtZg/laZag95Y9I/n14bB8+ZOz9+qyHY/
6Ht2GbRTYHmC/PnYiVCuySoNvv89m/3ps0ENoUnEUDXyDLRgfp8lXDWn685jSqjW
wZ27iGwJ5FxvcbCcRG+8jM/3p/Hixmyh/V2iYHhVZREX8arW/hwIVfk7s21rHe+b
k5eaGwjpOMCFB21otSBbd15zDtPi6NidXl9lyoPya5b7kIL2378R6OvaLR64iZQ6
UBZIouond4P9x8l4LhVmwzsDVOFz9aki8W3aOM3BMMo1S4qhKMonsbXxMvwprbVf
TXEKhna0ptroy5JqatdItNtHf7yQz8CmUf9vvDKN0krUnBHkEF6G8NpLFLDHgCMa
jdroSav12AgAAe9ZjZyxOHMrytT7YTKldhLbG06u5p6FWy+eMhnBU3vz6h3LlfIn
RyhSVpv0MDZVeUJFQV3CdQ0NDxSRXEMeQXfUPa9daIFKLUzBtKrrnTSbZFBighrI
lwY0WHlCKFPsWFE9FGEsIWleNBPwBFTux4KI+wMot1YvVwT+pLUyhwV2IiCEh/fz
7kS9D2hZZWB/mY5hfdpP3yy9hO99pyUCAPaU9Yt+4zi/xs5Uare0REn5Ti3m9Yy8
2+go6FsPbdPjOARNI77TEyzv/cho84Tg10UsxFZq1/nWILhE3YrVI1WiBqPXL3OX
Nzf2vtGS22Ke4Cq5uwc5wyo0ZJ7p7Zjs6drKkRuqahvZYPvnka0sriwe/43eOOrB
aZU2lcdOaFT5T36oOK/vw7LNya6biKrx+XP+COvA/NQJMhlwIpmFhHaFC1Ig0pWJ
337NmkAnsxxQ7fs4zOZDHSil0cu0HFyfrt1dDUFL0EZmOG5NFLbkMZyfixkxgbfu
So61Z3Ou/cNQIUEEmd+yU5ULgs91DN99E2l/8gDUe+Iiayi8mHglBvIc3pDGd4i/
2VbjRoqoZwObgBNfp0LXgtwXEp95Vo1b1nYdNK+GyLgknO8VYCntwF8hXErEmFfj
HfNCoG4xmTti6DfIRHHJn3WredyxSEPkmbrgy0q2UQ8SxODpZzaZDv0LZd20+u1r
9wXNhcdkGiU6bWZbfvb+q90uH33RMrAlV3LW9HFVX5hhoAVeffOIXc30FwHGPeyq
YUij6qFsVMunCxE1TLXXJBW/7jHdWeCvA4G/XlGhRKkymO8qlDP4OjXO9iTHKoUV
WA6iQZDYfgRnOlpnGk0NBp3SWQAQlag+qwfiFMzrwXgkrO8eDUtS8H8Mzkh1J8KR
WVtBk+qpHpkPWU3o04jRcm8V2c5156ZJs1K1yHmjikZDPDiMM1fIbde9IQkkB01v
w9LT6NpHleotHvhvzNPiCZ+8wmGEM7rnyBpPVJ4B7xnOexlvrwxXiRZAgOW+b674
91CgDmpQSw8+TEi094IFtTdYBINH/obiL0jf9jMdy9OFR8dEaUhN0Takw5FhYeh4
VrbUH2LYR4QRDz2+qmnjDTAnqSzONPycwAmcqLeHHQaJRrfjIBf3ehjuDo1MK2zR
mqc6s5Lpzd0g1LM9aBoaXf6F+x/WavkEuE47mLf3jd426oiAS5ADZSPThylE4PQJ
w4AiC0zIK+mwYd2GOlzwl0n9xsCwCzEQLcCZL6XBU4CrB75agKBQfPUd2s8HrAXj
VKQzGsilr6pCJq9zftkrMclKh6+VPpTjTvNic26i3uoLqSSpjXOwC0JiwdoCEh+4
19Tfsp3jqLYVyXa9nNlcWH8JaePblSK1t/wvbWFxMQ69KlYrr43OyIhs/QnGzScq
/Hb3w58XOaqZbDmg47TMivgDaeYrUF5UoDnCvwH4Pe1YIvytaGrOUtiGCZeHGbb6
tNq8RLFCRZFXo1OR9XV0QDmKVf4JykCuEk5MWA9ppltG3PypKFKZ0Etltj5NFEBF
RGUE5FPgQYSJmgXhaHgLP+afMFVfq8MBA8NHYn1kFF068Z7O+GmHs6lcKgW09EZ6
S5Y0g2PMgGxLVbR6dyVWMat1SQraOiGUFA3hj8M78OMOYjn1HADZc9BpRaWKRpwm
Yf87j2FIJjeSQgIFet0/TvMD7RWdM3Wc91rpoVgbb6Sfvlv1gVXEyybZqufICD+9
l2OS0pLSXjXcrt5i3OGJB5pkw+D2/Q63p5fed+3hC61/36CfdCZXxVaWDsWhKad2
gFv4x4UZKZeMMIzLkkTR1Sx5nVk2W/RHotYpVOZzvakk7miQng54OkIWN3SzF+B4
S5RYJqdfnkRLAnfvBQ7m5mkMWuFz7XZ8V6lwxJZ5uFmZr/+2sRl/oZGjbdgLmOD6
sFLfm7AQQ2Su4jo/R0DMyvyAlZFjSZRKtHO9fGj7zhBel907Oy8h3LgTPfNNq8B8
M2wFJdlAInuDw4ZOWwa3DZR904gcSzvg1tbK6iFAe4+jPx9qIxeJq3YynOjVrxdF
pGy+mPj07+2KWP+JlQ/bw8r/jbTQToQB8Xv4BRIkGFy+Vp1UJh5wF+Bwl3aFtf7T
eFcNOzMpamYmTZEdrYJPDYIE5+ppQUcrs8foh5hYJykxacj4e+r76a3JlMt61qge
s2Xkd8p3WbvzxRAe1WWsEZZ/rMDgsE9YPGWB8A6MuehC6I+ZZJuYMZVC+eCkSF3d
AMLF7Jpg3jw7zjucxUGN/Rcxd9SyaHMR3WIqeqGu9EqFu1OONfpmJOMWTBlApFUE
wNknILcGfMBKcbg2i4Cjb0DvejgotWvHQDF5VtV23oOUs+2jtWS8S7sLrbQaBB9+
ON74LDEdM5RfjEy+docoAQMYRXEA3kJoSvq03eRx5073z0eXdGuVsVd9TmwW9rkx
qWZ2+UEAgVAH71/NzbV31cYL+03yx7XkAEBrZmVxwWGkHT8A5SJ89qN9RUTELMp6
D2XeXtZqdJchyeE+LDQJZikjiX2tKitDpnzJSeFI6L5PSIq7xaOTgq7V5VMWTyNp
mpznMIiHh9S7ij8B+h4PrVUrIsJPNPL8BXa8Zj6wSgmzD1EqXdDtA+E/+CE2VsZg
x70XmqfDXG2OHQP9HWoHigK4F7lT4ZVOSZvbOzSp6YB+K7RcSsnFp9q9ZOeum4q2
KMFfw1bpIFJvIZiDbanzjijY3i0/44sToSrZNm8YD6bqFupQWnUQDluU7WEHx9fS
hB2jZvy3wme0x1NOqK4BgIbKONFg0tCaD7MDYkJp7AsMVsGqVvHkpjLSkufSKKFF
J07CFBwmVQ/m0tt0z6ecpMyXcx3znK9Ah29udsSIN4HDtBWSncW1UfVS+jV17ESa
pd4yoj1+dIlIoxUSyPBBqGQDsDyeSsSifKXfmUa33VV4xkeNyLKTAF8eznnUzhjt
XticTyyb3U0pDY7pSCnLkZTdWAaq5NbXVe3yPalyX79s3u9Ww28L7Hg4Uee0dB0q
r+SNgXj498nGkyNaxyqka4iMreAEj36dRiK++AGYp7gBQ4nGw6ah9oj/RwdiiV1m
hCawGZpo/Bejt8fUCV8hE/lub+4JPlkFa1JXKTH9bCqjJE0hoz6cV1Q06OldwH4e
dcvgSk/rfa689zAScJ5MpDRW8NmyVaeBM4cLLtMPiXYtw3ZBdlgnKnrxbykl1tZx
PLhtYFjrp7T0NuKtzB42Dv3WQfYODZ2A5mxNBohylnnxtOiM6xr65ddNditVoG93
X77BFkYc/kHgxqWriD38gBTqflqbVfDXJLaQqE2RMFUHIDkX1OfcDeov862xCrNm
pAUSPV/5rRwSBBh7tWbfI+SKqduGGqlW/o1xcTN0wvVzH8RN/VVraI34giBgAUzo
2Q6ehOmOhtoJqtR/eLt0eyJhpgZER+t7eKvLJr0noqbQVYTOIE7KB/xw96Ujd+TA
Db1Upq3slr9LfiIxEmx5XkuPvKbz7lsDaEgzdI/RjfLf9B0Nr7PnXuTPXThqRAwf
OYg95fZUfej0oXmWHbxtRvjfs8DsbWkegCS+D5CDveaqkzVbVv3W6CbbIfcizQF4
VYlIz8bKRVL7HncaKl9MnexLC4EF80+THwMRG1OX3FhEIasuGypxpAa5ixsgLIkO
a4b/3x6MEkWwY3+hLoOLwDIfyiJxlkra/SWN3GWdGOeg58SqoCvAP+9E9gRQHfCY
yfRpPpG9wfnIVC6csp3AjW/JHvffi6fXI5uYTgNLg2r+/RYbNamL0J+qLMimNTwA
FKds2wtCYXCGfsUlcggHeBUlooyrXW2Ng7uTbZ9465vaE1AXsWYjfq782D7+kwgb
71q9H5KSK7BpKzhZJmUF2DR1Cu0Oi8K/KrTYGztvzCSGESdJkNAsfCG1te5uM9S+
Yxa4MgjA/0yL2Mx4Wxogry3schdBVYTdvSZvAVFmMYaOzwGVt7Ga0fIb1UA20heO
WL0oKYj4VNjIyng3zNrDAuGMRNsmH1RN4eOTXQFWmK1RnlEJR1EQXpg1wXMuG84b
hfSwa8gI/7WvMe+5uJFAEEoG7qdGqtJ72lJo0Ko8EbdPDNF1R3Gm+GwSC4TD9WpF
BXfcCk1kD8lzTcPombP5NBxwo5m3IO12xONz0NiE5LvPZX0UidxEthPyZdOn0NtV
uYioQd0m59NgbttRvXnW6hLI+oGLsWib+F2QlpJSSgK4F0VohIhWkKzIVkPVBpPp
lF/XXU0XHVjjlmMaLwO+43Ujsbu/OirSpTnS7v/YkrvAljuHz2CVOAHbV613NQqL
FHuO6fh+0y3W9c8j6Cw7ADnf7nD9UKXMZ2E0Oeq9//8hrCy/rHWb/RoPgz2/BMVn
PgdDDs0m2vIgYZ6jXHcs3YhlZZ2TUgBIQm7tspEpHZaqjcdWKLxN/r3BdjWu+GhB
pB6MaNqWk1B4XjMqatxC/7+0PO6Z/Sf9w2Abi8LxKpI+71lEvtJUblNE/T2vi2+Z
X+oSwyFkIeONW+Ti5+8kGH3Vfx1F43I5fO6c5n+nZpdvNLuEIpAiNQYTvWwYdkOG
FK3vyl7QnmRU6XoqFU1HkEkXmg0z8wabVs8xA/EFPNJuCdVxDbd5jh33UfwZctA5
pw/kxYXMLTfPIwy8BwbpofRJW5RDKkVNoYTBlY3hvs+lNHb7nDAKmgSBeLAZ7hMp
f3j7BCmT5WUmskEpmKce3fUL9Te3XVSUyEKeacWjh7SlzacQy0geuyG6DvqkJsOl
tihNQo7qZMR7u54pICiemW5e/96+aysUxSmLM+LL8kIpxaabXJ7IJlQJXaXqElDp
SlWdC59tChOpiDEON3XQKyjXRxpaZ8Spr9FQ2JbAJAE+L2xZHnNFuZYcFsXZLiyS
A7rhR0PBvfNYBvPwa53qHRuzvNIWawLltPuwsUWzubIUe4KoM1Nn876GNE/Zm/UK
BRuUktmVDp3e/czcIO4uHweiBOS95CjDlClN/q3V+pFQJYapqQveTnq7Xdb5TBAP
y7eUupsz2na6IoX0MTgSw+46TpFWNWydy0ML8Vc3o8QZaIYBxjWi3tTpudwthJEz
4rqg1wjrwPa2v5OFv+QziPV3KH4n5QvGhr3JzB3H629JGDPvIhrgdOpr35wpNogV
+OC9340y8dy94hh/3XEhCSdjUJxo7/4dQ3FjW9lYZYEzcRLCKbi1AA7rDyHDBtY1
REzSimygchm+AmOgngqBjHVr+sx9GXN/X77voGAJJmyxA9pbYjpm14CboOWXNg0q
tEpEpdWhw7gvLjyApKbKtbY4w1I/l2/Cw6y8XS7U97tjVTxGu5Dt3HfAjVi+Gik/
nin1ds1gnNip0B+mI7Hcs/8Crf9EG+hkc5d2SjFsBnXXJa4CvRZQgUncRJOM8XQI
fKwoopcCC0ZUB1WFsJpbmHKRe0N2Nxhlzxtxh6g1k3KcG/ze3UDG1mKl428wMXNv
UZ37BkcDl34CZdzCNsI8csQWgQCNPYlPP5O05ypwnYCyGBYFeqNRxz4QyQryBMep
g+mOAIh1xgB80YOjXsC38hhop9/sFR5wQOcOhsEgDtQPP6jx89exlUCrZ5EvLtVr
m4ZOd/xO17y7XOxhNTF9tXrvEaVzz7B7/+gBksxGmT1RSyrStQiDYB1bf1J8MUcg
CVd5qEZV0BtlJENyi21Lf+M/m3SNwYXtLQRGaFRU0Axn//Lh8jk8S8BIuRoFCVxI
pLrdustS3QVklC4kL9czhqr8lkqIwZy33Z09NWeIHiVBJTbBfVvSFTHiduRtJ7gG
3ehXda6eRiBDZC08iA6hqhh0nUBSX8a3aYIPPNU8zD7VtYojFKjButWzyYzZPWyY
Ys9OB0bjgTJBj1zRAoOLQXk4wfy2bAKmi/2+enU9F/dJ555bN1SjGQ4M8npYvzjF
C/QlYy54wnyz/4UEJjkXsEeCYVsLlCAS82uSNnhbXn+Csn6xMsVuyfwngVDFVnv2
sXWhzpg7a2X0hVDkKK+SVO/Q7XCCxgNCfWhD71nRly/z4q0nzjpOCSb0fG3PhaQ/
8zzHHqPokBSexrp8vyeycnSNZpCqSaEqyVEqo3ph0hxr9gZXyLP+JKme83RRt4oU
giRR9hXS+FAwdcJUdB9zLLrGlX94QhElj6PTA8NXIvHKddHUOQq/Vri9ZjDvz36i
sBFR4XqsXqbKGiSmm5Z97f9M3Z+OM0rgI+OBrIxbGaGFSj/18fKjouOdNzcxiHh4
tbFaRsv7sms4W/9s7HntefHSU4o/yI1WzGOovoe5uxjbUq3cTJ/KH0mrKMjtiuLt
Q4bev7pPiMnfluPsmlk2Htreph2JdWWCKzKLJ5ohnRuuk23BhxWKxtXWLwlnt2jb
zbMxkJnhrIXsdSX85xpH5u0fdQEAoBa2TpD42FgGacoYZP1bS3NB0FnbaSAcTr8z
to/PS8Wm9QYgg39RgyxaSZqu+kZubJjs+NgWvzvaao+7+1CKfu4HfMAljoqaV1Y6
H0F3/xQX7VGuvLJovpXbGXPg8jjq5MPsm08ramhyjM4ioVoQX6Nk1pHLp3Lokoq8
3yZL5kXO3nsRpCpNZCTYRMyFDELKqPq4C/TZX7gWrrxZzb7LOBdmx+HQuwQFfKJS
vO2NvD+VxoaBGPBGYmNZSC3Nis5w1CXU8kbwpHvtydWKCSkhg5+bDWMWC1G++vxa
BAp0tW5nMT5JXwKzAhzMc5XCPvAT239Be0mP51JVWbzJ8QVxwdO6aDPBcaXjQICy
kDZA1vVy8JgHLgmsUaQpxQFK+PixhV8en3528e+WydmWuFoXGV1XSN40/hkSBumt
h07ds/4kp/HctFwVUHMyye7zIlE4X3a6d1YOPlhloGuSGtHVgY1KdzwTVWzQE/yq
59lYI6MIOG4vZrQEqM116XZStuh5UJfkipJI1X+qBr+p+2y4CiY36xw1LSeSccj7
2MahT8cyJUFHWJEOSL/2O3dYPT2WBPSxxmbZzkpqV4nK77irm+qQ7gD1/tebHgRV
nYR7KJQrKTsGxHUaJG6iqab/PyCV6wTSGJdqhiZ9/ZySwSHo7JwFQ9AeGyHZ89LB
Oq/vCBwenqrjFvi7LSwnIGzKWvAMh8ay+W1U1T7I5jASqKlKPSg3kpcNxkIqSTPV
rKbwd9TCSF7VldIcyhoubH9+WWr4jZl5+PLOzqqOu9a4JAoVpV8VoCZ3rnPSR83d
2FLVzoBxIxlUIOabGsrNE5BGIx0HFuQr/idv0E+wS/okDcO6bFZKLLdpzNaxB2fb
p5Tl7a0ZHLJcyCiiL6QA+ZJ88cMi2WV2KgqsCUYfGFK6tSasYyS0fmdU857ezlmA
YwFKMwDllHa9pHYGxf9sMtzx5HXbB+8O17DT2KBEJKJGM7v+jj+Fx/je+44ydCnZ
diWjbHn0+c4fBL/ZfMCMWVFHCJecfnIbljwlU7AWk9O6IB9vyvPLj5qxNty48iSp
tgDa0rIF+r7NqV1oXAk0q7TGvLaKZMWa5BWbnRMpvPYS9wGWWgNytbVfj22yjPIZ
Y9cSqvv2si5ULox2LL1uhd8CEK+fS2tAEIpMBGzqnlPfaIgpRZuVEqaqhPRUPL2H
LxXE2+SR+pWUcQJLTtL2agOWD8xzL9aanud6+ehs5BZ+EvfRL4JEDdVlkWlowfqj
zq701uXz8yvOsWcq4tGaHwuDW4l2ndosWxoBDNKTAtgHS7pnt9wa4QlBneCBJkeu
D65NtlleSem2s4yCAjYdDUcXzpMC3cqsO8svHEkB1OgFVDwNO/qAu8n5thfI2a8O
p0MTAggIg3VAMBJsuY50AidjYlFhYncyHnwcL6nQH/nljSR+9w2EdY73kaB57T65
LsrRFhA46La4kElbFm/r+xg6AVcJsPNPn5mGTDbdBHx2SMC4b4gn0z6L9QAYV13H
eYZDtiqT74vKylTUaQru/2loFKqhWjAHC3cilcUG9F2fBcnXMltvlBOmRGmpXCfm
tzqYAKJ9Y5RcInPT729WJ7Yb3PfaQ57blbzHWx9kvbY8FzmuViSK8mgH2Ejm/fKr
WFWbLaEmUX1ng9ezoaqWsAKaYjSm3QIYUK7qPTDmQ0uvRRPAjaIKISV2jLKo80Gp
1iQpS2qwZJ/Z7pquS9ZeRGnHUtGJfGs0Xxz5KEPBrp0IC7GqiWAcQ9HQPZZ8r7Ym
jSj3ZDMpXEjWCFhQ66XpwKPOm2Im653zekU1VCHd19pu2VJr+mgY+Zdfa2dYaIIR
K56lMv+UEDeBZfzTpouXN67wxpyjFc9qYHSH+Qja7LV3Nf0Z4FXR1iW4Fil9Tf+C
7HvvnjL/ybSh4epyHnLLdV7gxLsW9A7FXdrcV1fDcGuIE5QOkXjebJS5m3kietjn
R8JY0TKyRSFysiDuwt23YiFNLtVSWsi+6RSqmM+A9IK4gIakWnuZV5ouhualbXHG
9sxW2lLBXFssuHVD2Wz7inoSIgSPDSts7Duyi6uBk7n/XXXsO4B04trPjbP7aLBv
WgOYWnrCr5Tk6DsVa/zCMR9f9qdNbyyZkOOAuTClu9RI+bLG5R+E6gs96khC6o06
LCQCT1U/aHabTwIjERBoZDRX79KyjNkszEH+mqz9FoiP7zxH/nAYtQTtO9yhQFNz
Rw+VSqjJwk1aJvpwG9L54o2h/GG/MY//cou0a2ss8niMDC6Cjm3EpUVWutFPdwOY
BJl9lYvdZv282PB4IB4yAy2GeZ4bKjS0VIqvTxTjRD4eTIxdRCKIfWsT4Cq40mYo
7S/imSsML6ukSmd5wy+9YX6ez7fb4OmnlJHTbH5rhIyCujYvyP04PM2rPDAGaFLs
fRTpvXUkZOi1yeDdAQ522VvZa63+xqa/jgI/m9PlPP+OFCRKNbWV0Gqv3CF1PDpa
hZPNUDg5sGcGziVKXmovpoPf5OBxvkIH10Fh9cuZBJJyTiVhqDOCvIV5ffS1vLB4
29Qu6RpCa4fw0cohztEDwTJAf/rIn60OKvmwlIkhymOvMmDJgw86SOu00x4mwsyG
8MjJw6tHdCTck3RJHKcnZ+9dZUKk3m2v5/PtbJdkraWJ4TAwB8S0SQLRIQA4vss4
IttA+hd9daBbpT4nRAGQQlcJcfMDyTcwBgeA5/h5QP1KPkXqp/Qhr3z1q43KgFbZ
4iNZodpxvrt7/DeLvXR+gJmmVMH9AxGI80MrXYj11HGRCEvzv1ldgOig4TOzxJ5I
gBguGXdFJfLradRF1QXI951UQaXpyekiG2m4kwZqMmpT0dUOTbdoxCQ/ViBF+XsS
p9+loQpqi2bxFC20ZkfvXZdspede8VOUh3T8Inw8HVwkM8J0szJEqaIwcEiodUY4
4mXm9F40n22XUQsq9/lRnQUliSHvGK2jwyk05eBHtdThPUCdgjI7h22nSnumV2vR
BNE0eNsu1L5fn/qmTdqaAWNDm57/fgBUUe+ea4JBhvzV2k3Z7qbIIYbXLYXooDow
frzvzP8tqoRGVUkCsl9eGiSWBqZXfPkyC4fwf9PEenc/2seBA3TviHtPJYlAsVB8
NCKhI+PoxPZ0p7N2ntrjpNxrMRcogzEEEvCQAkLqx+5NrGBqUDQgtysiJv+uHrC5
BzXx5DI+HI37NNkWJCM/G96R+5IDCuU09L135Tot6Y5Qll0MRuUcyAyej4lWZA8W
KgGXVG7gUrnebA5F71aZV5yfeRWn+hTxQ7Lc/jS42XhoPnMewvJOUGHCOplrHfhz
5ycRn4BLvVm8qdezuo/oi7VS9aExXUc0RtIcyatm1KdjlXnXl29/lGMBVcJiXd2q
fUuu8llWWHGYyMHF9rdjtATYqHn7ZPjI2UOJJP09cCMhmYi1KzExtvR/A6e2UZ9A
TszJolzxpKpTFDhSM8MDzXrAHBq9m14Cq2Tp2oEm4OJ/T4bmm7BMSrZ5ZV0fmc8m
V/Sbgh8GCYVtJlvh6JvPjj+GijL6KX7JM2P80N0Fc58GkbiKOh9rCLAmtMV40kS8
34KuC9l5G58ZJp+ADIvJns1rU9hp9F91iZpb2mKfTcBYQrsaVb/NzGMqezMOWvmp
4A0lZ47TX4bDCFK73nr7/VcU5bbnO88aX8nH2Cu+O+rw5c7IHnl1NwxofGQRA1VF
gjvO7Xqzu8f7vbd2xymPp1AEHV554+9Q/rBz6LCaLYZq64qrMvraFLL6xnw/ek8Z
XhMJLl1GXGG4MIDBvRoRfrqlPAAJZ37ZVhm/+9r+ReGYKDi93Pg+sFXj8s/chiOt
MpwB3nYF5iTuhHY9s/oCLmczr1h7YAy3LxBMO8/8RDuTSQH2EXlJqTrtHYqJdaNj
oTtFf/BWhuFgazAKgofwZMFPCV8nvSdJFaSqmPXhacQ+oSlJqk1xHKz6yukQt7ve
Fv44kojdznguFMlF6zMs6O4Bla1mFKifTFxfPLGX39ngGAXnPNL8E22bKGSMjg80
PYHLS9RHviQ5h3nToJEIRoyThT+EZcXlBZ/v05FchUPSrYMisMDt6KBlR4tKt3Cy
W7tUGxEQ/yvjHiLW2NNOO9CFKCKywftm+St3WhQn68QYm9VhvP3HyNf77WcxVbun
7Y30aRcXIc2J2ewz0tE7Gbq11NRh4xUDTHriTLtafmRLcTWFEyFXjqmdwyt+qOSP
yBU46yWfIveBvqmma4IVAEM/VsyVCEZe7GS6MT2CRF+DHpAEyTGpj6kWYaXXiKfv
KBifzXSFmcQ8ikKApJeAO85oaboVSBDOzWcUgrIoKDM1sB8tVYuy5V4NnBb9RGtn
P5I9CeB9hzefbikAoJ1XgW1f//bRe2ca85FfF4ptWbdLrwWKqi6m+umsX/HXmiWs
YcTxt3j5o6avs0WsudDw5Epod4e0Gc/cshfTRdGOCPvFiqR3gOkzM9B4LX7xL9P6
ME4lS6Padlq1Dli99misSmySQkYuOeD2HrUa4O+iEGeMkx9FsSv6oWgT+hbGcyHr
DmO9u9rluKegkhYBBaMIY/YzwROlgQSPq0xktTNp/LubhBCzKWXjF4k8vV8uC1wG
gCMzzo7UMNrGtmRGPHzxohXlydw+EyN9+LpbxonMyw6BAhHJKxAFxbvQ1F2RGf8G
m/w83KFboJmbvfT+T4aSFRviNnCljZECa1fXwjjY570qUL74mdPEWZeYJXE66MDt
kzAJTSHKRdEKxH7LhqpkaXJNXauOS36h7SMJhwap6LepEj0eJJ58scqG+V8iUCJ4
sStj94zmN2FAcPKnwpd3Od7NSt4QwtMEM9b2JS2m+5mLKkInColIqybxCQEFbZKd
iHg+SKs0GL9EQSzaHAunHSJXQ3dSz3KQylA/wFpb4hQmSw/Ut2E8yeFUyuCZ9iVe
LWEBYbjosBZ6g4HUsIxPWoAxAiaImGOND4f7oe3uEXiQVuZtsShgNj2+j+5e5+E3
bnvxl68euMZyw0s2Mo20I4UKqZFuS8pTI+4kD+MMng5iaum6oJpg2EtCqROl5qU7
MWf37EiVxca386PfKK9vjlt204E851QdWjGEfZmvHFXccCrhCtmrDx3sArgrXttZ
bFo/JjLbo8FXcKK10gptHGAYOG4W9q42VHYE2cLsZQhhFMyICCM2tQd0Nl+pVXMY
WIh1TTs23JJ2nl7VS4D9/7PEvlDuoPZVfFuUZFq9Hv2+oF1YyDjjlN277OfEe5g9
jZa/bE7rOl3/cKXuAa8sO71vaAxlpf2D2KriXAhlgCfRfiNObmDXXAFUaiMCYcaG
wNr/QRdkJSI5YWB4EXmkfFx6rZz9lrk/3tlNUU4KECcVCKFssGHaznKcDDaMHpQt
1KmaMwZXJUNmOIpuSC+ch96ocO0Tv0evixBRxcEgXOp8yYUDE92fkJ4z+7RtNKxC
5keyogQTiMOB5OEwSMERTUJvwUTstQdiaQgWQkcDyVUGtwmgNbGTR898k2sME0Jp
gTeFMZR5uEHqh8vsvaoepjlwgOOC7UZWxNxzwbZjRHg5m/jTqKdKPxQmsHJ/bH37
0BlCmiksvVHrAx2ddt7DsQw2PPDf3kzivUslBsEiHmD3IF5nQbuUdVk5sWhMgtqH
vPeExe3n3Yy4CeNpvG1jMivMhIlcawnea6rGLZiXhY5IFn3eWiPJF1wzpY/pdts4
LwVUZ7Bmw5/Sn1dQ9TJPIu2KvAtHA1xBheJyyE4eKBDKsLXBKf+aD0JEqwHmrNW9
LWjeFDNK8VrKXxN9RoNcdPFji/WI+34SEIPuoPQMNuBvoULN5VG1maCPAkdRLBFy
nGJmAlIvUAvVO6l//xLWghExr8abIGzMjUPockf4/N1vHFDaEDpxKwQHBaqcrJWW
9DLJ7lUKefMjgviAEs5vZcIRZsPtYSEkU3vajiECnO3gH5Ar4Q4DCh7u/Jr2e2Dj
IfkXAJ+WRRAheqBFEpq3w2GxggXPURAWTZmv2bX9DoOemflcUytTiILJsEVq+ipZ
rvPawBmcG3rtrW2NfzneEstTubnmDoY0LIYBarIz3VX+mj/weAjiCvuacmNprXUI
81WmIuIweHoBZLcEQQMYwCJch0QNtM2zLR5EciEMli7JcJ/Y9HzQPTrljPAdy8xS
lMu9883rm0K9rniUznql8Ztg638Prh/ueBwhFeMzwaUd6s8o28e1aifveaglLxwz
2DL0WJqCCCOKomFmLd50pGc9ssxjyIXanM10KEwVrEmrXmlPxeEudVImEQCzliKp
q83B5KlAyQGRC7THdEEVnVB0FebB9Wj1Mf4iKQN7Y0Vx6A7L7en02lXXopCBJGVC
3fGZpND4Z/d2y6y7aqPMD7DBcz1tuRbbk2jTZkohTnw5VT1jcfl0jqEARoAjmn6o
2rW1IdaS68xgRaXTB3O87U3eNp9HvNlViGnvAwC0HpjTA9QOel/fZkm7YIpN4fKC
00e3jRm0+T9l+BWvzQIuJK7g4XbMquPq0LYiLVRK38qUkI6FBZJajB2yY1mmGqBm
CxyZ0+hE6qphCGXbpqQuqlyIdfk69RlQ1aDR5dCJ1UTfjZohzdrstPlB7IlalFr2
1pFGa9xsYsqLFnZevb5UMNRlo7TeYCsTXzc0EbRnhfEaaVvFJWbGsWwVePtCsF4L
b4Tj8Hy8DJj1FdSuJpOYedDdGw1is67gyOnEQHTYqTWXLJUO2Jyeg9w2m15tAQ2f
Ci/f5PHpYEDXd3Kb1dQwkw08gRdz1lC7xznW2Seh8rxPWFiMTtcXnMikHzpj2yhR
F8auT4jIJai7D7FGcIINhN8plB6+eQhfJQvN5hq0cieke61vuwq2LgZJD6GK38O8
oZ3Mn14fmC3nVXSFWvHED1Fje6vvLRkCGh8mae4ikvQb1RBdMI0YyY5TdWfY/ifP
PgKrbP7+QDBtrn7ZVlCFj63CX1HVou1BNuCZra1j+9GCQAl76bBSHSeSZmGK/T2t
XsXUe6bdKAGjGfSAqPex7aia79A1utxaef/hZ+XWk/hqPqxVi/0qJbjpjxK0Y3iH
XIj9nKd8nmqoiKkyVhHwF4RRrCFspofCiDWV6oYRaHR3zQiIe2h1AZ3CNf7+iG7A
guRz0rKS279A97aG143wTjMpINplGQ2XZO5vLmYfsnb+zJpHgahEXBrQUCPMPUOz
LQoZ19CKEV3SguzpHfJFY/uhf2W4Uj9GJjkqAxbnUAMFfTgq+CJ1tGPr5TjNL+lv
l5FbXKzbzZfJTBe1vvcAPV4HSf0p6Ehsp5681F9SJQXiSwSvfrlu5HsV4f++fGPa
vh/g7M1n7Z9nKRTxMiod4BIJh8QAMbaf3SsS7o3/4ASFzkiqJGCaVQQIDFNLQmgE
SfTKerJIIRwtJ3fBP/pJsTkKAJ+gqmjFOpFcG/yMozeBUr0c5KGr/JLAl36xmRtB
3MplUF0vpgMNdTXQCi164Ypmxar/M6uDBly9dXlWixPswCey5UDOygFbOxGsTvvl
B3VSNewOEliOpqJekp4Z4N41PtlaxrEXiKViN2cIksoeSyqtoGi5MJ/WeUQDLqZI
kBh+pcLAOOyJM0QDff4IQK6NnXG+awJIuC9jvP9hU/LW1hJSBY5m+K7lcaq04W+D
0fGlyZwG7EEGVlP9YdF7O0HU8PMoBb/nNdljWv+2jkVjHe9J0A9XMPbtZ0RaynQ7
dPmPk1DPkrjk6Vl7MpEB9DP42FYJW8rAJKk007QesbJNifTH08hzu85EJ6FOml28
3G9VNL6Yd0Oxlg33MfuWC1jNBD9jTPVLqShyXW39IxS2RfiHvkf0IKl+yYqva6vP
OZBAUUTZwianvXIjtYGbMket6hGaLOPPb0AUYEom1di5tgIrlpFoUv02X3R62r9Q
HxtjZsu4J7GlMzGHFVnmoCbgyvKqM7oVilhLgOrMiYof/pFGtmixJt62mQRowr7B
NsJRc8W2xL6xBiJF/MFGccEJAvNTkvV7S8nf1oH/iD9hjbhWcV0VSG6e+aOACWEu
ocHbzz9+L/S7h+UrAh0oBbcAJqsAohJGDaS+P5lm0fZpomWI7Osrm8BkZTvtia3+
sX+DnCkQjQUzBfu4cSES7ez8+ddwLevPoZpTFfTCdB4K5/IEkk5oYjfFDZetrXRs
A57jwrAd04AiQ8QiA5f6tc7FoglhSQAcG2ICLSlv6UgYMNDNY+mmVFLn5VVdufax
uhXwRugUUoxsNsQpkSGLvaASSGiGJiHMO7LfxDuzltNnGB7kfguzFMOuQQqvmGeO
EZIHoMeeWXUinidpuWE8ppk74bJJ0+qXPkO04KwcXKXDrb0gj+zRhDWeP4gDDKGP
QPiZENmFc0CWMykQYOwEhUsIhnMWZFOmokZYCJsFXUvniNTlri/PNTPAaEdjyCBp
t9x+vH+RBRwi+Smlfa9NVlXrSnDqYp1FIwJQpJAbv0ybxhm6l1LyNv2+Nl07fZh1
Bxlmt+AiMWMmG+6IHONq3lzDatx0OFqSwcb1ke0tbtbmebTvBodDDZl6rf1IIUGO
F/YDyIcABefyS0ig5yfPa7dgU2mpDo31/0Ip4YNPbLN1Ckl3q0dMEBwqUks0nIMV
eiW81l8vORnqSg4/NSL3g4c3DljZKN8dDTE/Q5zhbvzZetaWMxQly7eFRLRFHAIu
S1s9/fMqqIPGs5FagIlleZMX7F2Z85zZR+MbBkxCMZ8WlbYcHtfnEec4bgPChjU5
lkFw1U6VOMF+mp+tQlUmW87t2ZWO8wnWftG5yAb7/yb2aE8Ogr4tmp7Jj8Inv7ug
E1Ig9fRvx5C8Q9kYYetQ6P0UWUw92zW4qeEHCQUI7PBIUdlrEPNov3QbIEOqudHk
MTyLjh9Oa7VlcFMa5OC98iEdXUI1nZJk3OizZhu/SRY8HKznBGUxFfxIc+nzDVuL
LDCoazmwEhWHdwqg//U0mEdZFN/AmJNc8B9J+DMH/0wvk6Su+Pmc6kkwOh8KBJUi
4vOb3MaKoaQJ+ATtYRlGKxq8hlg/AnWX5OmllPOs5/ogT7qXGMA6FihOtM2IIHzP
dLcjfT15ZR1a2PeZroK17pGwtYfpNgcKHzGJF0u/obUGvwgc2P1meQYi6Jw2vfod
51/aeJ2u1uklETG+KEv3edbkOzQ9mKRZf/hrD4pw9Iw8htY+cYWjSSc5hUR1tB/X
ZVjYtiRZxDG7l9ILADbBGOXT6FWkfYrqMEYYlZCq6ER2DSDybyIahLK8kDBdjwZd
nxVrM8czWXimhVs6wNoYjJgOjG/MwBg4ECDAekSKetuyHzH8tI8N4s4qNVpKp6iy
W5qKBf8coLo21h0xVnre0PrPlMN6ZjwM2QCI0gamUOeM0MCgYYKA5lGyZcb3Jk4z
2vh8MRNXjpioL0A1p5S0ui3Nt9su7QMX8tf3hsB2y4iKg0SCPrWq+8KXvdNuCGtj
2Yw42c8BFODs5OodI9foFAESs2Xa4DGBnQt0+xXTU9ydXJt01M/Y7V9uX9S6F3rC
OAd5BZRr9sXeKkqP5c8ekegKle7lIbJZmtSjdCcD3vyF/7ssnYR3J19ewBnWqMNy
HkJBaelHGjxNAtzUNOVvdGUtizmeuRo5ECo1IAdQt4Gqjx/e2OuBz3ypUk0L66bl
oK0quVnXaBLop9e8jocxctYQAK7x+A7tz42m8AHUDEG67qDw8M2828PMWpEDTsmR
dcEUpd4lIhGi8nPVKZFLbKhqIBDWF9JZI7yoJU2WDQvxbngOWY0ESspp95aYr1/s
gmd9sVQh/Dzn4Lzqj2+heTSEsibLiBfI8vWf8Xsqzc0JH3uwpx33VD1Rdy52YIb6
as8MLRinWqfZs1hwuN1dIJWeL4GB+IoEhWbAOnwSGHnOvODH+b+OEvWjfGMSlrTy
mthGATynbinYuTZfyUM0iRiXusXR5cR0vvzwnPod4y4a4qNQYaOBEy+rv4JoORgD
9JXjc2IcP78Bgc6EbH+WG+5bok/V6MpXw9aH++PXpc8NSmAgJX5PmvQvLiSZX6xe
m5SI2Ia3JpsBQrspJCXHTE8dgFzaSbgbBCd0DouMYwizKco6vBaeDVqmlHU2dGci
+rGjNX2KmW3Ul5xBmwoNYg78VfUlK8GAF+tyhdCqxWWJcnJ0DJbK0BlhNWbOm2CM
UUEafvqA1ki5raXI1+vz8bywuWCmlR/so9TpbjDCYIeGGagJsCwf+TtcRlz2mFHL
4TC72tpAqoXsAdvonPc6pfPwxazf0SIrRep9vkrhqjr6M3OWR6MWZIjgNjCMQQFi
LLvzz/btds6IbmStovjNSqLPOUCAABf4hqSBXTxVdIeyBNO3HWkhY/a4lmDMYHJy
+ho4OTUbUeaVbID/J/WM68E1ghbhDodXDlC3cENF5iwX4t+y7I/XeU/DEiSuIjpA
O401L4sBJ92QHgUH3T9NI2h8qjDyJtn9gSpDUq0Is9bg2/ol29drA2DYGq9VF0XY
Qrx4fpHvrCL5PZrxCdr1YSXX9y6grOb6JnTkFN+qMaT2FiW8bCKKUyPcT/C+dIHr
YSbtgx0uEsEl62MnGShjuGVdkp9AFqzEgKJRPwsi2qIWXCKtWIwYeFxi+WP+S2K2
TJHyAaSee3n+uquYeYEwlSXx7S9z5XOc/9ojjIMSI/VOtbMCsnwcKjAAcLGLyyxk
GRqqJvd9MpU2qj2UzzRG2MO9pCG4CmDsIt7A/0NVIeS4P/zq0jEhScMVqQE+Zx8t
YgVfO+8YZ1mTez7hLAjySU/2m9yr+9vbZT4KtwvqqKfvzz15vhMoYfB2nMsp7oZS
tZ2pC37zbOCu6mk+3Clhb8uNjaFM3xRI9wjYjsYqW/GIfzMLbPp2dr1bf1j6j198
V0sRlMr6yIbl38AveFjwMhUz9qiEsfhhPn2YssbGefdQ3WHlXhMSuyGAdR4Q9oR3
+PdVwmA9rywFvwyNgBSdU2Sn5u5RLDwIkNanWtL2fAucnICx7G6rD1cYe6khZPd+
D6hIVGssXexCjCpJZn0zdPTf1RX2oiSwIb1JulYUS0WhK1nyFAw3cb9ZusPpEkJo
DBM+2ZGMq0ZxAepHvDoUYda5WYy3/llgI909q44cvhhKkLWB3iUc8nOvY0T3qofB
5REZV4H5feUJsvQ4U3akGt8W5LNJ7AVBJdi3H1RW6e5fLSJ9e4unT3H6qNdRQZkm
0IIWzMswWrXtreXTnSiSMoq8LE6gzaTJ8IYtM5Yp/ZsYNXWCh9s+Q4z1IcCQqIma
0WwsQQjRecGgfROFXpJyQMbxbjqYNKdzrlQAtqdfNXyWlo1tdjnl4jvSKuKbUYZB
ndaoRJLe2o6b5KRSjYklD7x082SyKY9xIu3ZiGy9dN9PVOr8AFecbZKl5AlyBWfC
TtJLc3LfhaPLJ7sSOISRvaNTRf0+t8H/CWwKjxdqvjb8tsSgELGdvmAB4h3z+SqL
U4iqCeZaeESr7T/eW5XojivXX9THcwuiEeSKon2jzVIuuiAGn+fONMYC3c9TzGt6
5gZydtTnPX4UFhXAFxgTmv1ciqAN3nWY8NzvWPfQ/5bj1qe3gNQKaFJtw+gqH0aL
Qmbo5Kl15gJgjrUgjP8xsn8ONGznHGcKl/fPO1RUFvJuT5uNvEv0Z8rdTE46S4OZ
BSZURts4YmbVRu9nIIQ50r5zfSsRVxn40VRhjYFhdw5UsKJWtBtSjvT1qQ4Mwqk2
ymjGCmicNck8U4EHaqFiGy3B+R8/XMSN8orHSoiGsuCE65jQC1+ubHsniadFvlxb
o8r4Z8ykg3qKF4sNBEXlczSLWCcqGuJjWYWVDA+oaZRICxGn5Ask8HyxgRPcOlT6
ibhEtL75pN2ea1fdnd26QZXLjQIpbmIdfKF3VevG3TeyYW+ZVocUFdhxJn757DMp
FJIuIV2oXMVo03pWmY4fns0PErOFBT8jIm5S71FRl5eB+esg3ms2yPBL2JzeBu9Y
hbradbddTYRyCZWtYRjbJFRMSWDXU1sD57r4siOW3ufEh4EsnAuwrZ9+zPnnp7i9
KDffcip1IOdI2KzvIHcUcpXQTjOoxFlaRWyEkKkwjnAF8jv+pQuriEiWb9u6MXUW
bQogxc8rGDBEHWCSZllrtUmqIuCRxTZmdhJuBNS2q6zurU8QHwMMgxxXwC++IHrG
2AyTJmOgJ7IBgTT6V4cXozWCwWpPS7Gh23kxMhIbrUAfR5h3cjnrJNuuwkGKrwbs
rnOknYefMFclbnkwdWXU2v/puMlWhM8UrXAagf92iaqN31sZeSuBZls4TnTBDxBS
KGERiGC1CGRrNLIz1s6HYSqp2uOInaZeMqTUzc0ER5ADmx5qSdBLs8g9qDtcn8NM
yIQyeV871XXgKyXDXZDokw7S0jZfH/mIu6mG9WwTmlToL9/6xzU2PTZMyFLHtSnM
pzyMfjxuIZB/t5t1Ul92K5w102sBBglJua9+7b8UiAXGMNKkRItNdf8oPaau7haX
kCeZJVaGHha51kjDEsoJ3xUCE5QB64o8OEpJCgJOIfYYF116WFkyDJoObrvI7Nmb
3/4mAFJcWDsC7iVFEfTjqSZPIPQTPRm3D9c8Dh4JXLTyAbfM775VNDtLjrkP6kEt
qZOzALyNQ99LSwQHBc9AcRqPLjRcev4Rv9WsCkD4P19J0b0M4fWVzXJLx6/+XhXm
QSkfcXYbzjndPSHCbOyYIi1j4gtmRWifc8faOQISuTWhwGJcdZwDA57W7NtliERk
ELMRkDUboCSx0Z/zFlA7MUrTsQ/QtZXOFNPLgrA+fwlLzPLjrIqmpNs605VZ5wQL
LMNLWjy+ZZBcieJZIOyVvpXrHh0mI23xCSUPsTcIlKfCNXVYqJD00oJx6K2CbvyW
tRRbyyl0ydaSjPzwB9wEJI81MBzK+qxKd/fA0tTmT6oS/tMYBJPDfWbyyt6h+Rjz
OA/lFXxA1UZ0qSa+uUSM3CulOQlIvNOEfdqZ48FkFgcE1IqsaJ35HsrapJiKFeSK
L2tIO672zVCi0XAw8X/9yjO+3mfciAnJd/K8LT0MewTJhknX5z11v/x3S5OMFxOs
pN1b6MJbeNVFzo0R12YLjuLt4nOuA4dD6XiHYFn2vP25A4vheIoZmAZBDzURnaaO
I2OKw0ElKg0hnZmR3y2TdsNpMSlwg5dG2DXIiePqCikQDNlHep09jkWlVyyuRxAN
bRzfB+pdVsNY6MmV3LZZPwAjdg06aDq7XXXn847NsgGMFHC1KZI5FCayYbssIXXu
cyz4hwgLZ1GdUhNB0rxJa86dllSUxJCjhMp4CzgKTPp+c6cQYyFM4g89BlVg2265
FlwWgxrN46cQnzbxY6nYv6sZKnuentdHZAH/qMbZncTp46eMrAURCY0D2r2fPF9Q
d0/r9mfaQUiJyoWcX1xAlAoM+7ZLzRNJpEygYXy5ZAe81PNcl5aVnw3369N702Qt
s0zNWPFB1ftxXBWsRyI87Cy+TbFZ42C6OEQB76yKBAfyRsSvAdPTTbigLjGiGIgF
0fLnVPO7vbAwdKrH7dAXdvGU+9GgTOFxtvtAVvSj+UMYW2TsRvHOcCFQMtvx1laM
QE4vi/jgR5v5SyGNhJ7YLm0/vOQjwYQLIoCwOSOjOZpAM/ZzZ0QWDKNQz1yg2YVW
Nf5NAU6zCsKOCXVoeF97ZlJ3sJP3qkV9sjosgn2uFMAdao9NYw8TxZqhi9jFA2Jx
HNQjgRzAtYswt+BO5FSFDfERuZI7UeZjT2gknIl5mzCR7EnOOQSAwvSw6/qzoQiK
DSL/na266sZXph9TPHkQq0XUGt7C1S/EsR45ZJe1s09QzuY1w8brFtSF33JMKLlV
nrkJnLDli6/aw1Tuv26pfZyAWTqoi7n3y2GhdUerGVkMRS7Zj0OnnZWMKUkdAciY
OhFx7IUG4rTcSRmZBG5fK3XXhL2Hvxji//bf+2rUgVHJTHmTEf1E7wgip8Ntjfzl
ocEk9miYsxmrM6Xtpa1V+Bw3Zz6JhX1usNu6vhcoxzQSEYu5xFe/Ghmybse/eyLW
uJxBgSJ4gAl0wufen2RzNf7+YfpdEl0uOVQcwQJWluPH/MvNcqin3Sd7lIIS9KP1
F8QXxZn1xP8nfe587/2gy43nnSXddfe6sk+mE65auuN5IyIK8LtQnNAB6rjQfnXg
qkq5SPochAa8F14rmFxoVJDyyvfhx5QasW37+EXmn2gLdgL9d2MAWoRBDf+PsZ7Y
uSPe4cNXVI3M5W2rpSQl5k2Q6Tj3M9pgfTnjjBGjMYxUPCJtpPX214TCgNSzWmKn
MF0Xn5isrxsAFzYG1KGIKr/s9F98W26gx39rDAzLzZWARzaHQy02fcbZoN2uF9SL
4uPlL3BX6IryhY9TuxSY96Ktwdofvo87XhXmbZpttLK0sS4NmSf7Q5GBKf4MMJ7I
Y+3lOsCeHT6KF6BwY8iKWq319d7GiqV7oNHb/iz+5ECuQB3W3vV5jlZ7nwhUgPk0
GfmO5Zh/o3ZVzkU2XK8EzR6jcyrBRbjkgw5bhHkQGCdvh3NWgWsO9JrEvh4DuPck
7lrKKRwm4/nBWuCdBJtibYJmFqz1QFUATgJd9FOSi3KGCKJxSXCOVlO+wOhuITkc
Hzx0Zj1AtXa6G26mKi9NHKnMblkakAtmuxH0btkO6aKzBmRCqeqlPOcmQQAu3CEx
UEi5Y5ih9GWUDO6jQWucfKsUZHYSTfrDyizT5gm4sBIquCkVVhj2B0H+gFtx1Ei6
e0I3T7+WbxAVquWg88nA8/jSO4xYFiBrF34Jdzv8dNpuytx7wVS/da5xjgdevLe0
K0yMnFDfX2rmcAwH5hi1OWdmpEva9Zh0340HJT9XOGKuYallD6n/dxATdmWDEXQt
8+WAlUHCi3IQsAGXLHLyRirylMTLBVKsHJaVnldDmL33zwSfwpNxmjJepN56ECj0
XVJS0dQjFuuhgVB0dT0qo6ICgklj45iDhymmUG3EfZpubx+smkwney8xxIe7OeJc
JcnXwDhDbHcbAFrjFou4/g/kyUMC7VeK6Xvo78pakED/gvqJytFgd9lElU3kfAqp
WcTefkbGg6dmrIpF4qnjmisj0h2Ia731jYTxKT+sLQUryfaNk2sXH8xxMRFCZNKq
oz6yDTLAyq/oZYnkymjrUwHSx1WEs93NSfnl4MLfphFp6w575zUV+3mNoR53lObU
OqFPGnU1RbRhuFbN6G/HxQvbMLOLBHoHe6ZBrwvzOt5mRjs3pnAe2D/Ya6l+e7X5
IxaDY2IYGt74aa2ndaS4wPAD0X3FkycvRu/ThkXVigFVc4eW9MqPmiPp8nNxS/HG
v6ev+x6eDt5y/rRhNuj+1cVv9URWvRGwnis+6z5IWBWH9iUu+rV3FEX2730kV2EQ
jMBlBm5dl68FwRFrcigpg9d5IB9Oi5OTIhFbtyi+tE0jgRu0GyzJzEk6Lslx7l1r
LoCAkf2+hlFpMW9Lg8N04FLSM/4wLIuzy2nHs9VKZC6VlPX+RPhlQQjaZatdwjxt
aT3S/aQOR75pQr4wRjFb4W72sY9o3dSERWjgk2fzlFdbIxtSvqGBwBbk4535xS2N
7P6ewHqtexqQp73AJHIoWyD8ZLY+OYO3QnVRZIJxgvxYOiX9fC/Qdm00HIfmut2T
ZNTJNmlslvXBaMXt4h+4t18vR8/PjbP+OfC2bty5943KXmH1B0l0oeSb/bRtZIq+
Yq1RKKlAczw+u02CkJnUYbsG6n0mv3Kr0Q7ZGx5HuGzz+gE8cPDo6cxqHYcYaDl7
+oNTtjkf757pOWkT1WI8JeDbG4+goT00IDUtcC/c00hYNhS4JSjEpXzuLWFwVs3I
K0aHh8zmeH9p5q+444o+J1Feg/ee7+oQmHnbMWylrruGanPAiGwFdxHWTa5fhk/b
UUiaatRpMHFE5skoM1Ee2WC30mW9PugPXkP6b0hP+ZJcR/Pnf6agmVi4vqMFzT46
Zsx7aPKdGCujnRhdDWWuvqb/9/XkoqyC2QHP0Ri0PBQAI4KAn0hqkUPu7cRc3hik
CWamgz+oU0s0M4zJnD9hG7n100nnqWdoiwHU18vbXqw6srX7bPqtVK4ezC06r6c4
aOSZpaUnyPEl1oxPMVDYUpxT57naFkzlUfKYjcwftO52WG4V8oYWPUnShggVov1k
yT2HlFP3pAw2MPU49TjqHDrbsCv0YNiGvYn34BOcjzEQrosNIYAYJPZ81LlF/Xyc
tSEXsiORh+MdcbTWNfkjhN4xRtI/F5xgESeywdeR6TPbNB6RQE9/MiRm6PwEpUny
NQat8j1aQzOIY30WI3b6p5Nlbchqo79hojCxafmO59f1PdpmLSOXHDrmfpFRDeLf
Nzpqvt8xyjZ3bzFkr9CYY6BpeSANBwbIR+Pg8xR/USpNKB8Qi2XLyidEMw9xmLmv
RhIzmcXww9xEIK99Q0EgMFDRlONcvvcvNICdqkgO0XiNAwCXHEGCXwho0YOlGxF6
YZf3CCvMNkeynS9dK5WE/c0KdyTY+nKuzRc0J41QgvLwQ37zw+nkRtIzLRe2qaS8
DkWoART08fMxr5atPuhtz2R47U9V4lAGFFvhjiVSnLXfFQNf11Njkr6qIoj16LA+
HT6tk8PZecyVKR2ve0X1emYNG5WqASieIjTB9M4k1cvS1MIneb1dR21BAHqi68vy
SACr8Tb1pt0niduMAImw3QDY2fju3lOzpEKh0xArRXD4ueAZPo2HCur5wNaWflPD
z4ZGd4XGmrALcvxbVJhZFzHWItJUkAFetAGohCrvVfOS7G+pnkHVX7U46GNCqmCj
b3JUJ1p8H5U7HQqQMAvZc0GmO21Blq3kHdb0OreqcW4kK0GsQhz1vJY+tgEhi5GC
B38qlmU+2mXxziscOYwfq6mNrDS0kHMXrQmKtmt7gZ5iIX3MUMmraYThkqZj5WBR
fCpRuOow5QfSNYKfK8NVsm0GjuM5hYeTtI3Ol8M8PkHsdbKDjOrktbAb75WaQzys
IcZJLmLEs65PZbWDYIzPB28FfEBAbrof+E8arV9s7J/oHR7kqv0wsp+IHyGcZYbs
B0K7gxD5guARSTrQEIYS7yTrLRi6qH8mt4KVnissq7RmrN8IS6lo5mcXWDaDgCX1
724DsmMwdfglM/D50hgoaH0jN1oM0+zHXoH/iA38cwqhIdIab4Gu8sghk3gQh87S
q4dutLBmmmAgqym7CHaouI/9qZ5Xi+DBNzB0JXH+swoPcLBniGRcO5n0MaUAh24z
PqFWlVszf8ppJKjI/Hqh0e8TtEbBi6HwBa2k7VFEyv8roJ1sgKM8h0g0dvBDG6Mp
PeJEzRWmdr9yfFUMHeopNmQSkQ2K62wUgAXJFIl7hReCJoL6XABOwstFWb2/ycnD
6/5mql0oSb/+79r3K8VrQatVSLgJgbyLy5c8pJFv9dsr+8yHll1tKrz8Z+4sYz8w
BZMXrCmq3B5r6fxkDnSRjq7bgqCkvybcsZr2gy6UeGBqV0XTXYj3QOhy8m5btZpi
1Dgz5SmdxxUeYpxNu7Du6eTk9jMj5EUBcaRv/kphSupjRxVTOP6yoGs6e3BRgKRR
TPe7vllMxd2M366Awf4/uVe5s2jfWxG1+zduzC6rg0u4qT67j1cbhptzhcAOIHd/
Wjk+yO2DPKLUNBab8gdFRrQ+S88TvxKOVkECyy/OF+js3y6EZLrnyCYc45C/e2dM
nBlmKg8gLSwA8VovxKi/qmp+RE7TqXZ3wPVEbsm4zPEm4W6px/FXao+BShAKwaGU
LWEjHMp8kvRHbBZerIXhGG3IkrFE7WWmaGgLqlhjxs99K+l8L1zSFpeSyf/7Qjsw
lkXx4+bkjqH7JcQ04qnvYYnIbBDHggVOfJRv1cSoZ9Lbz8psyqD9z9VvZgrxa03s
ZlaWuN+aOeZc5SE3Lv7KxH0LPrK95Kv69qPnLm+DH4SbFxGU8+KumbiQ6B0ruZgZ
cE2SzVpd00fh4lbl/W21/97ZwIz3vqBxYfgHtpQlppFTJVQNVQqub4exYuhP3ckM
wXwgcQKzoE7k7jkGFFBTsFwwxOnNEbh4R3mOkXAHnmHRkBWUid/PzxUehlufVZZ8
iR6tpvRJyfTPFNzAbi8jlvLg+nC4PACWkW1hbDSoeNarysxknOCcRPl6wsaT0gvu
i21/9o1qyOjxICPHrOGDB4oTifEIH7A6OvF8B70cSBLampSy9p2vl0QUnYM72duC
eXEJZPPzhHoPVncuWMQhiTeSI91zoIx4vB5Bp9QqesBCAS2t6e8PrJB46Pfp69Px
ALEY6tv6Q3yo0IHWdL4P4bHnHRCJldVlQZyxWf1IB062Q6kTeFqqfDShUpkcFDnH
qMPvleYRtcXniPhGp6mhk1pukW+yjpTZ+66IDUOSjzHmOcMf7r5FA6SC3f6pn0eH
uvSNrkCn/YSBGCk0oNeOqpWapu+/M2fRZyN9TSwf+0p0qzC668GBGYIi+dn1M11d
lYlLxOF6uS1/jY3a3XswwlK5kTP5VWVDI7OLvbLjmUWJu3mSii0bVonHPno3S5ZQ
uFHcggQS8t091NRMu8Egc+qOzDtnv1fY3EooLGk3p+zfairH+wqoha7v0DeapO+Z
8XUCqO7Y8jcnDQJCrtg9WOiYJBkFBglm84TQIEgHcAgS2+cmSmplfhlcXzBuWf8j
sW2OhJrKfulPAwWAjWWSSWfXRnF6h91LcPe4IzY+CwwTeFIuBv+KHPQLEz4a23aw
xvsFU6kMFr3ZCjSxUsM2uV0YMj8Q+o4M31li/ES2sYqc2vFokBCA5ZeY2otKohMd
bB4h5XTMImhxI+pUCWDjf3tHSO45lu9Kg7RPsEW/ZZs29ow7Sac6jOiFp6JOypoK
VvcXkLH9x75Wkzv7gXBckhurZGn6ZsUXSptxAorokS9Ct9qU+L0Umz2hxmpXmsY9
+x/Q1u3pQjBbkaOtcPYpH0GWsMEpeeOLO0jmiNZdEkhCbgjX9JFIELTvgfxPqLCp
qkDmojIq+VTubY9jOkk9RfIre3VidtgsocPBbYjP0J2eilUBBtHMi0SnjVewEl73
iCdGAlhN+d49RzA9WFPQ1g2h4Al89DByor2IUqSj/2Bf4QotrdHFtc/KXP8w3fZ8
J0wA9RmJrZO+Iad4/a2RWC0a7Gc2UHl3CXRBG5xvglr6m2fP0HtqLbGiDxo381ZN
wqlapzeASg33rz9+rDXP88AmNqE3DXUkytVrj4NbS3BD4OSBb6pavTvBpoOy1o+E
sL0zI5JzmHkc5NZ5sG6AUFQ/rN09yiLVy/POxZq9vDGE9u/kj2dhj73O3qYhuJlH
BR5n5SxBjFpy4cuQFksTzEo8auaAjPhObTfSg7+IMcLfi8EQOioH/pjhIk+bRWlM
DGxzZmCRcCpbjuSwUzHebMna6Ewdcl5Onb0cSj4ok/i9lehtS+GE3KFxl8F1rfKT
d6w46InJybimIaZBnmTwvPJ61BkBZNDwH4+CCouJ4BWrkOe+4371xOWhkpGfIcTH
Fn272nW/boe17LeqvlNZoIHX0f3ir/DqXYjiCF8b9ujYU/ZZJwS7EOJv4jmlzEqk
0o6IiIOEfsTHLrhqcK4EiHOy5KIb3Coeznb9oIMFGYDxViGUba+Wdfht4QtXYNGK
A45UXh8qQ9q6bnjl7DxSOxxoFIR9RO+oKPaF081X+RtbzRS9z/VBy9nlNFnmAYrt
zpru/nDZTWngHgA4h4MuSxoMRMpFXT15MPAcSidL5kkr5deMX42xjhZIKqEN8EOg
ha6Zv10FiRSvz073uPuUa4v9AARZP5ZYDWgKrJxpcC34I8LbK9akcS1oXmepqKPD
BIPpsHZxmePxIqZE51OZRKPFciEYYqVmLFE8O+k78+s7tGCbgTfcCxak5Fy2fIJl
MDjRafY/tEhqyWX9HkuDC8vrcvIulxqWTiLLG7PAP/Qo600j9SQEiA8yB9niMQ0O
WxF1r1DNTok00NjoKJ/GMOiJABQHUMIDFRioQ97ximaiOoNOXmmZoOcWr2EpC98m
Y3BkJwNg9J/2EFuvo/tUNaX8tPKH0L37Zii5Vl2eEy05TnyevZodKRbn7PoJoX8k
Zh/5+zzK8m834jR1etDyw6R/iXjq0R0JQj3N8lh+t28mwWwXh+P5HGVjN1TjTI0R
Y27WV2n0V907Jnic+UjdU6lZruy82H2VhmvkPQ4lr3lCgIWXCGaA4ns/Jm1lGwaY
R7zY2fGSbKjQ3QgD1EtbTCo3r3YPk5pT6Qb0Jjl/6EcE9yTfs4iwIiryAxef7HTO
Wvjl0NK7I2lZqLvciDfrl96PnBU9Uxoe5qj4E7kdI5j9PfIN0VlLg7cCYAThzlwI
3L09Sz/oAdxFflde9CaDm84Wc2IHi70LI6mjlkkan8g2AVbgDiV69YFkMn+YYD6R
sVBnASrUmIDy0pir2um5InNAj2U2NuSqCdlUfn6SBu2S6vE7p1eLCzLBBawKf/IF
+d+DxDSXOKETHnXf56qHxBTy1GIjjG97BT7pRmBAjL9mGTOBsTbepOggkGHPQW2t
+Ln1m4RntWYoaRrBqniHLkJNuOgIWm0eF+tC8kG3I4iy/PYDv1rnBjB6RinuJZjl
czzNAQ8I4mlraF+Wle8xXwk1runMBkTZKbn2a1RvISxgOd6Hur+V0UDl3RsFlDGd
RsCyV2lzLUIK/J1M9cNhG3EcozSSr04RRc6e6v3AIn3fT1szMr0MqTzmLmT5OrcC
GklPd/09NaZPHT7VNd6VIs4U0zw5rr2A2ZKvneWaLRE3La6LMVpRXtaSZ3gL/4ZJ
gfm88rfAukK7FJiMaDk6A+EELvlO4uM1ptpBUMsV2FTj3CVSVsaK+EdJ+q+GcPK5
GQMgeA9GmEgLLTwNBQw2tzq3kjOheFM3KQsuPg4zGY+8N3QDmEU0B/kwjI4ja5KT
XunsxqMgnvb23D/77sdySlE9367lKi6yZbsispIT1oUKG8sZeTeUIeVPDLNLkZ17
vcUy6q4NaLl4J47KfguyVN0eBw4XBXHoL9aWegJPS8yS2XKlYt2blL4zSLXYW36u
SX9YUI8m2yayNMuf0KSUu1Rpi15c7inmH7y3zbD4MU9BX2u3vic53npp+2eBMb9J
96zM860thFmZ8NDQ7mDbSGNLzvDcJ21s1DfLmG/pbiWjWCHolx0YVcqfiww+5tqn
fscGaWv377q/XIt9b25Vm2iDO2UoJm1wm8MOK25jfJt8ALhCIkl+vAEpFhWXOJyY
VCEf7xfNSVgkBjfY/loBJXA+WOlkdxLmsP369zp5/SGoU7n1NBjG7eBpqKjhgtsr
dvuhTStKqU/QskW6nh9u2NPSzwrtRo4JJV1OIsjR4X3bFhkmLFibu1Fp2viQiCMY
oK9ciDZAa4AT+ROcdHMbkHCXw5mKJ9Q/pMo/uUBK0/hZbal8lNJ1frrqJNfoSwWV
udASxJL/yWP4QPVG+rNvDhXl3HH53bUXQNIHSJ6CXCiYJvhF/EuybwivF3oKF3Op
/XFSXynZCc4j5RCDctCk9NKEpnOh4Fq6QHHM9dKdkzDhPmcKOJMLOPezPOBLN9VL
S9Mg5UeWOrvCYm5fETUz06t4EN0pHOxhKuLc/bjVMkpw0zEUUjmWJgT/wnN9HSB1
lpfhjEWLRANNJEA2opOffGPzRt5GTmlw/4LRrradOviKYJsE7J7l1oiBr2wkrjcJ
2cv9HWeps5CfO97L0dYraQ0sQ8JtadXuicbusjvN60rJfknaw7IJgSvJjaVBew6N
QlLPJkphd0MhVOg2+v7LE+iXLIQ7U5hkuu9abraLpBMmrQJdwyU1fXlW1LHb2xZ0
ifRVZUZkGBN+E3+AKCeUu+JiM92GfqfSxsXDkaf9Lru2MZ7GEshj+CTk0aEZg5e/
pBl3Z5LAlKh7tvqTPB6oIR20EUjJboH7KCDxk+ue2HugsWhC16Z4aywQ7in439z8
6OLDnlsFi0rfr1klDGd+UXzjEo2+NQgbdGTesK/hs8b1nL9K9poBF9cS6mpnAYeX
DWhzMixDdgNO1JlJUzCD5Sr5nxV5DPpy6SS1osQvRv4x5b43CUN0fNvZ6pYAYjMa
Wd6iqSKYgF/ZUPeMfFKFTAJIAy/a6sU1zyMb8s4hiQcFhOHkcnl859X022kQsC+B
9yYEcdgruOtybLAyl4rt9J+2HzwmK0WieTJcnxElSNVhEuGxerl4fJUKzkGkKli9
anFGjRaOfW1nf5KkKWcl+novNL1SOj1li0mbL16UN+t99GWYYN/gFr9VJzKn7wdP
ie2noTdelxoGm5+ipG/mzJwZxGR74dIZszLALTBXV1UWbrDoVH4B1b4EFbtE5mSR
h3upX4LfvbPf8qLRe+5yaUlQHFn024rXCrnGFOEGX7I2+ZElN8n/IpR8cyktl39u
cg1KxBxh+z6DF0jkn49fxJbf77UcDmJjPF8vstPSzKXfu9o+EITe3EsR7cqLgGfi
wKdJvPxDXMOWlj3EKVPZ5Eto091e7x7pAnz2Gnj3arnTsLsVrwrEnT5TseCIvdGg
Xq21o0e8VVDE/cEJc9pCmN4CBIXSaOWRqeiKEvkO3nrSjZP3W/E4RGsQe5C8U0ar
hMDrpt+SHcKVC8H1+jip7hW/R0ksMUhCNe+b8Ig2/EOmkYV+gfoQUYZ2mSjlbsna
AOUbJqcS0MpxkDrTwLdwsfQMT0R+z8mx7GJd938nzpKB2hSL5e/SuV1jVVg1ZOtt
xtar6ziUfywB0nBi/ekPMFEKa1aU2LXjzSlnQeQxIGzX5eO1Gfzlu57lqywqRRDi
2KlEmQgjuFPjIo064XBiJR+bj4Qm9ebYK3GFw716lluZd/6burLl+MwmbbHzdv3X
qk/W0l5cngcfbidTD6HFqtJNOXb/6JHJboAYzonQiWTwe7WJ2vpwPnovirDMa+O6
jL6E3zNoEYfeDQeFK/n8o2ajOrty/QSH8qk7/YaU/kDgtzDPMnxVE1R4vgW41JxY
r3sR/bnkweLXR2IkF6uz6fzw2FH5qVkyDrf2fgCjAWYq3DZ08IGjUWgp5WAUhdWM
p/oD4XQeBDbjds4A0DKiq9paXIjQG9gq0qT3WgOS6f/Kicxqwv48ivks2QzLIMB1
RzYxDJ+nFalhllOo3V6PyX2z5V7VXjUpljeaLjxmkcaIfDYsZcg4jhsLWeTNN1hc
yAzvc8i2JhPqG7Hci4mac5dS+SrdLbDTQ2tYrSV2BHMAX5cJu1hwNqZGQDf7o5iH
STp1ttnOs0cLXoFcNCIiVFf4Rs3uk+YsHT+azVStN4oWYahW74r0E72c/MyPhjUL
iZAH+JUmWWTxpCrK6UJx+VYX4ilutPOainSntrrCzOkSZhBaRJVYHWtGv8Iua9pl
Vx+28WZOlhXYPq1bzLTPHzMCkYBunw82Ws+FJz4Ef4jRKcwkyCWqSpTGpNZk2nkI
QQn13PhpYUtynwJHHXKfciOXK9sRTrIhmy1+NXzzuzXpsZUhb/sTC8wYtrSWn4Dh
7c8aMi6GE6MlQCCr6dMtu4G+3oS4zM6UZ01YN8jR8l+r/Bl/P1BxRoU3Be1AOp3W
FNYSeCVoUfao9ZxduD14tH4NebIkf4nC00qV1Z+sl8KoVNQK6dnWdVGl3n9euqH3
Nf0WgAZcnpU61CVv3pRYqnLRSS3dA1ueHRSeYTL8aIVtpAf8SNDTFL2/Gm6ekaDY
8rCuWj7bALlhjDdZwSSqM375ag8YqHSmXAL8EoVGzbdudix+2LCLfe3t9WYASt1r
LJJMqzjloW3AvjjbjRr7cpoS9oLBTpt5gOJ2yYD6xjJ6sb6X/Hb0r1MmFjJXmqwB
cur2awLZMdnw2bKzp8w+MaC3iCKdcansH9JYOuxj4Zp3aM+reE7YXvbEjOsPpjBg
yWjKP18j/zQqMgnqVIQRLfVrNoLemT81IBI+I2nNMU+Yzj0j5Qg6IlsW0s5iZx8U
eTuzzNPlNYkWYhkulhjOly2RFZpFDK8gWw5B/SVqz0DtYbRP0WMg7vBxPlSwEaBW
YZpHOKwjWLv5qr47JuF/lkY7ljHFh9TffvdNgulby/fr+whpwNgzGQZgi1AhQrdM
r5t3bkVeAGsXdxPUhM79hyOWTPiECx5InPI0J0yGnFe5pOD7mgCnqdcQBEG2mQ5c
VZ7k5jIkKbyja0w/6dK04qb1RlTwrEG2FXlEyAdwdT6sW/8QEuepeT0iUo7xtfS4
8L6A+Zy8l8clDF/evT66Li/QvDgu4VrSH3zrPTiTabdgJaH1HMvuJ1m4tjsNSKqR
O/IbeaXuiG8BcB2UWPI4CVegQ7R1Z8Wl3RVctOv6R4ygZ0blhB5NEI5n1yfOCpUx
GPKfyJs1vH2C+5U9OPvSwDedO4/0KS7SfkCS4KiVFIdkce1lg1SMni8gnK00HX5h
OUdx/hZthEtfkkHijU9OmRJ39KKy70R9xxuVRCwMdlfttpXXgZoju0vm60biZUFs
rYeekayX5Ra4PBjh0D1mPZlh3UJ/W2M8Gpra7EboqydGogFOWqZBdamrlorYd/VP
1uWVmXCaxGzJ1ITDZg9WIML/u8NaFPAUnc5ovNWWg9Rpovaq9w34cvCoyBMeMgpd
XIh+HId2R3PD+Ob3bo+6Qa0AKojyiHoM2kqsC3GA6L50jjYgGJXzpPq39b9VNMGY
9yct6KVFqOagaXRwhSdvYC8KzlPN8nIrTJ0DE2jFBFvKPgMC0TFAZAQBLIkKtmVq
fd+VcMNqvH5N8Vf7kyUWODtgjiUVT+GFyiHOmlc41PsanDDh/Q9+9KpYLNufaKeF
QjHkatu+JUqLlSCwpgtlGspxSCwXv6yLPmAh4fTCegYZw0h65J5z7wwwnpBVKbDc
sVF//A8E6QNoja6ugpr/2vbzRFAjvRaYmlWW6oCdy2C3cm2ORhzfKLT/tZnedd84
Qr1zWOszpSZMjaWBqHxlQX8wX1sd1hOTyCIa8+fzrxtnObcleK0MuN1tZCVNfyat
Nt09xIhP+4pnk5jM6I3w+SkfsYIauhoh1SiSFJx/g8XB758ZO7kklKPCH1LPxksi
zXWIwqYEW5EMcOCUrwvT7ZOWj0pCwCDMhPxfjjH22vZca1zrqwaLmY1pHNx1yOn+
upsWjnWCrSdlj8niVJJ+2XbDJyBmNZ+xTEt9SbYkadyptq21+KVbE0jeTRyT15wa
zUlQiaomaKpUWvjPQgUOKN/TWSyFnRKuN8n4vm2xrQXkJd6idD5ote25dM6aoW44
lKJfJe+iaVRGJscTpELZdqxQq/9+r8Cu7zJnq6KpyBHpZ8IfYxuZMedpqY4b2/Vy
tATMA1N7xjOgaNb6vOGVcXtgJFCMBeX9r8b1zUhS0nksEBlhcLxjaxKoiQzW8UDw
A8cosnPdwQWs/Cy2Awl/TVFgxX+vQ6AyKEpkwZqcyL5WhW+gy7QwS3dYFNZMs1CV
5PDzE6PKoPODTDERht/9rnyq1+/XrFQc2NZcxmSAbdzTuBytph7tEPaCUywKDF4r
Ofka3syIlJZfr75PXYtYrA4Yw+MCJkbiOCeDoH1MlQmgV45Bycl/T4Vh5b9C3c4m
MQhLGguHGVsPhwlBScFYhSddtFUIKUOXeN9R6Ha/IQ8rjgJMjNVoZ+hlNYbP+Xgq
/wI22MDsg4K21ppFa/oRbhARlZZx8EBzqFiJMXbkpLUw2al2fsylH1OpxgZ6SFF0
990Xman2LKv6GOWskWx6XfoxBMKsoWxp6XuPqE69SmXqxTWPKf9Sytwd6bXCbvTH
oFOjp2L6cbZGeQ4rHk2dg0c2hcam8wruN9h+1LbR+kuSWXiHDnE6gWTHOtarDtCS
y+tZemz33/A7q4qVOHaT12ClUUbsDdMMBzHNPS07XMV4Pt99Udo32l2+10u4xu+d
bujko7fH/TDTTIYyIO6qip0ZyLioqQr2cZfZZqd456pRmWSI3jttzqoHNw6OfCwJ
/QaaCwLXIJnVsOW6GvQbWbaJQCP5y+qJVrCVSMjPF31axhu9KvTSuVAK/YrbV5qT
+lc56n4YwSZwZF64zv8KwckdIpxWfK5GF0XapcfqcAl7mePaFT/OcmT7o10R2tlk
rcG7fS+ze7sXf2UAxz4Ryu9RGESo9008MaqJQF+tsRLVQNcm3Fmxei1x36TPWmmc
TFf2m8+nup7hwkZbCYtESfAzloJvvvN0MjGm+7xPumFscPvarhN1u+43vV7ymSdc
lzskE/LyotA9kCtexvDY6CtGsqnHb9Nw9jr9pA3WhhDvmH9PX7LA4crt5No+3VHq
jzEI86isJPSlQnF6qbFuRi80XLD0g8NVsXOY0tLQcKcAKUXjTNvb0+vzg+nURcj7
LHoz+yzWB+GalHkiM3nyOj9SuSu1bA9ahZ9sHgolYfe8mHd8OhO1wCMGli1Gewj5
VIsdy+JlE+uM6UoRP+wDlI/+CdUzOf1FD1hba0RLRVMJsTvEcsA01d7K/2tuttKx
9qB8jRu6ZmP/kp+A+qvNKyf7b5XBtItEFYCbf5cu3H1cbJmXlhakvGcmlKlSHqNs
0p2IYHHUc7VTtGFvBT1MzA9ZXyW8HlLkUI+Uq2AyT4tzUAbnxQUcddlOtlXem/Sa
NxajiIa+CuXFe+qIcSuL92wOE5fK3yR1ndJ/rSeKNL6+2zA8wFJxrhriiLLgg4Tu
3LmTWNdhSpCq4FWvsY2w9+Tuja9tU1lvC9/Bvm5bVKGWmdUXjYF98H5mbAwSx93R
9KG70OaZYJfJYk0B5W9lI/D52uoavjg/JkbTnbNEgXxDNz/GqVOB6/8ETN+401oK
2y/rbr54aj2oYwnJXzNjRmnqgijgqdOHcLDa7NdvSUxdoNI/GRUAJjNh0aw8LGNF
h1zjEv/S1jZmynEKYXplZOzBpALUvZAZOBBQ8XXq6TB6XuEfCXWn8Z2fy5aBOBsy
dcF+/ulgXJXWAc1JkmS6pr+OO/A1qFFOHG9yhQR23mKDesqz2zvLJIkzX8QRuZkW
ZeAyNz0DOpHPIe1R/DNlF1MgBE7FA4IuLiUWAO8xAy22kyD140k/2Tfz29lBOJAI
JHUbocb946n8oC2FtRA/gj+yL13VdV4qfz9nZxrXwkPT7FhuY7PhUWc/hQ81WMSf
j75N5p0+c0zYB6/i220BHqYkoHXCiXGybNDYhE6YnCzvgMToSdPTgY/ZHql27Nj2
okCXyngyc1fq/NtixYcrCb7ymKRsjT9u2ilOAHpc6NChCxLw1/gKVYbPv4ObJcfL
Q9r63tvI9SL0AuLYWwyn+uXbkPWRimT8NHV0IY6MF+Xb4yToBn7mfEm/7Yp/FnCK
zsteN5nZI+VISDqWR5lRbfChm7WRZZs0/KIuu8CBYgrZv3ZMhehPueZXECtY+74c
nwBRJcUa3GTOwdcznjk392bTtjmVISTAEJ75W1mQnkLL6sfpCg/Bp+5q/D4uzhq0
nzkbNATZpZDvpLXKU85DuorU6k/QHfUTzVtgmiXBGWVXvcMhs/LbFmFfleTO8gzM
WWbJFC/1oChNdkdMq20WEZgtRO1Wp4Vdl8GWi+35LbqcMDLrI9e1rxzdzNzZeeiI
ZjAN4VmWEzM2huZmAxZeFWgLhY35QOkwCuEBhUNe1fnyMFKGrwwNWYALfbTELX5s
96pEV7GxOTge6KanlbXE5NQr2DzgIoLfyttCDEhWc9BaOlIxJQGhZegOVEIaYQ/z
6vYENCbV43uGvpqImguUDNtZs3Rc2L1vZ8vPuM1271k4jD5ecw15ZmsaerMHsDyy
njPzGWiv9nld7/6WtjrPOSEKHcAabne96qWfYQHiEhFcdnIlYbWmu6PadqBYChN1
WhKSUTEr6EVdjTAUEXBb1hNG/sjORIbWV9rBm8rSQ8PQiPt8ku8i2psGW45HRO9T
RxD4grrAES6YNVUqMWXHiJfFfHF1c61KhhDRM4Wyu+SyeOFbKKUbfZYr3Z255F8U
8p7Vz5m37Wy3KwjoG1I2OFNk36bu/VNZ+7MEXXb2/+6cJqWh4kNsaBlKVuvEjSX3
avEpT3YxXt/IjJHRkMgKeaUv76QGIEqL7I4Bb23rYvXwCATsGGR2zMwOGiPhS7rf
d99ZCLB5hcxU7tZvyb+LYv+NNjtzkUCTxlXOrzBtpz26b06x5/invNCIE+s4HDme
+gLfDXPqT4Fx0xYscHRsnImRVp8ZIcJIp7Wnyh8TbFiUEwfytpuN/mWxFBsI4IyI
hKZT38Jl8M+myx5DMxF7AGoc5FpuQmQCtYG8lbtGh3XDjTjEAJiQZC6LkOWPfr0Z
PvoAeNnBM0FIaPNOHfgYFmxLDp8wkD/S8GYgRj2I/TMm6pb4GmEeZKRRRVKk0FxE
Xc7FTR9XJN/MEeINkDi/xZBmKnRw7ls1A6SrYCAnRiVXkIk+9N5C8BjgLXx0gp86
jtANsw08TkCBBq0ek30fnioPq1UuKOiwU1B11XsRk5zRROsNIx/G9eYJV+GPQMHT
k2PSPwvRWINXwvHDoLuZH7ZLzOBHXftsAxiqxheY61/Vhxb/tCOBAQctfEq/WELG
Mk2WS69IBvaHidJB4ewGOm8J/iAKEwUD6ukkb7oRlrBRjx8SsZ7zOixhUPYKrqMq
PAAis/TyeL0rQb1VDPBGABl7kKwzey0UsXORqbSQoDCVY8oP2HhUlOZ7Hmr7Yaz7
tjJTuTGjB+0u7G0zed4I/wqtbE+X6enO60lDGoiP5pFCGGpXnKKr+tb0YBlltPCr
uzp4UmWsFZ49z1ifVj7gSP5aEWkOgkpQYT7ipSPnVFjlmIa6wX8XEOZzOb6muK1z
YdKtriDveF0sr7P+R1LH4U5W0TMYiwhVmw3NC8elUxnkvayl2/3IKfnzCn54QFHf
MeD1ROBkbojNnLYU+eATXKOHeWW+/1VfdsbKUCApFMyYNjmDhyuW1ZqeMHVBArK9
N+PtkufUNPFcZJVmuQPuLnIas88iOsouIqP/1FZYQT96bKzUbfGzUvPAmeaOydKS
yldxcLBxZ26z0Bn12x1avvmb8hE9cSDGz9N9La9E2Nax8qhODyYXEYoSxkIWU5wa
n2rhoi05aUkvubAS8zRQMrvO1yMym3wYXXOzCwb2gIKFPnq/ZglwsS+uC+Cp7vk0
FGnAgDr3q9qSfOXEm/FF679EDZwdNitumOpDom1HAa0ojfgcF9+D0PFV2Fr6JRAY
Bd/X+A7OLzhtPfMfprIE5EUw3kY/fmzGomaidCe5Jzk9+V4i9vU+K37387tSwcZs
gUmzK6GosM3v4IbGICaE3KAebxKVdJsNjmPfFRqSHDXnjor1JnyZ9SI9EUgTu7da
x5crYFOYkFrJaYZhgtuKhPLYUm3SkfzqwDzL3jOq/gRg03qfjSadGri32QLdzb7U
r5fMWUBsZbQNb2ODKzeJLVDK8qIvtxUl/C4812yFcsh/Ven9NgMj2uvRo1pjXh4V
kwgdmdTBjEMCEew9PbSDDza7Ntuej6KPIFYCvjJ7bnQXdEyir9YXeEDtGu0OSZx2
Ijc4Xeg4baBZ07uFIYqPQ6u4o1/7W5K6djINza9TGDLglbN+/NETA3TaUH4eu991
3YPkeeWjycsghbZ9LqVvvpwjmKoQ0SbKDTzekKvbnm6kbrynwK4FoE0eWZSdJ3Hl
Xy2aFafInc3PEIQUyjsGtgfNdxyqgNgdMgHR8iGcPDG0BmqllibTDmOfhckkK5lU
YCkb3JaJS0aiH2BOZQ5pa7wjZ4bew8vVNpsUeSa5WcRRMi3J8JGEMnr5b1oJKgez
LQ8Pys5U9UGDb/czHTlRvn24siWYhV4akv6ZL4Lcrh8En1qYz28lW2Nyl+14CicO
IghjxdzsB9E7gCPNzdjSvJTd7UsmoO5R9IMj+rFzUGz1KlPNo8tKnZlRuJG0K5eE
kb0Jt0JVbpaSYtMGjwHAOtLOIntSkfwMiR5PncpZImVsQupoT2Lx+jXVebY51WpU
JfJoKc8Nd8x5s9U5HDP5Qr4gMcdoPNRUbX9+XMDYjlda3gfoPKyg96nnyEObumLC
9Qt3rdkgsKrjxBZERXbw/e5XLh7YFYV4gJ42AR9lryOSrwpgN8iIv4SgGxxRxYJV
Zra3YXWvrRrkEShd5EmDChxG6gX0bBiUB9afN7oAa48RD+xZmEygfVMMwsgtOivM
WxFLa8IGCQY9A7W/HZScSf+PTA+2zyH7IMS2fe154j7dB63RqWfabUfGe4/Ruv4c
rQvpoxpgMYYTbqNlScQLABgtnIcyxOu2xKSVkvTb0qOwzQiZpBq8+CNjXPiWBE8+
vP4rmuXNNNSet8HFWftGaY5QdCT3IobePBhwXKhGFvOfzA68Nq7j6pb0oeXaYENk
NfnIvWcwTMmM5fxdTyhsgDgBW9rznSPh6Bpf0JhGBEMIsrYn+cVzMfJGewHFf+uZ
PaO5Kna/VXEJ85YW8OOl7KQY+cpLv8bgVSYIaD5IwjLC6/IFgrqJIF4rBtoXsWNW
WTFKeJWVeSiLcviqtrS6mu8sNGW2KJMzfPcDxHqfEPj/NlzP1JiC6pg+3T4sdToW
UCMM1LZfex+PKbpSb8ka2rsjkDYt6LYNQasPoIo62rTcdR1AyIyiYqULfe1r7rzh
LicM5c4q9l0r+zDsxrI4LfVVUa4qfzOslkg2UJXucNU+pSZJCp8srMDtpDZWGdwS
tOVzUdTWE/CnLF7NyX3DDNF1meE/KhCoy5UNd6baAmQ6ZXXByLQPBz0LE2irxC6W
jIy2A4VgtJ926j9Ht8NZ9heUg1FWE3c6Ae8hunGvApQeWpLwLkK9M7dkXXF3f3CY
KzMgu1D+qKOO0ohCFVlLJqa/PqXOfzhNtaic7yUVZ0sloFRNL46eBLragQjcI2Kg
7A9N2TUxTDnY7NjtDqagbK68Ht5nhl9SAyoby8cSMax/FEMIumIUHExdoBiopaDn
23dD6YRlry8bOIiuzP+AN6XzS+mjRLZrrW+4Kaq1L8vI5qyZsBSxk1nQ0QNuCuZd
HgLXpE9xaVtqZlLSImB9jUR0nRb5u7vbiAysnZ/ELl4zUb2Ifnw7vqlbKNFQ0GpC
T9NhhmC+jW4aDWFpAwbqYHhTJ+bnmmUkIFMEf49XiK/4oFqaSrTxzQevgx5yay21
sV6Zjc5Jdsq5apwiWS7jzbTcUqJBeEqN+dUqscj1FZ86mA7iPOPVzdRuP2iG7yfp
teSVQgCxZ/2YtFsXTmaqZM/7LrN1G2x5dfUMCyUGfzAW0YFHKLTi7h1m95V/Ajku
wHtyVSJ9eVMD39gQvdyobSlOUbNQnpn0OE0qxN7q2f9TMztVosacxdhWF6h2sF29
MCSdNx+HmOttNbXqjd88s6umB0Oz82jwCAN4CoXDO/FtMtkI9//HS2enwtm3SlH7
BSkC324eFjxjVGgpdjqsXhIM8d7iylfS0dI9yJt19jJeqBpCF1eIlguW4Sp830LH
r3U3OwLmrChZoOswuxdbxf8QBBXgSDY2+f/D31zp/MiUWKsnE4x6oiIHaGbZEjo4
96VNHVkmJYetAtO/omKcQ+aa0Kc0dI6xsvw4ZFMZ9J1/CgMJtFEunoBec2UhRGCp
qt7sqrkmOqbJ9f5NI18qwG9Mlny17hw/F9VVdoUjGQAQI+pZBaEG+lj7KMQotmaG
xVKDyrnjFMbUFAKaMgHmeHq93d/7yHYoVnsIO/9j9ZETgf8t0SB7hHAc2YfZC8Ze
bfg+zWYZfFeGPxXixXnqeTqOsa3YYx00k8hO2TTazdWbcY3deakiNpTJCFZwq9Qd
WhvcYfxwqffCLlMFIlq3N2jdmYU0heRIEYi2d2jD0iBUzykQ8PEyTah8DLZ4AYkv
NxBHw0oQgm9/HEAKCvEaBJIVj1vhgRBT9RONQPzL0aq6Hqq3WI6j9HGRlzB5pigD
dYxkNP2tFk6x0KsE9zFZIW4KjwH6UTXw4/qEuAXHEbImE8Dsn8H0QAFk9ndjKQpE
JAo2n1ao64fuNDYlu4nvNCN8daUmOFXQ7zlUQAEK7VIOArtvOYUbuYI/fP52hywx
1828VA0nB40U+2IXtX7jLTqiYV7o4llmZA6HleTa+zCB6vaGdq6Um/Ac1C7bULrX
V9/dgF4qc2Um/x1qzrkbHhwkPWQhXZCVMktcOWFOvqBzntmSfEkGIy4y9EN1C2o2
t9oSm2uv+PymfU+2adI+Z77A9WB6GdnUKL1nY7IG9Tz5YB7gCCI+axlz9Y0igBm6
Ge1mV5PxTQ4eueFukSyq7N21och5vg/5LUlbVwHTRYOSmJ5b1IMp0jhEXGUvfTKQ
awgcx0z/el0AaF/B6KVSo2L5NG/ZWBoe/Hm0GjSVCW3p/L8OskZ0T3vWctI90Dk4
vs3T8fxdDbj/lbfIobO19TGGFJJc6620OWQwvBusz+1DrpLjMCFh+Jxtt8HjZQA1
jslBz1+QWbuq1yoTe4XEGf0T+rZ4cF8EHauaSRu2l/5emBXgMbOvy3Om3cedP4/G
6yIwEgAODReslBqFcImz1Cpb7JKynXfIBob9KCmO4McKk+MkspPCt9uuP0bYL6N9
2S78ryF81tWtQUsZevQJcL24EEFzpBnKwbRorAl7x6cuv49aNYGgDpT3QnJVvbWf
42iLF99YrClyHOmAoC5JLLuk1iY218K7ikDn87G4U8zAb8eyHVGwMf3PqUmxOcNI
x8myPL3Uebu3MwDtqQ0c6tnyn//wEF/7ZioSrhCNMvAbEtOap8SlZljCM8sWjTBr
Mh3ndjGtizO7+I3cwGwwo70C8EInQqevslBWhYCGpYCgvbc+zHj39zSEQj25o5ak
XrDUHSEqNhzn4duNdZ2cv+7J+T8ur09IZkVcoYS2uOU2Lr/TARkOwIJ+8JQsUaEJ
whQZRkT2o812wZVBzK9C0rw9+Qy8EJNKapahOckqB+xr2j118donZ3fjGSBTFpU2
+WNMAqowfNpQJeNp3zn7DfUATfXA6xHqo6d38DwHQXozNighhhE9HnWCAgCpkwYE
6pfp8NfLh6m8T6dHYsNk6nko/pG5woPuyNNOQyoznAbBYf3tW4z48+7/jKWI5f2e
9RP+bfIZ1Ny5qENkdlEDv53nFpI6+qMaVt4xZPAMVoY0mClcOeI3nefChTHQVipo
uchS4+Tk2sVUvWYoDOkY8suNc4KJDBZvQvOgUK1tFdBvuAV7TEp0/NWbCyy772ZE
yKnOOpX0jWop2cbkKs54lrZA5t4DE9u9QXSYgKgozWGFkdev5ABlm18YDfS9vcuu
RwwpVaTbeC0BsEF5PHtjccGjnooEh6WA/Y5+c1rLRQCnP2cmVXeS+yBB3L/aDR+z
DJSnxeHlSTedTGl03yvp/r25pitWRmu8gfmACcKiZTvEWJrFX8lpePkXRgjaviW7
bNDYrkQuSj93dQo3rCtBpxPVHDmUcfSR7VMYWkTF57EgQu1X240b4Vh1Xkyp6ccK
Np6bRrIrVUnr7JgwOZxp/iIFQTge5YKm7ZFTCrEr2fWdxIMlLMDUFn23BXnJzTBg
wUCQxY0NXBoIknGKG0a33XQBuL2s83qSZrLE9beh/c0scDHJGrqP+ELswc0k+JJU
EsirqnDfb10qwNmyus083R0pPaYn0ie9jH+2ni3SR1mP7GAWzyfClWPNiBc4AZxF
ZfO7dDQNTq+ZQd+q6l0poL4ZMayVggytG2D039At5Ydx54T6rqbvzDL0DQfSr3jq
cKxXKC+5GDLhs43BZGwP9Qk7gMYdBgGMuymfrbbUV7UIisSVQixyMCf0ybDI6Esk
JLqbeSDhGVm7JY5506ov/gYO1FbHpGqHKU1zQ1Rzn9VFbKmFZ9stejz1zaLs5vCW
h8l7huld3QITFRjxVUbZPu8/hG73dp0hLXoYVOPT3t/iS6iejkowFlKMFtCdKyaZ
UqXCV3nctF6aZEo0rIX0JdoEzatm/GMw0zUuLL54xrlyvJRGUOBzltLufWMlDFUw
id0wbIQK5rh5kO92WhQfkQ/iNQJ9SkXwKRlr4LzmSszqbBNmN0tWHKHHrRStpWRH
2S6QFwEfQyXYJK/BE7pbeE9oqLMgSqKuG31cTcQTzODVcuW4rRTI9U+3icGCHYPX
ALbLBuVw0MKUfZ0EirP4zP6xZwFSyajVn+azYUodaIMSGyLa2rHUwBa0W3SEXwBW
6ATBErFGjBBvMvHlTkU8kSbmdkJE4neO64OpIMk97xyGYH/5OFwgxtPc2av18sDl
5Z3KddQF+JC48SfxzhxoDpfWwvXxJpKWgNOB3DUSIm5Lv6lAhzq89DkSD4SQHMt6
nUtU7UfyHahLS2GSkdMYLU2yLS5ltq94stI3IeWXYXY+eyCOrv8vQnVEOfCXtk/G
S7hAGLQCiTzHcQu9yk3Tc/vd2gftnmfzCzF7sZGX2IhmETdEI0viRONQymFWd171
W0NHB3co4r/WELz9LC+FxCyW+fIdR3BhXPBR49bLdvQFJ2HZ7SpZ7jV54dzIDo35
1Uu9HjivhV3viQRG5NVZ3taZpWL0b0tZwCjQEKlL684zLcIy49RaLng7vgISum9p
Bus8toC0WXwt6tslglbBJGpG1m8iI3O7RyzA0Jfx4oiIOH/76ADBb4n0yVbOQgxd
8Ll6Rz1QtdcbBT9husIWSV4lbIu4UZIRBTVz+5jnyQkWrwUNPD+zXULOFvCobdgE
HYHGiegiMKZjPlu8p6CCt/cz83G42d6AyYRRTPre2wHCBRM5VC4uFSVvrBoBoP9w
WR/GP7MBKClLsepY/5sWmz0/17j9C/h9kzJioUkr6NJ0VgcXl38oml2NMbQVIbs5
nCP3FesOFeEvNcVNuVD/pWlgI+N26q3XKQZNEGVrL6TdjZn9n76R/MK/0zLaP12y
CS6Yi0lgyS4UfBRQn/BzyG6gmRgPUOrkT098RECq6xJkgLXBuQBIG1AUNXZlgl+C
2bcQYc1LNMVuyYpVl0pVsWY4A9J4GRk6GOhIpur3fHPm6rk+L2+Sa67cSc3uUvaV
aZKGkW/Vx+DAHBZeDNWOaekMGVVSfdGDxcOJJbMrPUWAmDMtkFP342OZ/62mhJeM
00TD76NIGSETY/6kTqduG9ZiJyxj/edG2jRqzc8x+i4rpbE9TjI4krgHekFdGtG4
c4IYHC8gfQB+2Ua6p9EhsU7m3/qvUNETTDRdnl7mt8oSNvRuu1UnJCmz4LaTLF0t
jUHyLQ+HjREgZBYiEOaypA2tsuryXe+8ZmsrYuMLmDB7e21HbWAkAqqjbWHgqN4O
t7pmApvHwOcrJAn7hAFG5rnHTkgJGFY3yReBEIaJYTsiG02Tq8GDsJNdu1Fs0kIj
MXmiMspMsgvKQVy2hWKJOZ+9xM26azcRNTDdymtkNzQL9g75dtVZsNyleFqanbUO
LznVmex2dMgK29+0Om4jicLva8NvuQ72I/kuxhLT1dQJCSHKpY+FFWH7SmjN6BVn
7gstccyEyzu4xj7LFbF6OxXJ0EfNyLsvVmRbCRT7Rid5xjjglyxApCCfe+Ny7euB
3DE+m83Kul2uJogo2CNyd0pin78a+L5tOlFVjWeHGYGH8LSHJUDT31qW4oe0zzp5
qKghzirQW/mlMBOdyJU+8jkxrGudZY+POnBoQbxoLA6wpAGuW4Tkubg5yEWftEQp
G294r6NcqPykVpfSc8N6XMUtychQ1ZmBmCPONn44oXxqo6Jm5s35sBPK8f8rgfaK
R1T8cmckfF2snW7JdREFM/54P770EIZC5HIXASxD8ZNEcLk4nPcfZGjBtnhfDFLY
BWj2jJKfSpacG62v5Qp59tY2Mmrkn/OuwKCbysqbTvnTayMaVEdBnNfzPZwurBmk
TW3ZU+4e2jlVUdP6atPX/sOAZsRkGa84zZJYzRDG05SaQSGfW49QM/dYIsXkoqir
+rEBzfkuOcs+3sfpSU8Bk4CMn3OWQ8D0H+F4tpLAYkAmM988wByAdSyPP/p1fuUz
sP01gu3G/p57skbPmwENLN0OpId4JO102IYiY5mFv+KLgX71Xx4RLhF0BY2BFeW9
I75kJ1YLk0hd7Tw9SepY0TU+U4bEXzrY+U+Lz6imq6xTJ506pSMVZbwkU5LpTD2J
N6orIp4dftlcsENjLmpMTLUBuizySUblaS7ILN5e2hF82TRFmQWKQgOcJjVUY7h1
xKy9H+1jXkD3GzS7vhIo4hAObqazgBFlxb5SfY7o1K/uVUFnsstmL1510zaks0eC
xBCTL33UvPGOWLo1sRA0O7XQ4vCFmb1DBYhNOR0BNPCmDYnNIUrJs+pXYjavQyuf
E1YDMbel3L3V5sTETAB2JesQXxJv0kyzefNNCsyvV336oTMH1/e/tv5M3phdKLT6
uP2s8eNVMnixKi2es4aQOwoY/AY/ukW1vSganViGtnWF//OyRvbgoD6YFsGnT+pB
VBaSSvd2PihG6qvRu/oxGjn2WVsF1y0m7pcPpLvGJb/Zi06lnAh/j6spRAs9ulgD
J1kaMCEWIniG1ctD7mpOrlB7CDqYr1Jwi6cB5KEu4uVmu3TDak8+31mTpWPrfTUI
Zbe+UR4MKMW6wwB6FeaUSR4n2OntDr2/KQMOVYFPrSY0nYY4zaIyYOe1yW9iivGo
XdKyuHc2q6IBxedy5vfu43Br+YlzBc3LqA76n//xI/vmB8bpgyosNNlqOl8Zl0hs
DRvK/iJupdJOMtrfOXm275WVIFVpUryJgKHFeKtMYK9eh7S8H6VtqAAJszqHRWJu
9jIPb0u2g+O0sNgh1l/3Jc33Eefl5EsrTRqJFKQfJvbqEVLR3WVG9XePM2e/AAFx
2qwcVOEdmYAXH676Ki8p10ks+QRu77+Jkaga6kRYG4+5M2Rn39TzTf4E0cwo9CtW
mGw7m5s/g3h8M3wCJBw+qr0JHlNO86WJdJKLMf49vnzKc6YAR/U+GVW/gcBVeUOy
wU5nBP37KlH+igvTm6RdnLeEMSBMhFEGMWnanFtj/fVgMvVQmx3/WbcrKsvhIaWD
4bCH+EkSDOaTr3tIDpYRU2wubHYvlde/H7okxh5XHKl7w/2p8x9M32yxAQM5Hpsw
Tm1qIyFXncnTT7UrInHVcb56TSqTE49fxJ222+R5ifm1CJOxWAP78uKNYppX+sgH
Zw8fCx/xbDw35gTLeSHvkRqGRfnPH5GV4nY28dYGqOaMtTMnhNoK6XmtMif3RpjB
UpDLmX8RCg/iv4uaT/aKfQoMW9S6JbAaZwV4C1hKRDNkCOEeQyeD27EcWUZ1b5NA
E8A1OnwxOn0VvhV7vm71YpWewiSO1U0pz3dHXs3lC4VJHBbSRIZ/zro78rguHdPy
EKfv54qgx7LdKdBntXcsgMdeZR3pDLROS5I/v4vN9ZJrd2q49oixumfEQneTXLla
/gbnRO281jRQ0xQKd5LawiPb9TqRWD1yYsfyUqPY1Bg3wDIH2iljthAJqRaTtgSs
jpf48HKKcvUWWvzr+v/rVuPE9G2StwMbwLBVsrsytOc6BUuBqpvU8BUKfkqnt+5d
VJuLQdWxiTYjI1rdgkF0D84OE4It+S9cSfZzOxE8+SKNMSf023O0mxKq5AIPUIBe
rBlR2Ub6ddjM63lor1M9xAitvXtThmjyODa7MCdsZVexGjDymWeyhrpAtwIwGwCQ
EXVpmOxS8yGko52XdVfbkma1l2E1t9YRtiZz1O3hxPL6eri9jJR7jZFAmZPu9OZ6
+17yOLMP/zE8g1My7L9rit/oDW7cT1cle+Sfvj+IhgUytDTFsY/yyFoUsm8ki3+N
5PODiPv+Xby6sZh5oOV1c8NKFM+jft9j6zsTSAHqNvFPH/+3cPZORszSONp8uGkV
kuxObwqNKZ/P+p0RTU03lgTq3zN6Hg7NcbMA5XdQ+hnJh/A6LtK3EdnQRvAx9Au2
jXjDJh2t3vDrlJ5/vEtuVsON/ZlfpmwKqEAhnAVQV7T1Z4tQF6e8u6WboVTwMrfX
pzclVvmw6EJjg3dD7CCzTOWzrGYQhXA7bS90WWfhboEIc/bt8otLxghqHLi3IQd9
B86LVErRMtwoQFO85e/V95jC1tMPt8UFG5aLKSPUQOmniZhAktzWbf1l+HFQI00E
OTLpdvli7dAnjYwkcudwlgkOInN9cHZsSwv1Cps3psg/T1YF6JIeM5nTjegvQ+He
x6ZzG6t2VtgGyBSkwKMwSdyR0SIlGI/OgiX1r6gHWwPFKP4o/QghCumRaa3WP2MH
458kGa7c3/5pv1b9qwyX5rzixqZY5G6IDoneaMnMtiiL+DFUKfUaLID2LHj8o/Hv
kkGRqT2bLYWmy4mXexMrC/yuITG55DAV3SxNOyebNKcJW144P6/I3KOzY96ZADeL
/nWnBRYlRFtHviaQ45GqqekpvA7H/4k42Z5iTf72eHW3UPbMND66WxdWJIigN3GM
Qn3AGBM3TLRWGiXCQI4u38og17cIrCAWXPZcodfyCs3loKg0vYzgfBzf8sp1Z0uR
U+9Rol+mrdQYGnVjz5tDxQxr/YH0+ZY1Xh75aae+yYOjUObbgf2SYS6n0Ge8hy4g
XwZaKbrdTgMOB68pIN2LXsbeoIY80A4331LfqPQGP8heKhS78eof4xmtgL6OqXaO
8ieGMbyndyslAoZJQvqcvOi/odMRQfgO9EHaJiCncwcd1XnsmatxT7uw8Pbbw3Hh
njC1eQDbaOzWk6qnPBazq9wFJPNtP46iL029S6htmld03o1EWMPBAgJZImdXhENQ
vJCmL5AUzXRgfgFOXF9pnaAkgRYBJ9OrDOZP1fIurKzU58W+DjI06i5TU6zJzazb
R9ua+DxuJwb+9OSmGBN85OSrA74tuoe32hwWSsdDlH0Ah9fJwRO1w7CSYXtHefuH
tcQS/JZiOsk/tNpqdGh4M5QvDfQ8h6jd/ZJrgy50bPzc/rDYd4OW0Wn9Nyq4mPmv
RbFjKMLdHeS+H3S6JcSSyhmTwFbnRfFWK1XcvBPZei8kb9KhV5XHQJrSy5XLLkvB
6tAEDlC1Irqw/fEkdjIzjZb1yVPvPCT8zlygW2BA65rSCRsrsFreUVd1neiULTNP
qh5tHoUKCO+Rt6mdh9YZCmrz08oIYG+zZfkBaaap6jkoubLZ4r2LvlfiLFfp/GW+
6pGPKOmqy4RvkQCJsrdPxTxFtjmJJdQ9/tBI69raT9xXvPIG5281CfNnwvE5R2pl
OtIYVOXt/suaol7MTRhiXW2bWJvI5fQpJWsxVY7BYxFTjeiYSbDMB+0qoB9TLm8m
Bfn8SGN7R1fiRvG51YEIJlWHs+2DWzQ6DyXjGVn+Fh1XtjA2i2Tt5wQoudy8zRVA
cbKSuMCdJLFOdwi3C704gMDJaKbuILsaGBIhxY7OSg4FXuCrVTHraXHmg6aboS3k
cbrZp4QXdwtbirKV6c6vAE/taaezJOGP/vY+dF5zGe0hDC0OIZmT9+QfPm27fi3Q
sgNnB2U77AZUm15Y2BvCZY9rC9TEEhFoJCSZjSVkkQqecjm6bs2ReHBdDxHyTfUM
jtp+7OYuGNDHmilnf6X4JUPuwpfEQM9BPn7Z96IVP8eJQiXX+viv6oOoCVD5Mkkm
Ap5usx2mKcVccXmVBzirEB7NGaHu47+cOHkSMhoVD5b3drMwFdN4NQPMsiA79sfO
8/CA8DO2l65QlCdyniGST88r8lYm/w8Tc4tUiX5UVOgPsWVltCXElkKMYyDfv/Cv
IDVT6p3YGiqsrhKrTFt3b9ruoQQ4cBX9z+UL2ey85TCes9XpFTLllzOECSkfeZIL
DS4SaMDC2Lgrgek26MMaZ5JUlTzgWk0cYLisPHrdoAlXXlKla6ipvzuAqfYqMqdG
fpXrGznRubljzH+Qc7H6OcsKlNNlEVDu/lKLOxpgJ3JA6WxIYjeY8jOrkbeoUyRP
/c98XvoUus50RkEb5lqP2r1ZUYi/nwTCtH+uU5LobiEMpwNGySDZOTDqERkWQAb7
VnLpXl7/p/SX2gFvq4VjNkO2AoqUJ35OLCo3Q46QVoJus3bRxrqQOZtIcjPtmjoo
phOi3CrHp6HtPoNp88bi1gEWpVaOJ0IrGGZNCuImJlO4Bj+zY7QrL9ZpERZa6LWb
1Q3pH1gkGnYpwPn6GBkwaFOb4KCADR2IILSL9TxW9hP7tGKUeRDt2LBse0HJqDPn
rQzDzHfoRam9I6EQYoST4WhNNUU0PEWbgkyeklr08M6x2WZyjUKeB6GnnjJeBceo
dPvSYxDtM/kafChqfkFLAiIk7yJGugQCHeyERfim6rku9XdIQke0AupR4ZBqWLiU
Ebny1yRooP1FsMquXXO+exEO12xRKMt6i8ekqeN9Uj6YnpqO7QmMY9gHBNqkRCJo
VuRURz7RR5DxwpMjS/kL2MB5e5u2R+XkgOIemJZd37nfLPMUJjVrPSL4UVNyZrLu
gcadSrwWQUtOJK5BVPSxgFg2i7ePwV8wIobTCxT5JByb6UtqK59yOGDx/e+F4kby
oVAb6fYSvl/9wcniYkSQA3ub/jASORGBmkywVROI+04iDlOk1jI+hCgSQI2UxgrG
aT+Fso53r76HbCzlKK6Cv/wok9HHuDnHdU5tD2yaj9edZGiL5OKGiJKqh6VYJBXY
Yt/zvM7JHLKwL5xl8CmnPB4IZz7tWo04jcnNpVz9yV7O8vZ/pEks/3+kHr2NdJfH
Iu3pP+n2xN/Rb4uJkBXWpAK3we7v59T5ECHp4Sz1avk8ocvqnxERPriR+UbkYAU4
3/RCIF/ABT7t5dTMOtmPSM8WBQwGUeLpf2N9r3ddMVBlyjQx/60tIB+t5w+XBIYa
iG+e5qnz2EX2YxrIxtF6Hr6QS08LIKw2RaEErFqyv8tqNifbQwe1pFm0Wp8gueiw
z89mdfV6j9m2NFGzXqcT0dOaFkwinK1Q49cNhpR0bXDZ3zxxxa8pZUwlnB8tjxZh
jqt/gdbtIKo2CbEOTTzchQKxSe4ZdBDIWmQ22mpRsoKlGHyXiHKl4LX1RP5kFA8a
XVVPjVt8TMIQ8ae8tXEYsrbCh7Q4Jxh/6ItiJMFRUVDTE1ZLpYVTZeVYreb6PnCw
wSHBaX/kNtheJMt/uht0MpceDAtH/5hdjAjT/uKZIblanvfEMhcC2nswWNA8uZGc
fT84fAbHrNlCdls1u9LTByqggfSahbPH07j4pfXqIzDuoxt1xqwcaO5bmsTtihfr
BtaaMx8q5SoOt3NJO3nyQB6eebOIgmqHtV9l3YghPhzfcYL2XCdlvmIan6+BdI8V
J0+qXEEg2hY0E9q+IFb26qf21D9sXg7JL7x9UpFLlsG7GYV1IwP/hHHrTcyznLfz
T8MwJHj4GaCYQPa++9eplj1Wkr552mDWqvV/1m3YM6wtsW0ofOIWstUUBPsEKykO
/77lbtrOHztKpXCnDgAgksKL4KYQ7+qvpzD5UA0oN6l9c76PiMY7b8eGjsQt8MgA
FOW9un9VnQtOEshYJeMME3hq0aXtXRiHm6JXwutrBz23FDaThwHbW8S2dPsZ5TnR
twpS8Ws8T/cEVe40BPwKwI2UOhgpAvIurjts9XlcT1SRGyDhGuhMB7TyUAnU1Jh9
rgKtcEyR8slbbwwWxoqT4HMZ+xIifh47N/l354BlZvdoWJx/2cuUAQLgvG22mFc2
bw3uJF+m5Z/rub3eh6W4CWxYm9kPnhfrzqy0VvwDuWmEs41mikPVOhqGhusxNMNL
o/7/lTMHPm4k5ze26DZo9AusOsiz1r/LssUCLrSdEc06lRhr3VXkoEXClKWbIkqx
zMLZLLF96LkfayzXpsDy3nlAt+ceop9DiAKvvQaYZVuZwF6rpTH2oLWz2hv/jCHt
fNMSm5MSKDsnCAwlKqGh2jP3jhQXtk9KpTd2bFhOf19IKLvlIebCkLB0HynwwINd
qgYpsHSV4Rh8UmFCqhERcx3XcSWw5ldDjx76IPRAdACOK/NvguwOLi0MP+H9h2w8
CgdG8/k660xIXkS0KCHgLll3uNE3oauImIMIraHax648U6ixRfxt6hFH5wE/R2Yz
4siW1EQTc6twE4505ujFHTtTACyNZ8OapIPk0qHkLyM7T6OljpNniS0BIqwz8/yL
XSFaN/746HV8Vue3545aIhm4DvqBxdKrzAU6jQUP6ODtW56LUii8mWYBNz8GuS1M
Ef0bbpkeJM2LVSdnjTJFBxL/oiwI7CyuG3w+ZplXY/NLhhybPn3dzzJu0v3SK+0B
WHjq35LEteNA5/dd10GAUKqwgUVcVayK60flZka6vgEMbTQw+wHw/dUYEO37KEPA
y+mIGe01/ZfU8TeV4SO7uxV5XB3gbebDBrGNwisfHGif/aAqxToF107YSMFfTaVG
K8qCjlfrT+z1UYGEA8/zLIzQSfi0sjDf0rhHMstfX1io6ICAlkxApxEWDXdEWRsI
6zD7xVeXW90FX+RROGZroEOvIB6lSM3kcj6C4ivEXAVRuQN46ISngQKT8f0xoNpY
JTpVmmmIT0xgH3dkHEsO3cJt11Fv71qZ5ZcjShkq+69DtL7GwbUTyljPFs0ddlnP
E6pPH8t0rSHYHNcM1woJDU+66h/waQ0Zlfa8326u9zltr4LGBEr2/D31uN2hoAjI
I44gqtvRiH2xkdOqo66btxZMgLxAnxezxD8Q32AphyNl5WZflHvA+0o0yPfbJWFI
EtJfrgVMagEbUA14amYkIw6TULG1+xHDRtETXPMCK8UvY4EkSe91a1Ou6J4CqjXE
H9gSX1kBpbwdXzYwqw/PoGDw2DhEJ8Q6NwVHMx5IXgLqWkV+23Cg8mPMjJue6SOK
NuBiZZpqFyzUJWLlYAFBFtdV/R+Rp0YqeHiR7qxrqkJKrI2xwRWF2vBQKOxy2r6d
Yut+Ek561tVEVh9HVbJG9j4ZaN45RcSfAQUHa1fe69mc6jfqQihbcou97FdxpbGg
LfjCsFUjrBLUWRlAS2mf7jpg5PC/BFcurqDB3LAcd4z7VFiWQj/XOo2kyAzplY7j
tizq40PCdC9wMzPwJfMSQPnlYlDqM0XtFy+E/pSAdWXqDSJO6IYFpDbDxi24tl5a
loYcBO/TG8aiB+iAEwfmdJtyePA69vm/WO07Jb8UfBAEHLO7EFMBoDLdSho+JNI2
sFc5llc63QwXoJAGcaYr+IjEXoVq/0ErG6vGwRFb0iJ3pqhFAfKKb8jO8iztuYzO
InV2ar60p7CC+oz7xLPRTIhbytkcW1JxJGvuB12ykuEY9gmYOFPDpEadkz04UwOl
SP5SK2qmsB5tNWVAAkddeBqsN7UVdIBUcPoFdF0gkOZ7S568Ud4bKdPeTkt3Wvg5
6Rng/IzWpRXLFuZHGWjm1FJK74QqgjVV5uIvyh8Wh4U3LbH5zydvuQDICwS/V9YU
SFL7TWmlOnwgxGy2xZJoxrvfiv8dEIPwQWiOtWMHpf1IyA45Ynt4ug0gXDKQz2A8
Ky91KKelF0tQKlNJ14MebWERsUA+WpdWwpoZ5zYddVrhhfT/6c3yMUKWHg/QvWQv
KaV+2RXTpACHiqyd7lNevyqh40mC3V1SPAF9/4HQrDyiggs9gDk3GE0vEG8Wv9th
pjKY+rzn48WySh0RJtZseCE6LQ4+vMpfoA3I5A9yMUeD5P+D5XlOnWajWZSp9n64
x+qatjn0Th77HON7uKtAlHutWV+U//x2sFB9ubVNiDbURDqraJEl8IGgoUNvf6gg
RxqyDt7+udH3Q681Rz92cMiQ+kgJogxCDKFz+wXCr8Gnx/0qwcgZREpm3iKBA1ez
FRO58R0AcCQgYzbO7g/iBvwa+KutN3pX0APm5YBeCI2YMi+SaF9xqLJmiCUXRp8l
6hsuUuRMBuiJhWdPIPt8mKWiffDl3ee0l4pXPLriVIwKXjqTm6uwiylkXeJq+C4D
aM88RIeERvwzR9F3uOX/IUW3FpB2HTXrbvUpGcL8nDakiXpPXJFClQoPpRJYT8Os
RsGMRfoEnoS7b8hqGkgHrogKQPF8UEAeKxR36JTHpzI91nqHeD2XUVHDgyyrqz+I
a6p0jtZBl+iQyMiOzSrXySxjAY8DQvc3d51lY151tRG6eXi7VL8Pvbl9x1v5mhtD
Y9oi+4FTQNzMHi3Fu9g+YTsHc31ZKNZw1HXRhG2VBuceA89r5wchmrHZoKgGsAvS
SpJgaK4rLzUuOseqajsW4yNfph2xilrulMv6TZ3+wGtOzxFhD/RdIG2nzRd4lNnw
AWKngO2V47e0mlqAuT7BvGKGT84/KaQKJoi5O2a7oxiWvZ4K3oSU8SEEtSA1Lphr
vFDBRAySuUX7ic70XogVNzgR8g6SQ4GJBDpgGFHKKCsUi3dkI9Wnsh3pjMZq3+1+
h3oYxK1mQtzH1VytFG6JeA5brtA1NpH2qJ+Zrv7DR7mzCZEG9RJaZuZLTTQkX/qc
n2gmLtv8XcsNd/QiWzffLzAuJ2gxufv+00A1t58R7AWBQizMXx2+H2TVrhHWPQaz
k8djt6urXUEB3wU8pTw/i80vWE3L1GlvJnRbHgv2TDMz8W2KR3e+44tQjNmhnbAp
k2F3T/Kon14YiqdQ7yw7SRDRoF4m0PcN65+DxRvN12k6iDMxmjs2RdVmapZBpxyl
rbdcVBbcZonFQhsZQxnLbj8hOC0gp4DJ77van7rJpPZV6M7wOAdKW5X0y0uuE9A8
LcjRQcuKzLOSpsazSz5AvjSoDQOd1Z0pefgF89jsk1otH69WZqtmC4zh5R4wEEti
3uVsNTRXY31yKRZpL/2DelFm0MDSM1XhdufVSfQP4hYxTa7vaOpotSpS2Xa0CFtR
/b8dT6yD3xrbtKri7ZJ6PYj1xpl2BsIVsOxRxwfox0FxvCa8bAV526n2K5SQDsY+
U4V3ODYJ3ABBz73rjMAjyX4ri7rnJX+Z3iRTNu6HbXQXSv5LQBYUdZL9XA+X9Dtk
saA8hx8v7YGvoPR8UCAAkOO4wnub5TgQIbRzHgI9PnMt47HJI1sCZ0ar2IRHQ31I
58KU2Gj4LxdDkBwHEkCCdGWxh0B/LwOHB696W9D+7u/VFEgfVSh/CKwqxcJDbXZC
vw7Uhyxq8rs7T+P1Znz34Al6bbgYx1SmbbbmsJbWwXxzCV/PsCOQ/FvvBZERT0/s
HDKwntGbND1Y0NGjgB2XELZHKYP2XxsHee/TJ8SMhTxbo1/Ei2lmppL4MmJyAHRV
7+rVn/suxmhYbAqlzOa5QO9if9dAM2tc3JL4Ee+GgnD5aEUpiM+ex5gbr6OziQiA
2/fF9e+hf/Iu+xTlJ5WgtkmbLolZtA+QY7G5hnQ7Wr339G7jwGc43EQj4OvTtJB4
mDnvSRV3CaMPgCfeND7cZL6WMDTIHrN+rjsNFGr9Z0pGDtDFgKPLo9eRt7aA8tqu
8Ef6FAzSLbbWavzARC56AEm9HYapnPQJN9m3jxX+Pr2ATmlwUFfnDS0C5Sz7jsqj
YF0D8yXAM4CnpoN38zDFGp+hXyHtaK094wLd1dIU/e4ywMssN6dvRfHid7ff2vCV
Mae2xC/aDmefbqwKDNSTOT8MLNOSjJem8I7jNljgdnHuECzFxo9O+LSkJky8h6XB
PIBJJZzRdTyaz28fAsFTUVDm9fx6NS3SEX0wE0xM+DweQAm2Ju4wkaUdlOOr6cIK
/d8cdVArL9ZIpS3Fkb5Kd43e95k4GskocFSqE1bHr3B5bXfEDFUIdIksFWakJnqh
9K8Fd86VVBmKnEy9JYBzuMjNQ210qViKRQTsWXogitUv2ZRMR9npPg2ou9Jxd2uW
2EavsPEkbnrvsJOMs1T38WDvb9OP4Wy5FAuSDyfQ2RCFbfyBk79Aej0X/bEUN0jc
P0PPEof4J4koWwrhJ8Dj1+KRCfROWt4stIk1Rod7TA3o73ogmx9MYtbFwC64O/2B
M6yB/Zho0M4jwHthP11r2ghyOz2IM2VjajCMYGdlqTKlNX7bXVM50IhXfAKmF58T
XNwGjqulj8e+T+BYJt6weEA/YDYEaVF9CNOGqOdF8IP4L1fUfSWK9GlWwFfklTtI
onwDJeyNPz64x3QnJbG5XCdpAupBIrmQdQ+YMmsjLw0lCj06mEQJhRfrBWNwVYtv
77kSVQJxznHkBVVxHIIleCGL22DJ+ccYqxOeWjpOYah5iuBOfIIVbjCN0+pjpSB+
8M3YBQO5IMfIewp5f0POKXDu//XGyyjcdDLYFmqa0ywD5q9EcXDvkV3wgFQpAJgi
rPLpKa71vg23rAB3AOAIr6RCG4lRJ8tCNRO+BU0uzpuD58gOh88ofZTEPKT60lEH
HFam31UIlJafutygR+bH2jup9KUOvjL2OczMz/uFn9zWOzStFrXR+ZhTppMGObzd
JgAl0LpFES33MGIEc6u0HDNaABaLXH1aiCCZueNJWENB4tqiqx0qdLqy98zIgnoq
5/uRXMOU86iLKrc86+bbIXD4Q3uLlkJnMWxVJ6YJSVeXjRi8RABkHu6ntckv2BZu
WwRxWwWU5ubKbx/DiyLGTenk5kyzPN16YOKQ3BL1Xsf61n7dtbag36hM1WQuRaDS
leFcyBCX3q7Ev3fMz4D7IByk5xsttdDPBhaXUmm6KhKxmEGWH8beHW/50qxO0imc
ngiulnIAPz1Lyt6DiNFj8ASOvkPEtsAPqEZ4Da9A7D+1AZ7usXMTVvLeU7gOY3cn
jf0B/oSiijJj8q3IS6rw8/XnFC5Xs3pM33JEQ/JLw3jAJ/LcZR+ypDc3CRnNa6R3
sdrgEeQ6u8tLGmdz5eVk7JMLsCjRxtNhMZRI9aBPASOvQRpcMmhqfEULYgaJAhqY
hzRGpOy7gNlIx7bXaaVMaSXqshZtXEc9jS4cYitKxw/RuUS8hPGZ33xAsAznkDX2
K9ABrQlQHlxAXj9QNqOLsVwoWv5cSX1GBGLpBB/fd3TpEw0E1XPjhv3ZMORkYEDq
kY95DG6Py7gr9w4zOWBgVP0E66iPC8LyeUeJv/bXGJe2i/wUtB1Y6E1FOhJDw+Q5
XaEFGOysP7ZLpY1NXzDw5LKgMVccw/lqFKQUSU3TFwJuvnVc/ndkQ6qp/ZT/BcmU
QJvtR39JDrTlOSfHK0PAcND+0ceYELRDa/RR6JnGhVi65/Q1RwviR9gtiH2gHnLV
gTmuqGd5iGrjThXACO+61qdmdKxIOtRj0Ch0NutBPuGVVmWd62OgGZehzThr2sHN
imCZ82K1MgUHunNkiTShHYaLfcjRHnXOvD74s7YPFgx9ecSvBhZV2z+aRJjdLXjI
jJ40HAZb0QV/jlwa/CYXNuLcTPIdukwCQA/pt9ByvuvY2tyHy9Z2p8t9PZB+hpup
VOIWVh8fEXpgY25n7XvLbbOSIWMcxj6ido15xflnRJkWH3z43SMvRA48s7F4Z2SQ
C9LXvBqXR9pq/Rx/3K7BnMLDQSHnecYUyy9ufIuQpBYKVVhMNdU+c1dJ+OnnIBzy
KsRrr9zosdGXGbfxgQ4gspokZmhSzC5WntaJBtZ7q2yx3mE3g5swVi0H1lvS7Bqj
qhZRgJbfTdkykUJ1alDLdkaOX3n92TH80aI4ll5Wsw6fCFuA7wuHZZnWNY8d+SzF
rgqIcVUJUZ9pUu39GjAPTjZDZI6oe/nL8Vy9xXZwP8mEk8YuXI/fw7jeMau9rA21
hprHMYLB6+JUul16XmXRB/1WBDR3dxF4BR17O77c6gCa7rqBJyRLK5qY5z16Jz+U
y2V31j8Vc1sH7z7vqQQFXATx/TAiZN5v2TohdCeSVrVsmSkSM2EqWF1ziTCwh0s/
NqWfsxJJ5epvVm2asBkWqJOZZ7DwCtSvjPMaUUDN4ZSTGvQ2QTRw8s5C7CTxHmhJ
qTWW5WbOJiu+VKlaE+wcCNSqhrDQLX8mEaLsSIuSt/rfezaR99MHeF1z+Qk6KL47
P3RmmCjfUc87dn5M+Z7f78SPj+UvFtFVjRZO+1VADhZGQY8+O9m93WlbFEpqzj1v
HRaUVf9W6AGCNVhdeab4lZbi/qygGmsQr9trTVJU6ktSAVVnL40NA0463CchaORt
uWdDTyvbR0PXKH3GwvCytMawyyot/7i0LFcTF9noGIellZi/9q5FE/edKEKRrotJ
FaEik0xWFf/tIxD/FYmkKlNat8uv9nnwMtM6cZiygQJkWPiBqD5vJxR57YdtBjG8
G3BBGlp7WaAXyQ63uFfGT3Kimz0tmIMiJh002O01kA/T3SwZAk2v8zbhEm/oUMVt
cSueutZ7pz67WUv0+GmsUwUFxJEsbewT0FPZC9ldJU5Q0hHBqSN6Qtzo9lCAB6KY
a2T3eMadhgZYXoEnypb8nT8poThi3iZ8L92znSp3SMHa/PR58e0NKl1J5kukI43O
QT3SZN6gBzdwRYEQukmdki3rCvmB/Ddy0Lk58Y1LhvJ3hTR6zIua+hBXujpgMAUn
PNNI6VBz3uBSRt67qr7RjEVy86BAbnTfTrAQBHgVgpa1R2fkC0UaigSWhr5p2sVk
XfEQexz6kMlmPuE80gqOxNKiF8vJW/dY9Mlb5vAubJ8GxrCdW42RNonyeMiiMUck
e+ny/YIxRHn4eB1iuqMzJf+xwPiaJhcC4en0s37QXu9Iw4B8nV2eaqEuaftBKQDg
tcs5jnKHh4uJgcylsCcUdDJyn7Sping6Nm00klWUu2RKb7pV2Ryw5PQz57504RBc
WsxQEEqLz62XTiqQWXWh99ANSJgd1KoSkfxLvD5eE2598P6FNaU1KSSkVb5YUqvh
0HzT8cg0BW/pipGkicXpHYXNJ5ld0Yat76+OixRL2dYHT5nQtlUAceiy68h5cCcl
Yl8pWPtn1SMiSDfAM2farhRvdCntVWNhKAgPxoE7WHgUImB3N2Y7f1p/hl8gixB2
8rO19i76L0RY9kRjx214TMCbPHXVWitHkutqUN1riaWy0B/AnkYpIcnvai1fw7sw
jqmxGywMo/QbGlQ85k+JquE4x8jHnMax5YIMPt6ktWaIFYTIZZ0hOFGfhfKnwDti
xJWyZJom3RjqJDVP9daU1Yl9JHmu1Yi6ALbIukVSefF+oVxmy2+wnRl9mxuFX4lB
m4nkNOEliN7KeOWg2TRy5fW9nr5nKDHA0rcBSj6lQxfHSpm4ab3lIanG5JS3X9WK
B+b4/gF5AEuSUIx39/1o0CIGAxaf4sSdh0Ze9YiwEjnQNarsXnjEy8RKRVNus5aH
M2fbg+GYSOJYDfObOzwa9EH25xuZ+ACekDhwwbxcBb7LR7ug/1d4ttJWK3bkaoK8
nSB1XocRNA+/lsnxfxxkbpMUUew60i48GzDapI2uf3Cpqy4aC3aT82VJoen0qBri
0oU6cqskGfcaEmZl/kB/gmPW6dbVDRWxLMDfxND+Pwae2O4UdLSB8R0U7UsKh2m+
Nf4IigDqIU7YrGu/+ZEqoBxEnA7RmWeFJRfKee3z0wUk268WdFS62+pI3Eref5uy
iB50On4JJOGTBc5mI5S3BchQhDH2KEK4Mp9B9rFRLd2WlXZ05hF8NfZv2wuOZ39d
AsNU23nPzJHFP2kNbKdIlWc8NoxHsYYaC/hzykIdjDzl1eiEfwkA0GFgAZtG43s+
oLp5Jyatcp1uxuZ+enr8zSR3tqZ2ltN7R+mQDWv+Flo5BUnptxMU1BrkVGF+M6et
mHvNoYJsJpYEuDIj61NIMmZGibAO47vYlkpw474fqXsb4AssPa4UQy/UPlM5aurc
74GNhNIqBB1qY+FPszDJoC6iXW/HAAU/9rrxa0qLeGSMbJkdhU1acI+xLIMArzhx
pOMjlnc89l/H/LU+kDvZb2yToX+TYWis5lmVzQ7nlvjnkGT7/JzQb2EFlvJtmXjp
2XWloJCJ5P4VHzYX1GNzqVtwkCVxQBoQUta53rWTCDWBAofPWTmggZWZSXs+ADug
I653dKJd2PZbPJ34+OY/zQCv6/3Rav0b6VuIXje0GFxxzLMruqcWBpRu3vDZ+lEb
h5l4ngTgi85okYLeev9HDY34ULl5aeODzlilbxDnTtWFUtAA3FQ8AS0XWpG+NM/0
C6ivL2oYYx5xBEKz2AcTe+6RDQji6G36T5D5h5HxWG1Gq4F7aM3hjPXumodMamWw
qLAgfYcqToWWIvfyfcNu8StigDlNZvTVkNK5ZfvedkzEc5tN0uSlixYIodS3P/Cb
fB7RPvhyuPSpmzt+w5Yfhs8+6ytUuJ0euvu8nuf3lu/udOAQMB3JxoabIXMwMGn2
peSvlWdUbek+Qi87hFxRMD42yH9AvoInU4d14lVwNG/WW4MAbgJ7qc31Xct9FVoQ
7uRfVhvT3sAHDPj6qqOSKE5BKc4hescptHNWsIXbn6A0vUlZEHhse2uGq0DVb3KH
/RR8q0+x98UJFYyfsDLclAX79ZfC8YPiiX0SxTEgbeFOHwfTjD0i2uecaxsIq01/
DaoOyJgSYoORv6ox5ygPaW6NHQ6KOFHwADazk+CVd0BDU/R2nocSOlvJFv6ZO8dJ
ZSA4Xpw9eLXSebJD7ZciM/NmBMvIOFxvORTYSqz9HQHu/92iGosteJi/bXd6riO9
y1a//e/eC/PvHlMYWLHbT5lEQA9wpfHDb3GqaQwLqB9yDlvL35FR8BHVRFvBrwYD
dnPrVZKu8bOU2x7EPYPt5T00ovY45m0VYqMBEzKOUx4CzZoDQCVCOazK6uRUtGRE
dABTkvGJMzVJZcsTF9985uW2RC2Stb4Wj90nwwbNyAMhQ/+DAW2vY2Q6OZoIPY7P
1R3ML85HDR7ji2zhFqRvBXKDvo8BGC+0WC62qbK1gyEAIxv/+hEFkCnzaCR7IZJn
9RTbldjbuolQz/J6U48Q2kRoxlpuxbmTV1BexlR/ulJ4yHoJd60td2WKNquYEDqA
U2+HPKfZ9UmkChVYveKaIIozbOy0oIjf5JE5Ax3SpzzjMu49TY8H7Rojdk0tZWfH
dfJAj+aqDGWMBuX/eH+XjCefaKGUn5IO6r0hYWXjoVqWbQKUobFAAbiWY4G72hz1
3HQyrlYcxyA1IRnCIMKjp3rbmcU8LY/PjiYAX1MXuqOOWKZRik2qGNv5Hv0Xs0M5
frv3wcKbINCS+V7LgjLxTEw+kw37onz8xScgYMmes5XrgFTXesBNJ12Db8gxVf0S
LF7Hic7G+pXFFTjGaKv0gGo66V2aahyy8nJL8pXNz1lL1LCrU7BBpxCwBBwN3Klk
S4Z+2FBt60eOmVVFlMtoxng3bDOK1tfhr1yDZxOsBqdKTAUzz1oheC/0YpYydq/M
8wA0AdsxGNbKDH63vH3q0quHzN1ya7qHe6bcvP+nDJeCv8APcnDXwNQIw/czH0WT
xeifMNmfyXgfKmgWoYhQOSzWb02W/CHSV8sS6lklC80rwXKWnai1tg4iwXhnqaN9
zCiQUFmBO8VqEMddQrfSiRC9z9uoy8BYjLUx0R+COv4PvY300VuTMqsf4fSPQFog
qzw/ZOnKw0i4OrDCCHQB3vNrH3hL+X1Id75V9iuPvCqqEQ+wUF2cm9g4cl9Cv/Wo
IMzr2zp74Ny7JwLedYfENqszM/GAhwQg6K2KpCC/jUCGtK0l2hAC98SAyo08klZ5
Syo8X9LT7SxpsAw07DzjP9ppQpwHserNoNXiXJBzPUsgimNHiVywlYZrlL+CQcf/
ujmum9+5DS1L6W3fI9Og7OeDZl5u8f1eEzg+8ZNyb3nD5WTqq/7j28KfvUw1+RCB
ZsBc9KKtdr8qQOAm3oJ+h2P1XPiBAMHZO+fMmY8JsDNnBF8B8y5ZqGEdqgCYQaJ6
1QtVV7bDX3eXbdH9Couq6WjgakByYgTXnQGpn7Re3pYHrfta8FWa+lyuaO+CqPEg
YnlmAyd6Mj9ra3fcOxRQXiOuU0DamBObVjtqO76N99LYU/mzQ23pkGvMZNwMqnA2
N8G0C+xlGY5Q9xsRngh+0uCuy4wt00IIaOhFYHU3rLZiBKfO95Njqmcgyi3SOBUO
bYTp365IrB1ntqVrD2JBdx/hY5ynDSl6z1JXlnGaV9RirxT1yWy764NI1oHAhqwd
+nQIGJQOfFtaRk170S9Lchp32M1livQtvVjfJEab7T0N/pWZpsUs9hgda+BOEgk5
UXkodwWQdYmkLh4D+E2jEAWb7627yhyi3FgA49z3XtY3Pj88GHE8EBdRAbIXxg/v
jF03FZogM/a/ZrIiUNTUJ1f3OnA++7T7CafdEyWuCmFE4XWGor6bSif/VfLZkqZo
Wq839Wblj4UeJsjE9e5MVxVNnpLcPtoXc3OMSAItqeBIrv/DfCWoDfUMiGGEtD3k
T8oV5OsWIFxyNvc6m5NZFQH7G6sTqjQIGhpXaNAORz8RpVEncaQdjC+jnQt4Kib+
jamQJkq4teHAR/yu1aCS6rXKZZOhm6PurWH8zOmT05ycbYbIZU5NrilcSfuZ2/DY
wDuUWoa1vwyF9/cMH6PA3tU4nF+aGOVO59IuI0LrWS+1jUtmoKCPeLfnTFDgLtYw
Vf0gt9i/O+TO4s66O+e7rsPSAmVK2tJTcIL1nKAKwDlHbwx4eJ74KnzQtdtvTG3Y
kjZUM6n/jPitSKNNqhqHMr7Jrqig2Vm+ixtL/lGdxttH09wiOa/PCJNh9HnKdn6r
wrZv8hpU5N1rnEn7nv7b+Eo38GpEIbn6v6uBurWy0CYGHHdhbLL4Q9EdNrJV3G3+
dKD753TVU++eCYcGkf4qqUfR1fk0eg5rwtVrrgIKK/oX07iqhWZrErNAlJKoxkSo
Ie7XDSz8hZXMVrwt6nlgivGrlBDLPKw5ei2H4pLV4EUGHjRXHOTzL+db0t969fVH
8Ag8vUcwYt6c8KMR8SbsDrys3yGIWytR2tco65wbR6jYNyw1A2zUU4y57FBwZ8Rv
AvcgwMX8MxKmAg0sh2jTmBZxiYDsuAHM98yandMYvlkTJjtw41efYIEvTeD20ypz
ab12LKB+GBbWMA6LQE/duttPiKoYjOsWblnr9HqSWt0clA+qrBxEAjhqgFfJhbBl
pMyY4DyjFEY7D4BhOq59GdIX/IFryiFbtWQ3cPQN5Gyn6i3nD6wkg94lJUYFLmjh
Q2GTsHh304Yk4uzxRD+4h+2LiL/NjJ0qobjPWAvYhmrHrWQLZ+yD6B+63+xCq3r4
4bzmnpmuC36O0C/8Xg99yLRTzC7DYHLUpigSCsYoVnWWDDTbdE3wfAuzHJHEDEM5
xAHZYcEX8fKh2tncCfh8n8s1M1DP3XLJNcFf3TtBDSq90qA/tYg71qV8/AhAEJm0
RBdTOYL8B+uJQrlNIReCzN8h6VRlBrgwRx2om3Wd483VHSx/bT9kjKVOLTAU6eGH
OSxBk5NzvcUHoGSnJ6Z6an7DLrKgIPTZISUgtvTqEIrJGbOcaKO7AbjshQcUOfRO
8zs1IzkRovEvcvvWpk+1+zQul1a/Cx82vPQMI1RoWekCy4dgygusxSWQoegrO9xU
xTosq0lCEt9vjwmXaxsE7D7eGvr2AxShFOBaVdgVIwdlzZCMLPY2hoWN+86P9xy9
YpJO+2bvXYD73LjaK4nWAX7L2EhfUgXa9QlIyWLP0yRm03EB2x/Mmka7S27J9tkG
t7bzucgtYcHc3IlbvkZ2ZqufhqHc36GjDPgS4ZnMU506Lb7568ln5vGZwp3relvk
nu0f2lZWIsK9T4ndRSur9EFxv5+dW8u927bmZPMMH+csE76Muj3S2L6bbe9thuDZ
Hs0msbWp5M/S45M/MYICB5xYdAnciiLSnlxA7jYJh5pIWTcGYvtBlnkPYAslDWbA
sDHnCOf2+tjgK3YJPXDK2UO/SzCObZ7FJNEMjizzf2sO+65ahnLnnhSdd8U1GIhA
p9ZCluQ2Mhmf+XMCHvvCuzrZVfsbwyp1jazBSX9gimeWkJwLAuBUy6mF8+2NqK8E
swEUdjt6l6HKcJJkfBtpjO7nIKdoekFt6I1gZhSnoQ18dKedolepNCbiN5kGZodM
kDdb/NsHHETuivr6VqduB9ZpyMexj06jn1T1plNAWegg2ygO0EOfyhixBsBsCb9K
Ha8bCqYuldTPY/axhfXP1r7AmmZSP8pJT0yNt7IM1lLtkfIh7C3yVmovuTO3quBy
bs8JIW8dsuxgARkgsQASYXJsGS46/sNPapI1+4mBqnon1LE7fhA1ESm8+qusxKyh
zVwlcd/4C3ujS+wBCno75X4P7c0wzlWHirsw2KT1pR3gsxTPq/UIuS6YdWDlfs81
i78gFgOCk55ZW1kuof2IY8KCqBguaN7IfKNGnYQvHtMSpoCaXBdEsxbiw6h5hssJ
C3OcW1C8fZKjRpctxA3y0duuqvsML+G8FIw398Nga8ReOmvmtwDgkh1vIeuIztEt
yKzj1d1kdElyAfO/GJQeJFV7vBrmwnlhfsR4q25n+UvMg+Pwk1pTH64uefWvAYET
hXLlNErSz+PQyb23oLBz14l9j2GGIt5AqzfOZFysO6hWFOaInemlQle83u5ckjs3
FiDRr/QAKhZaxK140qlBcJmNbmVC5HSzct0DUe2gWazf7UDGJdD/y95aAc45zqxf
scY2sUgR0i54/k+IurBZXh8PqV1Vbh3W7b66OYGQObo070LziVzgpBrAxEoBd4hV
6z493+Iss6trVmvQgoFARE7Ew9wmBLmNLkkqXvLe78IKvgArAP7M93jP5Yn4aB5s
vaoQZx2fC5/IQ+wMowt6C2MQC3Q7TzPnhNDVCPTllxqQML4hBw613g104Pi5RM82
Qz6OPmXbLxgWaFrgkqoSj0XdAxxFtsIaNElvtFJdVfoEdc3ZwaR7ZkBI0ZztcghP
bJB9dKAtBXwqGQK7Xuy2utlmYvGebO7NhVhpnrtdVt9G+mcMeNJEpyxJBMoH5dk+
M15X78cnHCbtzsBjW2UtVB7p/kM3cw5WqrS/3GAInBBeJOY1qhNFB3ZB1TRFi9B8
geeRLWEFGzMJHQfHTupJ0zRodqjl/P7hnPjzN6COL+hagnqDzWpqJ/eVS5w+lT+l
rwO1bMzTfcS/FMyEQw+W8N5Em5wQ3ezaGKIDgtL97AwtGfwU78tjdBXRk2opMirK
elV4pVDvah63LkQ3y82mnZMZt1hNMgHcbbJ/Fq/96rt8Sa7vB6wPZRSqtxmEf49u
vpXiywlYPgWK9sR4hW2fi5592aKxVljryPfJhqfeW15Nc1q1/4SaGlrktGDsAYna
nHcpHFLxBPsaMtNpcKMkcLnedljUAWQff38Os7pbwzm/Cprq6b1x1MzvNlZywLhS
ijwJRt60BhTtCuSMRgWr5AlII5qFs7zbdVR7aytzbY06txMgazX8EN17Kk3gzwVr
/4/k8QslvtTNQl2Mjo+LkMNMJ31YRjAFHUTndOjmQxUwUg4yzyHN+GfXo51DYNbP
e2lI8NeNzycJ0d9q7/HOM3ocxgTfG9A9A9ygmbbaHAEyXIdm/flfLZLRwdwliMdX
qNKCfnue7bWeOGwKV+INuBssbce3fUnj5XQtwOJkIMWNdDpxoQssF4Gi1Bu+ZHuo
toL+TvYJxyQitdgNgwrUKrQUmSN4waLmDBBXktzDdOuRWCtni5WHUysWWQ5yLZ0H
eJQ0v5mqDq9PlvE+/VxtHLlBN7PRGbNB88QVCSQ4U2YNK6CmunieM0UpuRK+P5Co
5QPI9nybpq8wZd0GYFTVVeTP2mzDAjnH3/qDFDVZoKerqHm1Kb3pwBEvY5fd0uk6
kuNjm1eD26GCuHbnNocW5uPX6mvMCJ21wyCSSA2B9hW9e+1GNT6Y9m0i8pa/t3xU
mGd3eZufxizP0eyRK7nKf0jkkGdaolfb0zb7akf1EyfdudOLhxWrbVgOr+etXzFX
5wAVRkDgqW1pZ5JzbE+bj9jy6onfkAdR6ndovwJhU2LBT6H+UJntsb3rho6p1iiU
80TeFpjDokrSfefWxE9amjgelevIkZ2JP4ETovrxHNct4oyvcF+NN7ra64PJIS1D
DynMFkodxLwBwC2x+Ycdpy3sx0ZuoY+zxoqiuozhvXMcqbr4m0VSjp76Hnrz2iBL
zzDkogNpqhlR68ZUko+Lnrd/fNz1WsVcuiq6oZOi+jrySHlgeRrS8mI4/bHFgYqv
d3u9/syaKWpXPCtYo9xum5iyW5Y/UCIpDZmrG//sG1NmGZ48mepQvw2Y7DY5QeRH
eITjC1S5TyNri86JnevVWMVgnW6CQMwgrPuRBLhaWqbpEt/cpaQwjX2WwGaw3aBL
E9MbFgrtjvUVypfMc7yTSvKrqhLP89AJtKI2qc5b/XDTjBUK/xKwAOhWQopwRj19
c1HYaQwegPnvEsZr4caqnGokjUNiNJ0HjtDlrl8KZQlZduntoUmKyhfELJMVUO9b
kF87kPveOixCH/BwXBHAnY1R3yqyJYy5hJobvXwMzwVGiT+T+UVbvmUUVMdanU9o
eUN7zUXRXJk401G20T3Z1iRG0bRGFNojmAVzBor8NwMaKW//ikoXz0dNiiAURQ85
60spnS73n9QlYJUak/SeWtAfM8l03Pppv/0yJY45VSQl8bKPKr0WgnCLeOpSAYPU
phioVkibm4RdHOF/TW4B6mdBPsWt7Jl7rF77Zs6Bcg7sm14dVhxuTZllI7jrbGMu
H3tpyq+ipI1lY33NfVoe9JUjf+xwixBpwCJhZ+9ATGI0tKyRcksyTunh89bNx2j+
wscYdKEo0A/cu+IyDHh/QZv24t46ChGojfZM08Vn7ECbQfk1/4sBhL1amHTiELU/
IdluQ3AKo7op6B6ZwPCgoXW96vuDAXF3fvCdT4k9HKzD7S7U69osvlmv2tWyQUS5
F8IFLE2Cnhmg3VwG0mAePrkc0lxuIziKKZ1X5zwqVrf40bN80vn1HXXNvIypWHIq
KIZxYuAJYBpXWjVMu0o1rtRgwWsMZYhn67ozQjQ2++rTmVJ6ArO6tHADs2I/xFIb
8w9+dMGhZJcFwmo5XSGRJcerqnZ9bV4kLg5j5Nx/AkW8DZfTFaeLEgy0iKue/QI1
w7Hn4N0pKj+vYxX/1soQ9N0jrz7/B3qVzNFQSfpnpd/979KyxBnUAil00wLsm9na
jTVOmU7ozdsBQRdPDb1RjX1LjpJ4xnlt40WXEhUjm/6120u9Lucea+JzgBwBQ9w+
F4TQqm36UIfFJzyYzIzS/tSrGqnrD17Ft9xwtKeucEoI2K+smdhTSCGprJpud1hS
stDm3BT/xoLVCwnXpoEFfgClBQj7RPlP9ne2bp+92bc6nE7nJVcfCv+RZm2nJuDz
4A7MzgC2jMKTtqLsE/HTte76DbelKgtuQ1rXURu44jfMgUe0GS0PFdx6MzAsuZle
yuH/0cR8VLatC/SxitEoZedt/mN37LBQYaiFg3tamxMjop200E6jMqY8uenLsfSg
ERyheeyuheVcwka6dckqkboOcnu+jgZC6y9mpM0aMi1Ms7yCNHawi3yE8E1lyFQQ
8oiRAolYwu42S/KmtrHQ7RdVoRayhff6nxFYnal/tDgA8iiUSNP6tpSag9ar9uBT
34w23Ryq1f/FJSuppuRwR3uapqyLhQ0UTEYrFSQCjxx+QaLZOwbdj9J3F0i5pTxL
BR5A60SjoJlITZFeVYvoZIn8U7APqcehiegsCupVMeu94m2f9D69NOpP/rxeeP7R
+UCdMVzdS8kOu2Ts7GWzNNtaqNZI6rycJsz3/olhF9SWWuu61+VkFHb04LrCmPRy
L1usv8pSEqOQiKoD5QmeHQeWNSicJZwS44rqp/f7QYIUq8SCM1I545HgVyANBme2
TU5TwpWw7qD7qsFwlmZXZuY5I/aNF5l5ztRoYxB7JsB4X8Qv2gRl4kBAkB7AbHYA
m0XWHisQGWk2l1Dh00xyq7bvzVw30wBEvL63Am8ou2N7i4ZTnTXuMqSAT2gXR7gw
pkLwJTSdWC+ApFcBtEHxxsxb9pcwyIArm5sB8LCDZiW2eo0pUtQXw2aPRkRSqDFt
d2FmA/tEtEIiF7Cc+Z5cdJKAXEEBSFIv7hWIewFohHl7b3KiGjK4Oi+4B0bAScwU
MXbyMFk5NwORYxqKwH5Qe59uCqZNRfqW1jVAvGL8mYAsOfMrUBaffNAH5ShQddfw
XIzDL1Nrp2mFpopv5++ZKC54x1EFu0BeHaqwOfPkWgD81K5mhVK3ZMJAJH3nixFs
c8mE78eM9SmUI2zRr+0zkCTcBhtWhSJUgKY2/ItTZaeEdkFTC73duWaRTIgdYmlN
h8+H8Zb4Us0/eDD88Yv4CW9ef/dVtsR0WDhWtU1i+vmXKftubwyYyVDic1UEb+c7
xrg9YpWT7q6tuyCsL0mxdgyXp1earbZftyEcud6Qw/Unz0T6KBkCZ2EQoe9P1Vpw
aYsV9XllMrrkmot02sx1Vmnou68UNcOzEnQ2R4b/zT0A9cIz4RoD7JzXn+BRJJaM
IGX8FKMbUX9KiHItqR8sdZmemodnEHqXmqZRkGTuiQuNqAcmms55mQOXXSyZ1D0q
D1v8uS3UNs6eaGqGNPFR7JSvdoSvb9WVO+D8H+Nrgh/Sy4V3dTdc0cMrFzkYkwfj
4RNienM3g11aaLYVG2meP9/IIvkkQ+msnsfEIuMRS1Mgb1PfULgr15V3TqwPbStw
Tl8j1vaGvf9OwBUDatGsams6j8UDaI/9Ffl0Alr6PPlCTfKoTjxmi6H31+Cdwhtw
0D/TIMAUknEEXbwddNky/0GJM2ti0uxT+6ZIJGMhcR9Q4yL8JnwDlnth6i48Ib5E
Ur3jKJa3jx7gI+Wi/aUmJi1pQEvmgUWD55UStd098eFGeSW3wbANHeaVDck0JP9p
izLTCHkpu8hKI4ZwOGAP28gKkFa/E557UaxfXmDlj2rbwVkM/TG3PX8ZrPyq7aSL
hCSYFK27z+kYeJlajGrifIhG78kAiDVLJLHFyEtclY9fhxieL8SClqJmnkND69OQ
sSFJmGbNxuCEdeTa50AHox5DgkkLbys7CAhc+rJldgpjh0RPHXsyk9WI+Jt7iXJY
o6PlirDDtZW2MSUVxbdhmHUeLDUSuoE+M2J/8EAbl1mByKKqLKznrkbol8YuPR3f
1okcqEDpfab+lxNQP3wrRZpFr1UMYJ/Rj/94BI+4g2aux8D93W5AgHmKtAhD5/05
K1/0UwcJm4OO+e7dqQq+CUEWudjSBUnpyabJShTdM/PsCEfVGj77S7YFB/V4gOFY
ZMsvVlHwqP7Y/faFyzQmijLEWGAJE7xUj6lPKMig65gs2W0edIkVNhJyroJA0V2O
roMP7fQZ6XIPcRwiz7GI1T/wMak+a+lHk8XXZf//E4+F/NHFEpcEgAWBXzLID622
OWvzhJ6rbGbVvEvbUEaQoMJcrgbic7j/6LTI0Y0uhtdiWiTpiHd0YKXtAa70nNT9
WUX+k+vAg92M768xEWVtJHD9tiU/2qeEZIghCQc21E/sFzA4KDwDHUX77bnSEOKn
s7RS4eexzvvCQ3kjN5Lk/knOvw5ZairJspLfEd80QE6XBmlbpNCSmM0tav94peVR
GSNqp2bu+5cIDU8yAUkCp9JRBwuo7/IyB8i0tGqwl+Ev5kUTjuV8siEN2XS2G5cV
gM36NR52zOsbe15t6Qtt9JkKFXnrYfNdiIw+VWBpthfImeaFp0JNrOgbUz5wdMor
u09qB/zden2kDvP9H1o+bDwS4hLwJMzc2HZ9GYFtZDZ/Ltlw7smC6/7UL3UcGeuq
1M8q2ceF4ZwKqFTIGNiUeWHJtbunBDYHXhnmXCAdoi54mvVcCN/d4zGyriC2o2pd
ofK8o+ljG0DUByJ3RpSKVm6FRrQylUiOi2xxulGWXxShZY8a36XMNXUceDsmp/vq
q9PMbJ4bx0G9gY49ysOqzOhBvv3wjZtBgq+5fo8kAIO1TbrQC27H/tF0FNXgqbTS
4ng4bjyRYW4hgif/oqOy2Ce7rsrJN6mW3abyj5B3J9hBnsQEvBYSMlHx3KwAcl+k
wt52oOIcxhrMwesY0PC7J63crKSzZ+li5+CFmZxE6hIqT3Nav3uaNmvfBaNxDBlU
i2S5d02KJcq1hOKbT15MzkE8zU7JNt/rNwO6dhZ2E/Anv5AsCepyvxMV95tb3dW3
jEXEoUMnKhwwxEsI6NwvB787iCIJDGTgGUhj29k9qmw25OhQxcf++tD7Ys4T6wbA
oDp0dK0wy/v+Cl65WfC0qIJ6VvBwdNc3Oo4Isn7anLtHFz6hM8I4D5EpYwGtuuz1
y5AHHn3sQksK4RhTQBjN2WJZBOrw1Gw4Dy5qFUC8Tv3OwQF0yzPeh7cNQdvER9vo
eDBhXljq8eT5elX/B6HvyC74hnAcgJ0xGSStZW9GWQLJB5/M+5g5TUhLs8diG5dq
L+T9b+xV3PiHFWVy0lJBNn3b9nrlZ5Ha23z7LIqqII8pvUFdN15R0rNNYiDEJT/O
KB9fI9n3BCdtBSH+7eTxho4wuhF47js5vpubEw1g/38TCpG/x3IC4kB0X4/O9Bqp
9A08Q/ZC/jAoib3YAdh5ntfBQS8vnDl6oQIPXsMg2C8VVeoEbNQlZ2HYbPrY16/H
SJ/aG/CSci3R0fDh0CsHODDfUHaEm0Jd10YqAAloV8DIilPvQrF+ib33j/3LRpzt
2QdPRm+W27/ZtopQxisaWf2+dFgXcTxSUrL4xdkQreWmMaEBm+/Ux96Vzn5jEbAE
Fi8LzyQ23C763amCYMwHiCU+gkX0vXRPRt2LkYuOUAzKMGoSqhoVGDUdHMOiDGQt
tgyYClCsb+ZKBg1ZwI9Jq3H6Tf1i49G46wt27HxHoMprcvAm1AeKEZga1m1n0ais
VMfr9Sg1Cv+4UMepQW2tPo9n1yMoEdH2+UKoAyL2wusCk0NoEG3rmhCaBpxfJMJu
n/ke48sYOlQiHIirN1W5tQ0RyipkyT9T+6npH1pgy7ajSYzS0S784gzVceIYIUd+
CUs9umeble1LJiwbfPp4nRtUKEwHT6n91933D3P6e26cGTGSzWSS8UMejk96KMJN
/z5e312l23dRfm6k/CP0Hge+7qRb3U9zfRv1qK0Yf619/pwtp9g7Yv2yHdyRssC0
Gm8zxagwqcIhoiQNo/8vG3Pzh/p3IncFf1eYceBTJxDU4VzlSgGjIKijz0G8nWao
+SFfGUfspCe5ZXBzUdalxscpK1vwYYtsAkbTsF5ZgHMeF2N0+oX19jaUMeyUufZs
E3RYdmw89lH1BdTupZ5TXMoXED8KnJ+FTbLQbZoyhI3ko6f4SfHL1UfbJ7Whz1AT
d9WMdkW60nXDAENa4xjeOavIvAw/h//j2bZFbc889CnvAbhdHnik41b1TOCmUdWB
niwxp/f1Gqlv5NIVgApXoLbHadgKEweedd12QuTMa/yPg7vOpRJ8+DZqRHdX5Jid
tWN3iBd3U3SRC1TK2ci3dKUxCGdSGA/R2Zj+wpN8XF4bMZvbnkh3vDYZBENVeY+i
Ia8RHMKHmjW+M0HOGDe1B1JjAvQotOSpfqMHuUEcUZfc8uG1citgiU72GRRQ5ajO
bTcg79r25NQprfuka5rG2edVTA6otUl2Ril8TqvVdgVxd0QA0vz401wdHLwdrgu2
Xsfli7gfyugPK7iRQIppgK7DnuBbxk+VmUIyAy3EUjE96SKrMJOLd2OlsHSenbeY
bJJApEzKKPxCrDSGk8e/AN9MqZoiZByn2b52IzKSL2Z/c3uFtnOYPJqjzAnDA4uX
L7z8kGDnBc/ckRQc3qUz5xRO6SbCpZWMp6Ck2+ku6uqSrf32Jsup6J3Q3huqQ21O
JwANllFidLC20BPD+dndZM4gzqPugfIykMGpikKJucMW1zT/VXAkJjgCE++fXkXa
MubPHWxAWn4/wSj0vJkXKRrvsOWUjJvxp67VLDU6TniZSuZ0CmP4FFmifROaUJel
ksI5vGXt1tx6Rgj7UFrUkojIcPuH5LEbjm/RopD4YwOOE/SQQUuweqi/ZVcHpdri
yBGgD04hTQjUNjtOCYoPW8G1vGcXSp/8Q2R3/nxXRVUcWc2jQQbHueAlYCJ5UstX
g2afX1tpkXBgTITp+tQ0s+BKfP2d382f+/PhQ4CRSHGjt7kRiE8tq0q8xbikMtdI
EGrdULED7x2h1fPrxh7O4Esi32bee2Y/Ochul5LxIGOde9o6DKEGv6CP/QQ0XiSS
mohAAuFwaFMtNygjSrkj/PFPtrcplMhzYka1rl3Ca6bqAo422wWSMDSASf5jxZzx
PviftKL9sQcjzT/UrNzidGIKd47DeD1G3AUi+UOuX37n5T6v8fcZbDkhkkDw1X7z
LZRQwMtvw7orNB9LKdl9gE+bGRmBJXyxVrmh5dgT1ZPOF6+GiW2IYDPEY3Cb6V0+
8HAdCJtOjIdj4nhWvdIN5b69CCIcsVYeU+l764BepOwgYmxFtmIPzUqfDUEIUbuI
pzwl9KhsJxam0co7mx1A2ck5hr50UbE3G0vR+bBxNa7/PAvgWDlUhOyvoj78wP4Z
NJbC2yt7F8Sgx8hYC3pAOP8rg4ioxn5+ImWKAkF5hiBGqmyCUushhfKUbjWTn5nJ
MT/k7XQgHFbzx94vfUc9Mx8UgoKSD/Pq95LPKT9OnpjMHDcsO7s2RkO9CPUwpTze
VubxoXaq2AeUd5o/f/9JsnJPmpwZkSH1h4JytuWHvKCS4OeFNHsSKYHo8HxdW90X
yI3lfb4F2/D9QBQid6frJRntDStiW1TRsAIspbx01HJc0nx+v9SHSel0DDhNddun
Hmy+C3a/ctHE188YdpSrLlx6EwCMTu0Iuno5aPolZRjVgy1v9W32EQljPl0LTao2
wwyft8c5OLE4N3I2dxMUIoFCOBlu/EdsznsMWNFaE6R1gKOlCJETI5z7isHNwm+O
vggV4y6vs29DPvaBEcAZxj+6dDb9NJTvRvTrjNBV3llIXUZbt2Kuf2JI34kkA5I1
XKq07VURRCZMVc+akS3cD+wJ9yu1JM54mgoPXo+YTnbkkuBdZmsmStCcqx6Dnz6T
b0rKUni54ke07yMJt32/lPvSyM1doWV8wuJ5lONxmnvj4D5dxTC59Nf7EHdTxIWD
1bTdvg2OM25LlNWVziZ48taP+yCYQfSA9TpHMvLDB5RevxLy8XMuoob8uyGzCDCy
q7ImOE/4yQB94tcEv5JYkVat0wPl6GkwB9Una0CAwhLBYY5lfdQtUbOE6B4FVtfe
53e72+AMeC61J2YV1zUXpVA4IjnMvO9gO2/BJks+IQ5AiWarXcLaz+qlvFqhh/wM
gIolOjHhXYRChIpuG95SoGUo+ZSNWTAt+FbYUihtCIhD9OxdToF9bTqknv8M0s7e
Gcbca968E8jcUuwQ1jbk8fClMvZVDW3NQ+2uF218m9hwzuYnNGziDNtjGZsF6ZIP
OfRfk3cd9vue1yOPajXTwckf3Q635GOmVqTQgHix34Xx+EFg0LAJZhaHB8UnGV13
xI+UVTZpznO5ZoWPpMDXLAzLkQIDJYp0U6RlEgwfcmIN1fhPw0hfizOZBQknlqk8
D0vZlm3kA9rTPGPD2xHc+PJBMTs8negmyQmtlLJeo0Xj+XqKWVwCalApfz0yF/PI
DsamfKYFWGVGkNeg1xsMQB7n3T8I8BbbOksMaWAq2OpJLc62KaU8bw69DaQR3dc3
Jcvb8cNqzPAUeRHXprwEkWprhsvYN4HE6q0CRZ6COf28oN5o14ENqo06iit+c7LC
CxuN7fQNroEiJvz/bpkNJcyTfni37/1CXzRooemKUR5XuILexA3+qdOmc48KXecl
yS3CXKcYcsJMLLMDwIgFqcxr9LGOGrB+pBwgXbM5XYxKGLGOs8l417Hil3ByXh5d
z8cEm/wwEyYrF+JjtnN8JV/gZWGtvvdLEV1vVLa6SnGx3OgSdfVajtmOagOX2sOn
XE5NejAPB5NZOeffWwZLzNdIM9MZ8NbY+tltw3KuljdGleBOyBkpj5V13bWegGSq
UjY3VTq8MgWlGci9Kw7/+Epyv8HHwlVAgql3YhDq7gYrnvfgD3KL4oGoJoBXifch
k9dKAROb4cNnAjWT4XGOzNZrabAfDgxwonnSTL/4ruoL9tUMRbY4np7hIcwF5n8b
vk75EhZxizVxi4xwulHgOmtGxrlnDqCnPQRNgNzZg8bfWpY8tyn2VfNtSbOV8TWQ
rthEPTLvR+LC/JSnvn++G+yynQp8mywuc2VdA3yluRzxf/aKU0SkmTQZT/LSV1aP
Cev1i7ynk3AYUTBQU5Ex7fv6Lh1UlSvHVTlLehi5qIwaJ2ELas/bBT8HswiIlKAk
Z03ubCnUAo0DkuQjSDEva0UunUYoLfskWZijDUN/NJwoUpKnVNfEkz7KlstQ4gpx
HuWeRiSaoP/2BUxuHShgjTtj7MkR7EOfNSqD1NiaJzAPhUtWB7QPg0HLax805lqv
t8BRZ1KUvzes0wHJHLjpThZ4DHP6k2orhfQocilLy0s0xUyabUy/iYzMI2NwQbyF
kzWRq4F+s+q0Qz9LWtiZooGRJLxjR6F5TeNXmcje3QRzqBOI7lVxLpvHkgQACVVD
cSP0IlCVOZuxunontrPC42951zcxVUUCNEOPRaGWaC0JdWyQ3K5d5+CBiEjx8ymk
P1wnhCcZjp82W/I3Pdw2QlHPS/iQDJoCbljBtZsRTKZpLjMOj2jc0Z7Ae5rYpG8h
wvQvUUC6OUQto5CcG6EfAq8A6lxbYpPT+tyiEoHfYbG9Cb9mZLKWCzx8n1K+dG9t
RjOEzgDtVhABU+4ju5E+QsRoI4027grBaGj0ba2oCBWQ1hYHjw3ASPO/9CYBbzQv
zmTK3gLEH60qH4uNAVHzD8XvaiCPd0fF5Lcew5ZTDW469WR5WKvsSfoSU1jEOBLC
oClz2YUh1lrKTFDWmmQ+xNosZIq7aDAvAn2i2ghw4++wTDOZda2EKQ541I5D6gQP
pXygukGPofCwUA1AdH8Pjkn2KxULONqsVnBsSBxV1WNqwtw8iWpJE7h7ygmf650v
k8CQbGycBargYjoeNJxsO9TGjnzIkZpTBcWfT+C5I1/J4GrnOxpsmnuGhRnC5zB1
GYXE8bLrrTlaDd7DN0SH/M4/nkEK/G8RZF8p/c95ITIU4uQD+4K34c9ak0dk4x50
8whTOsvZj4ZPWIIfi7jyeJA+06TnSMJrnD8L+3OTTJoMxP9c6OujQpcnw9XD84a1
5uEs/lxNmx8GHqpL2YaLOT8TZOjLoOR6nm33lBBYaoTw8ZqhagEmIHeusnOebhg3
cjfTGf45pcXXzwCOxYiWyjIJTWbjG3Pu/J6S0IODmmYtSiy5fmD2laSct2JLA36P
kwv9tIkJCun9Dy4RdR8wzwDwmeUP9Hr/A0ZpJWcfZip1vophqbCUwFSKNmVruE39
d94jlVVoraQJfZHfiniHnFLxxAthUDXYdzYvBCDm7fDkrpD1E2n4vJmfICtP8hkt
81jRy1Zr6XEhGrFS6RdOC0R4NBOJGT6Tlh3c35Qzf8dqL6MSJj9qOcyTNOAYM08Q
XXAxRfDYzXxnXODQsLkaGzIs93ks8EPEra6KMRNzltD7KDm0kS4pDB+Ld90Fz3ag
pVN+IkKWzTXh3YzsdKl5vW37HD2TvWL71Quglvv5kd/4kSv6I7l2Ziq4J/ukLhW0
3/WBpJunqSSv6f+E3RgSEdt5Nosn5n171np50n98SB2xt8tHNuafehquS81MveGD
7KWfSnH7wWTfADWrBecIYcYOB3oo+gxKRDsL8cvie3gJhH2R8JXmFXBWAMiiY1p7
1c9a+BBHHsOHbY+wfEB/+QH+dnNobinxGAedq/f6kDrOZWxgZ4n0eNUFh66IPAek
gXzy6CATWPQF9uPNkOB99YDQ7yXAOQLrgv0Upk5bseFy1xYErUP5f5ZgEIoQb4Hx
ySTLTJXErXeCfLLrUUx+M+pRnxA+ndSRgFbVxJtBM9i/Hqh341lUVQxmwuTI/v89
+aZTxCcLLtdVtSCt9k7ORUz4fBi681j72lHjZijZWrXGOwNiavoIL1AoffOjB8PX
cFpcaAm5aLJgIIO8pOxc46rM5SRA8wTbjl5Od58Yz5yxfgS03dU/NVxesjQFCH+2
zwotPAs72dAtpftn4oPQs6C0Eltjef0wjL2t0Z72uC73yoWlZNjowMbra+HB2Vm7
CmoM/o8vE9GHpg9crxpSbxYkFEowcz+Xvk65wooi8qWtXrr3n8licA+m9QUj0Qvd
4sU+Qpmr+DaI2iKHgF2le5k6V1WNR/zk9sOhr5TNFBdM7HG//QQvw14TSCLcYzFR
3ZXyvpOVaYT/vzv3x2IN2em7Umsgj6+wUiW1sfIeKaxXmOabpPyoZjLQCkTQLDlR
8End/XfYdayJIXUoSy9qyNKXAW2+fk5w3DhQhvcsUy+SridWweP40mSsgSnYwOqD
msZXZS1rWTbhIv+EAI0Mt/nea+hg5BHcGvUrRSfc+tfpSP04V7z3FmcFLD8+Jr9l
H/mGooknL6WuDg+CFiltUEI7lDlceLmDSV3RVYMwnPxEgW6A7YIO8ot2fLI/gsSs
cRJtdA492b+0nHgeecRzfJib7uM9dpVBqns4Qurr+0cDxroOHf3P2HV/YK2KJduW
2H8sn/UdnPa7mO237pzL6ciRBuYX/JZr6GUxstTqXfdvtkB/i7KiuCobMW72tD3o
9FF52g3cTnBu84wPY5RCIpH+G605KkPy6FC86l5t1lFwIomQ4uK8lVycUKNBlWn+
OTPrYJnjIybMRYC4pKi7X6nsfJCFb/B98soQCDRwDj61FC+i5wxZhr39msSQypOA
nRhQp0xjlBytJH0yrC4ZHIZlWo6ia5WGWD3JSIZRtUU2Q8JPHOMqQWbVG8cPwtIT
rL3y9NxSsrFVcMVkOq46G7YFZoATvRQehQXZ99lSQhlEycd+QUheNQC5CMz86z5I
OXc+COfyhwmUTo2vBMrn6s1YNreZry0Lwen5ruUIn+wYnIyOjO6De0/SLAsdorBh
SA2k0Q8bdyTHKHIH0rX5LTe4wRUXxgD97SxzYCmpoNnntzpXy+w/gFxpPrHum868
WWzgPMrZgpeBWCY6TNNuqXl5dFHga1iM/ld+ToYAS9U5/NtRI91TlYPVJWRMy6Xy
MJu+p1udK6i+wceVtM3x5Zs//qfReQQb/wbQqRc7Ku9RzMg02GOj8vp1ODPYZXOs
QgFwtyHRKrsPRcPmDd6DHmJdFjwMrq5PDp0c1TCUkfh9yMqwoEXDFPfZSIilZA6I
OeBxHdsAB64pW/Op8mtCkKoA97FETfkPE1bDMgBE5goDuZThBY7GZL+ZWYR23oOi
mCuBGcIRnRsXOCR0ft7FkTUxL+jazF3tNntKb1YRMndlC16cKmTNiYjV+HuD+x6s
Dn+Xs4xoBNeLkR8O+JjPNUB7kYrhc9KIzrhyRENDPHZvFlYxC1KH0IxiRBzSxzoX
joTnNN+yfucyOuSTV2e8I4wB5WJ9v5eHCaiP8rF/jtxn8Tx0VV/kGlQ+nDvG8b8h
28EWvnbtiQPPehHZcCZ2tUO8mE3AL2Yn2rnQ6PQAnPLM2F6y5eSUt6sXiDcadzq9
/igKCwpkWU4Ljulfjws8+ouYO7ttbZgjDaPH7VM3NcpOQeFY1utbjZoJuzjJkr8y
jQGLpQXDGTFUTkWT0ALIrK51nKq/IgQGGWb3rz6iDvwHb5/3Lju6sZKJs6ShupiW
zkNkBLUj2UWi2zY/ct65Zewuv5Zq5/5wwPLiLsjk4DmIkpKHROYESfmme8u6soJq
iXfMHRGi4q1IZTVgzBk0F3R3/tR3NjleHtpjViYae4qzeLQahAEn+kQstc4liv0S
bYY925B6HpGXQepjeJsgiHtJ06A9WJtgr00I9L9O3DrKiYBnjw9s0/0WILz/McIL
yEx8nEZnsgXC7Bhmoqj2PWWHgfvlgB6LGnXDl0GfqQi3QQKkO8yQWBJVjbv6CZQX
giaAjTmYrP2d/aAtoduntAPtXOkuOFVR5FXo8YjSxCw5brYhZPAe/E3yUejBJrnZ
oQ1efess4TSWAQoWj0EIm4tq3udNjVEtKfMU3o6NQwOYFc5PvgVerOERjY91aH5P
dPxseapjEA5hO/6MeiIcssPLdAnle/MzCXge0AWl7wr9xRbomEIysg0J+H4z+QDS
LI7ysv3YC1XomMgZ99kkfIGV4IS3N+B1rnYhTeHpkJ6auda6xX5qo5r4GBkTbqKL
LmhPQz/sXESLwV5rZE2sJqHYe0WSkd2jgThwDK/6qfXYgqoa4NecvPRY94mXDATD
4ih24Ei3BX9MefJiISNnGMhASVQbmBy23Ar0YAOIdl93RgxP/aH69AzWzmzM38Ji
KfhDYs41PNcVk3fnaVRqnHgixeWqrZRR2SZLOmdgCZ4ndXiVKWN4l6NNx0oulkeM
zI3HEdRk+aZy+cKBYuwDkodYrV2IkkPkUEpKZtNXmpF07j2ASjAI8P/ug3h0fW/o
cERi78bNLpFHXDZxHJ4BXsYpd2Ik1dQN0fZxPMWXDno4fKqw7V0wOkX9aFyT0Pf5
AJS/E8C0cfZUo+5K0TcZB1FQGkJw2CD4iK8rcdLKksjWK4rtDAi/z4gAySeeM9TQ
TJZ76972S8J0fD257JS/TChLkHCAhWJ4njT1fQOxK1GOBPmD7nRZELu7lS4cKcdA
kPM5FiTWWePxzsfYCrbJ15DwRCwF5idMDQP9I0W/iXy+sNLcx4XibKckTIIChlLP
LGJzwCf3OT5WGV+jfSixrIdB/JUXB4thxO/tefk3V7Una4OdJ/tgrA6T33A1ciV6
DXLa9syyvWk9CAVSdeBjJ5A4qkC4aPTJsbGzd4tC+V8l2gdRKNQmmTVEspcpTwI4
3m52ibifO5CGDvPq2SVU+ToPhWtkKzRtTYPy2XJXwQeondan8G/gj9hOkH2Mg7oM
ND7c4z3yUiO1IIOr2s72XGuO7Az4NlhjmxL8em3f3GrKmVs7/secUxIsZ34z9g07
zJMAT08FvU+TZ+ATsWC140KWhlhEJu1OFKYbyTpuhVMhlr+ilpx/kVpo3uKjNNhF
KZH2CkSJqwwcucLCLLWXR0aOt+wES6fg6/gbW+ruMQUCAqHiIxXaYaRNFRR+ws8W
FVAwvruoPRg1vUEBie1+jpVqumZ80LCQ/kwvHHZdlKXmCtFm+mGLgaWCwKIcOZ99
s33pgE9weO6ZlA1sbme0pTTMxp0u90Ugrc2r/8Lw/0sssYCZXMNyWrPCaBQTMcLf
O0scs0k9d/703gLU+eDRsTAbitO+XBPP70txGiHic/dU4h+mq34o9G35Wxl0R0eQ
IH9OOsFWfZq68AwQE5q5H89RWyWcKSorFJfDJyt2cUtVFqOMxq8eqx7nunVyXJkl
RuIxtWUdVG60GJ17c780R5IOxyKx7uM4HyivKAAMDQYC15GOwnFrHR9/NQ9OntER
3te2tQLG72ncTTakjO5xQ+b4YKBSDv+VAm+ZkSF//UljcdI5khHiak5Z7InSPeaI
XrpjAQ+pqVxixAxeXM2MDMmX+CbZBINYwmvEp/74KqON4oXSyPvU18tsJNNCMk3L
juoK4MlLkGFLeybEJN14aWE24wLl0riywOQMbiJ1pPWCJwxF5GZvCRNF9V8HSBpK
wX7NEZpUEyLQIKZrVvshPSClqDqHWY7C4L50Zue++PWqQIxGVV24MRXw1l+BOkRA
nGa1wXJPwkFRIDr/ihICUBgdR+QXU7vCGETq9wfRIWPcxeoIpwZSwxZhPd8DBfrJ
Ucieu2JYyN6W3m7CNE0Aa3TwQejxHHrPw+AWfgILARTxXZwgB2y3QW93/CkGKAIu
Y2wqxtuF0siFWFp4lXGKXLgNJTxFCa9R12F76fqn2YhRBtCGBgYpxjZZ+qNYlVLi
WQ0t2EBUib2SCuUwFEcOvGcCQm4PU2CyASUYS/Xg+8jWu9t0uhDZiZXkShTH2/3y
fJU4brY17Oz2nNkLHZLmZRvf0D8EzZLn2mmzPHeatpvd/pvpN7YKfj5scvs8dfTO
pNllFnnNRq9R0J7ae2owLFLF5oA20JgGwtdVKgpi8q/2RPbDIbXFTGa7MP/kw7aY
grw/4rtdHKoGdQrEoru+5SuN/Al77EzSAIxv9SBieYVhMEreZXFkIgzALpp4hgZb
TRl54T+9tjLLMIJQ/syhDj8mPWwAqyXH/TCT1thyr2Uznxi/JC5purAHcPCHbk4I
lH1l20/E5SdePJ9fmMn+VnmzoAvbM+5PY6447f953BmR4QYHrmKwa671fbp7+fgF
wGYpMTsgm5YSrw3wWwTqg85wRmq8AajOMbPRYk4N/YswaCX4FaLSQ3h8jHuH7kSX
nmyTqDCSSD8yFgWluovG4qX2lTrqmqVUlm3PW5qVjrK7LCl2hv3b5KIDnyEwSrqu
RBPhXQ4q5ojZJfH8IOHPvMl5TbtbGHQI4+sp09lEP/8HIkqceYI+oIZgVt9RjgEn
XszJlzXBAIuNUOZ9Vp8SuvDF5gkfsj3MOYgUZhlcd4oIVWxshGgx57F37hDjnMrt
oOVZAnP5fKpULACMk2gXo24JqhCjER3NRgJh3sJYhKBHhx6mncK/wH30ejtAaqqH
qWqCvw5QBfiZwbYHVGc+DJFaKbVtaYAq/DCsS7/DLFrr1GRcaME/z9VARjdPaENr
f/nlPjeiFcdDxPlD5qKhTv0NHuCWTLhTV6Hz8HInIbxaL8MnVQZoBcz+0yt+n6jo
c+bi7QrlzKWTLw6hyTq8nHwBRyUYeV05zkwelfaI173spEYeR+p4S6XGd7Dyv5lO
thVJwInakloVznKRUiHLUdcaG+Fu8Pe2bQT7WhWODZkJn9NXpF9TOaH2vZHJhC8h
LslyuuNyrpewPZU4Id5YEORDxam956seDiJ9fUAC2p7TOaKolytVgrQewnMzx/Mb
tBDfCii72hoti1sucKyluL026NiqXtMypVbADamAF5NMsMO6cKIX15U0Nbgmqx0k
HiICZMy+bsURtUz6cCDpBVyfXsnGw2SyjmX8tqn3VL3CyrwUmE3ogDO2FsX7Zu/W
lvbEuwXc651F03wR+BoMUEodqVn3uUMn6SBA6yPWEA+MDxjxRj83u/Fo7jGf000F
rVYLaF+RooKSKztZN4I6FlpjU8tDU0xr3nsfIuatkXanwnS8uvHSwIoe8TYaq8wM
JxwdVinYCBI4zar4WNqR3RJn1nLmATtFYHNAH29EiC0h4chVQZ4zUGeGBF3FYO52
F3jTydGuMPqvao1Rxl7FSSSYv04dCqJpHoIwVctnal/I6rBKXC59CQIm8uEYvx0K
12o+td3KzsQh5y4O5vQWdmZm9y9b7RLwMrqer+sBHIAoKgviHOLMj+TsYHHXk1Sg
xVClRcn4i7+r8poagbjzPdM0P81RuhoOShn8WQ+N5uh3i9GnSn3dkVurQG/bcXax
X/WSTfVeOL/gy1GQYqZETqVCclhaB/gZcINoR9LPwxCSBAqGxCgUu7jpi+ybQ9aZ
L5I4iT0ncuGdIfwsvc7y8xpDeHRr5llaZeZNnF6KztwPkEUj32FcwRD6Z34vAQXT
ry4fdBt8EGlZoWO/pSk/dEQEJk0vYvWzh9UMRmJHkq+DJn+4hMu225ksF0XPl83M
cCAVLLUUDPOUuww+ZB2YJJg2d9/1U1pSIl8ldJ3pLAa3tLEdqd6ul2zFxVyJpSjp
1kkabXptmsXHe12T6LzHWqcxSRjvPMQtXVH5Wk/E7w8Ye7/UTEFw34x6KsSyC0wZ
82RolroDtw69nv1RWKe5z2w59XffZrN60OstW1dBAm998XtJwWQEiM3V3Sxm6AQF
pkj7/7lSNHICpDQ3am4+w8c49SrnPyK4mbe1u9UtMDAqOEhSHAiZTKbm6dyOBoXg
p4Ev31y3p13DBlBJj79j3keohyCskXVzaoMbzY6xtIOgqqyrnfKvwG89KRcdGXMZ
F6lYYiy1SrEYpS6VjHCwtBfaQdn02BEFfGLhU6Lxj7ER4lHcf7XECdHmILZJn8Dp
uxj4v8yRnlk9G4dE+fJtsr6UA5rQzFtZsTL31LBrEVizDl2romid0QGmotupYq3i
8iOKDBuUlNL3Tfm9r5H5Wm39EUSO2sU915S5ilwv+GiuEAG9W4LHcba8tvEszdtr
EnZ2jQV3wt1dMS5SJJIvZU1KAHKwH67ANLmzO2suuYpakfCf5rxY3woHn5uSuQOJ
fINNezkk94viAkKIyNXzw8txgcL4zxDTx7McXHyhalgCTZA5NqRaGUQBjThq+m8A
cefA/AfHQzdgG1T1N2BmkPIt9grDhOQlx784O0eTSoJXvnpjY5pPrZBkoceXeZQA
u4vmR9Gv0NFJkM7Uc3KoOUCAjJwiG/gSJEgzhQzWUglWb6fP695V/x5OHKX/CqLd
7sOc1Jd/GxwKEYZBAfMrtubKtaYW4cWFhMXa9v4Pf+vmxVOjiKdkFZ8T+4kbO30X
grnvIF9kAV/YFF2agg0BhMjMJm3an7SQT9Gdl6AzvTRuj7FMvM2YATOt7nAECeBT
jk4Rb8Il5CQ5q2QInKCeDPNjnWJB4oKrt76rsXacp3FQLZzkmcF3AVBKAcouvZXW
7XX/3LqqrQXUcHU0ngMDj+DUYDnnQt7FZZo/BXexxjYGay5WcKjfnRrHMxYG6Zme
60E8Kp+aEvEjMZ18PbhwZq4uEV5H0oydPrQcGKQoXP5wsnM5zg4Ejy05Ymi/JwpP
kY3JglFD9Djp6XiLGtRXGN5JM1+zoN+pvd1Lj8lSIEUtkRq6tCMLl7//UM0TfaiA
DuHbmKD9VtQJ1VZUP8dKAVD0H+avPn2ljBl1wU7NrxAj3EP9+Q5nDuFxUXO3ll6o
a9WXhyO7cOE2owBjeS7CwYGXS2aVn5x8g92s7DNXG5EmmkJUTDzV5glzIj3ZDaSH
mwT/u/4vl6YdzjhIVTDMhd6hL62gQZsYC+RoXlBFycEW3vKXOZ0e0AhuHiKIuEsS
roPJ/NwGoD2yBE95ocQrxpBgaf6fHnVe7lFS84h8/Cpm6UZLhP9i2Jcquacylj29
7ADZK5fu7xjzjQMeionnrWhkB9cOCWMZykIRhjwnQ+ldoHUD9FbWx4uOURIvmB0S
G4ueWCEIzw36krHgs/vtqFjjDNGuulOObxomOQ4cWx+9b9y9tSFzzdw3xIyiUkmp
QK5S5wBT5XVb3+kdy9NIHIjqlZOom7PldoRzSyOiyEwScCL26XsAhIGkK9ySLMb4
OxLgVasOoUCDIAaVojQiofvTcFY/QQXo/ASOiyBW39KdJ27BoV0MHfP2nmfeWtq0
kOo2oPFjG1G7Ru0azYxugOsBMKUUDuPYyTSI8iQN5DcwqhA0hP5BBizoj2pucaIl
R01UJ42IFdaDl6DJBsMbvbwaTEZf+HbArPNHGe9qiqg7UXMBDj6uwi04/NL6e0hh
jxqPBxySQGD4V2lff8pgL7ayY0G8PBkQCnDX469XueqhPNAkK9da+igKXARIVqRw
I4N0i3D9r2R3s66KTZiF+yFZrZkTdS4I1f8SdLAo4WNWEi5q6AXNrc1a8SRpZt2u
pspTFUPaNt0u+Vui3PVXM2yYcwZXTRRBq+9BokHHH8VV7tR4ffV68b7RBW15oFtc
Ug0TzK2gdRHCde01IxfKLyzjSR1WQ+KhgYx/225fvyJtjkIAt7kGDyNYQENgGhOR
Y2V/3PiPZelHqH3KJLKkFBAkqowF7f+xLGwhdVvjuU3gmP52LoWY8REEZ5fexk5V
RWhYdevY88Efk1iIr4+G5PhLB7KuAflBLiqcyN2DSEhqryLoIEucpQu/2uyCJ5mu
5GScTjDQsmzkzPLgbrlYoPp2zQdGog1UO9QTohQyqzJWAui9VNqdFu01AoeDVZoB
MK6jfyz6hOlwhKNo/JPENL0hONiO/c8bi55liS6PwdrgEegSQbYCt6lwPWa9MHD1
1ZUl7gRAaSZukIB7ej7XMdEP6O0e8boSiNlrdY/CXRYPvhBWAWRrGNz0Q1PyWcef
vJmZlL7CXS4ruoDQCVy/2ipnbidgVYVbesVIvYqr1UIYY6F0GsGNhmCeZjQrc5qW
4DCUFvpsD9wkX5NUPemDsOGG7EbOIA4adm9I/1pK90l7xWU8u79SBnQ+w9CD+zUg
BMil8eAuFcMhGmbqyrAQ+rKz+jVpg4eQXT6tK/DnHh0T8TMBzGcwMXqTIIMGaVMn
a7vFzglJXCKe31eqzO1BwklWIAc8N/eMoALy0Q7J5V1uMZLnr9x66YL2ZSF7CTEC
iMtrOuixhBk15njQW8pLLQCLgPBJMvdPY0cevkjQ4VtW5uWvwPA2JLTxQJkW4npj
ED30M5l3HldNvtRkIUZhMhbNJNd+dhtIOUrhVuSOQY7TuhOspuk24HcNEnB1fwei
2yOZyjUima5W3BQ0BEFIQnjDg1XIFsr+Xz/hF4vdWYuJjfLsnIdHxBE0apeyLa1Q
1x3zcBlTPgLwWhtsCE8NmJCK/snsptt1G3zNRyGNDlzw0xmYgeU/HmAwfv0/Wpkm
fLIsNy/zjywkr9AODfUZut8y6dPYEVpvt4mZJ+DLYYMnJwMqApS/pgYCn3UC0zsL
UfKpQGNtXpC5DFwKi35tDRFKfeIDUEXK5leKLJ164hi3p7Aof4tBEA/u6xp/raQ6
s44ISfPXK6lIdwY3W/29hb8MfpknMvTmit+ihNb5PWrBGEh6HQc2Ayde+v2JoGC/
kPhauJwn9s3q46/TBY7OOlSsSZEn++ro4GMLMflEofJDd25oCAZ59ZIVjItDLNPp
26o8uu4kOtL8Be8bNzs3R5lge3+UKAeyMj4R4q815ejRnq27gP4ltrQfiUPleBdh
nzFe6F4t+CqxtUgRuczrAv8hIU9kS8kN0WY932mRE3BrRYJLhw4Q0kn2IUScYFGT
w8132mJZzDt5od5i7ouIrSCQFzjOss2LGBx6OLacaQuYaKAqscmaigprswK5hU4N
UdImveRVKlP80Bv+Z6AOboe9hMYHqJaMPNDOw3KC2p4lNQkFKwx/TJlzuVJSCJmS
7zuqAeBaRz8xojo03jq737I1cS7TdlKJKDWtbBws3PDZ61TCfC31YlhXK4cBZ62w
g74xz2a73duIhCm5Z4J8dqXv38koSh/mdMQuWH6tF9o7YLscgDsRDrM1SW8ZOl1+
X0ewYS6EzUY29xcIq/uj3pQwIWHNZ2MXXn/5hAmOyd1Tkz8mukprVSmmofy+b9vQ
JMqMt3sCdKJr/tAs7gCoGkYFhxk/63MDImyZQKXpbWnzEoca16yaUjhNqilGRcEu
75w19YoaUlhtwzOI9Yc4yEd1BYXhQr119lHS85CYn0wtlHoceMY+IMwGU6GKpWvm
9cFgGjZGGR7lRkm0EkasF2hWD0cU5DTRJCEaAO/JWhYS+5AQI040LDcJG0KKRl5y
kY2c1Mb1Afj+SkP99CozTn8yU5RelizzVo5Ip3ZqdJnZcFZxVi4aPLM/aD08eSPn
CoUDikJawNTiBeekL/MeKAJQnrOeBFmQne7OVqEsPIbLMvVncVwp2e/Xuld1Cv5P
2eHt3K720q7k7lHyFZ3YMFtpfJMBQLlVdXe60Onk5VCp64aB6ByyfzNL9m7/cOlT
+A9zjoIHb8JncNT4FUyR4cjuR3coePZuwZ5rW1ZETJhvFsXxaRz11Y+1fAOUks+h
2Rujgy32WOnkd2tT3fYvZaO0ZohdIeh86ni3EkaGbpDd1aLrPFT+V/202XtJlUaT
qtjHcsY87dqlVgqFdDp4SxmZlRjppPEsKUZVQRIUfIwdQr6ReLUNUTnjCQ9LnUV/
Zb4c+4rI37gXVPfLeTARbO3tFBxf+t5FrNDY8YpilkMIJsb39efKfSCPUJAxmR+3
Dzg8vtjrhs/RYGkUSygQb6I6LSlU9mRAEb8skm3c5bsspA85ux2sc1+kM02hJttj
jvdnBNypkCcQY06SHqpEwc1i9c7Cw6J7auMNIV6uXxq323d1RuxWvQQPEz+/DaVL
mDqmfeU8/LULVb2WsthaJT7rtoAVXnCzwKE90Sylr+f2F8be/AYxcJJm9I/L52Yk
ZB1ieXr+kyQ1abh8pqKoZdbip302HQRdWnDF7SupNisNQwHauhMHLLOvdbBy7LmF
TR64oPTH7QQFA8WeKrPwFOj8ejk+Dtvv3BEdykPL7BNHTpEAZ6KlEWg180MQmje6
ZoFA327Z133/cDmgEQz2TQo7bKQcrnG0SvNPuAgDWg/RzBtiFDxf0M+ANES2njXt
Mmwo6x86/SfPWf/YNVmG43dYdDDzDhQ3nmrqxqEyUL1VWnsldcOLiJxXmORW/5ST
NB2+6Fo7UPLhGLlMWZOsxyB98zDpMlLnuceSyoZjVgVMui7zJ5HLCLxdu3MnlbwK
xMp7kXSkIdjw9yv7WkQcpnw9YKRWiFvTJToeB5eyxQg/yeZOGQ45yvgrfEdgzZqO
O9xpdso4t/V+BpTGMg49p7wLXCE2vcTOUYF4yaw+QjEeJo3Jup/LTvgm2+lRwqit
ymvXTS4gC/zyJ+rDvF9TVcwQ8TH106mdJ9ycTyW4+SNE3aAabRzk43YrtoLROEsz
qr5420ZRsvCUp+oAezAx4jG4dnuAFx37Z4Mqx2xx8GqdDTb5ydif48WpTVpIi57N
yM2CDaIZCqEcJu53opVr2Iyy3TVuex18M+u4oqvsza+q9JPyNClv0IOEstR3fCYF
I9t8XW7x6WxlbaNq4Tu5PpVH8kowb4BIaPgZ2MndjIXk8AS+9Ch5XrtUiXoWRJ2o
Ev51HXrCNgKl7bvSiRnM3ytsoCJ2g+gUskQCrwtSzTREBp4ZJs0Z1ofPVcHiU6Fl
yomW4LyLuxDgEPPtbtKQuqjKrFYjPv4VEyO9vEUTVALf2EyaOTc+yxSNGwHWdYaS
QAA8ric0tADm7hRVt6bL3YxdAq7X/p36g6IQg7VnVi3mJGhUwGM0ArCnauqA6fuS
rlyq543BWpFSMps25upA50NFOEzlUaVexozw07LHd5pNMQEzddGKMfKBDZAILO44
KQou3hw9u0rAXs/IK01aFO8QP/xVdkkg2/sO/Sma6/TZ5UWPRGl8OgADIB0hpudF
k/nI60aUpqZs7ju/xTGuGwvF2H9Dd15kOEfo1DeoBBkPfwBzW+5biIA5XlKqXXbY
+giyKhU9UO6zLYdUcaG+wZ97K9aqDm0xy5LwZxmNINJ24V1g58bugmhBalf62h/f
fCHzrW4xDSZM83rRazx9d8AYIauOd3Kl/MaYVrX7GOGQ3YHJyPhdF+clcgpf4spD
I3ThE7R7RyQ4EiW6i1F4yKzR5Ipz0xpGDsnnpG8KchsC9cL4l7Zl7famw6Hlj001
TZ4IgfIMV7mkfJGsRxu/dgZvzLPRwtKR0e7tJf422uU9ZgOUDW3dra0pfTIuT67T
VNDBcP8gosB7jV1t9bYq51wE/nQYWjHCOg6ujEMElF9bygUerPs98SB2Q1pdycsE
pEQtW7JcrOmlPSJd9F7rHcalrJnQOiUnXMOuIib6XsOAGw0pJLpATWGA5ys7Pmfh
t1Qh3UgVelo6liowp3g+MyEvZHdQuAc3exfD6FetVH0INfRUdhM272YRjfMs33ar
ip4FrXTeyl0AGoxKqKrbeHqWGTftxtrN9feiW8VuOSry/1tIdFtGt0pVCUrNI8Hf
15P1Cxrm5Bvp7Za9O+ic0V0/3uQMXwZ932wOsB0VW/8HHpPddnvt+JxFcBpHN6b2
NAVy3Z0dizJzJaw1u/0V88f8r92pAFe5J4/0VWDof9PprkhP5Mgkc+vObGjAIPf+
BBIIsSdulDWAFhgRQqgfOaKe2UMAlwQ3VGZOsyI1eAjSnjKMwvW9JJhcGt1eExGN
0hmOQA86SCSnX94eiVQKAHNhKw0g4NmwEuRFbRsDvOOjJ1FJjWbS3oSTTo+rEHOw
893pxE1sPO7GDVo/23gbGYhO6uhqyyq5F9dIDt1ts0sSnp9FUkVMrlwQEzyVG8u+
O8/z7+87XWeaDssbXJPUm670sHYdee/ll9Ib22ViTtL+xNJVV5MbQ4g+7iXUjmWG
vOUwuZ5R6alv9krEvWCOYq0bGg+p19WoJnlIsXNX9bTJz9TRHuWAu6Bfy92tYej9
pH3X5wZbWpzRBH9wI8YdAGmobAW2hULSGtQZIdaud5/kbAS4Cu0F1Ae1GMhovYuG
bIWYuVqskdd2E0lBADZvbLW32DhfaHFxHQt7ujAU9ATP9/wWFwB5ny16Ftwk83c7
NqrcQ5SNbWOk+JloFyhN8tZmFEFkT102z8I1p3u1eFz/PkMMDvIPC0Im0DtdSW0w
/SUr5mhvwBx/NSOy3POtXsP8jgkyccQ7Fu+EHfC1KTqO/QiVNlGeB7wMUXTcQ+ki
IhGUpOyWqnwtJqglnHrIVMb+sU08hhrQc7K3VcHsvxRW79l7d1jw/UJxA+ei1l4Q
/p2Teba/vwtMUf6UZCP7rtVVFlzoPU6w5Nvk0ZAjLK0838xnIeiq57JczkC394TN
u7cLQNZYFpnJA4CGVV5bl9uPJGDBuquvMKTooBDTgolQCdNrxBEB6LGm8W6Rg3ug
mhCBMMzVLuGGTt6IBzeP79bEMmm4+unrkmxRA0Me/AULdPL9dMA+t/NwQiw0YHwN
IGD49Xzcd7hUmbi0JBFBrzvDcmXyaBqgBgfpWac8il17wbc6vloB5bNvOz4LBwAU
pSkjNMCAu4jCtUssS9iIiXxXYydhzVWCQrXf5CmOqWhM+lbYrWz8LdR7llvaUb7Y
4+6ur21HD5KJ31ySVv103Cl3b4EMJvnusFUg70f5RVv4FMB1Ppx0AxFU4LmJt5sj
Q/KsSCnpOnnUVeC0qz51snio3XOs5+UDe2KCr4osfrDMHxJexr+Y4b27sdxwioiL
fRbJ7Oo5KieGCAu4Hucb7RKr5PjRAYYyws7ia46/FoP35gMZv9/3tj5E1cmv6cNg
1bOpfy2yezMf0qpm9X4McLfFKzafEuHq29+r9co4r5sLpRVgUi/0g2tnwmdSiK2N
49bJhckJqirbTMzSL8ogZOX/GeugTDHoJeB4ip8NVvbXOgdC2lbkYS6u0lQ1uUm+
6wJhbmD3vTK79ItYB7zm+/s0yJqhjJXX7cnV/h44xZZ99wg+wnaVNCgd72x+elnu
ufMWaVj5ZXqBgdpjrV5C/DK3SjbJHeaS3edPR1zd8roNJR4P6mouNIGdzh6CWBUU
izG8DSejVt0Xz0sqGZAZin4XP7z0+0IPWuJZKKwtIBOhFDLCXtc9CBXr+zfVPwTC
RaQIxtluuECfRzaXK/WBwErexo84RSN4vE+6xHFj2VLRuQxH2eQsfBUADYa17tet
2B/Xl3aFQX73rr7oV/GGXsF10XFo2d4Cx4VDThctnYSzQVqrHzbGJzvNLOL6hhhr
kI8dUP5RatJ1sEBnmYFaCTGfhPPxVG+zBPGXcVyCr4KCmgvPQdRHDFvbkeXcbCXY
Z6nnF/yyzpFNF765D5GsgxSyQKryk9J1AwSnCxUS17+aXiqmSmwax+dF4vyGSU/D
XwUQ/YBGrDqye3ytt5NEPIK+X9Xts1FU9+ZgbZo63NbYIp1L48K+CgaW2VjQDn/Q
hyC6Sj+m62URjHsqY8HSOowjyeuGqK1QIk4emltfMN0jakHH8IlmsTWmYw/PeD8I
OYIFEdXKpl0tlx5k6ludRVeNrOWlo3r3KmET4/NTPZw4HIK5ke8Ybkkv1AXijNka
FA9Mts0jb+PVYe8ARhwzhEeJOlq+7eIbgVRb/wJeSBtcQzs5aPA4INsrZNNtuANt
Q1gXQqyWBhduboL0VbhT4HsrF7d8HuPqZK39oy9lhNER39zM1D8CWAUPg/gxIYZB
6pKoGq+jv5e9IlsmIw3xASv9WoUM6GZMaYQppAp4PeQijE2SBZrkitV/U5thkLdR
FG5+9NeS9fm8eXUoHrJMtJWiJfc587C+hqTv5vWOpMi5z0D4/VsPpZzvqQ+8Y3HH
bdF2h7bB/85zHAEme/BjtNSerqkfpXfpTe70blJp0MSAW80kVElpV/51epSghmKz
nC41SnyHV3tPQpCBn+c2oJzhkTnFDfALweBlcgdnYdyWrjqoMP4UVKUXO8BODa0W
c9O6Mq/2wI3q1pOUsuNjM+z6eh6cM9ZD1suZHMWcoj5CyL0mlVR5+WKby+W4iBZD
h7XCV5YN4R8WXVCVwAPhWEHs3HSPgnKBgkVa+F39vtleUiOlUd87JAMrIkcqaEr0
oMBdxSQe29XTej4hTQnz79b0Gj3ZJwrU/1lE/j27mWby2FNmBqpGCb083xr1Nsqc
s5SuyXPW+ncXEyftPE7L8GoR4FlIcyd+aoBqLXt04IF1E9WJXVuabEy2R++saTzI
d4D7MexbixonqJEbW/1FArKxHfdoc4JnS3YXZSxockxkgwI9CnmbcRbfqpn8vOuY
xxaYlFbH4HjViZJaXEvJXVzM3ywcR583gDjW7jcBoOPtWv3Ifx0AoWwrprmht6tG
XsPH7JDHij8U4w6FErGbUWqETzh7Xt4DWfxMTPnvvVprPxb6/S4I7S8BlQe8nCUW
k2eKCZPcLBVK7hqEnjKhcJNImnz0dBc97rU0MiBksC1gPESIwJzQDrrY4gRa/7mV
jhK5YT6bfmNv6oKBoxu8fKX2Zgo1TxW2jiiD6iPxc6LC34crsFXP3tDnG37feMva
7EVKiOHbRs8PlXPJSNqXdx+ybiLk/bHR+rTwARexq8YnPFjsgX7VPsW3o2I2nch/
SXnCrDwrP5PWaQtXUoD2GBXEhlQ2hO1YQ8d18StNyJU/75GdKUqWtB+M59F7+adW
PxpL14bkkYNfbxxmM8njKGoF0Kx2Nb/v7y7K4FyiZU1oYqvMGmpWnFHanD98mF/G
AYn/b6Lq6H1Z3D8AiqOQn8s52f/vxebe4cUmQ18MstFnjoPvr1pm92JcDdDUl6FH
+1fGChQQIVVNzvHfys3TFUcUiRrX4Vnw3bhn6CuhxUu8iK6vwvY/EXr0sHshEs77
3PJvMckxpQ30GZBdU3IKi63MdiVdhfwBWpnvJU1FTgnHj9pzCHFk/eStFg5hCDUz
FndFB5jxZDEDfXwo7W+O5RuGKQe8MDZZVdeY2aY/I95XkRrdzLGHSG1V5YOfyDZJ
uTY0wewGjv0FvZJ6njpDa18llhaWG2eIYDkToI+7J0EJ4NNF0E7TuuJMt+XCknA+
cGXtSktGjd9tg15NtrmvXKKQ1AeceFXl1DycrLr6zjmpJjtZOl44wA9ruVOT0vXt
dovmL8GSW1t1ioUiLHY7zAXBhzMXdN/QkeT14LzQw5fEHtChcUjGlrcZrTnKaPOT
cfwx9+4XP2quDpFYRQ+i1SuYTrBeT+VIDIkdJW4UhK9rD2GpgJfWW+UuyIkwXAmA
lRFRkMihcx/veg66d4ANiQyisDjVSrKRMlyt151dLlG1sLUKWFM/OTZrW2+qUwQn
WtNF9Qf/Vo3RpQsGXVpbLY5H8tyiTTg8b2KVSvA2mqGEjjLpbY9vpg7ufgq5/YHP
E2mteZNLBB2zeqiGQ4RZ3CCHuxEIaFVJ6uZGvAqAqpfiiqG0YJdm2mtd0EpH0aIn
zhJ/hvuIdhnHos+CG/FhCyzD6AZ7ShM8RSohRAvgL5H7La61f4gn+fzg+xcKAy6h
SBtVYMC2toI8zElsWveQQT5BBcRdI2TyGd0qlDBOpLKiolwbbbXdiH7OyMeBv0A0
xtsF9AHLZMtCQeKtE6HtbwqnSnv+J/if9sY24tjo0vw0luZLVrbOH13AfBYc4V6P
6ZqJgq7FIWXoPqsvC2x/o4t03e4UisvB57QQ7A3PMVcs24off4Apl8ctx/rQcMax
gzS0GbS9Qdb6zA6A3QVrYZ0ZBiHcknAIXLnjSPDw6DFDZpU2NU7KYqd3GXaEYMz2
0GH5/0UXchCiYelPv32L6N9cvmgY6JT4VjWxvYdoLNj3cvop2dJ9r1J1bl5t5Imu
dgjWS6m+ZRqu9TS7B4JzcZiqgUvg7Tsj2bVEHc52YVH49dxAHQiqJRxepLk+3MjY
NSc0HFLSGDOA1BfnDrBqw1v2mxaySBICzh/XjPeB1UcdfwVBZHupXQ5SooFdSSC0
Hthmnz7UaLaZWlxIPrnn9LUIyrkSiqiDuZMbhMC2V1XRr0qolMxpbgv5GXfm8VhG
dFBoCPiKmXaO5ipH7101cIfHp48M1MXHYshIYijzlltb9M6E7idGWm12hpKey/6Y
pX4s6RhOgjLSp3XKl6hzFqWF5CU6kiebelLs92aTmhNJBoK5PP4mwXsrGsAskNe1
BRGaRezLgztfAxSCsraY+D7S/eScHbxbJIymSA8KAR0PoBZCeqZ7eA0bgc2ub6GR
TYhgP25gWbCsNURYcHL0QD/vs2VEGyOsGXlk8Bm9Wh8XPuORO17oxFsa1qhfyGcz
1npegzjiF+Pa9cWseT75l8ib8l3K+I5OlIYxROkQfdiiVN3CJlGJtvHgmaVQf5Q7
CCo6E9HhrLEdGgfJRubht5h+fJKVlKOwg+D6Bu4KdOK6QMm5yWoW9/po6JndkBED
0kxZxFCSaHxSxdVTkEZZ6krYhhFHD1DAQ4vE9Z9evqgJztbU4HT47+Q+qqxevHiD
v70BgA96mPvEQdV+qW5nnITY3QnUuY3ZBFBzsI6tsn/9Q6TpJjgC7N4fJWPdtr7d
dW8taHea9CDw7rX8CrkvkIoRA2hClnqo3jcjya8qcg7Ej6kBFpssY5j0YbppCKiz
mZzlkOxyrJGXEV78UnjRE0fHq7hv/AxUDk6CXSsTyCSWTmTLkp3IHZu1Wel1ZYBX
i1/QnkvE9TILobZyB5Xl2m9EbiTBgEslRp54WahnbO5LgUCCLAhszG81Q1RIXP6K
cCbZKWXYV5rdisTB72u8GrZbdGieNpo2fnw7SfleSZe+JHKVowsRNSEp5J7LSb8O
pj2rON/9vaWDYgxrGPTRrl1vwOqG9yC1Hgvq5xLDebk+oYg0HFauLVz37bCBOm/v
48JCzq20EwNVlk4GhEQ9wSHECDmdRlCPLUD2R1+9EYFJFpOSHPPFeICVUUHy4njZ
7yyeaBKVzvVAZwE1cM6A79PMTZdGjn8VN8d6FjY60UpDpcmf7DRYBy3+i4PqqW5v
OZU5PwcJdbobLlSjM8JsEnjT+mrifSFtniMnZ3xkMYzVCmN0SB2NyaltJpOGQxhT
/3cZ1BGr90726lCm7nM/CqyICXVzWR1QyW8yaGlcxKqkDN1PKvWM7uR+BK8LtnGl
0RChsg90ALlJU3+JaHG+12gaoAXiE7SSvnntoZ5IxMTqDZrxit2H/HOnWPQV7KBy
eMMbPGz97usORwbVeZTBghR6FcKCB1c9HSeRmWJGUe4cjGqu2rbNNnK1dNHwMPwW
J+WgPwmEcBnKoYbZp4sp74gglye8dE6R6HJq1kCApWG9m9soZA0sm9jlqUCMwnOe
7pvOexGhpe3/pbsRpd18zs72ywQyAN0ou+POmYS9oq1vKMGtaVEKjIEm7ciKLuwt
e+Ic2enUH6fRXK7paVrB1GRsYcA8tlY9gBai2frhuwi5bmV+D+oQwOvMRgBMJtoj
yH3FPqEqA+Z30XSVNJ4R84uryfX9/BBky1ok3KyIKaAM6gnE10+K4fkjSRV2h7gn
Xcsy9R1A4ZqUpgg83itBy+vNClf0n70a1RDO1Gp5PfGNgEUN8sbpG/w+lS6DVOtG
G8J7ylJdrEN2wyI4AmT28vs89oL4nzO5LiAZYQBYD53sfnsSsb/Fee3KMgMnXZK7
cWL40nm0rLJmUefDVKw8/tlIwm9ByQ8nBeTEZay/XxpIG0zYdEy8TRL6iSG/tkHT
qzvNEa8y6FcFimvMeyepz3BSECZGVu+3PUQmfCN+G08+FQxHFQKob+ZB9oyfHTen
I5yuFC8Ei9ZDUmObDfkq9X3wXbLzCIpA4ctllhX/nU0TF92JXBf2GDtDxmM/em3M
bIdLun/p6GTPvLIiAfag+C8In5dyqopnwIVXbgDcTf6HZ56Ee5rEq9D2tGxekZcD
aHcN8YuXzWbWErvvHH0UpdwF5a28rcQ/7YJ120Cp8QC4ANAg+uOkOxVMoT4kCuqH
mBhAoSsahtaB0rfaB8wPQliU2WyNZPLpSTIe/x+ROp4J8ZnI5SfATtRwdZNICTXb
AHcZELIKjDMDsVyNjosHizPffZfJmyu34gpJ4sPLTg+SIVBkHn8QJ/+vr6rKBstb
OZi/leNGPIF4GtFX8Rp76O5a/8GjMXgTEuBDKicfS0jGlMzRtLb3ZcoJ3voqhJHA
yYQpeUbqfmLVY8s6qrPxsY+ZNvrectrjKIDzGvVr1We4JPT7c6xdrScokkMQ7+16
nxC1dy9HjQVhlSdLl9p52wZOw+0RvpXrm8g3BhAOzLNp2BmEP/BKpm6dtVBrojWC
kaJmrzf7cdZBtJEEjEtNKlyS8NkSRb7O6ObCx4UNIZy23ZOAbgqiy9xm34s0SUwe
s43xJgtBpmDivqpJHf2qWb3Ctu8qXYOJ+2EKSczcdQaC47so9riPjR4t2KAPbemS
babwlx6MXfxPVy+CZDd73hxwul+0pFNlZoRRaVmXtcoSh6nscbEf+C91J3fd+GqQ
8/a6f0+swmmofdrDF+RFxuKE4bH188lovlcMpXewivIhGJXl9PK5hvcEXs+rvw5A
ceg5+KWmgvX2Mo8iTs1hovIyb2l2zIbJUEnRLTYotvVcfAWmrKdJ6qSuEf7SSZSp
o9USMjWMIzygoE+AfwJN4j4Blg/mblGdz7SllZc2DFYmwvR6yyPaoEG0NoNS1la9
f8vcMEWmOXwsPZ48U2kP3FHDyF21HkbwUrNgNcAljRKqLqgcO76Dt6+6qJU6IYV5
KTblgVswpIX3/NsiQTdmnLvIkS0udCyQLBlj3HhPgDG10BiW8K3yvRiXuvFf17co
2VAvJP3DwTsPFJX7+vvaHqAHYSkdk667CNtNyrQ2AOiZCjZLg5cNP7UBQw0PvDbQ
CM21Ury3Q03VLeTs17T3FA/q1amygjQTOYhJmMr2vSc2exvILaLzK0ozaOy+TI8L
M7IEPWUGz3KX7/edk3wwxL3VKm23tnTeRjV7zNa2S0KQW/AOK8+t/vWZLqT11qpL
yAHzU5HB0TAY0PtBNrotz+3A4PKizT1o5RRsFQeFsa6Vj9duGDxjWFMPRbwfWG4Z
XkyiTmiUDwNW1vXgezumLFreO4BZHfaHv/7VUam5IX5t77JpvQ3fYtt89+OSzRBK
n9OUAchBmzkFeDlNwDb2gg+PAVpquwO7HQNThXAr4Tg7b9ZDIJG79FgaxcyRY7mw
07xC7wvl4sR7Bt3rzI/7lzne7cMLXwM0hIUX4Ra/MokR89K1JbYOhXnTR8gJN/32
hRthMYwWxO6+1MWtIfkUp3w1h1cIYFOv/6c34CB49U/KpCxMCja46oUrVFzMLgwS
xYSQ2q5lEhvOIp/MpHS+3TB7c/Q7KSOX51w/e0B9FNWYjTagBKblqA6vESc1G0VX
4pYPVRKH/5HXhlx8xMnqUN0pfQ1vw/No4nHFajeLHSz7WFGKumUjS+3YUQIcUFmx
vOvy52x/uHa25daOJdr038BlXmwLyCCu7tIJWljqJvo+mcw4R7BnGzkhDuhp20G7
FtfTI9BwJip/i7FOkKgZM/rSjDGb3bTtoH7pRQCpyZTR1iXiaGpNM5Ht2/jf1qzf
dn4Rv743Fb+VLRdT6IFeGXu3xKcQO2leOzg1T19k6GUfa36fWlqZO74+5J1f0J4u
rV1yYFbACgehH75fCcJLpFvVytwR7/BVm6IWkvT+zE4iaSa8GxbxEnnJR1qVOMuT
71FHG4E74AZg4SLFbJKwjh9yrDrBVKdDSkeLHQWVxMWtTfdIFigPiaj2HRIor5MC
Ke8IRH/lFXreUdzEDEv1YN1tiy5eBVINQ/fV34ge8gV2rygJ7Ik3t7tbXefpwkHk
f5QMIvUKT0JwBW3/pzxFn8u3ERYmMr5+cfYPEQjzq+/PAUer9nwgkhlM+gWVGPqF
i06BmYgYOkMh4h+INDXUefK2l3DWQ3rLMZTFkIi8ZgQ5WW8+1u9V9o0c9fxoAiwD
IPsGG5/yF1H4GmiZEKjAq0DxOAg+mh4iDStntRSCzxvGgCfG0kLz4MXTaRCCzGKA
nrSkTt9uPone39Z7VjLnyexoL10d3hCiVlRnqXGpZoTY39cskVJKAxIZMaBVsuG9
+JiTs3iPBOlI3ZCgP7UWB8Gt8X9Lab7dXsl6OhlutdBcMi746GONqGCKGAKqgyri
uOKQpdji1EQZzg3lHloJ1lemIdTUPFEp/YWFuypP5EEQWuH6ALwM3UB4A+BN1+qE
+7TyNiCV5681Qr7nO+7jPJPyqA949iQJNPOxkpVNwZ6zVGruoeEy0V0a/0rvbf37
9TzByLy/GruvPhFtkoFYU1eC7ZbuDM/4mRRpcu+6dL7+3HDNrqlgoyW56dzjMOng
Rzrcgb3iD45j5u3P96pht+Z4GgoJTK29MOwHRlolMzIrvSR3P1YHZ5s5LEhVOrfj
8EkoLg0hk0R2MicIMt8SrffhVIHAqDTR3YgDzLg2sfGSJeI8rVJ0Hw/gywheDToF
cMSBlOh0KUUXifCMDEI/hIvf9RBEhlla+cZmf+rwAU3sjaxqPB85HGjHsJZUbXnf
uOYe7A9rC3kR8oNefzRpvwOuF3TWlXtSSfK2NK5Gxc9JihUNDRI2dhenGCP/ml8r
sb/YadsOpIDBqH/rl/cjq3Lu3lKo3OmI0SMXApfoPOBvjRzANp6J/DVJwZvcd6fn
iIRjtoFqaHp0IbnDeIf16qXvygcf0QL6FhnYuUrUiS4YxaIfhGuvZmBbFPgXztW1
SMGCStdIJ0H9ffRX2x7YhZZrzVAXUWNCs75VvqWAN7H2WDtbAEj6IKysVDygL0Xp
48Jhsc7r+HaoBCnqsVd20bgvfagDpl0v1htiMAgSI+u4wNGTtLDfgh6Q2sgjPP8+
yXkYquW/sza/fGKzqpKDCL548gEs+OCYBMJ1hU+vxCEId3TjB8nxw6qSVfh9SSn/
hVj5QZtDJkm69mtoTCYEeVP8k0102mlhnpx8xPn+3qNe8d0hopjCBjdN1EI+1bs0
YeGC83dsAl4Vtx3tbdlKox3uGTEKJYx6fkd/EOShkhoTchSQRYEBrNU/kEOpsz9/
m9opBALHdM/1ar9UWU/TF/ciut326TNmyhlzBGI/XBVNRwJtYf8XjafyVHoyOrQR
Dz74C7d35vazp2yQBBF3HH6GqfgL8USpmiOyMMR2FA0JMrlsUjMGHlAKEh1oBX+u
5x8y3gopHiKj14x+/RCqdIoPzRRhGkc+Z+fwGNL1usmlPgF8iPspDtdNGRwfDk6c
Qc/qJM9nTk50U+tkm7in92KbSa6BQdpq3LOkcuEOc/UUlrXurvaZ//D/gD+oX1RW
oELb87uLCTdMliv5Ntlvn/rRmeIH0oVu/VbMyj/gTp9lWvSV6Y+RgwRKki8n+jkh
fGCBG9SEn33CdLi36I/gZjOqmMEE6ym6btdijIvP40QlbhyrJSMgE7yyuonjZeby
ALkgImDkFo9LdN5+uV58MTArMtGvX4wwXSsWDGg8dgM2rBHOPBvR1iG6/DuvOXmo
SIdU71AW+UABZTdq7wWHoVey2xUtnzWYq1XvaCeMSbQEjfo/0Sgx1neTzF1vfjpq
tCTYcgBU2oYOV1MJ0qR7xjxLoqLGomfeaPsAH1TdXUSBgPKgRHsDwKXVsfyJia5Y
3ZHah9m0ywHNgV8S8k4EWOrlG6NVzmPCPOsdUI4d1t+dvyKD79k4u9e4tO2/McQQ
407jhG5XqO++VG3eyyEZgnZbZ0meufv5/CBm81ULK+VvcWvpHcINOQ2PaAM63JAS
0rGdYm5OzApdeXPj8kn7xtCrEoN0pSdPh4YQEvn1Q3yopq01RWf08FUnGBcJ8rK9
NSOK4ZGWc0xmqaxZm24P7IU2rj/4F00Yppv3sTD3neopSaz66KIlgKxG8IEcTgBM
QZ2x7va0U94fJ9eOawlxrv1o8oJZOioi4XGGoIuac6qFMRBQbyjppD55gKd7XA3u
FvGmTRPAWAkPHw6Lk7ZdGyoKBqzuMJ4mtm82WGeoOxrXaZXQzbYJ3hOH3ylHiegy
DRxYM6wf9Vz/QTnEEl3DxxbspyW/IpG4ppJAhSGUnY1Ps6B/8NrqwumOI7RVCI1o
5ev8rfRU/E6BFgejtBWxInmlSTpJlXs5sLEm20hJDFa6eji6AZ7S0OcGBzgPUgT1
t2JzhNBLPy3MQbOXkFzwNY7rOgDDU9OHIe0GiUxrI50p9fOT7s86sN88Nx1FrAbJ
zAE30BzD5E0aZnl6jcnSG4CeBJH4j3htrzKvzyLhdYqOwu/qW81vwbfX1QV4tPCv
He9DTe6MQUe+oVHAflL82fwkqE6MJbdGfzjUY4wFtmeqiy0fpw3FqGEdMnxbQMV6
mST+6VHB+kJmO9m+UME3jVbcjYseT17MWoIGRuUjpUJCJ9oKKK9+i94tidoBFwML
Vodu0cMGfqOJVEbKXsFiolvUeknN9A0PMFbkYlt0ePF2lXTwwMv30PEdhOoORKuz
U1z8mQqMTwEeaE0VjmQ2X5cPxvzisQQayJwaydnHNdrsw0gQGsHsbQmpZ13IvXz6
TehzZX+eXceX+ikpOmZcB32OFdlVHlYfaO88Y8JmqrFwTNE6gLoBhs1qJbA5pMp4
PxeAYJDZBcDejrqnQXS1QNAUv0eXbJJJe789DIztqcZogsY7jg/7ihbXuE/EiF9v
8mRR8fuBvs2w4sQ9lb0S18oNbz5J9y5Og2sxzopqQZuc0AYrKA5so7dgQErd6cww
AgwaZeoPVAtOpJkydRGiWwaS/Y6n5sgLPBZR6aXE8+UCoFBCFv7JDHNseABRPL0v
Fbu7lDSRwR0l7pGUPC/Y5ETuEu5t7iMQWUPL+6v2JKN+9lgSPubEiaFPU9CCe6pw
ZgK8mIdOrUvWipoLH4B3tO6cgrWWkKRGS2d1+1F+BoH0SuA1DO3Jc71J9AMIVYN8
MN46dw3UpkcKeUnAdcuWhjfgGRiUHDaqRB43gRpijdeTsksCNVS3f+4Wp3fuyRY/
UCnTRT3+ZGbYNe2ksalsgBqi4DSgJiD9K2TWceEUUGS0FFgRZpS5PajoU+kUt2jE
e50rA2IOQnB+nZKDdrM/y7ErK5oxl9g8KcUuKrJYznwkKdKb7MEgeVlem1zm8Hlb
hrXz8rec9gdMM5ObBg21WciNC/9mGflp1HjmcmEAco5y395BBbsZmwhlbrZZQwDt
pzvBDue3pBtpghxNzrrSmNBq/4NS4aBS9bA4/KnxzllxLuYhy1ZADL9GSbdYLlrm
sYOp/E1qTynN/rH8KKtq+FZXsaTuKjHRs12K3j2tOOwSyvO7+1dw7ApTfHLkA+SB
uganesmIiLyBaVBBxKg2wwiJNBCwRwOwyDKp7Ajej1ypl/ijHVO/dzqs+W8gencc
PTV/31lkgN2WmCL7UmCVtantA6HrZAEMpEAkJcQgLptilH4ixAkc4W8i3BNXFL7I
c/tYmLH42HqTnKMAnB32leBdCMpy1nn4I+pwbVqXlAOEVfbkVI7afaBmy10F3D+B
A8CV7B0MFxE/aKOZaC7w/VHXjWYGueIDpRhiUR9ofLPVRiO/phw5vAc0oolfMERo
VPu98RwJ+/rXrKTpV4HpJGf4J99KYFr+m47CrVL+pG+czFFz0LdTsoU1go3SxA1q
PKJEymTRuba+KwwmWOuiQ+y2iZ5kNluJE36rhZItmNFw97LXiV3spbZSefrPl11j
fa0fOS6P8XRhU2G7130EWXhEARxC9uDNLDDGXAqr8SSibIqZUcnOAAlJVN23I58a
jwl/TqBm3AVl1Kg0STuqHB547KrUyj2CO6FbBG/91FAV2aTYtlIQReu8nYA4Qggv
1NqLjw8vQTOWCiRpJb+n1gVeJskEDaJJE75T9Z83vM/9cwZhlGTS8oeX7uflEEB6
gQmA7bjP16fKSjiFqGytX2PIWZDyfxkTSuWoqKDuVGWmFeJA/sqFApWB78OeXhEF
WmcjDrzF+HVa9YwFpg9lHakCFcKm7fCbtUtkw/XTdtrUX8Yy0q0f210byX7nGtiz
FIa0Rk0h5OZguqw1i90R3nTgE/F2N7ROzVF3c11p1QUq0Vrl6VhzNqXdA/OSN8Ls
OKr1fgQK+XIrM0O1Ta63+IZwpf50PnPEwH5oVKPTDBu4anlb3MyIoz2ChSZt3G84
KkSksw+re+8Qk9ebdgNf7uVg60w5Y8lD09SLvO0BBXoX+gmy3WuIYE5BsX863jK6
Wnmn+LfLqmDEp0j3KiLjakDX+vVqZE17sjt4BUu+RmtJf1CpyFkKisiBFZRyHx3H
1QzME5jKIgfu2eUWDwuroM2NlSHiwgZLHZA5QHryXfzsosl3kr37s4XetwwiHA73
EeAO/+wu9XIkBNA8FC6tKvsJGcmi+Nj8a0n11KoUYUbdoqSLA3VpxWS8vWfY5lWQ
etn2mWnAnWTEoJIpwC0WwgKNjrxhK/o7onImQeKKSZoKYGCPcM/B+MyEXiiW8C9g
Km0LelkcbTN5tkzf+h3/nTL8ZPlLi8HR1L7hKQV+jSKbpCIcPLlJq6Lq6TxIeaiz
GXQbF2nnS67zbQ3WXXtYUUtrollBzHlzBdjNK/GQ+ZF8Dadoh6FIt1AaZUQqbdPV
iwgHuNKHCTklmrg5oFiHqQzmVaXmC/5ojIYXeQYgTLB/SbAZYBMUrzgj/t0zpnzB
Dw0uTQQMros3G+VRt+UOAjl3L2ZJL55b6VlMPBF1vRXPPGZJpl0xVGDAWRk9COzy
3PC1YDKDJOu6NWJ2KBGWNk8idoXZi0o3y+7xLGuBd8WQTStoPSRlLtHXZZo8sjFL
Vwy38G5fnrTIPdgfRny1tcD2bXg/FVQ0BF3ug1KdUKxsH+8p9WC/g9WWxzFzJQj2
6R4rz5Sbr2GCynyXSH9/pGkx3zM7btsr2AEr8OFjKIljvVf9/UJa8x5p3d6YLtf3
XbUDGKwVhMNijUd6h0WNsuAXEDL86ZhK/+N4BESFesMUhrFb2adTixasROu4RbyS
Wa3pzgtHWIseDrveNRlwmiYndLM2YPBJPKy13JhVe5qpCH4EfV3sd6jFThgLeIW1
UYtM4YGNL4l170mXHvpLRppopLT5+X+dU+IstHVUgjwSiK9xOxoHJQCpX0VFrmd/
r915BaAq0ndPkVdOZvBEvD7EZL9fEXteBbMNuLjufDwwnd9PDys2pHLsypmsvBQU
UKPhlVsNQ6SK8TJSBIyM+dnJ6ePhcu8kso3U5tz/rrpREePRoz+EbTSIQBah+ZSy
3YkICeUOJYYg8zuC2N8XRGlXMjTD5boQAsg4zNnjrx8IIgZSZQBo/IRbITqn7+V6
jRWL3ZhgBcbTmqyVQCpcj8Fnfxeu9S9R+X6IHc+VuPqZR/SzncI6X8MQrzpHQX6/
riJRQ0ufLxlpxaTdwkCqMqmrRCaOXFMFZBqRiVOaOqJ9WPEGwm1lOe0VOjdFHkor
mlIp5G53znBXCdTC/rDxNTwkPVmqWdcR4cB5ucv7FE8pOS9zSpgPHpvyWcrr41gY
Lcpqddg6GJkzcHQ972DkWjwCQt2KTRc1wbAKuCKs4zaxCWgwlUxEuR/Wt/y0JS9n
mpzbHCMbyU+pPuxqGYsIN0nGgVi1I15x7jmfQAPp+Y/XfwzWaL4XpnZeRpjtDiDH
XTgt0PH679ML2ljbwXL5FfvLB2eJk7V4zL5cQgwXmn9SSA/8257LQHa2u4yamksN
6qUUJzzF7CfhUDAeXhRBDCPW0vc7VXmHQCGjzTgC9O9Qh1HFCfMWijQ9m3X0xM2n
AFqV/HaRGaH8ZjDvnPHiFoV8gwy5D33U/OcJp8jUZhcEzQcARIGjsRBBdbf7VSPc
iMffwJ8rk/sOAiYW3ql+e/gysX004QxRcMcrJGB8L2eUqXWeC+xzvkmgHVzpSiM1
dDkjGPdLSRfiytMfShCCw7J0rJBpQkBR1tg96+77BBxODoMN7d/eed+roPVYiqCd
ZBVWgOuTwkmp+E5aWuFz4XxZTFfDZR3DGEy8bqKWfeWGbv+cZja74X4D3D6GJuNC
nfCep2tkmMUKP8dAmGkYM3aEWut2cHIx2doRcxSloLcxUZhD1JZcrxrtdOZvNzoD
Wc8Y1m2FuNTccBrE0GNk709N7XwF3uZHjYk8fxxMYMs4gWtumj2k5RkTk+JbVZlm
rNwcq9NxeqHZiAOIToe2SOn6wwowJPEJoLlx726xULXGMD+IXfOnO9oqFCJQyVf+
s1i8P9ZAFKhbXVy34C89/WeAza0mfG/2DS77NARMogqq7Ifh2OEzJLgMzvTJjM6u
HditBnu7olHE+A8CjHGqHepFodNIpd2F4LUge3MGqvUngz9n9EBAHYc9SL19Ceem
CmvLIrktr0MWCFTA5+89mHpU8Eo8pLdh1ez4GCKLlXRy/fQTXXRUllCgAiJqIVnT
zJgBlnhulZBt0VEzJEtgcKdDzxCGcZoxgzT955vF/a0cqVthkKy02jj5VtkWlYpw
PCWUFsn0zqfsFVIeZIu9+WAAZs0OBojqO6VbkbbgWkoYM4TcByCj6VFYzXjPLQbw
eXIf4TfQZeB7txk++8AYy3/cOFQ7omsk2qN0tI+XCogeyTozWz0H2EzCrMTMSyGp
j+qLUhHPRHc8ayttszo9m/S0Fg1D3DI0Tfrh2oWiirKsWjSkmOLgQ9FKvNmb4dQb
jSz7ub0/m3T4QtnjaJCVvJNivY7j8iOWd8yi+t0DdbL+7fEax4dzBhcCNM0AleLH
uPcz0Vlb/KDm5ochCXAdpvpPXuUEUyEgWhWC4TZ8c0BHAnBiUbiSJFhSxAhhjRXN
UpGalha9wjySmaZHlbE3F5Z7FmhfY9rtapVW8pbxGEXuvfvRiNGrQz9Ab4vOdTM9
zpEP5UHQIV9siYktCCLZtYTxVgXFwqJzXmRKds49S9VC27ZJv0+6Y6Ve8++1yfYl
RuYBjl7CT1MMe+9iWjb3jVAiNPvPDnE2pD02RYFO8dDFvQUFAK7VLZe3BjSKNYaQ
BPnKQEShCAMQ4yk+cfSYkdSMZtl/5tU2/ajTAqY1n1Pha0ey772D+V+eqLfDWfcf
WTh25UrFDEackymCOlmbuyUS6+RLHXYcShZP/PFsWPYOJJl6evs1bYSNHKZHIygp
jxzWzJ88uDVpwTV0zHuT5zbwUVNadxV/BI0zmXEhsPn1XbcLHhE6rMJCzv1C8Hzl
roQTv4nik43Xbzkr5m5hg74APppFOkCxOR1IT5RypHOKVLarO53G1yYYpozbhoaC
jvXmIch5B3ID1o0iNk4BHNepXfXEfGpzTuQpK48myI9Mgjx2IBZc67KwmhOMVojw
YPdLVlWJH1xnL3zSb3tiMdSaeIgzbBwplTDyy9Vj1qjojsk2kRJpGU6QquJze4hH
wf0Iz21gyZ0xA/PuFIL2vCHySpuHgDScbbI5z3ukd5hOXxHOr6/Jk6jDgebjWqiE
5fs1CWsOc7V10nY2qhN1QsAT/8QX9CIjQox0lhul34Y1/OfBeMKYuxcqJ9I3Wce/
+NL/ChrCESwi0piZpxRph6Ue8D+Lvo3GbY2X8CHFUAcYO/aOPV2P7GO4WkHyiChb
8FhrZGDFicN6T4C0Ra+Mmf/bl5TKYaPpRmfgeCqa0nnHope71aqoOfs112SCcbF6
wg+9nn/lj+cMOWBtSgRscFXa7GKx7w6l6BZdqrgsivVYmLLudnowpjl9hMdS9Pc7
pT2h/MV/LxhepT+am1JXAy941Foh1dJlC2EO8O+Q6PmnnQNguEEtldz4x4Ig+dAp
Wif9qAQTlkit/3TsWpO35iclVzAVtZWUNSIMscXwtVm0ZFT8Qu7ECSXEIuBeYswg
wuoUVvlYa105rPvlhuC++/ijyvZyzpgQ39e8EXCpLz2Ensb7okUWxGEjUZpriwli
dzWyMN0o2+2xE8FZD716IGrqPTe3HAT9CpM+FDEz2FnqqIBVcx+vjtESzOS4ebY0
7uUaeY7QvSFnkq08/1I94L2eUGHdazIlZThwEpLb8RytFvzuY+V3c6zA/HSSBcZV
hCA8/+eYCxgtAlsDb/eBjhBmKe9kMAYpBr+yJC80iTMvsGGcD4ppsrd9eay0gDw2
rdDfbTFDnpIpe5usy72o8zECtwwL0AZAJ0ANRARoWRd/U9QvuWSHxo6Yo9tZ8Rn9
jRoyDBl803KVqleuJHtrqjmdbFLCvEQNO9pE294jIE2waoXf3i9Q+aluhZcAmYvB
tRZtO60oF/6Z79PR+xWTNObBlMWRyLMEtBEsAf8tWklE68pQSNbcFR9yQMB0zSPY
L/mQDuRTE2Rk/8DM8TQhdvkqg8Rv/ugSWee/AIFF54fhOpB/nALf2pc15rCbpcHk
Vre+zru8ekbzuQ3yJBAG1ggO8+wbWVcwXe797aAH3ztgV3xuC1x3Y3H1vcI7qsgU
ZHM2igsEqIZVMrYCBz0OzeC4YnsNcnL/k6KA962GwGSmOj8OYKMN6DOFldNB0aGG
yOC9UlSIXQh74Ec2ECyAySMV8VdYaIYgjtOoVREd1VbdEKlSOct7wGmeNfl5Ju4I
CbKzfNjBOThcVUunfF+kf4JpExLKqczi5Ux4hnfD3Zd6oY2LdBy9xknkg8RKnJXu
32n1IeFdJsAVHpElbpdw5rPidx6gJAS3x/QGcAPQtF5WLwA/iuOfIf8IGi80x1/r
vFjm7vqky0lzFVAcsr5Tn6BPhjv0d9zBrrfgj/tfZS4MiSayPZoZx96TjgURdTEc
bDFYo7OStfbRuv9boH9YLW+WK6UoWOTp5fuA53UkuXmwDeV9q5iC+jLhkuRgm6Pk
aM4aqYmkxRw5DEX8Hug+cYcPTJYrenW4BWrzOqV1brTGa0qeH+rY+/11pED+DC/B
Z/33I5+5awAK8IRPkVlPjwVh+69252blKYQoY0RE29NB7jja83r+C0F7aMUB0WpY
R10z+29xJOGPaaLzdp/Djel+6VEqjJu5yH+VIKGoZCaO+Ae3ILJSHYaMOJw8G/04
gygwf8Qohfa8HIXJU9giVdc399FuHrpY1g9Fo6cIhxN2bcW93vL4bDSCTjW9P7fl
SzInfeEBcCI81X5zzY99QZdkiGW918gXKyLxrQF5R/FMvMpdFY6B/QBCL2Ig/+nY
gbRbynkr3Rbn9e2HU2xYFElCtT9kF5Ub/Nts0dnl58Yrpq9fSEqmbAqyJ0gOV8PK
l+BEQEWzicrlI9kjBesuqf/zfWcuZMTQeD4HPU7fuil+TRshKF4z5MgCTYfx0buf
nVVLZSf8Wbdne8wP8lquC2CQ3T+FdjwkTJ5YWMQYzdm/AM6lbCLQtBsv83zsnisQ
71oBmuu04qsI0BB3oOyxfcj+snZPybZ+yIAOOmPP95kmI4coUz5Q3sO0DOqyXDIp
vk0CjCN78bs8KlYqmvnTmIRc6JDSZ7Q7ekyl76fYr6qNFYad1CnZ46JhJf9AwpBY
JZDUVefY90Oqv410TltY2pyDwJzMluzJ6FuOiu/O7Rm8cJbeVxDSxaIvtIGTluYw
bgNZDAle4iSQxGXlWhbceadYnFvvNL1gMG4UXoIo1S+7AFjUCNQI8keCnLYNDSIn
+5lnn42XmkEz2cR8noIOXk5JGtUvkySYRqzJ4nR5y30ODbdXZsIzykJHxBa95ve3
tHOXvKIuwG8BO4H4IzC0QOGmd5Ejbj5q6K5WF9T5sGp8lVFLhFV5Dn+rflpdsfaN
KGrZzSlGGFV9mUSmtlWLYkVFxKA0wPdJ9Whb0kZaMjGmAijy+J3MEkdTnsQ6U2MY
5zvsck3D2KIKvTM8v16lVyMQwjdZROdRZiISpjqQTXo2jx43/taLqygSA6GuCpKL
kGKAfienxfTFunpbwKEOtYotbsermO7wrZJqcV+oCzeJ7o30hmqgHf+FHiSKO8yc
f1dS4Agir1HhY2W7Q4WGB6EP2WNGGJqbXg95bV1L7C6hyRmRUjOHL3saS3gVepTU
wFKAdsZyJra8QEkTgnMprHcHav6RejUJzy9+wC9AcmQ0Rc3KpnHN0Bek09Cxw/ss
qTSnDq5LEJiJkf33VfcGcJWrHe6uS1AxNC4CrxCdJZKSIIyXWtjXtOwqW+D+8tgK
zT/+PCg8SzIZLxDUyjquO5+hNUuIonLv2W7H6AGwG75UL8NhabF0mfTL2BY/elBA
Oioa3406cog0kcIda+7tsraCjNRG0ogEVtu0vtBLHL6z3slOwD0O3uJOMWYCcKVN
I0+trRbbuiMTO7CEF3jPwEpExZcyja47EweAxjhwkHVkFLN9T9eRPYw+aRns81DA
531gf7uBjjN/AZedHgLSavNx66nilydPUhoPm9gFdkOlY/FKbEnzxevXxwuvTREs
7WcJYJw/U76oWgO60SgVRDC/j38uTzPgt/xDRaw/xKB1VhUsjCZKWE+UtRQGv6QX
zvdFQbGE45o4l4vpx+sv3x2ENkhWj6hoRgF3AejuSV3FQsPF4NvIhxEWx/Sez7GO
sKxbtm+QoZgd7/qHkml1O2tCwkLtAkrfSNG6FpumRq3dl7yzufhBZwJFcUnI+2wG
vXj4yWXkCeHF1HvUzIaQ0eXjcZ6r6SAV4GerI2IQILE/7SrFS8XTQ49lIz2Ny88F
4EN+5mALVnIOJfMnl4TvTgpjwYyaGAqrZsAjluNf41iFCqOZOLOMiFscoPkDsoNj
l1k1VqBJK5COk1uQp/IqO6OOZ69y5jltFyXLpPV6PpoDRl3JuRZd4As+/0/s5yDh
ZDc9B1eR193+XZjQu3+2IKgQvC3iUflW/Wqbp4jANvYW9LpOVghqQVeRHqg5ncGX
1XcMpM0kK0o6ojDbuQa6Vm5XFWKnU/5IbXSyiYvrjg8ba90fFrLElsR5iBFkAfkU
O6RTWdQvcSKNRnvQke5tSLxZabLgL9MfF31YDk3ZXTel2ubGtcAR9CDt+fcdytEa
ZpD/+YxXinuRWof0LOFDXFyFSDBhus8dZquy6jHZztRAA0Nl83/EHbeNSVKtmT8G
eFpMRaGGT5ovh51taaOXOyyo2rZGaqS5Iz2OuEHKCMLOjZ35RSyo5S/k+kTx5wTr
verI5NA49zz2bdi8KysEqraqi2ovLaVlVLoTJ5AiQyiDuW7gJ/f3jywj+A3OtHsf
hHazUWV6hncnuSvgRRNQ4c3IQhMAjwvkH/+uE3zZzBZ864sE2cPYnjMilUQsL7dS
pgqUhwGYxlQVwU7C6M0H52dLYxjhFqFhZbD+zKEteFo+bzqXaEiJeJteEe30c5A5
HA3tCqeRD8cdbYTDrQZLLj9tjKHK2yZl1gav39R5aeoYTeJIFo2PvJBmnhjlrQ2B
f3LfMEjUritgTPCAmj9BPLy1pKSQ6CwLo0oGGMDJKuVe6auW86QQMzbTLt4O8KoM
VeAuS78fgUBf1YG3KONlyhVRxOV36sxxA+3VlrPhYeSyBNY2Kp0aW2RwvEuIkUWk
K2chgdmqJCX1HeHVQCCO4D3oHqXfghmpVOzyiyijEbBCL38Q0oNuCGB6IC8JDBH0
JW5IwAHehkyNiLzoN4Obibn/IHMeqZ7EpC3sFfP1zeNGPTrnFuaV8Q1XNyCw2zlO
2ZAYclSTpZzg7Z3rG4cheygnFkSPe3h+Rm+ybs+lZ05JucKyjw2EbiRs63YW11TS
Al4xGK9KkL6Zxk8k9M9H58G6UB9jKK4jXvMLOT+HzuvRauJJPQ6J2Hz2pcYnFszi
1YUTGqec+wSwfbqfHZyBI78sCUb80/hQhWBpiZdiLUYt0PPKuAR+XJdhuiCSkbdF
Vln8aXQCMstjIYqQK2I5Dm7w4ctmRL7Ioz5JGmjSb/0NV5TVKu0u0iWx2ewK77yE
ZGGVHrdUpuLdR5IdQ/EHbZ1KqTAnlbPe0UvMTHqkSvU+SE0Hodmuaaf8z4WQ9ydh
JDJiHiUZV4qjbjgX2IPjMcPLi9fgZWjrsDbZ/Z0l1iNNSBjC493jpNiYc/mcraOS
nHNJ2WPYcRwdW9rT5tnt0WR63hjeQQEPAKls8dZKnuqtgTJR3c02qeZL/kotP+9s
G53olJ1DHdZ/Uwr3oPmduJlI3nuJkgx0Vdm4VEzkcTUClVciyEHuNV4SZGS0VZT0
J6UmTSvynTEAG81YnYYmn39pk75Y1EdZuJHlHOVzM5ZHRdeGU0V4N5XmHmB4xTVE
t9kgg8l+WMhwo5b0oXCVYUK3uqmKOd4C4eHMAsg/y+sShU6DAGCJo7TvLN5EslOy
9/33lsPp4hpy1zno6S7Z+mubSz91izplHVZJK1M+4Y9IWYrtINLrIYF1I7Rswxlr
kPCP13bQ9VhkNvdiL1P7qmidzQmrsQoMac0f1JmZc3a8obioTpkzFXti9O8cU+hN
xfOhF1/h2bSv+G0s/GgZVg7tSZt7FK6G8fg5GUScyoa29n04v1mIgWTr9TxMrrQ4
VyhP5rfbXmIuFrhLUcb9GU6BtagGGQ4lCB4obkymxjVTZqi2XjGccUnSKLHeYriC
AC6RHRjKLxYcZRrkncPfGP9y4UGWboYnYEf51se9BPWxJngSHfV+bZ7OWNjXKyrJ
A92jxyrmKIwSYLY+mLJNLlR3Y6z16whdyj2abA5YskJFniJ5mSOQugCYSEkiYZuN
zqF9d+0HG0JTaRxhbSiZx/rxPsWmGKBQ5JFbPgPJvMUB6xa2rf5n/Rdion4KImlK
MmNTfY3mYNMSZPPYBzeFiUqPbzhK7pjywF+tyzdQUGyC2Yn4ylXZ/fPXb8aKPcw7
OFCvCblgFJE4j8OF9FQtKXk7/Xoh25u5B12KBmzlLZbpwPsE3YVtVC4T28ZJNTkc
ZU1XacOqtB7pvQDgqIqN0KcziNV26g5QzZQuPOvMvjDMw7Sp8n4WPPDYUje4vQCN
p5tMw1PyUffPjPKIycufLG3WVvSesSHV4tXQAEgvbe5WeelW2SiRYdlChY7HLDju
I9l3tdFgWoHE5ZblEddzOhQWFjX2Y2PnLbX+s+GxmKsG8I7oSJ+GtbjLTmoxLS0/
kOFEKZsDVrHV1sCwrmbylZ/Cw1yOTbzsXbbvVnrzx79Tk6n4VFUPx5EE6eMS58JY
y3zyz8yHdpEEdWA7YL8eed+Z/wGdJ+zbEVhe0lCeKpWLGsJldfEDxjvX+UFEMU32
0zUmkZ49HIBxBSxvuFHlIeiQYt9OwTD0op9jDGhfkhaxVlmHmz83A41bQCItuK/x
/rDwa2cQfjSJQh0HvgD+FxDU7d4mFaQqvM3q85MRVL5td1gkR+oCVw2P/1+VR2yq
yJTVSc4wBw8gRqCmGbdChtkVkdq1Ws6NR4oUMjuOBTQ7y58ZFZCV71prfEdLJ2tq
sQgDYPfDqaBFTyQA9Ab43Tq4zC00crTM+gCUkucPxIGW9WCEB7cEUBBIIcmaLrvv
XI7Ur3rKbfKysyk5/Bnf/dnOdUoad2SIG0yx1RnJdKptp+QfeMnZKuo4YDpVL/us
dK2ju99FxDrVyM6Ef4a0FJC1tuTN2R902o8tS/GRoFjGmIjT//ATeZmkA9v8lXdY
B9F+1TuFj2FSNErxMEiv6QyO2vB88AXgfZ999GNuksDlN+N2iCin5D0B1whOcMxx
G7CULP6G7rfKV0+JuS2rqid1zf8ahm0boAe58GIoZCY+yZ+m0HkFJrw5LxlZujOU
Pd0Tn/sxGKM9h7ntayYBT/7TpNaGBocpf8iPEi4kcs+FgUKp+WFbNtYEetzxzVT6
/t73uFYiMB+wnPu3n9xOkGIIPniwuBf7NxzVrBix4DO/60nUt/zsDSwhmldPi77b
qvot8iUpSZRnivpmdmus4leNMROnC4j636lp1X//3p9Bzunfn0CQCVS2Wdd+h+Zn
z9GO05QyBaLvHNi9kurMsRAoZFM2j5cl2XZw+vuJU0cMsebsWFEAy0diuV5j9RGd
NxcvXiR4Ka44MXcqzbvSmkPPsu7btn1Ch1o6Fbs73fbcKlPYrhTNrzA5J/iq9WOm
dOfb77aj40ZpaXvj2bIlGShGJvsLIOU9PnWXz/PnTB2YiAWef8YW+/U2YLkfqiiH
wYT2H1ndheh6FptTVwT/pQfccxxKh3sOG3REV2QFS+nFV/M+VAddj9oda0eU9/bH
OwU36NQQCPf0XddsnaKSSNHcMt5i2qfDnIU7sNBmmLTJwVkgRCaeDSCSV+fwed5F
MDXyQj9sPdGJzASYA+HRFQyDteWBqwTUCyr+2C6xdmB3LrFj/GTKg0FqOSe1wCiZ
1LOYaWCTxrL46/Fiz5+W3bEny9WwhvSh6UsPbT58orcEV0Py5Pbm0nCrhkjtpA/R
VgNGMty8q+y1lhow7zyFQeNHtWoNuI+C+H/UZCdzel57PzReCXmmdpcdwdTKPppP
tJwMSfYPgqDqpC+wY97eIK4/SHYKSgmDUU4qqSZhJS43CqsIPXsUYaPp6nt248D9
Kq5vxMl+ZS3la2wogBGFDelVwSEEDsJMaeMnFyAiJxDWCDHldAQKuj95ZpmCD/K2
/nhPuq738VEZSAvp8otqis2V6Si0T88z3kxe1/byzy9QXLZ7x8uuCPo424owqBOq
I/7mK9K7xdSzuRfqUdLZaKWA70XuIO2P/Vk91EF6ZM7eF52vkTyITRzdskEixyyd
fC5uvEDF1qnY9xdj9RbnJfK36GKxSr2SiNDUl+hnBh6kyBK+Ao4rUY/gXX7hZPWQ
RAcAjOVlZH9eyXRPwBf+7DiZVkHl4vSjj9y3xFC8v52unbnib9Bsii4OV5p6YaFI
Dsm7FUle1RopQUt0RyWWU8U8HKez8aX0z6fc1VnX5NKzH21dtICquihIKT6UzWwP
zr/f2kUb/VxgSmvYQP6dxaV+kdQz3I+D8dQo12SMcXaz25SdDaBG7vJ0E2SOeZnI
yV1BI8OpbaybiBcB2TvfcnP1XKnJFRQFklh7nfieQ+iXx1oKBA3pvfmCg8ad9/Wj
EPFxS2Xzn+I0+j070NtG4ASc2AIQe1HOWJYS0keuIzU8yn81tIk+tjZVrK5U1rin
LugKGibFccR7rOBesaK5aoLIWgt1kEBElrfPtnNzIoSQ0P3Lu42MvcWo0xJc8FdH
gW2LhQvA1fRfvKu1Cjk00NQXzNeEiLwLb8q/GTPCuEgYs5v0OoX7fhWMPDnHjP7D
b3xJ2USggZpDu3TNcvzmJiZpVYqYXAhtA8cKDOyFXqlp16krGNVdiEW6S4hZeYhO
ym4YA9K9VRTLpTQQZUdH1ioewB0Pj0xkSWFawnsw9q88a0/7Prqn+WSAl/iQtmCv
M0nt43XM5Q8cI3l6KMmF5DVmAL/zEI1Ehg79TgF/NI2v/XBJ6q3EgRURBVKrmzcx
WQAZEWx+EKYCatUOC6Yyu0uWb8lgjkRzWCMTvPNcz7/Ssyhl0+aqywBIxoUEwy8v
yv3qpeUUraZJ755OW86UtQAQ/cSV/mdSgP5oWm9AXZB3SBoVsD5R4PwOBZkTIfCX
jxJkDLzazOaIzPwjJsXAhufz9a9S/KhpvvnFijAw1kAQP/WAPmF8Lqm+39F+LHAO
AmUlhHrcjjYEZTyvvzlcclgRUx5D82ucwEI/xQugXINb1gYLjkvR67FoLKwwefkg
RfUpNW2zEw/cA6p1yH+dLwe6oA+dT0UmS4wWujwtegTDuUOQclCYhGdhVRjLDODl
CiW29a+7bE448jHf2SKVh3wskVSTr6VwYq/Gn8tqf4bKBq9Swwhrl/tqsWoUkM2Y
+ZVAUdmbKb2iBxB3hg2WuaL20x70xZqqG3h+2uHwST1qF3cT7HsU2Kf9uJ/ruhSz
NV5H1EnxqXZy7Aw3kY62hYnx579/5Pd0HJqIz5EJzMXZVxiILUuhmSslVu5A7dFs
loAFGWXWgPdqouMM3x3OL+PJqKjZ10RrHAbShTgp5eR9x6tgQd+izYZGA0d/oHkg
5Pmcc0C4cCeTQFt6nW4OsY0QU5eATXuwJ6OcmLP97uNWipGJlRGAz4sneqKq2GNP
m4B/WKTD+CKSaIJbj85zCLGR8sh6E1M3ca6yt29Mc7oAyqQfauoPBysv0g1ZVljg
6uaVdkAIO+MlrZa7rjGxLEbOUtqa3uq7bWVn22DcCcaCmA69WKmh1AgRJvSz3DxN
O2CgxmU3en+uWYbRTTxEeQvwqqBUUgWCkHHfH+sIp819Wl1K0nttoLvnemlj/+ct
ITcS8MVxsCCuWRfDDX2fHeU8ocFLF/MnoXIhq+Bi+ioyiTGYUb/2Y0y1Hf2UAu/f
DyJV1vmDAM/AbwoD8VexxRF+lR+Uo5z8NlIQos/xawL04ldENM0pETKi7JJZfKqB
9MB4UU7PmLezsL1OrxDLfdHUpfkHKDKUuXa09HGGOif+Gg1LQKrawTuYGqGHA7Fv
nncKmVvPBqfZHRwNQVS/WARZtAkk3zlJnkTNSpNNwuARjMqEkVkZSpuUwQDCiC+Q
HaYC+aldq/nIKodV1DjZaeqLRxUGCsrny0eS8RsKjScCk7WUYYnqJJ31BEgqsaRj
wqylUhbgPEpc3QoYHd6yf+XmNLhLZdPX00HO0IshW1Wfc9XQWEl/GmE8G+l6PtSw
vAMEDo4YXZX4x3gVYoE3BZJNWRdMOOfz4i8fc9t6uPt7MdGH6473IaxZPGIXPMcq
RQXHU7UbKMiJkU9c7hkIXeY/38nNw3xb2ASrZMfsZc8GM4DDT3PSZRhFkY/sVpIH
V9sR3bDukqjHd0tnlDkSQHVqSZ8QRXAY/+dwX1du3XA8vWT18y1MmSoiwYhALqOM
qyfq2rGw9rdWR0XTiVXPJ3iUzAyCBaHdFJEXWARE7TuzmfGkSIKxwufW/fzz+2Hc
Ea3v1SCO9qXXjFHW5C4QatoWHpgfJQbbdJxu649ftVLWZOr6LriA1wKPYna8JYri
VrVlaktoV+OfnaRulzzumnSQZSK9jvYh4FkddnOW2NR6ucAcNsAlcSkcBVzlCeOL
j9gvNIqRqMOdWsdloyR58M0GASOrx0oTsygaNOoCUgkDJW7HWzP6RocQtZ0LJYEf
JB6FIlQbG7epq2pUHf+HbqobKBrC7MY0TT8KbmxXWEZO5JhYu2QXmiIE7I8b2Avp
mSf86n3UDtbYfKGL3aKTgoq1RvzeaaV7Ymg/KHPKlv+jMNG4Lvsy6LQXI1diYfKd
dRtcbEfUYEWzLPeovdK24ApJGoyNDzvnN9Y81nPlmwIEhJNjrBFUeO8T3VNA5lFJ
6IVhzDmPxypo0TC4l1r1TdvXINFXKcqU0hmQuVJn5Ybnn2bJNmQVztTiv8mqaYMv
c42J9GZ4s6FIrCbCYKHDcMN1ReULtf4xcGX4xwj/Ues8w12AsyiRMcggGO+ENdPA
yK5+QLhQsbdhTSnv/3Aa+kUEXSQgIFf+ZaU8FFKNvnuPn3UjOkZOWgTKo6ntsYUT
ml/xEXMVVyo2d9qMauf50qNLlgvDcUFKNaNfGDzrAdPTkD4fy+Mi2wxH24BK9H4/
fEJb6xCJVJEzZpDctYKkjC5N73wukA5BH6FC9mBHPNqKnwd8v2ficjgxD2Z8nX8u
brUivYK6t2SuU7ug+hf+sh3B956q7g/xaprxqQMQqzZx2+2ESPf74Ss4yjdTmeAc
uCtz51pcr3e5kJJpDDT4CSG556Vrpbwwq16RjxM8sekD5qqEMD+KTRBVI3Re2bhJ
lYtIAWfbEob7s8NFF7hvSiT1mdhW/2YJK9pziHUYSw7FqZLMe+DRPAGMMLrTwZ0B
sdVJfgfT1YIPDzVl85/4mPttISz2rpYvc5CCNPS1yGDlLQZHM/+qwhuCV6Rp0UYf
lK9DCnnmhhS1h+RUIU/DqHR3doqncAF8grFN1gvTbN2gFtV+mXtDUooTpe277H3p
WuykLql4WIBFU3mvalBMb/71yT+YTbMJPi6xmZhpm7zKSkBqp0BotKmJQ3JcmDwM
wrAn45VEDSKtat0TR4wXtXPDH19TWAhzcYtXjV5LbbO/d/c2XgdUpYvOLFxeNlt0
4algFMeeXoA50sfVLRqaWd1E4GR0oODr8MTq3vsxM99EYHDlRXsnoa/0tDvig0qs
sa+vh0e13XkNiPux9ONOTbSC+184uqRUwSWesc6VVteEVOZoTHs+9AO2WDo81jli
qdAfD2OTTABcqeZ3ZdLRGxqBEbzQ4rIXlf7B/LIQwIkO8XBfO+16DO2YuoOn7iog
r5+pLmf4FJ/0JiSC8Fd2WgBuSispMYkZSO9Z4IUB8eX+m3QV3VewmyxGa8R1VEO6
JWV9FfTVC1n4fFtc9ABV9E8MU0gEHmFTvoTEkXBdRSLzfoPn4sJTjAtMO3mEmEAp
ZHzcshBGzKPnCjP8GLjf+zAhA6UXjM2kKfLBkIHBF5W8BiswAsxk/UMaKjXQE4IN
na27z1wn1YM99ZdqRfoyH+n5ySYuIKsiUJfqR4zgAdWldwV/n06wPbZD/EpZxI7b
81Lv5VWQPTSjNir+6chh5mkEaBag2alLkQJmTvY8czaaAbNz5tYQFUOfpI0SlLH0
i+1QpNl7hdpPOH9JJjpOw8DhjxT70esX2c2b2x/jUuAsdxDJuuhRl2t9fOdXUrrE
s9E73e1SlPaO+onG+g1O5w1ij7xYeLd6cav2+GWSh3Ji3DSRoQjBfguXaK4fpz1F
/Hgux9beTCoWL3hShRaI/tFZjF0kmgVJEUfjycyiKdL14Ia8QVec1JHIghbQth6U
6NqY8fnJfZpakWXzuULHf3ZWULuiPHwQ1Ahl98fmeTYilBVbnKDKyU60s4QnQ4+0
pONx8pHdXIxQjgjt62NS87eL+MgimQJuoTWUcG0U8nzVMRozvuuFz5gKi/EFaNgM
LsKEh1LI6SisVWLI7ZsjbslqN7Q+FDxUTjHCWK0BtKS9ggYvT3tlb8Dl5zLhdWvr
nvt6JVEQ1ZD5WyVIV02wfmyKXKwae8wKqSO9DjBGq5ETVsa8wLzOTJVBAmIiZDQ+
QpfdMWfPaXpAknTdZ9nrTiQ/a/QROgbQvsMll4hom8LuFK9BYIqpp2iTSLCU3+pY
87qfssaf8ZSIWIJhFhdJsZv5TGq0p31SvaS56ZqtxQ5IkbWNcFck3++h+Fwns76o
ztUVZzBtM0DcNgy2yBLxT2q4av6mHUDzOk/AWl6ytFkqLOAK5OGRShNLqcdeH03B
ihrtsqD4FN3THE9O2PyZBIs0Y91Y7i0zBIovIIqkWbljONP330WaE9viM7WvVHQH
tIK84WbuaYj5+St5qOcaphmzZwWMwC7wu13rsw/WdHu1IJBFH2x+Qh2je6mk5Qho
L0fZtYcfLPjIPDGc2mcbpdNcpBX4z8Rsn+/7STitSRfW2L+Dbg86yJGGXTCSYKnz
TY5mjhyyp/8CwT5sjihumyPsEaIh4MIg6Q3qkLJ7dFHsALpj+CUfGAm5ZwUvNWcv
bVVZDhBX6tTNfOySlqnLRiSIzpiapRFOujnJR932hgFwwh0kVFUxrJSXl9E67Jop
grVUEM3xfI56Vb9djtKksHIZX7p1xd4x356G/6+LRJbK32tK/OgQj7bnM069MX0O
b6YGPMq5ULdDCWa9nq8KBkH0HvFwW/lKdkZwCbOT0NjiHIoHKAuSrTMa1G2NOo/U
Rgtq0tzbnRtgzkzQcfAP5rHtMBbyqKp4l3vMmO8hWHsU8j7g4V/H2WJB57UzkeTM
4f+GsbkefpMuYeU+LlUcJSSIHUWGqYHgTLAMZxi+bhkP7p/IPnk5Ri4aQhbn1tKq
fpet1xec43n4RdikwDRCsSjlOI92ocvPIIloo02aorDiG+PcmG3cedDjeZG63AUa
91PDKDIbZO4vjaSccFx0K67X/NfQzSvLeR3p7GbTIKR5xVvXH9c7m1aqIwH9mmzJ
BdKjwGHz7Lk/Fs9FNu3OCgMcbWcEuovEvx9c7fjVwIxDD95DAbmojqPg487nAJeB
2jo4Ix8Rrr1qEcMVqAGelmbWZEcbNOYL0I8GDc2TeqcrwRK92l4CaalfuHG2HHNg
9qU6mi0UInzfcs8JGB70p1YgVNfIJedd/X+7moTaCB+VwRWYJunOkekeRCDIzksZ
7+fkxFcVqI5ZSHHjqPUNANudpSoZ9KwHpPQfppRWYLVR9gOMoYWVmpqXR4f99tiQ
rH5EvjI9IKQT30AZjxIXL4AXNza+nJdiCfihqxzYsH+EcJqcwrOJdsA9SCinaxcP
udR4IQzolsKhzhX6KE56HSfL0C15rBvVRZdZ9APU8sOYrKwRAhI0LoGpb+Iof103
uXjgLnPgRjAcmedGcvPSj26Sp2ytVmzSFnIaSF7B73SDISHnIDyo5wNtuHkfeiTN
iVAUx8XYLL1W+HY4prcgCaX63yIlpjEWuQQfKs85jAlsDuoqqBjc3mDsjw7jcqot
2RuhkvgXUOsDpxryCLo5GAyOlAWAsp3eG0n/FkhWOs4Ya6Dh0sasDoY0V/VGa/j4
ejsHYbUucud26VpyRqyMr0uu1tAf4wb3s3y8P9kT2/4s81p9yDXivulaMd0SKZUi
Ud7LKCYVi5W2ajFy8GRCP6xxonpnsb+b6CBlM70iA/ZdRE9yycC7bqOtGF2h/Zeg
f6FpAl/mdLU/v0TLkyUMJT2Sm2A9N9+e1i0dXpkT8cSR/WdhFJwMFyEmne44L4tv
sgCBXq0fNg2g7xlUTcjP0BUXw2pkHID8uFCTjRYWYQBmB9bV9CXAK6wriqE63tAz
HsLPGYnqMcUectEgbOZqXdfEaI8U6WGlqzspUuDhzdjV/6yF/ZfMWslUQVgEkDTA
0cfgdqy6sGhKQr7ovSztXP2vC1U1UazPR24jevYerZQMNXLTlH4D03/X6q8Tv+9d
k2GiMWMoWU7Y7T21Tk+18OPEXScMIG0CdlIwDbdHsftcTcSfXdLQmw7Frpb3txvb
dt73t96CGgX8ww1lXvLuMhdcTKFk9AldSrf4w0U4xE01c1Ai6Oj6SUM+i9MBYhXn
NL+u7KpIOiBr0EIHUEw1qAWxMJ+CBVbcMg91oLsFs032Z9oQeHgIBTRCpDHaxX5S
NxFYEP+pBEEIrNw2q+PG9+MlQ1ATYzv4hw8qUSjUpM8IN1KiHSeYvyMiFP97IJ/6
0KL4Ql3QLIK1qyzF4evrzdfCNukU8/bdEjjKrC6pYUwpbMPvB5D4r4735tpSqOPb
IJtSnoY2XYEHPDD8dPZT8kkC+rE/aX6dW2XG42afNuMntSJnsikzPPWbSzZAVtih
I4ujyS2jOD4/mLgXhxYX9KjQpvm1qF7jMiRvDhyPQivkxmsAVXY/OPixUR1c1tdC
z0R49QJ3G1rM2zEqkmPvjgxZX3uh20bjBPt6FyPm4lkvwwtuCcHXam/vArboiDZr
F7VjjyB6Br245iylInsTu60Q2+Nzzs9xeyCgvaOP0/Hg7Wz/Ds370SlqOQl4xJFs
6WnayFOy/08EfHrf9fDeafBbye2/S+w2j7w3qAWAhqpvG8BE5AOGPIf0FSLlyBPN
XG6n1tcm2N3NmzJKNtd83tWbW7JH+AoaSxymkWholIwaizCn+DTtpfi4HCwOJvDc
XkcnhbowbpvqmlxBHymQFrSuFWsJBgT3Kg6JO8Db5FjGY0ipeS5EUblavgsIFjMB
R66oE9VRQ2FucO4t2pmYDaCm58a7z0HOJNo75BgvThxb/QFkbFIOUjlShfiOVzoQ
GvMv5S/VRsdvrXb5J8HCAEp3WS7CgQZBiD/nK8By4iWhL2BXV4BxOvftEDcjhut8
H00XR3ztPEFXAl/jN96i0qH2560IVgDq48xV34JSvJZS2rHvVMGZArYZKEcWTvs3
q0VJYnCmaLXVAMOFFtF5kf1PfV5pZ4fwWJPO0dGrI2dBHn9BoGONXuAgugCzXpVz
hL1nicJpVV71BtV9J/qQiFWpHiU0VmQ20FGbTFUu9qxOUZUgoboPBhGdt8raYh7+
wdQ1M0YmcOub1TRnoBM8UlnXY1Z9kkAnE9hWySAMfLqZA26eWodwH/wVXbjSwUle
NgittEelbTS+VpXG4z7hYwrx/i/KM3zjDZm86JNvx++twDa2eZkBPiJNB9L61SnX
vMLE52BkhdgsmeeIXvnQB9wvBcxLo37338JDj/cn3kIRUYpyW2Zg4gsaS3Y3fjEx
JO6NJHyx6W6Twe0BtJLVDZAE7byJjZoeDp94sArSwyG/Tcyrk4TsQdI1QRzcBtgp
pBeurIc9lp9FTHHersESodYVhq76HjZVbKQn1p7BIiZJ/laL6cFZaCFmN2DhzQ7j
+LlIk+lPZIGCEYUuSl1EO3+l79lJL6Jq+rkrc0OHGX3CWR0rIFv4PYKDurHcbM0P
ZdySAJV70thY81LVdwqcE/oLWa4hxW7TtbQOOB18iIH4PNOmGb3MvUVoQM4I4MjD
E5KprwfebGynWgQz0vDIGyXSbVSvw+O/VxVrYc66xt/Q5toKucOa9EvzljqfGYVm
3rNRQwbKGMJ2s3/NiD4A99KYtIjBoWp7KmZXaZT27GrLN6HRmziyovDkcL/rbKXS
YjvqrWZvs+6S2my+w0qceq+d1PiL2Bfr9qETL5GKDu3sG7PtywNiPTZIWUYtva5a
4v3VtqoZnE4uzoNWVrzs7MHjgHlIa0fb2bFUCfqrfrTX+SEvJThARdxJdbkVWsR8
y42J2Vle/Yoy6KNfrwzDg77yGt4ZO0RmCTboKDBY82xSYz1C5wsdVPpowh/wWOBJ
1OuXE5WKirangwQ130HjucEOIsxqHvaajiUBc5fHexSxS2ADWkGam/g0sIet8ng8
ChNrr1Qu59Ag/0z0jE4s3a9qF4vFaodDnM9rnwKFonevMoitSuhv8tuIIC6irJeB
yI3iKtkbNjwCN5q+5IXtHD5t9K2OCyA3t6E1IpJ8LRySp8SLjEAVEEVgmY8RiHYF
5Tr3T1aQLx9D1QQCWw36ufqOSV9bhvuFZIKfK7aGJUvDJD1jDobp636ZmcL/Xbu8
wojtm1kg2pIO4QRedvIYA/J7caMk/gHjWZwTVjHu77FBVl69YvGZsCzrfFntsI29
Q9E0VSW98Po4n4jP4iR92/GY3/rdzh5ssDrw4X4lCigU2utTutG9Qa/Nrib4Ag+o
4PYZ9msjafDBMnRtGKf6d/t5MeJqC+x1ISVQDQNiimxia3HuGesQOc9a5jX+BOx6
Ozj1UN05X94LgOffZ4DCV/jCOfNomwcUgfZ78XmPetfoXsGSncFt7zWjKfKhaWjd
+y8OIGQNhWlRPWBM69dsZpuW4biWkrNdr/bJobB1KZ93ctmdtIXXpTyl23O3fYjE
V/1zRSwd6vfz5r/kjY9SYc4OFrQoWo4S5STxkWKbywPHNUXOr4alOGCh/34glxs6
m9lN3umF6+BTyCnhRmY6Kr2zVB6CUMZeXtF5QodYSdToYz0AGjenQ76k0+lHB9B7
UmLzDPDsPxXvdhru2sY35dd9sGIaQ152CdQ1UE1+1np6fu+z/kJoPbbxetcImQ0X
u//POK8FW2QX79gHkYW6IV3Y9yQLc9l58ombRnT628N2TF+S8fWWRJKeEm00USIS
ATr168VmAb/RmqZT6fk9sD5Prly8qVYsURGICcyOWiCAKZ52OcSkGxpmI6Zlzx6d
7Ev4VKANKJRi1PVT/c8TbF6h1AcOHd/6MjVgv7aYz0voPe1lab1WBwUG9p+aeTIS
bf3VGx4PzLdl4zIwlPzPZX6p9TBAUNTz9Nv83nRdKbxljTTBe6/3hDfJ6b/hw8SN
ReRpJAHF25DqbU7vva8W3s5OY3lCRoVbBsFadqEyqDvetpiG3vpEg02+s91fairc
sFdOzrg+4FvSziWGVVnN/ifGOeRdM/ESA4i3BnTEWlXSUfCWDlp9hW+Sid1f2v71
hf1DDK+7rEzAlHrKSbV1WcE/ofu7lo/dnqkYrs+TQrJezxQrJUcqbl1TKx1IVBzr
Ry2UvjTQm3aLFcRzUl+Yxup73xh4Tt4ilA/WrD0JuNV9IyNAYBifqFKDDpSFo8HB
Ubdgrn/SS9ecTgGx6Z7xMRs186HWR5eXDxzPaZ87mumV5xXTPwjcg7BZCAGsbg+3
6LP7soGizzfw2/5zFhhr2mq9WTfrGzRy5xN7zR39FFGPm+FinL27sMmu3c1rP0OU
ghBzxQoUIikixpYZSvH8t2zrHCwjaaSBDMVO6aJP1yGYK5YtpQQmYf7h5SUdIlMX
KmtDpsmdc+HNfr3Ff7C9dv3Du7wmuM3h7f3maVwaC2f5i7JFsDpCcA4w35QHQ8G+
yLzgPYTT7CVlUSZ/47f5MRJGDXBoLOhHmb/lgrIofcran72gDGUPB8pbFyzbgl4a
8EQe73WXEazfdYUY7c1TlrM8ogQNBdW0ifoPK79357FUzvaK2hJ8km1JM6VTYhfh
FsGQ008SFoiG3N1l2BQK0SqrW5pmkC0rgthgd6TJoclUP6fMU1rsCToG8iJ6C8Lt
wNRM5bZczT75A3F25wHsvDeeQ4gy7stw2rSdSq64OUPDk586HuV679roHurmdPi2
soIgba2v/kugATjqLAGzHSe/9WImtakiZLqkxK0rsOlv7a+lGfeE5ljlTkm78yFw
iDdk4b/NrXvISroC86VsG3pCMPGO1bbqlO4zKkXKosXjAbwRLBi0ASWe0B9eCeTs
Lugotc/35FA3+lylZ3MpEEpi42vGYg987pUsMXAVB4t1Q4kCnUbQ5+8Nc3NIZxsW
jaQL8hUdQtrJbO/Kt01hi65jQI/y9PrdKesn1VBZv9hhdosOn9M7DNfD+AvYbGnj
BRD18gaBzoYcimKAoOBy9ZJWPlQjpdTCNJKrXJiEZKJOJaEClUIZIahrlVgTcnhs
HeyM0KAs+0VIC0Gm7jNfNdOjvFN9k3OXY4SAPFs4s0GozNhDE8Vc7wS0SUdzMkn4
A4HfN8W2fFk0ujxfEk1Nf8NQbRToT7ILff7Hnea2RGaKp2Ik+gw7CJ9GHeL+QAQZ
Gz2hJ0iQ3XLFDEHMtHG/UTKkYwHQtaKIa2I/VSX1hXrm8LrGP2CwjjCv8yDV4QuR
/9yLqK880z4VxSfvQuRI+1pm3pQFwtRcgdmxxHxGV+DVJKCDPDzuPNSKGxbGC/oy
9oBwUNKjg6ujQZPpzDtA/Y47CXToOeW+Lm6MUuvTLyS/kRDmVUy6eMcvtUEnYMzB
MeYNMfEf8lkzgoFdTz4FGa933+2SvYdiLccFLVCsV96j+ZgVaiuOXXF4WDFQadl2
lr44NIFEnbjECeiZoG+UugCrqU8EN0aTqIZKhGjnd8BQtTCIhqL7eDatzwatp3kR
EyU0TyODlG3BnYGeEJfS2doi8ge8NZcYmLMzEkCK4Z+Nn1tnYdYS0dxOJ8s6dzV7
uuNr96yENYGt6sk/V57Nv/Pnvnc1mfjkNK9RV1KmA9svMZDVxOYds6qv5mFySeAK
3UBEGscDrDHo8MRyky0NbehFoLfLPwzA1oPtv5ut2VZFxvuwLMfbKt9+Lm8BZYLw
4Iyn3nb2qG/ZgZlLTRjeAMPDh8pdU/3t5PH9VfrfNkTktsSH7SloVQdId3J8Oo24
5/DfFFeaCW9+z5gGq9SFawijG5T67GAKlrlaqXnVHKDzt18PJv7kCq4dhUK8Fe5w
UMU/zCtWqED2pfwNHQpJNwEGroAgnVA9GBrmtBwyCZtdbbpSRhGzxZU0XWalYdVZ
+IMobng+XgDbgBXqrJWjxIq6gvsr0wpPsofxltaY2SPZhGL/jrnzZ8Ej7RCYJA6/
BXM5Tly1qVmyQyUb0VwTkhSRqphtUyq89j7jJNk9uhNhJZI9UVrZ7QP/B8LQbvf/
WyJzkyyf5rb++tcLXM4ngrNNggvDDZfcFc88xR4/4kgXERE9SQG2o/scmSRZkuRw
0b23s8hIdYx1SywfMvH0iQATlym6ODv63ODvIRAW2j1iLF8NHArjHOHwtDHm3shE
OHorpfRIBfl3NSy2Lbrrqkp6PpAxaHjqYyOK2+YwuFgVsyK7+LRZiIQC9Vtg6OZP
JQFZhsZO6knS//fER+JKIDy/hbV80VJRd0AZeR9mKgyb71kGN4tPDWY44+Ar3Mf8
vzr03kTR6KfdkKjYkZQYvxQc3iapIyGavcxahWuuKb4B9GPzR4S5/utnENINofY1
ss2J4Doh/ed6YfN4s7azGbEFlN1RlTCR85a1CJJbg5Qc8vabCv0DtXbpvpaCGdcH
8BEgXS0+yWMTc6SEHxOhpyPIpRThtqGKSztO6ZiFm1u4aTtIwuedowdcCsmOKpr6
o8ouPiUcZ35M/3Qeo9RMY1QVfpOqEEhVYvCNYyxTLiXpe6vXnevaXUglfHhTUni2
p9emkfH776YVv79aZYduoeZsXDorcqgV47LBsoo9IoTEBXvh4fu5sKVrmHccOhtq
o1OFKyOSDGgKSfvq26ICwBPSq8HOGddXNbtgJuCMagO1TDAo6CNYUX+w37QAgHn/
oRs+bwUhUvEu0UkGOzwh6aJKBzCyGLAjJUYmq4qBtmeLEovaBUcnSMiV9rO9JXMb
pmBmK/n1v1nNIQxHZQCy3v82S17Zswf7fw0GLFVI1HLma+S9plBi1j/ljDbTDOYL
uC/un+kpFWUr+LGvd1zP+J21YPvNVRlAtpueBS7XeZAXxfrwsl2KHD7Qoo2OMr2K
C2vs4elFLK5uSuzvizjOIS93tJxZszRzfPkIt06e0snmhAf0nQ+jxHwa7nQiyi1l
EomBwlY1QH2J6/mDthwHVaef7NB7qHJvmhDCyel8xvw+F6CSpvtXIGo1o9GhA2jQ
Aunjnx4NlHpp9ZMl0u+f/3PdbQ080fCJXnHnrhX0oBn9s1tBkL5CFeIbGeiCY28g
IcyDnuTWF0sPVQzvYpZStamd5r45MYJ26xDh/Jyx/lF6jXrPa82s613jhhlGuaxK
AJ0n8PbAvx8iLZif6V2OXgn8MjvvJE7iDTjMTkzPhWGu4HVNbn3QtlMvgL9CAE+Z
L0WmODL16y685NcMKXYO/u0DEU/fnTbCnEw0+Mi6urYQJfKM61PTUnbO3/pUnDN9
j4mlJaMdcFhcbzwXg5ZC9TTHcnINeKPgMe/UngbuiNebd4J+Un5YAVM7eHluuNa0
V2wRNHrH8e5Be6SjPsae49ujK2zwkRJa6fjNCIQ90asEGDa19MAzXD32O/iRKt1I
7BFosHuwhSngl447ABRIQIKgYSXQlaZPb3TZyRr1EnaEFEqTeF8nrDbYAyMrdGPn
mkTwADNcmUFaTEAjUlqwe6MYmPf3oB28U4BUUzcOfklM10JQxWAkWN/f8S+x8naE
NgBzNzB8jZWfvTnleyVtV4oe8+wh4Rcimwd32ztwdaldT68T5IacK2NQux3FKBN4
SP3aNtRM6sWOZt6yS9tTfHafOHS+WniDKE8MxCM/PKYthhr67JhEkS4QSbJebKAb
SRZoz1kjJg/QjhowFhTk6ZRSS+CB7aziBXmxJAhwXhgCIld+4WKS7Y1ZI1CkgMLb
P6fuqTGSrE2jEwTR8qF4xIfImdQybg91/axwlfJ+tYekVfw/5f/auy1+yy2t08y0
NAYRx8bsc+kAOHPsc+EQFa7VamE8AEcBP6HF1JYzB4DQSEoZ+IZgbWxr4GmsZxkO
xI3ZhalVerbqW4YiYpuF5okiYq+LBfSjZUVev+OmqwfpvAAuZ0n1W/brKe0QzC//
yN5PtKEyH628QNhQxwCpYImtPdOwSoI5CBDZMB+EXXVSnsot44O97zpft9DLtaA8
pjROYopsiMSxYum6TNnNRa0Ais6ucSUABgvIyM2JMLuVuAl9C0iIhKGOlighh6a4
Jgj/fmMwuzQpbSH8X9fgqQoTMs0hzMjvXpt9j8qckWxyulkVM8vMithrykvr7TXH
VD2gOzZbIx9V0hAXgt6if0fN980v5lt4DkycE0IPF/5dnS75G7d+IYWfLajtqANv
te+1tShVCP32U4kc1RZ8zIbUHdCylaaqkXToWpkhnntqfptHDOp3XDam+rfRdHA/
cWjEBpptTOE84dAqjl62aK8OC8U7DilY48T2RsAd0WoUJCKtPWd0c5bB/KJsZm7t
stmt0HCZ8j0knuibEfo6baPssaijpqEKAsZRZRSJYxAMoW54IewF5ELF4DnHOVd2
o9mac+w4fCLxwU4Vhjcz9CNMWFMpytFhdLHxGWJGoHUnE07oZNtztg+o2BK6uzjC
hPMOZuY96KXUivTRzG7K9Bm+xyp0gXZMMGKfZP2iGfilJuCEtNWX08D1W1mhFL9w
3dqExv8E07FgVIooGi1urXg8dfe2GHFpMvLuk962ZvrYQuwnRogsHkLSUnEC8LnV
57hfze5/1t9/t8UQaEfld7nUHkFpGUaMTmKSq/56cHKiqUVYnZy60IXberD477ms
9OtHuhjjyae7l3kc/Znrlf3d02JqBibkOJPyTibywNMEc9MPtNBxWPuedlpvnUrr
Txf1TANPfyx5QJ1sGZua48MiMMJmLcdVb11r874xqNRoUEjkMRm2+M4jzGjg8KVC
q2FFcU/UINRtMV1Z+ptwDFcKpjYCkNf7XSqlMA5nlDFHuvIhYXU5PRt1dWJ+7GIt
AkIcOdF65/iRL5hDttUUX4N0zuga+mflbOWfG94OuvlTk80rdfaALsuHzVzN5HbC
MLQ0mvX61jj9lEIR92hRKauIKoqI61OoGkizKA8v37zmKdImNUSGrNpFiKTLeaCu
X4/5XyPF13REZEguSlQTIEJtnKjTmZA4Qt1ZL71B/egHqMH+r6SSSl6Zikfsa173
EI9m+j3KFgiEziwvVIdBQqJXH9Uav6UtXC152y4RZp5QVXSRWaDSDLEjohvJ0QVp
gnzrj+B3RtywrbDRxOvLBcXDc33VLcdUBVk607kPTufuBL5b8jGqTqqOImqeuiZ+
uVFKpdi3Z7iSyuvUcPj5ccB3Z3PEBQTyzdC+scdNI+g87xkR7EnSkorGtSPb5T9/
UmCZzBvNlh2ONG3Wgm7M7I/6Wmpi2It/qROs+dcgf2ROhSVENpVZqPod7TVQL6y0
trZxK6IjktcVZWQUVKLiFFjwZWdKhMUBCvz/ei0CoqP3hlhVgcOWJ9yevXW9BQAp
IbWzt/8rhYrVry3riFcfW9X4l196zD3+3SuksAG8zBy043SXVrSx5cgyMdeH0gNx
kP2PgeP+6Ash4P7lUN6Cy/4rdHlZ7BAgiNlfVwM18pFLbbaUSlAKn7bQXL2k2OrN
srhC7gOX5wHFUlOfGvcV1Xtz+y+XHTWteHImenXE8T3JTYUvRXccs3xApKumrQ4P
Fwx/hHBRHjA7PbGngSQtSk02k8fLgQiyfp2SnhSkGor03sK4dgmNCY2bLol+iF1m
L5nVFII+Lto2doIyeBnCZgc0YbAMuuD5I8Jm7OoVxULvwS3pKXNHoCgTCzrtOZzz
RF3gQzf6mHH2/NecDTgkhkVSHpMJXafI52gONpGhgkbPYHyvpWkXGdpNNRJIXinM
JijoEL10K7wi4qSM6swrpXJ6rQSnFsWS/bad8ZqkGrh6ChCZgW2WL1MohMy3FiUU
UFpWl9SVl8qPx51Ik8fAq+gHtf3iBiPiE1oc4qQDDUct2MZPYy9uMWmLyomSVdcF
GaAJxzcMr0aJ4y5aCTB3seay5neyoa0tiL9IK9suGMNVS5YMuR5T4lTyzhbj0SLL
j55WpVX+zEv9fIAEZ2dHXJKkf0IM0nqw5qZV9DDyre7AVtCo/GDPqFkkYtt5Jk8V
EEIMm8gu+FDhEZmnz5xf91AqHUDl4+2Bed2ZhTEwNd0AoQfYfw5cZmnnZPBm/La4
8YWa5byR/455ijJxfiBD9T0QIv0LUzGOPsSLG6iruocdF7v5a8JRz5cNPPoVnP8F
nkSdxJNmY07PgIhO1NDkQPz2E/9iZUUHJZChYCrQfmBQDZ8ISdP2Ckr5Cy1F7AOX
BN8hBsIl4dT8PH4boz+63kWkWD5tUqLSosmdAVJe07t4m8ZCg5fYSg8hdP40yO5c
cqMfNmyZtbZeVIYbMTYztTiwZJaJPIWIRGymt541wFyQqp058xWVLLLT18AzmRbu
upxaCOY3IJ3U4hOzH7lX1jnU7PlWZ/HBJ1d4h280k5b7xWRdRIwNSsh17q71/Zgy
gf5ZlmsRe5EOtvGArM8d2Attopvwhvy9OiE9RCOz06DVRHja7kgLOx8Mb/FINNSn
DeyZJG+vxELG6axJAM6wzm8Qz3LCYXgl5h5kzEZ9ljI1/Uce/F7Uj7zD2NoDKeEp
P31LOWWznDasd9w1sEvJiW5v4jRhAiBUJxT1/HXnotJfKwllsRb/Vd6v0YjCUmUj
Qda539hNikFf2+rxhVYuPPHXWLeAJKxffBOFoIGSMN6AdH7pO2ZcE6yJNnmnEDF3
pUv6Pd0sfeWjE6H+VfJ9rwVWlhDUuuORXSrz9feQbGW8IEpGmZ7D3kj/Vz1Lzrr7
JMbIUvzcHy964s7Z+J1LLTh5gDUoRobGPQUTX4d/AZ5Z/umVAm272CFSNG/ZmeP1
Wx1ad6ComSjnXFAv0DYATEsTX+5uv/mguFg0EAGceqGseXTWsPXh7IAVU3eylP7d
e1gsVPApYgH3xZ1oqP6AVeox6BCJctyiM3MhE+M0SV80JxDhAGZTlPBl0u1zFg7o
2iEswLnYwAnkst60xkUUz3ihgmClBHdJNhbg6lAFEq4E3OjSH/02fxz3sef7IbLv
1skea6+aAoRUrMQ0z1+18jqcOZng0I1xY6+Go5L/BM/G7ZGbCR8DlDX196USx9Ta
qzNkBqyF2AqPsQI+ON+FDjo0EtB7psAxqC/vuq9liHYS3R+PujCf3l8I8lLLJnWL
BDBfLWSuTgWLMAziOfHGu4oQ0KCVbyzfSv0pbxHR6bkN70poMSqeJDE3YSIJaD/I
LNfs8eZMxadOjwVVP6bcyG5/HPLiL+IMnPc/8JGsdud9e7VwEz8OcZrOiu88pdUg
/9IHTFC3FSB1bet7cW5kGVv6OlB1YAb0LP2AXyounrzfTGbORyK3FtzHgbo8kyxr
nEKCS8znIqHwszeFHXnrHvi3kuA3r6c/ndE13/RBAR9xlepsYNDy1nl2NHOXBP3Y
y5MhbxegWGaNYDtCkU1Lud3c0Xh5HNmwePpu9GEl03/GxEi7VX/HwDPbzAwrQP1o
QEcvCCPbo+Mrx+lyV1zPqQRvvtNg0jOmxNf5oLxSylpW3kTBAlrEX5w7qQpAyLA/
rMwbmBe7dIIiAzioauBA1Wx2VLAVfN2emWHVXSZf2m/dFJcq8+q/Lq0r3Qx5S16v
nEm/0WGzswMWbdUTfcw6XIZbuuKHThRy6tj1I0XG2aIsX29nBLviqz96ti/Iholt
+xn4NF1C3QYRBZVjbh4QOspbO/g+ap/dGyQjtMKmk5QeyipWEDb0gCiaCMDdQmfQ
KfpPz3fMTAEp1lsuj+eeubWFzblrvzr570adcdbG1+MT+S8URm60RqQHvpuS8TXF
OzmQ27yyiSQRcN7Ohw1fesxsvisNycGC1KJbAoVamgKVFwgiJJBGsG7aZ6YnTepn
X6b4NQSnu7AM64FaSF3bAbppDG8R560pnJLftvwTDpIrMS1Q62uDaA7Nd8X5gH/r
cc5E//ZFyUkOO4ArjPapvAOm7XHA3yflabTfH6ii1rokcs0TKj6HmZx10DMs5McV
PTtUbBZ8XhBVIfYwlm0Fk0d1pv4XoOUtPwvDsJqoiTmmZ2mIIz8qaJ5QTABPfuIP
NpN9gFZmUyNXVxdl5xKkloMZZlDXY/PWeoisiUtAu9Ag2bP4hrdwQaO60YJnmoA3
UZrT9x7uKW9c9aAQpQYbDPgtHVNQjW8BGuSMKz7E/JgIUkobYwjorgQ7bJnZjadF
L1UMziE8A7B+Z9O9GHZLdM4riv/ZBX3H2I8LoHSyp9HQSWuXFdhSu2Uu/tvBLOkz
YCmIhMl86NLY7DCFdmbGK8s9QXHocoWYDeDRgky/sB28XOh/SgQ7KPmrcfVwDSwg
1PEUAX7jyyHVp7i7sdSejWjQ0ItG4IR/0qNFBNYTNJXEAQmUHdZ0l3/uFdrzPzGI
6U1LrHpYDB+f2s3KXCtgAzTa21KCfjODNEdnqzj/aFIUOeIwBoUzqb0nH2SOyTnr
ABGESTt8uVPJfvZlioIiZsalYFNdvZLhgEdDAY64fYPzZPOdH99djPyX3JrjvoCR
qFUmrJT4IVLh1u9a6tdoe3RVyyUyCylXHwhp2AQ6k8JOMoeDkER0XLUjgbdfXJNt
W0hMNcX2TAMi0BBnJ4E+FfgLJYpXHmHS7SFgjUhbK4PaLfTpi/5tjocEd+OsNElm
VamhLq/HKKiLyPUT2EtYg8dFR42e+jek+Cn8YzkRqtxPEJ+itF3itoLN6iVe/b1n
hGb8ibVLavpeX/cU0ayLnK7m2IRkG/Posd+cFcYVAAsWWMsHU0hegJiwea8rqLR9
XyApdhKk13DD4zaDZ4dzf90EDen9Cy6hv/oeXHtmSq7jP75jed3uhSfw58QMLjlj
b+CikFNJ6YI+1MIlKVt9wtX5DHFdOlC1JMVLrmoDaSpV/lBp/PhkP2Fbl7jO/GbG
ZomQUXFWdoDoMDRMb0wr1XZh4hPSGuUXgJFbQK295UouU7bO3enfeRNaBce9G9Pc
NCZZdmk9sPhrfvytxQk/qUF9qVrywsVYeCwJEaObY44Iw0N3q3RFZkJHLiRDr2EN
p25qMQ6p4dkinrNqGSN4ozlEtQqF1yug6nYS8gl7DRSyxX8PHUrP7vuOJbZY0Hg7
7rkENz8jiRG/4knVrB9AUFPbs32jrJqzKepUqhJGmr2JDRwte3eTRg3G1HqcNKIZ
LNHI8pYcFs++DA9u3yNcGOsjFFy17ndKFCmJ/rj4qLKb9VRntw6ZiOfiUbTXVi0O
P/wC3m5imNcRShOPyaGx5VXLgzhT/9FVlWtE3NY5U7fmyoIhJh7fy7/OeWa5vGEA
eAUnroCQNpq2KahQ/QWbL/EgHJXcVuQNRbRTmKw43wZg4fDtEeCQ1S0DEq8miVtX
T0kiCaSKsdhG+piKh5SycA0UP5qiTzIioZjQ8tcKd18vN8HF/N/rsn/JW1Omv5oh
8K/gvTARcG/Bxf+cCLbYmNlzdJo8J+V2fou5u75QOFiYeT339xxRCU0GSS3Idrzk
A4c+xqqytFt7P3gfFt0GM/nQ1pM9W/sxIRFkaionL/3bif5K3dTk0Li0ux6yp06d
2Le/uVaHEYwy8/ZC/VTskB2JVU5ls1e6f5RMBPRbRX23Eer4dWAmGmYknOyv7ixc
FyBz14mGK/DtIYMmtFfbn9hLjHAgIwxRpVQo216BWx+9WopR+LBrT4rezam0G7br
gIS/M31+4cYtMCd4unga7TTy3Qrkpq/O0S0z2oK82PaX1rM1cxTNw9n/3fwradUX
idjU34GSDJJx3pxF7bk7CmPftGUDYuzsjjIhQu8gBW6iSgD5gXOwWAAdPa8dTy1j
KEvsa319PO0Vu5sjROwEL2j5g8mO/zTQJPdaBobJzd6BmurBseHggrYDMumUc2fw
UnRdQ28oCJunJ6yyaoxnYrzUhNHf6KZDHuWFlcvkolJL4wHAcDbi9YUolsr8u5q8
v+z6ZRNyanMiOv3Vmm86175HdZ+p85T6yiAv676xlLr32bbGaosZ6duYyoC722eI
G4cgEfarmi1IwNi5XUq0a+7YTSY5iPBWaMESlW/s38f2gEEeWYct9yyP3rGO5kan
KIIhMYAywrokRccNukZhTAKRj8gdE3R+WfnLIHjmZbTsW4o16sBLAlTa807ZwXzE
J17MEJRdpDX+2AHkhafMit9CjuIgyWO/EFlgdWRM860x19DArQKuM9blqzA9JZwf
2w5yEqo6nerpvzLHL/QIc+QwI1ypyEzcxEBDgDZWcO3RrOf7TqB3+RBnqLwqRtlU
EF48YApNafoGStxmg2cdK8e9km1nPN3vXn2qHBu1QNm4FiOGkf1axrI7p97wen4A
vJGW19VsbgehCv+/NertyIZSYLCGFFSzKlp3Ki9JCPWCeyC4enyosye0tpcKoN8s
yT0pHG+enBpkm0/sJerzI/j8jZgLS02KKpOPrAWrKJLjXjFmfcoKPiAVKMiGGZg9
n7sVoJkDnzbmhatG3W4UsDmhDgn+zLLuP6tciRnwOs6csJwZZYrZ8srLF3VYWJOo
b6/H9a54RegKPDMIqznaXZYHZTFbi3D8b00T+/eZed2rJqWEdJ4bH45pj7YAYXU0
xdkMoWqcTy0InKWPoj+F4cSDephgaOB/b7o9IiBbHzza+in+1mbgKhltbm/GcKuD
AiEoZiz47SbgjUD6D4i9VwIN7r+xUU9Xu6dJtWd8spOHpLKlm9CM/d67DwVyVw/T
T777w1H1IgeA04/OswtH31tB8ZgR4Lx/cpU+TsgOclBKYaaNIvE6pwqhxBRMkNq5
Eb1hVTDlRQmOlkiZOT3IHDCSKAptZTz3bbEPDLBpCefqo1FWOSzHwxeUrUt8BBvY
glVsR6r8/HF9bu9CC+7L3DAST9XbTQqjB/4/QnocSEDewuosjXP7ZPb7BVyvS4oS
5Ab/7pSnkwY1WLEbJd3RV76hP4nEJmEU2lW2zdBDjQBsFqGYkFujDniAq7inMsSu
deshl9ukxFAJjmYbtvYnQ0dK6CRx9QB42egTE20MK6RD8myPVRXQoakEx1a/sJNH
h+Ayy2LmK3k9k5wiJjU8oFovU0ixtUw9gNNyBa+1AfoXex/RLzOuW+y3u6DVpwGg
/IiwYk79ZvQ6EZcJ/D5OlHcGNlyneRocFgQgHDMcpE4P9rf+Hi0dCUnYhp9GyYEv
v9865UWh1kdSCxNEB8aKihtKiUeS+U4O68iKKxWjY892hK7Mhi2Q+rLRWdZ7BtNE
DUty66eR+J1yDIUUrlx9SC0TDAIyQoE2IWJg89zGblGLZmybjO2SEJtLicy9ee5E
gNIwVgWEp9p7KBmN90NrVe69XlIjdlFIuWx+EwobKO/e85fmAGnrzxs2PLyaQW5N
qCZ7+5ptgOlfpxinO5F2rrUXrX0fE/8YEL5dTd6XGokKaF5991SF0QqdSrXOqRYe
ANyENHJMNtdSvtvkGi1oUEKt5TH0lTLKcvooTUdWVNLjquTVm8irhN08Pd/XILRv
/zFVUzW+llnbmMudxqR6L5ytCGFX4Z319wdU/WPGnOXej5+FF+2vVcTOEPQ1Z6oI
qR9H998wnWXXJ/Lm8N06IpUEf+jChT+qCd5Dkl9O7oz1yRGeBKo4ZdE5msT9U09g
Swz+hgU+0Ni0DPp1nf/zNamfnvJYumustFNTHPf+MxDTbc99yMp5dKnNhCu6OAA9
E2Zy5PYsUp+xuxcPk9TE8fef5bICWqo3zk4HnXE1JW17zH8HyFKCiRUMrdZsdKq2
odhQuMhFXdfgnMV0ewC74T+3FP9Ozg2os+2a10HsDCTnNFNGZpL/DJe4b+x98jAY
+VimL2O+Ea5MUL8cVMtT7a2DBm3CRBUc3jA24KySuK4CTUJQu3+a93994aIhvwsd
muEPJfRlF2mCYhJesQl2UQz83Y/uSA/HxG9Ek24WWOU4hXyXo55qJb86U8OyxT8J
tBN48yvVxEaozVSn4QeZ+6Atm9XMRvbJADqKDVtpGDE+7vNLzV4W3SBOHrqRbMlQ
K5A0WASFIRSdKsR1BJ9eNYepRVMy5fORKBY7xko4djOBXxjAXRorkJnedCbQekFl
c5xpCMrZOt5DF9UfTI3pgywa10t6geojUSlWbJ5q9K5q2yP41Fh+vmHgRp0uz2qv
485cwixBGLbTiCGJwgyTgoYFb9BcvhBmVl7y8lOIhIsxJtl4dySvMjqt9a4U7yKq
rqoPH9lI9nApFoI2pbbaFIRLLfr0lwQcb7mGmPEQ2QuB0ZnGtrSDnaU4cUNOQS8b
PjMY7NDH+53hgqibi9rRTIsxkh9NOKk0dqRtb3P/WuMs1J+ghWk94NL1zGLC/DGB
akOQzzZeJ4vPle2l8eG+7C01z1CoX/yt2QXc0zio60ddNzFmyt1LgskEU9Iy9po7
FZlelOwhSQdBZtAzF1bBfolhKT7FWLSurwHFrYflnRS8c7AZ7QQ+Y8z1A8NZkb4o
REXxStxk/wATEd7UPKnEFCdjKqNNez4owXF4jsi9Khut1wUGZwxw+CQMELaxAAOh
QxkawBuhquiw47uA8yckKQ4zFuYe1+zsBhFP+N1HsDGbcjLe8vILl8U8+g+UOF1r
HCCDfGjTaa4PtiTFWadHJRbT8LX4ARGx0M0FIyOQvTD7kN+ou2rfc00cl0x0oiTv
aEyc9MnCdT2T3mjFWmxXcjfo+MKuKc/a7wgDb3ua4OQTOJVtenFxeIUPq6Pj65Z5
zTLcC4GH1nTLeH28Lz2lfGSIv/I55/L0uDiUChwUXzT7ESimLaGATv2aWs5Zx9L6
9x42FABi+oPH46Gk6gcFpO0xMuHKGWPr1T2wJ3Tz3ZkyKPU9R+oKzNtWDpVBomWM
6T/W5z8moy0G1lZoOveRto+afv2tNlXAw4H3PTGC3eJF5kq38hg1XPdI+CUXrCsd
GFKyMZgx5Mgm6gZmDtwMXbVPpy8U9tcaXb92ewcmpvdoXbeGNS8X9Sat47tUKsP5
pQ/XyPOtZjoC4oYY3zkDgztWmCGRKYc3GSLl90WyXUpjZGgZtkhADDcGxBQN8hXh
h2bPAjoECXnanT581xquB0WY3N1oVuhFHoI3P7smL1C5JZA6OaByd/ar/izw8swi
VxU0YNrzYRRgIVN6tJDg+nW6/W1yISsngUJRPO4aQVYIgQ5dy6QDrPUAI3HxYL8j
2rsJO/Ce0nj6MkimKxcB5TLr1oZ73FFAwcsrBRc4g1tHU4qaWlHCrXMxjR39cPdG
+ZGPxoCc+5A8Mf8rjLzgf23D4Tq7l/vef+o0uGh2YJTWOhFfbEPBrhVjbwgbMKdI
UgrCwYcUjAymotkGsZm9dsbrmgV6d3bB7ma5QlS5Eykrj4IaN2V538bi8ZpUxrgd
56CSe7rM6dj5k05d38Q4Z/mjZf4Ggr99vdEdK7a1ENjDyMpspgWpz3dE3Evm/GdP
hwSvOQEfyKFfGNGIPHsEWAmiqAuim+zPMqBATiJBq4NPvBraMyUAziWYfLqJ3IjR
wF6L3PtxPrB7vjniDE8ryLr2KyyJZz+wczryds+gNpYoDL1kZ2ImTjKR4hVI0ASL
OCWN7M3vX8i53n4fBLMCQDHLVBrbTnI8rK7KJqjqjPWk+6O4tnG2M27RYwEV7OX1
GLPfHnHEtPuGf/0hqV3mhfWQqyaCwSZqT1IMijF80BJ8QpX/5AWdA6/D6uCaJ2ej
v6iCXzTwmsnkNDukdhyZ5Fsc4j0fx12nv4L5PEfUbUxQB+ogMbIDdCamuc/r03o7
bxHuosKN3Iw1psVIcQOBlW1ZLS2swVKjXUzRMAWOHAmw4yGphWbCsk75J0T70QoM
ZM3sKvrRbrqgFtxwCiEqktp7reKfX8ap+lQ4VLvz0vCGajGUtVtpDhzD/fGk+07I
fo2Ei8kmqSyjczHrAlC7IZbdDqPKy10t5jdsDpqMlxHug74ROPKmgMKDrY5mp4wZ
hWXwDF0nZ8Bjk8Qkeq6+bsVt6Hx7vsKd9T9zUwsUE19TXfRMNUT6YZ9/VQd95kD5
yGQJkq8alN1UDm2S3vY1iB2gn7Beu93Dl8s9Yjvbi1l/F0bEXQBrZ/1CTyMwnWnT
pdjEcmUb5sAq3DD1ityrO0J31UdkdiQeVh34+1zF/ePVGeX2B77VmO79hiO5W0j8
JkcFDNeg65vw8KP+Rae3q76sYU7rpXdDpCO6WD40Q4bSJ4g/AvDGP2jMOMqRyO49
xSc1Jia3MsgKYPaoXtPoQi3+hJ6cPlgIWAlV89BCmDi0dWpDeK2ozqrdP4tPnSyZ
V7X+A1MRHEAnzfLJrPoIdwP151OgVJ41G5W/LmJnJpkijtsBZ2xgqxOTzkEmrtlh
0OwPZUusEP0Wb9bjmayR4me+Qp1PoyB+vJRi9G8YTpgILe0sM5Eddoaz/EHg5wh5
0+4P/u8BtUo2jN1AuaysZ9tJ5N44PwyC1eGGaw8f+r5BAe+Dq+t/ENElZBZ7+m+7
OxF4o2PKOvNQ/HZMVdJNQZyYRPxH1QMPS55JkpgkvbhqmX/uLa3k5tSV4BE/A5Qc
ugNY37sfL2NLObylYbDaHIgAsJSW0+T8WOG7h2cKMcDQMY22C7g+3E2gvAULK0zF
YHNT8nbRSibScSh/MqrMv1LGtvJXmbnPa1ZQ4wg9g/RKYdRVZa4Sf34dekcXE3x6
dNxa4bN9h/PImFwuPbTye5SwHEZ0XwKxL2FUA85VfZzRobLvmVMR+74K3n/ElVsi
dEJQVNwIVo/hqWIc9xfWLh26VVO0drtZzPkzJ4JonECX+a/1m00qSJPIa4k/a2zG
+xL7KTXcHfjybd9C0rXvEo/BUIJ4iu1r4F2ez9/zNzlW30Xqd+EIcDZEKoBPAWJ+
0j731d3Zq6G8QWTnZL5laAfb2v6fd2SSCL6hTaYjXiaE0QS+4eIATfAxIXv3aSvZ
OMv3p32qtQrBk//3iBpFiO7hGSHsaXskOEhAj3eJaLFA3JBMmBKu/oLWa7uZiIyK
ngWpBQddFFg06HEc2ZIBC4C2UpRQ7NdhBzflKvJUR+iVwAWTqfgAo90b7Vk1FL/f
1tD4CcTncdzKFLF2yLA6w8y0cr7WwXG6mejHlgwrDs8LQRyvCq9ky/joRWvbzjCn
AAFFmIdJtQN2922xJNG/S3wiQup0gFIjNLV8m0OVJK451cTNnhNhU81AOgON4/gr
y+3nSisUrSCypO5egY9gxWbXvs3uVw3NCGE4Bs3YW5cB9qsAXMfLW5D68Rdf5Bpv
8UKObRqHaix/ipvCWvV3beXB3dkUHh2gjU5ngibLqdNypJyJOWUCesIsxD9voDVM
2jlzeFGYzHDE6VE9/vPewKUJK818V92F7nXrjoLDn9rV6Ih0/t8J8TU024UZexYu
BzYYtbd7exhbxTSgKDeYabNDsFS2sIckGqgBpEp1N/tokpkgcW0Yq4Dz2geSoINO
3v+9jeCqOkE135s0uE3ovmezGYk7VA8iJ2rRq9Q2NFtXlpBR41cUcW/0enwHFyx2
F7wP5XRvTAD5VVsw+dYOCGKa5fl7DWusM8pjJ+GUdn4JnkAwKPc4pI2r03FQzMWK
jIkKaOvd/BVN7oZzXTLhnkK8rjNxgsY1kSkp55BCTWjtyu3thq9cYk6BDY7S+5nu
4nMS6Si4/F8ItjLH7aLn33GScseWJpTDV9syi+6lx+g4nUutRseBX5G/7JbLg0x/
DqHEJWHsertGv7ao+zoNitJhAUbVvst7X591oZr7J81Yr23lf6M8WLx3EeRLtFWv
NwLWAxOa4gHk8IwZ/Rb8egB66ydjhSJ02mm81DY21iVKc3uRcSmytkVEnnF0vl7r
2LyKvV91S6jCyTHD3Yt+TDO5dtSJLeomlhLUxG08bBO3SQTkWlZoXFZRaXwJXsdn
AfeeGDHILvQMCdYWWpeFjwvSQkrHkY19x1FHiJGyuZ5V/qcXR0sOteFeQ0JQ7uTe
5P9wVaZWDYo6Sa2HChGhBktWOokRfVzEAceOHPlAql04cM9Ks5SouUJlRHattVDD
UrBp4ttSK0KaR0ldvxVmsaGkIUKPcOHCfxjpIuhTNJDrs/b77YH3Jy7Jg64uzVn/
UEbZ6Vln6FjU7/3Zwa/HvcJ+bj25zogJ3qcExQGoGRxPaMOZwLIymxGayMVM65Dj
gtbe+EactHMSb8628+CrE8Kb+tBNq7IzAtux0j0Gc5JWqMg8ryyW/yf2CJF11/Ru
BGfg29jXYUAWXpqccvsE+PH82WPVI8xueUs8llXIMYY1EBBMmgLtE8RqOBkE6QBR
41vohjoZDvJj/ZQwHlnmhWbm07H0YCM1GmIXX7bvJT2YzZj8vTQqLOW2NUZCifay
TQD1UfRHPhF63TLOfvEH8hgpkJQhBhoO5+TxIN7TfPnjNRCSlWLkIfQXFvFW/i3D
BMLULc8haqfiGl1/mXQK/aNIC022DkFrjiQBvIyLJE9xWiLoFj1nroptvZBoBASp
DIKocWAmEyHEuPtLCueFs1TbPph/9gjE+3p2IiBJUeV3oFDSuDdmZJIMPhxSSHge
MWctr8cfSXdlArADYnzYGZQU8VZRwgVeirTDJgI2sshMP8UdwDJ8Fe0XLvcJM4nw
xbenIG2g0h7lllC2JnqYGPHlaKjSkbbdWoJmowUCr8pvcw23L/zAxzsOfIxyoKC7
bTOAbnpQeqMdUysGc41wGJ1r2aea5A3ltYLJRUMYkc/y4uBddJ95fKV/aj3oLYfD
BhMpJk6ywxTm2ZkQDeVBjCWZsP7VI5BgLRYdGoJqxHmubZrE4GJZTjDrDoWeYclX
B49rOjzdw31XMeNWFUa1Vlo/28jCZ5FLE8ZXhkoWwuSout1vGlf4cCBnUSAR6Ezd
uKehvYQYaP9J1bTi5YPzNgVTVIueBX+DNgKIc0F+YTz0N9HBz/WjMxFSIXrHS2DC
wA2Yd7dx4c6MgJUaLyTIAQPjRXZ/2BjVdrE0ZFk98hoIFWqKon3DdrwSJpciWQgA
biJS7TcdvrLYMO7TQhPABlHbxXWc+RwNu3vzz3M8yF2ruVC6dSkt8zgkkrlpiLCK
B/FRKlFsZgaF2XQxvJGM53div5zb37wa0mJa7H8+vvtQPl/LhCApyDcYhBgGeEoU
aFLOl7mOPJmgLLKIaAvB37XUJt9oc0lKMC1QjdOVChx4qx37JCugSzkRrcxrNB7T
nYMoCjIBvFhKElnfvqxF3zy97iC6QId0sjCMQI7rW+VCidryfTGTwxUIYpuAChiY
1l7zfWAREfPoKmYeunqIAAyGt8sVIaS8PPJP/RnOWKgtpEYJSJI7yfI5RWENHKVN
O0ZW/Wbz2/jrjE9+S2DgX4eM2psbFLiIy/nYNW4M4K/t57QkxqHmoLd28aBamKn3
RSZhQRnPCffV64jJjxEJdCsCqofSDpn7nlc1+JIFpaHLvYQutjWjtBz69jvqzvsb
m/G8fmVmA/dKedrB28fOPPBziHxpEcLaZv78gD3ARx8T1Vnw9+S3NzDgNH/ErzQG
QXLzKxSF2M2jTVQI8uhgMlcm/SjDOCtT3EQmXlB50hmAch/BYdasCdWGH/5XT4+Z
NGpJaEKV8ex+JxR8UO5xoqfDxRDJlATFP4FzJSBkuIlktksAiX+7lREeIul337hw
YHUEkqmn5Zlq6MLdbJmWtuiwefIUUI6ji5rD0Uz9z57sPhfP+L+WIXvXHzpVwl4Z
zaAz6IvwZ98Hb8cZO4KymlA6I/RFYEWmvJYYs/4RQTCopqJG8ZC+aBgAVSEfzLf2
7nQNxwb9a5e22SEiUKY77FCKFZG9omhas/LS3PcLtWONkMR4YhOZq8aMKPqD6vcf
TRHxYvzAmZE1uCjL2NcgaGSLkqi4tq2vwgvTO+gxQZQIIXMzSGa38UdDp3uXEbN4
Se2zEt3HGuscrmFKoLoF2WzLmwSGheCiMf+q/acObbGHIWh4CLPFCzd14gcn7fS1
EW7on0hNbSPEduWRbPxrS5cF6Vl18OIPGZl3tVbNsONtzhfZHjlPTutlOC9wsrR9
OCLWRhWodNktUX1+/4zPeMAG0FEp1B6xciEI7QSS8wbDPfn0/TU+GXQgZBkL6te+
WiLWA20e3G8vvWUEeE950UG2EtcFhKPnAQuGwnqOun2dFGBEogKmr7Ruomb2MVfI
+J4g7vSSIxI8JNfArWQ4x17EyTh5+ZAHuIyUotQpKPFpNcrpWwWv6BmLWCTePwMY
1dcgIHxmLqRTGbS5RrUiN7ThMHEuGeCqZLJGc6U5SNpjPLnlneaC1elcSR6Bj2VS
jrNvDkMZQ3SUW/giv/yPCaUm2BJXsQ+mAgYaUYUlXNdP5v61JR8NOqUzgGV+k0u4
InEdLmF4vnW8xLUSSKVrK7Ffg3IYqqI5vLSFQI1ewjo85WXnc8/xITmU0zFLZdas
7DIjmdDBrqPdD6zGm6U06F2tgtwxaPbF/yzUILUN0e5aur+lGqx0POpySDdAFLYV
Qj7n3Ocx1J606CJvTSwgxlipYVwU7dxgHJiZBk5ku2tfz0sh9E3eLrXOYYL7/24w
BkpPytDqDRr55NAdZ+AZR+6ixnwdICPfM/r5uprTx29Zddf1lQmHBd12Hlsjgi9b
2lsRYYVe9M2vsupAgX9BhYdQssZvl08xr4ONRDH+1cNkgMaAsK0WiLCZZet4AYWA
2wt40ygWOTHc3xVYaGd3D+W19flMZ0GrC0m/zJ6k2wW/7OFdrY/S5CFr8S0jAsIt
+mdtAZr9vYLTWOE6WDh4NNFcWdZz8XwHmiprGLc3v44/JsBWwxgyD7vRWmkiXjuS
3UIM8mUNB8ofaFH+3ItbmpUHXHw5+eKmrRforFgQAvfRtPc0BYxqgBLZdqXx+dNw
k6nkZ61roDVSF5Xk0Tc50gV7sBXf1DRo3+D1YR+E82CIMsRk18OJdMUI3yw+ysBI
dhyIIiu83MjysvnEVHYObGV3RP0BpBn5c3jFGg5h5b8y7y209ImFD/4dknhb96x3
/nlw41SbejLa74dtaWSwGICHcE3iL7rG9TZrav+OvIChHUBkaXZaU+t4XQHqvQiw
4BtkpKeVcJRBDCYNd51Tpmk8UBsoC+tWXhFm0o0EiUWjEIzhZ69g/FOFLuyj1QAA
/1oPDMtKGUEUR3qsAml9eolziV3URu9/p5Cmax+Tmh8gU5HBHA1sZxeqDvz0PjA+
Wb7O/D/2e8vZ5cJRyp3ZLXcgOfLZarffRQZmSt65+5JZt4oBLt2sKbz6q1nUfHFK
ci8BwMEt2jUpjNx0rJBwJenVqNGayKrKxjfGDMaRQhmVYicOtYtMCKDRYOY8vU43
CUHv1ElndBOdaSinozROshD8pP9tJ53qIQyMCtT7Oh53+bp14ZUpemCqrK/OzQ2q
JoJl8CBGfsakdubkhtcXXt4p2mLGUa3sw6QF9A0M1JPbBsFXBkgrh3xJ4Ntc4ZEn
Dl9RCd/qdnp8BUjnRunU2ZVL+7KEOzpoShE/k/Orh8AmVCuyyQpWlG6zZrM6OW+9
7qSxi2MhUh29dLnPVvjF4pWJPlWzEqqmwA+RWU1ltIxmtTua49z3TqaYkttYj01F
YPvGNp5OVgrph70AV0DHYGEAUSvsdYiHpYW+FhcwSMKgFdJAX/+MRw9g3ZOZAB4B
iJ3g+XMo7zpeFUvB57hgfdooEZUKKlUQUID/8Wm+8WyWK4bu1R7CsaGvwYb1SugR
6Sn3SoxhoA06bPHZYawr7x+C3+3/Ix4arMewj+CPgjWgqrBt4yfHctEdZCOZ5upd
CjyEAfPSJlKtxd/aRG5O8aomCNxmzDvb2Fyg/iv/L98aVSZ3uCbZl2qyAWzq+VQX
u/DUgNVl3eTIN9SlLG/UPKrevkAbJYEROfl3zPzke9GeNGU8Rr7uuI++U66sV1wS
v0GxDwX4yz4ne/OynePg6MrVe7f7W0cUeKZUXtHtAHzkveAxMp2ZL/GQ8oxUm2Zj
KUkhBapnpfPHOsDXHhMoi+xIzY72Jr+3vNPEnspJdBt/b9wXL0Go/7OMH3CuMaxo
xYm37ZDzJAd0MjHjPRuJj0aBqXWyoHIECSfHOtSQagdDHdEgAGUeS9vK0TOXW+/m
wsQcAFup24EVo5s9lXzRd+7C1FQLOAy4v1nkVE0sYi4eimuv6XeROxcnKoTGC9vz
CgN4wgW5sD3N2uyysqXI9eVskYBZLZoxI/XefRDmkNbGD1SuyulRv4nMk2drFpw5
c5CW0aCJ2bDO8wvhWLY4OllIlRCqDQMgW8yrj6W3llHjvRhIth0GaCPh3XOgeyHV
7rwVI8GcWHieh8LeviT/SHeB6vkrztPKbPCocTk9BUvDfyrJY/U2kqFmRw7h6VZB
pgrz1L1kkWtBxHqDDEw5C1Vmehqnu1+9oRgX0FhHLfJVVbUH+8rlD28YVNffV+k1
lqx3XflSqTGMRVtY2st4s5Yjds7LNdbl96A0CAZHroEjj4a52JAQGVZ9ljISx02k
f7jeQ+p/mgY2SKcBIcSujlqKMGur7w4bEeOSLCcgqnEKScIGcywhrTThA/btHUu5
vtHDMBFN3pD0cwma6jfHblGh+lyliKEi4GmbOD86xK+XC0PtXFpLOala23rOkaLN
kMgrYEiksUiEtSZX37UMJ1Owas11p/VYlEYUktEOIj0//KmOXygrBJvMSz9IkhD/
nc0mpx0a1AM7iB5mnvqmN86ZqZYHGW7qheQDgvTSd5Iqlyf5j2OTmHMLC4ycu1VJ
ERA28gC79PVWpb+en7zWg9P/LX4xOpv7MmooXyH4Z1P5YRHnH0erq+/2gEhzaPsm
CFJ0UMKChi+GD3WivrbV5VF/soMkkXHk/IN9OF0ZJNz1VoljLWp7fTPx36JitIVc
IbQ+CscumbuOTigurStst/ovehYGbHZ+7iGyG6K84bQn5fbYfWg3pCXZ9Qp8eHmd
LJcNMH5wvTQSsfXxnHnp5GrDPpP/VMV8TriOy28vcRuLdJLXmQfwgc+lwBuSmIqC
fJM4cR5sMXXZPxsXoTg0dsQJVIdbmi3HWzcBE1frjL+W8fksd/CgwQTDMpApY4Rl
yUoSPaGpBhHW8+E9Z7eA+O1W8X3A1rH6I4npAWGntRtzVvKtQ7MJn4CYf4zBx58M
kqUKqSlyooX7FnaMn6dZwDsIgstFIiJejr3UVEG4lmdBJFTTAsKfmT1x2TCUsyxw
M3mfwrIdo6jVxhZVneM+24rROZNiU4LlLzBWZhx1dlKsAHXimrwgbDfUXUbzZYCZ
N5qjc+IVkwfDDws8O3jT4nuZLBzq+Ix2t+HbdlicOylzJxdTLqu9t8w0aCADaEBT
3CzDUBcXW2OqO4jddMYpGAg58/ni0tgnDsDyw54QQT6YUWcZN9ZPoMHy62mHUasv
8uoo2mXT7+TpPnnzwwdj3pazaBKCzdvJ5gyVTmczFktFgTelM8FHykXsFdgCIY/+
9I5qVpg1q/AI7DNQYZvexdBYB5u5ndFFwAad5DuVwGKVES18NK4ZNxSS5Sn6r5D3
dGadYlAtFPeUBC0oomxOuXpSVUyPpAsSsrZEXeuAlT67zHS6+KeOui4soGzTq5UD
NztkdwHPqjo9pfjHut+AOnnXT9eEc44DdsmZj+dZzzLuCP1yOhYtsW7Nrq89cmbc
UEY7CDJT9svkWCcvOJiuo+r00h4DIG9Oi3JWMKNQR4Dd5cKCD4NAkbwCc/4q1B/x
DCs06VdDT8nzj1LHnCiuPOrzMjMtbEcUn+OhFStMDh/SDb4AR+2JyU3MLEo+c2hd
2fziE/t6lmpvqM4y87WhXmuJPlUw+K/5/dOV9NrwBdJ3lo4z/tAj2yePsHeBWqiu
RdIavKToWbxCDcqUblmTEPxsH4i9tWF3bcbeV3tqo10KmlMXODuhcGK8wOtrIXIJ
Pl8zTwCoYGV/uiU/C0YrL2L618B8eviDJqh6KpIjluMT+wxPzPpmsMjw91Ws59LO
aNEsUUvJP0DjE1jCm6P4DueSF8CJmvmb3Ry13tifPNNAgxIoDz6XhemZx3+XwpnF
B80z2izfq0VnIsbjjtrNILrdR2TTkTbc02vQyodHvO+MC5uz5aopnMIHheprQMBW
qgKLLBFPyucblNZdsgwjx4S4fix9pyEoAdDNMC6ByGMcv6avLVw2gCAS+46tcjBp
rkqK9sRpIV0sR1wb1e0gTHT8RTEgzBevWfYFdYwoumY+Rk1G3pQYz2sjew6lxbsP
XREx1fFiNof/JskUiS2Vis5uMQtvwqRJ9cnadPfVADYXxwkqVl3ZrH4kG/MUWh+6
wcRPBlIO5U7EByccKI9YeJdRQ51d5N9Z/iJTL5NdGXnABuD9+2VpkUVrt9/v+5gc
4F+XN1uaI1LArPKd9f9GUTDAhVe4O69Mpdj9Snw8VYiklV+pFtm2MJbM1VxJEZwy
nKezGDfMe8M0ZFDyeJWGphib7+ddvizDpD/A49++siunSJI9qZWE56FpJtyX0vQK
aF9w5J4uixz2ogagWJtcsN8pWYqipK88NWLVSbe8zlGN7Z+/tPP2mmLKLzq15P5/
8c3w0Ds3XXpussjVQRk/unNUhwcSSRZyqgkvRhz7HU3mFsaCMMOKzdvVpt9VN3tr
35Y4dvYa1epwzryd46HQ/GvbkAylPQ/ExTrMCXcFVFi+acZ3loyrRvFok3jGlkM/
uAwli15msCTEj6j8jUqkGb6u4z64L+m4EnEmdEFuYmX4E7v02fsERqU4MfvWlWes
tcD2VVLEi0zT3ErtiLZAUPgxYHmGbFK3ObCQoAwwemCQ7IwWLFw3qU9PoGPx92hc
IoeSJbn8GUMud4gOoBA+TRmFOSDwOrZQYcgH9hcCB2GUYa6keRvAD0fuIcn8DqsX
hAaiuc1vVuh3qzpSy5fYZReslydSI7XhXVT/szOiGg1ab0lx9LT97M5L7NbJvpPp
H3wlY1ByrUdJD5YNHv9OffaLYAyx/NZj3JO2SW4DroXAyAmai18vK2+U2jQrjjmx
mBRFctfjXr9q1bA0LETo8ys7aMpzjVgm5xWH8jCFkve/YKBMD2qNq2QZltdk0LqM
pzSWc8py6750udDTrk6XaxcjDTwemNNCvvShr7Ge6TY8McL+Lt8hQbtNuePIr4MK
cRxgg5m26Q4NDqh3kIJ4Zs4uVU/4D0+BLsyvKO7yg388Q7OEEH3aTg/eJTSKfdso
dC7YAZYEPujPRutZ3ZFU0CJf+k5ZPaHi1kzkOd8PXTJUsnJ8DGKNpwH+933CVvDI
vjjwAt4KF+XSROXOYQuAflGgeb6xH7XeQW8GdbcdOCUgUM1YazXbu94Qfg1J0ijU
alQ02HMvJAQBsyJWo7CBvuxZiibjDbLATZ7NKW/eR96uqgLc/tfkkGxL5zX2B18a
iTRxKAfW7ULRpaiy3+OJPFKPHmca5GN1AtgiEd8E8WEQ2wqL5SawqOOknwrgk9f8
PyL96dC5x9e5QXZfXbS5r4dz5o/qc8OVAuPvV5pawqIZxLqCH67leivAaydCXrOf
zkQ8Y/0ziweqacP1PZUNLlGgIsgZbvojJKD+jpC1jenhp1g5iErj0hwTjI/8R4EW
qFnzJ0BaJytZbPRzk5VxuYXPVYxwc8DHjSZfrq5QgyIqaLzBnoeBiWT5wFu/dh2B
OzMT3PYQR15y7Otm5hErJHcnoKQaMo/05a/0ZFvg6iM5BRMuEYzHc+oWoooika91
Ss6aCy3l2tkaLHOKjJToAiTZCAJUZNA3s8IsWdmIaPt/KHWp8WNKFGfqgOi3nwRG
MXieCQnKlmRwLJsTHUmF/YtCkZgUf6vLO9w7hh8aWCfmyslIQZNBGdHsIxtlk3fs
BkmBInz5kbAJiE4QfiJHOmNMMaUsu7KGCHOIog7Yvua4W513v4jO9HuBwLIlZ+go
aiArSOPu57+zzeLUYW+eBuc2kuqbS2Cm7hYaJDWfoPFpGxrRDwAFGmsk/P1OayFx
PokzVS091LC5nPh5MO/PCPhDsEQyzAA30wagdH+t6uXcqwWDXKVX/CqmiL9FNV4Y
dsk30/E1cLLVX35HO+Yfm+UfSAL8SpNBD0ThPXmEHTUBvqa9HFaWMnAkWvOFJtHX
JpmTEYmiiHvH/TQopMbW/D1+DInwTS8KVwVTYVYNDvIrdtnQt+OJhlYDaiAtaiHc
66SknS7sfSvZ65rA2nTsqwIYBlVY2hs03WBbx2kt6/ovk99kufshkXSauAaS2OAT
xOV87ow2GfS8Pp8VuSTj/nolJhMgUuoM4ix6ZZJtVQqaUNJ09xnvbOCbdOg2pL72
/5apdDBjiS2sDjbPFWdF3OKr2gWm9AFNksDLnWc3N1DRh6R4k3hupwbWHGsdbeuI
kpcydAfEnqxS4Ht2anOXe5mbY41W5/sxXIYy6jcagHhgfdTEGNw/+3DcoRlg/vAa
FPtL1JABotRjK01KKEkr1ZZAFgVW32OgFtIXf6VBpRua9qWRLrNzcSHJ1j8qnZFX
95TY6jU2l0foswa8OAd0z3WW7FN3ZwIRXffThdnkxtuvhutKMZpIxCn2jQSyyJ99
/nm/CL5TKVOKIQsEe5m6CmGaNOr6jxHUyDOfPsMqCzv42o0/bhycGfr9SS5G2N50
F4js01YYanxhsjQzaA1dFL5H/PCp5qQezSrG+9gVjV56OSD9OjMG/P+fPXgJ4Lzf
MOgtiGaJ0viMt5QW93+UeXx2eIdlaWdi1U/9Em/C80w4CbZ/AV+fynPkWk9qO29x
VzZKf67LcC+cG9upN/KAjHhAB4lXLlgveqQ2NsQellTT979jLjC38fFqLINJAcem
K6R/qq+yrBrfSHDkoH704+7B6ZnWJ4gQcORzZsSEChfLbtsK34cWgi37tjX9yEma
KQnptpXZ3cUrcINgG6fUAKbS8G3nHL/LBUBOm/38tmednDJf1rDF5ZyzD4dTrkol
rZ9HItT5ltmBuoRo4rWk6dH6d+hXdquOQiulMT8MDmhX5lHtud7zxHLHTFc4qb6q
BNjsrw074Gy2lJKPz9EsMW8Nzdi7zVCc91c71Vt2KfdKpwHj6xDqUYbKFyE75FXb
VRPKED4NuGliIYIwGqjSlfM5i3nInFadSs2D/JmquUAUieN9JM5rQK2dhPb2glLu
8Hxpdf4t3kMyuISWzmPyjY3Crh3z7L9+OuKwzsB9aTQwZafHNQQ6gfIg2dgp29MK
QNhRA3hJog3/qpGczV3KJBCtY9Wj6dF65OdbbTJvmh1/qhAHtNTeuPg7Sh5Fnwyy
nrvCUrVPW7w+gprCLOTvHwVpjRynhjReqFcwoM2Znx9PMWeD8Mm40SrvimCh3KqF
+QEuWcgV2jX955frJiYGp7BVc6+SccU/qnW911WtOnY+zmJ2oA6I3ne+1vCTAZLt
kvrZOv4GCouOVxMuuo1R7MU0rcXEu2C2LF9TBy7co4ruLdcQeZ48sNA1tuY57NfT
/SLHqMS6YKuMhgV9clu5phgtpk18PuCZO6tqGhB3sDzuvRgY+LefBYn1WMTs+Y9u
65SO4aOjV+y7jFCfYKW8oM++1YnXKLzfijGmpQXjVlvVVgn3hj+oVeQVtHAYtlfC
qq5Rhz7B5GlKjXBvtPxUxvcV7A1eR7dGFSzHffSt50YMd93YDDSqgk9Yd9WWGPjz
+V7sTtmHOOdvcqI8rc89KYnFc/x9fvif4Rk2WIE9afU3J0xJZof5LoLJJSePOvBS
iO1q62mmsh3tBX+2ALouhOfqqFiH7GuD+ghMSNIO8TfduBNs/6cm48nWw4CI3XMv
E3peF6f+Gvdv1vlbQxEV0MfIwCPRvznWoPBOQtXtPN8Cm6GNPrLABPr6kT5gnxDP
tsU88v8iGDHQsXgSdOe2g30jgad10M0lAdxKRWmn2ZfbwMzdNhwEqyzUzono0QVh
WaC9KisF6E5VQFgbREvNmolkrcCHgQ/THtVgHVgdPvIUWipoGkxFsV3CYnM7q/m2
dopF2ohKjRWBSnoc+nAnYtwCRgKeS7qMf4FQ/XQkMU4y3xxhNiKS0PiMAUJl79mw
mIhQ4vTCQqOHf88e2MJTmKQcoF2IcEHu4zkkFKCZ6rkPIpPco2WV8EkcOnrH544W
jZzQ7d+7qd1gI9FskhqOZ73rng8lOd3cJtIloh809Iog9moFjt4pnwGsLswNAGdD
m2WrknO/uNAXVxf0Blr+gzZFpX2osmZaDnrYTULU4U2iwKDx9sYqzbNM3bjdDeix
kkHHQr5H8ypo6pl81rKxVcAAbiH72rqgLNkQ1SiYzID9dp0M4ZlgGfWMtI9rTRcK
2qhGEQGYc+NTINmUJyS/2wPQvEeGYEexXSBZQKgaQF5sGUEzZ0hVabciZ0mSHAji
qjhC0lcFeflyOOIMqv1pSUSGhMMihuRBTY7XfwPXLfh2FF7sMwiRvZMvsMhvm+qs
3vj176Ks9EexbHAIKP8XpSR++YNVAuP+VnGvl3EeR4w3lOSQQAEC7WsYPhwJWMwj
QIYAi2wddpCmGrcDg3GWWFyUnt0W6SKgLg/hnDFwpRVndVKKJ+DTBSymA6N42/s7
sGjToB6dJThvzB7b92XFy8DZDMqFtu2VlnCdrRprt/LVD9OU9ruQ2B3O6Q6NK70p
yMO6XMgMTiIUedLUayLNKi6m2J4Kj0p9dx8l1xk7iscG2cjKvygD/UnCAY9aroB+
wq4QYls5wNaswiPwlinzsGeYi6i38aqY+HOBqzs2HJoRFBre5zXRX3huYYFWogPF
tPJGLdA84PupDeSnTOVCNxtY6ZXJ2W8MnxtxGsdSrhw5Elei4mrtKLBmz5KFh8tt
8+cQ1s30uSCSGoV3J4snuRtRuedD/OcQ0V5Ff+7cEG5C63cxplJBDuoICeVpwFCe
10E9RYcm72wecf8wxmdu0caijRMiDCiHxyezBcyWOuNhTyH8GP3szq4XVPqbXL9Z
bmEpXBkwKzrZH9pqvZn2NzSPuwWQYQvgf+yNLnfyC9KZ514Qs8Vx2tWTAGvnxknX
l2NPHx6GJmSuaocfwvUIo07QT7Zaje8auYT563L7i0QC3Tee7ytSysQnHCcraezm
ZMjhulg7k9AS3/u6uIm51utJlfW74jv3MgFZ/VA+j9RBrpNKp9Yvg1c0uMN7b+eY
SnPZ/4XfIoGWXvT8+aoQ6f14OPceTXtroczKdTYBG15jhy/s+sQy5lPQ6J1ONOmp
CwIjZAEnQye6FOIUl8nQ69P8qha2kxd2NmT16F6PrkI6TfGmGHMu+qbTYbr6tak6
18RKxqyNwoxPqb+hvBUT5heZsJ3Rs4YE8SRaKjozOISFPEPZEYXi9p6DqASwYQNE
fQkIEEOtfgar94+mZ8++8afbGw5y3SGNu/TwWzd9zsuYpJ6bYKda6zwQsKJHpv0N
ip6uouCAqXICBiV7xGncQt+fPIKxwopA9tVLCqYPl7cMvnLOSllawrfn7twQReSy
x+pL7vYIGHKYHsm7yY6qiLrzrIyBDWhCASYwEumO8mx+T9o5R7POck56pIY8aKjN
Nt/h0bWkXpZjv71BaufCfnUQD9brdzR0mK2fO0S9NDx7veQy9IXZPRMz2/4p/Tfs
+PM+qIBX615u0YT1lk5Zfy/QV7ljypCYGLk0bhpcw8v3V1wYl19oRVoRpGP9/7Ng
O0954bSlMC9IjpG2YJz9GHGdCa8QJCrSUBPrvWONj+B9grqrjX6rp6MTl9bp/l9y
5FYJmtGYhowpi/rwzPvgPQza/znV4egYai0wLqQ3wWTt1jULWN5mMvHs6fNS/DGa
QlTyHhUlp00KybXHQJo8quZsSox7DIZvsYoUNA1CKkomuorNZEfL0hlPBPesEDFh
rAC/HaNTxnI34yFq60wyr0zR5gnKSsNs/KCuXh3aRTCDKFdJptPhy4OxaV7oOmUZ
nwzDnWEfx9cE+qO9y759ELF8/yVIOW98/X/fY2vGPPdLz7KhFvTYxV+bZB33T3VG
FYDbJm5aLR3GzzXZvXKfAMwJws3Ujp4R4DKZSLaQ8m5YLT+wfrOTgqVJ+++l9EMu
z8oUOtF8/3nVV1dvuN/yBEry5X7QQGRX1pqiWnKm8S2ZCsQyMGbC+0iCJFP4G+xa
fvxA7hNxD8Z6iYEew7lUoHF8IG2H/TCkCeAbKmriOF0BMuvtLx6lWE5gpfG972kB
NBB536YzBOMsz2xTWOMm9We/WXyKvTk9AWBtv82F8rICnGiI1zZ+Tl7j8HakKxVm
4SVRglKesJCIbFjS5h3s8i1PWJQKOrjLU89hjbvSadpbSwmhqdn0kKrqC1ioJFJ3
G79DB8Dnt3/GTFXmEYImDkGz/Cl39K/YzM8NxLcDl4LUxnKdgGLxNf1mA0AXbiSY
i5I7r0KBUp8cMapPERW9isLd8ELBE4ka7G+Nbo3g3VroDcppUHPp8dKWTnVaE/PG
UC2oCXKIEhgMqnCmA4JzcF3aonJBuBit+dPmWFiR3yqLCpsb/ADicvldQZB2glXo
DLhbyPf+NiVZZ2Rjse/JIGG9saDYDTTfQEpVHY5tYQfA44nynZWHV7fvpVPCKdfh
0nq2RWQDrRHcMbKLYpcSSCG2aqzRP2tM/xx9gxWv9yIvH1+cU+Xh/1Jh+d5bXo3Z
6Ljswx1ZqhgTZG0ZTZYjl8TCZGruyZ/SiINEBlRyYuekIqmzLAhWYUwp3rrJDAk9
WOqq0hsSXSMTz124OWee3ST5XaMV14m0ZB90CBTOtXjb5ABZLPP7399kQ9FyVgMV
ktfTbaZ1V3Yj+Jln24cCJSgP171/eHJBaAzUvhO6J9VycDwJBXbQvg1zNle0+zz0
3jIJAJJLDaQQ7EcKRErIJ77v6d4jOJTtwu6U0TZhlajCP6pgLIm1+hJ7m6d96A2L
AcbzKeBujEynGii3D7Vc2bBmfkJyk1dxrb/JqyS0sLl7+Se2930+Xc3KUK6U+jwg
doxZacji5PUPGsVwYj1xfw7d6BrCGmuuP59dlnQke1I+uujnf8VyWLRlhRRR7qVp
b8eRYewTpkSeMlKBSaBvpWsgOEckdBdP3r8P0y2Umiby2DdSEolK72MWToWryLA+
Wy/nCqMYqacZotxnwOhasAE7/r0yuTYr64j4ac0vdhHq202EBHpprkk5bxapLKj6
4kizaE99FxmS5SLte1RW/r4DnYl4wwhE/aYEE+PzRxQwcFe5DytmMNM1Z0TbtyZA
dsMbqZI93qb5WpeFj2N4fgaAy5moVDjx2VJsRpIT3bLTZ1K/7FAvw49mDI5itjUi
fRUC+Khi3gj/NbHp4Dn58hxESbamTOSjM946ZOnj2fqQ4BHLB5t2UStRzOBfBYad
ObLjP+eVghPyKV7AAFQaI8bIeyYoj9xsjni8hHcqV7F6egMrnOzXgiOX+URbEPiV
IZRHDcl8Jcl6P7U+lw+MWKh1vKUMW/QoHahzXfbB8ay22DsjGPHGwjMv1u+dr74K
VaYi8GR3mI35FDrMgsyLU3m3ZKUUvDPMoT8uE/tLcTYo5Ji//qVoUApZFhyHjPKV
MGdhDEkNpQOtyEWoctKj9SHSoluoI7Hu/MndfuUNWOEeQcgU7nzsLrHCfrPtAwbE
dtDj3pz1OOst3lkgEM+akDqfTUM/E4tI5RldiwNaQzORs7HtcQdgJRtLwRAmHGTY
xOlVaRVxdbQFrLBeyB/Zeh/jNlakWlJ7uWYgEV36l5ghOmLOB+pVeytEYxPbOSDn
0Gg102GbZe2h7YpX/vuzrdkr9ERIez6En9gJGIOZKRQNCEUx+emcOXVocoH5Tors
14YD/xFuwOMRTAAzgflGvHTv7VIbYvNZFbG6R+t7paCapF1qQg8TfkC9tNgkT+ua
ldR3p2300nPHLYdJo/M3UL8NhWBvzFShyG5AnkZfjhxqQImiGs8uuOXBALhTRVIe
ajnpf504gyfFYTZksMLVgGj1Mbd8fBVUvk/1GVwV35XWNOTY5eh7rd/XJZ291Zrr
2gvcHV7DjX3srmEWf3BQX8ZbtEAiDFbVy1kkKax0qJh84xvcetjv2Kd6b6lASlCQ
BXMGngLg7Q4ad/zstWsosWhmFgwvjenbr3R8N8CW2a4IbJKUcf5v0JNjDRcbQCNo
inw1Pdnq0g0pvdCc+Wjn0qTfZnrBSE9ru14xxRTW0b50s2rvf4rdI+fr0HfVdRx7
JU3gblQgip94Capn9IZVCJP/yNHtKX7/aEm33kiMNYWEber1cS1bZChcxIwwc9Sj
VMRM6S34eMMKtko/CViacpPvljXMHjsfTNZtTdgPZqpvpJ/ZoLrn1aDT7ZromWzZ
1shlb/g9WTb0rfADcRBk2XAbAvcIKZvwJMzqix5ITnytsUEVldPGt/aV0Lydt0YP
zTmpJgB7F8n11k5J+mN2stbBDdjwO8bIOuMOTxC6rVj2FE1/fnE+ro11mriyIAHp
kWIkUlt0bysgL+exlGSk/Q3qAvpt7EDgxuXrQv0yNFUB4BkhYHOJAhtSeM81/TYU
ikQ5Am7Vks+Cdwjb3piaxcGhqPwta+cdZu8K5JvrDm9+qzDTNXSgMK/KuJ6QEWRU
egSiFOhxTtvbF0ZKhaJyWuz2owDQiBTwxu+jUJVI10BTp5MXsAbJNdaBYjfh2oRm
JlPGAXqEFa+MZalcPk7LNbz+RhUj4VCSEkmMec1yyAS/zGt18GkrUfgYemSbbvDO
yWZr6/msn/2Ty3YCVwvYobYAF0f9PCbrV0937BINF2tQoZE3uh9EksBReicBn5DL
1FgQ1v6rL34gaQXwKQziNOfZAVyS/lO0IU0Kt1HCRNZjHoXhFnoZfwCi5BoaNr+V
ul19UK4h5GmCZLVJsHZ4GppCLq5RdGkpoc4T8X/eoJ/C1RXu5E7T3a1kwZCck+lX
5GvtW20onpxINZJ45S81hudQbn2fhNs8/7e8Afi4JygNld/Rw3ny4/Qax6lw86Cn
7gjSx1F273qbKtG46kmJHfT7hel2jind6JEk+/N9onEQ4JIWyi3n5tLiOgjvWjeq
zOnSw0pAeh4UwA45b2R1RXA3cqOHQgizECQJ7Fl1Og7S14or+rRg517PqriGtJEg
PF8b9ZL97dwHZrKcWV9bBQ3t/QKIZx8efhVN+j/SCL+U7f2DjRIYGBaSJ6nu4LNy
wgchJGfsF1ACG7NszVE8oJqQKWn8RsvL+hIBxlm0J3nVH5SO2C2LOWYS0+3ai+40
0aRJHpKFcZ72YImZA6dkphif4AlvPB2FAVstJjWltUVgV+jKvcBTATmpPRuHsapJ
nu93Nrw1mXBInD11zdvjPMqZLWPh4FWfq+G2xRrnzaf/IqnyzErMIWAz4FZrBbl6
rzpgEtKKrS7BHgtX1RvQgB0y741XbfDQR3reZzb0VTl8zGlcsfwmepoV9/IlObyL
io92+TssKdPn26gn/uYYWex0tcurhjQxTw7OcuQjTuCrRwQ2iahTPr1UPCRLUSpp
sJgbQk/gU5CC908P+6FGARHSs/JfKWmXfrUwRN4u/MOFWiR4Zgy0K7w7lZVyOhnP
Kj+qjE84STD20VHhYy/l1MAgRTHmbf91Ohj8JBC1vNAgOpCxsEmsHxeGNHOS56mS
uqTnKvB6bmqQbKSB2pqbeu9Oh9XcPnimWshPIf6BcipRf2wBCgXIgctJubYzfJdp
cpK0D1su15P68eiOgSQav5axpl4NAafuoJERDTewqcd++kgggo+vRPETcZXYmwoQ
yLxJbDrQYNxOJajziBBqU6Djb7anarx6Vh4mmb67EquX9RXhnqlY89XbULkjlojd
960HH722DIS8jjyZss33Mw45yFwqEzLo5kiQn/ypL711akxEKNUioATQU5JDGl5g
XKIk46JJP8LP29eVWao3JzHT73WTGpi8joFhbO5U8VJik/VfFMv0PSpun28bnUQm
NLHIUXpnhjXWScdKEbLRQCaHiju730z/YmSQ7MDOATGvMDzmfzgxNUXQnoob3J8o
/kANK+nFiG5TUWF9FPVJFtHXqA++ZnDq8b3s6WX2Cv+0DkLmhXRUsx9b33i2g4E+
xl6Iy8IHZb3Ve1e5ODzcPYa/WxWUdJp/kry3tU+yj0tuoDbqT5gOxXmTuRRsSSvT
Td2UyL99ntykmr5jnCX/7FiwQ3M4UqmJrDLE11/GrF6PKcL+pv+0l/zKxHPscKol
pX8iNTSyoKZQlALbIOv2GoTvvMUpP45AMgEOhl//I3NWrTHRFRpB43GPiUVYAk2C
iVmtGv4PcHOk5wiKF1HnrqXdbFpbrX+oe63Q2NP9bYSpsrXDrZO1GLBYktqlfsFl
aZZA4oOwCVVRsaNGqdMawVBsdgthZ7ol/SI3l55H+3lFY0tggG4b/ZtDPEm+Xxui
3dUTA76Q7DpU0t5j5dbO7RenWNL1R2okJij8+tVFFA89GPt54JbGEKV8s7kZbxvg
iCk29DEAXUpZxoMkmlQRg2yyoLjYu/NgDK74IvtOAzls2veY4cY0+WRK+GYIKAe/
wWnFo+Qjdc9DmA+DYu5WoL2Zd2/ffRm485fvT7TFwaORkTaBUatCAZF96kwgQsDs
86pHwoBKS+/1Sdx+9HLxLdKZAYoxqz6pwBeGaQNCjxmD5wTfBshLwogZD3KxEajs
mIEld6OBHTLzpc3qYJSr5Ef8KHVhJFufQq69oD93lPeKAtA+msmsH2YnJTU9Y0J2
i5C2Pkv4LWckr3uPvRWsfWVFKJRVmbpPpzEaFvlzX1qc1CLgRtQeq1DxJ+dhmEe8
wSNHH6qRw/aQThIRJs+YGTuejLguSXJ3qA6HH+t8kLKk9H+JqwPAYaBbjut0ajHG
DKP2LX7gQSnNEJKfvOL8zmA1nFZsHATF9GtrDW7jJ4UQX0MZe/fDma6irhR6pDGi
vaCcMQ0EY9RgWsoI0jxqqt5OsYFPLKdnB4HjvOFESvTHag2aOQPEBzP5SRUuNYEg
zcl2R6IsKqii69SbKOmEblPyksHQLPwMUiAn/yhevVNHKii259OXNlqFT0xW4MFk
QwKcUP8IF8Mhxg9cveS0fpCjCG5dhXYWwzvKqjUnnx1iVw15tJNa3S7wqJbfGURC
wvwr4i0J2qNvTaphe7WsE9i1kb5ebxE1+Dwlz05yoGQ5pNEOwRVRnLTGhxIo5pVQ
+5HucGJue2vPMK68V6473nWRPEKNJkjKR1qRiYs61m6qLm0jYengnqIrlmHG6HKe
xckIhbG6F+mM8f+JQLcRMhs3GF35xo8Uc8oGjNnwyufMjPOC1JjAiuHGhA01SHp8
73O7nrT73bjM1rbU+3iMbkYMp9TXTWaeMKbwSe2wqmXanvU8OqAWPKXCVV5jFksn
dHAAn/35nXM8MqKpqjmCR+R/sXHO62pOjxB3Osqqxi4Og4dCiwhCMxKnKTTAtBfK
VjXY7z5BmGXCdmHubNfsARMHofW4+Owo1qA+nk8bM3deAqt3ulGuIpj4nQQslgjN
brkO6Oa/K+WZ8z2XqQP4RoX95Gb7j7WQR7W/WiG4dyQWEnhlqziFPuM50fAlmt7f
KsD3xIVQ22EA6tda6sJ0c0DvQ4uNgk5amHze9foJpmxZ0qaN6GSz1/s2av8B2YI5
46SAnsAy7fxBtLWR+9tboHhcBrbvRHD6I6YqNyNh+tgVjHsr7iLIjtpkZY0Wg2mm
oCPR+eUEZSbJTtLA3R2bbpxwIJ9cbePKnJbQ0qaM9u8qDtWh2l4765/Wxd11Ju/3
N9M03aVbD3cv1mcw/2DLSVfnoTj62hZfEhPMg+G2p21Hd8w+GqGlzUx9IJxVkqo4
6lOphcRmuMStspvBVCecKeLuwKRDlqGEuhWcJo4qgb6WNa8j6EUxfR0PHa37z9xb
q6oe/6dtLcjxh6t1oSRxAEONkwwSvbjopVZldJjurhJAfwhdLPYHJHdELYbHEbUG
FVhdRzY0HJcerPiFXZ3CeZt+6kFV5+cQWxZtMeXmdwCU1RjcqOZkpQdtKS13G5bX
yzQxbdpwYn16LhBU65nHaJhPmbEcVeZkvDBfGnR8gq4oIRvXXqHg1Bxtdo9DZkCt
+6C+LmgMp4mZ7nugv3PFhPsHzTdGoNHxbIM64sm+WkOQKEgWubrwKT5+RCgEFp7J
E+bLIi3AfztW/XoA+ogTl5zFVeyko1mIUA7JOd/MbY5r0VPvXWyVLPLbOzYd6jsQ
uIQ40OOGfIqRFQlVoQBb031gQVvivb8SzSxP6EqUs2OxfWd6tCTFJk/lWAQk/Vu2
C6F/enap4s0htCQl0fivlxb6/0qsWPyYfLmMDUEkk+HOiia+n8kmq7jOCkFDsvZl
V0FVgrkom/g3fI7MPtAR6l5IqEb2nOYmj5EwcWzrPInK8b8WoaMl5mA24T/Ke+ux
5B4PbNQUXuWdhbp3M08fa/QFnZQtOHnj+OfTjOTymmTAm6bMpstHEwnczd+QhJ1B
dKrUMhKeVnJqzbB4caHjp41ILkunLQ2JxAfgRMymprhD3As/fzQ6hGSMJjkQXojd
/JglL1Xs8H7EoAEmatNqf4W6k9IidoM4lo5RbdlaYnmH5zrExVqY7VSl4j87OB95
HAwlyLbyQklMzBWJz81ZDj3rftJVf6Z5eutyY5VwuIWRorsGa1N7Mm2JqKkeVgYI
cMZPtFNc42gt6zt66Z0fsEExp7AVb7Obi48jM4KYuhgazDdZyQ7TjSQYE5s5YMWB
bRddg0yNehRXkrF2Boda+Akt8wWt4cuUvo1/V0FVYyHJt27ibvMGAsswbWuQPwBi
xHes37xXdNwSx4sZDWJcDACP+jLmnNN4oicMj91lyC2KrpeuFY1yJBUB3snKo/mn
o0bnY3co9CPVmybUUJOjhf3RLFkGJoEVz+7xxHUmr9LMgSPMJFUy56ba1/rxRzPv
qXWuwpZ6ARtuNUrnrTwjS1H87HTp0oSdOsuaM+aiIJwQ3kY1VKV6v7fjCTu3qbec
PzqterEpeoJTeeJiIq2gq96d+bPRv6VmNEIKb0iC2lmWtO0LmkEjF8bONG+tN4Et
KPyZywgQdqkQkWY4snuGsxrYevCM/uM9MnKMbW3yXW+poh+etjV9oRdy0s4fbFsa
s90fNydkFXa44lZpQ9x+629qZs2kuITgK+2l4TCjI3WcOmhcSv8aj0N1L8/tc9Ue
5m5iw45sn/GGWpZPXXdutj6elhPqDBr0ZU+f76sPti3ncc3qYYMMShBSmqJCDgq2
JVHF6EXrK4L+F0aIEox1ORUPzQ3H/I4ko5Ft9/ef9JVJ0q7Y/FMv0ktX+V6iybDF
b01obHYCabcGPvB1DE8DfauIDfOEi/zWk77CKpI6KUdkP9clBrpHGwQsRUNWiPQI
hZ0nVXVkM+u4CsiRC/Th4kerCRwRy+it7WQy8/YJ3T0hTYvnJfCds5lqCMKL6y6Y
5Zh4Xg81AtaS7yuLM67xxKfb+RB30LdpJGi6O5k61cvv5DnWImwLnqeZjc7y6l3r
E3wUNQr8wElPKLs3H2AMJESATe8aJwB3hFYQnCy5TNOwt4EGECyZv7agdNaAbJxU
zGtrkvl4cWeQhbtaxp1vd4SE5PxQTt+qgVcAUVFqFjRLGwnmit0uBdDLjQTWkfL4
AWJQQ99KCVEdvwFZTFejRKTX11EwSPq+bA46/vNbtj5Cl5tHgHaHrckmdp6SC3qn
m00OMU70vUv/mFVv6JIRrtfHRymQqW6xLVdBoDBfj1HUgKqMUBDCrws72jtQpaO6
bmLBbwI9R2fg8xEpOnT6EmlQMQVLd2wYgAna+I/oavNOvg7HDeUH8NpqJ/wifNGg
+BLNkpHNRq5Nw9bQxY9ugy+fJP0NwtUQ8HAzI9okw5TlfRu4WTHfDn1ZfjsCxQSJ
85kJaNuvPHwbh/3tB72CBiCw19MKVk8dNhL0p4X9YgFsj92xm9Yhia6uO8Z0qXgf
JXO7ejF2KgAhKRuJDf4zKkRdID3es/e6lgy25msQAeL21a/ezMm4HAxp+UK/SDJf
EUAgnjVPH/1UPyhKQfXoC1F6zXwNd/mZL+9EdJUn58nVbmdOB8i5pYeniBCm3GUL
oQG/WwuRU4SJVAjCXlvXgHcFysrTUQS33WugyIoZCl9hjVBFNcBL4gg4CYhujttd
5MfLute7ee6BaMTxzJlRqDpD3aaXdbEGXB4iNZJ4ydYl+QKL/ab5cfYhO4lwxWQX
Kc91lq1pGF1r1zweOdNJgXDJSQQGR0TVnKrx51aJdNlul6xsCr40Do3SqDKMmR+e
FkUyE0RGUxfx3NvIhtZ8A1TBJ6B9zUEj2tTQA09GM2zsOotemuELan8uqEiKpdDf
10pr2EItIU7NpkwqW++MdXgKf0shL3un7INaGl74PcuYmLbYrdYTkY4RewHSLorI
DJZ8hKonILs33aT0UlGUsil/K90lthFn5UyCNnTAPUQV6dgjQtkf38IUjylcmFpK
x1w9qMjhq5dW1E6NXySOEosAqJOAhzVNqDvjK+R5vAD/W4J8UGJEme/QNmbfLyXT
+OZcrdm6o9NJslPajly3wAuozwWeeq6BOatDsgmaSGTQuIcsEgGguIy/BNKQK47z
tC5N2Tw5YizNsf3g0IB1pBosgwiyRKQjbhzqm/tEf1pyVT3TjFisEveVrokAQlZQ
vHSOzSS5tTPoaZjrM0CMCp/r76y8fp918oXIMQqLfGv/NuRW2p1uZT7KoJ6TyYTv
y8EUmThlb+XqU3FCF0UJJAePRhuTa6cAQwi/PjhYHHNGTsHsOrEIXMKSqOKAobv+
YqVfzgmGe/V3jxLrjml0V3S3XcJVYLNP4nSxu9dvjHf1U4j4EIUAXWMUleyyhlmj
5XWl0ZvikMYtH/VhGaAcbVeYOgc4MyBbzcV+DLmvDI7z+Lp0l/Ar1UlU3pFz0ZBX
96Y/mxDb+uL7a4+ZoZyvqArd01lym4eaUpC4gkcQBSlVkxJ0xh+aDvrseof4y5EP
C/es3dl/wKOLyDn3dExAU0vUu0QkPEic/8PwKvVTGb3nT7MvAj/PNY+T2GjO9Itu
srk5h9bUfRKLxRpW4fV1CYV5wzrFdlTseVUONtH8o0rpvJ8z8Ir0Xq0d+DA0fc5F
IFLhhagabeEEhurO9jnlQrgyC2Syq8ZVxMneUcddAdYxzH6mS7oBtccUDIfffkPn
RqkeGtaUoQnipGIiOSE7Qqv+o9VB2mw1Bq3uby7EqLFU1h2onD12mMeq+yYZu/Bw
t/qI5ib1PCzHPLXqwAh5YtCV7d9ntp8eOhNs+qu1pNsPAkMmoWrIuo9S/yV8FpzO
D9Yb9o4TFdJZtOEJEogopQXLQ/EKhPkeDeufwn95/YMNEsHV0XDoTgCbNRT7KoGf
i75Lz0nvF802wUOXoURfxzlFkgwRt7gq6bezvPkVKZiqjXJvZ/98VNC5cCSqqf0i
PCUqaRKRmjnr6pM9umQq7Ee5f2ocA+hLJ5TKhc46IxLnasZjUlmsT63xfQTzGU3S
qJr3+B++HuanfuDO+hmc+eRtlxCCXFPflWGexuqb/2fnB9o+ZA0PYaKvDeMert/k
xElYGyfzE1jYae1pyZRRUXP/ym6wyvSLxL+yPo+Xpol2kjal/9vhqaocvI07+Ppo
PzBMRBk2KrYcOVPPKRv7AAEdFyNiyKxMWZGtX5RcF9G2noX453stiH+EHz0pQRVw
e6mLlcdvTNBpkGrZ1qhR/b05YdqulVZ9LjoZ0vo1VviHUPWSf93OXnHFBq+U+lJc
dlgUE9m2P2GexYnF+Voen/cItqHZnDbcn8VeiKOUaXyVyl08aE+8xABBbn3t0bmC
evQFLPWuK/ztulo6GUIXEsZuEeDJxD0Nles7QuwcF0KLP7kOBaCAeBnTGbBuQGVp
SFdn1aPwLdVX1J8u8JqWMzTGNg/IErevhdEE89K/NLn6inbceuJ0noDj26ZtI8sv
+CbQpR9hvAzy1+IThBQk07/KVEPWrkN7zDfbTlnqK4T0SlArK0Y71cuIr1MRiRgW
2cFtQ+WBInbrt+EZ5o/MoJ9+s/KNtVyMume2De39ZMMlmSAAb0G9217L3iE1Ll6M
DsjCmQQOCdtAiv6il0LIfncer0ldIXtTqyqVgrk+c5JVpo2joXbwT42SjOFoimE3
y5ikYPsJ1QJj3B+rDesuqymznMjU7zeqm7cZkH7mLVyekHrR0mWY0w9o71yAsWGu
U3gttZ2ZfMFUDvXJfSAFocXq548tOYxgrzbJ6hmi+f/KVynD3+On81epHdWKvsWG
6n08b8CW2FjgIKukCls19KAF4vuD/ubr0PgdBZm6B2l0UYjT7pIXWVYjrunGOeWY
WlOF7IGpmQFtg4tJ9lwt1qViNAuY9f7uU2RJfKTvi2qAJx0qsqre8CsdytOxYZ9R
pHMyxEhBWqabBoYhMOT4CmXOSUuPipFL/wHOJzCd/wTm1QuPiJGGxOr+qeBbRrPv
7nQC5RHze4lyECBKxmh/kiBok9aNbPCMI44ZsoKoy0qqMz5QidzAjy9lYGTA1nV4
iz6ofOPGmtTp58J47UqYynbJdKBuI4+nwzkvdGxTo4yge1DG4OPPejNhAJxCEuyM
h8I+lTB69JsyjrpnDv/ML8cNaZEND+qSlmkwAqWshxAno4rqLx3w+zG1jfAw47FM
zmFnMgWuksFWiVSaz6QoECNMVi34ikxbORczGhZ+O4bcR3kyp/HqjHOrUHNQN//U
MiYs6MVxADpac7G8tG4Pl+1C79xXiHN1biHXB3A2W3UcWxtfBQRC5RrFnlu9F951
0mvfFGbgdZJuEQh+c7oKxHhQScFgZUCsjz/Xu1OBjr4F/aNAJCmL4xObxZ/lNCUt
moW2jFUHS/BAKU7QZLwbQcempV+J2kwanFJiB3zMOdiFCpMegWD1kgj89SeD/nbq
TLF27CqVReEHEQ3hWqfdgMFBIBMqRHsss7MOPREfLXMypf4/jHm6wEMayWztBPZ9
sQHH52fMx8Bqrn0M01vSdE5ABSOLf7Hm0WrjsLfSD1mDjpW4I24d++Nj4J4iGxRy
v3QP6txYd+ovcLL9DnIfjSFk9mgWs4/OrJq3O5OE3UWZfksiBmvhQRk8f0IszL1u
C4r0NpFcoZRcnKjV92aqhCRuNCLMBpyviOJRJCfREGsG3N/XkGGPDe5jIiJx5Lb2
0sMOtKt6h8tjBeXK58wWUJbEhSGrdpV4EF8fq1wluOGlT6YPr5DlLiKtYh6o6Ido
j+qlvFFp47SXXTd/cPOJ7ieGvbVLX/JR2vZkAT8R6BlI2rUN8Z0UByRF1RVI218x
Fdhth83AHAwiRVNTOeSAAdl4QGdPd9S5aZj5jJgShuUjLldpNMjpuhzLBte0unwP
OkSfBka0NODQh8eO5z2FS2KIVjW48+j+ZfDEQYEIbajdm71HBtGI9FwSSXzshhTf
OAD6HWN92IDT2RGo8idXOHBCt9MjgzwRh4/fIcAjXRQ+gxh8Zn5QVPHOTlswsP/C
awL7d38uhsOQ7H8fQIcxAS6PPltul1PrbFBkQo3PIoVZ2py29nyseixq0DxXsZnw
IFZLCG/N4cNA4egx5IpLElIXWYnANh7Mezi1EJ1eFpRaOeNZAev7jQbUaMLbLMfl
F7UzObJSdq2OLjt/vHsuCwfNHKAazUfZ7kciD557+1PDx+N+zF3+qOZf/AJyJd29
MWXEJ6a9Cf1Cz/mlx5uLND/J0ElvbC+KI9IV3hA67cyCF1grUZH0Ab5nHgj99ceJ
Z62Y23Vcr8YpjlBkC3PIMGae6ovRRbSm2NHM6DZ7qipplzJZ1x72XZFmuUa7Z4wA
m8Ctv98wLjIRTOWoyZ/0GHJpqcL8vvSVQZlbqIRACHq1i9WltM/3u4cPkKPTv6fa
Qcz9xyJ02AuX5MWA5Z8/C2c3DaAuOH19dQubO+g068KWo3eXu5w7yPFQYwzI10sv
22heTZTLN4490lzEozw6bVrzNUJjXdhvRXD0ExIM/oEXqPS5AU9d7AOLcn8AMByI
Px+PrjoQQeZbqgF70lrbiLXkogTL32Jy2PWNvP2SoOZrqegIudaJRG0mjPOlDflq
et6smFY7H3DXExn4WreLbZgwvavjk9z+ewuhCw3TDWpB/iWqMQaIJMrOd4jRr4RO
/x+GwVPEWsT48/DOpwCVcFkqL8DlQEwMLgRgLBRPxPK1cIHMZRHLWN+XAYNsQnSD
czdDu2BvjBLkHbrxqnPk8QMwNgsz3LoOGuXH/KcTBIzLeEXyuZmJXncVPMLKw2Xv
3g9FWXcAZnyLgpyQlX9FNSmlZsuVERYennUrCN5cpk3O024M/NYqgeJRHQU4V92J
B4ykvjnNgSy2aLmFQu/Pww6vDT7ilr46+pF30FaYiBne5DDq1sUJCrvBKzKZH0q/
R7uQNzE9p0ITjRSPwionRGEt0UiMC7eX+n2+JrQa9TEFPr2fEHreeKlW13e6UNHw
oMv6aShL6PC7rIgRcE/iO0aPrbK+f0df+O38j+ydlY2uQ3hZitfzcBAZCbdsRhwF
6V5EZt/67aOiAyBjj9Qb+d634YLMmUzhGBtyy1fXosxYPZ2JSiEWfTplGTzzTNhX
K5a8ddlIbQ4YsUkZ1+Ut5Gy5UuEHsjhvjS+KaDW8UdgxnCeI7JrKtxlO0/9zJi28
rYwVN3VOBv2/8qKruHfF5qLdnHSLge4FUcwB2atcgJUX++W1wgUXsCBozOTmXuDJ
7Y0vi4TJjqMU4pMm+OiIrv0vqmtc8jxVt3KCiAVoEa5IsQaIYvpVQ8VSzGhCO8Dh
ibz4xliEfZNGj0pcM+1G6xiFxFpo1rFlCEQ0baybZwJUhDP8pja2+pzmzU2F2sc+
oBlLJAY2oxT1lcPgk4vcZj/lOlL2tdT2xACW2U+5GDoJvoM3yS4Gvp2/uRQ5QlXC
bOxX3YFzwbk57mFOH0O2C//5CYqALOW1gXWqyTc0ck8VcNnD/rcZBHkEpNm7nHI1
ya7BMx3ocnt1iBTmAdNVpFHfrYX3JQD+41RYc2PYesk/H5g+owteZEv0LQtRB5mv
RE40TsTImPGht5u3HMJ6qKJ2m8sIyMy2/gtqOoRLXLlC/hcc+V36nHrkEKJ73W09
665iZFbnQFDIvwXhP0gfxM/FqL5CazWea7QQLi0pzl+nyh+f8jZcJ8p3+sinH6yo
kD01iL1OwQOCe9t9ScuPheS1c5HSZLLoi6muQU/AzQIZJuh3ecot5chvQUW37WY2
+BZPvtWfsEYh7EjrCOhamKfFp9F88zrNFzzUkGuXORbOPxadghXWITU0hl6UIZuC
3OgHI6x5uqhpJeitO+bJF45cGC17FdL9KvXH/WLRl9OtnsrzLXx04wjI9Y26CkLH
kBznyUm76WetEmJxg8EgP31I5m/A2T/7PuKCyHGM0XmO5pMRhY0lJUC59pxBjT6/
w4UVxGpbtqIBabnmAPRmJ8GR5he9cO1sJKeUpj953s3L0e5MHbOiJ+o8nYOLKMxq
Qpjq0PI7seCEzEibsuPRg9iB1KY+bwvd4dlN//f0Jd8zuOCorwvF+SCKXLCetpuK
C0AZWh6AFrwmoYobvbhTxGb4vJqxx14hv81Go0/JWXYhMsDI6WoCsSDd2j3JL2c9
Rr4/lmN2jABqBrcN0QYcNjXoUVrFK85qdfUvGycBwlu6H1Tg8xDsa2zy/+t53Fq9
ekrVtielETlKuP6QttFaDwh0015J/sViT2slBcSxV6bT0tgFje79Q6YcfU9Qc14C
77+msUnvq0LQnXukyJAfLyDEbjQWkOJVjpV8b67hNT1CNMncdSolWcF3SUlApibv
UUQCOSQT+mfCEQtoCQzFb2yOzcG6WPNDo9kmvPDH087gbrz97+jpMk6ImT0Z+gVi
/6rq9Ku2MToR7q/JD4BmAK0AZJjSC1jddm7uBtC7iJgvpC9gpE4NA9tstbdRcUQB
isbLUWuT95Cn7x8Kf1LQ4sHQ4Hc2XzK8j1a1EchjcBI2MCbyABBnGbQ60stHYurs
5k6g9iV3iLU2BBQZ/MU4ac+EsO6/nH0+iWjL/GWkt9UpLRSG6h9TVqFzqwjMZqwl
KdHYCi/yGlbPRFa9nmyViL+i5iV/LDx51C+8cWxQ7u3GqFEnWpwLmieT8NrqXgjW
V5VfgyFlVJnGUBDnsukYGE8SVV8X1k2Ukrw597n50OPA0iKosykbzLsthmGqg9hs
uHUnOx9w+vRsohPy1K/+N7Dcd9B7nAfe7RcPDXGgdhyBwdPMhgM2BarwgJilQg80
if0r2MDQixCw2KnwSxl2OX6G78IohwIESFStka7SVZrcY6udNs68pHGS3jCPMEkg
p+7ex+U0qwX1ejPcNTdzeyxDMicSmNZS+TZBYM4lnBvUwJ8vf4db3fdjjVAWZnEN
kIWedPYXNphE9xfM7nNcGem3KfR58vgcK5Ng3mmu8nEt6tR6fwFVPSjNQvgahaba
W+BKV2BPcxYtkd/x/swM62rYUuDJvrm1fl7XTK/YMb0nZzOK74aMbH/syP/NAZ3p
MUFfKLUf+tXKfQ1xJWd46wGv70bffDX3L+FyThh+S+DeUWfZ8sYi9YHiMQVfkGHP
F/8gIm9QndYj0Gj5eYvY3MunBDEfjdcwCzMqA6jw0ZHFMXaRJ7jEHr6hkSMWRsNn
rDvdPwPuZTf06VVKMIMzIjZvS1oYVDNW+AlvlzZorFpZ74HAd7FEsHTcTCehAuIa
luzjID0IX5WYnNfkyayhOTf0Q4zgKK1gYBNG4CmjA8EjMvrfa34uELfLP6dT7ACG
33ZAgIDDAvdSw0qH7EHQhkhXVlloKJjsNdZr9T9x5HSDWD0sDRprOlUUPCJ7KYOq
aKkU+Ao7D8BFuUrCzNyEWp/KMfbSCVTzmD0/S+Qyt9cudK/VMNw1WPaxOPHn/2Hf
SQJDjcSXGqRV1NGT0iqor8Zfskvsb+pxKMJlUSjnYCOD6h3Q6ZdsEFiGCt81Sd8d
O2ZbzTa3RPA84CjeNMpSBildwR39E1lnZslSjSKBepCD9o0D0EgHUlhegtJKhc3h
Q6TJDcczNf73GMNljPYjWI/vlbaFsJKEhiX6jr6kOgY6AY//MOuMCmhcOow5JsC0
855EvHZAXf1nA4Lz9K+miPL0AugKcp1xXESFKReBGFHDRy9oJVW0o2CxvMEP0omH
nFwvXBsvAt8iluvucxM1l2F72KTNahqgoGg2v8EReLI5DC2vz9xCDUMd3GTdnh5Z
736ArECQSiM7ZPXWJrL+54VOWbcuknd5bE8Ok2MGyw6z79qF0hXkgQo+fSKZBwFf
w3BXWaBeVBTCLSs9B4MXnelJQPNLtIESpq9ZlB/mitf/mmO7ARsqseFIS5CvCpCb
zMhqjrLBITuS119PW+Ra03i+YHUtS0wqpBzR8R0pZeU0vwCzqmN6huwCyOM65OR0
of8nTTVvIO3BgVyYLrf5bPUe9lOgG/hmfxAq6mQeFlC706RelfNgIgzjZSlJIdTa
ZTiyIrthK6alz9cjqJJ0NhWsJsBZ+Cg/iUTa8nGZAgThNgtcqONG0r3ptXx+wBBO
p5BXsT7wL8biiC60vjsQzS3ut9UPNK9lW0WD0PmRdlS0ZBwnsKKb6Wh/2n9M4xKH
Zu7tyYmZpyvJcwmOFkmmbrgGIFL6ipK3brQzxaIJfO0Zanc4fY1M4j/0/dVILs0k
3MmCrRHQmYtFXEWtOYRsuPu/hVd08/Wu+u4RC+nMiL580dNJ8yAV0Ik6VCLC0dMm
pAkX+duvJEgMNuq46h9RRmFRRhPctndEsHRA09VsQzY9RnByo/ubaBVRmtZYpNik
0QUGu28j9HSPEFbqEf+6G73wby+dqRw5TJhEajYOp5h71vMIGLf3uTID8Vyy1Por
+w/paD0F5e4KyvqXs11q2/fNrvoq2OgolkzS+/nlSv21tKeSvWt1AjVphmptSkyy
k+bQstqX6q8C7Jr832UwBrw+eT/3h0fpk0uRhRfsgSEr+yBZpBi25BCfWhHpcXSQ
gPbpxLDTf9Ym3FzDvlvfH25DnsO+OtmUlFbnd9YFQAqwOS0xd7BJcl6QtnLf2CoY
L9lmvB1bvzo7akl+hqfUBdaJjPnqT+HxovmOh7dKl0wqCGErtr4O7mYKSTuNZQdx
qF0M5UnjhLq5JMPZHuy2rKy9qkEn3XAzyz/YiUHZq3RN+DqgmJwXzPwQnV2qqp6W
yXllBNsVjTAn4NGqTj3ScAqIcKofQodM+uhaaNHYXLrI54ZTLnFY8EfP9vxPIEf1
cl9P/Tyb4QQemSBmGysIwj8ZOaHDBgv29Lak60gfIeWMtJ3tldLXqRphcQXsRlEA
kD1QGM+d1wbt8RjH9G3ueYwWXCvJBhj1MX44UVafn36WlwAYEk+YoicbGHqW5kWc
Rq+hN221HScAvVnxoIbWTEbUBypuctX2Cz4q78wijmUpNVAGvK06gLR1XfFHBiMT
X33HzHb47zxn5Y4pGQI+/ClPGREJfFYWlIvY964LcmW+zIJP4j4OC5HO1/Xkshv1
JO/SFIYD5vsR83dEbZUG31qn9RWLvlRmVT0yuJOtppMhW4zapA7Dn84QZjvsAPWN
l6GBfyjN6mEUJp6g5ZXtjbp9BvJDpJh4NGST342xcmbB1s9AJ1x7Y6aeAPTPXvwk
Y4yUsJLQckoLZvxSVySWUi4Clk+o4qpZkqZdFyJaRSUqxafXl7bg8pCicPxVYFa6
UMlCEzW7frdrSDRO/PTnPNegVQDVGBHNILW2DwVJC+hmFKrXatcB82MX1cS0ho8k
9jpdamNKc7/gbsiSQ0DZkN6r+hV3FLSgrAIMHHfzh7qZ8Lk3rAXLiXgTPMyQyYDF
2/Hd4o5oBP4uEv2ZFIlyOpOLyvZ8SEDEWNvWuwXqc/Le67bVCcwUzkZdYlZDTNy7
Zfs8TwRNE6l2Ap+RrXjW87cVXO47zrvBIzZ+SOu2gXnP2VjX/8gSuNlFuYFJ5Ogi
XU0BTpsKveWCPZr4+W9fsZs5QHNC3Hk5WK/EiACNffHWHpfzFVjOZfuuh50nS49S
zgNGRWaar5dK7roHrptV2Onxp2b66lr12UILkk0wqh9TWU0GGauYYDuSRHt1t+6V
LG1/BJCWVPbSNQgB5G7UuaG+AO8Ip1AHG3GUrEYymTgnkhoayP7lUmJejulgmqHW
Yni1i/uMF+kIdnMZhUoHguE0alQa0iHM/9w7wzUFYoVxFZBNpZAodZggSHjPx+VD
qvPCanuGa1r5xR6/5KuN5ODsjkrR2+m9eYmqZULkqxEX+wdJESoJBR9vNBMCVUwX
7TGs0ah+SmlMH1o3DTItavokpBX07MDELYO8srhy1Z/6JEtmJSNgcx8X8xCm1I6Q
JRK7rKJovlqrfAVqXGoDSbEAvhCuLTIK7ji4S/SJc8s9cKnMYuXh3wncro+ZyLkQ
Tiux8zXAKrsugEK6lP15KQc8G6Cv56EcTT5eWnOtL1HTR8IMCjCZjrG34DZ0xzHq
GgX3Y1UpfGqU5/rTXxQQzEoXzbayIUhlxd8Mo67jjzNM7FotvVXffdoXSskpsHgA
dgFUH41nITMfY+d7278cIuUaaS9Y1NurjRq9dRdTV08nqK8wcS6bnWKWDcBNB0iX
zxz1jhtYfBLcKMPvZDNuhgzETYsom7/nSI9BlANA0kFkIrL5S8SCaeYZ74AHoYW5
2jgbTIdKOk4V+SLkTx1uwYUaYvKUOSYaQLfqZRp3Fly8GLwKesVtDepOnsjnTOYN
WyAJPcT4HuzPdQDC1pkijd/4kGBdrk2Xa0iH2UH4pzDakqTsXzS0yD1ov+DWC9zk
OIm1gqNXoBV7K9u5DxeKLP0AMM0LvTc0gqlgNB5WTgT8BKaQbL9DD3nfD3fx2qqR
f4BlkHXNHTfF4SJoYhlJN4fvPDw8r18NhpRXZbUerC3rI8aCOM0b5y++UaThdmTW
kXnDUDNQCei56svZO4VWCz1LqWg+F7sxR5LYbMJ5gQ88MSKFZfiGjQ1h0B/R4HLI
OpYu4ZqkItlcO2DBog6BUeXElAND/ztE9/B3wpmXtZNrktKtz7IzL2rpXhQkgDM8
iazGhS15vdEJ5WNusLX3ZBRSCHkyiqy62wU2g3DhAp7AuiwwElL1Fblkfc4hXnW2
0QFXvwZNNs9A6l15al2CNY5urb1KUxcaTOlW0S+OPkrhk/Y/4QjQ4mgL2gOOheVO
G/GkqZa02Ws3KBPyiEQTwhYRZgvoeLcoTkV4osW7+DLDX44HpbeNuQ3juGoWk4sX
lEZPYdDuYm/SKN5GRvwO8WlSfWxx91UnU1wBjoqGtu90cwkzD1SbfFsKwUfyWmsa
uIKekDXG2lN36M3FY2YFek2JTzRx8Z6O+1ycmCmjx0kcN08h0clu62Vwrx7uRZG0
YecNMrDPYdGz48CYPIfukQel1cdFiNgVgnwnP12bathVBVpFls0N3+T+Gfm8SF0C
W73KnEtopHVWR9L75AhZSuGPm1bhjRCHJATz6AvsBWnNEbkIWd4B5gA1CStBroNP
Y7MfXAGQyakyQxAK3Pm47wlBO0NqfHsz4lgiSZ4XzaNNfamq3ylhXNXP4Wh4RVNx
ggO98jEtnXLQs8kg6qYGk5J7hbVW1Q1jxmbbzGELi5PjaBAkKaggjGxfiTPRRhZO
33g09XszNvFJSIPGlD3Nrx003ho6PGp9S6NsHxtJKmYCGMcsizmiNBLV2lea7cKS
Q+nbplMp39IblxVjevANYxw0BQTt2pYhpqKiQQWb1ls6mIkwPSVtcj2YxCoAj/Fe
76VnqHVb0So/T6Vxh37IMSsxZbT807PzrcPF8p9l+SvFxPoCWeI7TjIX4Y5NswCs
AmoiDwqQrScMnVbkw+N30lUhhqoGhA5mKqQKBH3z9woABaEWOH/Px3bZYbZhFJn5
j7irKJIyUcA9TQIaPajFOZrgIVze4SZlc6MgjIU3U8QJBUTS3F7Nq7xO5aim8t6m
WtkJFvwi9xvHThDgF37q2tBiaGZ0zPm6L6nhBuKcT8B/q1oMlbrHo3fmRsMDVZS+
Ml1jSZuQjB/H1FXBO/wsbLxFv0NNCFKhAX7lOA2XBstEY2ugTsOpKlYHz+lu53pY
mSlIqxZt5jtI355e5kSmF9hXCuVxx3emPVDPUh7k2V8zY5L3fv6kRdpq10fUtCaQ
N0r10oiZHn8PMdTnB4dcnWlH6E9fvHpJ716s9poHgBOfg+27AS6OAxXegW3ImFGH
DiC6upltUdpDI+jigFB6bJDwrlPrKX4g4AfsbuqNmLXRtlM9Kck4WQR/JmjwNgT1
OlLIHWfhPkpl4UzR8J/jaI54vBT1zSHS1UKS6d47WbKxk4lQ2KigIcLkiuD8OF8z
2QeNScwPEARhrrd6ViuSDIHlddxlYcFTNoL7Rdto4i84k5t3kAky1EJxGpG09mxX
aBdRee7uO9PmalGBYypsBptlzZjXNjHDzATZiU7zVasjVvrDZH8cjkwC/OBhH+pg
m5JrP9hBXJKu/Xt7HkweLpyPFDWcvuEAMlrvQTYzoEiLAychjGUaRxKwfUxsYUTf
ZXo5gOt4+ZeQWDz0pTjBr+iYLt8vfoXcRByotntvMN44C4/zTGybswMARuHobSH4
1D+z+3M6Hw8s/0+BLafsYQ0KVCR8FhcJ/NM1UPpzEffIu1MZZ4k5wf438nHVvIup
CWGVieeCMmT8u8EM5oKAvOO/e7cgJt+FAXVS3j8pmE0nvGi+USoh5mwbpLnxbAsf
BTZ3nKJphZR+F3UeATB7KZTdNam7zotPSMps5/6+eTSDFm2iyP0HiCPx/1jq8l+x
F7fI+HTJEzmYfkyrqKG5Cv9B/L0fBB7285j7BYVXWR26FragG37EKjX0BhckSNjE
Lk6SwMHi5mp7AkHqHd9e0VU1hQT85z3xgy9rvU4HFMb4kflq6tUDMRAT02fW18ic
bbwG+VU2slftY8NulxO7YKpBDhC5WGYJq9bwnmnQHbrfZGLEN//PujPfGar4qtzG
BLYWoQeXsTTgnhslcWp/oJhZVeuzR8I2AvcJoGMfNo5KQxYeBrQamNzFRv6Ijo2v
SMYmZr8Aha4gc8hk0Ux5dGCW8h1tdfc0SsnuWJQ+kcfrgF6KGMk9edgwLdyArIAB
Sw5i/olWPk2lBu2hMucO27zTT7bRJPVdIWF1YDxm9z/WFjgLnwaxfj7LHSpo32pL
8HOganNp7zbqhiZPSIwfrSEXv/gp7gMTvLkbAxLdacqciogvJR3TgPTLLeZTdrNt
Vi5c9/JE+4tiazueDpYozPVAblkOArMyFkoJqzRr0onvtkWdvmQ33nTWnM2xfBce
viGCxQn47hhTY/zj7Nys10IZEJGRLL0iptDcOOx/Ryk1bqKjgPTGGHe+0U8dkzxk
cB+xrH5GlgeM8Q3NFESj6bOsZ2gQzLfItsfNbpt0CF1i8+YV6LLfYjJBWMZCJO3B
UJnF+mVYg/5rFyvSSGvrhxMGR6V9zuHiyu8yRZjl9ib33sRut5PpEejwEM9iY3GC
m61UTBVQpWmpD+cL5IKO3DKmavFm1eYWRzVxcTJIls5TfMXHYrNAa7doo1eCGZ0w
oQIFtRjhYKmmdVogXt/yuswu/ybExXCqPP19bK7j5Sw3/zJ14VlAIjs5HItrUF2i
/9gSfo0+cg/YHlyIhpeK2vWREsZVECMgiaiJOVQGaRzpnMso5J79aQMWc0artXnd
mg+bNWxNn1wRnx5djJnrVxfvZ5qqniQv7nrLkBGaH42Ugm05F0ucAEkZM+Imskkk
Shc9xv25QbBbe6PKJT/7smjDgRepLJJfXXLIVb81uUK1CvqKTgfPeOnz/0pENyOE
LQNzsTq8ZEmSuydcDv1NiVcUaUNloYxKptjoRvTl7Hc5+LBQuG46kkhsG+k71Hxo
P3MoWLxX5gg/3jmVtQ9WWtn+mKOI6KtjA8ybCmbf3cc/2s8TAcuE6rcxD6F4qYHS
nd2klIXDTD3Whqt8jbpYV9UhzOkdjmE3Dkuoo+oMCbFIFSuJTHjSt64XOzU7/eje
vZs7aUSstjf1+thsZSmtVUqXY3hlMqNll8DhT3kjZrO7wBcIqP+3cjn9D8ujZ8kr
bmrGrXNTr5Qo33oqPK2EScBrOhXqigAMSdub87ELzQKcnN2iQJgUFrUYlcXHm/c9
7RYXcw4PES9SUTXPR5s5yBqSct+WPj8TaMEwxnt+5U2/rxfkJDvEkj64CbBJLx5u
c2hCOM9eWcOkHusI5+TZjzhejil0bBtoY2b9tAO19wT6EOq6kcKXx0b5w1pkNhtY
Gyppt0yy3r2SI8DL/AR1mMdFTz0s19Bpl5ESz8nX5I7A3cpWvm7TEoXJITIzI71m
9lsOezpU+kZq65ImliCIu6OvIHEhdLsaI9iNm4DciClOq/vRi0o99nuo/lSuDqhW
nEJMGXydc/MIg8Ir/16hUHVTaNqpz0qOv2OTsmilGTkdIS42trUqxwrGGwOVnW2J
VaRw49DAp7LS0P3RSG/rQ9plqNYGpsYAJNkKQdLz4099cjbbIsnJ/KNsdcGcOarZ
nuhKkeOXWgixYXOIUsH/9w4+oV/a5ZdnYtj7EEOJ+0iraEEnoSMw43V8uH3Koezn
KukgMJYI/S0W2LXViJdIhL0pdoXHbIoBxdshKS6sSqBfEZIOcFs3hbwCoLgamXqo
SqxedlS1X1OW++VyzTLasJkjoKGEK4afyAua7teO9DmcXzRQ5RXVQ/7c2Iey7YvS
4s+AE7P3X4+mlM32Zaad1oapwFory3cICYBpZzFDNWLoIJJ6K82WKwvuLV5ajVXa
QZTvVKFOuoDUVd5OmUFQAtSnTEjmxUgd4R0Gp0h90XJ3ha5nv6D97+ir0tSA/5zz
QUMdf4VCZn+HrdTVg3uaa75nHFAZiZpj9+7LXWRhCoNVKFIiiRZELMiaiFarX89/
lSRhChv2egn7gX8jRUwVR+PGmYX4BdYS4Nudtbvy6uWpb8mRdCLVeEHI0ae/BK3+
et9XsksGAhMKJYkJkSxqe7JLhzSdbtk7QM90kEk1gpQzPqF6QvtVJUUylyASa/08
wYS/Xx3Tm8i6OB7x3tKN7e/7meGl4L52HHmZorZXryDmpZ6f75JsDP70YELG/LU5
DVCHni+OLktqedbVVNCtF2DnDEFKpYNVXWpq8TO2bz/TT4ii7Yy0q9q9Tw3m086s
KKthHbngtctwZAamCEyUhUrxNGMxi5QVGLqKgFyyBsnmQwghPe+pfvdGL1WPr4zc
gBJU8tzgaTJto3q0Q6wyV0fUj9FEGwgyFyQLpyrpre6WFuLKIo8h1MYb4kbJXp7s
sDGM/5u1AS9LvSMqS0H7MDHRqsbtsvwNU8CVrLt7IdlD/DfAm0m9i7wOfAxfHtnm
ooaEC6vJ84kEmYruEHeeLqULjSYKNPaf7e7SHEO4W05/gp3+YEXZCZvUu7B6m/HJ
0Uc05J0qDhdIH8pKTraAOrtVs++yGVH0ndL39cflOQs+hEhwOnm/mrX9x9FScVbL
23WI8GOKMihtKAwrt2mtUZXYDY4UFGDhwdLp5kV/ZyGLBQThg4d2McuqZa/LKAdr
9y/2ay6T4Gwk8JI+EP9JqR8ve2AUxeYq/URqqXpl0fuyBLo4KZ5p6zOM/8MoeMLe
JzjwTIkC9nXnZfJOyC2GxtrTop6nNRNVfp9u17w4sAMxWfRQWEYOXiMd5nsUwX9X
DlPIuqp2i9L3UI9MjiyIxl/TtZ0cElyKsI0urJEU/7OLYdc7bHG3GKPp1BdySWoL
ZHEK6/pqXPRaptmWl7zhRfJ0Abthibe+sWlLA3oOTB/b/5XlnDIQP7rIMvsk0VGj
GXSnYHmV8jMzEwc30zeGJsqfhKT3EZ+qZE0Rwa/578WcnxHesc0CqGgybv/3PXCn
8cRe2lAbd4ZZSkAT21oZWwVQk0Zw4JhtgSOjpMB135F5TNjoIDylJM4Xd/TpAzd5
uXTD5w7FHq0no1JN4N+i8YxZy8HQ1myL/x7Qcqp1cSbBUimzhyX3qrX3aCuWgAFU
jXZtfJlqrDAyehrGf3zQgYAmiloZ8sb8bgNq/0Toz5ztBbMciRiKvfZUznlY7yiq
et2s43v+ZYjOI1hI5XO2Ws6mbMfXrpLSHBJbO8uXPonPv2xSH9W4gYcSImELggEn
s1BmnZAX6wiweRM0EAZUQRQenDjFDFZ378e4VzH+gAKYX4DJcaUmY8bcTB4Rc7rc
+tIxv8Mz3nl2RfuwtR68Z79YW8qK8fESvOBJOwbS+oPG3aKRhcZ0Jk2TZVeWwIMl
MI6TpwQFsQABiWO3VeSaNYw8ogq6eqjH+OFZBR1+BwdprzOGOLnSJAcFM/3sKqoz
vBOdVbPVjLaHtgPep39wzATqe0ke87L8Me9uMoo7oOgTdYljCK3MdDTd7XiH8hxp
Oq2FDzuUuqP0Bg7plrD5FWxWhN6bk+ANfInQA9uurqHDQqaLHE68Q0mD0p8Y7FCN
m0SISkgZro0D3kU8ISr+eSRpFbwscXChrU27S+PtNTKJyNPVF+MPgIWOZxeokCOp
cQ4Q+Zu5cBnIXHRsz2PUqy7mdoAxLLCgJMx0eJ/THWAYHBSP+Krl6AjHXqT4VnzY
igfQuEon/joGacVAYXDigFNoltNyjfKpBV47M/S8xnzsNXUmZcgpZe81Oaq2bwMp
7jcspmMO1Y/zaTuSwon91Oz2jsVMMWX/vORsAD+fSo0ZkIpVzMAJu31RfbkwFQmS
Cn9cs0DgXXlqM+yRn7KLnhyWS3DdfWV09dQ5JcpwkPRnaL9oFrAqB7D0CJdEi75a
cJA9IipxeQNDIdWitnMCtBvFAZfhKQRVg6EdjFuF2QD9EqqQSJtbE3NIHsvfhM46
VH2xwrnrYH/mescmu+FFY4yaHdtgc4FCRo+upd7gCmzGILbX6xEVszFFkcxMdpAK
OTbKCN4pdXipR6fh6Z0Y9pChV2n0ggb4WK41tvCuXcEx6AZ1d6YrU3iNO8v2O6Vd
eqSAWdl+7jwQWhf/KLuwijVDjGOn37FzjKPSKCP46wHK9ZvTXMXnU2YnLMNdi9GB
YPDYRHDoUoptNgwKkLzJtCZkaxGX3xqiPTKl14FXRYg6+knj9ErnkHEhFfMMaiUT
iweleeCyX1MfqNTSiia5z3jBwlDss9J/BRoYJwPO1U83FGAMpfJmu9kdl8xZiTmU
rK/6nnFQ1nyVUuxwcR1WOAM3epf4yXRwlGMIjNWMsbT/Orx0B4pPYuDB0JF0+5ml
c2xTouqatxUSY2JKAkop0Ag9RglONEOCkZ2JQViOsPJEiKwPx0pjuW9foP78lSqy
7kNQ6yzQCeW6k6nl+g5kpcdElg0AWLe03Wl+gEk7lp0hIUf+ksUF2lqAY0Xj9bmK
72ptusDO5y9tbvGT0SifuB/qotoPBNHLdgmal6on9lgbqFFdR1oW3W2PM1u07t/9
bZ6t0hGA4o24Pba4zl2t0oGInzZL2b0NSfDojn9tbGyx5rs4vBy0g2Yt/KgPxv1k
f3ndcBlbYSbNRyshgNXlqegLwYU/HmaGw3/xTyWi5xqTTMgEI3L39kpqu2uUGcxy
TOAbg+RKyh6Utrq9phx+duzK3b0pbGZUh5+Tl5RkMJMPjmYJBDaDJbXs7XOERAYK
5XF+LReRMu0HNpaGQk9eN17uS8t+945hNNoOdVN1fN8iKqSHG9Jk8UXEloQ7Ck6r
v3GS9/3TkXw9JRJWJvv6u8XV7gqZLuHaCQqpKaENkB8btzuKhC51O+o/zzYe5hI0
HouhiK8+8Iaq3RpkBvK/lvs/SRfwb1IMrIKd7M205pExjE+H27xkVc2tQt8PK5EN
KtZth9oIcNpBaOtJ6b7jNEd+YlTMqqlbUVNOPk6rptx4CrThCMhXjgFfkc5uNP2/
c2SGhsrft4cKvrE/GsyR+OobpC8C9pt0vJHrUSW7/sa9Q7b3URUXS/wFQsi2Jh7q
smAB75KB1cLqbDQk+Rmb2ROT2owowXjIw+kNRiD+UvJ535rN6AIv8jZdDYGqZZVm
Wr1+R7xbdOhQnD78jwOoRr32MqBi/ZIQrQJHytctXMk7bFnAxg17nsmuRrZnVops
L1FnM+CItQdZisH4MEJojpEaHu5sJH1bjyji/RCbgh8PciOTp+k4WcjczrHXiaL0
MrT9saFWrppdNYCjs8q3kQRiJhF5Ws15BRw30bHBWU+5dl0ds37aCkF53ZvKtBVq
7808s76ipI677xNyBtlYAKxqPzQzEveQOB5feTtZXFz8lba1zps/+HDD2XbneRsI
xMYhz2gPpXznNmajjT+uZMc3T7w2BAvhlw06xQuR1SffSKl7IVS+iep1fEQ8kkJ3
FPF6WUy06v0/SNAFpq4QYOVdMzGiRtQrE2XLfrjgXsHMtiZq6DCebjRq6vReadXD
L1kBzFK1lnv52LvCh9dcRNeuZcUCloadXXFwB9F7E2EY9ZMFTiS8oMtbeM8h3qwN
S72p3cnq79eS9j+ZdYDp7/XsWzy5isjPptOnej/04VT+CxVtkRy0PufWbcFmlOep
Tbn5TsWV6ftsxDY1aX7abTmNO+LLEKiFaaTYBsPhvxb57K/k2tEQsjl4sKlOUVv7
WLMXB77Hrn4a1ZnVcwRf4Z9gMPBzRlLLUHQ/XUfqqYjEWft9dGZBtDSj/ykkLybS
7TCyRnu78+z7v8prmPr6VuAgfZoodzM8i9OsNVMexSMbBNbRPl5LslE8j0wg60PX
vx2h8bwZUhXsi25Jv4gPvN901sd+GMcdFCvaZXaOPC/yoSLBn/HtmnXH0PoQ4hG7
HM0GT6A/b0sMtFG0ZB3BwCYYfwQD6rtNv6QMtkt9K4lrYbyO+iQYGPFdpWbh2UvZ
loDdMNShqTI5ZCLa34gkQn2LZzwDgvrGnPg2cXrrk8ZmbFFf69VSOe6nYafGDxK9
JZDwNNcXInlOW9A/g4PeTv6l+JgAjEhL/ldXPJi0oeqAd0Th/2gq/LKzVWwozNW2
rNSbthspvR7OZCfJIEzR838hMjH45V6JWpZkfIdvMa1fPtWbUPbbSJs0v/nszlyv
OwoN0pTrshGjxdPxWy7eGF7diSBqfhdPgUSGBybmqptN9WJW/Mz33+yVyEgOX5dJ
eGDbR97JkFhdVadQZQ3mSa++NrN0ZLHDKhw3HREIF34r9jwohH7S6bcS4t74CPv4
xJNScL2Qnb3pgYJ54z7KbpOs4NggGEmwE2A9Uo3X2i5VMG8VNuWuKFFRwabvkX2O
zLDHi1n5SbRbLYCFLJZZZP5SetSMq3k+EZ7E4+9NPWqyhcsDGwTceZG2uv4poZ9y
LX735tgNzXuDjRQ+aSjAcVf9ZaVXd2a3G2kaW5u1amCpDtzCBvA+iLWMA7xFRXC7
uD4gBWG5x5kBC3R2i92Loa4JPOPyJGefIHV+YMMP1oPTVEoO2Mamn5s9BZg5l6bv
boEBTPnSfLcHNHVmf0HcBP5sCqGZ/zqJbzNW3I36P4Xr8zqJBlV0Q9Tbemzp6o2m
RZldQk8N3KO27KIsYGgrXRafETESzyPplxtE6+uGph+HZEfUYW5mEX8sm2NOxCZS
eztK6RNUd4ihYI8x0UwB8hF0rKMRv2YKuxTi7RYbfrrI/uBTqR7iy5kDc0YLCpDH
2yi0pmrsEbmAGgu+QIXVao4xYE+fvkV5foUh2XXwPansLSNoDT7aGON/qjWuhHTR
DAgUpIIc1e9YNwvV6UexWFWwt0yP7cYbRGTSPoPrv5YHzvnDY3mxB55VIVqOhLnQ
pU4IGJDCtW7rXO5KV5iORPhCiwpNm08GBXU0EI8Q8+Db298GzdPpopdtP1htivDO
R8CWEOYakskaiNim/P8hBV+lhwA26RHhEAUXyM22nYyLRodKMWKuGMi7VoHRIDVv
NvJGQL76AsgX8lfV1ATkNrfH7KkGFQ/Jy61XKY2cdITXlerAadJJQwfVPUgKlOoN
m8llWw75HhtxpSYSXNRZCUFU//wd0h3jzTfWzydI0oKDDmrP1gm8+L7NXvJcsmp0
70DJd3kr3HOglb8GfrcMa4UCzrFdob0Xn3vLfXEFw+5+1zk9bddW9Y/h1ugbhZ2L
l2rMOYIfPLaZ8cwXB9WcbjQ2MSZXJ4tYhGxVRAlojCXtwbcFOejAEl39eee8z/pT
qeUsir/yidOZivvGhZfxoqcKbK7LG9IpMqv9BMwZqCnfMoQEGXKXaAxXEPxfPozw
Rj7mehLDPPLGD1SmZRsJAAmrAQGsP1IE9kY+6lSJs8wv1DQ/PN3qFhlRFRfAJdMh
kmrGI+HDP0jsh/zlrY3MjftlQZndstPRJQNRT0hcHTb4AVnmbjxAgrdynD7PWNlZ
GqQzBCOXzPxYswX6T+HF6IGH7GkaAlUKQnrQoEH/IaGUz0lbZawJF22rz7b/8nbv
TmdDN1HfuLrHKEf8K69JmatRvHAsImpPo0UpVImgl90fIdwKQhxT6PzOdF3UXniJ
7NuCq12Rkt34IRNnzyXoNK/sSbmRO6B36MrRFkTUkP3MsqKWFounGU8n3DpBcvO2
CQe2R8MY0sqDbI+tIEHgv6MtRfNOfhhPedmy4ytUSlqAIU36GxipUX8WH2tyk48k
rJVUizsRg97GS83/uJPsXObty6Oi8qtePczgKM9KR2xBToIdbXwyj+R8K+JKvSNc
gfFZLK+xCtBkSUpits8jq2yzmzqdISEPlLxK00xBAk7ZoE89bn44OuDh7RoLG2Vq
HZuwkSzfKyDgNcoaOgS6BpIU0B0Z1dYPbsgCKqukWMrnqOR1+zqC+OxozLXIzVEC
jpRpOsJsTY4e4MnfJroKP9cYv1+gKmSeAZ+pHJ44qv0pr4E5yxxCqxpTCC+a7OxG
p0zfNbCVtUKeW+Ey+hUrCHlULKEVIFHDjJO43GaqaYBArvUzuraufEv+yQ+3I49V
rSUNeuL/bW4ubbDYjAPb01hpjiuIOT/uL7ycPwbrZ3fpVNauHD8huNCNgQpEGpFM
j2di8hczgWVDQ0unwbEcJCAGZqE1cwK7Vb3RNYIKdwNc5kzloABad1/MMncRYUjR
JKnC5W34bJtxaEA8+sJyv17Hk5MwJ1tvSvcCtbxeU07uqzNMEX7zBFgAPZR4VOUW
Ryqhpiqq4dol9uYUAqmgXYO5IEi2bwLGYQ/71E7jEFkw2V2A1Mp5UaD9wG7tSU7T
5gpcPF9eOjRXBNIif8rKFQ17bhMqAarz4BWbfn4U8KOqar7Qd1kjT3Tbo34X2sMi
hCbxw1ybVpxnlnEeLZ+xkJRlZVNzyEDhfp5tjVrUOw+DKvYzWYx+nM5PUKIave8i
f7e2oWSiIP384QV4MH9JJdQDpLkKHwBrwW3MtAnsEiV20K+fGlfMf1kUOmgJbWUY
CaU6dj2HVqzTI7IvsBJkw2RaGdcI1u6YecIJqnsvt21u+bTWU53OrId2zrgyy+Py
zRgjr+6INFpcIchugFMb1PQY3xE770upcdeoINUbvP5+cZe3CUbJrnXMdc7eNmX3
Yq+J+l4f1+GSKPDkymSLjsgCDFVmovdTd2Y+4kpaVKoMn9H/MbW2Rv5X6Tv+mnss
CCeztT5TCehnZwvzQDigZrPVXLFeJP90ZTkHV9MunlQhhjkiTDcPmLTgd/eiqxUQ
lVNu0ZU52s3oIFsuVexoSrWLYjnMGVNe5wI+5RM2jeP3fgY4CrugpbIPS1Zt5llV
Ma1J40dACXUH/3lff+dKTyGcap9+5SKDIydxLJbmLbxxMZH86j7ySZH3y0e5DFI6
veHCIi6jAwj3DaVDUlIxBPS4mbhnhNjsp+Z6lgUawOo7mdCcUv3Labqbvxz9pWK8
Z5qkGBnWSGUa9LP7EQVFq2tdSxS5XxfWCbUFkXcQ4wX6wYnO06jDqvsRMV/WeiZj
tZAbKAJkolvS0D40r9EDlCFeFyaJ7hKdyJw6MuF8Nl6DO2YYkFWrxmdJderUHdcH
h1fhANGbKdD4/FUOtKUC3R7GHb4Szph3q4grpuvkl2CdooMuNYZjfk1kHL73Y0lp
+TDMkGxqgv8TV+ItX/B0ihnPszRpZWpXAr+RV9TeOQrRuUO3YQFOX5mFwvJgmtai
XL9CmrKpkk8uCb7pPQHTwlr00sC0hTgrmv9IquQJbUoF5BAOYyusLP7vtRhK+9+6
e/bBVWzEN/2tRtijbjiHAlOAvnl+t2Y0Magf4iGy0PGPPWLT+kur/4vaBSe/r0Mx
v0xAOp4qe5w9NuOU5tnQqDEKd+RyLWrFcnahRFd07fvVZaRqO/eAV/EykgslejWn
gd0Zs3cPrcuf5zfT+wQ0PCHJeNExCiMkP0g1RdMfWEYFM1pxKqKbHuas+YkLBPfE
AJAIl13CkfizbS06/czm84z25vA6inanBpC/0LFY8wEyMTz9VLxpkwub79biWkCK
nd/sG+IJwz7YQPU0FyUDbAlnhCWEc5VYxTB/pXtgmgDf3ceyFKjBI3yjUNd+JD5T
kZSOxQJwD3HnbS2c1vWnpTdF8gPFciz/fVjhhq909q+TI+o9vjw1bcc5qxixlzEQ
P28W2ygBEfmW74gdogg3HyEvg9mK68CYqGK8TeVJtIiENivWpCged5GKzg9fjtDk
dlGHV57CLs2zzOXWvqbOSV1iwCu5ch+srHgZbHr7m7Ga/bOVcwYoPklZarYu3cf0
T14QO1P92CEnb3Y3LPU1Z3OYCDU4uBm8DjgnDpH60RvyT2NSA+yovL4amgTFzKSc
wYi3NxI3iwDGygIX6UwDyLekPA+V3ElPMaq9DZTHboB8uj0aSHJAliRz18crVQja
tmA08zWJ24DA2chEU1ZxIYlb6+abg2gNEzjQEq9FAzpjzIcUvV0gbWxlLdFcnXeZ
jDqQoIXME6Dgrk9O3n131ghqgx5jrkKPco8RFEaio38pmWSPL2MNl/1Lorcwdnst
Vi9fKkA0A0CsxR93c6CvhzR68xCRrT9vJKaP+7JIMCJnwnc73f5dRMojbmJlBYfX
YhK3W03vFhjpfOjlUQXnlmfT52px2+BZYw13aeNqra1EWKDuj6plvFEscXPqYPqG
TvLStvbwbq8k4+UhmpBUCTk4CTBfmJT+TkKSKfjAZTBR8YOxaoiBXdSTBpbo2/Cu
r6AhTQflSJAaI8y+gIvP9txM+Ew7HilzvldEOvJsON20QnbRbQDCf/uwmewzBjpZ
ZffY5MAexz4uihr80d8J85wP/KoaPDNokMSMdlByWwRhsUB34E+eY2xw7YOxkSUI
hYh/8Wnz7kuHry/9lMFLJcBHDDJmzr5vgS1RtHvkk6g2zW5DZkr7yNtSXLn4YgJs
KQZzk3x3+rAse+VDZQ5EqMuJZu0dP949wSYy8OhYxYE1iXOLi/a/ZdMAMfJx3CjN
a5DwH/GiVw6cYm8NYuMqvObTQ1U5ayuWVpIMx7E/1kEsyHpUyrnZJD1YMEZor9Ro
LZMh4alZjsyOJMyL3WaX1hvx0L8f7ItJGoGi2dvz1y8OA5NsvsZjCLfmShy6vuJI
3v9CniKexAQLy8mT3MJiZFAJKpxFjhsfQL7yRSGfwly+IT9H0P5PTm00q9Rb4r3a
QOgFk209/jSCYc4rkwHiJ995oj1HfEQJpHvoneM3bD/L6J46YHv/RmQXVde4d3gi
yxguohSoZCP3i6ggXV/XEpqrGGgoQ9wJn76txRXljh+Jgo6SlnzNL65QbY0EFoFr
hNukaSXfGnh5AAcSyKMUqP3vV4I7Hv4VwdqbVBX2dnouknzzKfj+4pKbOx7FDW7+
d3uV5MyjUiACeD1SPDT8xLZ3sB8zMEYzETunV3b5DpHnD15TVYDNueaXeIO2uqwu
BVLFnOSN/VEzrdKNNLV4FAYs6CKLP39ogS4OIFML7w1jx4QekIBy+BdJqAC03wrn
oRNuq7Sn9Dbi8wDM4hQK+eS+xFP1fe/2/fpGZIfS1hfJCmXFY9WsS+q0srTtN+aE
Q9wU2c+CC/QS9uImVPdmZks41EzXd0FE5ZIR1ViY22BxnHOjKNkg0R6A7hoS8Hvd
YS47WHWKgU4bCMIyd3f86T51SQKNg9GuKDVDE8Ej1C+qggMTpaKk1z3TJ8voONEi
IxAiugONEGrPj7ExZp1QAOpg/jIrq3HjzltOxKOiV33Mu4Z5NP+G3dExybTq5Mgn
wf0VJpBb546kITYrQrvtkwcKL3NBLnb+s2Z5ipqHlcpFu9G1mQd8/U1D0QlqajO3
zbd42g+621dL0pjc27dI+rsXrtmCeUYJQhcZiCyCMtcabjBMC3XA1a6bhdzXMpQu
z1jZFrA+ynwyPxVZLLpS5KiefKGMot5z2ahWHLQYqoWJg0cmCYd4cxmdXl9SaV4+
cOofDr3q/ketNcXTRJfFPeHVv+nLd5TkZ2GJrqq92ABBEnVhjcFSO+2SZ9o9wZ9Q
i+OL+R0niNPt6OQFXj8QL1wNmpS4cA8f0anCAoMh23OU34qZv7/6k2/o9VTLsWw/
W0//1xKxqdbzF7vxapEemN/113Vcq5ORouo/9skjpp5TFLOr45ksF6nOqZexAHOQ
VGp7NKnlTfW8RONguY5GWqmYyU1HZJn35lbjq6rWQ8VTRbtgdVjYYZz33KRonAuQ
+aOQiVf3iiCUdiESDvR6kQHx+UQvACfy5dI8vJLc5F5FnBQnN9VcNcNJ4GJazvY7
t2r1fX+w9F5cenLPoUo7EAEPURoxenDz+DAv7RYfcP85gJbL/62SoA9Fyd7hnNQQ
2NzdKWcINg/9Zcz0VB7lwW+hd+JcgZV4rBE4MGsWLMSPGunBnlOX4pGtoj8inkhe
wFY7q31f/sOUCBnRc/hGMIk+SdZ4Fi7WH1dtcArB1GNTP69bVcwpuoO4tO3OXwSp
VwZ79/EksGnFpi944qAl+lFKQgdpBHzXeDeSNlFUNWT1g4OfvGX1BFh5ZI08vERQ
DDjCFAzkAhlhCGJeB5p0Dfvl9ebrNXi6jthjvStvLFoDJ21+9OjJDU4wuIZvCV6W
osq4B+zo723Qpzi4UXvfsvo6/bR7907ilm+/+GYU+H4ePvcyi1iN5MhzIyrp0USA
OXk71+TVXpKNX5r8zV1fe+UaYtLcup/wL4ardYHcQnWNo8/JKritSDX5gJewj/Du
Y0vftZC611Mwm80UAXCoMs7V8ctcV3tS79Zg3rCSKk/KWFamooA02MlxF6+NHPWx
1rDfTpLVi+TZn+3GwEbqKRR3hm78aDHSsNx6pB9BBI7ePbkzhoJLRPzdJIaa3kSt
gNp1JCA77HJJQQMdGdBxTVggfsRSAfAnNyuViMgBlOMaN1JFPsustMYkq7K4Uijl
3lVXRiMXKVYS2dYzRUe860WbNvlAai99El9uKJe7tyRtUEfFQX3d9+YBkUA6Audt
EVRA9n0BeG6NdPQ43Dp0UqN0Fw2vhXMeU0fgI8Ca4gKiDZ7W8xpC0wE3IHz0J6KK
SnxrGNESodr3EGMnSPtVL2TiW893m/w5a48/2rt0pw2K7yFOMqhPbwM8nNUv9bsg
KAGMTpxnKGXrlEgz+uIRPmptYY5JFW5ttLY/zax34xJYDQCaQBvl9T+/7YLYjGe6
qvZa9n7bWmI0OyBah35CXEPMXu+JfFYPJa5VAK7bfRgxCMyZNy2oRKqvdnLCl0pG
HsoRoQjwJc5bCtUoqlfYKBjC2b9CzKz63+pGQO53vgqD8sCfXVhdBiU1wuFFB/Ky
g1CTde0/FacjS1z+QVFMl6gOkdfxGRLLdprBXDgBxwOmZ6dGOuGXXOrIAuzUB2HB
mWUsb3cvwygMVVado/MYFwOsmxCgEKaGJCNC8GQdrd9Kr0L5UjSMIWxi7NTjuoGY
izdkQ0eDgiZovF5Nfr0LIH3eEX59X5GARQeBLGcp7FEiWJ6fn5x6YeTYTlnpjadB
8blnU3+A/wmP6dB9gbI5a4AZmGBaWMVfvWwRndQO1DwVf74+oFpzfSevMnvFSwWs
ANEsF286TXXCRMQhYe1ZUzTfcUd28vLuDWgPkv5I0oZrWTMi2lnYG5tpGiINv1Vw
sl4AA3jaz+HFGfccDGyXLbgVNrMHiKl39tEdoq2vME9M/4S2OKdSU9L2WiAXukAw
ejP9v2cMRh9ZIcEmMLdG9Sop+uiV7gyU0K0kvnTfcLSmDEVcEErpksWNvf/QlG9z
3Q03Y+Rr2BTdaGOqzqTho/2TLPRRYQEROipx6Dt4WJlCV7wX7rMFg4KERok6Eqnu
nB4Eiec2M0aJz2+rEIQO+9czNqhulmhjk4IUzw8VPPPsNtaKd9thhTHxVY7LgLds
yuTkjvJK5B6T35JKCI1k4vXrhUGswZTbh9CbJPT1WT5I3mPN6pW5mEGDgfRNgl6S
KY0bxL7jjbfIQFYG8zz/gufEtKRjRqrlznazNuRrdP/qaDAwnV6/SyXzK1PmDtXT
AJ1Y79/pE9fvTrtxIU4lNZFCjMZDTx9eiry4NLm5YzIb9w1sQx11ADS0SXfHdVbG
vbaeDhDZYW5ViX3vvk9iKx8faLECIB2PFUUya8SSy2lxDDtWBjsA0c7OYl6mVGq6
5VHIgl0Gpe+eNdOb+XUkgyPY4l9WdWNP/rWNxCZ5vzPMHU6GIlhsvhfLHs3GH/tC
8syCZvmQsuWr39NdkuHp2YFvCNP9M97mt3ueyIA2OhjckKRv94yq4E7daagJxlM6
HWX21o6D3QH2DPUxedR0awCSHhdcguwepcf2D9vNca34BCj1hW3kqgiZhLpr4JKk
dhiFSrvsbDNc5YID0N97NvekwABeRybvHSkQb/6l7oXLqmPv2q5UGNCb0h0iT3xm
naGEXFHN5fnlqoZRqziFK+2ygUGeMWg1r8tEK8ZXxjKL1egcl2MKtfR/48r+o/x9
cXL0CnLYYdp6ih7pjrQuSI4KulQjS8YasYuxeMmopvigt1LWj5YQoeHHA2C/WgBJ
Lno8RoHNQqcmXEzzdOc8vvr0c1Uc38jxRpBbCLD+unvcADwcjg8syhM2QHvVrHm3
iZOB5h/o/V1O7SYfJxL68BKHwBQbt4uQXhLFm6vzrrLfizyu4f7cBAwvZ/suYkHM
RHIL8WuldvMKaojmboeK36ElDQ1BjHXezYDhw+GuIKt+XIDhaz00OAmMD+7x9SWV
X12k9h2emYJZNGfH7OCpKsTy1c5C+IINddaeHcDXos19Z5577qZ/D0a2tNXOQJ+h
PjGO5Dykc7Lb156wbRhDmPQzUQl+RMZX0qTCzfC3+rqklH36NuS2KETUL5/aQQsL
yMq0VRQ0GjpV6ktySmt1esXqhzYwT9/nWVHC3hzdQmvl4Z3CkJI1etDpYiG6OtSp
QS2pqpuxT7s+sw8waRg2gbvB6sCGsnEZTiETBUBvwMRrBFiPKc9m9w6sb1E5eevq
sE0+I+qPF/9W35AQRQ7d4YTr5k8yQds35vUgEnhEoFqZFwGRUaUejDccf48Gdwed
DICzEV3lfykvajzhk0jSUrfE0vjJ0LCNfMfxCIoLi96ioxavb4pzLnFvTD1fJiRa
8lh4yNKB28234VlBGE/cu+KzmoMXtR2/aYxgbo+3KgaVCv8TF6R5xfJcyeZY+sv9
nuKwBXLAOigVeMWv4bNAE1S9o4+t0/a3mPivueXq6pRxbWLZHjsyG6IWlEhhqIMc
z5Tg1XpHfGm9REpuFxghcE33JfqgEqUvMSDSx4t/LqapjzFsAe5pbv3M4kbZpndn
82nqbjpZJJQRiCdk38b6T9aO5oNYreSoxtg6lwIuYiZJVr2lc/QphLC5jNTxoGQn
JbbLMflkXzJ2dr/TbtcHyWGmhbY3bN4tx5zV2huQqLOpp1Idhu0KIGSKY4qgyXVr
BcxzWFJ8hpqGmFcJ3xQQWbcW0go2sK3uJKXCFCEFmAeemJ7JOh99M8bPe8RWW2L6
nKtJ6lzDxE1WmrALfl3F/z8O7XrDZvlzgUde9vlrtCnwbdVzMzYLVrdL6yvcH6d9
CgMlCDXmn3D9FdCeWluB/1jTMH0RqJxs5sm7dtu51EZta9n0EZ+dBrPKy8+ShAZK
HyJuEv9EcBqGmcnMN195iQYtURbNPWg2iABlZ9QTaN8hZ3KPjny+SDGEY9LFJTSy
CDEpd6lXdZmeb4IZ3siYWeQjaRUQ/CzhzeNbqZV9G0Wrjm+fJdkoBH9oNoBDb1Vq
IleFYhTy3+JvI1kH1VRzv1I3OWv6nYPFjD4p4nhWyqPB+ZQ7MrAy834xawuFVEf6
itb40Vo7AUpc7cvdup47ixF+CRekINwP/nFWJOUCsiMOZJ/NV4APHOJmTV34dmTx
86uywaeoD+te/wmAoKhOFEornamK0KNteO3VbfNFVf2pkj+W0AEqfXsr97KJqXJG
v9nKnPHvM83um7GKT7eVfPcVznoeISupiCZ97ZFi4qD7Jj2DGSu/LoaFGMHHFaJe
Pmo109axhpWhxFwe6KZH6xwaUglxORWVKunIHsRqMo/+5fevRmZlTCwKuC9id+mm
nuitMWZYUXHqVsOHpuwTBBwmHXjDoMUgfF7P1DXbWgvHEadnbzJ9VYYX8tJ2jyeP
RRV7hKtdWkSI/W6T+Jsn3nWlSKdc3znm4DqiGzjSPT2DeHS7pncjCl2nCRHnfETp
Ka3jCowcNyU0JOG0NZ1yw6nNIDnSCCGAifKlj19xSODBNj+8ZO0+NpFGT/4UueNy
YCqyK8oPcPKDcH4kNIUSgFPviJsXSMYKpNCUlp44GvwRDLpWR8wHDweXsMAMvR2D
g0CxqtVCeOS0sYKgq/qDJ6+LQGtwyLfsI3qdp/b/FNYZLk83VUSWfSiSs5MbhuAA
jkWc8vAT0YsMepFrJ4Ua3UazgHGRVmr3uKJw7r/Gy6ChHFnpG06P1FCAKCEGAIcc
lBpDr2GCv/mvti2XYSmI7w1dQFiWkm/qyfl8Y3nD03irCL5xVWC4ooJzKxIgDpJ+
XiMaIdQQC6M8HteXF8fIIXbIbtULMWLuH+3Z9ZdN3jSuT+ZutxWL2ECDL5gnIElU
ZvbGsrotQ1yDrU6D00bdMKJjDW+cN+tfdDhYMDMrm89Xs40UhstBWppYvn9ZJQPf
X3PIo3NLe3IJBugjOVIwY1tst6NYSkRvAJJFksnrV7stsg4eBAXiWC+RRa0iJRyK
8RNTLa166foe8s54gJGZEKi2lOkuuKYU1AUIoAvYndwKi8JVo5fjhcIfqEYRXzNT
JnSyWAKyndGVUKTviNyjnDvkJpsU/4ngcDU1on18IWQlBx7ND2+vjv9PPt9tzUg8
KkaQJZcJ+U0V8UP77kcfw1yGiz0Exg1rnPPBP+pHsmBN6OPeZllVljlTeZoPe8Pa
Tifq29SalDvLipMl3DnnozW8LPGbOpRb/s7QYeXCV4q/8Hrb08qhAYhXjEXKuWeZ
3H5Z57Qok11h2rqMTcEXBw4UWiVWvU+0HV9xuy/TJPb6pNBihBP7kd6xec9LQHsy
JvXrE/LlyZ/pkFXQRouWKQNdnw/Cf5lWWzZ4NEkBmlerNQHUF37ZL/gD1AeaF1PO
QPs6Iiai2RSY4yahCVVcW0fAzm6Mr0jtLlvAv88xAgDSk0j1kQXn7c+MJmlSFnfk
G7yYkOpQ3krxlRpuoCrZvk8AeR2M6ijadERW/C9ZIgtBjpF1RJSwM8WdEwnznjMf
CP9YH/qSzH92HaSErvqXBTfZlew46YgwigOy3Ogh5h1/MgFiytWNborgGmy/ICx6
efKW7pGDjB3z1UENS2AUHJXmM+2WBBkNr181qYq6OlmkJicw0hqmqHDutqBwafy9
fwxrmlIGm0xxKJwDyzkWlZXjKV5vuAek6VjgtTL4DFQWKBKUTexf/aRVHNEPDAaM
YfkeTYzoZVXQB24NZou1E2WRBp+WQdYKNPtchpMW+CppQruB6HliNhfl7A4/oCh5
70rcY4L0fqpuQdBvz+H9z5X0wPKnmVvfOiZFln9+M7C71mZyt3nPNkLxq2Jz3+GL
Jzvz5/WVTDZ4UwttprR++7kE7A7teJy+8XfbaXB4xO6z2u/VFYG7qi1e2q82lJxv
mpPDNMh41rW1J/xTTXLjRtyVQCQ7FjBydj6zLP5KtPoOgFEMhEMcd4P1tkbCzZY4
U1DtFqpD4MmT32eaQ5FGCVEHwGugWIYOtY8WYn9ARs81fWdKKmNZSq7el62BFtha
qSPnzN6AJ7G8YSYXADgMj3JvtzcSqQLX6+6UCZUYW4kXo/KBcrulxVxrzr/FsvKr
wFzD++BRXuy5dz50tQyxY5ggEDWqYKkcig/oYaxR2lUYFq8pRKpg3bsJn6fMbsYY
0cRhjac4tI55gt1cichx0YPqLT4wnlXPNw/cu8XADvjRZN+Fy328Zq7m0IW1mcvd
Zk3qTJL76Qi48wJ6X22zGZBxQnZ1+MZ9ln8T4ZSVzgCZxP6Em2OkUjlaRjdRwT4A
brROTNaF1b9m/Z+fQdC+5fNYYdH/YDBacUhAnW35FWuEcj6x9pKf/IrG/hJ2TTVQ
BXARqfE15EGpsOCZujF40dmi/ShqXUU6KqoGoNv/c8t64EXF44q5qJhHh7GxyUUb
EX4Gc/pvaXUCCjU3PEh08GURVeMJ3JYZTD8ruk9yepHnhr+mbo/MjOTnwEM1utsq
l2NwzgCuVMTj9azxGrty6S32DGGjDZE9XlbW+F7h3kd2wiD7H5mvnomS4ZJ/DHvu
QY3vN0K5iiRX/7grPZfzkoNZii/MtN4pTi7LNbLQV4bjBcm4ej5Kv3jl41EDdgIQ
USXWvRxlvW7dchtVUnylKA9dbhflJNcm0o9soNVwVHDd3ik71/QkvFy0jk1a+3fi
oWAXkLFt5f41Fa6mggcivaSxMYyfUT7TLErSXNzDolLq9PDFPziIaILfbZ0fCUx7
K4RBwEYW1L2MosD5Wfdm7HfckCS/QWluSyOXWe3GXQ8ppmmTnyD95+PF1v2y0t1H
MTQb2wIZAP0oxVmAJWMGzzn9/eDz2GMp1G/R5CWJd36LTAePb2z7ArRf5OnF6XUZ
UKy9dRzp6+Mv4CRg9NA1xNO+cmHel/Oq0f3+//HCpOC+E3jUgoCuE+7diJFsIqRV
fmumZ2dIbm0r0rR6UPTrQs6ZtTDNEbR0Ka6wOg4NFhQ3RfPReDzByQ9GhFJkdtx5
1lkyXXvPsfKzi4hEosk74Qer7+QFm3ykZlcNGYnJDBCqB57nfKHqgNKZI9Norgwx
ksbUmGOYJl8on0E4VS+Tru7BMomln4MiO/l5Mw9WEZyiALRdeSlHEdiRy7kCarU/
+Vka7v0weOaW4AEjLglvuto46njJRkp9AcPKnTY8ckAOMDTKZhlcOpmv0hzVRGxw
u+rE0Yg8YNEfA8oQlvtCR4pRcLx5ARLENsJmo7MSUlfCcGoxP0CXQnD5egk7jZhY
kuRr2rs7NCNUxAP7zO2hHPxfM7DziVUOXwVQXYdi2x95wl7i1VyVfQd1YwDillZl
PuEQgU9J2U1IlOgjr75k1RDssnNGcvVaJ+uflpROwA02G2jg2C29CJzc5+yuRwds
5GlSf+GTlf7esU/AGFFV6FHpSwnQJTspBqbq/m6sowjPySEDc6/8K5zYBxHSiAJA
Mq3fnio2OP7YUuoruF2FXg+mv/Jgc8jb93mBrB8/gEtk0FeRTI+T3gG558dTk0e1
FTFVeo6t9MBPQ5ENXWCQVjfqxZisb+udCxmF1lnUrzfn9eQCQk+3Fx+bjkNbL1iG
mf+DauRbPD/xOmV1Rbahg+DaHHM9KrZTsm2mtOV6xoX1XxziYRDq/Eozrax3Xd6+
vO9/87OG6A66Ih0NtllqX5GMHh29Bsi2KmChJEDiWu3XBPb8+1GIK0P2GNBVMq+0
8SNXcCp3xpIYuqJ+1pXb5pOFnyRbTM8XHFiLKbqd3ixhfmrpoy35ZuXuNnqs5ykg
YZwdr4QM6uBQo2R264OscMhPRp5fj1vTBvMupqIZoN+VJ8mCWgRbicLKB2bqQouk
ZY8m58adTGoj+jRe6x9n/Nj1EGbF1B0/DFZ1KBUM1kbYueRxxNHJQOGJY/SfvM9b
OpPRE1ZqbKbb8X4XHJ9b1nNduKpdIjYa7Y8O3hD+Lkft2iuXx4C1lIFf47wMfEJL
NHMqpjIQcgK3nBIHqaT3e8ZVTQBI2MBtifvIhbwyWjSQnft6eaogho8XohlfzHfO
+6mYwBvcw7qFA0sPnmZgqpCDX+TyjynirIB04EZSEuEctybbe9WItZUW6N1s0/wO
Pxp0JBTDtEXFgdFIpOgrCtXsiHgE+dislbGvZ/52blCFxj9r+Q42/CGcTBDLrhLY
XaKBkA1r12Sq+5bCfnFJi98XfP+XacLWHwmAFr34xYz1HN5vOBHJWy9HXX3Se/2F
V6sCNbMpQovetOiO5tb6pku7YjLtmKFlpv1Z2W3xABsM8usFkfAX8zI5iJzCHSWA
hKdjy3pDOzjD9OPCR54Nbmju/2TBySmf7f/U7hbXNF7VXA8KSFbxyrnU2+Riw43Y
86sr9jTNFoleq8HIJnQJhciqvpNKkGsbhCUiAgrEhdyV7s+PlGiZsjZAFqsbPogF
yCnTSN/fpyU2FaY9cgLESPXC/wPUsD8foSYImg1X0rwtbgwsNiNaw2XLMSZ50J5n
+weZBXnf98AdCdNi6w+9QM/vZ55CggzJvo0igvwQTLT1OTEdJX+6XJyx/oP9yiM+
VE2xJOn9S3gIdBtQGQPBb+5c7fVP6VuTj80WRggSICGx9eKVlJ+8+Y+ZgEQ6pEF0
AMfWx1T649FTPLRcI6mSZaTJmArP/uFAIzUF7vorLR/YqDDSwJRNRGV6Z9PCDcCE
K2hjQGpum5sWsqxSBYM86YOpleGU5UbkvqSUazQXr0K9qdJimwV/OGlTD9qvLEsW
otYNggtpntxMpaMAYypJU77w0uQBKwukUTvQedlaDN3x2+mVeUEzNFlRyPz02TfR
0DJoXm2AgF8FhxpsijkJBxDIhBmtXK01rIZjTZFWx53vTfxrh8odx7W+I3A72AG8
OrJp7EBdLJORZUewn7W+hRFEUyz+scDW3ybA4xi9r0pj6yxOzY53+HGZiUktxg3t
PjZZOjhDBMuyorcXtYx5m68otT99I+OK3EyPtJk4FjadBPUjYjugeTjY9jM6HWc/
SdYCBRNaLY9ejQneI27XXy9pWfLfpj9tRM10QPb6rUN/QU9ngiCR65Ehp2oXXZTW
wwt9BKewFr59YSG9HuMcP/3zN9JyYBU9aFCV/0x5+mWXFvnfe5WAGcrjSJtSeBjR
m72E1xrY3fR12LYmDobvtPrSyJF+Pp6BdcdCeG/RW06FTsVSY1W4nmiQ4FNe94FE
QSCQkaJ1n8P5RUJXpPSiBTsG1Pd/bpvu8IFSglxz22ez9EgKYV1gIWQN9ucIonuX
uvCOsQYtCrSgfd0B7oEhYZHwT188fLc3uk7rajT6JjljqtOeguTi3dYBUtPXxrED
jXYwJDXMAKpSy7Bj+vgGunUY0FVJ4pSBld6eu5A3F6dMIZD4aCoqZ540mAeBL2c7
lSSGGj8kVNkJ9wefFARbHOym+VOJzUxieT8DtdAU/T9oV3bmwpj0WDYZRYGhSTAK
tFg4rty15kRQvwgAOLiP/KoBjgQGNcBeTmHsBJKSxV2ydAZpXZI9AoDCX0ujGgRO
/UieCPnvTGO5qE+cskGkkOAbkRz12A4Mq1GoUl4ayGXzduYubGWwhxzSfjpDnZc8
trQZRPFqWJoHFvX2P6Tomn0NEdFKK3FImnKwuqZzWfnIecQG0i3eF4NkpDhypUUe
nRpqydD31M7GRHa/GrkEvrkyWlIWvt1cjftktt0unCSo7+Oh9QXP95/DxmgwOHUH
2WBdc7TAOR4nzX+cZlj5cuiUeQ8p5qs2hTwun9yVdOVtgDKweyx2T2OJNYaSd6cB
5l5FE2pK+51H71XE+quU1Er7wSIHI2g7NQFV9UctypjXLGarl+xHIF6h+JKnWqZq
FKM950owcZxroJBxQYeMIUPf4e7W3wIqxmEklCOW091qndafaxuyXM9G8Ydj8kyF
lwc76hi+IE0BwBi9nnfBckuphvgo+kWo4G5tG15mj60PAAipcxVYAS0+jboqSycm
AmDNbqjgH55cMS/NAx39GBhKxgHH3nuwP7p0T+ulM20dnniw872pje4kTHbhpBpr
R/XsaWwpk3INP7YDxAn7KrmjPl4qIUgHPwNXTp2XVMsc1DViIu3x4FuhrNtP5xyW
YXk8d8EUjYbgcHd6HhlqobJmM5RjirATbSiizymvudd/2tIHp3Z2pL6IAEbzXgYv
TnL4l5u+MUMicM79g8+mf1I1uiAfnoFwfekHKswRyZxSPHVzaidpI2NbnNGvytVJ
AN+E+pDSPBmupKHrC9cLQaEaLhhByvZTNy6nWpIDajsK9MgNe9i+3YGx+Cm8aUdz
g3XeZJW68tV/TqZAKmdU6gZ8uCJwc/AfFIXFn2DvTw0V9KI77xy3twz3ug36+74x
yJp50P6pbA2UOc9xYydFKp5CZ1RTjnJfll+TxyZyZ5SwT8LIAD6S4fv+OSSZ1g2k
bG38DQhYRBCqTPkl5ewNHBJaL+n7HMT1S0c85aJrMlJNWvCqLy3hb7Ya5E/AeuBr
+2RZ6s3u5dI5ZVCKNUrCCrq4rIUSTbxE4v3vZKUjB1bccAEP515gdAuSpmAl0KPN
9XjhX8SiT0OOaTtv8uvdUC5svqs+escP46keS2V2JkJDHM7Lreqx/lrVq7hSHYPa
XRy144ASe9Rz9sjAvw0jNjN/b4+mr5eOf4TMbzDzKTgjWkeHqd4KKhHJkTExdkDY
Do26GyldOGBbqu8hj1uVxmYPC7zpyGdTD7lEzOBxM+Z9SbqZnBYQSVmUz4KLVx4h
140DVKm+MghoFXD8upfLrDXOyejck696O3GjIR6fellV2GeXVQO8zNKuezitY5w1
Ds5YT3tX5AX9PG9V1I7LrcY2Tp7qRUs/1/MvYpTCYX8ZvFc7sNVOglazZMg6x0gL
XozGRMX/H4MeXKKhkNtl9miCDM5+qe4/uheN9ORQzuIU0G58h2z1nrDm+DvTciP2
jxYTWwhcGvGVvgt1G/GB6oBjf2d4gjdWfiSaEn6uBjs1fU+7hereIID13BiCI5aP
5TInqIRk5i5AKSe/3mdtfiMXbUYhNxLPCDS0jVeAWLVI24weP6XPRPKUEUI/dvF3
vjxmFEWOO+fPX5uiMZRJXD9SPLm/ONYiVEOfGcxcorB2RTbO6+AU55lV++8nuCl9
qYMLrltrS/NSz9OVNuZ6gWfJ2SZ9EvvZEbgi+NPzB0MDkVyTpoGI1n1E8yzy8QMm
eUzK1pCCWXKp1RckyglzCAZXdgB/LSNc8MXg9IvvojeIsIKBJxVNi/hSOiHlYGV0
Kb16voPeK0ANTAmSKTRfFSygFrxnpzKrx1JQrxALBw9CIzAhEKxxCDzwzBIHFD5t
IbfUX4H/jtJYhU3ya5gKu2x1gP4DOFGJIUIQwd9ouzuLp52x8qpP0qNE+ijLmBQG
2WoDcoHS1prjBloErgbx39GKXmWHCbK0+SeV0fTA2Nz2GC9hy7QuP8r989uqGdkY
/BUHamkkmINzPYgeWNO4s3GlPdmWAYX8HVTQNw4W6df1/UCmd9lYzu/fCnNP7GIZ
+J1o+XbbAMUXha/bXDjxJCTzuUEaRdb8Ac5XQ2wKnhlrMEdQ4NvEqC6VigsDATO9
NPkzBEHKFlHTz5vI8ZGAWTTeWhqaKDm5jGr5TVFYXaUOlLMglcK2JznPN0st6CAQ
RuGXsPgvGHzMinUuUHBGVZRq9Pb+bHAmTg9azoSHhLiN20Kv4c6uTy4Yz/jc28/W
Q+KYUVHmSVDtrPkIyglViUj5Uu0A1T1IerLtDyh9PlvdH6aABHhQ4nQpkqO8/Rrq
9WhAvamV/aOXNDmU0WGJJRkhZe6v140a12XNYxhwF4p9AivJT/A3FkwhcICTluie
OPo1RvN9dmGzNFU9zTAgpGx3CiZR8CyDwH9JOJr039pMcXPhTavMmJXVC3ZDsLzs
jjLsq+Cxpq777R+23/oB/RxMFFLknj+zUT2aYO7Prvu8Tz017l2C1gtDnuYZq2hw
o+3wcW42OkORPyGogHMEUj7zXz8QpDd2O7Qq+svY1BUSmRSEZgJntd9jvkoiTD1d
NYvpbmo8gY5OPXbYEeECN5bcD6/TdyRdWkqEgIRRaF3gw6YIPowgfCKWuv1q2GnZ
a21c5Zg8S+D64Usjf79AaZ6wcfaqAAQzjb9//9y8QSIKGMRS5t4/p24DTbK06NR6
gLAiq4/DD6C2doMxhvxy1YfesIz3Ovb/s97t4sxgeJ73My1+iwQfzAnpp3kx7WP+
IVCS6OFzB25Td2U/l3QJ0wZcAPhrvGm59JEJkEeFIjDgBiqCszrToChqQHSHg/dZ
oClnCyncuEgZu/MMwBPxurmWbnp/it36mdAVHKlK2/nW8uTXQIf+QGCm9NiQpoai
v151ZYnj1unqGONky4o+2XJx3M1Q43xJ5EmvFTYkH5TVOKDiUNLGazDW9s2KxRbe
vEInRN/+54YhA69tv06O4QthxznGQXxrFX8Rd/yhRLII44jKCEVn4kTjrpXyvznG
jftPaxdAQmOunJnTWLLU7LoWnYE4ayiEj4/uFHrWlA5KQIX1z37q07HE0tf6lMQL
NcszCHx9hbzWpoF60rqxPo4WbmuYmuqGyrx898SHDikEo9fBIJmvzaeHQKcJzALH
n9qy4LMt0MC5cC94ZH0H+EbuPj8K4geNJms34H3sBXOu/ww41/3wZvQ+sHy1vC9/
2NEGqNiKKPDIiZnLSyIisT3jF4F9ZKIff0+Mw/rowGXSR5YRe3MP7qpTvafe8+o8
ILfpYpE/jYyz8aYH9I0tJWff0HojC5wW7NmLkzSUB7w+dOKLp1huNICjfkyiI72i
AiohYvOWgSjosTkitOd5IgKHA9om8sPoKFBaTprEdAmnntJEpUsx5wPGQ9asa0dg
eKXrN6IidTT18w+Z00EhR+pg37aCOfwso2spCAzxL/s6cR6hjk5Sn80hbUO2iWV2
7UDn+Ln6HjDuGDERisVRwNvLmyrUAOrATtwdcB9kQe4CtObOcaN504G+o8QLBZy8
gkRdgSW2IvmPgi11DOOqGQ/ctgw/iF3fYdnzhj5A0LvsPD/BMwBNXwMbmxQOCkPo
Cj9kLPfpUjL2T7pdQae5hJ+1dvWxm6pbihnlIlL9gqDJncW1fAPJfsp282cUncXS
tfxlWPY3Qli0J/CMp24dlU6+Oe40T2BgMY3rNNLy1yqi+RruYjusj24lx20ZS9Ul
b2XG8vfpiHC86tLPwlwwTUl6EN9jdz+PcRrNH6tbVWVgPTQMItQtsmA09ksQi1/3
Qk86ENuRD0aIN2OPPHtRuVf8zZDrNJn2bnVYMht+ddATPmuj+HHqEaqVB/aC/mhL
hbxfIRxAfH41xG9H+k4INWc83OSPgQCw2vPFQyacfDkkv1+taMepaybuFw07dHTI
UXjOoWyNsXRTKIMoKRt2bNmp7602bzHJ5qCRnNqRMU5f5c4BUqIhz5Pu9wYOUOuC
r0tot0pQq57YiBqUfOBLx547IxgwBAoarriB9Bcq3YAZZHJd4oE0OnT5uK+DagRG
xlMhPQfD3dKpMQizqxIY6GO+cV2bUwvBeYkLaFZ6T2Kcno4SwplfTScajC7Ny5Sw
SADjEk/+Cl9fN4tbB4CLS1dvcMddOn/H6No06LsNTFJXi+jULz1LSwBQt/508TKE
yW96skKBIbFOsWRos2W6HfcyGd5pLBId2EtgUdbiexh61DroSRdiPkw7FkW2MWEQ
UMb2tInlEk2h/7KyFf+tYt65ZWWBjZVVx2Wr+Ir9Y+huv/+6Gfsy15Az7oQpzUeS
viyHi1mFNRvyx/8hEYnueoCglE+DLbZjtIA6ebpreC/fsf6A5M+kB4+38xRtX3Un
aUD0lDUf7qnPjBYh3Qoe8LWpHKjXlheTKIw1QPLeKHbzd2gnmgCSRYQsYf+BRvmB
mjCmAYpRFKTkzJFzxd77o0VkUQ/p1U8jUNzkUTDl8TsuXleZ33uQqMg5kIk9qHz4
JljE67XhFSqfPJgoOGJku7IBuRbPQ7AUTkv+kmvUd1mngBs5c+Gf4vOlF98eTKtA
5zn18Md8E/pedl9ilqKBlBhTw7LH3stbsjK/VOVpkJCAUpNBxl9haF+1A9Ppz9v4
WRbF8kG4XQ38jW0U1c9DESUsARywEnmVcR/eWACSGr9Ov87h9rczZ1y1ZlgULMV9
l7zLZfsVI9MKNHlGaFvg12tr2aNpKc2+02t2GZ9BTGnth+uKirK2pbBnnYiGLeTm
wEyftZuuLCtHoPYwTsmLJdQZP+aZ+W3/NtRtXLW3wHIBtbrCHt6AVzWRJLb/pnzF
CLuSpHRZbBPoo6UGE9Xb1xdbWzuz4SwwxovvYEbxwoxsLMZ0PBvQtaUJDWjFS4xE
129Iqa8RHYoti0W6gMAJhfn/u+Qs0QH61zNEkaH86vR9XNPhG8playzSvKMRQHlI
f689TJksAXg9M2X1mgwerMCbZPhsyuLvIBlF+a+VLymZ25nO4MFuPEUTHHHxVzud
pXsRrhwJEtZNnCgHtkN/cmqbMuYnqeIFs6KVg/AlR9rQ3PNV9SXzLMmpeDNDfgeC
N5T2HI8DC0/1NjDi60M7NRyzoFjJFCmVcVXsUDEO6NYzJRa7tBV99jshHx7AT6Za
ciNSLevhr6p6Nzwlw/w1F4oSjTPkGget2ChaUxgEP5d+OH0bxpx79GTO6bnEnfUa
AmAZFKXtE14ku5emm6VoYqlh8evuQk/1MJx/RfZiBan/pev6TiAeVYbutvhK2wBY
H/wwngdcM7clOSUjt2ZOuwB7KUMIb4VbgrxPbtMkv2GytzE3i3+op8awa8CYK/wi
MWK3krgo4EBTXWYOaKQ2XNRg7ihiHe/uqUix/3Ahlm9OeW5uIspb0TN4Syx8EF6l
lGcMK8ib2e3zcu2+0VXDCy/6rIx8Hl1lTH+fqGWRe0RZFrZ+MJ1rVRPqDz7tNcGX
0w3pUeXk0cQvv1zK4RBlBYjeo/SX4QrsYKEic0GmbqRckWNkAaneQbGm1t/OXmVs
Ld8rFahMpBD8zO7esmf5TrKlA8xLqgykwFthSD11kUnRq98wHZH7j9hFxszx9ZGo
ItifFf0zuzM0j2NmOHcTDKm+dfDJbcXYiKnIJz40ZG/xiNkxOh8Xv8v92101xbGG
t2xkQ9f8gHmmJQUfupE+peKazjuKfKy1LZiQSkq0FuRTWxA+h5SemGtQv2/8wmdF
LN7deNo1jEdO8s4y/WjBlaOyYTQT3ffcenlhxHORI+q6bN5qr0KJjAYlpUOvO0vO
oq623u9grPFnbNoZNhrF3ZM6a7w6mCk4vFiIXYG/IXugQ1Po3Z6igimzi07q7xu+
w/CdOan6Z7jhZEaHlb9zEPNtR9Vjx8Aq89m77nrKOgRKj1G8dEndV7himtPlHXYs
rvytoL4FmxjAsUD3LS9fDBQVeyz5aORNwP5S8r4Ug0ugosdkztE6ZpYMB15odZef
FXAChuOtZ4MT9xOr1mefwueruDZan0XrfWlTaCQQSk82E7+t/Tnzew/Iwncfmtag
3dnmDNe5i95zhYJc3jhteyIMGWGfBtaW4V4gpjyoq57FGcEcvuX7NeLS1cRoPFyn
Vr8F0jEyDpphgzS0Upj9RnwZP6tgmENr+3tlcj8X22XMkN/VWTZgDAyEdB/4buve
5IGYLD9ZEcGcHmDtWT1SaEPe3lyRV1j86Ye1svT9XnOLOHOU6MxDiGxLyRWtUJ2d
IR4Xhe5k0ERCQBId/zevm8i13jgz6SApygNuZjKQjKA3MRGNjhQIUz423IE7xUed
QuoqJOZHU3iC3T/giTigg4W9WIgxMQafxylq7jNbs16dvemmC3dXQ8IxOSkcwp6G
s54bJ8YULeSDXAu/nNIukf/PqbsjjPl7wvL5TbRwBImJH7Fhj/e40QS00rqB0S/B
Ld0qORphBcuJCBwPgFIKM4R1sE30Q8aWt8YMtzDbNin04qCCBL4XExHP11Zl5UoR
uppko5yVALBWJ1zYswMTT1vP81AYvmhdbX6eVizHCGY1f8TVhlIBIB6l3hcdu9w/
Msfs+s7ImtLG/5hB5fgPI0Rj06uahOdK4slHmPuH13JIVvY9HLHG1Lcf9ZxS9V18
lyG+jTBekxhXY2ks487xGa6pgu8nsNQ14KPaCNsZQN7j13lHFiQpx4XgcVtk94pS
XU9PxXUaZTiy83LBYtHIlXjk7oCeQvTLUL9X/IX99TUo+99eD6e6kxZfBXSqRNdz
aPbWTpCUxuXWrSwlDMZw77RFfTlR6GlquVfX86cPtDVR3V1Pra5SzqkGdymeioP7
UySuuOb+wGIpgEMbYeV9RVc7nB6/su6bV+aNnrT++QY+28KFGVSY6QTttx/pTS79
JWJPZRGJl3OHuwR5DjTANUhnNT9fbwZNm1nD4CKxP8o9SSwMCKtWrFtQAYi6mpkv
Q3FT31trtHKnkCAFPOBNPRvhYGI1+cVVFe4xdygqCXm2xn7RWqfFP5lS/nqA/Q2O
oKCVAjVtds3zK6cWuN15e3a+PQF4zTtrR6XA3aTUgZX1UnPLQtKnOKIZdgo+fAlZ
twhdfNB1ilb1WQYA+TG5T22tRx0AXfXhJAbGmaVPZqgBSrnvvB6hylAvLKmRROB/
HvhXaNUskpvsbPsb0i0MjO9HxMhTYf1i0ourT42MZ0nMbdcG/xcXkrSPSuc1O6dd
yEDbocsjfmRO8E86D0RJUN3bserRdVjQY7lDKwv9am5ZY9ShjX36xwJ8r/HKaHS+
y5I+vDpWb4SXnZM9PMoC2Vpbug5BmK9aQrKM75FbiGgUkZ4PxxGXK0p5ZTSK2887
0/Y0kh+afrHJdbTuU8u2r7P20O8VFQlkBXWbqUDsow/pOkOh9UObo+GcHwWUKl7+
JEs7Yk14PDJXCCnjw3vS578oPwhfzcdV16SeChUWu4T94MBXmhWo3lGFtNQJoJvR
doesKOWWE3cyPZ8PV26ZgvR9OVOqWzOYDjurCrrkD25bPL45h7TG9mRQoU1ERA1A
bUa6iUMzuWZBi8yCdiy/U60I7A4GLNXVvpeJvlYL+jLvtqh6YTH+q0tihzjYfOW7
AtcTBfJ2FKClmJX8ev2lRDStV//Gs31kD3P2GUIBY38MSd4ZUlZcPivRa1sOWYc9
Z2hfPkhrqXGz1A4OeTvKEhK0fosdvNdLJQRT+62zzEA8uJA+Kqu2kDdOmOOb4f3b
G4Lu9fjRufaCEepDARM3P/OpGrvbu586qRBtMjoxi9wU/eikjmjf1u83gWtlHeP8
hvYpRaHvxVBYGuGtVCBVfVbpmki0nIOyXhF5jIkDpiqp+wb265iJP6mMK6hTt1Ml
jI60koVdvDlCerBxgcJFo2n5t/RkpuOOs0lRFYBhLhbXOm0PJlhPYoY8Dd9Qx1s6
uTr1yngDnzPWRyJ+E7y/29Rf45xG0x9m1rG/BE2/AZzsmiqD258GQ3BOzKVEu7gh
SPPMvTmlzsTehzAX7A8EHprc4VQ1Y3kX20qiGFryz1Blw/4oSiosDMQ8H9r/xmCr
/Rji1sHr1vCaonUaZuyyueHeCrDQ00EL5KPhUwi6bjA/Gv9pR0KaWieOMYvoVY5n
KmC44C/UrnoGqXMZijaoG85gGtu1vb3927tlUYDTbruNghL7PioJlrpVw0QYqDak
sCeN8n3kPA0uO1+s7Llj0oapmXp/ksAs2X3CJ+JH01iIgvAOGpn0bqjPk8eGieyU
fHVM93E5fgjHXm4wG5l5FaySFTilY9qrABLToZV86hzrb4QZQ0A78Q1A/3WzkKoE
LbXYey2uL6VGnTeIzSSCllD/3M7Cxyc4+K7kxT5IetSo/CajzDc7vCPQNkCyzuQE
BHESM26Q04PckG9Bf8s8FhU/6DaXYgXNcL+lRPgtAq6yP/5VhACYBQn+C8H5z6kp
zDAxFMdL3Tg0PdvruiQv1YmBatEh2jwMU0HD/6dVecSWDZdYeWEd3i5u+HG2bHo7
+QMoK9Pq2kL+FIV0b+7v+MGvc6UwwD1DSvvMFoOo0fyM+mdVUUGZzovupYtwmXiZ
r0nncEBOrqQ03q/tiudmu4GdB95JTKlM4nDA4WMnuFQGD5IGj0255Sld+dYIUZ1N
ZfUAo8cVRDpOyvF1IFlEr08FJ6ptMDfeJw02HOWQCQY2kPW79cxsiPfavbftoSjf
Cc8MRRkVBITbuImqYP1uvIdeL66gipQJcoGkinY3v8X1PNZUewGecvYeHs7FsmWT
b2qooPWRT8mF9Nn+06Ug9e78zQU4KOybbUxRMWly15uANY7PDdzDwwYECY8Z50p6
ZlNz1vIG+HX7uJ9aQs2dVoFOEgfhAZA5GgtEPbVH3BqaGAZKfgLeNLgRU9QWM+C6
elwffBvF9w6DrInKIPhbfWEDrjAbLkPkELFED//iRYW3Mrk/e6Y+050x1RFrZCbZ
bAXEYiONcZNAFlEr26/qTZU5MdZ5FCJN5t/eiU5sq+EA9xe4uKK0veUgz23Ldfow
5avBbIaLlAfa/7yvtHaj3MwGw+83EWfh2nnAQqyGh3zhgT1nih3a0EURgH1RONO6
hyaV9geWGnyQmN+qZu8oVdyp/9eR8mHj9aQQqQGDmDawSXMj8VJ3aoF42LvyNH2K
FGTstE6/lJ+TH4Ww9TvOQiczYRnXOWwnDbnqcjZOpzRB2lQEfClNQNb0hzXeNzEZ
bjSoymr9zltMO88OTlRlVUzbnxcUnxAQZWe8+C9sxq762vwanaZp5L8G0AyQsFSo
jVtuqwko8xN1DnPFeSv4b/6YXJ4+MiIX1XPrBSatxBbmE+1jyufDQ8ZtQsuL3Tvt
yU3OI3LsSzR6tZpFR/YJTLEA/H6UmNGQAi34Qhe36oLlCj6KmWWjx45xLsuwv8zc
FWk9/1sk2GHHSXnJn2Pbv0PAx/Lp+23i4n9uF6BDwQXYeASV1HLflnW4UzpDBRHz
qcNklN/pOvzcrvEL//mjS04lkrPa3vzMr1fFWFbpdTbq3qDsln7nj667ysLlUpMB
ufjvUKWIi1uzv1J4ICfuCYA36gX3QrN+eBMvFxBVtxHXKrKboS7OczuCSHQbuuZu
BlJRjLA+SQ2leRPnDktPrsBZWrGYMAvhozZ3p59Albl+hvbYLBUjA3YAnstNY1Wp
7lU2EgkGLQ1/qlz3n8Dk/F2BLo8rYQf06q0DdzjVhtF9+X2s8GgLJcCqu8FBNsss
T9S6sUYyEhRZ9KCsycD6bR9S6yLLkYiHS0fvQBr1qwxImyjMs4DcZcRpS0kMrBy7
9e0mEDgPJntHBGjSqRVwYlz9NnKqVcDwxNTrFsSHone2kI64npcuVAaBAdA3YHKz
D/lEcVoTTVt7gcslZNWnKaOL7zNE1hkMVBPRHXd6iXgXwtFchr1q/zIl/dBItpaz
1+xPODsb+okzBBTh4H86UOYN+QjGmz6IzowpToxG9bcB8R968tynHOrVHMcIG5Rg
4u6IhWfTudHDProfb+uafQipHTzR9YQlb5k0LHkZEOnvSmg2gEBSRQpk1xyP6HpM
d1kI31OuzsDgfeNFq18MxM0nk6NFI5fHT7ycKoXHq6rkekxw1tt31a3I4Ea+4RGH
cbKPeIpzHVFUNLdrTeNbLDhkkRQu8/MtVoGQNxRbHUpXEFVTCktW6wSnG3BNtH6E
Z7g5dbZ09Rgu42ZT7hESgF/aLVPUjc5F9f+LK3Ar1jxGAFlBkH4QYojamg0w1kNb
tO+QmlXRtJDYWkZ/E46C0JMFYmepgOH10tGrZn6w+zKrfTVPip/VnANSD/ZCYgi/
FJe4aPT3pwHcGMm+/V6Tx7Ebc3cjCv31mAue2VkIY2ocrwiUKIrRuvNcv7tUcVbj
jQYx2la6GcVotNj9J95Gd2gRxdfaTSddC2HwuBHwIl6x6QWhCbYp+gXMc1E6WlB1
8jLKqjhKEtqk5ERP6Ak15y/0IU3yRMj4Bdm6k8iOA1CS0KX4xwdbIKe9Nm5PTLaR
zJJZcDAdeUL+PTTLb/hcmXmm1aWz0mrrYEtaHXEmvTkSRHtEjo1PbgEFhHyW2a4V
4a17CwdOm6hU6wRtKGf/8kTd/LVPlxNP+OWPLvnOtB3ZHRMMLpikN2mx+Om6b0y9
9G92fZ80PvemT0W7/CAGlAvKmvixB2RBmbSrJJTWbX3zL2uIVyd4St8fyPnGVmAM
pNOYkWkTil1/9F1G6aHEXtVPdqmIL7SL77dPNgEy/r5Fg7Eh6L7qjf7EcjFxFza+
bWSv0sV7vx88ljI7LKom3btS2sNaTxqtbMv5Y3c34jIVoUaoGdajxOAZTusQCu5w
2nGL9PNgq2t+Du6S9EnujnlHSoCtc/AJ/4bu6lM5eCE3CpO3ApbJRtneOKjaUjtV
2ENTAoPVe4keUZgFUItn6ZoDYl+SAZSFz3TO4vRYKbnqYzTfRnbrGFH5IKw/oODE
pgVeYXt/pnIc8bsgOFW+J+0qdJ2awIIaubE2zkxFaDSDRqa8PEF2+3YEto0egtKs
L3V/etp1DNr8Xm7uP6yYsA9nybjVg4famJuY2eXe0s0B2D9y3a1hgHVdpBe9Ymq/
wQXlz/nz5zddYM9EF2TNLuHjXvd+tCAoYKQX21uCtMdQsnnZe/B7QlH/5hzFiVtC
iveYKy82uIZ83VqgIEgQXyfQzulS7Dy9OOuzzaX1YtV5rYbMbC43P0gpn3n4bBRz
JxNDdSxijtUP04C+S41+e4avFxWq6bcuZbgo0iMsU4kQu12C0yr6DhsL6L5CUfJ7
qe02D1G8z0TFAceTlKuqu+AvqShyCU2H8WG/iDJHWpVIggPCzm/oZ6EvLkQ6XhEI
1wNxfrNRFi3sQRryBtQ9yeBRc7PfSmVvxQQZJrpBT896e4noN1AS9iUPLt+21XfE
D6dlHh+rcJzFT4IUdzkuNVD65IQIkufwzxjgqsE0gdJVZW2xa/cGWFnHKgs4QcGy
weMnkppy+YlK/RcJ6dRH0lRcECqREp7VB9wJsY5QTGMTzde9J2SsQnO3AiUxlnO2
p22G8/yCEaPzYfbkSEJNB9WX+y4T8pWTf1xEKrR7AOo+99KI2YiQTMyrsGSG3VMH
mXYtHCsI5UgiOjsIEmQtS7icUcvT4uHmyOD0clQCdgVs3JKGhrctMj2cz/PWA9NO
OQXV6MHsg6ZIc71E7ij2U3CXnhxGAzzglxl08y8ZlEbNfqXSIixDmrMPQHcTy5jX
NQ9vtsfLFytZeGANP4IQigv9GzLFpBwZvRRVssArSosLs9xq7SY2xbKeBNbqe7U3
zxTcwc6QwMDarfd1nHiUBmPsdw5Cl9zRU0nJmi6kTfCjb4VXtt4UdqX9j2AGLApP
+qRvxCa5/iROi9CL6bTanM9PS5tvvce7k0HOcIG75wUEGtqt2PYeOP/Wi0Hce8JF
W2vk6Ni7ivhs/fnkfYDH87zw2FPo3NyqHR+iGyjvwjyltPknAij5oaPCm24HzQ1X
Yksq8GdVFWw/vAQdAne6qn0ozLICAxhxXCU/fpa2WfihYOhwDlqNYfU8oIr31FdI
KhbxDVUHpfokwzBZBXZjHIx13MHv+msLoVHg549+rKEOgKR3UqR08/2Q0ho90I4g
SFsjE50024qJlrbsQMAnnyHy+l0GyJBDk8I6izO16jguKx/gjBDCTwk/XVIBXJZK
EhpBi5o0BiojIRK1E6xCXJkNMjCuawOd9UH18EEs95PBYZLfFC/0a/wMqo/3F2zo
xFz2Lk0q4wF//lWsNZXTdXDW87RmFrD0dUO/lJ4HVB2zGxGAkbmzadBPdTOsHypO
lA/AYiStv9K0LhKY+PfYWpFYpFyMBDpl9jnNDBjVfei961OFIU/1CRPAqucq6ik4
Rg7EU4m9MaghMPW1lN1y7yJn066EsvXM+9v/nm1KGTcE4E+MAJcfosGCHp0YCC4c
uJGDzZhI7rr3egb79lHdW1buX652EbRRkojVaad6zeaISFqPeFYdlbMz26zgM/dc
MSYwu/4myp9DrHgTSVoAYtOAYi99JXMVR6qssL3hTRa9nGZO+iumooH1HRxqMaD9
zR06eRdX0GRf4Rh4XDjc5ZEVC7G56vWjAY6rDDUl+R/fkrk2yEgTEEBg/ko0ZngI
pmK1QnShrPC7b+DuxZN088pUk2HNiQ5wG3ZrW7npIJnlkTIefQRDUs7EaFrvXYNp
3QXQ/X/CwPgJ5r5QkTOSAM04DcTLKK7HpS+vCy9WsYBbk4ZJgePvjvQKPnZpc61T
Ybf67A7dG1AL3x/7u41a4AZOT8i13QtcZ2tdchd5IBc1Oo6mKSOr5Jb3VfLUtpCD
RRlknSx3YDGCg88dTw8gKI/ea6sXJSN9hOap+PfQ/1ZGMrp3wr7PQp9du/M1zFqd
0e7QHjefnkeLzivzG00G3BjDjwdWHN7sdei32XGgecn4neH+FXVHslXqLgYxYRQg
4x4aH3w2Q0oU9+F9joiLQexUkC3dDLMTagaUSQFo2c3z768/M4K/5IW0/AB/tznW
wnnFv47+aoozMyneZ2PMj6CjiCzzyAQ6Uh5GmDFBXdPsjuhIGoXm7ajHmIn1R9GV
VkNmMkvRQck4fn8yYd7SbnnI2JWJcdwL9RO1ggm7dffn8Z2+PjVQvLCu1V38yiWO
RPTeZklV+Auh5T35/w8DwnYhKaGfjXIDqswC8NTOPGM1y5870ZppZU72G86uWfMP
SgZnhWbShI3w+0N+BSIWa0K9+daLzjdoXN1kNXbtN08iyUIcMEyVewcEq8qP9ebm
XaGj+vLntPLXN++SGSaYwZ79gB311C4xR49saeYv4OzO6uKfoeP7bqFWVNfhhmv4
MEBSS7HeqwRoN3MqD2XJDXHz9X7K5hGznNQDwFUlePkqH0LVflAwO+kqica0snfT
H3KjmlV3dVc/cX5qtk51w5L41tT4lZICJHvqDd37LLHNPru1dxwEg/IWfqMbX9j2
obcvr6FyFJHfIYkCNUJcHcb2QvXSYXwKwYAKnXUYbZjH4/El/t2qnywTm2C2b1OK
2XhK7VzrLjW84aV5FmGVuum+hN+3QTuymiaNXYJJMLNQGRLPXhnTgONVBX9nVweJ
2EArMCvlaq5fnpWNSfoNsK8z5seAcz3ZMMpJQSGyhk6skhQfLbrtordATAG3oBVk
KKoVByeCYWkmJESoMPHtlCO3wbYari9zmdoUWU0BjrpmsBEI7f9Ql7uPAs0x6jFj
QMomXXJMRBVA2Ja20acNdlZsfIy8QZVmIwprtAc1kitqQ5Jyn9IIFCqLhwTEY5TO
vbqE1xhIf46AKzM/6ZU3DZ/+eu8R3otN1B1uj3gssKSVkwOzvUJShwQKv+qf/wJz
Z2zJcibotuzSQOH4+b3RAFPpS3HYpMh2IdmolKtz8nypl8ttbVqOEuJmhkTY2yk9
ec+ekZ1VilH1a5w38av84QBgaR05YpBPO+Crdf5y9eRgpM54oi5dCyFbOYDeS6ph
srcGDU5OqUH0P7OueL1rEaXAGPiM+7RCjxvpMUQaqLTpsM9RwXcUollwqsLG6u+U
aYDmRE6I8NEUo59Ez15oSfmgm7bmPbXGjFkcc9toc4uEp9lEVN2lC3DFwp2/Lz03
4SdlmsjUnsdFo4AiRjRPyp0xlWLdYfJtCjw88rcWIIuFoFSPQTdv+ZTyH/ENf0bX
hu/yWW4lShVkbikTBMqCrwPTkC/OW9lbTx8idyD1qXPIf2ckisEZbk0VX54TkLx+
kkWNTZVpSDi9JwRY3ZqYPAhEeHPfvRqxHJ563SbL3fPQeDKvmH30QLEkG8FQ6OZl
sxsRX4eAZ8aQQ0A2XMnwRgkP4DrwmAWvrOY2zZ4NEVjHeJlFNy2VlPmaWXA5PCv7
E4T3qyEu1LiAM6ztWaE2TR+fkGdwicNOqrruxqxXiESoX59VNa4pM940A/Sa7FWI
PiNUA8Eu9Vdr5xRHcOlqbrZOYtZ7MSqM4dVZwC2a7U5vb+deB6W11sqWQWmmztvb
Br9qCOKAT2obq2xa4rUqjbd3+F0NsdiDlC4vyRvzC6POdCoJFaNZVt/kQpcwfHL0
Sp48HxPRMl1nneSMn254aAoBmt8iPnqLoH5g89AeWmauO0b0o4RY6gT8kBB5rdZU
fgTUlUC+Lw9hyeRzZEAmRKZJ7EbmguVbSp5kFMmuM+Vud2ZCmh+M+r7/CDOPMyBp
6QKOlGnMpeJ6fwQvsBUZWJpARqO1c2eJ1DgAUYswQeJWrxoRTaSRANqBjJnFfvml
M0yWeDwBVpt/tUGG4JhOFJGOOGs0Mejq8DCQtJyTLDGwWMSzoDOMB1fz0LSgjbpi
+ODtw3AtUCog4+kYN/fpyCvDUwQ4vKhuNY5RI6qDb1ziJD5/eyIePg4Rd+LBA7my
LVZDmIEKBV4+8pqtJUdKl3X6WJ3wBHGvIt1Nxzze+z4u6Ejowk1sjoMjDPXx93aj
lOP8gmoZNt1qg5+UaBfsQ8wvSJ53WwBs5aASZKUGMSwm0S0eqo5TlcAXrTlB72zA
IJj96lS9CIgHbxAZtOWIZl2htwLp+vjGugF/105+7v6FinY3gLJdN0HrQZgNjOBD
XR3DUPkyyFIEwiBCoOyc95tssXgf3eJY0+toSYRTnb2CMnIqIHrnxvx0H1TU6waq
AO06pjz9N3ZfkzWyjB3U/4PBk2gDk/ZyPazz5lj3rBp2coAVekV5xh59fZKhOyW5
3XBMy/Zdymz0MmCJIfsFAI2zegh3R4w+LEX7F0OmiqQgf3Q+EJXmew/S4/KZKfIc
G9zPBZKlqzOHTFVuK4lKaQRTF7wd590oSQMIGlj3vvXJq3VcKMufCIRhUFFoBQif
HkrX6d2U+11wJ1xmdxMaHXBgNnzxCbfYmG4vLsnEcFU6bW5F5ePPJZKPZZXd0S9f
qQBxaUjkJV/WjkGQHhFUUkbke3OA2ZGF88YlVA5+mV5ChifIPgLpjLQCbbXMRw64
g3giAIuksKyBVVKR/bR5zhDPSlgjFDNzUuald4PhgLNuFugciF120D6brajWCBkc
Ud4cP/Vr3pcTDTieyJ9yD4OClxd5uZKI/qL3ME6Eqtu/AI65F4WA80Hdzyd9YMfr
CyAAIyE6Qp/aOFW9yRf2aPpnGyfRAtQtKcr9h7JiT/BSKzVKadEpcLuHpzuWIHZ+
ku5XBRDAcf0BCSddou0yYZUET8Yu5wIffHXTKNujghxsqwDpJcfkAymbg8+HQtEi
m5iBENTKx8wpfrHf7qS8ZV9So3CnEwHIvH/7goTkSbeT4HYVV28+fMXqcd27S5u7
HtbqzbsGkr7uCnxGcbfsljGs4/ow9XXKVjenbFwk9A6BRuWBEQbZwuusp8vggx28
zJDq7O976MBnzfai4bs4MANn+nIN3/UoCnxWqos2WHbX1uwxDmNcLiTSvLgUc7pc
CCHIUNelP/0MYv0ovJ3d4nZ5jW6vtermX8QJEHcIj/l3vwtknl6LV8w/1gyS6VvA
cDw5f4J9UAig2fF+rtFN0LU8mqpN6ZkcJhGgaK2Deco+abNK676oMcY+8dk5tH2Q
uQb6AUIg1nXnD1kit5uI8YULSrJ8w8AG7RCI8Wj5b7LKUQWBDFNdRnKhpp594n+y
VAwo1qXKoX0pgzvY6MCgsuviyr+D2z+C8zg7hO/A1BqS73qUQvLGjD92fMvz+P3Z
Pry5dD97HS1M/V4N/U14N9SQ0UMi+m6Uf8x/eZAHz1Ki1W7FKWckXjmeFwUscUsM
dZvVel+2tKsgNDJrKlqFiJxsBPM7H7QeLTJqmErabZNmV223uoJFFccKOhIrSPMQ
cq2ZP3sBf46/baeTwPUqr1LJ1R6ubnAeMGnDg1WkMhjrTZrWr5oQthwVQKBFIdy2
CEZSFwxPvTCf1LDutBH6nfiQpUAyFNtfc6TpYfOoomcD7kcB3UVxf2fhrELqceE8
wyEPJQU5COcNDMYN1w1OJW0Xc0gxLn1VKuulkepeS7RTB9dQ86+dVFjmMj2E4EiO
Qkef1dmC/LIdFklF+rc3N3N90/MyOPLqzvWkPcnHMpDqOtzTqU9HGVS9ydOBsWC6
jGbeYtRHegHNlcyCC2Sh5TASSqpcq7igZgnDUSCex2jqWyUQSkAQR3eGBt4ZKyG2
9S2QB69TuSw4ytQE6wL9LzXmRnJ1ltAzGfHg+At84MevL4+IB/8M5LXPmqOgX/Ha
v22idBV4U3XndQBp6ndWyrBvwmW7dr0Altf1uNGRn2CqF1bVNkPQYNa0+1+jVrBR
fJteyqBAgiBEm+AppFc2liv9g1i6GfAF8OIH0ld5iJzCWCwKaWJhNB+R23orfSmh
FfIsPmDsQFNkZpT0Y0WPOccZhu5czXRM35puwj7KXrfUdG2F1TQFeEXtsbXGFeWe
qIl722iJz/saGEAHPieICFFRZaAv3MgdvZc1b7/iUsVPINDuCJA4FsKdOHXH01I6
e5oMLxaRGnydOwqglFz9XjmIlDbzY+eR5+pbphI/ESHrW4RPfdcWXyTVXnpRI29H
//EN1cQpCt14XQOVcQj6vB4E/+rubV0wfrdSg06M3yqee6MuL6vWaCAouyzuKpwy
gnysw0DOt0DSWuVoqXnjczoO13HRkFqFkAoMB/zbiVGWWJz2cnZnUbmIC7LDqZeM
uT/QAsCBwVq/Pjafj3dQL3ErgIeuaEEp0ucrHPkbOloNgOCzq0zRqBZDIsh4kSqw
ImrX3wrP0TavAeVVCvKy3BcXMPwIpCv44IwabynWVBs3jNim8Gfc2LDXARvFfjo5
CGNPZ0u5LuG1QFyld7e7SB5DdQMHdQ+lUyCAbyFW+mR9lKpZgpf1ybU0lolmvadG
DzJke0lPGxZIIn8tTr0fzRLAX3NxyJgTVvFfso+2SE3n1WBkDqnY54xnkoHGRv7e
UFaxo+Gbe/Yx6hvjwc4ZrqKaHH/GB7du3pA4jVRjP7yQqeAdKxl9U2YMZEgm/oXn
D/H4bD71xPqAkwYXLwZplA5a/WQh5cF0M0qG9EFOqbJEJhGpJL9GUIO0+3c2A/ap
tg6NoDW7nISeGQBoBAYsayVcF4+NARdaA6F/ElWFjIjjBpH7nwxnOdAsyHZQzrI1
Efpt8rPW8lIBuHxLMZQo9INs9MB1V7vYcTu1Sv/NIM/5P5AJhnxhXzGL69S0Juhn
uNSUhYZBgpqWOy4v5fQL739RHMIlzB2OtlIJTvR/VB8BqENm0VW/BGXm4Q00Y34J
oLQVLTDnKiqMGF+VdG6ylVMzY1XFMXuRhYiOhR+XWSNpaYWRkDrK8uwpumM8agys
IDFLAZE7EVaWsOnNAw1wwzgO26DNYK7enJQA7d0v7b9q+iTKEV5STlJ2nIWKKagh
rEWxP4WZFX2LEwpwXSmrQk7BUb14KrWiRbk6kpfO5HSPPasedbXk6Zx2lFsETaA6
jm0PaCTopYcgk9D74JnSCwLhYTBdKX1KWCY0at1F54vy0wxDvP1HGfWEUN0qbGcn
n4xpX0/WIRGcZig1Nkjb/CHeK1fQ74jBV5BenSOjsP8GMo89hmD6EPhEVOD/bZQr
1ThBOofFpgMFDnnKGcEw9U1hS2j0V94GIOsIAdSAWt4igJlRYFnTJqkJaK0dzAUU
1twcT5MS4hhjLgwT4ejMXBzIqGDP5Ez8PMLYvihQtNgERFvNh8fZ9lys1uKVC5wM
t8aCocIxO7T8oSl9kUKqfX7YH2Op414Oak6n/iGyhyDCjzY6j0tDKgFUL3wruuN0
ovU9G4SjaXzqWjRNWpNBDZz4EuXKgiufxTs8tzH+KXCHjOqOXHBVCQrINbKLFA8p
qwmI68PS//vQIE8JOMPOep5Kn90TI7INhkGLQMRbY0F5pcFF0mXQy8Jj+wQL5+P6
61Jo0piUpTY0Cju+UCOcTpMQlloXbg98YA8RbMl7PVhUpou8L56tCaO03yAmEbEK
ygKuixWB+pfhDkNUQO6S+WzUzNKuNoEbHpeLCpTPXEJ1rPKdJAvSTff7zT66qHhu
WKSRweRrEJe/dJTDNly7Xb8kmVyMcY74o/Mo6UJtE4FRgzZsAMx4Zj/YhrJOliFy
5TVMrS6CgnVtf0yCQZ+F6gfgkSFtIED0Kollm5rFhP6PDWkPv+N/V/qlN06i6eB7
EfSBbqT9jaTO5RfqREwpXcebVGxUZox81bg9VmJ2NssDcQUov52Rui339VC4+KBU
7rBqsHvYs88FtQjDw40E/iTCykrs9AZRPDjwijqIT+hnQYXBINdguYw/iU5J+YTo
7pPNMagvRan67OnbwlIhsRb+hg4daP+hUs7i4wgFzYYLT9V16eaiJ/p3wldKPm7n
XJhZodCQHLWbaJ76BQFRPIPOIXnILcbfwK8UmzGXeWx5+p2G0NGISiYCRJYOKeNx
PsJPd4rfr4hFFjxWd3rQ1DxVlvWBXRSTrdv2BWvkWXiutND0CZlfaJOSPMC7mhtk
XAFBFotT67hQA+iqed4YUX6lrHK8GP76TttPMbSvOtHjlMncqnHQvJnpfr6BgzYI
+Fm/XlC0nytwoIPXpNjwJaKTmsfljGe1S+O/F6NfRkgU5dU6T0cwFkrp83F6Y0LC
5Swa9E7YFOt4vBxGwdUlCXk75afJnZipx25Ty59FknxJ/ZKKxnQZe1Kfaapk41eQ
ZDYOSZDyk23O0fWemRTKmDFuNWsYVp5RBcUk0DXMDU6hAWlZSNZbV7AQOBrDFgBI
uDGLsHoc4TZQuMdj/y+W4XJf0Kmp9JImknAhrAGg1siV630nh2Vqs43wDOCTWL74
PjXAeXv4uXWzemT7KnqdKb/OJ+04RNJc/eyh9kFbhmQrL+TJfF4bv42Y71h6aGEa
JA4qJNpok3bEBMd734mcaOaiGWne5N8tKSp2WMPh057c50sBYu1zl+UBjumKYcE2
XZSR9Aq8sYpZ6pIR1T27R/FdkBl06JcgVZfZu7mrsEwHvf0qN+jckcxc4oavxtcP
RrCi8ekdYHg8GTslhhPSZmEsShAaowj/M/SzA11gXeo8j6jUFlwjx6CdAAA3fUcP
KQfXyBtydJNDv3U6tTrCi1kP0SP/GWjiCAsuAGD9F/mpbfXlEE7BTzyV43VG+B78
m2NBxVKQDMKrEiuHcskG5uzOxtYilhJQFEuQ/sn20v+eoGkBy62tnQQXdbbAjzGi
ApXkgD9iCNnRE01Eyy4tKhG1D+f9aeWnLjIrhuH68QWDDX51VBmIVx0jBi1uS2qe
+9y2lEm77YVWMLsxTe8J1eTc0IjC9txjcmHYkPRyrqqTvguZEuja7hgTEsLFMqwz
cHKxWHIgGwd6uSpKoBXqAi/k85BAEZfwdw6O3spEQF0H/9v2wi2uhDwuqJc3QbK6
YZlyq1l3JqDpo8BIcLQIRk2+ihKyvyVf9PYFv15Fki4cLNLmBzYzWx4hUAoo53YV
NbuLFZoX79ogkKLfHKRS4d7YmYHveCSBQWqg6X5TCOJjSVSxZwaDMJ29mKi7KwZi
5pcVrjxAmUNjGc0dedGEfNvvEfwvXXAvjH6GXGFoSIBHY+iXPwk/Oek/29oFJMLZ
XoKHiKRQT/fK03jNw6WVam3fH2UtoFxcWkfn5/gMACJu8+QO2eofL3DUzxdB8H9M
v9CWzqAI86VqPYHH+Bxahxt1+7lLVfoU76OmAjwzA/f99u/zppwMKOY9084T006g
Vx3sJDFMtfCGOwK+KQonlHLNcKtRHH+IqktLh5y193gVgoAfUm6zpiTdMmD3InQz
iYMGIBJasrmw1dlGJlFxVpOfoATXLTCrQH6GZtpTYqkm+teqXti/6dpLtg98oXqw
9PNSG5zVrIAShpMP0KbxmFWHmcx3c9+V3KhBee2yQJRr571pB9CDnRb7LbYr95ht
eyoEwF3YcyqspN0qHoOO8FQtFsvzJcngi2XVY9NNZ522mYiZEoQzkwO1QjEnLWL+
gsBYb6Q0CF+loJUUaSG/CTn9Xgj82SFt4xtvhK7W0UHuV8prScXoqjQyXtGh9ywR
vp8RnhFmpzyxqkt8uVsOOTlGNTtHtZanI+UsqmCaQCJWHiWiL51r+HO/+DxjVKGy
19SWX2XDINikUdqdvfIrSIaYj/+x55ThOtyZPwah1FU1PFk36OokvMemUc4oXjs1
Fe56hbH1ML8NnLaFYd28qcZosEclaa34RDYwAAkrcxN9eOsv6NgCmBhRNyVXb97W
mdggRtZD4IyCGk7BUvmBmAnkjXxJNAgMPcdkUb5gdV+OMKORj1xPSf8FvYwYOoQn
WlcQJoPvjg8+qU2qxkuppVtHF4Rw+OLHw+kwTZSOvEL8hKorPEbqgghHKJVrSV0S
xTrVc9q93f/nURfWdh9pia6szuezEaluWJEMR44EQbZEPaOvZsG9YdT/a/eqQKD8
VYH2YT6dZBgtD0vf/9r004KUfxpaOiLge1S3p46vfBXsUcvsxQppPoWhTwEzJ5Tl
9rc0B+Wu0qG5KHshB8B5YZBg++WkxbcdLxZQcsoBNRjXOEW/MdvkdWy9tvbFjbyH
AbgzHdq0DPr44iJ8zTg0T6ggFeownSheeoWxhLyY0/Ia6JF7w67UkV1/OLYLChhO
BVSAlKW1BPMLHaq2AK63DaUPYaQc2zIXZqVOGZf9p4lcQikDgw220NQ5H1djSrbL
qML/55y1y94kHJ1bZPuoXNg0YRRpEtsks1GwFdQPIWVBg/lzEC/8Zs3Ile9XL6Qj
P4jT44zUIrV1gInMFZ0TqVhS4IQYWj5RjjahOaJ8hWqR4QsLNynFmEplAy75+GOy
gsKspYO3Cs3YcaCT14EU+eskkOaF6KkQdX099Kkgb7VSLZ1KwBd0+a0ALmVctroV
yrm8/jnFrTbe+TxT5CZhpAyhqe7rwGAhYnkJ6zCgV424Oz/4E2mciZVsEckfpaGQ
nDL6EM2Dh476rxl0s3v6BWPfrcLPbfJDreJsrUa4o17nKblVX1sB0+3kJU/CHpc/
FZSHgq/xG9tDsgmcnG/gy1KiPTU6ZhmEWn4GrdE20jLMlNqP3z4mEUfzF9I6PDlL
qLxI456JPJLw8mOGzsGW9sj1WHIp3u3ild9gLvzzcqTT/z6oa6tBI/efDjLJYtyP
7E/09EMJ1Nfy6v2gP872Nl3PzUrn66UeAl2B8UTOBkFdhnw3tk5utk8awV7NNFmc
vFT67ZfQJzJrCeHQlHOQmMWN/asWsZhSJDSsaSD4nklgcFca1uiQjG/9pJczka07
RzJohvMZ2xwcIFM0nuU8QaNvtmeimZsAXH8o22Ky+/CPKJv8r7AtXL2Q2kdWZbOG
JWAy0TvAS6WIm8ArEG6a32qbo3xXCDDgxr1dqJyBCYLfGTIBpBDWMi3O3zpdAjlE
aul5xdRQuaPM4ZwY0gt6yj/FZhrN7QROzSMAuwcv8l20BEmJQucbUgn8T9ik94fQ
zQkX6/1JaxGA+dOkeDK5dXjjPGR+lX4+p1twPrfzwd34cL9ytUNMvRCu/pBoEU98
erVXyblj6wSWpUJJCuxqUXDUvzq20vGV7huI/viNF4fYzmxcA/EIXnyq76UBaRlH
7wh/rMKX4VhYa0/G7ieeYk1jpSzVNvRR4zXp4SjchwsPWrsscVEyY0hEk+LmSe5P
HKqF6rwF4dcplgKCwF4X9d8cB3qasJ2PbvEX3Sv7KZ+PKFem0R/tjF415aQJKkF5
igDp7q1ZDeLDUl+VBN9e59sk8URjAk668jA2l3tCtzMl8wsn+Gpo3GGfoGlbQW7Q
AB/v3K8DahRYcAWIPiiz9DZc+2pKOLFgTtSoib1tiLdj19qtY7OmOfsQM/INuf+f
XI+cApRghcFVfyQOY94UtIlGS2yasHe7ioNn2iTZFajNNa1LbF6Uyz6Ksg+TJoUL
EZ43lCj1WWynAx8nH73ckSXvHB/Liq/oryzlQdbwTtoHNo3Y33xMx4v6nI2eIwml
fT+d31LWHYw7w67Lxn+hwt3uC8wvn3emQBvzYkV6xVI7jVgs07nDi3D+3MJJeHWC
IOmwZATu4zVbO9T2YeHLsPEYAvhB6O6FEV5o5VJPd+IouPXIHD3O7l2m6z6gYkVs
gqcAJWT+wdgyZPZN5OUJhrhXS1pNgL4OuRtze94RRyAODSFfcppceK9fqLyKagTm
XNZned/MEKFlkYiGv6i4Ev5ERlbkFeIzJu+A8ubQZdqvwmdVenu+NQTHqn/wbHjr
0CPild1elbffXRyCl4jZwsBlG0rD+wSCZ13LOzk7GuyaFWlsc9xnEVtLiJNOyxeE
Nd9efHHwEm+gW5wz4HHCGKekEtU7/tgNg5TFlosbDuP7FFKxjQv95LuQyGJSNpGK
QpXkw3iO0Z6c3v9hhamfuW5x7aP7HqFz0yZL9o3TJOJrrv2pvpCe0BZVhrvsHyAp
QZVzfmj4wlAYux6zCf3PD7P3lX5oSIPPL2NYKWGM/TyW6h2UolwY3+brt+jKmV79
jhHr/MXKwxCR3XP0ZuwBumSiMWtZmeio6XxAMkVwWRguMmbtqYpHBvkMPx1wdBc+
o6ddcwSlZHpdMcA3OSzSvnj+VOXAwpaeoBV/dSnqSNrIj6xKXX+D9+k6gzd6Lh8u
G6HGFcmBktHFgwAra3s/nLV2RDYMOilThXQkiyS2/Q8kgAPdCFVI2OINsgRm6bCb
2RFHqjO61O+f3oTFtWVVt+2BGF8TwryzHu+UzgW2evMIYxzEA/jpKI6CebZ1qHmf
uD8RywYryZhe5qt2EIuL+4WWJ7HJIqXmNhMh96jwcDtnJ+7StAzKD8XaklWyppie
imy0V/J+1JWC+P0jCjb5ELG4j6xryc3HOgFEVbeBikPvqR8uPF4cDQCsGWzOkYOG
nSHdJqlSgh7PXhKzrzqEq3Hi7AJWJECa++xa1oLJ22YCEiPb2X1xiQNaH7fMPDQQ
OpLbq/IS2eXnrFX35iENVdLOR+jV9u1p6wCete96ba6FdjXhw0k/ySsSFLaLdrDw
rQTot+BcLs8k8WX7AZXeeVcOzb5jP7qDGkbtPWlBsfhGjUSZVT11duD26iJivUed
OacCzYN3aYBg26T/K4LjiIU8uISXOznLPxtuZPhdRqSnknI45pouPft2JS9m9fFy
jl6sQsQCguW3MNSMkpP7wv/tZRRxBoA/Exc+nBFPLEy/ZM8UNLVjy1zH/MxMieli
AylfA20nBx9OtOhfUfcrpczqq1ewqvFPexwcLQ4G6RB9hgBbkbdWE3xqfjq/TQxA
1zP+3gsoyruneiWVRPmk/ZnFAbKPVRlJVDNMcS6hJ5w6r+CBxMVrex88jqT4LWzQ
tPBdlUlhT9/eavtsbMNcz1CjBizxYULR0atHE813HxOfbq+Ddt+ARexbyn7z8bhY
EWKuicvaB1YCLCp5cTHJUp2bMHe+QTZSt5uyDEJ90lc2fkLmNDpYxDEaLXI0it53
t7SaZVk4rgKC9VHm6QX4bDs+PDoJvPMcvASi8hV26gxC8fq0O+FUSyDRkmUNILIi
OgczAd60mbc1wNLELQ3Ph8yGuQJvApTowEkEXj1D0+Btbw3fazYH3Kml50OgCEhm
Xe6tgBaq2BGPU+FHiipiNlmSsq2ueR/7DHxo98kH1sFafzZhUZtGT0rG0xeGrMRc
10XxUKn7nDBx2bytMDgA1pPJpsyhcW9TgZX63GAzhiIZrUinBdKpXjt2xghxjBZ5
YzcyuXBn6r3m1z4cNZV0Uv92m1pthDPJPuiDDOlquhDP3qdnWTIXnkD1cNd5dngv
9S4ZYC5HmiL6j8jDqssvNHQUwClDUCzBNVxGkbjzMbgDOpxdqiKqc4IH3PJ02iSr
v9q5OtOyEjzcYzmFJK8phMJLdI+yIGvqpLO4NCNCw92/H+G6qegbS7CtV6Xffvxg
P2VHq7+MaBp6NoczuO5DZ/fqIejPxNKR8fK9qo+Bmmlml/rQlgEcaxJ+PsXgZ1mk
wo2EjyVcsnGjAkCIq68/1QgFzhMHrE99nM9Z3PflmIt3yN4qf+DyOCiCRo/JSOVB
Ce+RU/fpZZgAbGq4/S2xH4ZixG0DBH6B1HpgHtFD5B4hQeWr/V2HDiMqKGiqDPgL
1p1SQpGqNrfDGudLQo6KXekdmNnw82CHZvauvsNmEM2Vw4ENBIO/kL+1Ru/ocCSk
F+3gQDv7OC3RcrQU/m3OxEu6avQ+rkLN3MraZ6MOkiX54C+e6rPNeErxvZaOGrFs
7UsvsOg+YylyfNJ4dczu5szYvFWGMLvCzng+GHauXCDjGJ6ZR6upXKF/PMibY14J
gUCNa3khwh7F2f7BBd/r022eMLV4HwNIg5+8FOZieCiWmVE2ezuHkyjcR6Ob/1pc
0hMnhfXDfGZp9GNEU1/+MhfcyAabRn5NksMH2WR5vgI6MztuepvIUZXV1nJsiyAi
jhhowfQzMFPHuvnlVOEsAn+16jaWNqSMFwtAsfiMAc/ZykwcsRoWw824NTC4Gp2/
eUIE6oU7IHWiKwU9bt/S9WQrBs61BlAjB63htYjss/g0iunrEJJehmUlwdD6adGd
QDQ1lvtpKSW3igtfF3oH0bhmpSt1opxHVsoMm+umh9cIugGuI62Jvg7zNmHBdXVP
r6oB8x6AlwiSpBpmTN+K9bLj9JXDOJnrnR6vpZjtvF7VBAQ8R9uYDtaUjq6NQ+Pl
vo+ndEIWEQ6ir4FGUbm7r4rSmZBVGwecw5rCe03J5TFLkF65f2/m3O7J6ht3nJ2d
UowFeZSK/tfoevhDduKYij4Y5XuMOtsepUC9f88lFvJ9sGSNBLzGGuD7utU8lITA
RG9EfqmzqDlyl6JhXKzJ7QrpJw06XPgHSZ72sWUX1jVJCIXFeBp8nkBRJtgX4dLl
8vgEOwRa74WCfp8RoYM9KUk4rSDfUwZj7DfUjx2TxjpMFwhmn6j2oLwIoCMbpDSC
8CAaOINCSU/JBZbHxhK41UIx2mVxf9Cs3B0jPVqJJi6fjv94iRJkfV67HVBf5nCO
iSXaE5Y+fxrsJrxSLddIRJnHzUG/MJLA+1qTRkMeWjF5bMMfuLDCNyt07QB5FEbU
crJ9R3cSUpa6W5Bj4fq5Hg/v3oe/jgV4wvIvbQwAOpCZLKEZill84Ll2w0zS+ZL+
aEVnVWZjO0LzlvzoAuXPOtRdjphekSvoGZAxJJA+FMsL8azHJUNMnnINz4XWXiFP
ZCnZpB0YiqBGaXpkyfkQpenIE+D4opV1vmafM+u7DqUA5AyRo/cEBaKpaS/6PR4C
VWARlM1KynJpE+X0vxGrqggEvFhzf/ic8REkY0ePOtrZtg1UgqXfn9jfA8IYrAKQ
d8omID2jIa7tOIDdQaDY40SRsLlv2ZwAYKiXEMDaol76SQiu+z9uG7+YlDhAU/NY
vzXZDp1wvhhAXyolvDd+mWSwC5flKDVggMqhF8a5t1MyD2NpEfH8OCT6NjoanyE6
yBPdclU0OmsB4YDmZacTg+pkRbxEOep2SwSWGsy/ve8oS6KHFZ9uJcHwQZyRp1+w
HLW/tjm53donDyJEIpWmFscn8vTW2Qyyo9t8txTgBKIYKeniG94OjMLk1LhVGH5y
eKVgfUnj1Mp0TSkjPpvKzgq0jlB9stE2jxbtJunfkCfqukriCfsyDGZj0eQ2TFCt
UhbjqE7vYOUlHVUHcqg/SdtYGZlFa1JM6zVj9Zh2zQ39EmMjuFqI6/a8IaI642Qe
NhuSQ42hv+sGiFA2wwl7mL37lWsaFcQcipFAubjGJeWEl+C99BJb+GJREv0cmKv/
QtZtd0kaVr8ogc6n/22bc4Wbf3vfiJo0p8Vdu0k5+f+pbWXPNgK2dL4yv5YFA+x4
jzFZqDUc1UCOEdM6zCH3ddvueJl7keuAQ1XWsxHz8wCJ9Jgqe1vEwGBama2CGkci
Ax3nfMGh7db0/lXG5hROspHVCl8lTlmFbJ9EPykNX7klIy27FmMbAjEuUfRBxhja
3J/UlyhvcAk5r47yQgO8HTLOmcPALf/S5FLMW3sBRUEslSkp/djnosWb78vLDnyb
8XACwAlGfoHmFU5Ss71rpq379sQ4HtJxFREvMm8gJ612tY4hSZJuy9A9dvK0Nadd
JESFu24QmG5IS4lCog/Zw/+BNxjJcaRaOPbG7IA58T6yMcE64YDSnppHqk0g7et5
e2li+7NdcD0/VQLmV+PUqpkE/gNWA50LEItySYUoVBcI5KMStazrU18kn45b3NQ6
zYJb6R2C5eHdkwYYQsteMpxQLLZW6b/+lE9ulLC5WlWNr7VWEzhF+9QLKvNGPy8F
oF0J9USzskTyoFFvAhUtQsHmnYukjc8UPIhI8ccU0VGX22TAlYrsL2gXFFh4vf5L
SnnGffx++ZVi1lS+aGPwrPiQ9wP+dS4ziqE4rZFZz4LeQRIQrFIkb7Aj9jXrdmIH
9Uj/DlQ69LEtjntnwuOlqfkH0IEphV3X547RphgYjuJPeR8HqD4xp66fwkbWagrg
WNKw9NRMijJtTx0KTDVTA7OJrubbabATMmIVINvA4pxq5208jTv6E5Larh43AaMC
nsj0PGfh0hRcWcLx+WHYYdXss/fNVPuePsH+HHzGwMLqTWEIW99hWcCXMBgiTqKP
a0haYngbk5+Bz5JTTKmxoJsLvU9NEn4034bySKtm0Jayf9jOEpjY9Dp+o1k4pOV9
prvYbMjTU58T4338Y0m7naIHOE2DSJplTx6KXO9XZghyH5non+GyckxvqZpOSlpP
GLkPxFV75NdvfeJir4LejCB2wp+rmqLsWfuFvg30Huo4a2K1tAmAexKmZopOdNR+
oPTeNSs/D0oR1xVEPXoCrOcUzBByUjNIciuGzySsGYravTBPlYHpqanHfnVbh04j
D3WXRCxw2vpe0KmavMsgnfkiMO8ZhWPA+RwJ+qqpOgEKcLgtR2zXH2AhFrOV0iZk
k11IuOy3Rf+wkcnNUxfjUv7IwxbKKacAz06xM9rVE26JjfVnAfvUCvdZPpIxKZP3
YWEbl76F/4Xrx/u0CcgcxNUi2gJDhd7bXa5PRzUDj9X5xoH29qXyKJcN/12kDPsh
f6Cy3dn9uv4maJN8JXsg2I1tIvKIFwPM94Gf7WkDtVLtaabw0eHijgo5bi09/FE+
x/C1gu3ePUMH52UEWUFKi65gJcJqYbYWbrlkFZj88bFvoq4bcMsJEztQmNVPL3Zh
SWbOMpXPp3m7OnWjZyzSJC4vsO/8VCif6L6L6bRVjfDeld8kL2W23R4Mg2VeRxRQ
D5vBQNvcSKNPR1mso8KcN4DdK56qKiGn19kK/aUseNz09MSgczsOwbTHNzqR5GW3
bRXTfAmGaOCUXZydlWvIgsVtoUZ815FzXk31MVS4wN1UwQF7FFb76LAQtwGLb5qR
/sNET9mJh4pIcF9mrUBHcXpAUIxTiogbdGiggjGJVI6tnxUZ1RCx0KYEaREwxiF0
qFqzwG6SSHIzsNLOd89nWqDD0xA0Yfcd/yFSWPmLNmD3L3RjxbclGXQzdE/T8gHO
oQMCBCXMDACovdN7424NTj+fRDc/F6IqU6xNuRNoz5Hcfi7mJ+1Y4oOrb5BKagNC
6LHS8g93W7lIZw+9LhuulkPQohlIOm666Ruaa/QJmMj2/G2kgM1xHrQ90Ny5tQ2f
z1TaBnWsfgjb5iDIolOMbeQFKp0kMosu7M+9OMyn3BwFPMPxfdqKHI2a7AJhlxLb
UCYbP5q3CMDAhjtJubJdWtDH4WO+h6yBHndSBfXUo7tcXAC1bN/gpa1JaqOJo94k
iIwbQqT7LTLbCMAvhNqODme3xkz5jUV4UAoBbCKN7Q2xX8kC9UojbgYoall6q3oS
kPnTamO0utqHHl1gQpNUc+/EU5WpeAuXAXqEc6dTwB9PADYJ44S/xSo3Zy3yeuOx
jEcHkmafHBCaMSJlSrl/SgWJXSuJIotAQKjpn6Wnwtb0L4qIVUQC4+QXva8qrGtM
XH9Pc5Xz3frYc7SMHWkiMWQjrlQKIkWE5C8d04EwgaoauCNXmRUNICXluElMBzU4
NoiKxxlyQ6AnkuXRATrXa2KVLis/NiyK+yigvaO9srlMCik2ditFicsx5d2IN9q3
I7ibPcMPaL668YQBAkZj4CkD6yj4pcukMlSSmHTwD5sK7OQGfEHSzuWd2ep1eyzQ
pj17JYatHtPT8VYs7A8pjJ4foF1vGLfG4nVRfCLLnCPBgSQ3sx3+tgJnIEQAJylW
boTFA0bWNZc9/n8BO0sitbCsF5S9nURAvtjf5evJz7c1tALlAnupHLQCQn2gYMPC
tM3hGGMacVoeKd3dB51n8x1y+FqYI4ZfIzXsUCPyWLYgCdMyQtIEOnbabtazXLGR
cl4RdWK/HJdNFF6UZwpzfUiBBxB7wrnd4nB4ZOFDaAJ9z6hm41Gko4FyF/hC4Z+G
qkk5RaMBDrQetiKEtjcz2XxZx5+E6apRG1HYg77jRCD3dkO7KBWLxDjl/D3XlZKi
QjYR5vM8CwS3sElK8pPLb0/apnuTyaeMflnkTT+bvbENdZqcttYlzskdm47OZIB4
1LfQ0bA0W0WXf5dsJY1jTRcVR7zeBBVMcHg2V92Ly0m2eLNZhpojXJjQHLin1pPw
mAkqxhtWRA+kJ50d6YXOdQn59c+7eMDO4RfN1geX9gud0vgozc52M4uMbQ5Zz0PQ
TpdCrR/emqvrStr734YvF9WhJTAQTCJe0uhMAng5dH8GeYmJ4Li6jl9951BP7L4/
raxwz0drPdb/cHPw/LRXORbGcEfGInM84H+s7H4YSWl03SSLYg3j4Svz5Zd15SJD
FfyVWHP1njYfe6dCWIlYySprU1LiOl7/GuWY/s+C3KFe15KmE3d9tX3NCwOkLbEo
6py5JmieckUjU0QiqLFiZziYV7JlkA3HuOrV/nGTTvecxHYeeoBvr5aiVw0fUbRi
O00hswwCaZ6/s+DrYTtkT6qEzl19d8pXSQGXulAa5dxP7PMByoCM1OioyBwl59Se
00ycC9i0WViPHOCutXtHD1ICES/sNjwTdfU+fsjwVGSkwKibQnqf1Rpd0MyFM0U2
h4oFxixI12qrpq4AVYCidiNF/xjSublMeA0atT4B4GJpCOnjm5ZO5K3JTQpw/R+U
8bljw2LmDrqDU1O00Eic4W+uT66bVlnCxLmXM0uV5+Rr8iwTJziA82Ap0cCJBrtH
xDpgwiSsH3fa0U+ORtPu9i3disHP7VP+byDNSHvRjDtkqDFfFk3S8yV06eXYIlwo
gZlH2AZC6N1m+t7nsG0hbDJhY4N8cLiip4LpAp16E4CGeaMe3B0reIuYTv7BKH+L
BpFesnhIl7uW2Zq903fU9G8VRzfBZuSgm7C127wiMHx27yYY8L5egbDKYmnueGQN
e/uOQZOasHJ/n+asL3KBvpFCnyJjG/BLriRaDP9HHjOMUdptHY5wCrGRDxNLJkNn
vaEzvmdqgR9oX5NyK65JBcJjEZ5sPdGHZGYrvmEzJbuPtC1HecRUNJdOVGz9xnZQ
bI39bhfPHS6YupPTDk1ZG/gYJHDBmg2kW2ZJiUEcjVaICwOfYA7pEVluNbQs8RdE
H/jLsTvUIZMyC7SoYjALsjIO5AtrYRKN50Kpon/EX68rtm2VCktjlPJigCLBEUCu
rDmCnM0wlLnqRZLGAVPwEIKlrtK8uOOiXxYiwBzAmqax1920ARftgsHuT7poRrh8
HpiDQ+xt1XdU9/qX7I/CXXoW5daJG/HVQOEWY6mAA3XTdGXq1aW4g6ShGwSiKLIR
0tEnX/C3Xo8bqeMtS7q1mrZquK25zA81oy8zNunEMHeWqhKJURkFhniutZU/uQQw
OdLLONXwwPR2eF0/URGqhs06+8EqqSByS0t+WmQkV/JKe8MGbZbbu91zpkHUWxod
d2EnkDhDGGfVQ3oGo38bYvFgKolcPwny7at9xl6lo2JZxO5qjY8im9mcGYtpjIP1
SWN80JBpxlK3EEnJABMIwI9Vp1bE+BFvgaSg6HwDnnLM2Z+x2+wAMqXJeMnxUnl3
0AxMLL9AZ+VRoe6k1miQ4mQ9s+6gT/bIS7CRCrLlrSlZfnGOM0c2n+Fb1YEaLeLX
LK77TJeEFve5w628kE6tw0Q5nl075Kx6k5XvOeDxhDdFt/8xCqVgQPFtj1oG9lek
LZj5uJ463k1LXtwL9Jp5DMTNE718x65jGuoMGuMmYyYXTJjrXL3lDml5xuYmMxp5
3D30+IyA6VyY+2be4msyedixzeTyQsj3un1T4xo2nWMCT56Yckx/WPqcBTBToJrZ
hcqxGNAJq4ju79SuqaLznIEVEpvAhoeIYe0/cz7v4WrqZS0GphNsFsgWCse0eKH8
pL4Msg0FJ1hqRkaGVNitLfyKE7Yf177mLlLVQ/u7525Gp6Vo6+cws4dsTHxqdpvn
1x79RUWod7+q9eZ5Mvu1NPxpXeWGgOllpJUtlnfvbhn2RrgpwDMNoXIzHnRaxuXF
DstF304XuIO9GSbGs9fCud2y9nEqWmnX0+SB1HcNqZiBATwPfwmEDtZfX8ypMJJl
jGRAsQFfGkesBOmqTBeGFWYrwTxxNjQiwk39JNdvGeARF/fZfLchZe0/o+Iol0C3
Swzqy1DVignHD4kUSTqE+012OtrNXDJLuyc4nevOGiTr4MYzrkF0VMA0iVKvJlXH
RYTbqDnYiBehz2WZZRHpfPqx6Zs2rF27q6Y0OpZZfmD0D9gGJja5ULadkpe1OM06
2KgxpvT8Cu2nxcQO4JeqIzgJ5Znvu+lxpcsXPIgRc8wUfFCXekDHcuK6bXZO+MHq
cB1Lk5ijGunr3p+29YkMjIHuJttHT94Wb+O7Ij7V4IdxABqoVBLviiwLdNVNCn7o
EIcpDyLYH6oXHerc5EYSImllovD8s/zz4xlsxiLYm6PwA6MPibR0KOt74TKU9g7m
HRQEMzBrLf0qkFRU3Po4+76Gb3B+FB/qvsN5lv4PQRhJ4vRZGGZ7PJofzn7M/und
anuRrbBWvU30Lm7NIqXlxnLleFI3LgrGMpPDaTnVwj7K1+ii4Gk0cIC420XBgMbi
zA4jh4qWgfKCaTdadta2lvRZC15t9ght2JR5e5Ijq27tx7HrDWqQr4ysiVgWOZmw
py3OJ3f7lLp5t/m/RF2/9DQl7IjL0qFRBjbIhkPWYgWKW0LJOYU1j4iPcZpcecTf
dcgbS7tted4t7GNTd+wXXsa0ZM8Dzh+Z4idoDBYG0i4GXh4DuBHIzs+keLLhByVd
QJCYnjkE6ohZm5TZIws33VUPPiVAifjBsIP9BJ2C4bJvnJeLLOCXdEuqQajPdIMM
5gf120UzLT+jzH4ot+/t/Qt4zhhOJqFakvqLAEeWabgSuFPacPzADl83bspj633V
LI+sp7XFDeDXDb06VmUmRw949c4nK3zAP8q4/VjNDSR811+vfa7A8IWyi6cSOUur
NrH8xWpmZw4fKsgOQ6SYk6/ir2GJMuyxFgAd2T7kVYLa9S/7+xLQwely93/f5gDs
SBlCsplSoqI8cGdagzdmOl1EFx4brGN7yrMgLHElR7JYtUWxT2bkyvXdODa7c2ko
MTioDkv5s5PKaUv3r1iT/0nwnzpXir2S4wlzqlf6i+UI8ct2FqO7ARp7rQyRHfNc
wnnW5KUYH4maw88ifaTyDheF6EyTTeZdqluGZ9A3MCRG/ZginakdrtVeDeHjpKyQ
886ZM2Mk1Uv1EaZ92+n4UksNwQ9H45cwDB2+nZEDv7cJzcLIMB+8O9ABWF6H8wLW
Ye4abc8oqNf+TJMTezIJuj3a4cjx3eypcbpV9IGam5fT0m1wUS4hXoeIRqrQnrEy
HjKo7DrjO7Mmh7ONsWtviRvQG1QDDZxj5XKrBW57ev2Tg7A0rDkAPUKgcktPKOIf
FoqpF/NKlVvdpRvJYG80k/wRyAFIICFr/KXLFkCIMmm1qQzcIn6F2BgmjwofIkED
WyJFLjWk/ix5Hmlz8X9UxonRnAq+9pdfcEb+PofdkrTL9vEqn8o7w0OKF/bCGfuD
aIZJ7WOdmhNl6lXgxsZ/VZlM9zvYuzNiMP0FO6Vdj5RHStk3x8Zhjz+koOQso2wo
RW6/1h6xnEI5qYHAAlogy7NAQdSFfnMNGHpaBDZK7nQfEB/LUiqXNUcKghFLzfuF
OzVhso9aQAastyEUj8qtR5V2a7p7W30OW2CPbPnpI+pUyyPml44aer8o0oM3VDFB
E2HkzyAMxGv6nRCBqTqw2JtYUqZfdcHHVz1Ji+elMojUAni7VbeTeekJk48jT8f2
znkzljZz1s8crgX4NjyzQGzzv2OD5E5FLkBZtfmfSWMTXA3e+KF6haW+1zg2YOx/
xkkQvLPYOeaPOEzgMSLSbgymBy6KcybjMR53gceFMGW++elBoeXqLu7xMFbmjfE7
ZjmrCfhvAIZxzoJowsfyoQ8cr74xj20blN0iW99GgW4D2VrPhFg7hdt/mkk+d890
JpmSCipgEkt1qdeL/nzoEa5KHyWENQtV/TnQzINULBR9ZXiyZy8gF2O92HfKgBMA
nFGuJw6c88bbgSKE5k6cUGsxhPNyVzOb7XZ16KW7laE68yWUoxOSz7iOxvw6MH51
d6CG+BpWVII0RLUijx1fTJ4hWYP32MvwebOZsL0Z+xhFQQq6mB9NflQkIhZNW9hB
dj+qyivbghsaJpYlrizcVZmdE7XJV5BUNFfNFO4kXLHrNgI4QGEn2vYdGW+dIys+
k9bEAjgDiSp8k1CIx1achImz+XXUMlM5/JbPsEsI+zTAaxp+A3TblfKt9nfJ3A/Q
smmzgOTxRdYGUejqkEtn0VGYhvoG+RBUm2kAj3r65UwjFTb9rx1VKoZSxmlsbSiJ
FMMBNhIZxOgCloTopt8S5s2Nu6ejA3U8arO1hhZ/VOaS+ffR4V6M8OKu592Z7dNG
4X+iN6K++hYjlaOTNaCuXPvY5KFXN4lEGN/JEXWBJNWPlLngz4X1Cp4hz3FZXO28
pc9U4wtQ2oVO390tmQJxudpX1p2TCdPU9+nI3aofa10lEz341PqhUk6B3ogwj6n8
qQZ+4oRIqXrfn6Mv+xT7HTaxCJ2sWn0n3JghIK/YOD4WvCp87fX82UcDwrFtN82r
/m2nO3JjSEpWHde/4QpM6qkc5eGwjDC9gXp0lP2p9iXhSmqou1Ki0/bAfQEFBj1B
LD0jrx1KRPLiwyBv2R9RhnhN5XCVbFCCR0Gc0O7LvILmp7VkNwQnhiG04cdcJG6m
9/mhMSN1Pvx+F17BRMNXw43AEK9vNVQHJscUW7kjYZqnH+Kfcn3VtjJTZPAWqxAk
9+oqD/K+/66rdKv64hA1FyRSexJoH7eJ8h3GSOSWdj8hwmSHzT56I833MQ6dgpeP
wLzH6wUAsN6mbn5rB4AWURXtC3QIt1glF6nyoqb96xwmJ9kGx0U5LGZj3I1hD/l6
mRQthMP1YOO/6Q1yvTs70ehUyFxng7ec2ZBOY1oOb+cMoRXcwpziY0iJPD+osSsB
SFQCEtbH/LSoh2gvWf+knQMKKDta99cadhX5PH6KjnRVnpEjZArug7NgX1jkUl4B
ZYl9QBkeE6X5zFJLwu198yEat9sXOjOhKiU424nd9NoZ21nO6W9t5FRIjrSP7lkN
uI2QtzYNxUo3eOQJeTDZ7uhR4tMEX08SS2ZRZsWxOazXIia9QdRqnbtZ3l3q8/5E
Y5broxlGdTN7f7G4ygxQVxC+dXapxViclwjeGMn1mBgs+hcQeahwpiu9zVoS2Koh
HkTdsicT03zl8TSryJMd5fd7WpvwGayIpTlcMzs4JDAPr5UudC/NqfpCYoV+hhiM
iflfR/zUPNn5RZtQgGYsGsrsg8NUnoUXGbco+jkABaLOxiBv+LKZeJMh5IBb1WZb
72UGA5sng8BrWXtRNiQ4JHVM5896BajVh6QeA/u9s+3GFY/qCE7Uawh7LUWjKm5o
nLqFrjd8heuVE9KPxmlyjrMqLBnHmrK450kLhjzu1u/n8JhrbP56eT6TaWkQWZQQ
r0cobDSbMDhHmtgzEIoqa2D81uxgv9C+plTXaA7p+zLV3v4wl7fVCEwQfX6gq7FO
BhAmfOgA7UI1/HfcJEa9gBc1WrfReO3RrOMyNjnjCxy6b7rktG2rM53Sz0LaGo2n
07/xjynAixMPUBofSh1BnfKS7Py5R/Sa7l2Sq7EWe9MhIGCgCss+Q5TGSrs0IwUZ
dLUtkF2JzlGtUiGumkKJOai878b1UYlUgvsqLAcjf1dch7YN0bUHAsFdHF+yMcXs
oSi1NyBQG1M6jbZG4C33I3y9PnQ5vw5Hj2PmSj/gwbypeZB+yoGyDS/4snJrzP6S
INQ70q/aXsdTifeKAbICGXOKqwqgud6QJzrl7Vcp9XyFo+utq4aHePze2qfvJKOH
E2siV3mCVaT3f09/7SVg1bZlwGA9aA/wXPn8Mo5sn6e8owHxbO7BNM8CNfa+5//k
++eo2AtpJjXWBQMUSXbyEEEjEyLBz0xZH2IA/ZzHJEu28kdSExvzO71U+Wpe0RW2
5s392hUF5dTHf1iwdnCzhvSqZN5sg8fQqYxEG+GV52Y21pL5kQNkH94VpkWPLXSk
J/drOdcuqIVRQwJVtwftJdg+PyJQ0C4qtSnjWEsVlMag86f7BWs53vRjsTJlzKlF
jYwqJkpOVeXuHvTiBVqFTtemx1w1+hqjSmfRGdvLc6l6O9R5SRUNbkyjkDFev1VC
XgUZBQ5aXkBckqszWvKy/rhnZOy8KuDMsP2HYXa6uiuPvK1Y+KKkZ7vJK5ThTP0k
TFT6C96Vd5nLKp0Ktvm0UA2W745VsufTZFEXyC2vLa+eZORV7Ukhev3Ta3bMeocd
k8kvcEDUxO5DqT6yTN3SoTqKQ3PxMSZVpk5pVkosI5C0etaITguJ2TyPuO0uVAo/
ZfIBetqwzLe4g/Rw5Prd2EW61bTs8gbGlFme3pH2T6jMHwNUZqW+ZEF6BSnfTvHi
ZSUK6BnQzrypY/FHCNVtnkbUCcF2Z70O/jzBxtzuYavE8FFrCziqIicXUPvdxZHa
wip76oTtKU9prK0F7QZcVnqkM8vTV02QAdRo/ZRQRZuJ4oG/2hN+nMo0U1W4DExm
QtK9E8C98KjCXyTrHOGPMYiOjqPh1hmRmK8pKr0BjizVviSz8sCy5f19vP1WCJeU
OFH5J6bqwrar+ESuPPBrIn/Z1jDWRyZ3p/vPF7/c9ldI7MxewDtXUouFDlAsBrt2
j4qopuQD4CwVClkOkRqCOuN6q3i9oequMRw1G/9oWy4suLQalHD/vMH+u6LiHSy8
iqyqR8AR9t7PD0NJl6OBN8kY/R7SghjoQMZbfWgn/N9qlbN1J5oHQCW8CDkTf6to
aYuJizjYI1CfIpdkZL0SNjMv5IoT5sRIK/gR7+aDG/E2YCWVE3QQxwSFrXzokxA5
RgLzN/m0zAQlaUPHEU5ukrxhjY/iaRMWHiOJECrAhFcP+XYFPGEn9iZ+z0q8safc
R+mh/BXS8lEe+QYht4QwENfm6lH8+jPVhZgnuiKn7KGC/rXBYnzXj0W7dCO/bGIr
ZfIUCldbteECO9clWRp//kmXjDppYGaOZhdGY7t0n5YxeBOljQlGqP08nd+xcNEH
P2V76Xu2WsR98rMYJMAcQ3kff9jfaGQf2tQTFC05vT6rzztKKzF6Y03fL2C6sdZ/
L3aL1l4HiLTwf38Nxcsom1+s0UHWHybT/nc8fvE/dVWFpTz/UTlVVE9UUNDSQKHf
Lnu2GWLi1cbNgYwCCtMhgZTiRXdjvjbImZgQ9syF2opzhUflJ/7rJ25o2LkgXCzz
qJuPKpb2rQMPQwKwuDN0SRISdljtxQfM+bnhrHJjtTAXWoz4LbjqVh4IT3kuDeAA
siJZ/GSEFDn6W4cFJ/vXFjTtWVJS+kU8whsOuaKxQ31kV+A0pvXeWR49TTeJbq8Q
lF85eFPXjMrW8P6D8bkvvFRvEUaorWAKaqnuE++mmuYTLW6/3nRE2zOFGzby155d
qIdL2ykNfIsmfUQt5CoM6aMhmti1Gqc94lXzFR3PURzmFgrbdBfQQ3XGGB0SGQGz
BUIPgK33cF7FzIK3846vbo+uJg6wcg6G1TtTZ39aMlpjy5/xDQZBgQmjL21xov1m
oggksfGxvzrlNVqQ0LpT1AaLGmKoTb4xqLp1Y9nho5sLD4568qsvCk6b3wA05Apm
8dV3nqWxf1qrZWUc3Hpge+KEe/XBpNv/XxZc3G/B4ML/oAQ4D8UmENyvtu+2k9w0
yqu4oSdjE1+4IPyX7Ll6vgsz4PQwGSNWlNHCS6olcaay9aQG71nRS1SOaC/V1HCR
azcZi19yRnJypIuVLz3qpEFOhtZXB06n1U57lumrwKbqs3gieotsdo9AJuhSHOBc
hFOQLxq1OzJcqZRZIdGoAuzIkUHGvbxNAIWW4aHqXvXLcIr/14nDSNX33Qsmg/Ra
Go22CLonncDBNi+iYrb6gT3MgtMMT31eIgvJrUrxFJlGbusy3jrE6TS7cNo9/Uq4
dgGzUcAYLUE6UIBvnpjODKmQUiwQh16qt9i0+jCQgzsP4JtlqnT8fI7DZ/fqtx93
e6aJttnUhbIrdqRvIovsCrbUxFd/fd7vsd0e0URVw9mQELuYTlvwfdqzljr0HH7B
LxfJ51N5wmBoztc9xqRNNU2VAQHIY1ckIxBuq/ChM8SyOnG+cJHSTs9qVwjD9ZpB
go+TMt0w+DCkpH+8BZNQHzELJYaVrvmxquA+kOj7NLFzLXvKJHaRW9U3q/lbDTwe
wmXub7aOxazmU4m+Pv42kJlpIRX2Sh6PJ+DqfctiVsTHo3c6kS48copRyVLPUDCg
jwrY4WyWjdeMLfl0i4Md2W5ur4JLI3icxz2MFNHRGjYLZ9OQRicIro0CSL7y9Q6Q
34FdMjuZwJE8sVcO8NMic5Q7yhiTXjaneLWHejxsfdtWQYV0zFuFo4LxO7oJ3Qmp
kXCdwMGJCmRAn5cGVpTmhiKcpLlu5f4I+HN+IuIxFLxNABBMJXbPm/ZbOi1bu9b9
ABORXmRWH80vWGS8nT5C918qCjmJo1ZwwL7N7m5AGX7gODziYY0j2WY1ybCFwoQk
Yvg3UjCTiFvc6ucey5ZmOMyuGyeepkQbB7rm5t6wXUC0hva2DpliJfkzFJYypoWw
r/V92qgW7JgmlPSKUV3PAblOEK2S1g97lq+1BY8rfU3OSvR7fKg9PmIeEY2763E+
9LlpzkGEpHvpMVkx4M8i5+dJYSXZ5mqjhxx58NRo2c71CxT1DcROWApBwrIZO2Di
lqDR5EfcEDOF/PcY80d1wDRSKDY8CppwGHuWhN4NNJUoNCinIrOVjDdQO7zeFwe8
oHa7fFwTk6yHUt33i61HW2NBjGKMKVOHjDGxpT5qlyz3vh8ZvxnBoaQTqsjOtQc3
rS+t01+DC2P4yv5kOCLzoC9CVpBKaJlU6MDjvj7gjQHOfg8Xs4L9KxCllQ9Rb6yN
bAZtMlZU3awD3nCbsYpAks5DWwS82+9Hjh1whPY7gmfp0qc7SChbkwWnPcwb6Izh
eTzI8AWzyZE2cU4SMiW5xPKMX9OziOhk9fyj/+63kUhvdTvAmxXBbYLA9LUZYhrq
jTGdYNIoNed1AtTpp4ecsDUjj67QhNpmToPgp4mJBsWf3PXHGQzEdffDkGntVSok
Fb1Gq7CC8jhDKM4cr8U3yOaemW0oYDz8EWJuoKf9OB5JXCoCOfejFXsLJ+nlhUKT
2LLoATX6lHyb1KCHFKeGcuJK8cFVz6MxzqvTsgHbI+9Vbt2JE8dj7+ysbBHooXM5
SNl7u9VQ+MvwGRgIz2FJgKsCzirUB+T7cjT3HoS0AulKDLLYxbpUB15MKJujv0HQ
pCp8RF12XktNsRzaQFCzSIPV8xGy+BEagu1WLmUg0ofCFMM/a6/uEpw2TNI/Gj4K
xm/5orWQpH8jRq8fpryG0U+XB0QEz22k8GIbFE4oYQSb6YPLJJmRFI4NWRkaolMX
RMZ8FAUQ/csJdFPphV7FVfJE4lvYVmkwu4R9HDbc5E2inCk3XpQTjbUvELUmdt9S
0fbGXtReP+i3gBLBsLLj3dIZ5Ni1v4/ewvKOMZ6CjEzuWlgfcc/5RfR+VvNgcEqE
u9A2PZJREJwwy6OoJQulvcxP8p07ru8hiOmLMcZMgGM+lomTY0DI1VyXKck/jvxc
n0NqnMEHck82S5/HbzLX6pysNO09rCpvsBxB54qs3CFafs9ApFANWqU6C+S7fllx
L4pi9wRam1KscW5eVCxa6+MM6OeWL96ORZdmhPakBNijsndN0TH/Mhou7IW5xeS0
zhyaJk3gp3bOxqqgoCjHhns81sHkDvvfRd0RvR2rp3OUli1JUcghRttPgjbewKzT
DmPNiUW3uhDQCRS95hx6LMlY1Jqrvku0WD/iXMXxDoG8X1FRn257nt0smmlklYK9
uL5TpAiWrln1Klr/FLfRpcE9CBgAihzN2j9KeEMfCMMctHZzBQiaiqcx41BDvKG7
EddRIlXL6bgX/2aBZ5XYRilOpXfQI1Tzo0E0QPKmb7uN5pz6bOEsk2aryzx+8BD/
5q5lI1ihYpSvUr9Xdp97Iy8wZSkGKvH5quG5XdXEmANTRTRdB3DaocSdkXL3ub+h
+V06vMyNh88lL4aadkovct4eqppi+dQoUDccUIdzXPOO4yl4pblnl/f1HHKhJFNu
mediiIEI68VkNN97+tud0GuS/YPuAERTu+2dqj9nScUW2GjC+/ypBjJB8Qcq4zFE
5TUdX7p66JubSsKSB0QSWN7gXMUwWBPWSXjQld7V457b1wI5g8WAWCIg9Y4n0zPu
8RhLvcjsPJHPn2zAH6rYYmJvOILXzCvX3uSr7RRKtfp4eDI/WvgIbhRhbH0/vN53
W96yvyBh/fT68wuzwZGulYVrZUCB8N4ROPiaRtp2TqSqNhq6+cjTGvsyJpEbR5NA
MMWr1wcUooAg+j+MMvARd4TfJoPxG7upNVsGAbuQUoRQjKNDB/m5jugPwiGFpQe7
pTQ5+Ay6ZOjlh03+79FMtydUfERyJRxuv6Y3b+B6aCh1JDRSXkrufeaXLpX7EYJL
77aikWhz7k7Jghf8+CQtsVqQnMAXZvbdKRZXmOh+zcK877yt/IrGYDFHSfeCpnF1
WlB7NORlQIirJ8bevC9SWRT7/ZOln2vMSUgG22sp+NQPv2Rlk1nLmcU6T0Da9YGm
5au7nev5kkn336N2Hm1CVR3yN34AQCnuOFo0zkvngeceHXitwjm1fMC+KqTDqFS1
A0oBx57Yl0nVmvr5F7XjhLBzUkQT8shyGT36O6nZN7hC34LBbFsYONsmlA1/6FtC
ymr6TWBIXQLD/uA+2psHXHsC5Ajxssr75XuoXkrNmf5AJntKfPN5dhi2O+syTJFa
cVxVdm364lbzXcyT4m3Bew1BAhWBgFTcO3W6A1ucNfpk+OtUmiCrzqXKpGkaTirm
bGhe/deMkU9NpGxDb9/e2Obl+p6gjeYy9UFPpgAS3UHiKnXMBNSBttRQvKfXluao
giyKTJqcWnuTfv30WNMukmFcLxrdHhUSTp87+rNiELKxX4UsquNCCcJ3AT199jhs
iaI9etHlZiPqluFWfA0rQUM2wfK6miKY1mtiJeY3xU0dJqm0rtYpG01gphZMRnc9
7xjRZUK37BiShzzhHyOyZn2ettWMnPu6myUytcSfW6Dye9ExB9lQSbiphTpQgUiz
BBMfnK6awb8dhS7630cXmTIwvdV5SwL8wIOK5Y0Neg9DPP8oXKH3Phw3Xq3dxeQT
r0+IqPEqr3wWCpNavwET0v9yIVmNJiGYDowtLxramxms/R1Hbo8LsgHi3P7/8HDu
/zm7CyhrAvSxHRXhiOhlLEwb83j6dK3li6U6G1IswCCKE3YmpNRsMawzLxvv+GDR
a65lwE9lKiduDQzw4S3020vRO93oCHPmkldnHpRlcqLfOFj1SLqCL99QV1jmFFZQ
dsoKX+IPGBMBFX9FLJTKA4IRhSjdimXbbtxonfMYyQKqUGptrNRNKfg7jToOysA3
Q0H+kA+UeZJjTLa9EtEqMLoNNljyn/xqvqSyA5wTYuFWHGq8QamUvdeuLH+2kxLK
ide+Y0t2thb0yfq8rJgBVkaTCX6kygDuiq9UYbwzvSP0qQVjiwv7T/IVL72aghZ8
77b0dcGS+/C4nzCpuv4PpJxP4mZuc406rZUtkXL3yi1x8ICmwUYU5cqe8lVDsg0/
5YtimZ5PWIU0ybF7ZcIq7dI/5RwuTEKMLrXCAGkQUrMoLxufpWWsamXzvpw7DrBK
fBC9paZvBNkNqPHpYPMOX02uWsbofEGdW6VRD7m4hWCMUfd7iVABBKGvZKF3MVB3
aKPsYltBIKUjIJNB4HLRf41dmEFXeZg1lzQt/ujGZGBrj1JNuMFp/IuO9BMetwXR
PP4YxL7d4ZMI35dvHo8d+UlFa/bWU6VPXFmtxl/YPquWz6+7TKEN+yCo++U4bUVd
+uMMRtrRBAxkTesbPXXYzb1wzggUy+y5wXGvy5I+RMCeNtObbPgCDfuHEmJK55La
im8WSpWK7J/43Ry23BTrZx+4Uoi4EayxiGMkac5E3aVIjz8OZW8xMvBS0KRSHB33
tKSqljGjf23EhmepkwuBvYLk7ixBXz1Pzz7R7Z4+nDPh9cN5KeGvzkpnr/4uRj6k
lK2Ebc79HIzoB18/xGOUE9UdtQhzfTm0A3pXBgVNnhDdvA0Getn+b+q4Njb0fHmH
ngvdL//+93C5Sk/c0YHKeGt7ohtj347EWbOkYG/W49nsQqGUXkWbYp3srODBWuh8
THV15dN0xA+mKfoJ+rylWrihPKVa5j8YupD9dHotc8U02oqx5qIKPpVz0AiMgL89
7Ajvq+09T9DHULzVssR9N0dK1liYM3TEBKCCmtJWnNQ3gOm3eF+qt/idroLeS1Gi
6rQcGEfDNVyScFIc7P3Zr99Vl/nAtH21T49BiPCogRSJdU99wr+VexPuvenh9eU0
pls0kYy9wAtQGlEKlBh+s34+O5sZSk5HTO3Qn8hkQ+a36nk9O5wivoTicdfRln51
NkH712jK3KHyJVrnqQvfN+F6QpcGXp/JRLdnpEXUsR5NjvzOAaOX7JIaGQTy0s+B
JOyJt8e6vFsk+VYZItN7zQPNSzxqm9lScYi/6sEombAqH16GtG72A425HVMZCsxF
TOCEfso0YD/tyMRgO2LUwqeOhFsKoKMgrx82bbehIPzdXeBBFtXZq3aKpgNGTv/R
0IVENPOBthRlYhAgg5Ft+xDb7O4tpj9D0JDnNoX2rs03JF4Qx90pbzUxPPRJuNo/
1iC2ztqYkhymBiJJBFwVwYgWneuypn84DVIoaMBSEi1htlnUy8R9/uaijtMYN/Jv
5DWm6w7Xfj41jlQoHG4N77giC3RRxjOs1Vh/NJSSTMkKMINrOWL5/5MWng2VvTIK
y1iitpCOObCVMHZQyINOXzbBRSiga+ZQ2iIvw6xjbUtdEq+cibnU5+6VGtIbygFs
zpbTY0WONjAIL3OZhn2fvTJu95pEA5lGWiEpxRvf2utGH7HCaMabJPR3gycsFRwr
/nz8w0IbwV4z/8OSpmm7kTrJekHfs+rv5W6XFIA3IVMbj0DoAqOMYpOr7TX4oMYn
kM6+7Z8WZgZYQG0YYIkBvTBggZI3BqNrdHMyhkZaxuTc1MEIV7puv/QNpKcfKfai
TqjPsG1lIZvQa3lLiPoVVUp94qLYlUf6cpi4gc0lKNSmUFvN8hezxFzYz/Fm0JV9
nUsnB3hFoK4pVtP+haChouBKtmDXmgm9unrBYgQ36su2ys4M9nJahybQbO5ITJwO
D3wwSv1/fazc3FxN0E+azQey7FVGbIKXldFbX4KNgBMBeL9hCKXOaJwZMDzsg2sC
675zOIjdlx0fhFvRnCPHmm5bTzc0I643lpvAZbttmfz8df4otl0Mvm74Wtt/DkM5
cmiiBcHKFfJrWG/0SI/UerQ6N9eR35y1UqfMmZCgF5SO9rtfLUZVGO9H+VQwiqSv
DaIVDSjPDer5QO0uiDPWPZltwHnHoveKSbJynXkQ7oNrtbbbT1MukxQnRyNjaNA3
4DwBEOM7nci8XG/9GceXkJMhr/qDNF5Y2/gLnI7TW94Tahk+vGhZrT5VQaqd73LR
JFk0vjOfXSXymKUojjJSs1BflglyyI36xr0rLo/uShgzlIF3hNIV4HppQ8lqSWDl
AXdxKOCKBTYjoURV++iCZPQ5iqdXxPCGZofQVGoTaNOrC2hwIaDvurR/yYcPGfNL
Pa9EvDlAiZacDu/8G0bQLnFez9Te1aKk228xHZ6u9w0yww6SR7QLPmWqG80TM9sg
nf0MlPOFGOrt1gVuGYC9yx3aEC3i3sSnWoMIerrLNWDy4bM93S+jXfXt9NPepOJA
nnI++CkFKW1+kfJ9jAQ5e5a6Q2tkkTtSOdkUM4JxfSUjAfDvWa0+LvLZfm+1UfEm
rdrEm6bF7RUF1pL2RVP5ED0m8TeGtUMDfiVD43ol2EL8CxKRE0DVw1YjBIKHkxAe
UeqYs3Zy1lqJuqvws1rC/v9qnQ+D/GRHFVO341wgal6YiRCx9DYLn/OT6voNXLeg
hF9+H7gQLwRMbzElWMssLfD0+AJmoGu4WE8+7LiDpTIB0lG21oLvG/B7WgAtIUSg
X7dN/38oT/VqJn8w8n2QL90oEDakR9I18J8rhboO+IDJvhFP/m7/2oqsYCiRw6pE
huJpYEnBESj/d/Nt327lFfKmYh1ajnCbPqLIaTDliMBZs93gFFb/BVmh/u5m03mS
+XTe00cEMnHAAr/Q06/9QLNaBMSUrLBjg2CLECM+NOYYLcF8i1N9QpyxrAj2tDLg
Sauf1WljV0PFLgX3ItZwm5bOzEdi2ryMqoNcoHbJDbxixoQTgTdouwejRZAO2KDA
9pwWJDu6EG1POyG+ACn/1yMuGd1fRTRqJOI2FhZaw7e6G3mKLzXhVQFl9IaJWI5p
x47gWH/omI240Yic97xyLYgULn8HhsxiXFaOCpQH9mQ45gMMYa482C4niSQCjwMs
t0eT3YKU7ZIOPrGzyt+o6WCE3PGvC3WH6I2kN6GOGHrqzoscgld3dfI91bqB86yp
oJVNO6Qtl1S1SzodhDlR1UtYtkqlcusmV6u0o73BqZUqh9hS+2GVAUJICxA7bjfj
KeuTYt05DH5/V7ixIPhRs7TIthqL0rXig+MRgcD1ALEF/4RdhCqnfF44JX3g5OIU
agwwOA8IqOZr4+8ptQIY5BTnSAxxA/N8HlpShlRXwsfRimsT6laSgNY8oYSNKyxV
MC/vrINqnFZQRHIAYN65ofWNaEVLdjeCDfs3/I/TJm97Zq7UY0jkLW+sA3QtAXU2
bFr9yG1CGmZp42kV28RXkb+kWnEa2dHy2wbocycm4CoImPDN97V2zJjf0KwWNmdx
aM2cH6TteVqiFmnzGE44UgrVQKIRCuroKGCqdzF2BjePNuPY9rty7x3UC+sHJcxf
z1IGdkQYASDYUsbyPlUXifYCVvACMBF3SR84imSfRZDdal4tmEs0Onz6eu/kCemg
nWCfEZ0YeGhD9qWNN6CTw0P5BCFgUY9/z5vjeHZ8ndJu2FTKUsYiNcBawMhWbtYX
alIT4sR/GODFnBReVXTP5PzNVvgD9gGEmxCtve4hksbLw7GbzAWaBEXwfIyHU1jK
agohRQFZkqPoXyiSdMNHF4CIsedDihU4tPg9eAiCO7xX9GCPYbTMEQBIvS3HG5OH
XRBZIfp0BnaP/QxkEbTwB+sRLEg3/nQ7lHcgt9utSysN6RWm20uUhbWx1bIv3agB
XmeHT20pbjOwYE6k8w9B1oDz0qLWh6BdYfxA1lC7RJbvvW/3LWZSWbuyQv8wKyVA
NyOtO1ZCvk2OfyfouVDL4WbvsW0ap3gWB6jK6NGZWjCwWOPhfIeIISeBnRKELN2Q
5/Gk8W+opQbKpTGAf58U4w9N1D3lorX1RoGUjemB2DeYcz/eWPKq5KG1IrgqUADP
+k5A9+UZ0Ck4VyAzSm7k/nu57Kl8DAIYH0OOjw/o0NSaa+9jIEHvMnqsk9pgj8Oo
WH067T4mQ55twzVGErOi3nDWV1FR1OzG7iJRcVB041kDDPzoTy/IWrbbI1ld2MLt
i1ncaB6L1NIOM0ByrWICmOsmfT5m7JqfWv/uSqEhnPgmoA8Jn248D8UAVVPnNGYo
Qx6Lj/JKlFf9WEvVOqmWLmIqC7lY+UtzRy6mAuUE/yTAQT2PI8nqPLjvuHQyIm5W
Tm8yyMt/p/vzya8ouwB22t9hZ8KW7prJIAEBK2bHsuyLQ+qO1Q21GIVGkd+73OJf
cem57rGseSuFYv8sGlbpecNXVycMjeiiaxZ1x0GoBxkqlA85IZ9Kv/x867aulE2j
BA0UVMLEBEjNKdm/1lZJA8lADB7C9G/h347/Tut/N2PEMLfx/DDdzsPImmZYrzW7
878wSnpLzDWM3QHH/2XKZDkBySDggCsP2c5DK2oeKr8DTmEyBjzs4v8BzHiVVSsM
SEOE5ZDfYQmsf0PVxajXGeVRhLul8kjjo2r6MVwT/cQwWzIaYTq4KhRTKmJ9xMbm
K/enT8fMn6aCeMIHQaCIrblhMyXBIzWqG+Bp5S4NgZ3VdGl95SDc72D0zvOtZ1pB
VW9/TgDwu5OQZBXgeDYeEkOihVAlMKnvHKThBDmX7tc3TYZR50jZKbDFCgEslO/u
LN9BTMDskXAkxG2SqZHjtp+q1YiaVgjop5tjr5LCiGxstIv+TN1xLEun4UAy6hV3
nN4OHzkjOZv5uKuIJP9cRBAheNEtrxDtONOF8zDGr0zT+os4XZnSr3DRteGmRsk3
C01x4cYfRYoLm6oNzx2YwQgp1stiHfWIYuSFfAV9rs1sbjXJudsZR7Bkp2w+2N6A
+vWRjPaann8I8OIHmvQRMLvV02pb01Cku9HCC+YmAdfhepdim8wp1ZNQRtJrleQ4
6Snt4njJEzD54lXH+ay4yBIDFDeX0OiviSvjQPWNL8izmwQcf/c75TqgyNcJ2iIo
xpjiwYygve36j8XYIIM/4r1BqqZJ5fK9AD5tt+hc4h0moL12tL6O9DxRQWqP9wwa
l+eIG6arHgoG5BK5HxN91MWijTdDD7jJeBwVtx5bVPHkigRu1B/bryvCehS4Pu0U
E193PjRsMcGG31LJkNJYKHoXQDeaU6SaOdVdgsyEB3I9MjSa4xwbQZUg2fAnHCLc
4fAKyffQg6Nfv/KxkAP7UT76HzgUdHlKH4w4ge/zSzhsCpjYyyzXzd4iFKuohfUn
YEcnxTs2Kc02PyJ/E4FK5V72f3HIjXDu0nl5hpbZV5I1u0CpaxUV+J1DAyqqNL4X
9V8ygYXhzNOIO9bYlQshYK81CUOLFk8WUX1tkSAdd45AQwGo48IS4M4tcl+yriWu
pTh2B+pM2zht3gpvoRJqEx96JGa4BTRvhm87QpP2d7UFXDJawDp4vJ7HGSYeyVzq
AatLectNNyP0wGOrOqwJQdm8vHET2eaxlA9YqKW8r+q+DK2/1ud18Lrkzg348OJi
vWDQEzGkLUsOlDrVCkLqCdfi+GhX8pC/CG8AYOk2fpCfRH2NpRmBQKBE9y6ZYlqG
CuQnDDTDV9t2J1NpLJAXqh8nC/ym90kj669CD/UT2qMCZLS1dO82j99htMSIzENf
HZkhv5T7YR/YcipN8pK+FTksXwmeLJ/HE8AbmdRksT45HNNwOrHSWb48F0y5RXc8
M6lDNfKlRGVc20NNOOfBJ3LfkWLXwmleEfo8xWtiay0oLjkd+G/YJi5Z+dRcpIWZ
NUcVDGyid38+AplknlnNrIdcpC9nfoUi6fLPL6BFdUjcSmADf4Z2vAqx/iHJ1L0s
3nYdtq23rwiEQUf4haiS9czjCv/EpuvZpJWQPIsaJgnJ+6+eoLAdZaDtUf8xEG7C
Bz5uJkvI8p9uaeUxlnNDoUDY05y7XruZwuiuZsSOVFKxncK32+0D1O9f+A2qO8VK
nAlEvECwlW68ko2I7zlDvy7s6Q/iz7isD5E1xhRHjuVfqlxrjyXIFlgulLbBiWKq
C/f0swGEO3DkmwzEYuMXA5nN/NyRsb1BguFqSIVhDwNf0okTg/BeEzfw4NbAczJk
Wt4ISVUuWFkISQrBY3aT4nXDQPncAfFFuaSWkFaC8mXknnjiAEYDlAhdf9xPmpzg
OcPOSVSk8tfnwVZiicyevyhRJUsbCaEcq6DeQNWKjbinYSkpmbxZb7xm4gryRv7t
9TvEvQgPbEshs2gwdZE/hIDSNu6FehAFurYtkc7iRum14YQrBZKxTwS9OwoPK6K7
NEvvlUnQbWUyoseJ8qtpm2PjKeU7om29nSXO89BoHYCHzXdkDKB4FsbnCVXYiEwB
40hRU7k8YH948m38dLR+yIm4mQE5ITR9hu39yw+gcsyP0uISis7NBrmJffa8bG4l
7oRXfdN1wbTTvwFOGZVNQbR/sTE1I1mby0+NZyrxEYopDL+4xU5DGtrsyJoEdHzO
v9AMt4QpA2Xyh8+bTXsrqoi01to/wO7m4/d6vSv3PMsVgsu4KBY1DQ0MIpacJB1U
d/8I1Z5JKA0/1kZisSKhIrXM8KPBuJ1uzoFzHpGCh4DD9YPKRYydFBXkEpO/5FIJ
38H6PFpj6wMkXRQZbncwlE8X+oVkyin11vQfe06Tm1veATO+AWfNSDTFnj5OlsPU
pmur3/PHrAQZ9HDqvw4Rnp3NCSvkMPFk+V/tjU98jhwBx8RHVjeVLJqQV8keBa/e
o4PgV+ikh3rFiXtB+K1fSjFwRuGwDASdGU7bO3ZrC8GJi6FO3akHnYak2Pw+qKxE
CrBeeYoj+BohZHimiBMM5xoojwHdRy8PgChT5EgRQx0SqTgplp1l9o3vqZHq20l2
MiyXbKHh0p8kDyuLLdJpr/UT2ZnNNXpOJ9l/O5woMFGUuq4yzk9yva5m/X/Nvl77
IfxqW8u1aFjxSxvnoMpp47zdeEFfvqAJahwIz6V5RHvmXlsgmK7BKn0TKDf1TkO+
Oe/5SwcO3FHf0ypL3Vq2KwN70kXVmrvJiPpapex8ySkBgKgQEzNrTWLayMtp4UW6
3rr0zJMMJ0ZVXzFBWjanCtviA33vr0SNgd+VQ2HrtStUrGsgyWqjq9ldjykfd4TZ
WJa+ggDrnenbWB5kxDSqOynKtBcFnEE6UKA7nZAZYkRF8PXcDaN1a1xvmbTR0Udk
HgQsprxsjgR1gizXpBqX0siwakJMJ5AD4lNMBBBmlqtVn3I0niiV0G0rIu0FqC6c
m1OE7EAkToTGCC67SBYADdSD0VEVxiyuQbkp6AeBhULiEin0bs7uw9+lt6obA3gx
KwSSYh5B79lj4G2X1yfyHcXcHIJTHPNZKMgh3iGM+7Ga1qOoe3ztRGzF6V/hF2la
WbsbJ28UI2WZ8GDRZF6JrSej0BKrDJsZ+GqHOavEyJDzTEIMIDI4VU1r4GfKFOt4
euEOVoAY2H1WE7RkcEVPQyAe9uWGvrS+/bGlS4iRGMFh6PERA06NSm4cGCTXyDxO
NfCYY0Ko4ecRgeB7Em03vl8nhzYYwo4sY6WnUnjcAJZ0A6Uru4dRHis0YDjZlAS0
AJmqYwxRla6RmKZYqqhhkkLl0ACl9sQtQ6OHhMuHLjdhJVKTJPv3Gb6C/7K+xs1a
HFb66IPJ808oxIPmtY7t3SXLFScgHO9YGl0mvfkUmhF9GFTtg0B55ybN6CD60mtf
LJG3rUMlKO84bosV0TnOGt6xWd/PzxApHsk1fVgopLP2GWQVjMgsYoMDNI8zrfcV
Ji2AZl9q+OWqodT/6dyMx+FYsiPXEBHetQaTeKtMwDj3OBSu7I4DHIO2diznVzSn
iwc20epikiGaqh7gCyYiZxyw+dlVXI6wrThs0rfGYKca8KmEDZu/fyzqK5v1SbxX
w0YWu955r2cG5ElGBf6/z2ixgQhR3C6Pet1+w82JPrzuP3NpiK3/cLYzWtqEdxAI
QWfDLw2KFtd60O2FS2wZcywFy0dpMfWxlAwIbe22WfpuUC9Mpu2Tpy957KQfKO/V
0IPozpasws9mjJLkS+sDJyoPABfVD9w+IU5ixJtEVlaQ9M1/fVxtMqEpUlwnvtQG
Knx7Kjup30BVOJ9LBIHwlvwsDvtS2uiyTZIKKhiPO7+8r+89IQCJ/naBZedkslxb
62UxrzWsvBofuxXHh+E2FGEt6Re8n/atczVCFE767kZlZjsHstTNHFGWCBX0Cnmw
OX0LqGUi3OqIXZPalb99YFJnhLVLKB40hfh2RV5mPa72UpFkp5HdKD4LhR1ROnQ/
W6YII1GTLFHJhwi2mqWDmogHoMVZkPRC+KmtYiw7kfKmUGOXZDu8OpYuhvyELbIW
OgHDc3qboikbJ/O7XQgIUgxFt0f3V60o8H+he1TiEH8clAQlNl3xucg1veLSCI9Q
nMbeVjEvLUNZVjTaoYdyI1lIfJZDfRtJs90xA4pv2OptnO6eKNzOGmjtNsHP2JYe
5FSG7oB/JgvU5uAWEPhBYL3qIz//V7C/2l1Dfk5TFyqLSb9WeHuAtIB67vpOI9ps
7+L122E+v4TsqMA3zP1Z+B8lMHU3JrolCk+FUHgEpJqjX/5SD+l8zb4l6SY15C2X
5LsuMf/tycuywMfFZFn8Ij563fw9ROqjn4SzklimCxG41xFAEsyekkk4v1uC4KwW
l/S7+0BPpJJFwjr0rn94R5dceix+NF63KglIiHry9CpwYhBSo7CEUJONnX6VqueW
LoXwo1KNbA34DLnD54jzh3yBoFDwKfsm+Ab12oRjJqc06HQ3NdkGCpPgmp1ABF5y
BnJoFztKng75U7h7n519sb/XxigZdv2+AD8Jfsnpj/HAxy06+zTwtCFLTOXE/lVG
8uYFA8jmRwBMm9VwrNQrnk1gBpNU3dVrdnqsBMgasP2hsCycbxShzxJs+7QqYNB0
3/KzT2+DF+RG24XItDn3XyG8J/BNtQ27HKD7yorC5yZAwCVpxXUsgVp33FJtedx5
lSuoK0KacA4Iw1t0WKEPY2W/wbRNF35XZN/kbk++/4nvF2ARqp+J9fKCUYg0olUi
sS0Db5gGb6kO91uY2jOQkpSb4HKDhWAB0tbxBoAQXRisV7TbbTZxXWc7PN++k+Wi
Wjgg+M9AHm2+0kV19+lOpupYqoPuEpzQOuwCm0TCweNNsRq2iPHZjO+3+/v1gmuP
2JEdPUSR8QVZq57UpHjJZGlF5QsxtQt/3hTM5TZ7Sx1nWAss2helP6FQ5ZUptSwd
5x+/4X10/1cv22uQYYrq/tuLdX4OiWV+iZ1UdrOKhCVy0lP6WwVsmRHf3Lk5sTot
4AVD94EnXnWxvj/L7qMcP8Mq3NMPfDOEfUDFz0UVZDvjC0rKg1OcTxVgGlwIWz3N
6xnxCiA3rAc7loV/R3ZZgkpDbHBs9lcapzFTwzP7DSeAI5dhFqwc6ZNs4tGO/Arw
dLXlNlpxF8lwe7tj1lyhwReGMfd+eenmwq6lmTMW5q2TVrkrQFVU0oz6DSeGlS8f
jjtVc7er31pP+LwTq9Tqfp8fox1/N4VPOaEAiK36OIrKidv5jgTRcqc+951TZoNC
GdrUeu8Xlu73lGt4O3z6/xn9P8w2PjouLUkFvLIMXbbIdrxbCVOYvtoQCkw0KC5R
512a08zMNDSlN3aHXAwomH7YKioJFNmhOsxvYHPdAGmMobVWFTRXpyom2ywc96+N
copdRfmqc0GDm84rCfTOM7YB4sCszIc5Hnp4F1wla9+qu1WZc2J6q9GkyRH3Hyje
E/zN+MpR+QxIiS04rwmICHhz+Nw0CJcyJL1pzIQ5/yh++/c8EZWQAjGnTmgFh6BJ
ZhMZ8vOQH6KCiS9OWrh7ZM10hgdoJDvlAwpM2RddEjd55Q+ek5fUtC5kJtLxOEIo
hDHMxcEO9mm30xfaikb3TspwfJNG7fsCuuhwPvKD5kA0UJpEDG8JuTuha5GU1gtV
QcABHhUuMlulpmqUxFxsKhRyOYbHtN4eQ/fS/r2eYA9cOuSWRGF92JY122ZpYVEp
tvk7Es0Npkw+C/YhlYiaTYlz/wfKJFAxwa0T5DdcInkRWfFZaPImpDFdmEYWrSvB
fgvlS4cu8mOka1PEbpG+yS2ekwtkmL0NukcsASonrI9lA53bv3xMLochCdVZXKLQ
sYM/y2DL+Of9anMlQrp2KKJkyu4qAi2kTyTLRBrdfdnZKKU8BNeIyeo9Cy36eUn7
dm4aCTQfbZU5DUFRgfMsgrY84FJOkE4NtNSc6vVp504QxTGMdgLC1iOEDsCsUyxG
pf+RLthugkF/47d8i0hpkQAvq36tAVGtzYUFzDi3tcscp5zVChY+ne2wUBIsN62B
lA2OdqUg1V9ruStX2RPD2S73OGPd3gEvFflxtgPU8nkdw4Xl55c3bBV5VgcBlKNk
xAi0lzjIkzen9eXYvHfHnWyK78R53euGdSOfgLN+CGC3LFqTnrUcqMN2bIEG64UJ
NeZbvhl0N18l7AyJfY1WlSVXGL9ghMnoNhobQRfLmHSjdrvZPQ1F849D86j6ZPpS
0sSd78FSXNd7sU5O4jketWIjcYAMuF2qPd+kd09338t67/TyxoXCYJ/L1Ty68235
AW6drW9uQVX881op5Jm+/TKYLFG3EhLXR4vUl/P9ZrMKaX77BNMWqcwC/4b1yoES
PwCF4o7LYtaZxtI7Rkg64KH2zoQkD1IgnSoMAVGK8oy+KfEEs/8XG8XetWMTBJ3r
HlIXCw2YvlViiJKbruNj4KhibRtdyCrzF54/IT0LSd5th3qDAudKAMCI3k/wNTAU
eP0spkBBfyjyWVB58m6+zDa2LAkpS8jErY/FIz9TP+oIjS09HRLt9xUF2oZKfQk8
LZXwQybEL1ACoIQkIrCcEM3Qu4EnM79mCQeSwBYy4pg+8uuAQZKgBC7wVf1qX/Ly
W/WTy3W2MpR3whYR5yH70DrOecNahmPjp16F4dp3a5jFgbdS+X3MO3ABfOquO1c6
Ao88ErIAw1wvZNYDe6UgQncs8WpAAL40+c0Q388C3YrUsWLgl2AVIsgze3GRV+xh
LbIuPXCtG5BVIH1BgNCD2+dDiH6n/VTyZHdaZdJhE+WdQSbZahfnX0TV/OJLK5xf
pCUA1M4BStljNDnEmj9QbQT/SPZEeHV32b88q6RoKMPXGraerYEoh6sdMmrm75H2
sK7Q56zbcpzjiPtqkohmNngQYVas33FkL/SG5Ar802DRab0k4r/PM0M20DhEoloP
1UlM/68703nf90KjnV5kHtLkJFKIP96FsJM4u4kqtlZSmqBg44zV1qX7UO66It2v
V6m8FVtmIRKnGw3M8B5JI+kuWeDt7J5YiGwmhw3DAdE8V6mJWs8JNkrq+xIYc4V3
KaaPAgebrVe5+nmm4u8HfoqHp7Zrdv6NpsYzv0lwYepI4uILdPfiKLHWa1tYqJ7h
Ly+J+DYF+eERnibYn30JvdQQhKQIX8R7etRyr7A0VfvLEY81NC0VSwMwwF8CRYBR
82KtKNcvciG0kl15WQOVV1h3mrRQDlFXiSCGCi0D0FuvBqdg4YbrS+4vdwDhujFR
SCO5nwREx5CTfjp6MBn7RsZRDyPl+mPLk/lP/hOp1s1+nMns6PNLfPsB7z32kzmD
g/uN8yuXf7kKZBA2OZF2vVn61C/SBy+rxxI+YgGEAHgdOmvlT4Um6d1n/aLR2/Nz
7XbkXnx9AvuTEdJLs604jXBO+UTzXxTEvc3+OD45IgGmdOOxXe7vbiZvC3kaibMz
rRemOuDJoFK6wJFsi95D2iUyPrfhnXZ0AHZrtZbt4w9HTpgvPjssKjXVLSh/yPu6
wPAJFxZqIifqaHzecbjI7oMwRi6QkkffqamL6s3/ApHDctIL40YuY+tjE0OXm3ze
PFJZCfPfdxgZvtpp81duMlQDduiq1yIP2kZK7XRK0oQ9DJCTjSAi8bVxVpqMT+O6
31+ZA5UAyPhQUga5PU/06GHD/bwSA5cjotYyGWlPkhtPYru93oGXiTJdC1mmJ9dU
9yr5xZ4G7vnap9h6mjP+O9QIWJ1JrVbttppZXZgBsWnZ9CXdZS5buk3AmSa/DoYS
vJ7/V0I6UFmpRzH8ORXWFWZbU2WGbRuv/S3yQybvRSqOTB78NoTvPC28b8VBcq1L
/ZQNEXwoWk1sQzKkDTPIbvyAJ9o2FBtOYqmcPdEG3kc2xxNSvA/ORBHbrX+6Y25w
FeeXXPFBLAZHK+wTw3qkYFupWupnjwgjLz8/Jfs00rIcDdX6wl6Flc6eTsUsm0ZY
2i/Ji0xAUydoLY44csPDQ07SvewQPg/1bCfSP0/JOyv3Gv7eZs+qG+E7DF7rywnF
hEuBmnK08rf1d3wYOujrqwc5/DyyUXfuLgVnIW9Fya5ciG1BM6GOFlx6HtjaZDIB
GfWOvzLFDDSKU9qteDtJTh/5vJsWebv+hM7++efGzqp2+xZMFhNkCNtIE/VFsPBQ
WSl6EK/tl6FTF7hb33KpCzBaRgkRRj+pAP0ZMTlOZMXs5tDkWccSdFIZHqXdZoMH
i/9l3tEV92Em8pRR/ocpEguTF7auYOovjeUx2ICr3TXBGFWbtjJfEPVQc+2NGv23
SSySsTBxyBhPryZx1v3kNtd9rBzwyJzQTrYGUPRnnfZqnVmsgyDjFhLoS0N+2G1V
COmsyRpmoiRUl4H87k67Sy8fRu1L9aRzg3NEfhRa5TRqW3waTYoJd1XZs4j0nQK8
PjWQ0cVpreedpGFfqAZ5dPjFr2+Ep6Q6OeOsrGLz6JuCMPHTzYq/4DYjNDI1t/nV
TiIPIGkYJT7W8WozkQzuDg9BI67joM2wwwvHWVf/5jZ1sSu4GBt0TzqnAiF535NA
h+0W+ZVNKGT46h3iYqx7VPIluiBJSys8/VcgJl/X6iV8+1vr9yiOO4B/Jdcbcom3
ImodltYcMn1DsPZKzCafcYmbhJu0wiIWyg8hxERGSRL4hWoLYmON/6+CBwHJVU+b
ixHoyzj42qZqlLgXNyW5Z1JlPLvtpavYiUV6Lz6DZlwcbD3Sga3Hma0xInR+rOJW
o4n+qC/4gKizKO7n2OYJTaaAXW5Rx8NPS6EQDkwR+mlo7D+q12pG81sdj7rVJCVc
H4EbADDZpG27F3PcPR80dArA86dY8byVZTITo4/qjdOgxw8gNzv40oB1/19mWu0n
WNCztpTSIYltjJRKTkCRlhbKcIqHVFQXaw5nAForVcStpdp0/Xpi7H/P2r2FZcGO
0ACmQ7pDF1Oxrc0oWVJXq+iXmXET+jX7bOZoLeTBiWRe3ZrDa7QEb0PUZHklThEh
Dv2cgISZMljbHsYUMykD8UYRDanMxtjdf4L5baN2rIAS/2tXkJCfDcnWXAnS0OSD
+JWVrwORZDd5zc0fWqEzJWN1MfWA64Tuxn6bfm8jGLkLx6Hd1OyWwytmXc3l64NG
8zw+APun3BDi0nfdTlme1VCkcNQM4CiTEHfgrkH1CT500Z0lZylDPY/chVpHqooL
jzdjvItnT0N/oPaxkPmMNkLEKBRJRbbws2P/WSGJO2ujpW85Lw+VLHfU8gtq2Mu2
FcqeXUcWzpRHErovYCARgg67BrRWLBv0tKhb4M1pM/hSD4TF7DY4JYxFZDnrXgzg
5IPEEn4To6i2i3+2ffJ5L7iZQEFxaTEI6QeAdCgzPcqwuJGwMBu1xnN31MczVGC3
2gNBVAaL3RQAkGzFxjpC4NWDHEPepkCsfQwxBnmAqKAUs36jcnV/FYzrWtbx7TDD
o9pGYD3MU4RCIHUZrGf9KPBZ0e6QHSYpEGaO6agu+EFHOTavxyUOuuWD0WM1O7yA
WtJPXU5WySS8jcCtqWmkCOEhVHmMgeJKNJ8WpyPejO6CAIB6sfCfuwjJcWCVQmBA
dtE4zzZfhwPtV+1Hp0KVq4LNH1eyInjVWkemtpxweyu1+iXyCBcgjwXIXjPtl/52
P1z23ue9Pc9thTydepFdIznhdzrwIJ7ogiHQlVaSiAJ/nJGcFzLQFJdCpplIJQ5V
OUMlriRjmL9ooNIBIqGhaErhhFXFc26eS1TzALmxfpbjm5yiUjceerpNw8uwTpxW
2PJRi7GWKjE2AHilVd2TtvML4r4lmxOThLMtK7LaNIMOmNszOA0QFkjHCrkHRLf6
PAO2lBG4hjZlPxEVEtNh4kbLkYRaQtvSQp+oZS2eZ06bDW93tNkEvHM296Cs3/2V
/okmFpnH+EaFHX1zd+fDVd7jD5hSl7cMdPY/MwgnTomsThZCLg6zLKyVQWNnmq0g
yRBMkKOZZfWz7wqUnM0GHO0jo4AZf2Ef0gCt1TiZMHkeu9J7N2CF2QMH2OlS9BTx
WorxGekfNqCvd+5WvxLFyr57q1RAOCshiqCyAT/r/MgScOybrjLK76i4zyBlApyD
yEquE0bee5EwNSvteM+Iz94aKFL7UwfpSI/ziw/C0cnrqM5eCuL4b7MbFm0/NbfW
40O6hgfjtDgjgOZLf85vSGtf2yHtaxRDeKTMuGn4560XUo9r8oB35bnRNGJwpaer
8/kloXC3S46AWtPbYKfcKG+vgdIzgNxgmhtEhiB40X2Tda8LPFd2mDn8As1tXfD8
iDLeo4Nf3BHaekjWfbjfUIpPuwQ0uGJI579xqvX8q0YX7Ibk5KZALVDlR1EdADxO
ZtpMLwz1YxnqlmTDEVtseJutLURMzzvoPEBUzt11SUfu1mGfavs3kpbt7OT7Cu9Q
o/Gg/hXH4XeE7vQ0tZiKjRcSOE/8hvRbBHYDUlcnoTpQ436abx3/EnJnArK4Uq89
m1b3J87moZkp7kz5cChL6+ft1B62n6PH6F6D7w3tuuJ1BeKo2HzfaemUg7m6kfyr
2kqaNcwSeI4XIoQO7ckRY7jOIIPcJE0w4eQQ8t507+MXnV9IIHy+lj5RQMzc9faC
VVaxh9ak3fNDBMDqOee777OP/ibzrRIz/Plev9PvRO5Gzim/248sfH/U+re+jHA2
PT0aJ+iLUbaCZQRmMyDMt66fSEW5vinTEI7SUUHbhhVoVD0yf7e7KJ4ACliByPcq
sd2Qn9Hkw5RmplwQIe69a3Er0WHSVQjVVY7IVNwaubbUBtM+s9QziaQVfinH0F9d
2CGs6DKjKFvzF9YNmasikb9hCRZYfkzO3b0sBeZcnSiDMbI/N/dFEDoLJoS5bDtX
CLQ7TrjBWICiqC41snpDdI45yv/ZPsUFnKtl8DzKCuNa4fbb5V5+4SOA7WN6srLT
XU/w2r2SDjVT5sqTbfRYh9zqzln5l7Gkk5jEp8gLoQRFx+TF3EaU+1SM4QCyD2Il
ZBpGvNYnNyks3qXRbM/4fe5CEixR3vuX7n1o/BjMajecLGEpuhvZq77jb/ZXnfqG
ZWYnaRVqycWbRVING7jkNq4oTFQPGI7F6xK5blnEVlIgdzLIv/HfGw9aAdgCStRC
mCyMaJVOC0suL1Jcbl9n6+1pIKlgvNNDb+EqN9Os4a9iBcB1mctTKdro+jiHTSoK
DOnJbXwlxaPl19S3qUwE9vgtXU6w6eNX7M4+MSAs6Bebd5JDpkx1QGbWHM37zBVs
kmp82QbOvTuDTB6c++49vo6NSmZdJi41FrZZF4wzBVaZ5CKZ9q2pRIihECSHaN8I
HXyFYZ5LRtxCzYvoorhS3UfIh3qsXBoqypm35ZLA7RT1UmzTZvt3PKr6WkhvxFds
8pS/oku5qDcP3G27GzlRrmxcjannrolS2IjlI0qjCkSlVSNfDpIRNJNfND29cm5o
prooWqxlv/wUNIM73aoFBr4LXlV4EKDpRvaLPHBTLmbrrpGFQ1hxYT5Px7F/+ojE
azN81P6zMLBXM9N/2pTFVUGnXNsjXFbjKrno5Zoooj39/dhlYnWwLdLkRWURb//H
qfcSVi/5mBN1JtvV1a9Spzaoz06EhAjhi3K/FxxIHOVKFy6Am4fZ1IXmWY7dv5w3
OQ4P7G6EcLVNByeLl1k1T120s8R81buq1tCSeU9rsR+GOxDKobz6/B6lYJ/W8Upc
9ymBdfmwvutCND4eMAVDhJBoIZ02kbziY4JXzfufVHD/C7pe38yMRhzemoT78eST
uYpv/HbJsQzPciUDOGMYBWsMY3UwsvxOEzsLc0Dpec6PouSmhBSq19OBfWmb+c93
1yyQfbjIm6kUbGnyn9zFYxkWZN8JZyIEESr+SHoISBozDt4obSvSQmJ4mjqh8Gs2
J9I6+Gy4Z6kfECxCY4CPJH7HN4pI0TFdJGtNs9qJyVm04lXlNx2VudCCspKBytfr
KDZO9Hk3ERHXdqvZadOQUHhD1xAYOoILaw1ScwxlrTt2ZKaKC/X49GZokMyYF+6C
WC0PS+f9hNOXeL0Lt+EE014fziB3zH9kHsz+3tVSklL4+AJEMjAgGezdQdWQK8EF
gy8Ms5Ve3mUlBpCQo07aWJh8dsSfoPaFTVZy3lyL0r33H1naSA30plU1UaSHw4b7
dpNFAljgRjmYMaIdw/oQRzOxL3GCtltMDOy0alytfBZtDbVK95vlMT2kLvBd/egp
ps3gUhjK2hRUBzus0FfNn7YDNfaRj33gMDhU7JWQQTawkny5Im59SlMFekhfo/HU
aAk1HKLuo7dmT6yzs48naVnCDPQvmvoW0Q/qPvgePliVKiffldcDOArB6IZjY6tL
q3kdTtHyM3vqx+R2DrCza205E/27Ol0lACfIpva7rv60EYxRVwr/N1HVZ+yh6wkZ
LTz8CacYXpZ/2nuvxa7YjySJQnyglpDSdJnn9NnWFvRGpyYMAeTKy8vLiQTLGbCg
RFfcoz62RWEIHOaHvYumNx1R7xI1MxQCjV4XRYeLzIhElLveqPL+ToIkjZRlxyY+
X91s8vgm4IdY7dCy+vGbf8lX2BQFjuxx9s2E3LeUz2v8abZGCXlg7QhZUCeM0VUM
d1L2KOkBnZcCnM5rjIVGDm6C/+hqLt2GIqu7EQ6BlHTQwNjZBgsd6YXbenmk8F7h
4muV+wMrqipFHWrkyvN1ThPDQ8EWt7iNZ1PqXYmKTJTbqEWycHXGJOjytZTrbuXh
fc9QARcK6pv5ZHkCehp5q4Nk+E2AlNnTfVJMpTie/fgEaJBQb+kE0wfhoU6td77N
i/9Pc7WvPRMTYzWsCPS9TwtftQX0UV6zI5nxBb5GlQ0veW2vEnOxM700jIqNZuiU
1X2pl5u24UHc7wKSuHK1gtkAuRQCZ22lQcmnHWY/wvIbEAyCxBEf6B/mZo1dVt/D
hnZWiZuLaBqWL6u28ToSG9eO/UQH+bkDyIUXLES/cGmIK+wwxzNSn3BE5owTsNc/
wQAERg8zxSjR6Y0xPa1bH0i8i6O7rTSymqP1cxpNHrpn2qROZUxajcDok9i8w0qq
Dv9taOSPCkltTkNSjVaKJB667t2CSNykb5APPwBY50HThF/fJ++ATm8IQjGDp4+S
hxCr8TqiBk1cZ5dG/jQo/UdGyIr4zld6jrA5UPGYCVkfb0HZsJUIWFp5sZPXdU7B
gFMlqhqiUm2HkpSJdhO7w85pOsC/fliNJTx7JSBLAdFEe6J57i/GgifrhNPOnI93
9eWxMm92Vu3FwQGLxNQQWeyVZ9RP9NRw9x5MOuurrCCXq75Wq0IJUC95RTkUJOa6
dltNdWlJXHrkeO87RnPIyidiPoMPcW/HVlwwx5aiv0yKgC/buXuGc4llqdhbZWCe
Cpsctfw7lXucMh30vYJITqNyLwCwkgBePjb8AP40QfbQLfg2nb9zCnDsohGc5h/1
Z+DD0Dx1Mxilu3JZpt8vuXeK9jPtiaKUzh9M0HaEHkC55+itoUV3wHBwffgI+i5x
7CTYiu/fZks1Ck73cY32++T3wHwRZPmRRHB5To+WQ/Umfghj6jTVE7kb2uVp/Bld
LRHT2BcNSC7XsFNKsP3TOur5FVuqtWa0Zi/LvZ1lClxybPnvzVQmxFx5Y5p6K5Uw
ZoZ04saDITAwnFQd4coi50p/alJefLA2VVRq5eM9JK8q/UNeOVLcrSJTOlfiq5sE
4rdQlXC6s8tsAiU/LzXROzQJz9GsahlLdP5BAUaqM4PEgALCBlk0Xzaehen2wNlu
NE4UCrMxcJ5u+Sx24sMVXwvEnxLGLAOUCrMG4NqmjxVHTXKcs6NdPtFYyb15rPza
2IgVi/oN18mIEvMzE8ry9U1qGW1HmF0QKn/yUkT0CWWcRJ4E7xT5wMuVcjKtwbiM
ZD0O0Jx4F9HUWFcaSy18GzRIAdsJVjDX1wLyiX1bRFlzwwOG8FSRMEK80Fx/FCOJ
MZ9oSOpjwG1zmDoUSPZIl8WZOUt5qAfYw+L8HfxMwYiqcRJ7/g/cKuL3uB5vHAg4
auwMkNMNwlRDv29tE4XkCwj6BT3Lt6zM9W4ySd9X3MN8TfIz/2oAkXXdvzq56+Uc
PDweHtm6IltnzRb2xg8zrNAIg26BW/kTxtVSVJi3Ha+fCXCjWx0q+2nVzzaKC3mL
C//jLuj5tCt/4de6NZdUSULEHNTf6Zf+c7CV/y7wowcPTSnuY0tKBifx7qeNCMXy
+PsGJeXn8n4W4racTqc3a4QjOFNjzTqgBV+4AKLmmQYV4ood51ME8TaAWL32krhf
e6aae7gzxrtGbg9WQzIErcDT0Zz3HkwiUfYD0FX+mUOWzbMNBRXZUkthpWDpNeye
Ty+LzJd+ezocIG3bN8VI6IwcLiq9Vjky3GFaHc+P1uu7Sy7VOBxjkqAazKcpYFLY
cR23JbowVZRTGrivPL4iw7lXT51szgqCVd2uL4KEuNLOHRTHlGwNpebolc41OK9c
9Asw+jy86unDVN1e/InZY90zU56KDmw4ORe7+tRuCSs9eCHaP/k/tGM97Bk37uCZ
s88QKJoIauxiVle3qAgVmaWt9NDZEugYXvhlzIBDqIdypljyNTjtSpk70/kUdNEs
j3r8OnqhCt+5yn/FybZ4UAd+b8wWavpfHS1fgMWT2hR39P7X3klNnGGl8dF4BsV+
teC85GXqSwrscxhHxKuh1t+c1HNmXNAIiRExxkFPVFp3TyYbSoEhZysGawO+kGTY
l2rMBPx9nrafcIYuzSw+ijQBtsq1v8k09t9P3EVfnsiOstxD7hDOR9+2BhPJ/OtF
FkRzHJf6H6ZbnHatH/zr6eUpknr1D33oTHlAXH4sTFMmxG/tcov7CdbazkKjiSag
NAw8MFkxzqn8HnnPJIWpPPotYs4pPu4ijnx/4BBG8KxBAhr2QjWhDAvKrIwZnB6V
qLuYgAzUUyN7yO9C7W8rr9zmufKwU5IK1BoPEzDkNOE/VHG1EKOWEIRUrN1PLaRo
ItFlASxicqQ+JyATm08/FvGl1zzIw+WHK8M4fclDbNOJCjbA39kmKIhrI4wvJwrh
7YEg71nXZDxsETWYnUXxDXmBw31PuB9NYk7stFo0W0BIHbQ+qjgG2W6bXHohNdLv
5Gu4eQg7gj9ZtF+6kuF2GgSJZzQNOSlMcR9cF9hs47J0VXWz/5rEwPGuHKlkidz9
vKu/iuGqyOVHIrKaxWb5fe0YCXZlm/trG+p2pDXEP+OMCwMoEi1+ceKOCZtqEuUW
gmqmv/5iBvPaIEA/BjfwIjvvN3anh4plODZinILEaIw5dPDMVC/5jOfqn14oHS+r
6VICOuVk2mNmK93KqjT/1vFImfc491C59hal/A52yQcNdDREod3fVagqrHI7yrv8
Oyku7h1GZxNsb3KAp2VxI76w3GaseiLeeJOCZOPv9ScqP3qwTwFzVA9U7S8/xX1s
qBqg5GJ3H/jcn7fzFz6m/kCwH32oXnrwixfIicl1tTjQdylT6C8AK4vusoFUVgIU
M3VDlkAwhvIg4zawfwDFcvHHbmqAwSJDa2K22CgoJxfeS9P/TA9gghMyFaNXj0Rq
LJAzxxrNS78IwSAsE23fuZ1jXA9+YvkQIq6vJ+HtP748pm1HqQvrcrWTZ+P+gpLL
0+sWUMBw5w5QD1La8sUPiO57cWB8ybwGI0WgrhXxCUSshmilJzw5AUkRdG4R0xFT
rLXBmSuXqgKh3UVjR6LUwIbUGampZTJDjxXhp63dvUVwCkR5fAYymP2DvWb53gDB
a8mzR9ddb/Fu0k23RNcFGnjL6VitXFwuSXccyrR0jWiwKHMhr27MO5vchcdPpwuC
asTXyDfn/JjTRHMIvaoWTyKTZbdxzKqIVAS0NlrQ9omgpeTX8GHRZmLfHe2UFd8J
g2dr8aDbEfunW7mgl9v9eJ/QCP0ZbIzn6EzirZLCV9zGBRwDS6KFMKnAvKL+Q1co
dRFYNgdNAULdqwtluKTldxJ8RgKsGtOpJFlgCho+de1jnnLsy+dD5c57i9EVttRk
XfWP1lDACBde+iOLbjDAKHOGLBIUzXKQvD1NNODYjhJb4Do6VnZgqAk/UeXA7CDi
f/fuXLddBltv74lylBnfVhm06E+NWYcLnr9mVlCzQzpMdrw19zDFxKZuP0QgKosY
qtJhnOon+g4j0hOy1nzJfpo+Ybfhul6laFdhxfxzBFx18yLgVA7v7B1At6PpvPh6
rwOHm8mMs50oUydOgcPxYrJQz/6wy9f4XGitTKvD3oD1SHw3cdYU9lifUXWYTdZg
C83/OP4l4imM1sL033xzR06zdfCZbChbtVyoqcavLziz+FJU5eTRL4kIpNOn26ak
vuYsPsKWcM2YaxrkoFHWhu1yfp3IruI0PPNWXaTacEFevhtfk5nSNDfozeoTs/MZ
owo3M90w41t+XWVKMruc+OptHk26Z56+2tT5I8y+kmErtGtk1ZyYIhkT77Nusg+s
I+H72a4uvCxEb7Jc/3MN6/JLb/ttWbqqxy8mvRqvU5MLC/l9Drx4qNa/TAeI8sY2
F5ENdaM1mt5Uu3fH0h7ROarSZ5BMHfcX/fiGxHzF5EJ7dxuWd89ThuGJgrw+Jh0k
KeHQUV/IFejsMqDINmJT/am51YJ60RMb8v2QVF/4tyDw49huziTM+PMrU5DQLqvc
BAkwVxmtDE5MbXwgZuqgXMn3YC6Kt1+jb7ld7sdBuhDTol02lGgxU40MkvbIjD9t
By/3rwA1ZQuKbw06Gmy9rvzYqoMdbnCKXTjJVNwxotfPzT61gP4TZFWqTm2oMY/R
+WzThEbKCiBbVr2Sw+a7GBRe644YOo64zMC/TTN+O62hAtHjyHZGCtHczmyyC8iS
HoWuXJ/YvOr4+2Nqr8skk0S+roKftCq4jajr3rCuvCGs0HpNnoZQXrfQ3j3dUekd
ttTy4X9fdZkRTOQqI0bOLWlJnrGm7JI/+RLCUq1ShJwHZ8t+GqTKc164HpZ//Omc
PTrzz2xi3qcs2koocDG6TcnXeYhtooi9wB4sxsenHxzbR5V+/zH4IqxcdJH5+Wvl
7Xq3+L8hyWBrpXv+v16GnVatIQjeI/xIv2chR9/VMrZq9IM/ZD+8FbLxyb/kRrVG
qTQHoyHIM+J6Hw+JDAlnIV5E8X/gI9f0QKeq6WUpkgJbyS4yGwdRFSlTb7t/dsPB
/cSRacdB+K09CD8huQp+ZWM5zjnkYZSPm42UgvfAvp8a56VAFWOVI8Po3JGvwTRM
V7NX2mlau1HTaDZ4M/gsLE1apaZW9lgKf33ug8j1zlfRXZVyZbd+mBq6FNuKInlu
8aMBIsa4BBmjD/6E/GoPHXrc9nvRn3kJEnaU6eT7mt3XQXfFvMWZSifrtk2HegsM
0UxCr1lNUIHHTaP/KbaFnfXB9grO0dM6c7rah31rFfI20W4wTg14Ay9SFf/nswLs
zRDuRTNtKSwzA+QCkZ2YcXiVISbQXCXDzCit8Hd5f5ZrYtCfaFZzD8xti9+ceEg4
+0whAJZTbRqkHDk+hIL+qqIJs3Vx6J81F+mOHxRAosXDDvXboUv7cT6i8YBs0+1l
MY6zrmAk1ZfJ3WI7MMfVEoM+olvDS1/lC9T4w77vNZDxv+z7X0GWEoWJgE+uAP2o
SIgHbSrm8jjcCKmR7c1gjJu5fVcPzDPhFtRnCOV29nKVXMt05o88133LTMabFOUI
BRJn6VyyefwfnCbxpWb028+eFXBgZX2IfYAbOgFOEvNP+zjqX+/082o7IJl3KbPC
6Fb48W6NsC/eblFUOJKpjltSmilpZbMPAbTtqIp2NVwL5AFVhqwSyfn9uCGaYcfo
WARuWA+6g4ZuVenHy8xhiElrdnBewoSNMGIDjgie5uyat7t2ra/q+PrAgJbIvnTW
ctHgNovg1srsMIyrtx2eeqL/fXhAHsgEy55VUZmseY994Mr+g8LlERvQ/yEPplNH
Cv6u7IyV6exlUBFKPcwszWKzga0t/Xo2Ham8iv6O0fXt81gS+dQTXeeA2OnXZ98H
oqK8JA1+jfxMsocLGO+BFVWveAvEnFMcwnYZsnPjBlPrDroNwfKnR3N/2keh3GCA
BXx32ewukvjDOHUCwMizdZ2olInB6XcI7vRC02Mj2q5V0Tshul+eUTg91c8WL8fr
B9mFoy8aWKaiiYfMlFKOc13ua/yshzZ7qTO/+FJUKT/0hyq1pwpF1tm/OLQ/QcrP
nWRrppebliKhqBAAetERjL0dZ0bWE7ZI8jWbAqK4xB2KwvBaNL5oGkMuoDIdO4Bf
z8svzYyA2UraKo2or4jVsiPK9yN+g6G3oOf6EbhqpadtLXNW7f/kqi4FTr4otQWO
G+FbaPOluKjTHw63/058OgBCd3vx4wd2on6OA57Sq96CJSn8OmaerDxzLdq8NOYk
FEUdBExUfFaM0AxmJUDXhmABKELgd6BUJ8mVIDpAqMgpaXJkkmsEhgfaXxaLZzVA
hzXxsN9GVs67qj3WGrF2ivLrs9tD0LEasOaeLrcpbjlGvvBTJTY5Eof6TdH1SE18
UILCK3PRHdssPPAWqqCYv1NZaG8hhBhjBLqG6Xzue1I8Dy8U3ACYtG+aK6geM+BZ
EhOyPvP98oVTWj8NKW4Z/TvNhPHoQxntJCmynXwN/fqMHWZEGzZIyLHgZb6+eK6d
n1eB89HfdYZ5l+j8t3PrS+HW/Zg683f/3ZeFZUkFjWm9oH/Zpe1t5VHQv0smsS+s
yRKE4+Rm4sJMWEIuZRleaVvSftks2xj3myZCCkpNjSNaevp1L9L8Siz5IaxzXzlD
kpmK5sZAcBlQ2k91OjOL4J1Qro//+mR4Gxp54FVa73uCw0TGzQaED7FMSKWrwc5e
ZIM8kxHxURt0fNCN5iGknwlcNPmssI6YcZkP+BhwMgkUyCV/Npx+65psB0Fafc/T
U6fbXTKgafrnrpsNBMSvN3fu5LR9vMxGrrw7+fDZ2VhkCx/5ZvCQKrG+QLdz7vhB
3WBcYHYw77aaeIK6TBXbpmXbQG2sz9AH9LC08VdFjWV8J9/9f65db7WKwyvZUriz
aLBEXLjQm8f9vcN2RhkV2MQT4Vmz2cGPRFc7m7OhKgMqUekf/+6dlgSmuNASBe7o
65r5SHHs9yeoTacC7R1Gnr5zZ5znyv0RJkp/LwozXd180mtAhSCui6iLqTz5TuPw
HjlUmCrQkeRZUZT8E7CaB+F/OaIVAN//kHvDbg5Ud3Ssjitmp5oipvLeZo80l0O5
nXT7U0BiXLWB/aonK3fw2WH/802mSu0ZyBR1JyAuveMoAtAEf3PqR14m95GruCKb
C7IrTiBmm7DPEa44QOk0AoNESt6sPs9OUOVqmFUPgJnvQrt6oHjyYAM8ouzRgZxC
HUVZ150PlJvdhNvumvZYJblIwE9q8APoK/G7JNnK8drWTCurC47QKx5P0qzcNGz3
S2uWe3yZNC0ZIdXCOrmElxVFdxza0dkQmRk0i0wMKHff3cQ2fDos5nTzQMH6Dum4
AW8MAA3KSwhP6WXzW+PGQJZKxBL02UyNo9ERQvzkGTpj1MC0qLUjGzj9PRjYFBlp
+jXyWfU9Kjm1r7VQIkWbHKq0o/D8bAdjMcNJvZitf2oLHBSgqwiVcJaTnE2ndVNN
1q15ncbdksG4e1MUFPmQD6+q6NgYD7gF8aprq5NdOznzhazF8ArV7prHj4xmA1Vt
FRT9pVjrwVxN+k+1ZeQHRXfRI/ivmy5qxokdjeaB7c9A3xHfSshpsXYpKJgupVhe
Y83K2Vo0bTGar83rGZJGFzx6nycNNjtfEnvmiEtrL4WfGfnyCME8iwctJOQ3u2kK
zV6Fk7KvfVSVkyXEPBF+0ZcXxclrJTm03Wrkkd8tjwLlbiWVuOoxiOHCzah9I5oX
vxt5awtO9UOMdKDUskIWTN2p4vS5D8ZtZ/0RiGHsqNz7wEllzKlehl1/0E9+HZ/f
dE9x41B7TJZkJLWt3itB3m5ADUNHbaXtjoJ4gjPXtpGOGNtUTVlRz5Ptqc/pr9wd
YmOk9+GbAkiUy2RmWN3tNF3AzOcXNeBn9ohsVVrVBR8220LLZ+/Y3FHx80b0Qb9f
ms7MalNkhw7R9z+6E+pEITHdskZXIrBQ+HSaO+/wAuigPuYGG39RLQnRjhbVvS2r
tTsG1uLBcPRZVHCBPP9j+kalsKdJjqt9hjcOPbXr2kfk7W1JpT4ULk6lWHMZoQ2b
t0h1Aoq4YwtpW+Daf6xQECmCVJE97db69rQ77IREpxbLG3UBp+ShMw6XUqOoTR6Y
rHxtPuzfL/SFp3NyMWa6Nr4zE3PXJukWXLl1mQTc6isO1tPLLh+TvzEJfZ5CB9QO
i17dd1V3ul2+/ED1r/mTwJZXo+dHDjfEsmyTFDGzeVe5vnwNIwZirxYCoFkT9gcI
PPzUEWHNxCRoI3Ck/mpiSs+Pra/rQKeITMAb6mKgHeRY/y1Hxfz4MinRQUWxxV7+
CKUCYX0M7FchIg0S00+Ic7X5Nwp5QGgFpe06wS+hf4Z7VYJUkMZg+ufQTmuttk6l
VPHJaIpCFGBAcyYqX7lpfwob9z1b40+i6rTX67G+gJDiDXTx1A+PQt2z7Hm2Xptv
wlm45vzCEmlQWUfys28Ahm5hO94jOSAdAj/M+xK8j5QOfjzC6Nm97sc2TtcLNxmp
gg7l9MT/aOX7ytI2matHLEWdJcqGKsfVDGoRsMvNqVf31UMF7gKuc6LVuSm30W94
IWTMV0LUN7IJMIqHoujbgDCHVa0nlcl5TxKxC1jNdiawsa5Q717Ws7B5WeVEwFbb
fmnWafMOPhu70Lb9gbIzdTgYVS1QrQz60KaSZMvO+W5r4Z5Osph1rymO3lYUhATt
fEu9xDCh+IC0ex57DjRXgeNfizF0I/kldIWgC97nAFhd39y9yfMFvYjdSSqB6gL8
qd0+D4o0qi9oMNWRBYf3QK+ZBs/2UTap4VsOYGsb5urzoMFcL/Pu6LdtvBqNpA+2
VD01nAg8NLgnZiFJvc+uEbTNyo9h9Gb4S5PIEONj0FFKNspBYeD5u3/N7TJgp2hG
ug583+uO2QsK6HDNdLVybabivXCV02jeNz+HTTZa9aUzYG4pA2k1QthXzj/iFw05
H2iZQYxKGDfcIfqFyColBoMIP0IEUVYZ5GsyvfY2WGyTa8LvY2GpPMegNdR2dxrA
96lThAyqtfOeM/9Gu4BjabwLN0OGj1QMc4Ik+Ii1zAlweNZdgZGvfEamjkbOPzeE
i6rta0ZTFm/xWHRkiWZmZ8iJAMpaKjNqPTkyOREqAYzMYv28qbOVmFWNovJgoatJ
3klcP2FgkEioPbkuCorxizL+HN5FSgX5/Lugl9sLJjzIYqSkMe2gjzAgdLYDRRUi
7llk0lxMmLD8/UAFWoYIyXEhfdCLdcAv8KoAkgEhaC8XW1xoyrCXUtkeLgGcbqCJ
WBfwosCu4qg3hkYwjOvpiOHt7DL88B8ahkkZ8JdtRDm4YHTXb5WnQ2Iv8cVli0Bh
duAmTmJ6Nrha5E5ysz42xehSAagD9AR+mk/lN6ILLQYJ3Bqm3YVmCGZSzSSyv66r
K9tlIwboHz+fTzzOdiOE6YCkKYcGzk0SV1tdTuHCOLz+oyYJE7Vy4FGTP/F9mF6T
5Dex7Htp290PB81Y10iCix9Nrv71V390bLJ1aQjMnGe8KE/JXeydcqbgrdlqDUmS
/ILl7K/E293b0t7gmRzCLMfiY/4jhnxR1TNbwovxfoohUGDn1nMtSjF7l0MJctNw
lnErFM9xFjXDCyEEWEVIhPkVr9UcgZSkJ/mOqkrfmFj9HsnowPC2fHn2Yb4Di2Wp
l41UqN3h0nAQ3qT4iKi339FvrY8BO1FlgvaFfeOejLEbvEfxO7fLERdmMH4gX4fc
TgkSxifQX/N4C8182Kry/5ioclPJM9TNLa2uGrndIwgx3OIbwZKU71tMObkEftS2
oas9uqclKlet4RaH1Nekp1iwC/btCZ+XFX6ABltbRecNczUTxHVrtPj1dQ8pQ32r
lY1VDYzzMHIaiAePPTrewor81wMa3KipS8+6368JlmwugaP+kwdAQSF30jx5eZLp
Gqdp00Wr1BpP8qShixJxRDMv7Y5pYIjQnmOzjnAty05KmDdRPdZn+7KjtS/QIhH5
rOAlUyJ0mhBBi7S6ljRfkIrXFGNgQ5U9/DHwK3ROsuTyc/0tU7hm+I6l7UrYPuQ+
acT8I0wigGdwZ6CBYgqbkZqF3rFSGOukKuHnWGICj1oaqC2ZCe2Kaf+C5Sb53LcW
+t7JG2FoKcNIFYRtn7P0JHl2cn5WhFQ3mWqXOTL8YoarTUvsodEtn9R//heCxFqB
lyWAcnX+hPH2j/fWqslFsvBDJQI3eWPfoqdIGlF8pBgGOFgV/NPBFzqrEvZL/3DV
5QIhCDVh/m+qkFHbHQng5XE29ofZf86xObTdc2X2enEcfGOaBoBahPYZjQ0Zg1m5
jS0uyTxd8yr5CPn4Wgg+eLePKkU9RfBmFu80Y8hgbl8FqvC9E27dV2gIF3FfSynB
OTit9PU1qPCJeAp9IBXxrPXkiQJyhib1f5EtWiT81rOli6yZDNeXN1/jGtT4EaSd
Rj94su8juf2qjpTDP0PZmonNwpmUNeBJbPcfXtMnaPeXUqqBkbOez1m9IIs0v60j
On0h91Jo9hrI7j2Rs60w4M8ZDdf7c0bVff2skXdiTggsJIc+uh+tmUYVV5u0B1WQ
ir3YL0G8M35O9s4Hlkr5b9rYqbMqrRi85qWIrJKtf1QpBJE5/sDB+6dI1qIkllCX
JouMRe3pRWfBfqMfF2lc6AAi71Rei0lW1VcqO5TXF8n3qhaktScB4eO8j6Kb1Azc
snhwCTUh7lTeAhVjIV48NVDu5hOujInAQJupHJuiA/XnlI+0XTAy0aNOPE8a9vWl
5DLI+1GiHx5pJYWawJbUN+eYopM/P9Nr4Od19qexPvF+QxRgw19vqMQwaZyJGogy
/B3mxsn34ioJlhw9Nb1li+RxPGVeI1TE2ptiSZRGtnGr8URDOjjFTAogf+8+TiQ5
KEc8g7xy6KrYJthqb5bCVZsgcpuEOdtOHSm9G/RV6AvjajdC3arR9NL9yFGEwpau
KFR5R92oWsFb5FI4YAsA27RViwSIIMJ7ktRdpPAu16eN3XVLTh2VPyWvXqVKjxBO
kCcN0+u83sk5V2gIb4zHpILIMMU73HBYiUtFqBhsfy7tP/41OAHCAzFu1TtS2k8P
cYaMo0e8ZnU7xQSOgo/QVEeXUST80PJcNgasuCynFc41n4wlC/MW8hM84SelaHgw
dzTiiygaZvyWBl61ErD/oojYkZaXtrVxzXh3fNaFV2TNGTuWw70SNnhuw9QWTaW1
Q5duipWKXjrSMo3kwPOToRW0YAcLZAhhqZIpyItASqvoSj84f1qfskRegZ8jDQnT
Pn6uWdWFgn8qEYVR986P42ZG9Z5EQLyvqw/qKPUnYw6reJnm/38R9VdJFQWhzYcS
Pc4WDeXIqFcFIvrJlDdxEzUxsoxajcMaihVJkowSgYgBMB2p4PXjNYk3VP0Gyhfu
bYCHRyQzBiZwxFm7iWVIhk74ZCNGG5+4JmACU6gds0Qrv8cmCCbCY0XEr0PrxgVx
7SpB0J88EznkEk6o9Z0BSwKi0mJGqfPHKhqIbIkDnOkF1IbQw0znAEe2N9FFrlIV
frwPbvjUHNTFmtqgt8cfBY8xhESw34QNKCp1dy8RN2uV4Suok9HbV71G+KCpwdXM
XU8sfrRr/9wmKsH5TzS00WEnLHRK2sVM+14XfaFcULIdwCTg1Wiln2o02j7SmlIl
1Nqpc7THz3zsdHKdQcvnoquwKtlFi5YXoF2R6sXhPgbiTCv67DrtN32iS4vQyIT/
JJbYBhdLobSjtIOMQxGcim4GpgED3sBT5aVZmOleF0eYMgx0LLvhva94USyzy1ak
2yrtbydEymNpbN36ZL2Lxh8UtWLlRqk+gEBs5Y0uTVJy67ObY6MNJhI/4CbIgp/t
H9xv2raWeDwBiQnhEk3U4EkvYm/POyXpVDe9Os0u4xrzcpNpTJDfoW/ymXknzvI1
mFvWtNTbo0v+pOVKB3zQg4wBXkBGLWhtfiYbRVy5tUy0wQ2rxqqoVGV2zx261xLM
YcJznKorvIoGrAp1hjPxBx58mpZOuZiQQDE2Kiobd9KFd73uvL22vzliNqaFN+7I
UMe/wFVZ3Jg8DKvdGAlyUqE5b9QVdIBsFDyHbNQU0AfrhaeMdf47vnYW0BXg3S+P
L8m8bfULZGYejHCVTjRZXLV066zbvE+F+MxsJwRN6BRcjQGkXcxEogJoBBKcKPmn
5VxAaKJLuD0lhwsYjSSLdzIRBREjQ7bocwb0HaWL/XV/RmIlZi+M7eQR9mLFuBw2
zMmcU3Xk70SDVVL6ZiK4U3bPxtBtas5Fnsg20GiP984D1d8MHPapXBaI86ivt/ch
Aap505nHzeqUhb9GB38MAVdcKe5fcU8iZfetsL+FPiMwUx/xqHzME/nipjVEzp1V
PbSb/7QcPTMimwL8Q7nhPGGA6JI/1mzEdOOQzxt1btmLUWqpuvCT4Yjd1hJ11agO
dHi/IP+aVYYzH20z2a/YPOlxLsR7zkwWoQ93K5/hygzg1r/YNvEo9Qfktp65HWMl
N9aPS5gpElIMwB7upsMRzIWMDzDDigDPge3bW0R+cCUWMRRrgiz1nW/6d4iw5WJ7
MUmn6tFldaYQ0rZcYs8FgyRb5vTR6hAlUAAnStV64fKokt6IBTjFY8KxWt/7lEws
fYg5G8JOx3G7k1vPb/yj1jjQPsxzCe3l2UhV4J8D4L+8BJG4gjx6u6JJGI/pu7Zf
UZGe+OD/sidAnv7eUXe1adoDYJwfJldZuNd43mJ11lCwWUt2yxunB+xpHtxSapbS
Gg80B6fp2S76RP9cFGtDq1hDVHvzeG5P5jhhg/xs+jGBgtX9gog9bpwzb5NxbBJ1
gH1bYB4DWyjgGS8QFVgWs+CyKrLjvTsiFZoZGY6R1CrDvue2jWD1WGel5UZB1uB6
+qCmXVhS/13BqKJvsltPE5HzenFRrUHpd0tyPzVUjCA0LDKqgVyFV7YBu1F9juY0
hlgjs7Tpe0PGTiybfpy4C7nU3eHuazfRbOKVTq3+a+dSy+p/gacbRu75ZNBBsWEl
WS6KnW1dsTcd45WwaxPyS5q2tEavaDhsLN/0aVizWQWNfxQTlGgXyyReBs8qx5Wm
EEtvuzTWSXjBMo9JwvcwbClPpHfc6p/1kf7bNcgGMTr3shhRPUevZurop6Qmssrg
nh5NDm+j6qaLSBm9rCTz+ORWxJu7Y+U74FC/qkHrcX8CObQc0jmzzackKOFmJ5Mk
1pMJAUfz5b9eYD8kZlU54/F73JugY7pceUCgPMxDu8A4escQtN7J1QdAgd5hvaSZ
SXzwVDRk6JkNvlaITRNXkixg3JKpWsKD1n4zY8TSVbaPfp777WMTNehj0UWxSOt6
voO7jP9CFIbuZ6C56PYn+j+No+kzLjDNpAdEW5pCjjuT8Z8J0HryYMgBroqxejGv
1gaf9YEGQo7qbcAT6Fxiz3lANSk48XmOMmzVfWn9TpSn/6Ntq3/ZrdQib6wyNlcw
anSoByFutLqwnFQwmZlAoiznWvzcaYoZw4QFlgJTPGHjATHmrMA7BFOlPGFdq+th
IFJTaT8Lw2WANjs32kvwyujjQyucceHgquyM5W8bHbZp/7LZErwbunOKIVIvb7+1
Y9sgt5f84MBxoAnHTUacCvLzlUN45Ucyt4pxLY3NUpUntkmrs244Nekn1hMX0bxY
ZnBDZlW2uL0Ly06EQ5vS0CkBFn1glu9QWfASCjT2GQSLkP0usJC+LWLjJeGyZn51
gRVksRK9yEjIZodcd+SEVNf6e0Xp5lxQkL5nbisAKnwbHtOnFwb2iTKQ/UASf9O8
Af9fxd0xzHJcjz8kqLgpsaZXbEnfQ7If11kv6SqSQaSvIZ2nwcLmy9qKRXHMyKPi
8HC982KDz28613WaGfVzIskZafg9L5IOb37iDdg69jp8hs8+sHxJ/fLH5N1hThj/
Mic5pdKANirxkDA4E0X9uH9ur586BxukmmWJo2L47p//T1knD7BIvdnEx/gPrssz
r9zwRnqys6Lpn7LJNtODWbxy9EINZMwauHGxjpI9CwX8QcDHEMqoHd3ECSPSZXUi
Sy+//DlWz/R8Ccam35Qor0P3ehFEQ+uTUv5e8O5HTDAh+g+zlzV8ZyE82nPAVDD4
0R1KacvdDggSJSVs4q8AAKs4GObf2rQEs615phZ5EtyuS+dR+dbVTf4aok5nxQ+Y
tJwkYchugZXAO6AmUOfh830EQtCb653R/iWta8zK+kyEbt/r8+k3Kc/UyRbuq2xN
SVBF29SwDrGIDVa4HtLyyd1DVFgk1dSaMTwFxr98JlJJpHBV0yv/ijvoZY4bZGtD
KOpaKCvA6My8SBJ6l5GtY6TAQP4KzKcZKkIWcxpSJkjtyWDXcwQc96m5vz5a4N5G
x1V8w4jeVDjiHr6TEVtsbV6ZZqILJvllpe+RdhIXU6Bi52RhsvMopEY8KDIxOq02
CmGfOhlYibMQiuwStVs7K1SfQUsEyq7OuJRchJ6qzbzMw1o1CsWW3HGtVakGGZvJ
j5VTYyCQZhQ/CBRyeDIpSRtScjbYkx8/cuZqnRQyW43Aorspp2dElOF63cjp1kwv
fs258xns/kZhxOoT+PN9UCVeOs2mQnmRG00EevBBOWBigU/DypfjEdiXVIbU2qfO
1tfKZ2PCuZNo7ntKsolKXwWq5bW/IbFdrui7KpHvb8jAmDYe0b1CZVLkOkGyFuFM
T6jrQCjiqlqyse5074EUCCqPMdXRkziatZi5QTOikuPVVxLfR4ebKIGERxHhGnt4
bL9F3Krj2JD/T/XfEaOqMe6X2ECIIDFNtR4AKprZf6UVxSMB1zbE+Vx85Dx4Sl8d
Dxx3dYqY7PDB8mbfeJjcQ2gC2murANHf+nnard+RjtwiuYL8tXbSOO3i9nyIx0Rk
PnLrtqoo0eysWe6yFdtMaSegAyBRLhNSoebvzVukxBZ3AsCc86eLv5pALgcxn9kG
52vx7GXc/aRLA+wCxB298gdFQmN17nZdVxXe09Q4VyWmofFBnrGBCA2ReW/0ewym
iRvedk2Byfedmi1/Cc8h/C/y44qW4DnoqTQn0WNQDSjUVXSwxkB3J+QCoH956X+f
r1AgicBY22u9A1BGeMjMzvmoDPZ6gyMZZMzyBKtWWdXpvGUPo8y81Q0tLepyc0K9
2ZgSnMqQBFtptHWGzvTS4E6nhN+KdQA41HmuEetKRAPg8iCzFcqze/48ykJtXYuB
x3iwU9xFfffkHpuH3f2RcdYNUdRuFTwfnpR6GnwRKvs3x4y1pOFTASUT5wSk8H1v
THd4pYfojXHjY7rk9QPQOaW2/ueMPhxngv/o9L2zc6lHc1eYw+USBDwircOdf15S
JcoKJzjgM2+aNs5xekCSKIJ8kFGhTfZ/i3RKj6Fy6v11sXx0k9Af66u44I9PiwZ0
/dzAfPP3Kkxa4V+YV7Q3FdJy2dCzd1iL+4IWdKO2Lnd6f3I2TgvaqTU0uyAjjdlY
KsXtYX25izAahvK8giJQ5O3h7dt05eqYg7a3kOoDViTKCbZv0dvCd9XeYfdBZ/HC
buY1q76ZCy7NfVbSpDXjo52qRGACT0pK+lwQVWzfJ4STtgTY6Wc7bPhgUTYVA6jk
4vsvmXK1Cqdksuk0kfuS6ap9nICPRnqb6mE7VNfkWI7/XfzSwT77o5n+jaJB8oDH
HqcVrJ+NjPchhB0tmYQTSpeBwedFlthrRv6t3+RX2l3Fx7R6oICD/LH1jkKPwk+e
OsvmaJULzfXnNN2NSHlZOwhUUBNSr/EAEI4dsRiGYIdQMo9Sx9+0WBD7t/Bkflhq
KjPh89dhed0onGXDZvYsDCLsbX0KXDd+lCeK4/QYxDVCm7LamwWeZsHF9KBppU65
I7Cl//ykGRn/h/zb7hS05RDfZujSXC6jU2Ijd53wfY+Jg1KT9sK1rSRauFVATV2S
EexSc9Ie2w1e4izHMppFyNgUyOQiQi0BGUz6ezQ3xqiXapYBWpwWbqi+TZoseuRR
ar0lJo/Cq5m75hI2giGHEtmsmCH8l1XMC7S5a93S49HDjcQtdW6LraXXokGdc1oD
E2M8iff3HF6yILHRmDRvS31iE4HqmnIyZisBY7apF7LkjHK86HDbsoV40/nKwJAc
Dw0424N9vyep6EwUXAzMdPAKedud2wCMdeA9549rnRax0xvdpRrPwq6NASxZH20f
mhg1yP28D4p5t8iCPttEONZHYSuaQnxEECjMXuqAKSqBoD/M0MFazf4YaLLTj6Mz
EsYYxLOhZd+OymfCzUwcmlL+mujk/PchQ24gszTfrMKeQkZpnyUR5VUQGPxBomZz
esKQjPR3VSZRThG+lImDWWWg9OC1m07PcmerreqVCO/HJC4m93fX/1tU1MFOYscA
SamZ2Yz3y4W9odlkhk1jHE8PlOu3ukT+jW2P+cgyUD9vvtpth9pt/uAZRCrhWvqP
320LKB6Dlrh5BBiiPpdxl0D27tGWxg3yUlVa1lLlGx961hDugEidLcI6Eve2t+99
1QseKHaOVcsEKkwFRjZxb07ofk6eahc/+W16fZLMeaWmLgfLAEBZSYD6I7djZGUT
ElngiADi1g/AqfeL1SpbAVgr4kmbvqlTgI9bDup2aIFStTTa0jUK61Qw0jUwfkJg
JDxlGjhw2eN9oW3Yzn8xlbb7+YCzpSw1q1G0Zp2JQ006zGIgEgrkXZDazc++PcKj
nJ6lTJTVBLEXH0qYEPOsJ3GoZW/Mhe2pEYCoHqWwZA1z28mKclkuZTqSZisjpQpo
w3qwcaUb8BGjvUCYLC38okaFo6GDYax+d9OkY/0wCrbGoXp3e/uV8c71bqUi5mUt
8FGrmg4rswOvyo9pyCaRiw0U2bJx7ETChyHxaPRTYb+cVmzQJD9bK5ghaZjbSnvC
aOoaAJFIacJdpkbnLP+iJroOqSO71Wld0Q5nL6VAP5rasy0FTN1rVtP5GVgbpd1m
5LPVgkwWX1/2gX19OYU5LUcxt2eLV/7dO+pXiGcLHGNS72WYRwdJvDo+bN0P8mJn
mfChLvNw1Z44sq98bh0vx9VSFy8gydY3c9nK8I+36W6TKt5hNDnW1A9F6To0Khlh
j//NZ/J1sxYJB38eS0y0j0amWu1Cp2+T5Ir2OYE5sNxxbXXKjR6IkrcbxwDBdeEe
jD5gVVdUPi4QFWXRERhvQdBvdoqAsCCN1NXmUql8wqFwDpWzdksP9QERHN5nKWXX
roj6OvqBrtTa96RW6twlPhQw/6H163DLTnUJo6q7Jj5NTwGclC9Ti04rd/pxNBv+
cCAoJgQ10jFwdiz4aYoDXh6XZeutrROzIz4UqnR+d/flgoq2E0HIillZW3mnfFIh
jdqtXgdLs5lkCjGxggjYMLXJB/SjkJxuRV0ZH31oCyip48p2CwoUxqHT7ACPhyFx
WAwp9cY9oeHX/S8/fBjUUwdJn6SBreHzVcfhNJEuSeuPlUt0akUlYwczqd0G/P9v
sIQ4LCG9Ckw47TT3efZtT8or45YWdSVbqj9otkNQ22fSJVh5TijVslUS2kNP6RRt
XWOzLHlZLi+GALCxGln9ydmqxoCDbyDQlA5BxVCbuzDy0KXDwSbUr4d6IfvEeSjW
9N3po7IzPso8Xby5/SV0d8YCEcz8SVXf6lQJvXDdoYvy9nNuVZ5yamMBw3WiBqgC
YbXk+p4BbPdHCfhROKpdToQQa+WUclJSKGLVpEIN0vdsG4+ikGn2hI/TesufoxYn
FV0g5OxqyjNAbVvBb6QWTP1dxoQWKtN7Gc4BUlsbu2XfAcCpRCzU+lkLExED5/c6
WfwrZsiwVO5bmN8KR5RNZzhE6m7Z283V2hV2IYW1pXXz0hALNK8kDyPnIe6/sgSJ
cjBmpVKuqzSkIHbQzKZ745m+LFME5bqadJa015kX7qyRS+k7keBbbQvLwkadS2BD
stlF87AjTcKzSpzVvXPA0v+97bERNXYP62XJS6XLzEXABKTEjGvjHl93j8HQlSjf
4efRFayG2T9Qe12Ut+chfsjeglod8srp0BtWecbKNFT4PIczXHta1j7bIBGyBnKn
DriPOAvmfUvnaUmdBz4WziOZ0PwzoB/vHWeQA6XrgOyFbF9iArr/VYNbe85zyr/g
bJJIDoBtL9aupALJiDG8ssPydGiLwFZA5wHwJmxPXmav5hxcd2f2I0vAfP97I1fR
dOB6QWxBfbfwdbUplgUHIlZsr9eTm7j+lfj83+JGZ/kT/XKaCDaHeU48wJ4ljXL+
PCvkTC6DlIRuOM+J9Yacq/NsQzNVu9YW5j/gDUg1vneOmm3YesKn9Os1VKfSXdSB
Y7X/wXh27v8lYIBPwEmbHvCZRQ6yrACSdiN7PAlD+D4VQOWgY69jRWVftX4ZEMr4
KMDjDybJGRWzPUXPF/EPY+KPn8Zk5lmrzhgxVlpxs0xnLKMB3SO7rD6m2R8NmiIr
do9zyB/szlyopG2hotTQKXclPjZ2zb+eEnBZeNCc1qlX80GN7nVAR42ZozswIHbl
PeipFr7VsNXggickEYbOgaI36szl6t+czHBa22L9UQ/NkgMhK8Om1xfI9AAwHsaU
EoWJg5S7EPwJIVsjg5bfIlKEyDYrCjdkKf3zXB+milsrzyK66MUj0CTwlxqy2N/K
dCw+tvIg+DpPEJO9xP2uQbwyelD7+svnhuPO3M15Tx+PZY1MYMCSBIuGgkF+4OC+
7yAS3fkLunuAQpzfqCNH4wR/91V2yEiVLGvyErAiehNeJ85WCgWrjo50Md7BaQd1
hqSx9K0VzaE6q4aRfvmjJ+UWoUezJPwC9PG8lgIsL4hBQasSpRqNwzfiqp062J3h
nLloM5Xj7qDiqnQNEnll6UdIGemUwSag91AkUinfZZBZAnlJ8XNG9PIFquTedF66
l9pH/SgFZq5e1HbZ0uCgyVn81/JtVds19nmAPNVCwPA0qjiprqHTcPRXPVuadqJC
IDQPpEBjnXF8stZb03YkDqL/+BHeNGF/X+EvXTDq1/PuUghs/q639tAqOvJYhbFz
JIgp28AvqSX6IPRtm3qNojqtym7vTHFt8C9e3nLoPbIAoXaTLI0tPZBH5S3p8wzj
X+ai+1kU/QIWXfUYirxmkx9l6jhO/bOEmAAWyr4Bcs3t/sNkMmD2x+mIt8+Sc6Dz
RJfSq/CAfex29k6rNV1A3IZ31WwsJPI+zXSvqOfEyLe3ZedyzEntvcQwlDHHkxKl
1HJ4ibzgJ7jEAqIOY8Noca6PacbH+mIq7LoaIY9AlA2iT/BWmvSd7PYcbtSpDuvv
PB3cp/+Pp3q2/PhiL1WsyyC0LVVZbZK5/wuQuvK29uJsNzvRB+rz/MqTA+dIlrST
8gvRyfO3au6eCjj0sHBvQZRai7GyjyFR7Ty3uDR8qjtGr9m+MLAlwr4r93ozajPe
pC9shvQD86C94tWUpiY9UgbIkTKhLASJGJnLY2+d/qgPNGuBPdhoALv1dNnOb57X
nS3EnrWzqS267+BLfHyRiFg9jpDAVxaZP0gPwI0vI7hvhLIOAAJFgZWaM+K1upmo
I2N5ysTcD6Zj1CnGStOGwR4ZltD0AsNAyLpZW+urmTtWkWED93NfbLnRnzV1Ir0M
JTtdsRj7k15uTz9ZnbTFoPozITSSD26xw/MvLWPYlVb7AiD1zq8YONT94wnz2Qhr
ip6k5gd6I0mqD9ruxLaSzwX0RKHHzUmPI6L144s82vH9gIsA+og5yf0jsppYzj2Q
e+dK9lcpHeiASbde8H70xQYb/kALS7TF2+8uhf1rJok4+G2nJ0zxuIyv/NjXPze6
xukPw8g1Yzg0ZAxvZv679/ueJ8axgKvm0dfI7IlXzDp4hiVe/UQPYkqmH+FZRNvH
+66HR60PZwz1Telg6XRcDE6bTWUjf1hErGuPtFe+yVnsSlek2+JPywzvOYIipCJh
/IcnFQbJkIZLoWd6RAFXanemp2UhSkvxylJQEER381jrC8w++s/3Ua23sz8IvLtu
wZ6rec5f2fygBKJt82bQ+e5KkIlAQoU7x/GalbiXS6FRElwtWNbIGGCoVF8MV3ts
LnzfbGQ+He80+5eZPquVPO6GnLBDuALi0jFjyjYltL/wyn8ei94d1zD9cZIuybXX
XqSvnlglQ1hPMaetQ5Bd4QngdYHhuvE5UEqo+wCCObEGAtztgsTvcBz5cKzcKRpD
zowje+RTjS0UjMdxtIRmtCzgS+eoD0WCfIvwfcWr2jbNWYb3mGextFBaDyayOt4D
0/8MxBXlPxFhNe/6FPwzcldpC9XtJdcNUyqo8Wzro1kLr8rIAtXl7hOAvnbU9qS5
jBEso3QuicnBy7sV9kWptXeiDCetkvcdkVYwY6ha/eObtEsieeleWjiTTb6WxAdQ
oFOo5lR5KFKUo9D0iEsHoRWRLOWlk+pINT5e6kY6N57jGT7X5ClCegTpGiVCzl2/
i+wuFoaO8lm8dzpC1CFpbWZaeLohP2wXaMcu2pHvdTgc7Bdg5CgRz+BqZTa4DRgw
HrmSQMKNwUCZJAbnh1Rj7mvvNjZR5H3ieT5E7eTB4p5P0+qSYTu9lEX+yjX8kZuZ
1sm7yuQb3O0EgxImZOcn+ahl2vxvtsvI2mU/HSDTsVKrae7j/M7F1GHZ/ad1ACBs
eVLB8RPSve3RMsdq3UgTGvtFkUR7cy0AAHAbDNR/2PN7QJJqadI8VSH/IQaD+28t
VU2K3VITYcInJsG4Lv0QgvzLWTVFgYKXdMz5bdnTmWx1o0AyizIYxxDzjssE/pDK
YVXhd0MjxZEhQPZUiMpqUYGgs1+txIDK7DlZPN1PeSnDcsqLwTd+KnFk5yCaAdbu
NlCz9+uU5UZw4/COhpTk5wxVjOlXRzFzAC7X2VCJUGfl4hkOwDd/l004rIKvTRri
AwWf9zH4FpLLOGEZki28NLRoI0poWEUVMT11CSU5Ahcg7EorKilk7PgzvG0U12vv
Ef1Mt3oE8WZfOS87uNnyKt+iFKc2wB26fEHEnpAvEi2SHCl1Q5XAa4SmmpMtI+MY
Y/97AFf2CM1RQfO5omVNnEsfx9iVXIngLyg14agI2VclqLp0Bf9TWViSWA/djIdh
v4+H2K4RfBfCWlHzKFY0MRE68y07SI7UoANuhEYttXentI+5S0zcw1EBhJrjNYFX
9c/p4B1toegpUB0q4hmDy0UB2qFi1mqApdPYoGdmRwMdZ7k7OGddub2qkeJcVcJ1
NbQRdMRXNQWTEE5EHn6d2fL3qTJL2k+Xo8QSrwdU1JBj2uhXyTkPdyCqoyEII3wI
yLiPLGtpVDuPJkBwg/Gd28XpQqZ+xnUt1FTeGutSqKUvGAUS9CuzxfgrrVhIABWV
07vtaRDjTulX4al1NdRCRCGF7knkEzO4kb/yS8bTnW69Pxzy3B4bbKM9Nb5nMa/y
fJeXgcfOCafGpEDOWw5HQr/umsJiN/T4cr0ef9NVcuW6gtGHNaHfc+gUSGq8Deqf
snLp18AZ7y7k7wSWljyPdWqfT1JeOInKQu8ylCkE0G6EzYWqnSC8okg1nRyc/alY
r5AlvL+Av5qTntfPd7ABES5u1MZTMbLdfEI8XuzjLurgA8dZXoG13TQ2M14urfqH
pLdfXDW+zeUPxDRKregqDUMb9hrmTpnJqTIdeY+TJw+Jc9Lr2Qd433yL3Moz7j3v
cLEUiVvrhaHN2HgK3usOkHyI3rQrhLD2glCOOxYLtGLkVtPxW1I0wn/NEdZX+vYQ
zi0VdRTgpW5LOHp4CPUUYR30bl1GjHLPJK7NIRCcOXRWO6WKISP6VDkyeOpbXZW2
zVUvCLcl/UMFFnaQa90WdmpamcR51HmDm9QwO2vWwbG84BXs0ZzTKX3LcHT1PTyM
r5z0KArOUrnin/KXC7mP0O5+7yZJnudgFanlmJv4Ds81tNe6rmddz0xiQrbFdHUy
y71xXqNhPuhhj8CupmiUnZQoIEKXlYVTeIfV3YMqvfpGz6fuB1JILJBmxo3NdDv5
fDlKnBRfgnQjnXklHhIZjsBtK3dKUAwZ8NQt9GE8XsOW/PfG6N7edKKshlyik8cY
3ykjaE8XjTNd/UbQX/JzLhPPrb0qa1qvF43AFEkUVOhZlCECXnsr1VFcZddIqb8d
MGpWIDf6Xg6AZgAugl7kiakAwC/e3BuvQJTkdiq3aN/oyzQqjXnEl1kRKFaWcdFi
EilBAqGoDSywWCfRYdXQXRVZDEGTXLagFsGGWHxsTB6M0BcgleoNgnX9f+OYMBFR
0DcSSH8iG3Fb0J66AiPFqbmnMb+KKIU59L+PJgS4vJqEYg3VFG5RbAHgmSsaG7LH
c/1ibQxFgzJxRW6ncPQpRTQPhS2ZpUoSmz3O4NGWST1lb3TOs6ZYbpspqor1xf3S
hLlMW+fS9qNO8abnrbyhzICWalIJyWHME7FQDORwMI/HqC99If4azCOZCKn1w/qA
jAoItYFbGv8Z4NBdxVxh1KAxeEiYBKiLVj62UuhGnwVZMqknWuHwlZcWgWHvVUhx
HIc5J+Yx/ZnWBNjYVy9F5YOdOQ2mlZWZXv6thgHmVG3aXuCvUvgxpsl48lXvV89I
2cN7n1Pk9HOPsRXPYRlum5kqqmWBkx/UAE8ehzOsITggh5w5nl6RrjX5h40/AF70
SlDes8HYpIceqW6MhwEeoWoVYJETN0pabhkw5qvNh4BWtPKD+5JihRpR9lZfk9J5
9AdgctYpL7mQv0/TcmcnrRF4ZDfTAW8S5wOY1s+Umcl0FiEazGZt3rnZRrY3VtF+
40Tv1JLRu60tOJfTGCEKIq9mUrO/pPNDw5eb3s6s9rQjj2KTQAllUTpN6x7SZqBK
+etue7EKNUKgF99P41Up7TinU9DdNwrY9M6eq7pY5W0Owll+e5XUV7XIpy1VB4hd
gJ/rGf9DyaZRursYvGaBjQ6UER5knmFoTfHcOVuC+GtPiQ5BcZPSe6zcFlx6iLox
K1J+Aeg0tFwK314stuoTX/wz0zaRZcCkbSRfBb3MgnDkt/mzLyDeV8nYd5ofBbz9
m4DXIFQB+dnxFHj6kEwIYiebrLXJF7sK+ukloqmK44Hh7e9I5RXwAmgI9Mcwb7HY
ER4fTYg17O4cN8/iaFHuHZ187Ke1PY4bTKvIhcyBQKkt5UDhY/lw6ggZCcKg/zj8
PsH1MD3vo+RQ3HQ9SVxeHjsIF/mAFximnQw6zbHBQ89YCOqG98Q4+e89ARFpyLuN
N9TeY1eGLeMGId/A6lcRVCMZcwvMKJOReEZHlbXOvu8UHK9rUOfCvAKRgkRZRtaa
Jsqtg5yQB6R22oPr/GH6uKpbRwdunggDeeVwyQfLO7KgAV+R34uLVTeLr8JYAwcB
dL7dYHME73UqNpgUmZmrnpoRii2yF9/aVrv5lDn0Q9GJGchqHfMTXXn29j4FvpZ2
dyweaAcqv7jx2wJCZur6uXCOpRtr5KdkbLJyvzcwyrVs0Pknsk4O75fyoga3dpxX
BUcReXT9ybyTvk2aO/r/HI/1Yju78Lu3i93g3DbKvmMF81B7/TUqMQYVkFXv88sZ
LcXvspo+pU6TaV/JsfywYs7RpmaUh3o3T7S3uD6cuJzw164fAHColJGeapNkZm1m
yymQsqSlRUKHmgIH9FQjPixo1rhlmqxDz00BbS3KgF32+igYq6nVAM5x9wE4bPrP
usyRAU7q6igkZjVQ/Fac4BuBXsB5yPMpwFics500UKX67Fu4MfLWcD37BaBwIykD
omqgXOMIauijAYkXl3RIFnyrURbewNut8rZGyw/tPeOvs1gF0EWkYnnRo7ecDm3V
7LirnSbTUCJ2qwWxavs9ieHexalYYSf95luZKXUaINjOBu+3mGIT81MZgFqru6EK
cFzRheQRQKnHi/ciVlWdscMpK460CSyj2M/lkSLqFxw6sTCaAvKPs4zCbn3bH+ff
5bpXXGJNVlY7QOVtzfCJU5W7E38lJFzDXL0IvEkta/tOH36bsBxYfYoV/q8LAC0Z
MZSlG6Y5De0/W9afuVPjwSCiNA4K9w0hdTeeiGcJ+eryVOU2jy1Yqc37EOezSr2x
sIz5qk3nVu7RHfyuf1XWM4iXWWojTi/kIii+E4/RzU/C75jPzbPlrmpEJBzOOwOM
ZG0mNeIyDwgv5giuPR2Xrt03+SRuiBuHp2NoXmszD8YTQEuFbtuzequlYvvag3xa
6P7txS9X81QSWcqDrj0Kt7D2sBgRnnof5GRUZq2fQith9sDxYTHdvnRwcSzvOrYQ
lUGWfodhHJCUbyT2nygaTgIRImfwNRDhF9gxpdvIND0ZoQ6pTY7CjR+f42LPZCNl
4FW0VlBycRDLcogRXgZml0e17KiyRefpU7HsDnud2gSy2rGZjtk9SqBbwsrcj/EU
VGbH5YrS2GdvsaaKH9PBs129PhAvYUOIWpWF6rSthUeGgBBCtiusidtRZRLPjKiC
jrcAVfgyhCI+vR+dWmAYOO5wkD3Ype2nTT8V0hwH/guJcQu/fwSzMfsanFc2n8MB
8OOT+x3/Ah+psE6tDZXRaQVglhZ3nxp21Z77jsaSauDgNhsTGu/EuyEFLbGBD2h1
n/v2nP0kY5WMgxC+6msSewK48DjiuBbOjPafna8vWAQs2+jd1PqIvvsXpnMgmlau
4YADuQ+rxBwDLw5dZP9urNb6SgjK7eG8wrwieprSVfpQEB6Uz5ruJoV/bKKSpwO+
wJmY2ikPipjGMJHbGj+5nc9ouPPj9VUI+BV8dhmTlOkIcgGpNVjacJKvySMG8tOI
oARag/F7MNsJpha+TdIiB1AUfIdyopDBPd7zaMDcmn5iXkPKNdM6hVpvP5iys404
VA3l5J5s4rkrE2vLVF9RtcuIFWz4BWQdVCM/HgV9S1PrABpDdIAqfNFipeWxW2+T
sj55SAeKRdUCdQz1K1ped8HYxHUGVYQAnIxVZl2oLwZRqfm2IEkdC0DeNOHAseS4
6Jhazu+H8EOZS2OrmjEL+cbYW2DsTzv0o0mbBIy61Ubclp909f6EMc19zmbTYyF1
hGUcj9Ln8YSBSHU5uKOBUWZ5udg9CxHK4hfmw35LLvFxfP5tNBuKpP3UDPLZl1ST
qLEqHfxuUO1/HnSdtZJZlxAWYtecvv/Xx9SVEWonvcLGiVDvTaTXetIfNetNUCBP
Z7w5DOtrvchxWTBGzOhVKUDiNMNyIGNtVckPhlx7XfoXRw6uyRUaxZ2M2f1Qcr3w
bvXnJ2jCNjXYU1cxSwxtsJESz2l9IrEurDHqpX2uSNL64OrB4WxBI47Zy22L7Vua
Cm4aVcB0PgJfn/7+ffZlr4JTeMO0KOtmY43NTUBLKveQSYycmuNHxW73tFY9+5Nn
GdlGUrGOOCFznV10WO9xYFtIfrEM5dm8v/xHfD01Jlp1o0+E6n94Bw67UQ0EeV0s
nVg1CO1qVH9M9i/8tYJCDP38hgUpGHhG++XLo4Y4mG0rhkWdLjzyqdXkwI7pmTen
/AqaV0tra2EwEoDyilluTacgx7lSSFgcin3iMqe+yKMBvIA/TXow5qxM1dtrZ3EE
ZOpOIy4/yPmXt+Gc2a63KpCi8XXtLj/ln6qtA8Wk/zefcD9SM21CWqYf93/BCbAp
M3F7/Nap/YH8vavReDPrNRm1Rdmx3WnTSW3+IhZHSsjnScy/H7TzphyUSsJbUYkx
yTwFgohvPZIKdk6RQ2uhW4YhdyiaBGwvQT03qlNKAfdZPqoGAIwZ/F5mggDdR6bY
o4PP7+caSpfVe6hJgIG5b273muehCpv/SU9SOhY1NhHfe4VKNLdpI4rF2GppKrr1
ccVTfQwqWXLMUFWQsATB12enr2/svXWHAxWW3+DvtP34WfuNrb8LcQZzxWcMCHMg
cq4MZEA8Evly3XCmVT5Od+1FnqQ+ASx7taoajduPIW3tMN2xdLMTsFGSm+12vTJZ
6y6SaVuzbYeakapuHrVI5dYg/0ypwgFunouUhzSNzM5SnCs0wHGtfFuDyFy/uH4L
SEw2XL5U+V0C6NqE5gaNbcwc52TcS+7HQ3XnaxpJzggDgMNEJgDP0bpzxFLYYxF/
MnxX1iUt0KCIXg9HUoXo7h4oUSt3f5FQMsPayj7hIQB+QwS2FYzmZkwUbGMYnFRx
YziFykFtPTKmM3zP1KQaa3QYrGkdcxTZsNqbekxxQiIo1aEiWoqVkHMdHL60gJWb
PP/FVw70dgwy6fTj/HehT+Ej6tzVGa5IAXBNxCLop2MmbEcam+YnPQfAXFb6ZKmK
R1kJsCrHSyHGvS1EfeNyb54+Pd2IszIqcgsJlhnwTmMRq0pRzYGmvBb6AmqG00Hw
VFVTVtUSr1lAJbqzr4TlvysqBnrk2goZKJxXPa9yJZQyd6rfv2qc+t4AlAMmTIve
QQ8K15th53qxp801ht1f8HHFEd6NpekJg/xko2oe9YzUEz25vNOf5GdFnxGmcWAa
aLcA29vjckCCSZKid0qSsM7HyWvQcc5aQuDe62tSurrXSYleJQFabpZgJoGmcBnx
0kCeNk/E+eZEJvQ5cvmZdihifu62cwMrJK9GF8NwVik+y223bC6QvXKpbVC81kym
53Tbu1EOrEVnyiusLOenjW7k7LP1o8PRzgrr6VaDVMjVGmgSkUIScJNk7lGZ5vZB
jwIf1ZB1CnXAvKhkjapyKC23bnB635P+UMJ15uARJjJg5gCgErc4ZeBU+p1/JDcz
uWRjdpDuslc7wzVkMfSRBABpYytRrfCeqk9dkHZjhtrwApDKrSnJ5O5hVts200Wn
b6I4XyjiwRpmoN3Clb1P3mhnv8N7p5chMoQuIphGFZQXM1wYfSY7Deb9u+YbPf8e
CZLk6mK30GJAv8z2eBsubAAhpH3zfCyA0XceTa5DBxZ2OJhOXI0k/Ep6oc61lT77
WTCJfGPLOBmoOCEHzrf1ceGGxwoRKhgfMm06kCcCjsjJzQfaulc4lRjKUoB8I6ik
+pt0R6JFE9noofiN9xCxLSjKLLjj3gkF5iAKCN9JYKNp0JTQPiq/pdUB6vrwyki8
JYtqX6SPJsLzuggNXU+yRbmuw2AbFUoAkW5SqYg8Fjiix1dAWaFaeUKiV3JJOjgE
t1BFqPOm/wrhnwJFKZgVGJ9Pcs0EVgYa+WwAEoI4F7wrSlewSX6f3g1GKi/Z6R1s
/YChMTE10uq2BwZk3HHf/FAP3BYInXQCB3xcjWUI4Bu703Tl18Uv+97HGUbDooJM
B1Vn+R6sJEyAuzbZeN60ZR6wL1AW6yciMtextyHLNgXTtvgT6jtr8DLPXw68oZVs
0PRT3mikGAptXVfcHYnn03fJIOCf4mHX2oXxxVDmxCkvIXjUgkvmwlLqELUKNEIa
ZN53gUmOHuBmr6L2hDTCZeXMS3F3UDhyfF0C00igyXHxlgeGRZX3OkULmE3UdyEY
22iBEHHnoGWI398sGIzkxkpDgaUQTY/LnkyAQ/yMyCrEChyYHy9qYFklIpjWPgWk
Da6/bf1Yr0MsRpuNH+tcxt/fmJsZAOliCsTzQhoryL0o1OSj0W6+pqseA4mC5TDy
hbNzCgF1CjP0IOXT+YoxU7ljYfkrz0Nmond2R1uAOTn76/+Gx81IOltZoXNVuucj
jAQo3y2CLv4h93TDEIHrnw7+D/VZXdfHj6HoI4Gvj/XrRAEqudGQV6Vj8udmiKbT
zAviA4sFVRRQDcbo9+FGVHEssK3QIlrzs5GFEC+nSCT5m+DCUA7XpfCdrQgS53WV
XbYCQ14OvLFZhxK/Cx6cZx9Qs2TbL6iSsDL+yaYMtZfP7Yx+UQ+hp0KXbA8hUnNQ
MHWEN9bhdjKtWdkVyF+gXkgw8C1WmcQoNjL+ILvCI3OdvwHs9JNndlk5PWvekJM/
jocUM620D8Rgh6en49Ne3ihq1LLYnHD/zoWHt8bAokr6Skw2WttBrNfTGHqKXvuy
t9ekk733MPdCNO84g4lL/g7nnQ95oIGNduJWmwIU/QXEJ26y/H3ayVldk/rZRPPQ
TDfxbyr5H8IF0XgEG6A3xlmHdU2x4daZIR1jxz0jR1dRJCFlg0mSeCXJRw/3Z+MY
Tv5WfsR8e6KKKzD4V3651hqDXoTm7/Eh2CCU9KhWAQMklhKrQKHPkUanFVWWJBLy
EOueLE535H4tUCw5Mku1Wg9rAhtaxFBeIbuhJMDNLXvR8VOUhEQHYNSKLDZFoxUo
TUHA24iIBGifmTM7B7OqQwpGFzp3a9vJM+EoCm4ZSveUzr+CRW0PB0jl8wWI2mqq
dg6JEtmuwI2Eqk27UeXMwGN2rBhGITi+4WrzL3ZPVUtAJvT6lWrSQict9lN1KOS8
TFjE9m9QPVZaEMMtxLVL3D8uJbNHLSexswIM+TUrDfkn+79ap0LLKkD7xIfYzMEw
mZozUGhclkkoMI5eHIF2pCPWaWmkupfXIrufwn4E2AV/p/xnwxK8DdvnMPNuFITn
h9zFHCcs1iR/gnLVKgx1wPQ3Qx83vtjivSLWwq0jzhQoOZ3zZbDwGISSE/plgSTh
SkcimT3Wu7z2LtOMBDmjK+AVKEvx1LLouB+bNMEeZeqh1WSRkPkJc1q8tjHhOABr
I+EOpWBBGlezEoeHS+gCojvNeSLKmJR/86LtmMmh2Glsa8s/zG6ObLsoUY5EHUT9
2j2LuEo3alBAMfRl0x2xEpYMbWabz3i1sAIB2/hd3TCxNkVeVYG81rCI348rnFz1
aNy6xiUustdZwuquwVbTdy0Mfjfew8PUPuFaW1ABSuj9FtS9rXsTnowoob4HlRL8
RwbL6bJyTeyP84KtmE0cA7a0epCRLbajnq0lUbml1PU1+55k5OxMo4A3I9qR8QBE
d7QOZ0FlALoGC8SoUZoFXIcJIotcozqQTgXKP97b130HoZAS2m+quiRtTq/WmIgs
PvlgIbt53dJhQUBMJWe6pGBSn0IqhHKmMMsZM6XcoWnvoJLVaGU3RVG5JFbOf8S3
laGNSEZBYhTEc30pzC2WoZZ3p2a24Y3cxUXtW32DnXA+8+Fk+tO0hKj37vP/T+5B
23nc/ETj+HZkT7ePIf9bHSpAWHt95yyxTp2iR7+HvAGZ6Y2VXgJdD5fptQg2KPxl
jG/2iaw81bapWVrLwBi9jWjM8ATbGPjov7vre911VNifRXwQRExfniwQCcNE+Alz
biLNbnZ4B+smVZ3hg9QqMxb/vMzBtgJjncpgaQo2NlBF0kv5BiAU+eLhKoI9AUqY
6EH6OWABIP44cvgnrKm5fAk76F9xHtlp6LPdzwqdsOlLETGpDqEjJ/lGUdvcmTYP
yJZ4GAF4ruDJVlf8anc0gTg0gJtTnvI6kTOujCuodEtQ3uOEfl8wi7dJPm5EASNy
c2bCyYh4mzsxnl119cN7I2zDw2XSP+rdecU22Lh+3UTBziJrLn/pmoL2rQJchyxD
saVx9ReP97AFqngMyxyxZcjnr4J45tanmWtXqjxlLfOzgVao1SQPWYwL8oNYGkjF
D4zJEsQCfb6p9ij0Fj80THAsOMNphmktmoj9jGeAkjFvnaYuyaDaB5SrEisTXWJN
Uql2unOMzCKdfiQ4pDeaKqHfwCxEwdgankAndGxgTyXhcCCcnPfY+rH4xYFssmge
cZJX5csNjukus4gU8kMsJIeOI9moLnUH7WbPQq1P/yYoTF+F+2KWG15mZvvtlqyM
ZXXlRWjRvGP+YZGZIf19zQsnTpx26woCcZvwSCxaONUhiVCZDnK9VWQ0w184UlIh
sMWTydMDiYNHqqTJH9AAprSvVAcrPpK1mNfjT7Sa5YL7wMz/9/eItdhGixiQz/Ng
v0DEwlF0C4dxCkcUhbhvYU4OrQ7OFkFiZ1R78rMeZNCbT1yjTfJfkBk16jMBZhCz
BWUP78I9MO2G+3EL3qiEPiKtFirLDda0+Hwf651X+ur1O6YwOLCDdy0Krj+jEDcy
OMAY8a4EdaKEExjb//OamcCLDqqqFaWVmchEuxXxkP+eQswCRLH2GJcv7a4mT7yQ
k6r1vfl502fQQ8o/uN5F8JIMhgFZfWSnrDgnpIFJrqqcSYKyB4snzWraDDpdXxY6
mEO6mfVP12rWHtc5wCXl9F+Nbml8DbcF4RwfG+5HVhqVmdDdL42PdmzqCM1tZFRX
Qg5DXYv7BcxIGAiRp1O0lp+m9VqUv9wfEyKHGWox8FbrKs+4D/79t7SebNzIv1d7
9+q87OqDf2U6Oj4zJjoWI1FtzDEVUDfP/jXz55mMz1AKSvrf4det3BPDaSBiLvZ+
/gJ7ujzCF8f6RoffHx/pP2CK4pR22O1XUt+8RlZPTp6QbsBI7H+jNpFNYraffNfH
cSuWfXrGl0AwB0T4/8BJHkD496O32Xxz5f1q9cwfDULoyULwpHCGt4xrHqFIkGUI
Fz5v6BhZ2g1fb6EFfw8QnKnZ2AkNGqCu/N3iYix/ibPJE77b4EuvwT70xCWnIhdP
e2CCjuJD/K8nFxpgW5wKC7DOYM61XV94Lj00nhPXPwERu0qvc8rHgBe6rF1KpsQZ
CjpZgyBWgtyfkQflQkUbwMcE0Ls5S+xin9vhB+WGn8GJ8RIS6c7qt9nHrRIdJNAI
RthQEiUXWIug8cKN5Ya461pSHS7jWIRYvbWgJj8Un+ETxU9o2wotY8iwesQ//Snp
qA1daJeU48ion1z6aAubAx9+UKCl4k63uKJO/feoud1bAK5paO5A8jtFWVQ5+ds3
p5xCuhX5nA0Y156xnnVolpJpgVwzxoFY+5LmPDfZr0bH969DLX/NhC/OUgvmVeJv
D9//1BQrfugDyCnay0Ozl4WLlsayM9K4hmfTW29Yi/11Rz5Jnr6eZ2fD3r4eZS1g
EYk9w1n2FsZPz0rl7x3QrKE2vzmIfq3Jxj284Sw17YPDzTT1w4VZjOtBD/65Kydl
1rOoyIm5zG9QGj4nINpHXPeZ0bpHfbngwxlyL4ohFqdLGPoQGXbbFH8TDuwyUlVw
iNTHAh4OfJK22hvf7fq7jIPKzem/4hVkTu3TNYnYa5F0fqSYXKfZYRftlhHYwyMa
Z5tMSQHutRt1PIXHwW6OI9CU1w2szDlkCiLbBY7y/udt+dkdArNoIyglVuK6IqTG
Cd1YKSU7bRg9WvdgpQWH4TEScidlg5fsvmEZbBmg6hcIWlCCa+GSr7N69IcRI19d
KzX760VXkK4lXviwOV0MoR7+1VCcs02I7D41et8OiRHdXqqj9+gFthJBzhzTiq9Y
AqhuLe3Icw5EDrzDuUH7mtH8zSJJTXpMNg1t5sloBk3Zbo8cPT9eFw8g/Ia7qfVD
gjfQnXN4aoA1tex1fIhkvxS9kB1PdfVUO5JBjESlgyxKtkzZmcCK3N2JJo14+rwG
FUzlh67pyJ3kMp/mcIvKfcix7ONCD97Hc1JVDUcg2CPHUpeoSYbD6ko1fRpmePvv
q76bDjmxF6iiwuQgeqdAkMH0aFapycMfP6ASHG+wtHf6mlC+lpQUzusJfh+yYHi3
KA302R5Y5CXq4Q7TciVsxxsI3QnAa3+qNag3twONH2q9uUOPkmcLjAb5Q6Ly1iGm
ckyPehlwWHmYWf3cRjz1UvMQ3dh0kVZuW1yc0ZU1VnVA+snbxf9GzAwFd4AtWK2T
HOy8gawx9zC9RBSJz3XU0pZDVPPrScKsb7Sjyfw2dsc4Q4LxeUW+ltNC4Gy57Za1
NzyioXkL/sCfhFm6gi/3gk2TcW+7Z+Tj7ZQE4QgoCsoYiPUSdMWp90H4bMES3vwo
3shhinEI+JyLrRoo+I0E8SMbxG6rcnlTlE8mBYOEi+5904ftBR0TCSj4gFopLcPG
Iu+ygKOCUhval/cZgfu4BYIX7SbakgxbZe6YphowOZesKSqVEu7+iizLqKERC6sG
ZMysf89Vc8SoiBBySuFp89NDvtR8kCHP+0ygbBFV8wEI+sOJ6d/BfBDpSeyroLU2
/tO1v6s+mXSDSzLy4nXo/KXxR/irlhLY3h87HONHIbW9GPyzchZ1qah4IbXKkMsY
gUpiuqkDsJ8f+ix4Gn8fucWmY1aE48xWREBGVCtl9N/Cr26j85iJdGFAuN7o63Fi
LptON2cMc8GgYsmbug8T+7+R+j2D4lcHTO+UVSxzM+nISI2yG1It4xdtCTj98kSh
eNA6gJJL3MWHubCpsdsDqSSnOrssw7nH7vguC3XImeoj+M5gi2BrvjY2rYDkl9O6
2y/+dErUz1fpuxun+VppYvty0hKYbXZPoCf6hdzpr+cAi1tsdVygbCquvBe3T7Eq
PHBOyR9QVq3+2DAK/E8U8jkiSkbRqlH+ZLAV0u90EA7mKYIAJuPT/wF2VXtORxsk
aTUGcFjHkgS2g9Jks/GR14wzm6IsjGml24vqEvLxPuMd8jD2ptVsUNU7R1HYT/sq
jaoYIMKu7rtIVJHbsy94L5dQR07y+Wbzm5LsuAyrBZk22t0DJfRoRO3R+sgwOME7
JThRIGVi8B4Hg45gPHeyAtfMpXIBBvUi/1TmQVVKz4v4pR19bp22qUGBuE0d0Ucj
vsn62GbM6bMUE3YQbUS9nz+jplMcnqpp1yp4widpwbIjKwY7ns4gm+RSoU6MOPjd
rk2ZURCO3NVhmFtBiWVgqYwkx2TTmPXqcHfSFAnDjFLqWtGQYNvnW37Uc9VlxWFg
MmZONUXsXsmcjWVBodKHRGLJXuw6EqHM2nvgskidoKayxrenCGxqEVVY38pPANUC
JPUnCv1hUTiAeac9jvPtCKiYQ+kgP8kKRfhIsR+glmZtwL01SX2DRpwjyw5OjPre
+aek4RH7swP8ZhjZDn5uyNzDd6Ck//XBiQtTlDQRkpOfFgrm/GDNUIGkyjKa+78m
VBHez1dhJ+FxDiI4SkvmAm/6RjEZ0nRjTKAYfO5TN+Jcm4+5A8pUY/Ood95wHURZ
tlMd6bhlmoIL6RuFmOoSH8PVGvniKH8752oC4ONKpUnRHkRDDp1v6B0TJD1Zc+0N
WnFIR8r1lChMGDkF4nYeATkR5WYczPUkTMOL9hk8FVZ8wm9XLSNSpJWWVIQh6SgH
Kdr7QNHl7tK5rAy5W6ECNUb+owG6N5HBHveX1oe34XMGLG583NRf81cdnaG/S8dq
otjXE9EKoJTltx/5Ah1yRiDa6EDUUDZuQ72hDb8Z4Dr7odJTgtGwJMRS8/DGsvfy
Qed1MI4Tgvk7gZfPu6Z3S/0L3t/OnzhVitzrGwKkeJ57PDMwFwMc3BLoCXbM2Jza
WMne+JbK7Yz6JMQNM3HVsmJz9WXga7yObGWqNARZEaaQYIAb78srpTHhwAcSDJL8
nzNLD0mlo4T4SIo+OSz9Gcc3CVGp/mJGMYTGn4VOmY4BeGlGhuOaPTFH88DLHRoA
74Q5FTO1AsvsjticuYCnNsn+CnKj3lFWxgc29nQhi3uI2AJDsS6X9PCR6FjBYJpm
y1xA5vi+DQKuCZQos4Amyn8tQfcdAPSWs/FuAsBHuYz7G07ePi/G0Uw/3K+KiG3U
kXcR5baIZaq8HqEA8EJ48Ql9PojPP+JLMmVYInjvytAVPqVW6M2V2IA4v0EMP6Ng
hNTHiyiLsbXTzjjCLfmVK5snLS4j9GwxrYscEbiHPwjaOMac3EQcqNkpJP/GpNqP
8/g6b5ClYTciR8mn9/QTV9/XL3Q0xIxt38lALlj1g8mz1hNEL8mkYUiUUSJQK+o5
0NXl39DduKurTHYeP+DWTUYttAhXVnGjE0hb9kAdh1J7Vu5WTkaXGj6UcxjwQNPk
e3d/kP0a5t4T8tP1Cl3XLoJlcErVuXkwcGxBEjBBfneuySojOYJHvDaNQ0/dwjyF
JxBIbTu+sEPkm42pjVBp1q6JOIjsW8m5Z3562YBUWBT5w7GLGuGUYNCxXDuXbWY/
KnZ/ylbzEIMy3RPZWY4kbSRDPy6sg4K68Wo6OjewygStD3JERGVxhfNbmb0ylV6a
vtwlq9UPwuSB0rnMYHjzYpsuVd8yQsjMlgTIgq7eUacDgIAZ1x+5qxxCdglPHQZ6
3oW9zT48j05nk1NfpBFh6deKUhW6VclzpKT2cbgi3TCUOhEpNpMFlEowUyK10qSx
HgICxMoQQmuCpu7/TdpoI2neboAhcwNPkuBbUiGWjxqc9KRRnxBn+ABB9nWHM94w
reBGgG0rxmp27wp33LpE2eNhMgVDc7W/qDN5vLEd7nGhM+534KEKpY1KMkS0xdh0
LlKAAA4XVbiP5nugCHwnMFP1kGbdTj5CP31IB/5m5PWed4DbslR/ZABvBvzLuHON
3bHJXgdselQoGIjSBiFiO6jOBAVU3UHFPuGEwWaJ7TYqvADSeH7ZWYdLIEwHoOwB
The0KdHgYKmUkx0zJ2/1gvUjgAzYXtDpV9Z68mw+/xVV2AqliDFjuwp+/+7aMcJt
VA5Q6uGgBUl1zP1CDTSlBRLgGBk4yY1cOLAco7k6QYQPdq/fPE40k7We95w1CzCl
9xm12cvt4CH7T4kSWxp/2YEZ7C1gTQKoZYDjgvc5sMK0c18dumsTOAUA9qPCU2BL
T45jEgc7TLViFchjb/ekppd3lbsG037xkNgyOjiSCZC0Jyuc5Dxa3XY3+skNrudT
o9vktrUbG/rAvcSNUXEpXA1S00BY6P23HI3krxylPtCXhGwaGb1bnrB6bqWiC2HX
4KA24vdgDFnnrEJ8qNYPRcpFiQtS0KeIpfv6ejh12BAv0lKfYUZyK0vOB+4r4c5N
ND1+LnenFG2SxJTKkiF1QQ4/+iw3U7sdrMIqVM5WWjNz+82EsbYw+0dr9P9fjdtF
E/qF1HRTmRD4xJZh6Yd+7cMeNVz3AX7l2gTxqJIBXcyj+2pdeyITNQk15MTGHpjh
CUFAkNsBOeTaOqsQfNVpKWgav8BKaek7q1HO+MTepksDSSd53ZgoucRwpw+QaIVF
ji77Y+sddiFBqCxE6S8Zd9EL8uBrrGFmKGsP464r7cpP0iR0eW4oSgPIInid9aHJ
+m3Fel21TLdq9VJyvy3FsxjlaSZU6evTwElc0Gbr5MFI0ImRj0jYQGg3SH1zUjZe
XWHtPzrSwPAixmNin5jB3ABcld2syWZHrTlqFMVX3cRhIZa3FdN8zJE3V8hA2sPG
l85YqPN481TvD5/AK/mbmVC8vPK7yUqtKraqLFhUyai21QJ0lV6thd1JZGNt4Ssn
dfIqUH5PHss9KWRkZsSFTrachFs8JzaJDLsZLsrNjyuvjx2wSthwBiA0PTHQW23q
yw8AednamPO6MPJ9CmQ6OvFBHmBqMFaFaeoL2zSV3Ny9+vZGtqufsFts0563xXkk
ZGth85RYM/hHbxM3k6U+6ca/C9Fnh3+jlVOMKriG3L9Tc1BcOOZm2pHqHHK+6zgj
srJ34m/cbU4tbFy8EQLyLKiFeS59nUbvISafV0dJkSLQWRaAhwDJx57ETp8eAvom
i9kT9ry49flARuGSbYYBt2ig5D5GMgvtZ97buqs8gnQ72C3uHDYnNyKmD5GjwTEZ
r7TknDlw57Ha0Wj5mPXSg/ewPaPfgS0Pmp8ApBnVcPcJLa+jqil4ou26gYofdbe6
OI6GVMrSA9XYd83mjJKlvhYkXv35BLbh35UsPbdlVtdV0fZpuc0PsQtx4qX+x2WD
SybY0BeiBnPh5xT8+zkC2BoJKDq9QbZcDPSWffjU0Mh2JBY2Rs/NuYvf8Poq3r9S
lZB055uw1StShZpvcvku+WZrTIt5geuZYTuiApwhdMn8fLFItmDrEQ8cVKxnBGRa
DILKDj2n85Uwb3Gxa3glhPWhLnJpBFrSLUtEIGHuKHz8jxDH7uiK7LlDgmmekMrH
rXZZ+GkXiD+OZ8r7T8XgrdO6+pcWJunab8zMRaZUmcVNCfLXwqeYtmfK9xf9lv01
eNZC7yQnDPDGR7uBqDiyOwwYDqo+fLqgOLRX1aiqNx35dvC8cjnD8oAagBuLQrPX
rHxFAek5vEOZg3/aRXbp67ZKy2Tbnqg1jsTYQlbS2MAO8s51tNCbjkQ5BuET0Jmh
f8EL7DcsdqJ1cklsqo9zQ9Wsh8p/kcS+anTLYbZCy6vPh7IXPBn+eX78PA49oHof
t9VePEohYxy0TEGQCEQZjT+vUz/peR9bqNbtPiaJc1u2OsgKuCApYp+1LQpIdAtZ
TbYgxF0j3k0tmjKNCsqboQ3pIXuCPqnxDxhoZa0S1gxN/C13zqVvIpzpypSmiBan
GB8kQPCyfn1Vu3tFNTiIXbyoy0K1/OR2I9WePHlZyHbhawmFjdkjBJmA3uWAzRZf
8knPl2uef4y5TslQD/2pfZ9f0M2SezZ6oBrJiEQ5y77V/YCTf18FJ2SiXRTRQf1H
GzMXdkt/X1pdikTuzFd32mgnXkAJYuP1sEnHWoa3uwNT40387sga3vpfBCOFz1mB
D6DpZiCtMmW2OjB+EjY8+IuMUTJQcpocwlQpgzQ2/BKCZMi+kumF1GnRhbSJVAFD
rKL6xYbx3wWp8+UT4xCC7tyVV7aLBDOnT5bXgqiPw8GKnoZznGIdCu6K61IR/De6
1cKQVn3XFgPhYWXWNaRe2+gBv5AHVo1+JUlAEwi5iyC4NdUtbmFqYWa+dmbtNRtX
6fam4CC3XH3I2iZf46N+QWCo/eyMA5ZhCNiJMfuGXkLnrTo1sMV+9bmPq4d2T4hy
yqgjYWJabqlzBoZxUeLmFsrwTPx/yAmc0C78tqw7cQEtSg6Yp3wwy7+uAjwLCT4h
arDYu39DGlekNphb03Ts2aRf9w/47YAr9jAeZL3ka1cQOH49nutIRH6XWbZvuq/b
jXm38vk6rEdd2Jet+mAnxzUZXY0XQ4UHpd3sYSnDC7ECSwSDwz0qSFcLLc7kpq4M
yqahdLzU33FaYIns/v2QtniNUR0G09bnIxoMDhxNjMVBBO948GmIo/mefyhWq1V+
6D+WzJ/r+U4mVRV73upw/EwynogfhnBQnFvGFJtqiae5NF/4gDveqTjPsiKM8cXM
x0OIWV8XuBSe+hkJ1xyOaCY8MgKGqrN8cKBfdMTPbK526bGjyA91eGM8iBkR/tEX
gGXEmjoMhiLpMg9FWrMfwWKru7+Gsl2irM1O/qeIZlL0zPNgZi9bsXE0VdHsSPd4
LY9ue8csPx9/qSAgFJvyAtYraq2YTSz9MMG3MTKfHgEUO1Hp9eo4mk5ovLFkYJsB
siFf1hKjLbjBzPOFV+OKe3vO2TrXWuKBc5qx8fBXcwcLSGU+fotqqeWafkY70/0a
6/hPsCsHbQ9I50SvNqJoCfao3LDIm4D0/mR09UR82gLazWtRVEpt9DsmI9xi2mSQ
u6xHSYqEutztH02kgB5te7zO00eGM0KNt14aZHg90eybx/0UfbCYUrEqUm5HCsyA
xxF8Z/aZrynQsbAPmwmUKBQqAqekwZhW6FouZ6fXC7N4cM27rmRZZH8rq/wGhHId
uPyqzTHQuODw2WOkB+oCqji4XAqwWeHjVhEGssx56WaQEwje9VrkSr8rphNumRD6
5uwT3jHJKzf3qe045R3a4fdSIsAwgtxSSNP32WyzmErAkSzcC0TZUcf33u1YH6s7
iX3Qap0JNALMm5mEB96Tjes07SsLt+xmpdiHpuuiroDimxKcjYXwicROWWTAqrbu
ooSqsvU2Rx9oOoSp2GuXZZSA0whjB8wbGYbP1HQjNgRfUtUyWKAFkPjiJfcjkOnW
MUp/5gE5IpASOP49R5hbpT8zmV8PWwn6g5UwBVWec+Mh9grvExO6aIMvHVhTqMGQ
2wjAiiYat+WRZ7OarodWoo23zyFmW4STvmnWrgtO0dTTaW0KHFk5C8DVrbUvCeC5
upZiW+yroSw2Mix365FS8PcRUbLWPMSJN2HQeMfik6fEH6+LrPTY5sqFh1/WTJF0
v9dtWVUEfY5A2omXA83Vvmbuh2Y+NZB1CyLBz1Ep1F2AN/ZZzfw6jdCQZ8bpu4ti
qBKoLPTCw22XLbXhhUNJGVI+wOycIYaNpEDYx1BvseQTzJAh8TdyfSYwWLIXZb/Y
SkOEAYZXJpNGemh+D9ih9zdfF6gZTngGwoK18IL86hghkWVnejsowhDF61ir7fZr
FIzqxyoKrxt3A5em9QY7fwX+e3Lymm99CwIQJe2JdjwHNUHEqk65ZNf342qkqKml
JBjely/5rWfI33gt4M1cqkH+CgyX57uNiUhT+aWq746G1zIz7TKocnVepEkF3DZd
pulFWvFwq7e97+abIACRDXCoaIchDdFvhTKynJX+9uFr+4lKA2/2dd4mneyp6ocG
NlZ/f6wMi3FN/VXPmd8IIaMgTDahdCbMoQiz2Afnq9X44Xptj0SLCsGrOGlergBL
3Ady3wzrXCsrAxU6oj45TrKrQDz/WVcJu2WNYkEvNVXPIJLi/A5HAU2SdOt/PV4n
h84NkWNlv/CUfHeI/67bdbmCEekdb/aGmoL9QpQiQg7VgCUMszY9G/1GwZPH68IX
hXOLtbN5U14kUO1GVlNrJ1epoAS6EdHwpvlnOTpVJ/UJWMQNcLJuzhLUM+v5wbY2
t3jehxyLHXyyy1zXeJ+yOT+v+H8KPyJLMHwGeG/JNmH8+CYgo/ntrnC6psTmRrD7
tEtfkIO2nFRbq4ERxL5D+IcjHBq3L+iSXns7LqvXkwpce80/qEmVkh6UE07KqL7W
aoEwkwseTl917jd/JL7dcU+kgPb2cpaWNO+BbmUqMc3QUXiu6APBcU+4+mzilL8S
TrKsNF9C26A2VHax20rrsTrOvMUHeCwn8BzoUa5gAM0J2rMDxR5StxDdTTyIR3f6
emLtrD/aIQLwFoCaRYcWKDvyx7TNfZsyjSuezqunuLMzaXe7/aKZNxwZ17ksnCuf
v/DbhF8j4XC/mRNZRYUlTYt6Cn9aH+m7kKQ1LoQf9/xep+cAwlZ5J0aatUxiyYVI
qN/4vEeDqkr2YLQZCVevC+FPV2k8gyHS8uFwmc3ySJc4I89eBxt9VApPyGfukc1g
r9GMH8oBg/MumZHr8/tigU/NnyfNMLbVMDeb4JUbIZ5Qicnf/0PPpGA2eTN/u4sU
0D3SOFYXQtEfV48T7eIjpZ6yGvhnQoFfbOa73F9K6qkc598AhmesLp5nrp/fQ6qm
JC1LDufEzjks+uUGXb9okzCyogUY/CaBrgIbA2ddC1X3aM5okEZ6YWRLudNeJxM4
++Tpvp9fOtam8XyREj6oJaknjs0dW26NCgcuyi4sQsIxap5Z9dzrlm2K4AXFSNOi
BEkDWVZ6fANVmIOa6G9f3zcN8caJIUBAFlE1fp4Axk5K6A/3AX1O/Jalb1a6AbiY
k3yimatPWEI875efRTGdVyxuT/Rn+t0cEk3fsTSxJvvcAJMp7U4c0kM1Xc/MaxOf
4o7GDPwWB8+X02jlpP9BRB/+I+EQahBSjvCRQPyAnWmeFcWTgcut60o3936i0YoL
AaEspy8EOIPQquMFr6mpTpltFBMiJiu2z0HtxAcrOi0LYlw1S7MGbU1/L/tnpIxI
dK0nJsKKpGQzvR33WE0V2E5LreZS/OJi7L+pD8+ie619lKaOuRDAXQj8M2EW503y
nwXJyRR20tooVt78x9cBCBZuOgxMcnITxrKYL9hPSC1uDfO5x3N+Rgp0cDSFBMhH
QK40sGaTuPa6M5lEc2G0XZQIDMPAwTIZveC9GrUcMlnUL8ttavmKfGoGc1697zdV
THSDHLWa8m+IZC2xumgxPxyXYk0sfhny9jojMCnbGTesiyTYPlXuqwE4wjhH0Jpc
/u6/csYD9V/RZLhrCf8DNQPXMIOzxFw3yEQi0xz5v6+AjZt1wyPLSR1NalAOeHwF
wMjxHav+lf4G3x4IEJ3zxxwkCqaeSQwgeTl8vQOmApBmaF/n0Cya8BMVyhhG7Klf
RAGMTL97zD/4Kfy48s+g8a1lpbxWnRR/VC2NKouJkqedvWa2AoHSo1/d80fnoWLr
r2HpOS2EG5jMbsht1zJHJdjpVGvZtHBbpHm4odi5IV+PQjscg2lgCR5ny0JtifXq
7DDrEJbHBMex2bap6qskO0BtLn1YT2bTBoFDWxfh+Gu9PctnYVzZFKhORGedrDyp
nea3cqf4g6o74qOB8tFyVaT+yLJejzG4Z5dX9BgI3KTzGsirtxsiOhIevbtrq57k
KPtSlDFlv7WvxvLA8QVlN/VkY9Wc6rzw+FYRs9wn4eJnRG7JWCfECERAQDx+se8X
sd/q61t3FQHYxz66kVyRN8/L5Pvfpk4/+5v33blR4eYCU/YeGqyHje4xPRxW8zIr
qc/Vl1L4H42YTbNzioJbdbhkw/xCflNjpV3PMK6yUeWf5hEpTHFyxlAAHWmfwNE4
ahrhUE5cMH6bKoWUcnkmB3qm3YypEpv8RHMqeLunQEYzkJtjy9yF5fLS/leU4Vu9
2BlnxcZ64IQ2xXyygRWp3gjUWoWfN/3fhw0TEajxfl5wH2lZ3XETbvOp2lR2+tlD
9q6KxaFeAyxbPnWoGD3XakQl/AG2rflZlCxCd5RoJSdGWpZEaIEAX21V8fYslwOt
ey+chqxsZOE3vzin7DurglxZcTc2yDRgAWWJSxMyzr2jyXrJgg0ACjF1G5BTuwLj
3TmZh/ELfT8KXpaaPs2Ns/BjKSbCRnc6C0exnVNVu5dtVXKbrNu9cr88i7q8QdEz
b+1JmhIZRzOY3MH+iOiX1RhgU6QMb37nUqnfAG626gdv97PoFyzobKS6365Lk0PK
J8LXASHcRahGCVzN2b482WQkygO3nKMh9HeeMwtFv9c9vgrPUvUcjNup4U+ADqnl
vIQdCgNQgsegOug0p+TpmW78G7AFVxJ7JVLb/2Qy2hO9yUMTwywQwaEmtyS/yrU3
EpANy6xla9Vazm0rICOTrk9gqIlKMeYwWXODpjPd6er4KkYRzSU9PnZC/5XeVCNM
0xEWlZHyYE3vaARmUyT1V2AhFdOZPx7w2+G5QeJdg8CQTDF11JR37iKExPCCbEsu
X1I241pO//5JkwRvQ1N74J+xOXaKZxrpdQTqgsIhb3usX8BmuoqVM1toPzEKN7P+
NLBs2nS7s+cvv/kNyBwdILrDh2DWHjBIL/9Af8yD+2QbuVZdCbyTX0TW1gXwK5RF
WRI3S9wi/5J6Z3DUJHaagaq7xI+Rv8aGJe9OPg93EqorRAUaW/d1xXbPlTUWzCMx
auxmtE0FS/PHCr8AJ20TSdULgo5gC0WG3DTSwyLpqnaM8Hv20wiUN9cCXzJ/Tk1Z
7CetxwESZhbU/eBbGj8tkyt5jd2C90JCDwgp6dYKS8hyDJMzGXYA5nBYvH+wJtVT
WUstvzW12zmBh8kbmam9Z5cRbO2hNzEotpBBMMMnP78vcY0Bwxbz86CdcHQJ+3OY
DicebBOV7mse3iS5SP9YJdNbwRqOaPLw1gC7IsMnjOv/oIQaT7SSehGa8MJ79tdt
TDStBTRHHC67Js5smD0rvEbkjFnbWvm9LdMP9w3KosLdQjVD2f2hDMNDsPyOqA38
gapk2cB1azqYbugAFzRJFCyoZ7IpT/0k+hJMucg98D5yylUJz/HjNI6FeWOC8tbq
4+M66u+GqhYOFVYek3M4b3AAPqP3xldkax2YP6X+aaROz12GhJNoQFYvLK9ymlYK
sTWgg3e6kl6tpUC829Z4E6jrQiGj7hvWHeWW1NunZzu4RmL9+5B1zubrMR7UEq+1
zWVsP87Nj3gnP6coWEtICzHF3wVrtTj4Y0l7I0SphX2tO4TC3XhElPSk9grhgui+
nozWrWq5c4Qmqa1/k42Cksh8shuAbhunMWiUz41Ep/4jmCz7kgnFY6s0JWqHHaco
o2mcSFzH5jSTEUgV9SXzE0U64fURLYNm0qNQpNaOPx9gJ2+dDOTXPVywgMoMFZWw
FsmAELwt0B/nfprxucYqG2NSXdJJxh+tAn+KPp2DhbtZCKmUMXwOBlEZGDa8cIeC
PP/g9ctysf5WzC87hY4RuOZS2jbSqJAqVSqZHcrTGbTjV+yTZUvtpWK2D2yXfJTC
yQAqJ0tmC7WAfVnc3bs/EKqLHdg3iNDmAfVOXFGpcVW03M1Bnm0OjufA0hFsCLnA
q+68ARYoMYZoa1DAA80r1nZ17s5P6AklTM0akCeVv49etT9AiTLdEsbDm8L89StN
WTdktbf1VRW3RRILJbLGZCr12OGENNAqbJtSn9tS06pq5/MK5omOAra0mpHfxx3w
r2hRD2ufuLJ0mqHeg2D1K2ycn4ggjEgel5DeNK8BcNEaMzB56Y3/zWMTbJ3Lt40L
EClp99Ltfw/9pF0x56Vv2d5eSQ/bVPJshVgetYUmtpXMkWtGOKE8/tMQ7bNJBnf/
XaViZJBVLlWj05LHbFwVfgrQCom3dnhpNhbK0znyPd94V+ryEb3LKSgxfOrBGhMY
trzncbCtjbGgvu2sPeblOu4NMnjFrEDYkyDeSWC7tAske3cPEBpDEC9wNW5fsslT
aTemEc25oOklx0YPanonPsYlYRshcOpYmqxIEtFwVATKD2OXPPMxVEKXVXnWWYAc
nvUOc9cVQ40JuT3jQLxfXU9j7clYMR2zr7RBODVMJn5s6qFy8F+dI7QKfAFrdBq3
CNunljEvxkSww24ZCuFX7vwPPQHiCMGLCsprwp47WtJPwh8ZV7nzWPt6DO96jZ58
tFbNKsVd0TA/quOie8YFlMNICuVW1BzwgmAz8kwf4bA1jef3FlOKRaZvohRfdUh3
jkcW3DmKOOP0SU3B+teY+hySdIf1cBn6CJJgQimXpK6NaElGLVXBPcyDkD1swb/j
KoOJaQ0XM/uWHerG5nAiSaM13tFrKzV7S1AnrAzP6RJnRzdD8QkcMWySg2eGtIrw
h9q5zSwYILEMZ3sLXx4O56yDtTqkmlYGAB0m9ssxAaYAK7n4cUBjGv4y/KUPWcWq
DhYui+uWnv39XXclL9S7aV8yNI1LZQcM4xQFX5HVm20DmLzb5/fBB6X4hDCWxofu
YcJGUihCRhDjq8lwRowp09yIeYaVXoJCyT5uxFK9vgQhYBxLxrlj8hdMGl3VyQnp
pNxzWegAW7kX1QIMdEary1I/+MCQOgnWHWjrcr1SD09hlwUgGP0EEM7zFDDFi2V1
lThA7qPFItcqcXGlsAuBGSkPBidmlYVEURYI8oHn15JEHicJGLdTkTDFy+ELbk+B
ZeTWC4o91irQH4VWMDCmCl60qZ0/TK21wH2G93XMXeU95Hlj79D78bOSwzWA9UA+
Jn433QSdu79QRscypq7+fu//VE5//eZsiqDF1Q4ASXa8LjhgXswWUicNaBm93m6W
XJW/xCdkuA6YyL4Fk8HGoReUyPgwV6eN7jSPNNvgQGAIS4/jdmjI3DINCzJE4tUw
+XbbBQ/iOsFCjTlRKfnalsSW0jXS6IBZocJ3iY/+YnHuFHC1bfQqGhP7I3ug2z3T
bzynyM+RmpiSgV5ZxGoQ5/WgxxfEredTEWSkCuVPly+ppPTkOftmS0gi50NMDD25
jTichBgB2d0qbbiaEnS/iCgEy9uBFp+UG2scjKB+AYxW+2Z89aHKmcOyzG+2n9Zs
xcEKrEz0kl4T7z01NUTsab/5J2lcq2u8EQQP1bVKIGt4qiY/KSYZkbqFqmGbxxQd
Oxu51Q3WOXM7vPPvzH3CTabOF5q817e0AAkLG66UR86rK/pXcSDSv80ea521+MwO
LBTovTA0wbxzmTPEqAlqGF9yHwQXCTYC3o3ruo7rxA/H0WGI8hC4WkzejajuJg5y
ed72wCFjQb0IeAi39KUfC9Mv1rdyrzgPSMTFXWug3i9CbEfGIiHchMx9ozmS5Qko
RDH3KSN49Ch48p03M5tmnWFLK9Rr0319lZicyLVaG69CU4KElm7TIu/OPnyEIz0T
BDsBYLnY4LVP3BzKkLN2zVR+f5t882rnNCUBMBmjGPmSebD4Cqyg3Rv08QVzBogO
7sunEWgZKJwh9oAtI6wxRfPc0sMxn3Funs3Coxg7cS2pXidj58l9WVzf7Pp/5aM1
BmJmgKpWqlbuTPHr4sUOYMVapE7/zws1udzeWgA7ofH9HwaHUBbdoT1gMzh0iKFG
Y7YGU/cXOouMFDTBgWRM8w9taz2HmojCjqEUGUyg6ohLHt+ySfuxQgWn8xwDgtzz
PrcqcckQtdENMUfYh0kJEMpcCquxuURZL8u92lHDte2k5Ok4SfW4uimcPCTHq4Mf
pFun+l83t8cHh29N+b6/kUcaQd6GOVsfDdoON1rBzqAJtOgN2qlUny5yJrCbKAAw
IlAeNutx9h2K0nKUU6X5Gt70wPTYbE73f1Rpn40l7PQL2/qEN+JagSrtDlSJrZvh
HSqUi8WV+f5RbPzbRc0HTKCSj0HYI8t49crUPxUzHxYlETlB7AKEJHKNjLfuGk72
MPf8zbwASE5eqz0xRhZg9cDtNrgGfaiiyAdENcfIvEpco21yt+/C3YQ5Z9/iDEbU
D7Z6OJwt9Nabk/pImSjszPFv6MQCir8g5VB6reI115tiGvFAjwR3hP1Y7UB9H07c
e6n7yl+l2/7UAPmzPeZrmIrMWzkM99YoLtsrOteLTV1VnNAnjRfFW5eivaE9j3Pe
1pnIYY9dINl6sm4aHQBOi5g8MWgh+9ukPsAiuJXx/yx3gQ0YiUMgq5/OT3uGsLEg
WEuTR4k+1Jwl4GcnJPj9utLNp7ngVLKMNEV0VpXRK3vZsboXCGyGNijzgXxIkLew
Vi9RJfRNPaEcWqentmF5RAKrE7THw/oiqFg6aV4Jmq5z9Racx4Mk5V98TRIhhft0
spUBU9Rk5JtYigj/RRhY4WbMra+WQly5na1yLffBVaROSz9dzRcite9EfoLAphLD
Hth5sNKcS32gTzjatRbO8NOEeWau42J7HscXFSA7oc5gp3Z5mO5Or+fBcqa3XVFT
VeGhsqS29kq/i8ipVkyTARCXabFe5um+w3YSgKaAudxn3YHy54cOs0oc0DYfDYu4
xDMpqah6fblH6N8QWwXNQ8a01QEIHzH3dDPVem2ndZlT1tPbG/jpcgmzvr7/OE66
tnC/n2m3zqmc4m/KsAOM9RTQJlat0Xe0l/Hv+tNMZ5KRQEmHwgAFwOZPL19J4Epw
h4SMAadg6vAa+BK1pcrLApmLU6YeFEqczbSfsve+thPdzTYTpLDRu0DJzbKKQZh0
rqeACPpFVyzHZ+U8aZFUcjrokJv3cyU6lw4xNZgcZRwCv3pMhMltnIQE3iXpsCZZ
p4WHeGnu7JBKMwfOMlL+m4MHQC7uXN1C3pFy/iluNiQsV+YolqDg5kjMZ9MaePuM
Yo2rcxiTHCqzKgp+gvnPeS4CNCZAZqqCtbzaLN/Svo5ossA6N5L5G2sz0x4Xjku5
T2HWHhTW1Q97tC8Wm4RLBhxOH2Ht3DXhMc6HgSiVbDpglrKsK0LDmwgI6U93B5ml
aW2x4i0iJxpc5mYlMzxDNQwGxyhekO3bjaSQEYm3doZltOkbU6TOnpj70XUU+oEj
gdqB8n0ySwpkXRII4K3Av0rj/9PHaMxBfAcdjcNzvytwSJ28t/es5jl5irRx+k+i
UjxzGxQbprt2C6POGttpic4b2bETJ+qfk925cj5kFf7joq1GeYPTMm6gD3D21Gze
clDHGpSSZaAV2wbwGwlk1IrTf51XEDCLEfJgGMO5Cw7Kt2U/h/TMeWF8zvXAFsze
xbk7TBPgcM/pzu+7IhuptUUysc7QTh2UF7vrUmng0RYipK14bjH/j6t2F3hIQpQ6
dDWg5/GVvmZDQE4tLd+IPBHsbalq2KbiL/1b6DZPvmEWDsXjQ1blZuvCaRZf8jqJ
ZG2+cSJUV4rTJo023MecZrotirB0aIxEY3s4hBi0u8Fz3qlkeR7e4wu96i4oEtQI
2v8oHA7V23z0ukKKwXudbK7k1Aq9c/AyCjcRf4my0epOyFNtWsdGGIiAIxNOjLN+
uQcyurLopemVoTi/vlFj5I32FlxIdX8X08x6qIqgMfMSAH9J18xzeOHumTh66zY+
HDQXYZny4nUihMGyTiJf93bdexvPFDYeSPhjv7jdVtY4VTt6bRCksru8GxJ9+dKl
YoLjwTS6HFZLr/YvDpevny79xQLcJNPfpkcGsaGNM0KvcuWGUZtxgdnuu3ivfd0T
y/9lC8qv7uNu+2ejYpAcLXgmbvgxiXdvEysBqYVUfb2bE+ipU4AnTA0fuS2zFp2/
MNuy0GowVwPzFh/4MFXcdmaiKx1tKHzbHUafgLy84uajm+Qx/IhexANHqGr5MWDN
6S2GadTaQb7QKw4ciHfFgMmDb9+cRfsszqP5LpEvvP1goHs5b9us7/7CIbBLjsAm
ywLVd6vsOKWh4ESyDSXvyNJkr0ackmcXaaUI9D/cyOGegqs+a67WxEHesgyD82j/
GkowQfshIsxXMr8h1Hy5MugN3jxXePCzLvqvjPTeR0WvvZzqRNrbrZsI5u+1Sq/Y
LFx4++vFopBnhTnrPyR8tFlievTM8qSb5dsoOEVwB99tjn+QIDjHVwFdOqizuONh
JsV4O6vxg/WxrSsUrux2/d03Bpmi5F6vEKuq+roMeiNbC8O2aoTcxA1uOyfINCOP
t2I9RYqqwZMgaz+0lSfLCZWyYXjKUiFrQHPhXcB1sRDIJm2WfSdtK15pq79NU4ML
7Pq7qZUMCUHycoTOhIpJFtWeQ8s1UMhAWZUqpJVXFYOXb5knN78M20vUZy/7orZR
X0urwZSnVzHsOKkJjEqYb57+L2aP//Ga68hR/DEC0WTMergivcLnJwrmWgHe1BBD
sNkmz4i9SAwupyYLGBZGJbH8PUyo8mm6NGD3+Wh/rPx0bNfpu4mBjArl4gMm+ncJ
h3D3+tuOL0Nd5QDsg0mzA3wMJ5SZwumsFv0rXMtowl7thMQs925acxLkpl9Gb58Y
EF5NjXbNYVz60Gk9dPB500BTmsJdPfuqZ7IQDVOY/WQ9q5bVKydKZyt3jJ88tiVt
aUi/aHW6Hihm1W8akd8AhCdPsB//f67BuFq+hMdJsaZzmr3AorWeDBOpkMuM7Pr3
gyePtK5gznbwIGKOIp6v2SqJETeVH+aTIk5iCVvJkfLmll80sJzpKd0oBK0icUDG
740YKbrPYgQQlQw7t9sRMgYi1q2UcYaCh9FsUyhyQEVwGhiz72ynHMO4F+1GX6gX
AU577bHMYx7ExNKMmm1AZj8UoFK8dVD3NeJ8ArwXXt1+S1H/33+lANT0prJ6lVq4
OwhSK64vjHTog5HtyZoy4Zhfs7WloN/9kg2GDIBOvuh5GfsFmP7iYm0/7k/h+OCP
F+bmTVEweZUbsfYIatdIbIZ68sh88uGfHm/C0d8CqGcu24TTKvdDmJG1soN1zOZd
sgn+5iNhpeB/0+Td5XrSmPrH2zeoAdPBXk/LBorF4LcR+VeP3Ee7/58sQa7tdPMN
q+cc0m65sGbVgWIssx/CBq6FP88HInveRcmzHrWUiLF34K0DBuR878Spwp6FgdxH
wNvLgw+APs8QwAGJ0dAB114kxuoDRBEYmYeuL1vfeps+mYuFeqhUbKIYQwfzXG7v
uctUFgduXJXVGB2Urd+6x4f4+OzublL9eF2nb3DupQbCNWWT7TwtdBRpIO/6X7ej
lPjjUo0EW9wjNLLnCnOZ+rLrGGl6ZIjNSs1sqIjS1C2q5FUORR0TdUd6r6gOFmuA
c+zCiPLwmNDcKZx+5hKKfef3q3PAzkmKq2cGobndfVyKIcaXPH1vmLh80llY9kit
4qEOt4KbK3BzRt35dOa3hQY4dtutaIE1haM0dQBa8kSj0BORBUPMYVaZeHNDf0mL
jN7PcMor1KZx5dNcYuvARrZOdqrkSDh6lzsZf8OCj9SpBNPuer6aM7MqSWY7FqCR
OXIoHcFRIKeOn+7smYCEcFayzvFKeNNVNUMNqAYBUqzicUqiEVBkeQN3UXaHFCzp
m8V1hYO8R3xqBSAnhDBwqnPNhpk2ibc0aAgdWBIeH59jWcF+XUgoNMw41eZ68cWo
81JWTOs3dBzYarD660XSTtIEPwrHV7+7y+knT6c2g45E1Wf4iW8/cXLyfOt5mLy4
voFxW+ICEJStPvgMSxO2IvC2t1AuOEAT4iX9lqJzkofFiSp3ZHSpOvp0fIf8+Qz4
G2tPwmisRoNUvyMVWPVKyO/xneG4rkkrLLu56ALqTng0S25DNZcIxsqf51ods66b
v7kzYOvWs1hmFSUeUDZqIqymJN19OMpnjm1pTwYsn6zR1NgdOgLpudr85tGpw6Pw
a0UH6oYXWl6E5kswwaKKbXBVl/LBHI96pz+RqckS2RyTS87noP6GxMoI/Aop2oqG
BIig8dpztsyB8H4b4rP87lwJyBhtDNVy3+QNoe2D1Q31DOM3I8GtbmjETUI1APtu
4f/KiwVxU/1zjTEb1Tqw8Fjl3sAjyirdjIPbwLlJDAzXRd1WRWJ+ISUYzEOnaRtD
mm+Sh5NbYgNyMKMwkgWvWXqfj4kLlp+MirKGYGUoku5a/XpHBxee4ajeO2dlkrXB
ZwFjvwF4C2QovvUcZG+wE0n3RXcPcMskQTwdDvXbk1I+LNUuu8oxPx1YuJF6HfIJ
asyoDe6dA4BPqmF7uW9d0sIfF44eP+bZpJeE2VzKCeyxgVELwovw3y2OSkQz9bnc
Yd7lE3hSlFgq2EgAs3mFoDBYxZv3MHcT8k+HvzuV0+iIZrD3Y4NGLyLT9w0stebn
08Ms2OWQVc84OGlQ/0u8FeUVcs3UxrIPyeHZdH5/Nf9X3UCXxH5Z6XOdUhGeLYJr
4x7J0AweLnEFiBgOijsi8hatyBxdWZ9H2oIANDGGqhQIsb6BrrDgA/rKedtb3gXV
0FLh+9m5ug/FEEBFwIRdaWdaOmaTzyf8597GNliUSxNR/UnfhB9QhIbisnrdlMHo
hz5eiIa6TNnELz/ekI0D4TvCylQ8XwQImi4/JRo4vi3xm6ytc79zq2gshVnAXAqV
E0QDUNfpIk+deOClALUqqIG/bfZg+PPhpuanEwjmg2ejzacF/B8x1sJHxNIfnZVw
8nkWsBEHCjljMzSgUsHW9np5qOgTkje9hmAIxsLVx+xyJw762j2BpcLDF46oC2mx
SUfgNyeY4skiRd6EBlEk3bpjEYMzM/ESyC7wU4iU+BQDF0iIRlcxfeMtbeKviHLG
2wbI/s5iizQnbq7OthFfTT3qN/le7UZ+cSwihIDxJrC+VscbqrFmO1A6YuGeVyiW
qpL9Zk13txbpgdD9y4I9os1eb1Fq1YS3rlBUtW0qRHXHKefErzukzHcL47mJkNq8
y3cceYGBD8wb39Ca9zMSIoA61awuLA8/IM4fDQHGadRCESvoBiGYHnIqZXmlgaqh
sNWU1B551i4UvyCl6HtWN3CBW7SUOkL9w1wQu8L0P4oP7KBY/Ei4eo8DJTZAkTqc
WNfek19q8a+JbC2yqYg1dMHLNWgMkGzIY04ZG2F20D9CJA8FzJlaX3bTLVzY7uYv
Si7OJOit/3kFdKv97E9iw14LvNRX+LkD09Rc9WQSqVyMDU/eKqBjDgSLlRd4yzgt
hUnNh7ln0xoO2lym0khTpRLhRKftpqzgFpTujpGRDj/Pe8k7xEiMJsMYg1+gjUyl
SoNhno78stxLwcH8AkrQT6+KYJdP5umHK1q7BJ9ws9lqOUXVE4ilXEQMQBoIuHH1
7MBG9swHGksP62z9bF8ngIs03SF//LyBatu30LIRbJKj2xTNsMc4Z9rXUZtVvnlv
OFqBpCfBrR3bUtcgXmJgwYLnADnLdudsguh6kkgpUPlNU9CnH2RErhZyyKgykfQw
ue8o0v47fk+Vzj4DNAnS26mQ9W4l+EoXeZXAO7VdyyxjgZqpDdQ5ib/EoCxZS7ae
J/uRDeHT0cM7aopCpq0XnG0yFEWWXy0eqCSqKCc8euvFY1ilOInln9ucBcBemrtl
g6bH6qYWw/jk00APrAOpYR541GfgbitVglH5+Y17bxj9V2M4Hv99smhxfFCh5a95
HJJIWU147qbnUOsnjyqbrgvjgHLDwsBqfeOx7rkHUoqtmURFmEU9N1HD365CwC6N
klX9Qlzzdo9AiWlPsQK4I32dAbxj0wKgQuYmtZ25dXl3+09YLyXgkwMIOypQk4Uj
QTdx5PkEljWnWneJGBUyOOuH3GWwHv2su0icU3zTKkc3wKbwTjRsiQ4YzBRqTzi0
bhnvqBRA/59ubvZIRu1RzXoo/V4ka/pRZlxRKTUMcVFROnPGlOmkEI29bhwId/xx
NZMCq30u3qX0dpXxfHcsL8DEry8K0FODLj47NnjNe252h8ygWILGilVuH5pOTAMJ
BbcjFnDUkMuCfZ+xIboE13Hna/GzcroVD3rqbiBYR1poSbnTB3Xq1/iKdldBaPUu
aL5+MNb9SdYPc8ZieXOQ9m22UfhdxjUbkM5PajbaA97IyAfv9dLW9hY1NC1wpjIK
k7hVR4r6hCcsydNus0OvBktXoVBekyOaiWov4LF1qHoLECI6hlAy/VcZFvlQ8HAq
LwAAsLNQKgU45K1I2zXAumpjFRfeghtplM22nzUicvPkyWUynsrIz+0wI8x6rigG
ExWWahZUBpXeChkG2YKAfTEkv1tevX8loDA6ZpTPt5QT1+sSi+3zEgS1dnaO+mfd
0H6TNCUDm4tOH0JmrnCwK0ual/I8FOE0iSJVEl6V3S3QE8R9d7kSA/62oNaDXqN/
oCHZd5Oum5dY221lZP/jdsroQ3Rm7VAjSVyGuaVYJLNbDTyhqabOpuhPCMo8b2nY
MNYjApSahFTAuouNjFHKbOt8dZmKMGIdT1pFBnKBQAZDPafYArxS1x+Aam7glwG3
mHf6UafjBRhTm5ZDrTvhknPoiAGoaK9L/YIxst3+ChgEysDJwT1BNfh0IdX7Svk0
FjsUaUZ1T3Fl78QO3wDw5wcXl5+KZ4T9nKrXEbbs5DZFylVYoABIH8bzj7h6xI1m
9rolJIhbp3Q6bJCNYERAkrQ0q4NMg4+kXI0awIiI9QYY0/GgCiscvXRWTEQBILQj
ItFt8RI4beL6WtpCIYSl1FMYAC2dah5uurCtg/8Dv6gbfK45cDSa+RtQuZv0iBdT
o8Klc0wbuk2wkIAnB4aflB5rA9Ab8ax/TMLhyb4L9dUuQ+MkRawz9hhrkA391Roe
RhuWYBhcLZhIlLhfxLO3itpRwLXGBMM0OwZQqK17LXMzTIrgvS8MidQvay19/lbt
Ng86AvCL9iKbdAZvhIGp3Xzf34U+ghIGT3sYAg5ihCxEuHSYUeoJ0XIKKJcF9qVx
MlO4wLWJiCPA7eAEsW2CKUKzHFvj/IT/x7ZSHEBi3mxc31DH17oKosqbj2RtT6a0
/P1Qp+6KQhPGPv2hsrYp5kYqRrYu+/ydNOH2YTV0uZnPFhXiXIvo7QiTZST0I4D6
oVUOP4+rmPApY1rkrJE+ZECtDdtq0zo8DxWsaaENXfDiZKLPrjhBS4xfk6tD16Dt
pQnfiGWrhFs1rHuPFEQ4R7nDoHE2YrsJCRSxLIXrD0rNUODdWG0v/zc1BSgLIel1
nlSAKvvoHsIL4uMP/i51y6r2M/1rqK2v/zVI0BW5ZVdJ1xZLOrvGNk000LdzFAme
KyqJaa+a190NMKgwZM/H0ZyE35Fwr9FvSKl+pcUNVFapLz2QWAat7CKm5EEAdyQI
DboNyywiDeOxAuE2lGvK8NHaHV6P5obp62lRPNDTGI/wFkfYdyRTEjkCORyL1OwI
WgUv7gJp7qIud/hZSJweKeuPdmvQMBwlSZDvF9+PKyypWu9nq+zgHwTWOI9HY6gH
esYd1w5+D/PWPHjnK0Dlk+WjLrk94wq2fFgARef0lEaGrNOdqrZ6YemdOVg83Aq1
F5ZqHgw41iA1Nky5ChiHs7z/5ufWnLHSjak+xMpFpXvvgbsgV/hFgyB9+IZurz9H
waxpH37dgterMtBacS2IsLFXzAcUDq/cUQ0qNiYURB/j7JiFKNx5C2G2eKlVrNOI
pF4dAgFmN2cmZ3IY+/sq0EKeha8Q0b5ooF+IFNzO76Qtrz3xqCOihvkZjknT92gT
EkhL2hUnaHY6EmEaDwZzwA4bkUpjo8gRynZAFCvaPn6C3PdyQXggr1vjPwUpzUbN
7fzZJzE2rqJZXyUz0zUzRRmTXTJfqWtQN/5qxdX88FiGpTjEveN6+pyGaYApPxWP
zF2RQ4mvPqfHUyWyUAPU3uJl1c3QN1KphcQ0o1dAiEOOsEGGkc2roc7snHJtUXoI
HTzPW+/DP7bt5OYxaCWapu17z/ro7dwRKBk926sUMK+ZtUppKOHQsoj7lImWXUbu
vgKXmzgGYQLaGlJocUtfHsR67Y6WhONxHovxZJRBsjR9LkPxngeAWeQl1jXv9TO4
jk2In/xSqwoG7S1JFSDbvhR9Cu0CM66URSpXWMxBgggybNnywwZC6RtyrZQmlN2D
vZ8PfrQ/6sJJ/+iURz52QI0AXQK3Nvf4bRVcvjBBkXN4CBiTLmUEvCoaFapg2fX+
5+KCEu5+52cc1ecs4nav6Hw9NRj+kJxBYIXt3XJYR31p0rHn3D2onCyk8Ba5iFa4
bhJPb7UBGurxfB5Cubk5ArXYoE1AYw0Hi5i2IHQPohN/BDyYWouzkjI9LfNZ8On6
YAmlkjHY6dCCW2Gd4AKfWoCFtzOi9FAKUTqk9hZPHkHiraaeYfRIfM75uNi4rAcG
QBE/2NhEjJhHMihn3+Fj+8DSDik6l6uilkWeIdr74bX0Va72f6Sa2a8Hw1SFKB0b
xf9TYJj6opaVjALa2TpWhvk4v/5RRaUxFxizVUo6g0VyDWE8Uazj0/VupUjeQCh/
TbbmmDjd9tDHsC3dbjnKOmFLWuyBsgaRFKkJ5sJlT4Ou1dDH0SrwHzu/fLFlPzLd
6RsKoW2+vJYBAkFIScnu0vGjI3oJDcXL9Zw2GmL9BJNDrScK+Ln9lnQG17C3Hdkk
1iG7refH3mAmiFT5hEdMNGdNmgmRODXD416i7KXV4dALfnd2XQumLHIhTnTIUmBe
YQWSF7+2gptw6swfnxjV4rjA4fF2Cxk8I+ltV3AzNSzytPpCp7LLY4YuHso7deT/
nPq53fU4jpklqisasQ63tzikAO318lEr7Lop2xGfqHvxu0O/FC3rUS3x8wKB6PVi
ttUwNL7ScexUiMfbM7d82TU5fnQPnKQYfcfxJRTik2kfdcqszvMsdmkQXXEE8eXv
5IJ2riWJmNcQGGJ0eX6/rJ/hdCLc3ISijeCzbEBQw2GKhIa1d9cisFVnTYgZDJOJ
GNCA8z0w/l2Ss+maO5NKHQ5TmfP+Ldq5unb1/+3HE8n+X8Bwc0rpbHiTMUJGpfP3
1XNjK4l0xAN4iQoYfAauOZ5xmaBpqu4CY7Z7gahB8WJ2cwPgQwTHwQ0PihZxnRaA
RZYPvbEXmX5oFyOQS7elHDv4eXdBiUZRrP7OQH4t68Vvzo/pEDzTnc0Rd1+uDmWU
TC/h/3MMeOGbR6iybKstDARZ9YfuLqg2wERmDthzB4jieEPvfMNqGMbtnkAfXLz4
xm9gTbLzqNHpmFw2vZI+8WV41MLxzV0vE95P45eIJJUt1HLWIS4AzvPWHE8zdb84
+B7D09C4IHlHkXC0ypS4aWtWg2mtV9wQUtWH0qy0Yl//TfMGlw/QOoIJ4hbefI6w
LRZuw+hCBOBzUO3Kl+OH691HfCYDuMmgwir3q9QaUpqKW/1IbhZA2EIhNoinKHL3
TEI71tWmyg5RwUOwjxRh0gzwMRYy2duhGn/BiwrIpPkYB5RZNdmSy2ZHAPA/DR6K
osWJs9Qy1dsiCIgpkNWEJcRT9gfv9+r3lk6dV7pROqMK4sOk6G+bpSFdNfBLMSQl
Rp/Jj/AnSHPVnnexBEuiACSA9GXAhyyStanHjteT9eFQmKdQwjDwD8BqQRq3Ks9n
XPCP1hnI2RWQfONFiCqLeYf4JZLnwZPtT9qqLSod3oUP52jmfVTKY0Xifgvb1lgE
MgZD/PcowOianIhSMK9D8lQBtvxYZGAZHG4eE8NwR1p/cDFnqMHihfLShCIcJ+Hw
1JXbgZGGxL7DS7UuWxwBFWQQz7MSYDxKI6clhbMk/kJ2xUkUG9ID5IT9UzoTYnyF
y/z+KJ6ZqrHBVfPTSB6TxmLvaGMCfuUxmD2LtY6SebSWHDtK/YtFh5QegsAZNTs5
Wd5TE42+KSJbLBEqfbOIOmuzlmLDESucaNRrmHNX68dLy1GO6JeeZLCAcJy9bXkI
75P3HX2AzuTetzFIwZLtbC6x2H/09Rf3rJY3Gy6wFGWo5Z7rY1g/j3ET9e4ap4D5
UPEZ9e8cuxpNXQWyGFCarkOorOlK+bOeQwuupRR5ONUm5Xp4w3a7e29XwOsydIXZ
o32IpeWxKWGBrPyqh97v+MArlvkr7XPRE3gEV1hw/sXxYCMmyMeulip/yr0OwTz5
LHIxNaZTrHzasQ8EOLbHvImS5wbZY5YxX4+QsXGX1JZCbI/b4rqalVYkrJ3bq7Cq
0PQCqeSdPg4ORhwcKx9EAX19tRqvNUEfuFUMZetS0ZAAODL1wlILgvywhVYj+O+r
DT1Kh4FPJM+Opm0yDZ7e/Ozikr5yCsPK0+N1fzbQ6OAOPq6dlMWj0Vy/zqviBFL4
8FiUYYDjYP/8QpiUZ9rU2FJ6fhtslzyTxRk07uYWh1cirf7gvnRHuRbhr1mNEZWK
+I+dVw7eIzCx872ne1OZg4OPty8yu5aNhZOktz70YoTpYVDrjl7Oy1RKaxI/ukN6
eVwE1Qu7T4SFuuCiKHVV21tPOJY3HE4u8ZESC2/IlfIpnq6M8pNjdu0skBV0zamD
3CZq02yE7jgUb/nFk/wQr38pZaXGJlC3AP11XzkCxMBwvvbLxBtZY4o/4mO1b66h
QveqViF3mSeuAhhA6xO5cs7fgHg6pZQyunWGe5Cj9ZeMe5iBS1n8bbI05JdrTOw1
Oj5KH8ODnIlo2ynITz+yY/ge+e58u5ZkeLN2lKXpn4gQaAjooC1qyUqUUxVPmBjP
ZtisFajyJrH9wrGTkVp4XKzFTmUnLL4aVKv349tEHQp46/MM3eybnf7aRnfICfsd
LtYWlVeddZv8lhEvc6X8A4OaYZsEG8LBaruJ9Cr199lyoHHBaMIB+VMcOLy5QxXO
ma2W/3AxoWbvHzwGsGM90PZsWTwkrweyJGL8Sj83gmjg6FYwXYazLfUszJU/OCYL
z2IHVZbRIBGLtKbcEQc3MSqYusenIB6hZwkQKohPpzRy9qvJBLoEr5dDFIMg+LTy
0v+w4+Xl/mEdL7v6kUCM3efhL49Fy/IzqZP5pRjF8kGKRrrD9p51mr7nAPBtB22P
Lfs6RTrSFaeZPLzga7y93FTH1SAWtONy1VU5juMl1iP9Cl9BoNtayPAcHtaaEafz
yuYmvtM1hHxqtyZ7FGF5igTZXa1D9QELzFOs8go9VSs14DprS8ZlpF8CaVI/sM3i
J7uFKpy78GHAiqQoJXqKKiwiWOYPYgjAY5qKC6B2GmyrtHKxeXMYdHwQPlDFEOLL
5p641RpcVubnyRHTlmfdM7NphTOFpPNGhnHw2TbKrfnQpwhjn+QnuplBe0JYJb1W
FFWMO/t/HO+p8lqQp5qMtqKMqqzQdFQQdOvp+gGH04D3RxhAXWLws5qI/Jenc7fs
CLGgXafpllx0OVtVm9KkipTQlC1eT8yB1TISHCQan9fGm00+p0Qg+F6uauHp+CP2
FsBnEl0WSe1qeBpv/799uGnjgHWXV8C/nwJK10yRXLnTyafYUciI/ADS5yeV9Awq
ObUsy5Bc2MTg4ESeK5hRwzhxh+2ZdULGNN+WeLKrOgRJbxU4vfXa9esMFiOIad4n
wUPStOkgv0ZV+S4hyKY8DuSU0UWJDQbF37IRO68SAl+ERE0b/xOe/SWCXkvq5s5F
l3Ek1pDclmi7k5csoDxuGXVo/M8X3QvoG/fgW7SsYuNfEwl2q7QSgzMSYrFqMBjs
YUGtt76ASVVm20MenrPppxfkNreguod5ikusbFI6ns+MxM0QAbrG2wYvdqHe7qg7
Mw8D1QvJeoA8i/VFnNFF2SSh8tGtTY9ti6496sOfLSf8WwPIFQwdSdwT8hP3w56t
RJbl517G/DOSeAC5LeZ2QO8mmAP5wA7d95fHchXhiwrTatnAL81d557Z448I1cxv
/3xQncu41sNSb0gzeqBlG2EJG1auYt5+Sajv24/u29R19tuMt2XQopbadnXkEe8b
a/cF7bkGoY32xfk4bojm9+mqU4ixixlKt4FbbejWUPZVG7DQHpxOld5ULJDqbFGR
UK3p6Pj+KLXsX9JBbgLFj5kkWdVr7pAnQQFdcKYeKSgbmGT9MPd0l+vfU22g5zOT
mHyamk9In0KKfht41V031Ew061Wo0tTKEavgT01VPaW8soM1If92TTUOq0r5GW3w
jA/TeWyfTNb2fguDa2xee9wu8PO7bT4c5914vdvu5r2J2x+4iO5uzCHQQ9Ujdpbj
3PYInJwPiGBkoh9w20Dy2vgyeUgfPcI0cN11F4d6keDdlbDUWXKA8inIGf3TXqKp
G+7DnWW92zU2coRv3pNAg8fzlm4sZ3h6VNziCefWB69PH6b+PjAnJlmOFnwO0Q3a
cfb94ybAJHrI5WtOu6tpmHD1ySHTpaJSP0xDV7Efz67mOXqXlCFx52jJyxyooO7u
ebgRMJpk4IWk7s8507wiXgKk7Yqey2qvk1SDPvdiOtF59zsHhpSB57eykbPGspYy
hGoxzl6fYh8CNJeV1YZ1OPbelcbxYER3CMYUODfY/S0Qf72Wg4xKBFSHHXy4mC2m
QvPPf1+dGOu9xJ58I44m/KFrmB1AzeW9462AUawxK/W7CdXrwCYUoNDyjetmBsOB
s5h7p+pHpdODAOBJkPx7wr2JiJ3WP30+PRt7/78/68xOsOBugWPl00aFIebRkoGP
Go2B1tO6WKlolPgLXep3UHQa9Ph0bqqC2knnHpteBPx3xBmPPuEalsx0I/GVI9+i
ywrIMW7zERnXVrdDAFVKeA/UoGSmTj1F4gvcBGtm9001wNBQyUaunCO7XEWGDwnj
7Bzi6kfI/qX+CWwQiBGXKkllIPEIE4o98ketIeyTWb8VSfUt/elii2pXNVlt4Ewg
lmURAfGdZIT3R7DaZ7T6ChFOQmxxKYQQKlgEFGlHG/RT7aFZ15zRO5FBrUOH9AKl
I/VEe9dqpeo5B6YUqG8DdXWcPrReojJIX/sO4P3kgVqMmsUcV8oa1/CFhB5U0x2P
vfbrFv65kiWxEOuiKkF+PspjEVgrqDjOR9teb9pQeWcatcpf7MVRJMBGrVfN0Jfv
wNC/cXlONi4O81uR0y+lRbDDs5Oa9gtNcV2dm/rcjZVMH+G6rqHyu21Xv0xtIc5M
92jwVIXEX2k7LDP58ImURdLmmRjYvVAWhKWAJAcsa+G2o+MKGHesUXXaITdWuK52
/U54gk/HUjKtyurTrF1COHHAfLvXV3moLUit8xR6iFIByfXsgE4JpslOeBxZAr62
vZTiRfLb/Q92rXNCezco8UtgI4XI0kup9DgNr9VdAQb4PbFjEhhw2qwujBukNlwq
1CeFxNxbHvM6HVzKMsDFp9PgwzutdIDqmaewwOgnQqqlG/moybrmgtUZauJZHDT9
H9tp+1oFJuuox8IJ9oWHVrwuEidz2aJ1CJpyYzpj3nw1gHImF7dAa1sFb0wMg54N
lIi+tgqS8xMytLMHGjyKkMVFATs+suaPIhJ+mN5tugFME+cjfnN2xtrncFpx0UYD
lLsH7OKuDqti8aIyw1VFL47kYlPusIJhkitn93aG2nUsPS2QTXyj6LSkHFeDTO1p
vDwFGnFQMHbjLhK7PyKNKnOsyJSRFkIhgNLW25GJ6gqNHnLf3AQ8AsWLMfFRCCW4
Tu29mGE/oKibHqWHbEoRF2+FMcHfUeLRPi7bGdIqZ5xLqDJPFSdRrCM/eSaJH8qr
pYpd3iM0nfjS8cn1+f3ibq2F2G/VCqocrOfl3Rf4zT4zWoy2Cm8FIeZv9hJOJloV
10Inb5GnjVtpLUnOOY10myxf1Qfezw3hTG7SiGbfVUiDjVxxGJ0lZWSxzQdGsz7d
Lf+l7IEc0xbY+svb9Um8RXbl2A6Ki2NENVBLkOLVw1Bh8kEdnRrBWIaSqJhXrEWm
Mbdp8Jceo9knv+q0B06Vm+33TlVZ7bxMKUnmugpj0n3hfReqHWQtDEknVpJ+XTkt
U1OFrhhcwDf+g1f4E71AY3o0EuLEVBTZMcu5NRDP62ixl2ZIX7WPkdQHldUHsaEd
Wg6v+H76UP6+/SdypIAvRS3NcyRhfOXmzn1SVCGF27pSeE+P70tiw7EuPM7DX6vK
iqd7GibRJQsLTO5tpqmUX8rT16YAfmpPFDEzuZu6VB9QzStmCnzyeBjYZqafTtt8
PC2qRc1gMvYJtAl0DnmB1ReFvB+IVXf6GU+WBl3wqvTRlXJeTRbMDA0n6PBFgNKQ
GTt9bS4RhPSnFsQh9yEfIcqeXwSm26wndqR1VgkQRXpL174y8G8JbFKOC6i4dUdm
m1NgSL+AeE3X713EDWuE6ulszxy4u+6nRRwYYIDB+Fj1onNBa7TgEvu+Us1ZOWD4
0+TjEnanlTTzSxJ13gnf+SiS7+XeAoE+PtWd3pcnhv/qGhqje2imMfQJ3j+pfr9+
BKd6e8NVL65dzoFcXEYGdM2T+5+OYRCUAVUFwoNIo8bPn5bN1qqEHxK2XFqNvo7c
gIwIuCbUJbH/UqfRLxIg4OohlSFSNho9vvP5tDi4G+G6ncgcSrh8bTZd+qpeRdX2
0ChIo6o47zk0iPbYIAlNU1tWzx8D8Pn7RwQAKKAAFd936Qykn4p+PfBveJ2E324I
Z1L17rx3tKIf2qt7bhrgT23Bk4m9InjzNXS0g2sq6Nw6Z1ZXpW0kBLru5MAfEgLP
0fXjSSYanDxp2+xktuMirtqF9n9zmJWwMBLv8by9UKWQegqtdeImsdsewzOZ1l1w
Uqjj0mBerOqr4+mt3YXEJYxwC+tUeIKC/rZDsoMRjU1iNxOnFmBfz0c3Xctp1rpO
yqvS1sEpOwBRKRH9dwgivPt/AoNwvJtHOFWJ01VA6K86iU4I37AwHeP14p7BOF6u
zLtBXnmQ04r75R+fYL6Nys2UxB+Wv95mMtvPYV34U/PnNCoUWDmM5lKFuq5D9pcO
gPLRiOg2AEo2RBOeuZC5l7WXLRSZDgkKNdfMsjVxCAvG10UKSINw4rr/hu0UxnJj
nxyWrTBSvh9wXjDJIdDCVgTrDjTDjiw+zdpgBNEi4fm2hcVjplliWZTb2r1+GSel
oiHKDHO5sosVqL6d9oATBAIfNaKfmy/ActWXi0opbkj4rfJC45iF4wN+t6XrktTu
BUsHj+m5pXWpU1tXPC/obVog2UpiDxa496bVi98DhSTUJqdtCj66CGKIgdOxEMNP
IYOae7xQFExBJlc6RpoZ0Nr83AVEbiQBSl3edl06j4TtGQoeNiaZi6B5c8pyuKmt
TjSQYY7AGdS4mXiteY/sV67sbs+H42HNhNO6BvucxKG7FN0TNhsqahyu++7udgIo
Pj7/KnSmJmT6pxEsYZfsQlE65hZft3UG9EenwhXyw1L26ds4EYSl+WGfRUKfd9Wk
m08Q/Q1QDzxPdwudNGzd5tAIT6zXlTLDnU09g2MmD4mpqQYVwgc1i717Bg85hBmP
Kf+Dvl5zooFm5EzhHCZ4Q66vV6ZWgtpElN9s485dQ8LLoZONNxW+Oz0paCxR362A
Ht5CqKHcnMjBqssfBqgySNGxQA++Sl3Xqtp9PHTnrWC4G4zwiRsu1GoFnU0rBYci
6CNYIZKtKl6pZb8qEGzPVwWgg3D8s8ZJZxD4FuLSQcEtUecNc4sLHrERNPIg02gb
mjWd1Q42rs+GihYLHHoHgADugSxlog5YVYqJAGL0pRxWm0lUlmrTT3wuSr32/7ig
WO4OmEXt5DATKZL/3jq3sFT+KivLg9Fuujh2gcDQw9I+XavY/1UCnu0XeVX2Kjn9
rrCBj8mnQ9QSyaoVX/WV12SGteOX3A0y2MAH8U2tqA96RLEYqMEqk3IS6ni5G5o/
yoj4zC9n2xqfoATXHiREqtMibhz02qcViNnK82R6dPrr2/VhfHcDv1W+n0/kxqgp
aVpLt9k5WoL7iYigudzxL7W9OSqxFamVcPE//0ddCfG6WRnCzSKIVN2pfNrNMIii
NDhw5XD+Ch4lYQVdztf8/2jq0aQuPgEGafhU+5mFkTiPHXU9CT2R86mB6OxVsMxZ
GLXhir7TlH9sOkum5IlkMOxt6ijKu2Ry/wxdSzpPHEuJIzU0Eg+L389hRWGydeNd
8q8uD5TnKTRo4gpw0Hkcn9UzKQtCtRn+IwA3G51ZTODdKUW5khNBLyNRBF+S2Hos
Euh/AFKD8cgqqIElXuZ6ThqjY05wPBpGbLlX0GcJ9GKo7f394rB99/seGLOJBNxR
hp/EG/kVbU2dVoqW6MnBBU36wEGIPhHDUvRc5Xx4CICAvztW2itO3Wj4yhR99NYW
cVxe2XPO9oP166+BUfRlfZ2tgBM8MbLm2LBjAb+C+SdityTqR+s+O+vmM+e37nq2
JbeNYjw/c6e51s5ZqnUuYf1fF1tyJopFmqLieP/E6uBZjqBMfpScuPSyuFO6/na7
gmp7RfipY2HI+qlYJMYjX4QVTAEYrEpKpHRn6BKt2PK78pkitEVLm9ygpAtGOvfo
42jobQhA/VgzpfpjRBG3oV+pLMepQEDtP3YVWxEmizMq6iJUm2LbUdE8TMqhi1s8
2YaBnGzFLAHxsT/lwWUHkz7capellV6D3nG8pNoZ9lOwopreKyimIO/TldNniyCQ
D5Fu01ItHWOOaQyjzf2PgiP1kaPpOKesYPiUJYzHmmKthAOCuIfAssbt+OBTjlxn
LC+7MOVpdu9HSBols7HpTfNMfMCFoZpO0480sjlIMkgWJ7Nompg5YE6cYNxP3ofY
7MbdPw99VBu6Z7INsGGsRnUzCQJaFewumB4nz/y+0xwE49uLju8v3Kqtc/EQSywO
cvRI2fAy6/8wLN9V5WAmmXxwohfyt+ow/lPQ0pApx8bd21ytJRJdt2tllVsgF9wJ
DGGl2WWXOy5f9FL/nsWf5HRtd1y8eAQHe/RGmMKOetg8xewvlJVP+i3DVShn3uZe
nosYDGrKh3I2stGOLm45Yl21DZn5UFjVYQZAk1otbOY8O1nwONU7AzqnbFP/7V8r
ecM+XkgAu5Fzxi6bivd01lohmErb44pAlhpbEiVB5DM6vINh3X6YOzoFoU+LHwbP
zTwnqNoAfdGserDaNjluP8WkfPw1awywQIuLx+nXYy9LwknQjMRHv/wbzZ1L8Oku
/G24ZP0L+7/kSoHuVgVJBQwlDokSNOlcL+66eBN48+OfX/Mv0m9J/YCS+wDKO2kD
DzarUqoHN5RlG9liqWL4G94IYHF+UfLGCxBXQcvW/4UgQDsfTDFa/NYk0pByKHiD
E3iwv2+qVaxvHgSAuB7i+PW20qBNeJMaR6EwwnsqaVh6dUkyNNz4VykmJk5pp6vB
RsUJ+fA8WPzkassMcUUB45sMdH51atocxj1CBI8TsY+QxDOCimUzHVlTvoYOHLa6
egXF0TozAdSF0P/YRCENmWGC4F0i8YXbSOU0JeTELQwEKIsroY3nawNT9qch7cTs
tVACr6VXKwnNK4axHn31OuVY/Nf6Zz9SIQcwEtW0yUjrttMQZuPxIdFaReeZrB4O
tNcnJx+5CwLxqHwok+tQGZmkdckuuVPFy/q0fi/XPlG1j5Bk5NMSVcTErpMDdyVH
9Frgl/1Ke0lcH2NHwo6W2fv1zMES4p9aFPhO3hfJeGfkelc8KvflQR+uVsgWr6p3
9g3wWVhQEEjyNuyoFyv9jjwYXEZwf3SB7Vqq3srquXsC9VqTF+Jda3xO9kvsqfeE
zL5VVMCFc1VKyehAIJdvmEBvAO+rdkt0ziHFLP1x9FCEmmzKYDEv98WAiQJnsQx8
6RfgrIPHnoxi2PkNNN4BNVqS3BIO9WvIizz2LCpOTR/KftVIYi1hd4Dr7H1lUZDn
JqFutTar2rqPd8Il7CItemN/2pMlGVu2p/nQfHpPeDDNHNWDWf6Q9s9ilJlEU4a/
Te/rIpFcR2RN2zipQWi5cAwi109Cljf5H1cYyVzEABNs/FPIkKeJkWg/jmqzL8aU
Zv18O0Tgx6pRGcNYNzvsaUfg21T818qZvPHnR9ckFbEEvVDD9Fyt+QAEiCqK13KC
8M//UToZZJsnno1sMbSeAF2d5r1xzeigTQR00fKa8jHtA0mApbjBh1RI8idkvnpM
sw+lUIk0a9h9wa35zu/Qw3otbwLx/Yj7JYBvBJpTbfICvPKBOW2tioPi8z4c/yT9
YkR0Hq2Hw6iUtTP6VQiuCtLX0Uy8Nik8WoUWBqcSeoPsg9k3nZEoiae6vojguDfx
WqyfkCl7NTMRmTiUSufc/Y3moarDEOUOeeKjeH2oOyKZQkLtbuP+DskqLKscY4tZ
JcrW+Bxrp1O6eKicPj/WUI9/vhA87oHWtOBo3RW+AP2gisTEAxKbAwtnAQGBhbcj
oIjxi4+zvTYMZmPqVuwmPDxfe6QheTDHGNJO6TvTe64v8CiG7qIzUdsftGkX4SRT
d1dxvKMqRVE6L081ftLfRSk+3lr4/taveAOGzNHYO12EW8qfOh0l0hcKbWmHBstV
yG4vptdSxtMhoPOgYPlzxe8xvxVuZj02B/Vvahd8P4YJJpTWp4KbZZFDX1Tu4tvr
XZ7qmv3uwf+PNZIvC3euHRDASGNAb+HEs3qHg0qVLv3qZs9r6Lm5hq6z1mlQPqhX
49VSCL+dbnyW+NJQoukLt4qmhb3EAxw1hbVzyldvjSC7minzT+M45cQ4tiXFViyD
ye1qTUDxm+oYf3NOw+cUd6NFmeH1eOxUDV75soJ7MJOULXCgbMNeUzoRbPYMRMiY
Vfvg+wAS6LkD8LLLC5n1QWNP9GBwaSNGQm5Qf0fI/A5ynBQ/C/ifTlE/p8O9gcqz
SORaEJoXW0wOmHLzw8qUCtI4abppHwmF6QDMSbglaXACsiEnsye+IriBLBEzId2l
9+xsQPFeRpxldr1TYhqrV5n4TStwvNLKsTSL9LnhJAVj4cz72xG7PicI8VEzUQhq
OlUczPQOHAurCIdLcV4+/VsHFNOvgP9Ag1zW5zrFkb2U5HcFngRvHhC7gDURaUg7
TLhVvExqKjTomYKhj+rAUq0/JkniZwF/Scggd5DQr6bex2Zj+yIjH0i7rVqlKav3
ViZ2lj6QjqRULUkL3g0KmOpbXhUxbOLpg0g6RxgAkzdJWa+GfDXKWvW0JRlNsNvF
LOL6OpbLBG1Xx0O/8wO8iDgFC9qTg27gfFQyzBrE6V+0R+NnuLKxGtwWfoM0RuMH
2jJI3stVXEoS0kdS+GndHHcVywJFNMJWj3PMy6gWwABhrbmbrrZg2AHS+zwUQA0Z
Ini0ZsjpwENsNLvte0oue1OX59mQpAfFWLOkMy/vaox9gn3ib+IIg2yShvmSNnHj
zxiza8WBQY3P1rmPF42nCjB0BqcnqvNsB2CWSNt1Eo3ItEHUV4PhOtM3Mg9xtg4g
d3RlIoCpVJVeDnnIh46ZuiJigk39rSv6K8hKVUji0yulC9/L8V5oS+LYwMFc47fF
+pOn1KJt7jN9xCvCqJTNKD0dMcHrJQlzxYhyWIRV9izSaRXaDXZRFzYcS/KUea3V
9rRIoN30M9Rzhfb2ayH906vN4PtKsBZ5eL9t0s1QjxGVZ/ysjn9TgX+CvE8cg1H1
xXj28YAckTqAPtkd6rnMKJAg72ZmGERDrDVifLOOEZSsHvj8QYDMGRWAl/Yawib/
FOQoQRQ1sdqxjMQ0j96iSmh+IV0JJEHQ3t0+cl7OwLZs1yfJxvf6mSPyOEvjqNS/
UT5btHMmp+IwlF4LZLsx7gFefHRYBk2NAPTI5AhcbsEJeTM53hbXP3vpLitKFucY
/JG3fgRIMbLPs/1pPXf7uGK07SMnh6S6Bdn5VhrVThonv1QvXyR1Nck6MOpaKehU
N1PF2KUcjZvGq0wLiqLptf4mc+IGCrGZo7BmgHFsrYWTBuUiaeIeXAUX/b2IuKtr
DmAlg58Q12l//sWoFSq72xR23ebptMFK+1t/4flGJdVka2GD4SS7tMT5gjyL5aAC
dF6UHlYnmSo7CN9zI3BLUraiJqbjhWEIlM912NmXLwSB/TXxmnpFgSfsSqmtXZXO
05/UsIX0FnP/m5mg8Vs4de478rRDLGV26wCfcJzzg0E7nWNbp/lj8OCu+6wDmD6w
OrnBQv5O9q0zWyFK3tDFnsS6Oo0CnsZDTW0FgRr19MsJ6bgvLlflItmclxKzhCeB
iQF9Z5t/Dm+kZtEH4CAgSoqpOAKbD9uU+kF3YYLtGWyisqNJ6t0TPC+0apfkbrYv
9FaQzAx6A0RC7j5EhacnvcKGHIma1acGHH1zcqBN5RN4Shb/NfLdtSx6SxyOvrGH
FHnWOk/cDoYjFf4qnMRdN72BxKNMkxvMrw7SVoo/LnXNseWPcbaA0od9OuDRopUs
8B0zAQhGKMhPMD6AotggUytSysMnkChaiBdrnHWvZd/eT2pfYzG/cytHD8EOkc40
cHwn456Fz0SgOJiTFtdmiA/okRURX34gAh2WHmCY8HD153bRlWVOEsY6d+ujW+uL
t9J96er2MAJV/pOUDzewTIq1TibdKm246BPOY0I3HLg9ht9UahH7R3Hz+h5ePUXR
/7CHb9Ny4T9h74mQcrandrz+6RPngkhIV2/UoJzLMbkSZ+xivItoSmtyhAgNrBZk
eQE7yS6SGypv4SXzuOq9U34X6NKjoeRVVZdNUbLAtKCxvTvNgWK5/BxfX9zzyfG0
OQw952AbwcFM2ugGsNDuZ+X9FhH5EiDUScnY+ZwLd/NoU4Wh2gQWJFxN9joubefM
/YtO651iukEztNwdvu/OJNnJkKrN6eg7c8lImfzhoy2agmlakjaNxsbFU1Lb04x4
Pu9TMF6C84gm6o3zWE5vF6qVYFX6TKmegE6qAacnB6U8PS4WVYYe3b7l+nI1YrY/
G3rCZ+d2UCiiksYDymtrwOXQ1Rv7gcKustNP1y+41ZlwG4oes0eo5SXqAscE7NuM
99x8BVlxux95uQuBxFWemJRWzVQgFMLvZHjyEoULrpsbqi+pB13aKrHVJog5rZ4L
BkynWq7+8Mopt2m5ZQqe5txHL9HaHoKrIqyTGeG0N2GS1KO43QoN8VYSiO1Yb5DU
k/LAyaqT+Bl9nQicwSsJIEFlwaLJ3m2+fcM/MAfXgn8U2aObityEQR6Jyb6/E81i
SoU2bEtajuS3R5WRGX7Dht0Cy/zihCBk3ww6dJ1xE+4BDKWui9FNkENVXqp02ekb
k42sMMIG0eStsZ4JPwr/6d6BlP5tp6BFque7Ksv68NJRhpYTm3BG/JS5PawwIOwi
YAGEZsXAwlfNIlZNk1k+mdDxOtTSI/dOvvtn/7RYZrhGgjrpANvQouL/evTDrWcE
inJS1eAzBTiqGcyTKk33gsE9bqqsAY6PluzGkTEWn3VMrmhZSF4fD6YNsvoeVPLO
p3pVD3ZETZWLBJwpPHeQ5o0HaTziiR9UycELdmOarSr0hs2ryAN42/GtMNbzktje
sDovavOxVT2H9xCCvBDSYKuxVezbX6LYmtfLx0IaKKheVhAnEy+LHXwWrdkem748
qub00xEe99/M/jdLKLShyuG6HyZRYTEvRKH75MuyhTGVkkPtDU9K5O3t+jRVjYjd
XcrZ8GcLO2uBiMfMfj/dpZC2LMJ0UkFKXVsGIO+pv0ZL6ndUaROFf8pL0E9YS03J
CdpsGRb+EgKj9p8FCpavQYqkh62SCGrUZWPU//K91hn0v0azx/QdeIhoxbFZBn47
YsDBUOJQDWbk/kuIN+dRr/wG3gfwsz7swPo8iAkrABM2rbiwNsK+VeRXCc5esQab
MXxZdZ5B5hm7J7G2E2uCL0CE7SJ48JHFFIo3OL3gpmLeE3xd3Rd+bmo71p/AWuuO
nM1WlhXnED50rYQgEpzBtGxHYOB0lBioDCSG4x8eX2KGSeTfwzq3FWrmObJyLpjQ
2NrerYKfv9V5Lha2l9LL2S2l752mpUAw9pzTYoq7HnV+WbquYgP0a1nQ43W1Y4qy
aHexFCW1XGHBelexCgiDLXqvfSKrUSWkfCLBSlV+04Qooh7AtPwryHFrmkBTFiXm
vfxJkhgVTSmmTUIfzzFr2bXzYJYFplnbmV9OrwXnYpIUfXv3YLqyLQEomZXgmU0/
vD+pLDMswrgTZR8Igj7ak6A3BR9oaQUz3oy3kt/PR4P7kpxVXoFkoZPEPR3YPQ+i
HT4uV39QWa5andLNtD7pdNrbgrGMLre4xnknbuU9TxmDKgn93E4pj+3HRZ5OkpUK
ogN/tZA+MwhSjD2nigFeeEM0G6qPsWHPknvEVKBHlaz4apOhKZY4Jm5a+JwlQbKa
/1dNsRk70vSH0pbekPzwx/tIhVsE/RWwR8nmPyWMB7ePOKdGoBZv6e1WHb5a9SI+
x+7K8s3qt0myDLByxK2EdkMkAJ0Tibnmx6aUDvI1PuzI3HH9K/eWxbrvpdVp3/9x
ApJJ6xzs5gdDZK49Q0NgWzEyPI1h2ZGqqVPsNMWvGVH8doZHIK1CH5UO9LRpPSB1
upnWy9EpEDD/ImaRVTTD5RmeSUKlzWJ9e1eSzSq5Z6cADWci8ZUw4rQxQ4cIhDpe
/VUO9r3KHt5JXCEAMFTYI06RIUVXJio+m7QPoQ2abDgjoZLpK1ScJ23cZipVrzPd
SinojwJR1t59EqVt7Fkcdnx0vfAZdxzsNwePOgZARHkeSgPJwjQhOfQtDAueuRIr
Z4bbZddl4OUkSWrtsvjj+KdIYfoHXM0N9PExUvLLazkgmnr+1RvFHZXHCM6wRGnv
3A6XZCttF8+KLEKcVPc2Im5Dfq5KOHr3AtSTyQ0sX+Dz/VVilcD9vNMyRlBCYhnP
HSMLtgsQKvEyOieS7oYY5QrdTKDa0espdNK0LThIRBaK9kLVV9Sksg5PMuapi4um
vZbadjZLBp0TSvMfroI1SDhPDWuh7nK90sDTbE9RErBjZoKjOyMWNOs5JF3Swza+
sV6jNOXoUxWeb9PDP+l4x8xRTVrdJhnzBArMre3fVKNn1NDDuZwKkb+dv6loMzGi
A6QFq6yhr9G/WkU6ETD4fyBNwm2HIpF2KYcfaJvHMbiEcKQ8C4FHhbsf9f/Ud/hH
lUvHrLk5DYA1jrm+bcozHdbTZj5ujU9icrRKK5vXz6en8srs51L0RkX9ClXE3Jlj
H+OWplskaFyichcvkBDCybntQkAs9lu0BpmIV6lBu3sW2U/Iv1Qembi2gaOiGlkp
C5VEtAmuGhg6IEQqdAggpFGOsuMWMId5eSEx+mWkLKXtbf7Etw/5BOMzF2EbLxgL
rQLrSuJTlW+3TixXHbdUsRqpJHoD67hG+VD4LvbAJq4tgQdNx40GO48O8z7Mi8dw
w6BX+cq71lV/i7etCgM49Y3KonrSAnJsaU4gFrpiw95Z85BeI8fo64IuJM3/+O7j
rH8shPS2Xrih4ADDmnoIVPutM5B68YaOx/Vz+Xxqu+hteJpCCHHm1uTHC7in4WF8
feyhBkRbmrGB45t+pLrJWT4qOcukyo01jX6s2qIBKZ8vgGv5GrYDAJH7pwvI9V/n
U6UEDZ/SJnSGZYwnOElXTPKwAbK2SikJZgh6HY6jtxNbzZseCB9VeLgG9LdwpeUH
hizK9KQpMyevl5womU9Llksajpt6i1V3SaKchZg23gDvnriwHgCItlIB3polwP4m
QhJ8IWEoE7ylNhGtgmOmOg3p2P/SD8L+ZsMRjKv+LC5XXFM1REDDC/1nzotgb/dl
yEEioYdLj91/QcMBmQxiw23pT1YIJZJvvLwStUYJmYn4Mb5C7JnA3ufmf7+c17Kp
WWTufeKVKxTn+vMDNE+uNyzx2pemsRflN8bHgEH3hGCSuDZoPHGso0+/1CbNXzuB
udQgPSWdKUP3AjESFPgYCXnFT+xWQEFN4OBGJQ3K8XpQLj8i8lAuQQ/7+JU922Jd
+gknBPv/Bbk77oZoENNLFZIagUBLxPNfxIeCDKI/3PrqYVc7/HlNT/bGPPWBY1lC
tnCShp4Hx5/0ZnF8GRoubiIBjGUC/DRUyVmN6vi8eWfa7HQ+QUvdOhjxCe5z62y3
iVoKY3N8kh5LBU24qz7KHthG4GbrELtL4EqQekbuYcFMGfQu4it2pp8PGkUStRdo
uixHsIhBs9HVTYNJ2GloskDgVCOXoA6k+bjS0bi8mrvjZ/w7/YpFPR4YKeNzetaS
ZSEqi7JNVAL5SZg9N3u2hOiOjZr269Em+DpLYRzGqSZ3Q9S8YWYy4bm6uBx1IMMi
z6pbDLhkRRX46sRlQvrzSFXkOZzTVa4HVLQRLdbob/bEXdYDpriWeOBOHB0Fp9aQ
l0u9S5C1maWaVoLy4l/wCPUgakBnOTOr1bwMREEowg4J8rkQJgcI6veGhVPTViIA
lTD8aT3P5AI2XQNckRiVuWpL8eV/4KUmXinFj/fGrVoSie1k7EabmKB8Yw2sH7hT
zmhG4cq+obLiAqmjHQuVZ4tqayhRA8BWaL9cdCsgMWu7MhRdQuEOGmXAKGx5gSjC
HXGFb/Hwpl9jQBFg4SXEcYjtS5UycnaFyUSPi7W4KnvckSz+gM9jQ9QGB/rTAzHH
khFYsCj7sfvT1b0Nyk6PjoSsSF9/vjanOg/kVB+/rBu5/1bqMtq+unTM9PtK25Hr
4TE9LCbabxvvGn/L++EqtNJ+ecruvy9CtHasXPxb+gc1xgFoBOZavTvvq2EjvHYS
UPuNHX5oSbSdmrOla4VzpAUIPRO+vffo3RC6CR5X+KWtAc0UxKDnrLqGGz+UMziY
KDZKQA/Td5vsgtAGiQrlcDGdA/eRsmHRWTFeZsAunL2k7haqigKg4rmUp3H9p2ga
LaKzB2/r8wxmRwg8FfbH0QsAdKxNX7HgoEDr/+BmnW/JnVhzmhbQEiXZTAIqODyT
bzZjZRQfEJvOLFcdUskW6MhMH7oHuBXsqtRbkG7LGfYqTsowxCHHEP6a6qEwC7pq
ynLKyicI7JKFLZYuFPlf+rERbumDtRIqPrRhvIV6R59AhE7PlExmBQMYmj4H0oog
IWV66Y+SHTFOBv3F+vR6biDE7F/WKAnD0PGrH/2viyD1ArCA3ypBUfab7usmuChW
QIpeJAR/Z2IZlkS2KJ8zVOLTShjy0iQ9+MHma5zVQmbte4K27MdVP7HtkNWFi05b
Sv4DVWGpOwsjmLuAV/Bcl1SJeaVRsQ5MkjGbOB+8MFqWdqfQ66VBJbxDdbf9vX1T
HCLpa60Flc9yi9WX6vmXpbtKHzwikyTp35bHsjFqWTT96qwFkCue0jyOVHB7SJ3v
anm+Bdqm+TDqdT/88ThYdMlZwZ6lKQhXxLWCuvHC6pOGmCnX77zvXec1y85pE/2U
dwl/8cXfZrx2xMSH0zOV1W7XGiHFn8QRoIbwnmDLCWGuenqn8JIEO7O83PogQS11
NGkK8IZZDTddG+qPnUvEHolkqgsmE89cbOuRb4Pm9KibSmDQMTO1LA2+HBl9csH+
Dmobm2h0o+cL0oS3nu2BySvVXzq73AeuPP++V694cu6INE4j9Ib6EwIAtzgeTWM8
ydC1aF8v3yFD02C3nalQKW2cj/YTR0d5cNKtJ9IRppTGhJNeaSSbk+YFyrwOD29l
tuCIXiIzOOSChQDJkAUdGq1W7fPrltzQUHjeViesa+1sB535RMZmlM3nwX/bxhvF
SQCAA06hvP8+UBLCyby1rUXwlQQA7SklT1jmK+/mwGChyZxY9ugzDzGAVE6JYrnG
xhtANvYdbSAq6ukvzcspsc7kg8B5A3sN48L+Ludfg1pjzfWFo7QMitW7t/kqetKt
SMfIKlYwcngmTN6/RrfDAeeatomkSPrPZjPJ9h1VwEgDP9OehaQ6iOsM2ONHVVZo
uoA+BPOws78H8NXGVfTPGZG9u0eg1K/smMS1/BZmIlUt5xaXahoOcXedfZ2dQ0Pz
53z2GTd7tvKlRZrBGofVl80nKKB46tDk6qI6KmzpRvacff43BOKPIopwl2k/bV9N
UzPAdoz5qse69KyWqMpOVaNnv42O1cuOHt4Z+zJcs5qODYE+f1VYYMYnpyWKRoSK
0RCEA/nYAYHFm8yL5zoI0lXyQEpDU0lWfv361mCnDHMJnuIr4jtSx4tJ3iCxsGy5
QE+673CAnQtsXtZBsr7OPWEeVhZzsBoY+o0viwwhDIZ+umOVKeMZfNjasfgXzWHK
82EpUxv51pyhv0BzoggTAXJboiwsPuCVgZo0h3SMgYgYesUQQ57+SlJ5Xy2c6C3s
wcf8LBjkkVqbiYmEBL23XRvhu7S8LzTKHtNR5p0Wh8UqevprKdTIPuL7zc5xDn7N
JTvF5/clfSrx9bsFDw54Tk6Fa+BjlY6PjvLSpvS7HJF+WlvL2V/cTRsvK5bNaT/w
Y0faUsXXsNVIdBGpjTF47ZDa1Ut4B22CX9qmwvdnWAxFuML8k7aRQEWc3Fs0Iabm
z61/JXnVaTlpi/S2St/+3mvxl3EVhbl8lYtrhc3BwLbD9rLfdAYnT25Xi52a8GLr
6ladQs1G3tXYo3ejifiOniZJTMVZ/CdmuiaTsIiMgKjoTtppDGz7cVaf72G6T2av
MEYQNoiWgrVJ4jXvAQm7aTnJa1lfEWAaOSquY3YcRJMUeC2/0YgcuyxQSD8iJ5yy
t5ieA3IStOuAYtuAlR9cLLGHqFhMtgMfrK2LeAZ7oCPw+9yVbRwdZ9lYXKVFY03B
LluGR8yg4K1AbYtaW5Srkwy6HsBgGVpg2Vfxp+3Q2FwCYHQOAGVlfSHKlQx4AExu
pdeAnysYJ/niFpN97IkKbO2x9Jdz6U7V7jPLX4I1OiEfqJE3CpPP5ibFB06OQ8rK
OL5sfXIVgeIqoX0MfF9Mb/v/2LepO1XXzqGwimjTLl43sFGoMl0m4e9zHtwyfD2b
fGDuVm4OL+M0XJDsdISci/5Syc5lfupc5JDtZAOn7FFqnGSOH70zcLvG42u+kLQ2
Nk9zBcZFI9eXBSU24pi+Hzfvtki+Q9TItHVR4zlviZKdPe+Y5nsS68eTOfx3Bb5o
YdGX2H2kJscUfNGNw+C7fOz3joli+Dsbo/cEG+2Hl9qi0YtTcp7g1cLNlFRtQl+u
Cl/A+e+ZagxcUifqpjWAVfc0XABBHu5eSh2zqvX/mdY9/ZURhVNUkiIGGaNtWSBr
DDDYPcsOkFb+es83HN7Wcjs0SzLi658LxwqCeRzD8b7YXghfZ/0CF794eoBEr2Jw
7oxAhqbNtMHRYYCANpig8iwdRK2YbVCwmuzvNr1PsZwMFMN+cfVKf84O7Q+epaAs
NVva3at1yE5DyjjeNyI40jUbIpK/GLpChBOsFa4l8ACGoU5NZCjHyFJvbuH7Vr83
CTTGcCQ+oX/pIutUSh8qLKETz9YTkDEE/6AsT4vr+6Q4Ec4/xwGJZJhoqmKoP36B
R1UBGT3Oe6zCVWnArNZECqB+R9DrBLT8OisxRZJJXMd2lUd9VkGopVs3sasYl0bv
LX6ELkbHSf8eyQ4b51SRe1F7ssImsfHX/NVArOlEBnYFkEo+FipDy6Up5szOPQ4M
EmG783tyVW0/v5mxQ0hEDLgtwvywSOUFIaljE8znGtAgy8TTFHpwfYrytC2narxL
EXzZOoL9hU1+yd2jzLvF4xcXowbg8bC4Eq43o8qZUbPVAKfF3mb4+FmTrryMqYzF
ikfOtT1A8WUCmCYpwhd8Ux0RiK2TeDHji7ymDy1U7o7tzGrBfSNeIrjj7ghQK0zZ
nCN6vWtAvsqxrQtLT9+h7u6vgNOzHbU1aIyMJYg44z0A+o4Pb5Aa4y0FTpGKotUp
GignQQY/F0aHeMjaxRsw2nfBkqTQmQH2Ta7nqWOHWtFkJCmLxHa/n9aqrJTOHYTr
hX0VxUoz+p+MVbstkK9fqwJGRNno4UV3YTxlSv1g9INJIl8QI+satv6V4zk8YlZ4
QOx854SdPJ+TKLI2jODxhLKzoJ9UKGhZNlPemUQ2TuhOQ4FoZ847wy7a/ItaGq4H
YC2HHRNc3vgMAhyc2kWZ1VHKtduL6xz289cYz1s1bclAhWe8M26JVNR8Z9i9ZvF8
wgOEaCGAiw3I5cg/Qb8Xt7FRz1Tt4wcO6D17ETECtyBlVxhARbCQaj1nKsvYdBrl
WNqzM6+NCISCMJYNn8BscFk3bG+dk+JhSOmJa9rhev0/CKRKfRgCYSrmngH4PaDw
a8BsYVtLS+CyW+mYxLASL/eDNLeWOVXdP+ZU5g0Ii0FOqSvK2cHOEvhfzvoK4aNG
sn4X0BbD2R9M7TVr2FYolCIcQrmsz6eruHYvKwWg6s4GURoVP2rp7eADomTIpGrH
z2k5NvUYusR6L+/eKoTS5xLV0wO/wibV8MSg1a2M6fdP6kMPlKurMJg0ncAhbLl5
Yf9ACZGxasIc4zC1XmM/0CFiAH4QnkwDgwluyf5Z6gAWr/KSWD8y/yel/AZ1erf+
11dScp3S73X9GIGlWioHyigzNCxaH/povOTUEYASnV7VaemxzrB39L5OH6OLcm/O
v1tp11ZZk838Vb3h8Mm2rPEV96nyRTV/xBTH4ePN5OlwkDSv+VQgxHZJgYc86Zzj
pouqmNfK1pprwTa+wyCfU8HV7uairT46snJN4qdSewt/DLTessO4vpHXrtzqSV1V
nY+4TtW/3ihzD8eRaP0Uxk0fDsxnP+wLKl40FqOjnT4kNqba7CYhySJQRAYQ2PcH
9YIpZ+KUGFE4CpFtfVGrbmTWo8VfjtI5sApt/xdcaO+Wdg5U0A2dnpN6VDrnI/L4
aQ3HNE6hhmWrqpKKGHqPSEa4ElhJ58hAVG17J/Gy5v99rNsbVHbaytvqb7xp48Qh
mY7K+wsNNrGM1wKAQSxHwXO9XWVsgNcJVZRAtn0qdH8cGtE8aLX2Yb2PmrM9g9NN
XndkefQrfX5JCVE0GcMNVBM6zG4VB7+pfncxbbWIYhD1ZEjA61qv/GNDV5yHnvL2
dWXXzcCzrtzW0mk5onmHfHELDAp9d7YAy0PRc+16n6mYHWBkjo9xsLzRD3LvDezA
KdwhErGxtlGmTui/7lh5dc+6hg7n89BRDv1Z9TdgK72EjpvElpBWjinmuhkFAV3o
5s6YBbL9rWQpdquRi7dYfXBAqCLLRHNQZCCaK2LXz7plFD0M7pcKifUqLM6tTv5G
2D5sohta6GEA8fEACL9a0/doOMUPv5id6U1tdORUM+VWGjISEzDeG1jDVKFrJsB3
AbAKiuN10MMSxso0CwuMjW2GpvU0HbX0JSAralU3oDYyDb9nGoJGd2R03cKFGK8s
lYKIc6hitzbOFZfAThz8XzhDRCCkd5vou6vQQW5Qwk6kAM8ZysUnZa4+bEeU+CdT
dfApGQRscrGRKu/ioatc9dp2uWO0XkSBb3VKlNZFRR2a79zcHGllMEVaX5bseyE9
T3ZTAoVxR6T+/G8GUk8lxZfZJT+l9DmB55unbICUiZWSnYQ1UdLwiJFZMNDWYfIm
r8YCguGy6YTHcTlUCuT3/wccJXU6UCa74m77emqmOEPyRM88z4cUwD5sjajmRrpK
/tQXRZgRadM9sRxslDH/HWdsLQH9lyJFlUzUvnpPvWa7qfWDMBafJq3Y+U2zsNuB
/d6gubSuJ2vXf839yG8VHhPQHkC1BnVz+ZVYiZ3671hTNybuU6/VbDslmXnQZyI/
7RLmz+vgNFk+qGfMckMCmKxvexqq0+sYlVLQEm0FNlFj8OBQBRzQk+qt5ky+x3xu
OQaW/X5Su8olkvVgUmkJo247ys9DwZp2R7gsB2wORgLms6CVE8UMM2X4fzuweODY
i+GvxBYS/nlz5jHC+qcgHZaLnhbyZWT7qUVa4ypF3U5RQuqz63mQC8N9BU0oNSGH
w27dgoS2rX9BOp+ZoxVY6kVHvYFbbYotHeZYxqX/DOopWUhCHOWXx1LhVnXzlHvX
ddcT7V/s2B+GNTVaS54dqJmNB537QtKHx8tTweCGX3AlxdVCacxlK12CYG6p5fbw
LlINNes2qFetwPmFzqjp1QC4PkZIBUTo7KQgSIjVX/IfxGnecJPTc7UYaFU2QL/O
PuJ4SS1Gz0FJ/nayrk5bSp8At+Cj/aF0/jPfrrn9l7xab+QN2xjH1/sLnAkNXE/z
lEz+UOJUCdQoOwjPWDcmobksGf7g4wX1IZd6kJMaPoUR13Pzs/I3JOPbniC0tR6B
daekteD23478VA7JJHxkKigutdywwI+VrYJ/TZSlNs6awQzmFOIHNB6/RrKvfYWc
lxWRXx1P8cFBosa57o7qyCK6O+lzp3mfZqMnuRbB0j9QRqoNdkFn3OPB6VaEP8wS
55jkRYsZroOi+XEpoyOvst0MgIvYN9GHsuBNPHGZgxf5oSjjBNcMNheLJhRLzG+X
TGI76l3U2XIrgalsIUgHqJvbq/cS9n5WllRjf5ewlqzmeTJ37IGnslMSJ9+bh6I4
EyeFimd3TEK0/q2eHrHYa7f6S9OONpoLcpVwxOdlgKUfGY9iOi3lluxpjFijvYdM
ZhXEujZbyvYqQq/UN/3sDA17g/CIfSloN6cFn0ifXMUAlFkZHEkyRB2sQuHVMVnB
ZI8NJBgGIzsjB+Nw17Koassn8kELsAhvoa68qwZ0tBf+w3OoYcLEGlqwDBycMqJk
ejsRaoI15v923b0Wz0yGynGuDmJrSLZOAhpU5NT/O4qothDgcq5IJQSqAryuN6zT
ISibyccAsx9NUFInoX0PB7T1NnE1knThP0NT+j3IzjhBB2JgaK9PmLRNb/eiPg2M
vWQbbG1F+tR+rQd9CQEUfysM2zjbULfj6+a5csxvBd0Sv+qbwR887/f3+PUpqfSl
DKwepCS2pWNY6XXw+4bKUw9RBCTyiTMw+cfPk97teF4/cvOXJ+K35c7iZ4KUl3rc
QTfDUL9LofgtwBMTDZn0cstxgINKCw6RDcp7sDKdxOtCKxBb91iMGNhsS0bcFdjb
skcMl/wSkBqFXQxNe2ML1C4KXe3pJkY17IIUOqYJJRx1PngzgmYRzZl/g6m1GOfW
ioFPfOHj74FPeMJObsbK9k+Drxj4lmlYxLBz57PRm+zl0M/IV599GtJz1D3yqxxD
Rz2Pa3ruS/hgIgqoJIk/EnL1WI78bVTW+gUG1vlY8DaKVRhjyFJjj3WzImnFJKqq
RddEqk1Xzj1DmXumvMw3sghplfc36nC2iPhSB43ptJvzPQ7l2wu/u13pOOCqUDKs
aZ+5NlyWe2PSaE9FXGG0h9OB+fuvcF4nChTXmDlGK4SvuJ9bOSYTfkll0t3WRIV3
FQG1JGN1iilBN78MoZJTbuEfGFMBZrCzKdcjTtv6R+YGEW+DCO4AEb/5Dwpy9RGp
YmYFjbhsv4+mwoq+1yBbO6yQSrouUvHnwMiOVvdur7Ab2e2YedKqImWBmWtLW8r+
fZpiA/uwiDuRZLAVwjTlPZROdLzx1j7c2qVZa9xFamAscZ50wYPh4CoEpGAwZ2cq
eyH45OaqrgIr5n38zSJZ5nR6urjIAZesTkCi9XMnQdGQ0Nc6G3kph7u4ALbMX3Jj
eG4prU06qJuSlZjDvbiZAJz1rBSB6P2RpAN8yaOTRb946wBq5JrXR7CzLguU5+y+
2pZpAle5g/5hlgW0/rDf8u0N7211dkUVfBH03ORgwlX4wMbDDBnZ18/PgKTrdehy
lVRs0TB86KsKYkSezqWLdF5fcUjrosY1IBpvA+IGcta5Io3Qdz2nYDufWBW/mClD
Lxqs2ZPg1FcIwV38TjQJ8c2Mt04tm9thvJSUjjpYgpZ8iCQa9hPnlbvTgxUPSCgI
XWckq2I6XL+ljjjaXMHJI2NbwfgilvAiJ5bmJkwQubzuVMA2urb7+SL/cdwsqExU
Z1u0p35fefZcm/7UPWx/tRoQNtuH1bf1LuaRhtugHYjQ1sa+wL011+x0U4lMcRUS
Bj6/JaDBxvnBoNXm1t1gXVfrpuysEx6+PqK8DtmuwVawdulrTvb0SK689ZZUkBvB
49IQ3F+pCuj4geftmfTHeOPgatdOQK5tCT05NYgghyh8fr68T9VNKAPgdneHfGob
5NBf17UcyjW8wNqY/9T9O39Fn5djOMfvcmSGNuO7KXYBw0pjfIYkqWgj0zSynsP7
Jj7oICkPH92OXTPubVzOLEoJV0g2CIsqDnyJrPiT6PDVVclynr1UkuFdCXHY/ifV
7poFq/C8Og8d2Fk0y1LmOiu4V0Oz/N52pENezv5ymqz7g4ifGHXYtaSa0NM5FYQM
2cVdhM6V/R0lW1LWDbuAq1ggDWJky+rSWgMhQjWKlsngzCDhaE/Rs2aYjEuZEwMG
7K9it0dwTCYXSwZ0lH77EgJ596907OFiZNQnhNCa8oQVten0vQItvFnb9s+XXHOj
R63jrqui4dxO+M3k/4JZIm1lQ+rcJlII9JdxfnhMqNsFSDIrQDx3D0boTBIg4uWm
clk++MrLVu2omD1oJnOjsUW8hFjxQ1RrQt7c06/gmIlU1JuhywAgROAoP0GlxF8J
oY9cdVsTmPL/0xe5gAOMW5fKyAgZY+SInqOFzcg2xG/bOSB/5lHe4/jp5AQJWl0H
mReknMU7RjaNqnq0+2wKQ7M+In5ew7y7w5qwld4F0sGO4NMxbIoYcULqOWotGKRl
kqOkU8lUgeN05CWKkwaoT/hIjbRRqlWSrIn6hbOs0Be3FqAIRsMhkNanlXIUbg7S
zmracFoGy4FQvfBIGOq1qvYaLlI/v/bz1nPi8rKzl5tC89bfW1s3/vA7nQETPAhK
J3NLpW3Nuua0Q8zq0BjnQAtyBZOrqqrUDvhmhMcS4i0ZLQb62aWiUL96GvTUJlNM
w82eAJnMH1EIcGhrsQtMZvAiGmG8VxfS14qHBeQYUIr2tiOIadVe+wJmZgRJHrOk
kQm690hzadb7Wpec+GbOk5har+a5LoMnomSwv0LO+M0hDhWitMGz1C28F6sHaf63
awkEE1bACXOYeUc6B9adzlGOTkdAzGQXqrMHH90ecJ/nJHOpgqmD86zUP11DVeOQ
hHkkAd+AeZKLHF+umyxc8D8k4gE3n58djoN2U2VsrPIdUpkEhqGtzIGdwj8i+Bmq
5oIMBmhaVdvD6kurvkLSMW1NhrbdMtbpeK9YBlMNW02qAYkCw4ZUYURbMHUS47J6
YxvW6EOihQ4LPVCXSIS+ANriShWzQOoag1Or23Vq2LlPE02ToENT4yZl2hrWDH09
wWAQYTljZ7MFIaNC0wjjnu3Yfw8rlUQgzRRUhOnalUiXRRjo7NPDmnUNAcGK/x15
icegBpMMt/Si3KhUOsCC52qaYPUBC9q7iFS3zVOyhl+QOgZs5BXAHh13pjU75J9r
44V6ONrQR62Mr3YwDlt1P8DlVsuvcIWrDLgmk7ePSmLR5i9CztfU06YINMfGvMUS
l+jKjRBcuPNHPNmKe24hbXLd4dDmRjNYB/fJTXC3i6hxLpEwPU9qsyqV/+pLxCnp
DhU9YAUTUAeubGWdpi3UL7iDn41j/oJ5oeCwc2JFoJ3GKM73G6HLy0AkC8eDTiot
P7cpqxrKllbNU6ep/Li+tLqo0EpJSXfQj+P2o/ZrimSv7jgJRKOVf5Z59AfjU5wR
IebLXVE6P7vADn10dmcCzhE2HNRqGb0Mb0ek8YiAVkOZzzhR7SQ8rH9OopsRgKhv
GyvGAI1FjbveT0YyA1g2UHUB+0fYJbtzivq/kZQK3yXqzyILtppgxmXOjKhCaTa/
heY81gmiNWZQzrL5Vxv/o1wnlZ9S9+OJBkh2TGHX/1e14ykg5OCKBtdt68xSXHqb
/KH3+QQcVsU8EeuRplXTOvPr7H4kUJ3mIcCPCHm+bhMG09ORRq3y/v0OC7xqhOaI
Pmbj7SjYvqQ6gh2bqnbqpu8lPyqMuplrcjLcMmeAjEcQIgndlBbsJck/ICouzyAY
LOgv53dmjyVFiJy50BG5Z1CiiadgQn+PCFpff8yO/t0Fegp9oSIXAO0lzURlXv/m
ZvIA32jr0fLzgQhhMcinqINK86ZC5GsaLsIOFEwagOUyqNsYEU5i7laamKytGtkB
yl8vVd3HlpWLvUjjUCiNbrQrhmzLG6TVL6fNzgnsDuE84PIE/RfwLmrxEQKMJGqw
Lt8xH772zZygsi7IWjVYPilBvuqcU8YMg4lhK+ILL6sOx+VGwqZw6o4Bsj5FFHab
J4BCN3FcbF+BP0UDssb4Z/RKMBoaxWQu20ceFy8CdapJS9+5bPRw0v8jL/IYCzHB
SyWRrRqfhyFrLIJZMc/sQXctKAMTJhi6yP0ktC2WViyJdOoKJMh/EGMFI6POB+q4
QVvtdMfNWLdN3Zf0EEcA/B2qWA91BG+Z7qheDwPycow+fkQfAJYGeiI26Zt5EOT/
iafQ4OJQMRH93kwaEVb6lrDQUeuT6AeIi8T8K0nz9MviAF03yqjl+OhWBT+WZCC4
lQtS7Lcwnv1cnzCuovyb6FXEAeVfXsts1yrv8GEt5eA7kMmAgv6FbPCegmDBWbcM
L0E12Xdu+muQU9TvAzo6m6m3MiY97N9C4kImq8xEutNHG/v2y2RCFgR/hLTAs/v5
DIRt4P2PpIHavqAgGnWzHnrTaltKqpE//eD4RDkMYYdJAcyCCdqyPnJuUrWiAMLM
cehh+/nD4ZSHnG7CG1maazgnESWEI49cAroRf5thMZLjX2YKrPnOYHTv2htE8nfH
93sSd9ycghGIn94OlqW90A1rO7GkqqDWjoYuYPBykPW6bUE5bgndy2NGMuecpXMH
a+4uqBnkn8NBKAZ4kEflR3h7aWqia5fzqjH2PZ34KIVGvIlOpDOwIuxxKYy7/Ub4
1pQ3HON8XpHJP9OMh32gT96E993uNVHClbU3ap9qQAjEMLsouNuTra62BOQKD7dl
u9+QIKGQ57PNuYBI6HdFdJ/Xw4EmIwYrCGtdjoz2CYBd+vuFhs7eE1Cpa9c9pcQA
UmdH1TA9jV+D9++QeTRxnIG3GMXlvnhkIfmQSxni5lQSGLH5zzMJV3NqqVwAnGxN
2A/QMn/UXFDsWRG17cXtgtJ69ZFadqllT88Y2mH7a2SRVpQjhIUZvSJtcH4FSQbD
3me77yWOPSZFa9kUrTiBnvuvMmdgRIVn1QKQ+zIpsjLb/wfv/26StJ/29zWiL69H
+zjmidEBb79q5xliTe8EnMuVspsNy//HvOthtC9ifq/Gv3YNRaSXNzt9PpBuaNbV
RYgq3MTysSOxWpwVxQy3Ct7dCKI+5f69WYud3zCtwMScbGKl+5sTwFHqYsgPnvX9
RGrFJaMJs3LI7GQ7JX5rRmpc7BF9qep7AL7iSEUhmAgTeBQYovYPsZW1vQS4JmUG
DobBdqhTd4ydtVABB61mstOm1Xnj9GsguXmakWrC+GqLpVmwU93ODJgBUptK4BML
cSDvNY0NPry83Thh1HBm7LsM2F02uioR1CEIqEEcIte8lBfov7cSf5u3P6/519vc
9k5T5sUMi+OmhESZ4QVQhN/gcXQ+2WS1N0lXs3H//FvC2fAKFXw3aM4LkftSmLdQ
vQQMaM06Kw/HxFTXAFRxOcMWM0LEl2QwCsvRimVBF1tyGC5vqc3/MeINqJTX7qb+
/yfOku6Jqyi5vFnIg3d0fPrp4DcqeoF8NzbEbly+zd/tD4Qd6sXyZYX6QwbAhgnH
eweJwcpqHiCDIRZ21omn8n8j8fuoPHRr+MDGtmr57kmYfCjBFs0VeCAiKtjAqMX8
HSfE7FfK4r91ExdoM1+YxRQyAis5QRTX8ayrcy1dkBQgqM+Ga2InYSC8rRRKdJVF
7xHXiDz4x7agyA69vqVgth8DD7Xwq6J2r1rsIuh5qP4sZ/I8uXRMehTGGTXvSA/H
S8vz/lGR6cJCj+Visic+mmToGPClKFMXam8AJTlQtH/b6gazMSpBW1nRr3Te+VsC
Rtl4Ip5DdaKnnWUdtzcQ1wGJuj9BD56nddcEDDDR4Qop453+F4DMfjbGZuoGjGLR
/hvDe2I0xpKg82NYTG1LW70leRaZuUm2B7f/aLFhbUASYYVCmE8lr8HCCPsvGwXr
0+UMcPYsJcxbIFYs3l29BLIQhOF0E/Zjg9YKUZuhpWYZselW3GrbB2hAnLz3BebH
f3wmA8Ymh3StV8QTwFBBcJ7clIJDaVN+aBElcRh0ai2lLfhJLxOCjKn07m+Gw8vs
ASf06tD54iTvlv7NJbU7w5HyB1ppvRKz6SbnGvgV3bZno0MZ/0Nfz2pichzBhknK
W+0cg2qwU6DeJyJBu9WYLLv7dAFP9NrCzaVEuCMyMczzmPsBBteVifemhisrz+Vp
hNAA4/+2hCRWEnBcpQrym+ENaQbfKI2OoEeUVhdXkkaYT3maV3giN1SDeB2y7pnA
BoXlN5P7hWzmuUyOKQDR+YrObQnXrR3sHEus/scoxi+zNyvrrsZJvmLaZZU/S/hd
m5PD3gk3UkCFIWscCxfbzbWmI7VY8mxAU0ZU678N5/9dSofl2st3+TIMZxgTDptO
POxlIG793uU8d6I08kA0trBwZYisrH1uvsPZ1dNGN/FPb5WYlxrhQTxXRXuvjrsl
wfBRZaCJlgH4MmJcTq0olBNudUwhZMlKryCM7QxqdualW8Yqdu1JqmBD4v6SOAv1
WGBJbnbj87B4QZtkDqVK0qD+AGNcOb3q6r0qjHiCrh0ny7PLqT5fyY4PKjIYYIUJ
+2JA6wqjY/ToWtkAKA5Z2qy12mzuurHPlxNCxMaPjc8FXWkbNnCyEgs1yT8/up0V
YE+DHFim7AROQUEhp8MnwR95jxgQeySJ/asuXLKmlAD1N05lbYueNfDdql/CIqeW
OL+iEL5bGSZAE49jZLkWHvjc1JMIBgQpnTbumEbUcE8keQDB9qyzxh1IILhxvzWH
8yFNTo23MgDWij22yLQzxER9DwbmcIGPeNzG0eNzxjwI0RlFLot1Q5OuYXhwIRVA
D4R+hwF1WPbGvWoMiV+BrQq2g9+Pzt+Hpjg+dZmnnemESWKGHb92G9ntoT7nd0rR
S9J5DyhSY1PfnulvP++AXEIqPj15jAOVPyCvfYh2lQvl4PwBL7LUZfTmEWEdjdM6
i+XQBjBVb8A2U4F6pjhA1c+pHIlgMjNahp91nr2RuD9pc2HL+/XVfAyBbEp8l2E5
wzifRrExwjJhIgFCAvXewbQrmulQssvhhJbYVu3j/mErz9vXgtBpdikVG2u3R0SX
sRYOflnZwqa/a2YrKBrf5z8QmE+ZXi5/B7Jm7Eik/Dp7M+xWFKgrz91KsD5Lig1c
VLpafupx8BY1QTW/XQ5LzJj0o64j99DnkayM1LZi5cr//KHkTgMR44yKlthBsAfN
+2FEkMulSQTX4yrTQNjwmkBHYYKeojI9EvWU4xOUDtGO2tew16RpoYDCynSu0Uj6
ifoLrbbyOmaX6zw4Cj2GjqWWPrfDNqGSuChQ7RbhPakz6TIk9AJjK3pNwHKeFyog
M7oSy7oUfWj8oKILjkHmGmAEwNCQHA86StWIsXzfNcb6yXoN4QN6mVMYes/1wv2O
YW47dCLdle1YP6Y2ho6EcR5v76dP86EkcVgFOevLQJUMpru5rlrI4E3uv0Ky2b0F
ojxKNi37UkTePTK8ymzMPBW1WIA/1OVVcDx0M+JZH6An0qjsUTxxjPE36aH+b3DJ
J0NgR4ahVvyDCHxHFcDwgm8tKOk3g5PxHsHQJKATPI3OJsx2uws5LfhF5HfJOl5l
cBoySkLQIq6D7MOil1wGcj3RlpNbeKlx4vyh1PT1H5p1WCJU/PAji9BFlq95OUbF
oic0ze8pllky9wzKtVN8WuFbeb8m82lWvJdHLnLdKd9vNqo8DQAKI60632EJGvWS
DcucZocZSvsy0Y644RRCdx2SnUCHMUVy59t+0B7JGoMiz4eYsByR+hbWpQ1X4yB4
IlVpKE8VyC36dHFcZIbNCkJZIjm3XSn4lJix5WldujLxcpBrZOv0wQ/ePTCaSFyz
hJFQ05BojrurhymDljhlYvuidCQV/HCW6UxRosbQQortB19kK5FEKH3kh0B51p4J
CIpGfIuDA/Kl//o/VJTiF1EqAybUCviZOc91/i0omKoJMXWf7RI+srtPS5szqZhm
QSoDBYH0g67kU6Dvs+bCmIDANdqEsB5gOmt3nnUOwws9gyeb6ZCtuHqfw2eRg6QN
gCZGX+gqyrgbtPqqOVAt5eT+ioM9InwJ+uhtie9LoqYeQH5RrYQ3DwW4BiFG/Ghq
bpGOkSbdqzKXLzsYsjiV0Aj3rP4WGNZHDp4RusK2cUNZfBVNseSDLsqB0bj/Rumr
JdLmHwlj0BCZ1Bf1vqYqm1H4hiyTpFevCyOixGhtj4Fc8JHwSr43YtLScqPafj3r
co+HzrWtRc1gx4EibuRpDYnxbdM3ZUj4QEx8bbYYsCFSWwL4fyZzJvqRXcGmLXk7
QndmPpy4jFjWnwRHEC6+iXAiCsRdlIwurmOBzdLaykRqe2P7lCq6w6gsfDf4pI+Z
5wNoTZTsKp1jXd4yoabD6RccopMsznPEqzJ8VEw8wbAqD74BraiE78rjs42vDsOM
78RcdyTsJHEbebYN5Q2EXd0j71EKb8fhIG05ONNVcoaaWvkEJem3osxk8Hrrn6Ks
Ffjn4Gq3nKAHT2SOmfRTh5XZi1RNaM1Ow9CTZoB/TanjCSPIXhSY6IogbQZ1vHW/
gN52Gmibpo98oKVaeKd1crcZTI1EN/EoihVkvgZ9Oj0RBRHR0RdFPWbxpefbVHfM
D6esM6ZVn/kutWzN7yomeJWVIwuHBjV3hhpmaZD6P6rSsx+MqBhYUg7pJSTd+dVt
+LymtHTawQWspG7vh5QA4FwunaZ4Ll9V+PdKb2U+QVBlcHNPhufLvg6pSWHxsqyX
UIooJejIvEy4uQQCHubah1JRpqO6ySs6KmW05F8Auc8r2lIkZRNz7e6ijQahYyp2
5hkSQjgZO2OKhgkNffk1YHsx85DVJP6vTBJ4DMbMijl9aGJgdXZDInsDkbWoUnJT
RqWH4InrlCDtvStTSb1j0TT4EzGidV4sNkuwY0f22g5KuiZ1pYi6lfa9+PhUnWJa
x+X+B2gBYzteS4feytG+9OMIo9jrO+4+Vbt9UHP+wO8sAlLZRFpSNN55JFGwfBEv
ZqNKy3MC+SU0OzKJwtDj2+QooL3xLhnTc6TN4QJ8WQcd7mHTmvVRanLmZLh44dvg
nCmLU1uZP5uJaARxNRK36BZI/PuoJNjf78j/HG5ieUqMCVBLGCqk1tdoQFNeBzOO
BvSq07wXcrj7y29gs5ckHbAT0t+xtiuJDUJ0SNCFA/YT7Xy65i5r1+0UtoiKuSC2
2Cjf/RQ0eRaZgDiRFBELkpDxnZlTQsK6PU/+YuWsx75KpG8n7tkxxq/Bd3b2Xf0j
qkN4dPgi1kYfVYUmes6c6bINgb5TI6AhoUWmCOZwLcDm0G+a6x+4BA1eS8kk49XC
9ApCy4ykYqKwz9iv7ohWYyeG6hxbvj/SO6ugoxdu5Nq9J80sCgwgO5wlE1cuUkln
LSjFQcO+tGMrungL44dVYKv8zVaU+eTPTzUe+I8yHqyemWgNcvUPLAGZ7hQ/LF6M
IT2fJwff0NKaO4u9tl69gsOjpPXhGeOiaiJw8ab4qykrc/4g3+xTgO89Go6LuaaR
6uBgfOc3ZbmKNmWL5fuS2TF/UfpeeNOBo4qKVslJeM03o6ls59qc/YXqudojxZXj
9GC4kiBBBlVND9JP4EZRFpBHvCQhTKX1gF0P5ku7KPLUdHNn+wvnKIclPJFmCBvl
POYEmXjtgod2j4EqKl/tX4noTDRztCZ78j1RacbJo+RD9yYGJV2MItRzu1cmzj30
EaFnaG+rb9/YRAuViKLJrJRq2uvWOo2/+xbXscDc/Yn0nJpn87HVNFMQA7M4fcu9
Y1KIOVX6ak5HUyKqpvZqjnz0KYLGYZnLN82L94ihRgAZKRb2zLu42tTT5WaE9LOn
9MYS8mpIx8wY2hqPRjvFxuGzrCDYrmvzFlRwUI832l0xPXtY9C6HmdBvS9DrHVjX
jdHiy9rXr6xRAUUhCisEFeGzACvSa9hQrehkPBkuy7CnrEx8gmx/0FGYo9mRNERg
iV4VbQq1P2M94J8529DZ01U3v2mXjWO3MRttlHl+d1KYTJQhuiIovDnNPCzdMaTU
NZYzuxxwybkGlkI+dVMQ4pTvunp0qE34jiz8VW8E5UsAe5l16C0s0yOpuqVFVLk5
JWj46i25ltSm7Uqg3Ce4A556bsLSx3oAho3S1LB49Ajt4SZ005RC6+xH7wHb5rC6
mcmMhjC7vyVnVlOgx4g07zdRsJognMfrfNsEXvk6xrzxI7RT7m6nmLFlCDhNOZBo
wo5g4P1E9ZR3jrcCxZSArdjgYuxj7bdbnjGVF8U8MTgzyFoFCKq0ie5dTC9drfAh
3FMsU2gk/rOCasQUh+bnn7BEvP9Tc/BK+zx5DHuo3VJcTOsMeN9+msaHMxqKiJIn
9Lu4zDkcbtK5qQ6nwmQTcPbx2QoJJtF3iT7zd5cXBWWrnZBGeAl14SL8tyLXj5ig
5z5DpNOExPMwCOYkgBMohj06C6p6hP7TCCc+67018fvwzBjvp4gGoWSB2eeCBbrQ
nfrT22hlljDwE2IWrp6jsgJWdSte0Zeoy8NJVSSSYwCexvQKbzenVH7q6vWnp4Ya
2VMcLqIDq/fh2m3cl6JXEnlPlgUWk0arV3M5dEp5SetRS5Bnhka9NR0OraQktp+g
mm8R//HQ6JEvl3fVIWxTLtW92yUNb6//R7l2J4hwzVzGb5QEyDeE3CV3uz5nmXC4
3HIUjl2tk24GUW8HCYSFzCjMWjhKx5pkXKAw8GsP2zzMbC5spA9K7Lv7DIpXWCSB
PPVZ+kZr+Ep5cuki7i8wVaynsiqDK1NYmzGHHI+S8pkf7q7XuVJHTrJ3HMCJtabR
hyRJrz6bfCgorVlmWW2iHM4Qr8Xxq+q0b31qDkCKvg7V+XBLII2733WiJVIPSXSu
QGtnMLrJ0ERBsy079IrBnUZkLdVWXSbFBxJTQ2/l1XWOUCh070MwwzycvuNL2x7W
hA0VJpcdCp6gN/eVs0s+WpuIssqB7QKNOhvfiad8HkniXyTLII3yrIgAV3IRyOsf
iBiRqjbgKdFZJnOGKry+0xKDuXTyqSHnhlxVSBVQQjKVpNirtUBiHXZg32AgaeNB
85VU9FG4BesCh8lNQDF5GGkUQhvoIq4zEhmO9oBjnq8RLZvaKy7aVmWk1eiIlpAD
BeDALSVVWxbUqwLXDcmvBITktXSx1cErKxcSJEnb6EhKKF4BeUNl5wEH+mJmbXu5
8q4Kh8YoJL3kNF5z+p6dausf8l4/6FVX75pCNAIHNqizYRjZk3gB47JdgW0VLx79
p/F3PFIPCvDBna1Vg1V0cxHB19z5VGhd+XLLxIgE2RSE0LVETft+ABNFvi91gd1A
Vt+sw+ZdDmahlgitcGQjEko4ou0n8Ic1elkVugrmgPdA3dAdB8a9c7PP/v6+1n/i
PiNVICXp36u2YMgn/sKy+4HQZSsomqFRRkFa+ng16vPHt+s2egBmvrHD79AfqzZg
o+bcD7YWF4TIQvmjYGpkEEACKnEuhFbzGnatoHfm0gDrJekWj7Z/6BcgRY7jLjxL
Mb2By1Etdt2kFykIyXzndvwyEveAtWWH/di7dgEbdjy0z8WBrheyL86T57Q+sD/U
YdL7bX1Z4nHM/gefZJ/oWZghFEZ6GnZuaFhqv2MxjpBAEtViV7jNqn4e9/c8OOVy
UQZzY76O+nXW+FMPvWrySDJTVGAZ9x1PtHHlCnV++xokqiu9L6lPTmsHczt8gJmJ
D2K+RFR44iz2hqPVdwh9stlEGbSfUvX3iksgojG4DEnDgGPUP3Hi7ny7ywhUGhJS
oOl57V4PI6W+oivqPzJIPuBFgyN4hDQsvcg/PCZhRMgU6sEnnSoPkruqeAVVle74
soGCzVIMe6i0Mhs3H+0CMVhw/9DkXpXjWw9YFcj8FN1AGFUY6GiZ5DSx1V0uarUc
ySp/xaSKkVoDD1/QkrBXTsaiefp8RTcXhY9Y0VIZB7s+vywEdohgQJ0rlIMInZ/V
+bh2FjVaAWYCtZ+nz5VOscJ1uXnlDbTgqiPBe122DwwWSkZM32zSUNRqihDq4qRd
uFDreqfQUgiuKjdG65fT/AnnWI/H7g+EBLb/McitJK4yoszAXVnAA2yyVKSMBKl/
0wV8dqAmDf7FZhR8iZsvyfj2ma4iFDWJV82NmSHu3kFQ9JRHe4EIv2FBlEvBgx4D
lLBWnpoDLR3ZqunhJBRSBmZx549VeTIbh7suOpIGIUGT2kixCZr51Nf0dt1KKbm/
Vj4s8ix+AMrvkCziZwcAsHlTW/xNQi8jLlQ1iv/91AxD+6I6PzN9S6p4jp/BYcW6
3SWpk8AZI46oT2NG2cSGGH29D9qTyzGHO9Nj0gwGccgE8bMNIuG373rRyoFWxQ6l
tAxjMp8CyIWWQN7P7wWymwvZJkNQEbzpylv3X4RDMR985tSAJeSq3ujpFrQWBpY8
Q8q2nqpdxqJ/+TDJ8LI4QuSgJxtptSKhYqsKHAVlSc6IT4GZAjx5KNMHiioI7Emy
Pz8L527p115a5k54JVkL+ayxqVFZ7oQ5C3Z73es/TUJijrjxT3MxKgztfuJT2C1P
sxTp6F1SOHPm/fkuZ092j+ZQuiPcQvoZoSgUelRkpMP0Wn9iUoi/m6EIjIXrOXwc
jayb1SqVUluR40nN38qGQZmRWwCEJ2kv02SPeNUezZHKdOYJycr7+dTzUCCfCGBa
WPdYoHCFH+BVT51y0/s6XBIMGeEndqYfRgoo2HOmdf7WJihpybLNPbENeo8HY5ku
nkJeTCWaqLqD8UrUgcQdybSP6cMsQTyEALtTxbcLZ6y+4CLXB5OSw8sb0bpvIu8H
mleDb6QzleaLtxM1aYULA+APFDRqKzmnIjDVvShZ2YL8cnisZSRPaAqzfVF0kAyK
wf0U+dAZifiLBIXuvqRLLeY/MDFOMLen5E/CI43rRuoKzuF1Ba0eW1HycXL6gtv8
U2fZnODlrgGzqi9UyshfKele0RNRA71qw2rJql1UczOTpitvO4N64GFtrUjQvLCm
22NsTmRo0cbKx6drTzYYl9lTZDR81hnxstzhpIEUPpJ2kkkPRU4QkmYMJlFl8hCi
pf+4StuWfJWkuWyYDM01OJfhg6buZxOphm01qEZT2tf0i4t04B17h4JxpmNfb022
U+f2XjzkD2KP9T9jViDIhzZvzrmOCm6uUKq3u3knAtZi3TyWYbObtS4DTqjE2qFw
g4jXmGQrdefLoHu+Q3WnUvP5k0hkche+0FETiSHKDPiDbrZmmbkp8mkQyci6jtU8
hQaTYuCWnK/jF77SM6z7UP7Tbi11yI5Lk/IDPrW0N6dg5zQPeKrgu3mlM+CFXHXo
w9d2pWdwbZxRgeIxTOjPm2chuA/QitGZmdhlYljhSk7WW9hfCsOyVkA832YHKa9F
SbNX+YN3S4gSiMLHNIqnwpyxVPuY6nOCdqKAJ3/hkhVeVsjSHWtrsnAWb2S3cH7T
gVQpJqsrP2pdWpCH8NchV++IEXiEv1PP0GEWQzugkbybzGMuadZJxuymgzGJgTnX
J9e4E3PumetAwMKK7/QpIatqWiMe/jucRnuKn9erZrxqroaOXlZ71QSp+2vy4+l2
JclBelZWzr12T74ZbKGHfABE90ly8dwRPQTgqvLyru6fWZ/WnaOMH3CSyc+kKVYS
CSK46uBZxzY6verPA3m+Vphw7rFZ3iOX6RVRLQ3XPHLHXhBrO55+Zdv3hTxT9Zdd
MDTg37oKZ4Dn2QBjhkvhGN4lD8gKh0Lu5cB9aayck8MidVNydmvziV+bVPf5FSzm
SCKwDQlfrjb27nEV9PHUAClsCTwtD4yqPVwklmf9u12q7kOqqzP5Bc2gBcmvn/b6
3uK8Avr75MN64Qn+TVrJ2BK4MTlieD8CtCkq/kkfOQj+DpHEeNJ/mBYyTHSj+h7U
QZ4NOC3X3KAXq4c8Vrk6mNs3YoGh7Cr03EV1TBgrA2mKIVISAPNVzP2sS5zp/J28
uEE1Sf7XtKk8IygpOQOAKNP8so2DQY0G19YI6JYCKMyUJadcTYHJtwzZF+FCv05y
YW0EIDEiE9kmZQg9mE3BOdvjgZowc6Tt/9cdwaDwSlskKTqf/IZjrruqpveN3hgK
Raj9IWZMGXpONzEtNH5gQ1EkLvzAQoNEliqtbeParxFdkTl9F98rnXP01paNejPC
kXLD5ry9VKanRt1d0Ico6GpBQcYQGY29XJYdM2y3TNwexa519VxOcP/1ovxyD32B
3o8LbtXT5OdeceVOz1VERhiwMAq2EJjBXYeWicJZrJjgdAvanHIxJpar3PXKqix5
G0D5dfffEHguzz+VJoMe+CvsmsFfCOV8b+3nsi3bMzRH76eKh86vTnR1XnO+VRck
jOJsoIbo6u2Uapi0FvN+zZka1nF//JVOnxzBDtvMfJiixOz37r19/gHJILKL+lAt
7N0kORKG9qxBG587FiRNWE7sYNHqXJhrsJy0S/soS/mgdlOCp/6NVS8rfvvddQMq
YqXqum0Almt84mFWnKy/xj5FS8qFKNeJdOs9ZIcjFL9M9XIzBOlxGWwePD5JXPuz
QYn0OWFfRA92kcTiWyiAyYUvWgqpl8XfF43LAxOM/7b7a0fl7iB4eaw5Ky+yVU+D
GphxMdS/smFHpC8/CFCM9twJ054iZZukdaS+LA4ZAcLhSS1oYO0ZR7IRqUs6j71q
6HeX8Ep701ogRYzPzI5Eh0chu2c/XV2OPDFGEol304weWc0PBGy4RI52IcfCw6dH
7rQT99YmN3KzD9cbdNIPOFfSeHGMXzz1ShdIJFwEO8r5c3dla8F0Em/DOzSoXt1v
aTz/+rvJZFRjGi3eBtF8BADAqi7+SB3Fi+NBDE+SN9T45Io0LB4k0JGLa1Dgzkfx
wtJQHxMXQYxjtme4JeQhHDYHNKzeB0Caaktuj89GZQybmrMzQy6aG1BisErq8Pme
rcTdRSwhHepDY+wkuY26DtVag03n0X/tPa0JuAiV5L9uOWWRtRuDz1So5Z5WEW1l
fw4Fg3JMxrNzPethWTLwNv0zpAnOXGIOodJY0SqOhMLOgkn/y4akPMVmkIkMJn+q
+M/kdkXOULjiB9/J2/fRvupeWtOAuDyU2twYZmtS4T31LvserepYtsGlnt1r5hro
nb1ng6adNUUJaRTeVSOgWXn0LpVSoxVRvkecy5+OeOC0j76euxvVEEhtbcu1mum1
/LLoPS+oGE5t9+ogOZquy+EE1FqNe/isAcT8O+gYXdp1voANhT61AFAVqhRUOaoF
6/gKYe1PEVSIte0+w6SGPXz69EMH/J13l+z2/vVsaE0yen0AsWSd3PZeQ5UO8+gn
0LdVQaG/ZImwOm4xqw5IXKISKMm6r8BApBlnOq5wiUn/h6cEBr88XL1qgqlVWiC3
YF2mzwZsizwt+jnzg2pK5o+RY5+Q6F2FZNmZeZoX50aU5Eah2ImupB3gUXjOtXME
CgQvCsDO2Xu0J9HkCZVjzNnwWdDXxiVTFIc2ZoII430Q2EwBXJCspj6eoG6e1c4U
JVAxH227NNbikkGw8BZGHFgvYE5yjjX4i2kvCFPNk/iJfe/vcbtXm8VtR5k4b4dD
EX1jePXMCVuGnBhV3OD98O4jtlBFYq7F8VlbLRcvTCx7ROT+2yzziJeH5lFnvDgh
72l2sK7wN/vqA059Wi+2lyRw2S+Dlzm+qFQz1TZ1qnlpg48Y5oJ1YFR2yp0O2gGo
7tAHPsEohZh+vEHLozEkcScEe4O79GVfbmBgEua1S6mNlzHEHgtsrVPQ5XAdG3pA
Fpo4aoERTbUyzhuGbiylvLFIH5bSzRfvbVo/843kHWQZwJKoWMZAZ0Y/YmB7zcXi
kxjZbtGYHG8uqufF9dCzv+1wDcl38OBJAYsvCMtjKurmeW0IonLRipjNGpfXn5Qs
RFHJ8lq6t7+t4PxJ/E8TvK/Jp1I++YffmvfUaURQhwkEJEY/kUzQgkAd55W4VMBI
hxG5LhZy7YFFtXwdcQFPSa8NilaYYcxC3sIKdh7HfmUNl6xs1mnIR4nbUmwxQ0hU
iSAP/by59FRu/8Rndn0dl0lTuQ/+Sl3jmDwbl6Wta2pN9Egm3hkgFafOxB3WfzLU
VwpgJiwPeSIXc57i9vu5gfmGeISMvBfPYPNubMCDIp1Rh1uFe+tGvmbolCKszGNa
/dLx1GW16hOQUMFk73nhAuofLvFO4SPJh1YsXVLsHYUM6ETF5T61uPJxBXETQ2W0
Jn7VSHRwq5+r1xtgdlmSdTC4UXmEKbb2mN2ALlp361RE/rbnfMh3QBO5ficTxQu5
pRg2gc+mOSy5Lft4OX7r+uDTb1XeVv6OVxnklXoAJESGsccoOkLeoNQBCv180y9h
K1b9R7O4FT/Mt9Wl7ISZiHfcC+HwBZMB3QsB8mwR4MKeaNUvyLdSbfe2/Lhd8IvW
w5njnuuIDvp83XHwAaYTyb7ypQbkFACH890FOgWOnc+JklITRcR8qY/zaiPLSxAi
eywCR8B6zeLbkI7gIk22olm8y3qINKWPXzWbvHoE/Hea9wkyzquYmYixNcNGPNgR
ob+ltepw1+8lnTeUk479xjxtmRJPlUPlUmMM2Lo/BSg7qjz136ELufyZwo4NrnN6
bqhASZsSuRhawTN4uKyFYGXprOeytdjRS43GAmioDG1xvgYAHGij0gLQZ/KCX6nc
3Y3/7dU3ZgeDLQCZUcKJ41/Q4fapuLYJnfpOHP5CCkCqFZkP7jcfigKoZdu69xal
lcdp8AGf7DqC2/pwhRRImyS/GYU1QexYOHcN05zOnaKEW/PRoOVhtFKoeSsHpdvY
h7EHOyoDKbvG7Rqr6qnMPoCMDwqBE5ydTIahQ34juCVaZPtEkYpqiuaAnzZSOc59
o9hzpITjo6R243cXImS0QnlBbm8NGaPnHtoq41Q8KKuY60PYaYRKw8T3Ew34ymvD
wIWlsEWC7szWkYxHAS/i7YNFfUXU8L/qtwmP8p8lkfdcogQioTzUq1shnPaVcO9p
EqI8+xgMh9sj5EAXdKPTPP2NtHBks3K6hOr4I9n2ZrpYT4VNDT2969fp3k+LnuW5
HSMkzmLcvj1pK78kXacMwUqnNvRinmfaEMS9ZbXRRGf84xSUG6R116RtUyH0VMIY
Xk/xxiQHSnlFucsXzw+ohWiwGqmnlMwoBC5FMYQTkOn17AB3dPyFf7hb9ixMj8fU
HNVhFoeGdFfSNlRJ8ggrG+tCb3FrKVW50+xTjGGG8K6geFLzNeoxbPX+qQTLeRi9
eCmOWp3OqiKmXKHVa5NWbxgy8ser+eWFXdb/BB73wejmHu5bMHge4muCiyWe/2E1
ZQRcQc3GvMjKLxd5Vjb+/Kd5yC93tJudwO985Ym2NxSFX2Uk00V8pvXNiDJjBWMl
g4G/FT+WcNNCqbJ8ne+bDDXZHkeaPJRoNHSSaDkMsC7IQ6jdcj0M49hjMpksrbcE
2z0BPqPzSpv6qLL0Yxc47DQfcyfTsFlssQYXJ+QjOWLArZbRnEvosgW2BmEXbohk
AQTqBfONpbJPb72cRHc0A4GZ6mHxzZJn8FbNAxiamTt5pRftQyeP3cH5Jj+1yC/M
4B+Tm68ghJhWrmeMAQelMAObvfah3XxBw3NumE/3g+Hc5ZzZQOxhPGL3asNAifVL
B53y43EIQTqC+20/ys47I0QWFSVS1Wkq9mtCTXjqiVrTd0FzORVIV+1DZezkSC4T
uYAqQCTs0IaujiOjIwulbeq6FrYYVzczUHe1xuQFkdYFP38Db0cV5PzTwkxQjjr4
czYQI3aVWciWqHCD8mWmsY/9BYvhUCp/CY134txxkARhjBeXteqEVJtFXPfEslhZ
3P6YrqpTWn4RAtNLO3OAASdW9YPe/VIJrz+66B3R8GFKitfqbRWMqX8cAetxdBQE
Pu0dCXj/XJcNkOlJBvRLrOJVPUEtCxU2D8TPUTepjTidQD9ddjoSOtNyEakz0M9k
nbA1Owxs3cNXmPZFbABX+IY8t4H1vJx9QgeKXuzk9RE8O5/abNidONfPt0d2CJhL
RR6jcOijEL0ak4UA7pkOIictaLw9ySgbKIfmMUUezrNWAmOD7oH6fEZp991YRkoH
jWmvXV2DuZQHkcqMPqi/dVPAqEp0gMxGzVnguZSDSl+EbT07mcH+iGkJecdsAlcD
69YCioY1CUpKCv0V08YPfZhK7yMg0FiregDxngQY8ZKd1xIIVba9olsmyFsQLxOw
0OnT6b8ukGPVnco7pxw9fRQj2/ZU9cZKxBFFh9rnMJsZyAX0ntGXANbL/V8RHXn0
o6l4quyAl+Uwlb+Tnk4qFIH0HfZq2uZYMqLmTigMSZPYbCCvymRCJd+3jkYDRTZ/
1VfPiRe5HT19pKRl9kOoj5PjV0UIZnXCcpHDYpTqRvyZAUQBgweeKbjQs2SeDgmk
ExHKz9+of6PsH2V4fsXnt+otfdir/d4dsOcbRRLWmp7D1Us0jbx9oABMGP36FTR8
9HFUv/dcwQRhzuRYG9+H4+/ZuF3JCqHBeN654Rdl6DvFLKSdOmQ9WtV3PWImEcYX
lpCu9NgHsrlT1Ly95ia7lfGDuuyTjugE2F6khM6U5pyKi7Tho4mV6gjTEM7DL1hv
otXjvRcAx+/vNL6eKRkusyiGCIyesnG+dVBYhUNwy4fy98FW9AeTS2zZRTtSPYZC
pknnVGYn//UdMaufFA76KbWzjgpiiRYM0D/WfHFR25ShJX/aVw1fZOBb/iQK/sDN
Tf7dB6pDKIQSuT/kem3HcfZ4uxxYjwxalR5h3nQSLv72GPftmz+3cxMzNBKWO9KN
ubsX821ejL5uUu7YwSeh/I5WzrlptVwU8q0KpM2X6eOH9/8gstRIBkYaKgTQls5S
sXn1YXFeoSOiTJ9Hw269n9Y1N0uLLAL0e+GFLETgmdQ/v8gXZtFFfcn2K+lZXfjy
olhxJS54Gt9TRsdh+WxGIUsbfLBM+hJHIXeiEBD9QYXvaV8Cj7ewL2ssFeJ5wN93
/nCfuYiPhYB74h6K+bviPVWNFhixPdaVIMBsyACL/GjHSYAuCxzFVXK0/Nv4hV20
KSTFY1Z+kokwJx4EcQ79YIPBH/9MAIRpOsfK8r+RMYfH5nMTNEt6LPxmli4wZ0TK
lL7R4snuInUlkBjE5SdZE91ubv1qJc/WpRwUedGz9qAk9cXMoQRX5KO0Zh4Azx1C
BFZGuXBWP/FREePgm7fDpFDCmK2/LiVEzWttmqhgdlw6bZQZ0Iw3KVzQo+jWP/jm
2W21p8oElURLC/YnkFfQPE2SRlRUFF0NykBM+TGxQHAnyOmNvlveuK+eg1I8L2OM
5clGYTzfFAFOEH7rKf1gx7ow0V7XjhH6n0+KT5bS775I4IOheC5z5+oTlmw/XmVU
iW5v/+RZ2o61f4AR3KQjl6ii7yhiQjsQvBsUoFESGPWjdou27Q1addfJK1XV8ZM8
atNPi8xZ3I0vk4zrkbgf38RY9/I+mi9SM7WFqf7P6/njLo1CCHYpK5iU6gUcqgro
d6zuv/JUnDJCKCPpsXm1Owlnf89ehKq5bIdiP1pevqcxYYrhct2Q8DMl6RwNah1S
yImvn+DDDBtLBoKShq/GVekgKHA72/bnUDCu6vUyW38Uby47d+p9ART6SRycc+yW
/M5EShnr+gu1l6W2718PdMCExmaD0aeUVWlGJR8pvm+XRezwuiRTmQPndVuI0BVJ
kWBPLU/yKZMdNd+ztWLhgeU5vkHEsu00b1b9dvoV0J5XglUZ7XXk5betaQbPiiEM
MFz/jXI+y5Ns7SuHxen/Gp2k0ok27zxrqQjjdbvjdRLdKNkVbscIDTCfLNwW63QJ
npphZvi4GMYRFYmLM+u0XpNZzEamb25FH74B2mDXgqGKxxN9RvCIfsYPETjStZCP
JtavFkJ5Kh7ocXbZ+G1EvOraMEhnLabCeuLhvuwKygRXthrBPPQ6n+nrZYtUaDgP
pkQKEsz44v9+qChdBsq5PGAk6+YK6Zr+apXTU58oUPd7A7She9RPhycOzxt2kIuS
HRXpyKmXRcw8Sx+5Zj7pr3oauKzB8zvsJdqTdDzLtx3FYetOeSg2HMymocTpSz+g
Z5VbDxX8cPfit18Zy8BBagtQ6kZqTJttRDsKMUeaqbze3r8r8HlTIKeXI/rlCoeL
vJo7KK5bIlGcOCVUgh7mb8jxZ3/UT2BL+1+qXPZEVQuJ6Bvob3KXnytSUASGQaHk
Q6Tvx9DXqKjKdjg0xZQRf1sM9oMUkqDDbnLa4BoaUxeGFFNt/B9XHsrEDlW7BWha
7IdRE1gOE1KuMhlJfZ6dZhOZxXsK478KuYNFlfY/din8NrzOetwy2B28nI7yKszv
Yuo9RdRQ5tTXa/tvLaqHVPbkQAFLDefsol8RLmJUkEzLZ/YWUl5/YV4UpHfx2k4z
ot3KRSLS29pjde4CpGEe8Zu5j4iYQqEcHilmn3rvnfb5K3jrWiU3yhSE2d9mqsGW
pToJl96waaZKndk7g1IVUDwiX4J2jwI+JNDR+uQWHiEY8KYc1Z0r9tlTdC3XxArf
s+pL15EqOb1IJiyE5E9log/L+NJUYZ/5OD1DAsWh3J3dyE/bGn8MTv5ZqHyZEk9m
P5bHTR67h2NmsUgtRHacnaAVgLWOzKHQYxhYBn/KbS/KlmY854VPd+bNxA2xey4A
7s62YGcqZQs6fED0TX9n0J8HA1cXd/p3kqUy+L1fXatgjgPzC14ZsxV/RkKwKEyn
MOo9qMcHNp+3AZUCx5siLHF5rxEoRvoImJPAEfvfo5kXXxGGePgqtjmtnDRlWomP
yv6Hsg9qc1x+JDjJWTiGtuA9qRcfnwGDolmJ7bgNLla21CHAjr3wXHpb+OvKj/ri
63oJipF92Cn+Y1Q7/Vf4fmT6dBGY+LgE0geyzY87sNkNEwtV4x6PKqJVQaALeLIE
JGnYQZZns1QP7ffTtiL4m3LpzyXaTulEI6E3zggCfscRQAnZKn7t0SP2VzOKqd77
p904BVJhXgwgdtykaeUAz3nnO9vGfIlSgy3CLzngCsWM6UkVsQKdETagSNDK5YDN
tX0XSPdIRAHBLOx8L2GVqWT9dbnvONCCD7lctbV3ZYKHbyk+i67nI3XBxTNm1j37
yevzR5SRPl9bpn09oS9N33JELRyZiWX+wmDB2gRoNg2TXYRsilnEqA7UlcWpTc0b
wZAnSYC/862kw+HMsK/nrhergLpeOXCLBC7OhdYETxnL1d0dsEr2Yrqqkv2BaT2z
mWTqa8d1m7md71pCWoMGHz0+gmQIC+a3qilgaSuXDuW2AEGMU+DyfTFKFaJiIhY1
gHnSrXuoBsUhUMWgmXNT4F6WPpxhB9wN0TNogiFTnupe4Lg9tzLSlEVDUgjJCRAn
1f4rgXVTqyGAcXHUaPb9Xw9cYvjq98gmfBpGr0ikIgKrCh3M/b8XrGZFtDcSvSgk
3cTDSTRZ7EepfevVaqDyGxBH0eLICkd0S2Tocsaa3OOK0CjmD/n5bVHVYSM8L8BW
AOeHsUbVtu9Ndd4ERC0nKeTAtpQv7Z6Gh8adprW0EZi5Di52eEw2QC01igG8eL5N
OsfGgo4/ZIknYkJlacfv975ZkclAKQwb+AfFBKoJSUB4uZtztlygYdYGI1aQonAr
Pxy0UZohqEGX2O/TUxWiB7lgftvupYjISWYjMg56K6u+zbB+b8p7Iz/0bbZMeOB+
eAjTYuKe2j2V/PnUG1JU2z+GCahyZrhEolm/W2UdK3oeB7C0jL6yeqU/Q+yq1T+c
Hh7Yd6TEfzik0pO8EntlVTuFICkrTYvQpvcgO9+vTOhJRWycn43kEW373HPkL6oH
76iO59PQckSNVNz1oHFfoy5EMKlnOa0CwvC83GVm3DGMA/v/8ijU3mlkPdKmi/Pz
FIq31cOWRMH8iAhV6mmXSTDclcOjUT7PYxTSZYpnCxcwtHvg36gpbhQEE+G5LqAV
ZBL9KWJ/GsmRJPiH8sQZMOMj/5cTg5B2+ypPDmBYg16eW3RtkvHaVafKNoBP2PLE
hxXzcb1Got5+hinlK2zVe8Q0xMaBABWd9dmmtWG4eFg0sjKvfo45Id2Ar5eMXoZu
k9SUOnYfbpnuWTIhxZ8Wu2EfkR8Ac607q4s2DYNVdTG6Rw2+PpngOKfpAWeIGJDV
gvVqIVv1dtuYQOPop+zhxdMKv7Sg/uQzE5mvVckaYWcNtgfULKj7iIb1qrYNBz0R
BtWc691TsKfo2v73AEti+dsr2iZdPoSwXt+Ab94SVXmpKrhlu8OYW3iuBwXolei1
JwtOlaqOsftjuh2+hI0PLRBb9q3xnEzgc3KwzltA35PCUazdYqVwfVkarGi2NJDY
Tayg64MvlfivcSA0DdsI3oLBMs6mw3brUAZ/JH6G/NtVoz3h+YSFfUSkwx+IijKG
hebW2fHv75rhEKv5w0HhPHBTpPxBN+IhhrjYJjWWTKYYb+sTP4mWHNFrh4P71YAQ
7+47kSOpG0kTIqKcyb3NlCBjSd6GWBalWqf6Em7Hc407L8gS7mdMc8HPfaobdho6
dMADVxqdP7NoiGxfsz62i75OfNcwK7aUjykG0g4mUJwtOxlBerwZFkKkp1+2yzc4
gUAuMWy3U5JMOv3NxkIk7oCyK9XUeeQSAIbdy+3Q9LXK+plPv6jlvH8G359rWnoc
7XH8kxvpa0wXQN6C2ISiaFWSuRwJulO7ddOajkNhztDdhUQhroSwu8JefXj0lI1I
q4IUvMOcK/zwYCn3oy0/J8t1XFwF1WVOM9Mod02EfsCZXYlI4I7BXwK2vKYEWAwN
zdhycz4JToEf1oYZvPUI6JRm0N0LlEkvoGOJmSPdebg6oxJchfy9QrHAAsuBn6MN
e5bSYbZvikPoMrJTTYv3Q4YJn4JXs01y2lLvJNvul2A/UhZf4Y7FxJBQkpXkJpnq
PyMNisaVR2liDG9CELgTrDDrYLFps34ef1vX27ZMaeQ7Vqbt8VabvF59t5Be4jy0
3gIYsHuMZq/gZW/seA+5R6ZmX9LLKIb0CDCfiVhwmt8qWPXju63SDOU0/E40aluH
lTuuX2JCvVGtsylGX+IB3nSbZDYrDUy20CvpkD5cSxEBykqVEfGFsAXerNNrdAPo
uPcfSNREfgV9mOX0uCxYKscVzaXSCSqKin+nw2hlsyErnQrWWtXIPGPGSRsOPTMQ
HDLFU1WA0IZthAHy6IVwRs/aa90ElMYMyue0lJLj3YFJkD2EvMGKT6Okz1inkMhH
3EZU1k4q7MNPAtI6kkpl5r+p34YklQVS/LGXIYmrw744V55GHMgB/IqeaBoKuwz5
7ZLYgSLPgdHV2wlYCjVz64fYi5K6CatHeOCgkEB1Smx1kXKEw7ox+pTUavSOzQv9
dgbN7nt7IZHMLt/udAe5FOcyhKPO6vqWUr5nSMj2ZM9M9UG1NpwjlvEFR0mZYoAM
ihEDfgS/17uBjkD7esZ3pF39xeXhxOiBVX9dVaojPl1qjScztOsEsEd30sf1fdUz
0cmR9P2lBAig7UZtcoYXHaoCWLTU9G/5TwWQgnZwTWvPJu18NgxZbTZoB+qN5NGk
7SbA5rGyoogXxT/OHKKKyrGJo+iWGvYnM7XxotcwXXeY18SDX5XbOOoK1gadwRmS
QdL45sICToq8Mu/0roK7/7Rj3ceQUn9VBDp/fNVsPDvq+DHPT0k4ZYRs9BH8NNln
60/fuC6+Jfxe0pXuMvCxoeiAvdEEzGbSFWRBThO1fPyEGr06Th9u8sLz+/Sn6TXG
X4sYbMZZ0XQyZJ0+kFGWCsnRZ2rDi39Cvl8xpQStyY3rId/wlCVtch6+4uGEqZom
VkqQGn3w6iGshM2P3j9c8iVEwTLjPtiTHOJDdhzLMKCC23OczHX+P/ZGDNBj1XlD
8GmLlO5EA2GNlDFvORDnWN3nyr9+zdSA2JZzQ7Cqs+/q4n0WVhNM+5dGhKlqINg/
7ZSZI8kEjlaMob3ckNREJ0OagQwarxPbJEHFcAQkmj01yG7hZfav/m8Uz2u1SOxM
EWBBun5mGPRFo8PfLsbfaJ2c6NsBC2Q1mTmuk1zgPYn/5RE1z0MS+sj9sg5g/qBY
9SgzzhLrC+EBOOyik2yzGkEJBtw+mIg8QekhmEBtQY82dGJ6kYOuMuFfwcGVlSXM
SjFcE7wpNPgzcxf+4GSeXfip1Kns3rh6EO1sW73hWkWHYG/2aSsQ/0ikkHpzIjzn
HQjoZzy3xNEjiH/GSK1pA+EAje1rhGoswiWi2Jp4k1Qgmi5cdBUtemEgzI9yY7dg
xIW+vfGOwasPX8XD5N45Um1BQvrOahOZvxwKkUyh3U/touPSPTmh0VVcQa9+4BTl
P5W7lz2lHgk2mGNug+fG3jovlCfZvcSvJA4nTRGFPDaqZI4tWNLS7ozt5T73a7lR
BEvbxseDbMtxOuaqNpt8vQz09gRLzW0HlzMMJZ1GeyJ0RKRq9H+v+JZ2UgqnUCiU
lryt8SCbj7K47kHE5Ni5PudruxoB+xrtVyY7w7Z6jF5UELC+y1Bqu4/Df9n4Yp6D
3lvi5c6rhsOpKhWjBfRFWicRqRvYYBBGSSP3GT62oa42gexhCdXZmmdB7XIrVN7h
LR/nklkboGIMRQs0uqgS89nZ6kw3IIPHd3qgwWgva0L9El7f/C8SaqqdN22ubuN1
4b6TbxFzLYh2DisK6eyK+ENZhHrSt8Izwu3FvabVOICSD9FEI/J3KQjH+jzsVoSj
kkBz8gPnZwkYOC4ATCSYCvlvc5gK+3U1SfbR8eIBKoIURkGl2R6yqz/6v8xJJ93P
AuxSNHoMTghRirn6eK+IRqG/ltbd9zr6eqwfBN1BxO+1HiUFQtgGLDSaR4jY+zqD
/N0mKqygp24QHrPcGT8fm+3DhpnpDalm3IhXPtDZ5QjHPWgY2KXzlT031Vwpl+lX
HU3qJY/UONSu3HjFnEthpqCXF4NGMx8AttWo10uRgdzx8+BbFQU4C+ci0GELOIYG
orJau77JhiwPp+RM24ns0iKALDOsal4oMveSuq5ICKoAEunbcMeiCQ2wT6GolL78
jqHmCZDRdMUJ/dd5HpkVapwOnidTAZb6Xqivu1/cwVrfxtHos16fEtUd/1ZQFLwV
LLBuVpoozT4ihujz68wBGk/qavovTGxezr0AMR887PDEhON3LPZHzEg7DQak21a3
pTrszb/e+DEqkFPJ3SpRnLzw6NRCDQEs1K8BBCKhNQ5KlgWahjE94myNqBrqiEcu
64ioSrg1yCyvTujO2T8yGVdH1jaZzeI3y+x0U34jaE52JyZEB9tR4WopjFfFnJ/s
BAgla40Y5UkxXE7EcRFhFAPvN3P/AMDnYqzxpHoMDHNWoXOXW9lhCIYw5hC5jn5d
HHMoM7kUVBr3OgyYR9NyKEsE92XZ0wcda21fN2zBL7J7z7ZLpLprtHUw9jHdP2BZ
JroDxX1CPsDjzS5GE/BENH7RZHw8/UCGQ9atKpniGgC25h6NI6pS15d6ZUtaiDM1
HBOi8M9taZSBQVOhw9IaGFVoAFT8v7zFAXJRMY9skvwX9dUTxoW39To02QisvFld
ZBIVVviW1gVaH5FnyKufAfmSMZut0UrcB0FfL27JxSNoYF9XQhuyNu4l5JQQkTi8
H9HIZymsbvOmF23qs4jtfBcVnyaKjmmjYE+Awr6mUPTaF+etcoKmRNVqI/DLT9UZ
fRBPqUGXBko6OqQ68XzzOxX0qCXFe28pOZuMVPw1ePrvSZK1sBgv145AFTEXz8jz
LBl+LqDp/G2PVi+ObK5Dj2lhZhBVzesu/3NqHRmyLL2FiJ/YTgFj7dgSmHk6buMv
FhhCWoeCOmad3IAx9T5u8nd+SbP/SoM3YOOHGOdXDiS9IG5Koc8V/TFG9HLRdvGU
9jlfnWfawUSTxFi3SMjdskR/f1hLWJlgIe5aMjod0MImMTX0DZ+vEL1hK8N+6PoQ
c4ese71JJdV/SHY7WToei7VcP6atAcldAvtKCvxOpVdhZenFUhdjOJjhgejB1csf
Y3fjdD3t2PILHC0U6uqCofLMgAyNG67YGL+cbLZj8zHlrZqmjAfZwiSDReo20YAi
hBsnAhTLqreDlCKvAz0xIk2JOnuCuQ6StFYB9cegBpEKUujZtZ3pNmRP3tfEFgRp
JTqOcWTU86FIdI1j/9PKnN2mACryp5BNJtSTqqz0uAhSSsyastb+IZE/9YSr8c2h
MJ6+DaWssCJXQD25IzuWV4HXbfMxaUiV0Fz79dEUSw3emW1DxJo+Ud8L3sf7RvSO
he41vjNHyhnm0yg1H6e83pWujnQ1HQ6q/1limZLqpoEHrkHXnPXsVCV0sjGzOljO
eB0IT1zcFXbtjyLvZgt51byojUhCBMc7uW68W3qaGH6FDTQWcTm6F0zqtQWHeoUz
hPjnXXam+wYPXZyu2F+Ttw4mDlWh6GqEMzzNiMBV7ta44lprigUiAHsh9k8xAKs9
h08uG/m73Qf9be2Y7W1OO7XOacV+MUkalhnWUrU9hbvqkuZgCQKoJ9dqNEKeRTga
POMJJtt4RC4B+QzXwLC8XMbPpCp1IEl+Zxr6QPMpctHDkT+K/23RPm53EryNG+Tc
yM6hZ8UmykfshooGqzXRXKeYoQ5Ojtzi9tYuKQ8OOttmL00xvBGzTPm0IXpqGvbI
nH29MljftmqCR/YnE6RRzKe6D6fqvDWz3A+62/QPTh05+kyCx5qo0Ju5AOK7uA07
Iv+wsfnprYIoo5Jm6lr3fhTXd4E4mosC1Lr88UiuEqvg8I7pbMAbca1XeeAK3Ya2
ZJiuQtalXpmYYfgPnRIdvH80ctBLs0+2xbVxBfO7ou4G6cFcqr1JZoyWt8XSfWPB
MbAOZ0WnnZm8LtiuQwIAC475rM/+PiBbTglB6oZIqR0MgTt8DCjXO1fGcs3bRRdu
ShaIANALCTQrLs47rnBYpdGVDyNa0iNK+KlIQM8EAOnkgmJXsCx/oDsJ3XRI8mnj
f17Qp7QLmuPB7kBrj63/uA7BoFSlY0F/lvfCUERQZqVy1jXNz8JGX2KBse4UhEsn
025GPGZ0Vf6RJxxYF6SLbW2P3VYoZvdKdo8RXttbI3K5hIJ3zO8Rj+Nhm/eIr+9T
bf0PnyjxGhQS0iWfq8XBeI8d1rChDWu/ZaI+fVGTMGGtWLWtm1Oy/GoO+JwfTkOf
theQQnx7PRrFYfzdUHWVqrgfsS3DKmSQN9EN9zaqob2XlWC+5Xgyt5rVuvJRmXHT
Z65sNRv0WH+ceQM/DhAzmZbMLjxI0mDye0DEbr3WjH2YKsnXZE+YuGEMHFhlIo+5
I/x0pmWelxFWrmD1rIrtHHW0vcetIgRATVeNRJgeQlADxc3HXMx07FPryCIXg9Jp
fOC5KaVjpT52lqbWEpou6hifFtaO3epaH+8Sfrs5xkdY7GY88HePyzWIrhaAA49S
gUuqlIZzVKt5BlY220Biz8K28prr5y1/u1KjUCS+2MsnJl8t6cRYTM/d3plH4qT2
4V31Yvw5Gwkm0B9cYD+TFr+gK+ASNtawzufS/yMFPsuthANPfTtCW7F0LS9tTfbX
/8DbJIqxxgK0hImbv6/S4jaI5Rg3EmyF4aqY4ErMs8Pz0C8TYjP7ULhdvypV2Lbn
rqqLA55ho5fkpVlPUrZQ4ulRHcYmAjVgg+76kXHuXD00KyZjizuHV+tGYXn9k9nT
up0NNT5wUlCH5/OzqlL94b1NJ53YNgSYk1qpGVNFPzSeC67tY1w2FeNt8Sfzw78j
Y+yTwAURLPvNcFjIKmSlKo93uE9rq8v4o8/6kqHpXyjZmqJXIGcSom9+g68ZeCed
NNR4ouqUbFcV2msH4CgkmNokaNjzPuB4QtQvi5B+vrvO1WiDp4T1wHwdGRbj80KU
xzCCbZegfU2Hn6jBRL3OivyoLqqG5HOyI6CzasUfLnl70eosQ5JLyb2OJ2AqbeXz
gBJ7ZiK2qxtLzQC4xCf3hKNRkif3h8ScfSv5anX60VePTsY6qJe2vNAc47mHcD2g
wM2WbVFZSdmNu48B9L5THKWv6RHteP9CWE3mqXNrxlHdiQh0vDtdsOlvHM+YOqoX
8U9n7uWqPF55wawH/virJgDWOPduux1mb5KbtnnzyZe2sbXwFdvoN5N+JnVXfSb3
SqMvpMpPrzLfuAfoPncOm75gKSE+qsPg7lB32SYpKfQnqPMCD+THdWt7G8R23Tly
bzkJ0GoMQTn+mNiAA1Fu5dLLoFQ7KiYNNOy593mxP10mM9nls5qS5DhDg4ZcHtG5
SV6OwAnETdxKGm2hoefSemE5STP1K/l5zi30tC06hQgDqeobTuknhx2/uz6Q9859
Z4Bn8sxgCvwHne8omqaeMLR4k9DZfqdQeOXwP8Ckw8x7xXpT2fTRdNk1uNoe/0Y9
WOVbehQXBBHHPlzUecrRlRK4tM/v6e1a9zC3vhRMQ7hlRkcbCwioCHiEndjZ3+94
DoVQVco0d/ZunQom+rqkbL3M0Zp5gtHwCYQ6CKw7B539s2A99wxLmIhVoWxcTFsz
cJPvJ6L7FC2xtqmIu3XdLzh0kGomQ+tl/wtdxdSLTsoV9dgSPLFuNo+k38LGm45W
jOTiFdTiAM+LtLNkfXtQa+NZzvWV9ccbMufdz7ACnzam14VzkfL2C5ab9CwrGbdL
NVIgpqtrzU61XqXdF6b539hMZAEqnhKvQtKGiEeEvvEKmFyw+tYwn76zKXziNwxQ
z/6QGHKzCrDZ+7yl5/2n257kRzOK5FE0M4qlA5Lh1mQ0ycPtTrj8TOIwOyatDSMD
zHpKqkpeNj0InpW/Z0FjGpO6suBNcdma5zqhf/ztVWy4iyGNvswPzihXGBAP0k+I
sgO5mWcbfd2+s1c3Y899L/65FPabg6dtjwQh3EPJvXLIip/2QZN9SNHNKRZybi4U
KHZJDG8bsk7U36CWi1OlZubM9Wqt3AU0L3GB+yWlfS3rgjzd4OLUzJHwYl0uBEmt
ojdkFnzxrG3Y9vE7mEpXm452Zz98r2WEZ3ofTZBQ6lLqxZSvH0KXkCMwYc9WKk4I
rWKSoNxDGHkVo33v42zqDNLx75X76WhlLVsRfEDIq1BxxzFHsjvDxsolfsVpqsQg
mk4OU8QFoeVAnXh1qsWgcovfhb95FNxskAo9awJF+p8w6+m9jgoXWGWB2zDZRi9w
K1A9Xfw3X+os7Nj4yjhiKyQVuEBHgGUEtqD1v82P5wx5SX/mcqvFNiZ32QTj58q7
/GYyA88rJBeUZPOkSPRNhX9lWopM76Pjk/mG4xj5H04GUTZzRWoiXOdP6uYH9y89
MxSzWle1443uX07p6WOCihbtmc+OPM/EoKbJhfDMApCalNOFMHuLumtaoLY14sRT
MM1stTMnuDHqhfkcmUBQ1ADrsakMkOhhy/B1ve2mrR5qjsWWHNuQnlqfAOeNjTUD
pWV280yKySkNTy35PAcggXvoUU0FUo+T5aBcYfbO9GfqPFU1WhEQ8/ld8jNk661l
H1mVGftFREPKYIQ2qnCHJzUAPKCuixwo6vUxw8X2XFgwAk/66Hkkc08Ts8BjqlVN
Z/A7cFHbTibvv3jHjZ5AHFANbyH6/nmgDY4OBZXDoVrqwY5GFCn9iQ6eVpUoo7I/
5/1EJuqylN5D9K/h2mcpZWdrt2R0YXGq9obOlY57npL7+x31fpMgVyX8xxNzqJHK
dG5kf8RXynQkD5LlfYnDukVqM9YoiI4PkFjA2FJRURxr3lF68tJjxvhBJ3ksy/H4
YBehGGaslF1F3YHO0gNq2sfTINHZSKDgYrcEY/HsqEh7P/7y5GAfdATK5n9NFDwK
uHBuh2MIB5bxUOS+axKOFOWRKvuz8q3LNz/+TNf1DWTaS4qn0HhfFBKiJBpz/YVH
5VGS2LqL1Wzr8zWlIFlCpzw1e8Nh4xMmoheJ9IklKxoUuddrvrHAs3RfeviLnaIG
S5nz9XOAh9F9taKGOR3SGcShKBQuKE3T+d8b02nCyTF/5anpFX5HXI491Lc1WEg1
xA1lMNO1Im4+HGmZrtSn2hlWEe3zbnQzwvPVDOnFrNCfneYOZWVVo1Rjwb9hkxjz
T9D/OkC7694nMPtEW/Iccvp1M4myBzAZ/c8m545oY71KuLx76jnwq/SbC0succcl
excBB+Uw3ooWyXgvSUL1atNYQ1sdHDrwejCQINWQf3ZH3LQ/8PReLjSayNoNyTIX
yUMaaZ1UEg7XaEB0KbE7jdq1MTJQF32v6vy3ORlJrNKBbO1SyfuwA7oTGtoEMwgP
9IikfAplAA+gjlmWNXtP7ceyjVN6qfwH8/OK+6mZ1GgBLi7zD7Q3SA1tfTHKpEGb
1uw0mqo0vLJOUblQP5UMOYqCDU6nzqyRfL7+3t9SrIWPPHsh+mYeD1vfopbuJTtg
hYQGqEQovpxAnZ9++NgPe4aiBGCy+a9Mf5V/uE7LclEJtYSkLhIExORF+1XHS5ee
2+2JtzqLoyckQJetnVXAThvXl9Tu+UVxGm+MwRz+ZJaNeaiga1+utwXw85B490fm
nc/R3Kn6o6G/a91ExIc9aLLV0peuDmduC6UM5RYyuTIhyi4lRccy5VKA1hvfEkWc
f6aY3jerzJ9VRhCuaU2Kcd0l9U1lcTL2W23+E9395Mkkmlv6b2fhZ73UeEpfDXKM
nbU7vhmfJMWZRhxfPafSsZfR3JBt0lSyMyHWlxG6fZalz+4LoHfWYXdcRhAiNRz3
qUEryAoxl1v4ZtRW4GCFzkInAfbKcprGdIW3LQnBU5x2OQBiZoDqJoJdTZ6v1Um4
5KGnp3Q0x8QekRlJE7F9JQKMOHWEr20+lvA8TJofrV/N0otOEjh7qWRvrMjba4E8
r5hs3lf8wzWL9DmlM9xMUDEpwDGWViZ94GXwQZvvbCWiCVo7X65BexPgQQehiuW/
W8kuOqrWutV39nDxP3ceqltVdNNpb9LdtDFvIZqTDk0lTw4l4uJRttlt556IMthO
IvgP4UeGNWYL6MvEJ32472dpHZles8tLyng70oA+ARgku9EhoFA46xwH3I++UgVs
fUk3e+dhXClnMhperO31OrWTwIPWW+DT6fsB6qhCpmV1NHKxsaR7KnKJaBm8nTcQ
j4NlgaRGHz8yrpkC9i1JC/5O3QCCaP90ldQTptm+qcomtefN6WG4J/2C+mkl5/F2
w+Fp8uxnYEPcku61P2OzRfOsVpG1ij0fn8Xe2rPL2TtiTIOr2a7NBYyvexZ58rPs
do3usnnrRZG/6InGD81/F/fsO4AbdRQA/tXs6tXyFLO82y/GnXm9r9yJ7umG6QKw
6BwrQ0VmDXiGNNJeOhgp/SSytVPmBQ7SRtDjg4qaVW5YPhcesTGOvKesZx0Pm7dR
lunWlenxNoWcZ+fnBpbtqYnouOg2B7Qfb/sq0GYcs3umim6bRbigqZQTMXD7jSI1
5M48ALl1+yeA2aDkCeWKsRECU6Ts8h8BqhaI1RXpHl5OR/SbocSlL0Gnu69EH07X
Yx81IxDBkuBK9m52TtIVnWIdButLLhql/MQGC1b8xnkJZ9SIyfdoyr5bYeG510MZ
G7BE7BqgdnUMqhrEXqsk2EJbHkj+TuAiBuQFUNrzpqeOTEr+40uGbNw3SrPVbhr/
z861Za7GRpblvsbXwJj1v4GQ6SinzODRNjy/nNhzl8ELSwkLRGDgS1yQIZV5di6E
MBbyakACZ4gZcCky2djsPXjiq7/wa4B79+Fgga5JabRNum6pQhK4yX/4GMyWJbqn
dWZ+LEr+QTrc96wAZeDBKfiHTuH6bycM+zWAs2NvjwXpc/GvXQqua5Ha8Pc5MbG0
9ZFGAZ2d+Px4131fm/3mjtNHeDWTjVXu4P0iJN95kgwLjQ5NU7CRF2gpUEeUAtW+
mIX46nQ/YbK1pab7xHmLnUXFB6L6RRG90oixWx4RJ0cNIvnafS01HkhK/bp/ZKWx
EbZR/+flnAC8m5NME3RRGKjaPJupdyEsW08b79leOhP9rdDusFP4SMmIKtAwvULF
T8nO38JK+/HDlEWndL5cz+8D5QrPZ8GSHOAS7FZELZHRicPS+5aw+qXTauGctqCA
C1UFWpNDn3wC7yaUtmFe7I8AYYVeyeBh2KrAG2RKmBXU4+1bUnpRtbKjuWwUFPzi
iHXyswgR0ViPcikKpiZZovYdWeNwDf7wd+BCST+qt7bZ6DBOoiGAPjESQE+3muOg
levSWgsRFUvjs8L32wlwzkwVoXcZBBoFTIF4CMEUpRE34eajWR5p9CUL+AejRf+T
ed6kiz60CqJJ0kOqj9jbrX6DcamQJlTLL+8856H8Wp+H5apVYxnK/Zjv8X0u6ikp
J5gbsD0uE1i6JeYvkhUwbf5+6q6UFFUZNKUTYh94fVrRaPmBY19GhRLipldo8AqJ
T6pQlEajfLE4gGXkftxTUBoC1E1eddTObpbZTla68KEpnWWW0KsYiMwNk/3xqTOh
d6P/eQSN0a9QaAh46sfxZ3sAIutLJSqnFvg97zRfw9k7UNYwmsQYQR9Lsw7AgGJp
wgMkD28d34HCdVXfO1aGGE0ot0XJawyPB55ZUl/uNTP4ORB4TmkM+v4Gjzb1HXge
Gm7heoCwj23+yLOPU3070pmmpS6MD+wrMW561J8PgP6Bm3RRUrji9Hz+mds9//hb
yOBlzys3/xD7qbuq0TehLCc5SQ34LfRNY5P/dSIymF08ypKnHktRPL53VYR5jyvZ
eTzroXDwV3V8uZ2Hb1A9UgYGr8bsIU6lNwGTiebcHykeu/pcU8fqzqD+B4R9XulJ
nhvzxs72plgtfkW3UiDHxIFL0YzlLAZsFdd0CMXDzG/GOtudpkwXJrXy9ngaA8vF
N1uE+bTt+hnkZ3hw3aqx10o2D1B6ro0lDgE0AeTpv9l6t4RTRi48Fjf0B4AUvJ2G
WfqpSdXTOPduY40MArYXfmbPvodM7GvRbkeR+LWVQXfQUpWIuXjsP3QuZquB3HW/
s1aj2xIJ/qJfdIyg1kAQIWLosxOHaBGSyvt68YnKSs0asmcCLE9flil1Ua5g5duZ
OA2sb/WQVRHa3UsBQbTxiZnKm7V4Go0bbHgEtbxWbbyAz6wY0ctz84l2BHgV+euS
GrkEoKr5TD3bd0ZRUbD+NSoFwRJFjYXs0GSOw9PeTKmhjRl1YPZMYkENGNOHfApo
YhQLv5vWeyJ5jDQrdLTA38D98WsKSRVffK7JxM0cMdQ//Bxb2Ml8unIVgv82EFG1
4FMdW/otfGGftQS7Fd04UX47c5huMC6joq0UAf+SUucWvw2rGSI01bO5r9bF/+ZH
+J9qjAm8kYm+zrVCjktMuxCPMjIEYMyYklO94oUnTdu944afnJGMRz/ZDpxO9ISU
IATtVgUTB5EWgyhI8PYFrLFHwG1RtZ9NYqtkSEsnk2tFjMHOQl5lQmoqFQRRXv3O
Jy35Ho7s/lPyrhzFVB0MUGs/U3u4Pyw0gcyCe8K+OJ0saMUT8Gos12ztAwdANMRO
tejFyCgfe9NTyz6axYil2IRfrSpfmZ/iDv2TQmhZZbhShOycRHGCCpeRIk+pOwxT
7PfKyIvdT4wAlH3sObZ2I0tP9uh6wv4p6G46MGchafFFiBfnuPNZFrRpSW2UejYE
+cZw1QZxarBXOxVXtx6XoFJUminSaDaqDL2D66a3yuWBuD4y2olt6CHBFgoVep/5
kIOslIzeP2NvhgdD6osg9kndbu/6XALT9E0juVGoNY1nyTFsAXYAk04K7+KATEK6
daYF2/8d2jPZz2tLy0h311QUDwuQrbtSpWB6x0gouXTTPYkoj9u0cYV6lYalWrv+
wI6OmkSLKwWWIEfR/xblZxkVgq2aFItRr5tfQeUOmTo1hTkspzP1Sue8/QjsRltX
131R28ArdP0dqfhkSQgT4GyX948GFxLtkPuGQ4F6wnCySM5OiMX6/VqsWq+pWUeY
W3QKCNZ9VZoKibza1IfrPyjE+LQWVflczZppp5UThCAUJTbqH/33U4jNgz90Tar6
pi8QTXrnAFIhRu/RcPwY9kQVPecKZHNZ0XTOLnrZzG0gz0Y9OcZH3uoWPzcJqA5D
sBODfLDRnIorYTu4PIXWtrBacPUn1mqsbUGeRKrQuvBI3g9BoF0JKq6R242QZmj/
l7Ompo2qPENPEROEKfay5a1eARnmPFCdZ2rNOWpMeyDbHg9Xfku5qab/dPslwfKX
wBcZiHAcVe8cdJHJw3XSAhHcbnp/GxcrA4WYv+DADTT24dSQQJ/XujMXeRIxD/UN
koIfh/tyx6EF4NGml4WOHT+w2r91QiHzOLE4BiKLyuERCQut9EH/7kBCFP92DAIX
X0vYL0SxosGMF0Bbi9v+tpW6waY0sN9YIUuVOSmTa+FdJwiiVqQz7sZbnRqGfnFh
/PMtF26hHtq53SvdMLnsosAW4nT+nXHlTp66+cDPw/OiK0reb3LyeiL2rQa7M2XK
49rQj5dMN3s/3a5LcsmADZmui3AXZ2qaBHYxx+k+dsSZpGWkOUrne9q4B2jwm3gj
s8NNF6AiBsnUgm5o/0nYMaa68RHkE1vW7BwMDqw6nFjgd+bENux+1GR1T3UthbgF
REmMVJIdV5jOkycKEUk8NaD1NZMBzhY9GOKnjYqenqDQC2c7KJbNKVyHecCK277y
0gViEUTOZNN3mlJWOSM4gKEKPiO0/WCdm2OA1NHf77kI/ztHMI3fdCE0DXAJE+v0
Kk4q9HTP3z7LGQ1aktRVtv3DY2tMfQIwtH+poqmEza8mPStN16Wj4R1uCJvJpWbz
GVOreImpx6Pb6bnbGj6a1kC7pQf5GgUfcu+M1shCd+etUEKujoTNAdJzp16Cz4eS
qv9mrmBA/0yyJdbie6glSd0pM/1JY4aOXx8YA0OJKEHMqxiiRpCyDcOzPNWyoF4F
HA84huKoiuFIP2ILsXRMd4KLxerCOrPaHDUs/wZNVhUHyWk/5GMdxH1o67FgY3Qk
hz2Ht8ypS8Loj65Ag8VgQDBs+OsI++Knb212qV9ZsKqil/GnBUWPcuZ59s0bOQmg
xPDQmn2c5RTWi0lfdba+nkXYv5hsOarrjQOEBFE4xdo62FlDC/0jYiQhf7qtViHq
dwQ0275JUrZAL7T1Iif/Xa61af3mCrU5mnkE5Tgr4UDdJlNnheOoGlsr8LH9evle
uca16KPnC1cpn9I8LBbL8IWNdi3ZgRwTAENe8KJEu6fY3RN8qOCP8yTX8KRL250G
kgR5SEHZkG22/MdVwK8y/GvXRzgosn3iwBV+oRcY0Xjx5GQRtdkNlwyyz2ljpfB7
cSrp8f+t8A7YG30RQVIXrnzeoPaJMiqA4euR5xsjKzNEy2Q0qL+6kwKyFzXRdIQk
ySNYjlAwg1T/QvhwvPglolHq4aMZm0Y7gLuieAD3/yCd5+i0G2/43tJJJ+FPkpC4
ZxzdHZQW1a1znPU8NJGPNN+iM3aLmOBZUP9xJRQGN3dfTO7pqjin/DufcBvcDQ0/
qDSCG+f84Yx/U2ASl6DrrwGp50lUX891zA7VfSvDUOUkdoGS5VcU8rC5WtD9kgO5
7UADtOQseKDXN3h9U2SilgJLdMRYohK20FseHizPs36JuFmMwb6uZSXwE+JFY7Mx
ARUyZJkIKujYRFX0VtdcTfyqFFuGuJk9LGHtGNfamGa3k+/ZOgzPHCnw06E339Bd
8dZ3oA0vu2Jv2k2wW6uMocivOVAH98fky5RQkFUTfuGyhRam+loWJV1K6VAXGYrx
0QM9LRpg7cBBLb6mSmIcZKLG31TWjwELFC606relfy/AShWeowFXWWEm04ic78Jo
zH23TPu6KWhgNXupJdIPZA+7HV0o4+NioD8mxB9VOMA9YuCPcif3NPutaYsJFRuw
M4WUAfjG8ZWuyuIinh+iz6mBjrs4eozQPuC7I01KvnOLQ0LtHf2lmSlIz+8AP44V
RAE9UmBAkrKL971dBC5T04HEmGc1rwBFSczg+DG+jejoqeTRO7M49DBLKivXRl56
wqrRztffQuY+oYYy2EeNL39rIUxobrqmribujyqIbINtNu1HgI0BnlRKWt3Dlqqj
eIgwPjToe1Wnh4bBCcU9db4YGvIAMb+GfycLlDXBu/Zb3JpDleYvn0ZOoxtj4C9J
ycSLuUojQl1ACciHF16PjvalM5J1tXaFqMhgOnPUavDfyjS9wxPtA+mvzCQ7Hrwp
8LBQe8YY0ZALUUyvmJqj44oMgTozS+I2+dFc2hXt5QV9dCyGFCVBOuJEPzDx//84
rh79Ycd0tHBJv3kWrsxKgjGlnr8Q34Ce3JHn11VoEgt3H0CprGNYcB4TIGF1sO5A
gSkXQUp+Bv3eWrcF+on7yAn7SDHrEFwg1kYDYKdUnHj6wnbqK8dh/6bI7xaxw292
Qd0eI/wiqnMCMJM2KopHOyslyN9kx2HTxzG3gRANaZtWfI29FkxYRnEfLVeVRmwC
q8nHZ7TS+LaJbtV4LJTixMR59ijCo/ary3ip84iUGlXcPoeCPTR971TOuxsasVEN
yELUz1muQjXXtZNtK7VTlOcsAwayi+5Cbti6P7k4o1rLQrfQEI94GCSFze83qPoq
yKguS45SZhYDdDAp0Nv2ANlhxT0jLGbsRDHTfXueOw2F0UJpadzPIlb3etiSDJfx
hK5a0adHxOdekHAOaDNrTu7k7i8Mu18scsovDg6SNaU9FcFlF6r5w0gW5nTVj6Zr
UnkPucSHZIO4XnuBbAtJRHUeK2u53YjpTmn3tWwD5GDAGZA5oh7wLgoYG0Y3l3Ur
o9TD7INqoqmuijZDaD0dREakQ8BUwNqN8wyXp/nHW2TGPo4G1DFlsnif+dn3ZJuS
sq/4NuIRCIbeBSBuQ6Sltrtq4jvFh3tfbCevguWwPCylMicCpk9x3ZIcwKCLJJZy
WL3WL2e5DFasF1ivv8K6u9UiyfzmcfBX4vBv9qfHz1+o4YP8nHDIu5kgBSYar5EV
KySTWmPJlCSDp/yMMiQHK1nygbzOGxNvVieGHTgpK+uk0DdLGOo3AtYm6PSS4d7K
A3vf+zv8QZKNVFLD5DuEOuwX55AULey7E2PKEbSZZWpd8ssJblAB40e1Sv7baMJA
2C5Gh3pGXy47L+BD6aNj+Eqnd1dY/x+rA4mMGQOTsIy0j/oZZ964lOXTgscAaAEI
dvXEjX2yvJierAdsuEczEDB4PLDfhtYOW8TZsfb5IUbxvskkfJwoe2vyxbuiJcng
+jMd/cYvkiZ7+n0sH/8M48ZiZ4O21Zn6DOZ0rdyqxpaDT1JIIaRbvdp4vt6uEpdu
ERyX1TJbYnTGAeDXsyiExtqYmMyjAMiIjhnSuCRAMU08XxbwdG5SaouAmVjSTfv4
a0u49eXDl8LXxdOxZSCcrQ6AhTVHt1ShV7nzrAUbkB+VunTVg0H1cdxbPyvd4Pi+
DLg1dMyIHH73q5sbNiMuQne6QzgtMTsQQ/BF87eIw+/sqlljJTy+XlPYpRT8ZWBq
3UPAeASrJwWyl17GPZ9QJPxVosvToPEzYAJD4EM4TlaaF1z1QDoOYrpPRLn8f7CE
HLyCcQjBy9H+F5r46tU21k6RSZovIICgatmCpL3UBRaWGApmkY6ad5FiJB1z0xrJ
GBwrxU+rdNTH+HE0R5iAbontwnkdnuSvTHDziSxC7xQn4G7z+Ge6dWms3EBFl5Yk
fgcVUb9taW9KctVWXsbe+vrxBntYgZVyKeyrDIDNZOaRHUEmuym3oyXcDbDZ4RN0
XieJVKZ/dQjGHKaukRt2GkZF4CcEiUKAlES3rsQ2QZOmdf4Bt3QZTlQpkvOu2YAL
b82zxFJFy/Sd/yQLRKW2i/YkKCTQdiY7lDTgbaf5fNgFGqftOimVE6VbaFOiHoLh
iwQRsw3i1xa5h6bh4uLnGRHTtdlMnHPJ6GW+dvXPW3r+DnG17hGJoBwI2yzBb4kI
4rs0l5EEG8LLjKIxNDxhoLZngah89XlGZRMNX4hnryqPMAtDEf5qgSKpk2sqd3iE
HLjWh6gk87f/0GBoR/iD6U3d60i95Gzu8+iPYfXZaY1AnUvMPexH/JemQj52oHTG
EYpOB9Z1Xu/SqoNDaTTnD1yIdrKMunfg3H38b9EOEhYLM4DdarY6n9DvPA+0c9K+
W08ei52SvDnd07wVTkMD5Kv2Pdx4Y5qa/iDJGUYXw3soDFrPKkuRYRCCKzWkm+12
MbYhU97BDn5mjhKJrlKdgnrBIOdXnsZV+5m3aKYLC6KUci4+i8+E+0JhkXUf/x6d
NtBZ6HvLd/Y9MciAb1XngFwL9UJ+a6qhMaKcuK5urqqGq1qHaJhK3IuhV91eAfYI
pHwMwp+p9cyJmrBfVxjn5vgg8bIlVi9lxCRXJTNWppD7EKkZNAoH3peSGpw1HM+6
f6wkUht/yk1jPUOZ7LiC/D8TMtfPagh/SONfPqW8ksls8bVUKUiY9zJ2e3PXq74u
lD4ARBABx6gcgQU8oIYc/NHsg//9tbprHd7/kR2GRj/qSy8iLyTk9DIydnflKxbJ
eJvzNSKK0OaO8Z/OyXaunTGSULoZsT6eGllNTaF9TYk4IP1Tt4nPKpOLDnBmdXXz
3RuRqJQ/5Pu1OYr0zqYlMLkKU+Ad6UJCY6jsgg1X/Ydvk1ZBI+Y/AvSFDqXu7Wd+
aS8bJeWyXfhmygCHfo4QshhLd3fSgOwcW5pSPLViol8v7nYlNY3ROgD2sDX0AT0t
gf6NI4hYL8qqZUcqm+jo5ucJMU75xvvRe7GLJHJTRioiiomd7Wlg/y+OnITiVAha
sjyNphBXMDTWWIN6UFY2ijM+h7VFITVQ84HKVN2bnpsN3BTbYxVIoRzxMInkrwlx
MUtkh/jzNIVG8QBoyB33Bxt40sbAkan6b9u+rXSneIpS2Ek3wD4bzof20B/8bVPU
Zgif8J4OZ2UJd3G9MKFUCwqSME6Jmn2yVDqs8EZGZ8aoAymR77E0DkbzORkiyjEz
Vny6/SALtjeqvYfWEFdeAHaumCBDl/1dNM0KfBtAU6aPZ1H9aa0o/6X+Eze3RNJ6
zLuXFypGSeWzfFpnrk/4QTIiV66KsqjZiZcAT/QdYLc5Yn+HBajdjrgoKPaYlEMu
mJtYmMG4go/YF5STnxp11+y9ajFzH81ynECB8UazMaHtnVTMcJQFtEU5W3ZPPwzU
06wUMO9sFkrERvU+5P9TYNoXtgORZt4zVWDQyWXBNWyk4rXJJH124EJIcpvx/+9d
EIH0Ub59R3JFvQSJ1h8wpJIjIzsV255VSDMnZ7GLCvbm2mQBjK8z/fidSftD4t67
OFVLJApaCSQHhKAHIYiKh8CmlpuPWIIs61IT83vsxYKDIJ4rhwRA/TKFBZfRW6jl
d6zJf5x4CCvD659/3Ar9VP3Kz2OrLj5Rla8H8wadgr5UQ7pmzdwg25fo2zP69Wj2
fY614icbADRrKfT7gTsw+8/fIBZw5GY4LCpRp/f1+PbEajEpMed8GeJRu1INDc6q
C9Aw7v4LcQArTgBY58uiuBhwFJjhKL1EEqR4VTke/EoLOfNYshndYlqXXDPewrud
mPgXMIK6a6He39029293dvE/cqxWFYGVWajxDfMyvuFXDcx+pc0OEDCGOvl9aDmU
dqFDZMMgWRRPcjUAJc/J/mnRzwOauGcRF5Yp8z1f7954MYJZQ4Zr+Ewz3BZExsnF
ATj9dFG86LFTOeTiWyu6uB7D346th8Gur/C3xgOH7mLIJ/LN4/1YJ3vJmF0vLzBS
52fjgJD02Bk1pEYb/A63rHjuQWVaKYVcryXHFoM+gECbzD2QEKO+vPQTpYYy+fLd
TkLXUKAW6+RMrbMYLqhaZLIovTJcKkrhkSJTpfC261Bon9gawMC0F053QVeb7G6E
Sh+ENtv3OTu12RmebwwMbDF0C4zV+T7YWxxSFc3qXO7F/mlJWghaI9GxiSFsO3DS
lRNbjc0ai5rhpNITsEzqC2UDPQtIGDnwphhtPcWa6juII0h4xOOPoTdL+PnL2Zch
rHonJ5sD6gbtlbvJ4MtnD7gqM27jtaGr84W6AUv+9yAvxpRgUMh0HK80idyw1/zC
ESnCcJ0V2091Vra2uUmzSaG0rAYy0Y+5nIgt5gL5uL7V4OGlxHt7uWz3lLbAwowf
UhR5106O6uJXaorPCssEEblYYgoKaBNrxUXuoe3qaUOkqb/eeFm4zN1Genhf/BnI
mVqd/VzGb2aL0LP5ajulVrlMYldkYLZs8eNDmF82w4Sh8+aRoad1sCEFvLcJiVJK
CZUauwjgju8dJKCiacvXyzfDU3SAFVp23LdyksdktMLpHw0sXhIAvJ4xqpGoHG2W
9YpsdL91CLK8JlC5ipJiEwpZgZxdaarspqk1/emsc6IivSgG+vHv7O/glEKgWXkX
UCqP6VDO7SgRnBDLCTCUQzD0uKcA28CwmN5gyFOJVpLQqMfd3Dlnpd6rccSQEcXr
LOKL6oSgPH9jobfXaksjVou9mQwu0QvllYxcBig02tUa7o63pub+0e5M9SYMyRRI
y+6KsKMEYQ66eqxrVNMXdvamXokUVBuutAP4Gv4Key1B+L57W+2CEAWBY7VeTbAc
svRciwpFmqDiMtE9wfjKqk4It1cfs6jdLAr6yERsjdR7IAGywB4S1QLjhErnlH7G
n4hQPrAQjPJ5ld3ROWrQThQvpt0ovOMxAZXPNXQgRGCWtVnfPWnWWi0pHkVJn0Pm
XtwDfjgD8Q7/Aimv23i/CB6qmdpG1154YjF0l65WPsthSRwUSqY4/JcrQLLyaPsb
zvkGN81djCaMQ/XlVUKhOg6FeXIn4PAedr0JNF2kLrh9vISpuCrqT43DooxV4ZSm
WftAcdedGQBwUz7AKD5Q9iFdyIYdnEewQWKJZ9Gzgh5TLeblNWsU5KgySh+yMmXu
P7ITvDClAB4ol/t9l5gSFspxO4sCLtPOyERd40Y1UhdzmkucWOepjAUg3qvuKN7p
2soiSVSx/lLc1Mnb309ozh34LBoERhn4YSUq1tBKIJM4lsIU8wWC3c1nV88XRutx
7a0EkZ92ftuivNaBP+Rjx+L65Pa6Cp3p3uBOA9KxrvfOrO6dYaCc7x6konBOWN6U
ktxqmjbJGesamaagqdS8rB6eOdd6ereiEWwEhmQBkJSAvZT3AcVXnEPq6OyfH9Rf
TW5H9X91tnUXe+NyUyrYxCsgZBGDO2aGwcUIi2NVfUaDw49w/99DSC1PFkjNhWip
NSGzXMK3IwEmcG9hzw0L2/iFCL41GV+igzMoY9FCTP/pKSSStT7IDR+e9ViM3hvb
KGhmd031k+Rd4e8Cj47SPWHOPqMzQlslpEQCFl8wiCXd20sPJR6FWNkwrXrz3/HU
ywjDp3gmEC9zUbEVPd5z+WaXKCiIRiSUGKOE1+6JV/efhiZNeVSP4dHmu6oviv4y
e4bO/QaP51Fp4s7MRfc5eFEfMvpy/xKTksqVUfLkxLZNPrlPsfMwewlKmLnIeR0d
L7UGgG/atWQJkc5crfZ+QypgzHaehEh4RwQ4jXzHVSJn1bkn8f+UPgAxscoYis+V
CGxB/oBv/CvssxGjie2SiApVp1yxhrQX3bxNUqi2tQDTfwHqrQ9PLqnGERP2Ij+2
9K/CaC+veGuX2LRXzmOJPonxhWfJTy847wO6DrKGXuLw5qD9qQaBcDSDsl8YfOzP
Fpqm/XFtK2qRuS7O3geKuMQ6YAJD5CPpGWWoRv3g95zjnMAvOABrCAh3j5yiXjKv
QjOZ/oNFDz+O2Rdj3ePjlJSF+jUprWT4uHBsocyjB5IjiD1+J891041Z/TgU65kM
jZsHx0ReAeh0azOMsLV7rZ0azfJDmLeVNQNsvXuXlKxNbi6jHYG0bOSOGBIG7xd3
jkWbCQN2cdLSr9pVpIu4gYaibXcDYOMMCXuKN6qoXZkwYvNpgeia+pFUM3ZreoHF
Pb1y6Btyir6sVs2ly9ULuLs8No7HhsfeE9feXoQ3go3tLzy72oc6ixdH61GcSD3N
iSu+atI3cp0KKUBgRW+1DonaFu2Z+kVJzOjwbF4MYONORkvNO2McaGYWK39B618k
JgWY3BACfg+VbYMOZo5MZ7bMuExmX+29yu9F1CtVJWX1Jb9k+smj/7O24KdVRpwD
ho6erG2mWSMR8L/9dPKt2qiTAlBdY8RF+p70OiJMTizA7FGooI+YBUgwiK8cGiCo
T1UWfTICaiyuycwAjl4IZFoOo08hbFH0MDP3SLK+HuRRzULrsSAxulg0kmHkpZSO
/204rmm9qDqwpMjOC7CT5RzPDSGo7+kgv6FCG2N74ol0RoBqXcDl+Bg/wbXtDrIx
W1cmcbHptRLxGlsLXGXRtkCWkBUr9491V9gq+bVAViP3nMES5iI87EQhCbccYsOu
VDecF4U3Zjgz5PwVUO/j/L5578FqoEFhkgj7F7UdozX7Qx+VEdOE8JOhXM+PPSt3
n4azaKa+4P7C168IZKPKWj+mITZ5Ukpg88SM1J9lZDg6e+XT5pRkca3Jryx8MuIX
lVLRYAydyXwd1A8ulb6Uuzm9TFIrG/uD4x2A7Wnm0SWppTk5g8gxPyTY66gS0dfa
hWCQfc/3q87pFA0F8d7DLYLX8CTmcmSrKjD93M38mtgVhE17clJMmgIa7xJiJXT0
8dZxBbf4i72ub+ZP2xVgM5uf5iX/DlJoQkwT3Ky4uVS1ZsL7rKoXOQyW7Q/Nfc/G
4335PkZj0K0vFq7744rhjClY9tDXr3Rl4IPNPtt4KYZOwgz1I51ABmz3XJZcV7Ol
60vYnqY/53ZnvwR0pShxDa9u/PIQGblu5VlF50xAmkoGwkHGaZEqf2vZxLOWkLo6
absMU4zQX33JmHPxs/MtNAf7Kh7q8pqIrugR0z+jcOzOZHaYfOlt0BgFCOwHNvnt
RsfkjJ+iVhgQnr5nUX+LbGXO6IvH2Vz+jQyoMJ3Tex1F11ghPcZ2xSPxTKdGp3HG
XXBqPByzaZ91Lb1SeBG3Fkru4rnKNq700LC24fRlVZcigmYURroCiqak9a12JkV1
5V58J3Zvna8IxkpWWvQMBnPSMeosBePfZ08J/J2ji4T9gnhn6ykCykI7PBeZs7R0
723hd2FIToAAxBviigLt0/0dGf+BR7+mV7cuA1q/ryBN3SjYfDfV6UyiszgoL9EU
UH8mBtJ8bJvxoJsjvNf9lP6zc2+P//VmTsQKkl8tW0bifqOFNggZI6bz77kcYW/A
s7YQcY5qIndjMZMMnHMFhv3dhFpVvhz3MhJZpfDtRnXKCZeE3YHa8s6AF5UYOoE/
s5XeiFmvjkLuWBqRv1ki65ScbpUjcRogEpHC+zfneOXcPxMt5bUavnMHmHelniz+
eJWDbOX6/lSZMzvw6rTybz3GLcH8Q3gqmPpPFJfnsM4rFBXfGzJ2J6PRQ6XrZg06
hN9Y3t7WsLNpGtuvrKdDXQ+bYEzIDJbz+FRkuIWwigHhLk8xQTh1Pqni6KP8eTTJ
cm2w6z1ZlWymJkDjowNjSDdYGQSHV9NyVeJmZRmFAi7x9LKWGAdvWcmoTh4hQ99Q
LXSfYJ/KExBo9jNFnzgVjBermEUCUNYC4Kofbop1RcsIrmU10dFeF599OcctUiT/
OEYhPBWnvzGR+QboO7fSpR2c8bU8DESv8Msp+56vStJnz8TXHyxtBTdGV81vclXU
yeoGVwszxIJkWIIgX2iBWwFsFsxBBOz4Ey0L+HohJnKBXQSDwWjYSTzQi0dDdT81
JBZAo8SoiN6IK4ZhgyhAyzwokcQzkOr4fugd29FJQ0JBa72CUeB7OkaEkQzXmOaQ
P59tYtsjsgeKgKEwy0E0Gw7xfMU5YL6i/2CfBCe8EpuK7aquCzdk1aDCSDVKHt1E
BW/aREFdcCM67LvrGnNPxnHtOYnOpsrvWEP98EkUQKyjA6nCht+14nL+pK8/UHcV
/fJum2AhE3GPRj3vqpiMxcjuS+cw8jHhy3XhdzJnLx2NUmTPkQhu90juAK9zPxrF
+fc+NnscBkuGCZiH55iioWMJ56OBPNGir0SBsGNAyTq6jboa37ygu/T9KewV/or4
Coomo/Qm9DoecP0JFNCF2B8mWJ4agwd+jcodka0Ja+LsnwdcIZ3x4DCKUGzknncY
yRDQETxsrb8O/mhhd28tmP+Sk1QCP7/T3h2998SqnIB7gB1IXnjKJSSp+tRvYgX6
VA8pMUo+2bs+13nRZbvDWXyWsQN92eI5gUJul+lc/VJQSuI8r2zCAqiIMzfhKEGC
DPtUpiRfWh3BQryORyJjYjfAXix7T9HivmM4bPP0vmpwlq4zNCF6czzvGEMp8SI/
PydSXj1a96GkOhHvF4HcuxRy5oW9fRRKJqghA8JfmnqLXWCFA8lVU/a5BBO7T4yc
Rba7FwAHeXAzIn2OZH+A77IHUCwrKw5ZIWci1l7g+snShFkpE47KZ5wjux7eC1B5
E7QazQnyrLpDq+bnZLyNMQBfcaKdzF8kN5EP+mr5l9lHsF3Wat/W+3dkJMJWFslL
puQvc+r+wmjcUOoXQZN/LZnheC5UaBRqUG+D8jSX5dygQx0pU008equCr7u/FdnC
jS97NwNZuzdAbMa4Fq9ZkNlbPpcmoFockL3V05QTNsPEBT1D6RoYtCF8aAOvsVkf
YQxrQHyG7JrxCGIkLMBym/LQs4nT/ZYRRylzrywRVHmkzKb/UPplu2MAzOLeZ9C3
t2XQRCcqy1f/KymYB/BjiVRz1nFeNzS+8eDeksEaN66nmVhT6jQBpXFir7QbP64w
U9zCU08JzRBwedtSrztzr/6OEowQJ2907l31aEqQ1VuYXIdTjcC+svtvbKEg1QzF
3CPXxraH0EeRIVsNZVltZ/R6HH/obczlfkUtiSKZSyqFN3YFvyQDtmlgfC4bh8yD
gkpPKZoxMOZuCc5FtB8y+TLo4bLPi82gI/naidpWS4+cbAV50cEnYUQ0hHquvzth
y/2jIa2ZPy7HAHDUIg6XOTQ/1aqy3V6dBud6RIzmJgrYF4Hj+DYIGLCY5M9AQ9x7
o7dqXuNvoVvpjANlXHJy5cnVdjhK9qR97gxLg+YgpQGLBNsIyQVgahujutELQukv
ZloFe+LqVJ0s9W3/zyGiPeYzx7vrfscDjgi9+wKUbyUlwLegtEeGsf/0xg1xX1Ej
R1hvudltl5agll43NvNXSGE0gCQGnR3pu2XBEWe2Q3NkGSEOArob4GpMGA+sPyQN
Xyp6eR0UayL3dW8JTK+oaDnv1xKN+105DHF8L25yjSzAUp50Dw3tOdY56jDhivm/
MmlvNospgmCAE0z+ORto46PtPgSp6cEZFcoJ/WtS+9ffrqKwc7u6nygx8T14KJ92
YinARFpqC3Q4ZntIY09AqWkNZonOo75Y8LgJzkq3dFBnx9XP7ZeLRzQHRPx1zUYj
sSNFb24dNq3+6TsKVwZx41sdAApSAHxhHvNfAU1ONkC7YVS3D8bss5OFVTB6j+zH
d9tvdzMtOgTy9Hc/OZ2j4IpbNj2l4T6KVfhwzMucuY8VjmkXInKbJ8ac3uJzjwwm
gRNh8FDUtrOAibBowmBJIfE95QXpi+RaNYALFK7BathG/lQ91aD4m5J95MzKzgJ3
XovCH6sSzmUCd6kTRIEjdyr1hpd3FsXNhiis9Bo/54xHUp7FztphVZu1vvtxycGs
5+FayHOHN7KZRBDY8r5X1AB7xjXcS1fiqiKnMDA2T4hvunUts9irn2UPdP4LxfYD
mt5I22zPP6IRcq5i3sgmbdGFJZZsj4IXXzLTSjx8QSfiffGTDcJSg4sRhne/Xn5X
/9aGrrvbsoYcuBugf8uWizY2S2M/PY0rvnYJzdxAifYuBhg9e08DQCYpd92EI8Hf
WqKtkp+MH8qKi4jjK8dlRd21mz08w/sxIDukfpXU9i7F3k3S7ZzQBELjKhx7fhJR
xo96qKjM8Y0rgFRGHlcD0RtDHynVCqmQCQBfFJiNETSXd89BlAvjJplY0ZGbCtqn
ZQ8dvFklXAM2HN/FBfb1LmxE1OAuqrquTPh0kEXek6czvOCG59Dg8GE/nTj2CGRZ
tjP1X3ZJ6TDxvI1A2wUL7v3a4cE41d/4v5b5UM1TxO6v+8DK1TBW+m1MTSc/NlT/
i3dy5fHjg73x//0sR72v+BweEFIRejHvB4XzotGFxsvZm9YI6ZyeAg9Ik4JBjA/U
Hp15wQgWcnKuvFXnO437spW4wNyRsLUQKojt3xF6pjcYjvK4TFpqv+vUrpPfjpRs
59CcAY2XHjVWtSAO8+GOQ7TSmSN71NQQdJnaJKV0bs8H42JHJfjRmEaJxmSWa/Lc
yQubENWK1cVZefFWJ+iJ7EtxEjl2DFHt+hV+y8Juwij6jyAbMeGgRS2giruMkZDu
YVpQMd0Y7O9RJr9KbRQrwYebQ4Pk2TGckacwdGAyChXtBVljfXi0wVzibwWifB5G
asZtXVFj+begztWsTl6U8XRX4s31NpTqSB1VrStoyhw6C5zb48KK0QtPAnPN9d0e
CFC4IzxRLQzkRTXJLex/No/vjdmQNu/+DP1Yt46nx3UfSVed4JBwCkPyjt+YFy+7
PS12+unSEBDgYdwXv6uEPHJkxyD/XRIrfVsrD1FS3qgpP7Jco3GLaL7AgpLPkwjB
+i9uzJ1+YhF7WsaEsW+uYf844+MOAc94AKxoxgcvhJv9/l8fcFAnN3PYBTiVUmCz
ZID1aC7jIzwV7dRQlS+ZJu6XxriJz4opVhb78aBG5O2Du4ANttKc85MPiw5rQUFY
vPlPZH/pw7s8dBveC7n5qmoFTKAzHpCfZE1qvkLS4lVNqgGXLSm5Hji61a2nTpiK
zFKL5osQO7wizAXo9Q07vsbxVnDUm8O/u25+Lc3zQAg3+Jf3wlnwupL87v3bfM8r
Ql3Q+NfUklTsN2SzfvBwm2czIj5mcAVwsj7MANiYEJHUo2avrIOmoS/Ir/+xcQJc
7zBLr5FODctUVNJA8bJHZyi0rQdo4vJFJSpzC+DI2pv0xDp79edR04Wuxi115fjd
hjhuflpIlllbpmLrOBFGBzajtUBIBrohUFRvH4pYv5qsI/PYV8MKhHG4ZsJ/K6x+
hphXFz9QiW4kibp5i/4Q49EcZkZdIlnF47E1C1KtwET83h7eOUJIS6gW0Rtyr3ad
DgTj7AenrZI308iflv+HzNlNqJD3iM+pJpB8wOa0mkLV6Z9SbAc+pHr7xtFkM2sS
/u+rKCjQf926fGYo5Gqiv1NKSzOZIElC5hx0nwK6TAa+2Zc5EW6AZuChP51yVPi1
UYXDhRXfl6720t2uIABWf6+CiR7r5FaasEbqheLSz3/4PvJPCLyvhjiVIuHTAj/B
j53BjizQPQQXz5VpCgZ7tT5BAqhsVZIfHX6O/xUmxFqhK5H5S6J19DZRjQBQF8s+
E6D7eI9nFpOqPYkCwKvkzHU4CkQjWYd5URvBg9VfL6q0tHef0o2G8SMoeRSvZmld
2mMB0XdOCPTXtkSxNGSUCkXDOpAU1HCPoZsqqmQ9QujEsQy2xmA6JyPwkKwrdx2J
bsy4fHnCszcbwbFzlGWx2J98dDQ4PImAX2Nga9lt+yhAAAxw40WvpzsbNSVnVWMJ
tIu51EtcIJxoXl3+4oZ8jwYYaCiIydHBhg04YzaS4DY5cKQNfO/Mj4ZgA+0yENTI
ufHNi/pUfZVvp3lsdWApKVq2UKJyIKOgVha4OvGUQXUquQFRwuPftDLnqqiYFJzY
Um6T0v3y9ZUkOup510gPPK5Su5EQud3Rr9NVkdyF8ve9ZUWXJRwwG6txvCvgpr8s
0VCqLRrgfBEgAFNoeE5MhunW2bJWxoY1brFNQwSpPtPmlYqjNE4yS8bbHX0wg+X7
oTGS5IhwLXq7N27gWSMKM5VSQLpdHZFZ5OcyZFCxixHUTp0i0Il+c4ZGTJK2rJLZ
AHcfFezY4mLZYB9O+TGovbupapBZvWRkTCLH4fG+o0IEzN4Y34LkIRaTQ+JPV1Au
MMAubbd0v7vluZiewotrSJ1h1GvuOFwXfamn8liALFprXw83GOm1mRciig7cDH1k
8U2hdqnYAWQ/Yp80xb4YRV1jQy8VXMMcheoxwjI7nhTEMi6knwRzG38c81xf9sqt
VIHxyVOtLm1maU0UnzszRHKu+TZpOj8P5CTZ1EYADLGRRvkFjjdaeKsRBtAN1RW/
ElqXmiHMDczfPW3+5q2zKIAyKI6QAMtashKMdbia3cFLDICjZH03/gjZ516yF3D7
sAlBdzZsoVAMeBi1mJQwNV25k7hF6gxifIMzACek2DYTRlNk+QqvjYO5G19pbGth
rqGRUM/1pcUM12RiDol+ToJ2U63hiKVSQAJOYG9C2XkvU7KrkdgYTSjqYRs7sQAV
YdW2rZUYdPazSavrBFHRrhyePh/ez7EWFO0v+EeT3Mk8uiuoY6UsaVtiZftPCuKO
bwRwkbEtFMoHqbgCoEAierJCS1Ba/3EEEqruIA8PoBGHCjNtcCRDG8Xd1SCOmgFp
rUgFvRlTdmoIEWN7kAh4e/7HPAjrfGGsF1OM1Oj//RLODyeQOUmZkWLHYpcjDBXa
/nGT7BGqfBFhKryDcGo+jaUUPZCkT2ZgNZp527YCV+OAn4XCUhL2qXat4WJEv/hw
XbY8L8APRERUvSPGUnCKYroSdOtk2XT1nl+or7KFnZLDjovL7A5h7170oOUrSQQd
YTZsyaATjI8jYH4TuOJ5WyhzymXrtf9pe32EaKVRuLzEQm1exHwhB6uACBNHQPN/
ZzHfiMhCNClkh6A36Fpm1AdSy8qkoTGT4IM9Vf+UDwWLgSgG/kR7YejDGSAWth/9
8Vg4Bi2w7zEeuUg0gRi89kJqtrrF1iAvuNZnuhOLt0A75VwxCVI84PruLBLeCxyt
XRaUBP2RnQ0UwNWoWcdgkpe4rRIyNVnLRbIIaGEqTJl+GiBbYjtyEi9aPMM/B6l1
HjGWl8fDO5aCeiLf382x54ONtUJF/qTHcQDHdDKuv/kf09k7BRUU2QGiQ9TWOIYh
UnKTlZI/v474XaI3ugWwVofabw49N7tHPsPXwWE4LrK7qicBOFCdpYeAEHRdOSwC
DLLFyTDPC7yJxcU2204bdTJUHiHDl1ZzfQQDFWrlibYEm920BRI/hF7L675Fb7m2
CAq3uDIbMGPvoRBY34x1frIyywU/Z7maTkwjxiVd9ew8d7fVzC7MUCZUEyuwDVH9
FSsfUGvhhMbCaTw4gD6vVz/+gX4OlaB7uryBgS6XRVjfnqMge0j/zyJJS2mP0xVL
rgq7UlMcNPbVQo6TMBRNToviW+t2NYGUjFFmGxvVc20lj5OacO+XFNEXneD/UGE0
dTpZRYzMNaydJ0sQgcGwlZQxM5uDQ521Ik2U6Y9rvg7hd6ZffEjG1PBRDqdFIbl7
GA7ovIq25xEaIK4Vil0GuMG6LBLT/xMDQlm2npL33OdYPj/q5sya2TvPhYb47Z5E
pmR8xZby3O2T28xH+3d+oWg9V91+KLAqaE7MwyGnGloye+Ajfr/aMsJaU2gWAeVn
8+m9bVAFilKORnj+AfxvL7vdPsPTt9cMl7IUjkyEPZQxyJ1jV+UV7tlqDXNcdgX+
9htPjr6MReHdeP3Agy3ECR+GPPpptAmT3HudZREm8N0g/4GHJE7SQuXiNZ+VCjt3
rL5x/yrHr+8sdSl7OqGj4tevJf8MhW8hgqoNaJXHLM90sUk6/CjXGJkEiwp+RcTr
nDLIL6KDplhHj8MyKkC/znYYRwB6FkdN/4Uj1yr96lOilLVeEb7PjWopB7nchf7e
Atxc8u3zSKzhd0ceEsx/hxynbsJBGO7d0+O8dyyTwm0ZLtHCZ/aPlkHr0KYoV54i
Sj4aaDToOxcjmoaqd2UIWwiyF1ZZF64UEMvk3DdlATlkN9OtpsJ0Xm+F1nuHzCBJ
9ELOKl0x4JlEi0THfsRyQwYCtS2K3ktifh/PRxa+RGIxdv8zpwSTN2y5lXt20Mhg
14JFSqYZQGhlBb8Hf4Bng2pdgZXmnM5AAE6LfiSPEky3DNBffRMtg3ojt3MoZfR5
oldS8UjLD4g4d3PNW2hLRhyfrG+VtFV2s3e6Ay0mBNWWrKoZtqDnn4J7WPFbQqcW
JV3Zi9E9GIVfQ6TgLbyoHzmKAyPbUPrLnXKtNNQw1ulYisUiBHqvuhu7xcWEE/yr
W1OZwKHpVqE3Mkt8R9eHqqPtf8N83SXCo6MBVZerOx7j4RFL3DTfK5CuJMFNAEzZ
i+z0E7waoRR9DIIXSnS8QUEIzHvDUB87Zv3pGUSCbQkN/f4NaT17jf4xwZRyGZDW
5H25JJIY/WUDgaHqih2Uyiat/Yb5XMMKhvQLbLBnerG10jfJqaO623Xsknw7ZCRT
bmgxAnsM4yxen7mKGmrNxj7ZEEzgURgE9JdJOUFxCncwni7nlhCsVvQnNKml4bxZ
0tiamyW137Qy3zm+0B+RRDpY8dRIZqBePb5WRi4cteqDiG7C6sAw2w0X/NdGV74x
YtSpmi5B/X5QaGlIOhDKeAkytO0GN/Cs6Cwbp5lFB4j8oxqaYCyzKPS7/tRIqfDi
W5UNXi3u/3JrfWNVxxsA6s8PFux/VHsyD6qLbrwWrBN3JkqaBGnbMZWbYhatSmRN
T2a2G/G/UqMyIm6/uERii7niWV5Weg1RtzpQUMZRKnL3wSZn+saFDLUH1SOSD2Sm
DbIjSKxvi3UW9YqS08ftr8QehySUbEEyNf+KLAboaaFo2vS4aXddZOEy312rcPWM
rOCGCdNgk26yHPb5KMibR6p7eVGqKBf1wr1bebxERn6WNbXov9lCHp9X8UeW9Tme
1+w1aOLuEnkt5fDelxi/4MwZ4rKUSUX9dxj+yh8qsrFDBwlUVi60fkOLVt2ACBnD
fzUqrPOlTjpnKeYk9A7j4NCZ19EYUxKNS1OzVByomfvmB/vdfV9sZRpKsTL5Fxa7
v3RyTHJUsv+bWUkuvYhy8duGOVV3DHigOBEfExSzP4bb2ENxmeFqmA1l6lQmU3YK
3OAMaa0IAGpT8wRjiDTMT/g7AGDuPC4bdROpoUKdWOg+yJERAnIhoTFWhe6mzcQ/
eR0379yq9tOo1uu1YbW8t3BUnNZLknk8ziQ+0u/V2LhhcbUtoyvrFxlgmpW6OuZP
vVNTxyfppNvuzcNg0/uF9i2B0EdhizKzlfshqnM0M/GPI/EQmokOGOZ6woJZzLQL
WxO91Yeu0HesfdpW4Spms/fAh0fq5DHmT+RZLOmgSZWJHURtdY7e5uohJeFN+Rbr
hVOGh085vMu6odQ8dWppk50xQ4yQ+ZdJfdvGr9Px65u2uhD+lc5DG32ijwm5I17U
Jb9oi/3FzFzkOuYkdZ+FSv9TRdYrximwvv4YXp2lcVDAZJZ4yMxuZwSrHUWb5F+e
Is3XmYq7iP5sTdBOOehidWvP9vC4Yd5LmnhT35TfdFEdFq/GvbcwZW53NbS75dnF
TPHMurOtXbrc1u05YmstRYG+xB+wLOhwdfDGvZogYO0E/mVJiAf7f+DpUzI33KMV
covcaJzwRqz2IIep0QZWd93I/l5XXU7iIJlzWI7rIqhKfBVVEdq9gRNm4c2SCN4+
eZ7bpbYs1OZAcVqmMjfmTvXY4Y77yOHMqSFy303Mp4x3Ywcp6FK/ukPI6OJm8oAZ
QNoKzjqnSC9zzzDQOh2j/7O30k6wCfp51PFXaS003V1NOizoPyzcAbkTr6QHNMRX
6J5VOHbUGZUvDUxtUHs5/WS34txEnsRwy44LzYdYneMaCpsKNoy95FtXB99pm+/+
nL+J3sMnq266rs4X5GPmb0tIePaMQCGvyYIXoXollfoUDkXr+9X4YoI9fnvPwutE
v/E1V6X6hK4TYcEFLfFickWyq8P3WKTLwirxzahoa3U3kehtpXkdEVmcDy6yNM4O
yvaYoGQ46FGcLM7pucXpHJY/q57A2bHrLVBgbKsBqpw3m54x8t1yZ11UxiXokih8
P8XwntMFEiB7w08mZ6/uF3bjBc5lOoeXSmKwZIRsz2f5YQHjc1V5lGQcukeI1OUC
XcUAg4DzOZrxNdO5vUjOTyG08LM4hgTOElOerQ4zTR4rizMi3MxfCcy6vQPuUj08
La7rptmeJmwVc61BVSI4C85U1qp7PIvVV5MuY7Yify8j2yXE/bFxJcg5KCZoyz3F
Ocy4cwUC7JeN30sN4kAHRJxqMK240D/6QLoz6FIAoJXoUMlSphXPGSBqdfN0Z8lE
Be1eCmj5amgD1n7XkLUt54d1KmZLwvAp9fh0KJr1Py9N1G8/hSSIPTYaNXPqz43P
b93/C2IMGM9M72Ki74VKTzAu9fcTSCEhyK5hG3XGCfj9B5dA+ELJCGzo6ekREpIc
oOmWp4faIQLrXsc1gwFio9REZgtcnK69vGyLRUZf660c2OtT5UZyUbocSGeEPzxc
829gsQUwWf6gFGfRujI1CPgIgztutDG/actQYLe0g3Sh/6dqe20eftgYDAFT/hid
40pHnaIDfV0XCuIsLOkkAcXfREq34tidUVmE9mLfFI5BbmvOJIcgfq74t15DB5gN
ipd9xIwOWUIpnp1969q9pi16Mg7/iQkwJ8K6Ym6qQ6u87yFDi/Gj0fevy8A/z/PP
pg5SBZZrIkfR3al4XGwP2G50AnhUubxDx22wYrEsNo256jXoj04YrtLIcFPynbZv
GTgaaHO2Xhnr+DXWnNvIODOlBwxaKYXggx1Z/mNVrYWWS1fON1WBYJtwxRSPd53O
ZnLnVVUKzU0KEee1II+mAznGf11VgabI4F/hIxZUp10HtCtsxkksYVLn25cLsQ/W
S/bI3wSeRWDvHS3UGY1ix3R6UsdF5WyKyVBLmUK1FPjxiwAtycVMVQC0d9y8v+cP
ycSDuXBQETts8AmUuJrcrRYAsbtyF6Z80omXDmPHqNZSQgR1Jhg4k6x0dwqLb2jo
Qlc/K/iFi9nLpEKIbWJAH2gvKAnsN8YHXiBjW42fH0xPhQGXOcRXsNFmqfgb+Ng+
2Aruc67eS3WjmhbuBYMjOeoKx9d4XuYArEQEl2rW8KF3eTPOsY39xmFvEAHRPUmw
gRRy+sJ4LNr6XxQ7tWRbDdlQNon1jieiqJgVVnxyVFoWEq36+c2oR+0obXC3cl9a
m2ui+fgXGPRunbo6lQr+sJR5FENT9MGHfNmfpnwWLldqzdQdesyGPOwtLm/8dF1v
CYujE3meKyjxndrfHpKHZspTveS0uCIKOXdknhkVksMNCqy5wv4NzAAYGk1b+Ozz
JiO1p5jMEcq/qc0ulP4iaCwgJYqYUgk7XyqpxmKIe2LEDFbcePNKIf5dA8C6gCAe
Mofj9ONq1YV7+Z3HrAvtB8iYgHZcAGCy8OoMLyJDi860pIv44MHz/DEmkan+qK9t
bVApsxH4o29Y222z2GbHLxTTOoC5N0XeHeypc8dsvPiPwN1AukGsL7uBIIpi9Iu3
tipwrc+bqS0ZCAQSMX+ydZ9dfdKvL9wQmU32siaI9G7fNc5uQ+IF0LgbzlwOSR2q
K+V2zDdDgCA9UIsvnwpUSO73aOtJUC1ofJr6t4JzqodJbAQG94aiX19SU5CBSb+p
bqr9Jfglzi7d7uOROVlV08hK+jg1u4c5pce+BmYGP439jis5RNq8OrKxD6t6gK7L
01E1ecubGjQ9fQt0BU+r4jEX6U1vTLwu0MggnJXqd6XvplCVp7PMKMpw46On49FQ
XzRoKbeX63wIbyS231nfjz+XDFl2/GOD0BbvP0q5a83T3OSWYX2kiU3JfLP4GCHt
SqOgj5EoPvRBnR7TVZb0Pp45abyjfUI3HFT91G9O8MXUxjOi0Igc+05+Q97YWLx6
n3RMA7sJMZYRwqa5MvlDqTDL+xc3gVNvZ6FkGSYzbI5wocI4O0rW6OSzC9NyrJwu
9LYaTx7kYvh/CbjbZYyAgredBd9i2JVTjezEBpYsegHwQzXuLpJDVRG/+FZ5vTp+
GdxwLX4alGPDkZQMASrvKINYZIwJ5q2Fnc4r/ZQUE4B+KXHVj57j4IhXEI/feEWT
57ffPURVh67Z1NVfyVeDn5giozsvMgBiLGhn3fTmzmt7gcIetwDM/LKLsTw4vrIJ
F2Nl9gJamOhI1/grmKaepSnz77adrdl99hZJFs212yniG6jeuxqEWlaS0sexCIFp
rPPD5tmZiVj0z+PQo4lxvht8rJXLGLh6N0OZj4nEtk2y9nSZMnKFSE8oXFFB66Ho
7S3Xextj4KBlO15GSYVhyGuBXAYC7aFvygjWXSGyJ4wbTvsHD6qhimqDH5dDGt+1
0qsiFPhDvFWBRBv/IHppffVpS2pt3PRLfiNA98iK09ye3YA+2RwXrzZ42HLR+LbE
0VOiylrLI+iREJoWZC/ErCt2FuGOOLg2Bzwr62rDl5efQTBIRWB0rUJNosX12/6Y
dJNzS1Ktwe/TtSvR8fd8xsTDzNdT4cq8pGDWZPRqEwuZzaPGlU8+2+dzqMqQ8aGe
a+ORH6eNGcskZ66QUR+9/uwvzMv6wzWLjhkS2PM0lBYRrliE3vwY50aVzYG1TlM2
IzDwEw+7pKf8AKCHiuOUiBXOpp3hAcUeNmv9HEyU/LFA6FYzRf6nKOaEvrkQKgcm
+v0bSPp/n1ph7Fw5r94qZ4cSiRNgezU6vQ0ksl5cYx9pJtEanzX5XkYTLj57hcuX
wFWIUqL0pQWnUr1wVMGjsQaiJTrGmyMLyUG7NpdYMOmZDiF4/sIWcdG1UaY9J6ze
RQYEIqTjd4x07ogt4phYAjpFPe5ndHYZwFHgq8DM1qEDgMZ5w6Hv7xGjdkZQkqW+
wfjfznDHXQnXk+pSaY7TxMB623I06buphDWzRGrYKuDJTzzAesGtWgKwGuxrBXr6
YIKhM4aOKI5Frv0J9OfiTAc7BR+h7ny+yfTBtV4Lskue0hj/Cvhdt8IHDqygwwLq
rBezmnA7D5L601sQV+J0NfI0RVAlP3/QrnmoMoPJC0dLBBxVQu3GwhkiEm8t+46n
xBi41Y0et9eo4IRmVEZrYjBqWn2bBxkVFU682tueoUIaC22cmxjhM5eOdtumtvL+
o1pYu0Xv8k36cL6GiiD5MEif8jmw3XNm08ivRRJ93XDRaCl6e9inBhimqLLG6WVg
+WEINRCzxakT4Ck0melANM4WhbDKbDPZUav07ZSU0CJUvbN2wYjD+Sv9QyzRWQqr
fnkmS+lVlhfsEr5djoQaJD//QmmEEcD8qnPrw/R8C1EmU0B5YSOSyUFKDKFWLIIj
AngGLmbRnF0dL8hspIk5qXG8RTcWExtxhOsHMV7cDr+H9wY/7rEsyiDQFfHTaEY5
Ys8v5lMt8bPsXpXqGhChSJgtNFna/6XzqwKToihdhqMgkAM4d4dw3TWHed2PHH0w
KkzC76IFhU0hrGieoID0W5lACjhrW4tLFAlzIDUQ8yRNlboAM22Co5sQ98yH04G2
Qq63fkFsvW6K2Pua2mfygWyPILcOkMfV5N3cQ7rH7eW7ikNUHWYjtuDxbUVIsCI0
pQtb+0Rmc21VRjAobw9f7FQWuBfhwMY815hum20EVUY2JqDftkQmHh/R0c/Xbz5K
Bq8MAVUOojEutH3fcBoR/aR2/EIkOBAIzsgH6V7lQrnVpIxFZfVbG0a4xSyB2yhf
eU/3E/hG19xKVVbN6T+RcOXoIEFrl7BdNtD+BxSpSf3RmCP+87LzHBUP9HsUi0Xa
puZF21Bb5kZvgatrhOEgmkTGypfApQLQ4KXVWSlWg8583Cs6Om/oSu1W4JBEyg2g
qk5V2rlyzgoieCUMviQwRhI0IxlVfgQEBMC66wdfglOmzQhjc8b8rzjrVzctfMqF
zwNDQ9+G6zwThlg+5XpA2MwXb3orzUvNoTK9SwxFssaxOQ1m1qKP+GbrMcWUbwH8
M0ay/5lfG117IWa1UqUzCxLS06Ytl1EpHL+5IwYWKTvokoXQn1+zEgalLo1HZzbP
x+L2o2Ndu+ZPQBRvYfoDqaHE+e1CoyTXPnFjo2kA6mlrFiEYNLwjdvnMF38rV9+A
ONKfW4vQJhoEGVc6Dpid3S40pti+2MNbcrsKgJWZvzwcGFb/19bsV9IvcjdkIuKM
iyPWeSsqAqLdrgKxdb3S/TJARdbAfuxIkiS8hvKiVWR1QFQp+Rpmr5KESgu1GQcY
6c1ApkNtjebUQ8R0cCOsKAjw8FotZuCP2Ta5ZXe07EfZCEn4ZpG32bEM3tXue/9E
1d4OPJARsYN+ln1OGLK9TKchtC3mU8ziRUkn5ns361n8fnFVspWOeBDKkLut9kZT
UBFC/g8NfNak3Fb5PzVTYO65H1q1m/KKCMWw/LwX7FKOcs8b08ybmxm1A90ri4z/
IsevgZJhGmSvg/PXj6ZDFJzh4vf3v1bTXnZrSFu3JIVZW8sFSCbQ9Nd7qP9sbnB1
RoULnX5GOiACXqyX3MZgIzpjncFYUbiPf4MHcK9SqWrxK4ogk4Z1k+iX94CK26na
+K7Xhp9ZKsfjFy1EZWDk+taQgSEUEOSBPgyZQOEXkBaJpDYzmS0opihwSoEO6Ml9
UDoju2i+sluWi0J3X4nk6gXbgEEaIjmUNTGYhAb7C1iThnoSyjknzL1MM40N69YZ
lQKTgVOy7Cvdfxd2Nuusk0BV6l3It2imyymC9h1P5jdSBlTHlAZBYeg9ygSe9WIb
5Lvf+7sSZU7UAAD3V9yneXxSiEw4W2GL9PzpUFTECuvYkDwNzyHjNXoCuuEekPGg
tIvbgPNkL9V3vRPNVZ50i/KbWeKHe6RVhOeeDv4fNHc2UPsgj3MvGtNaqq4czTq5
dYkIfPNZl80+I1TQuW1r8Z3Ca78EberiFWgHGBBiF1bTRvMV4hbs7UChxs3TW/Uk
oOAAVaYnLyum8NCfXWGSvywQmmKlOeUv6XcgKsIzYS89P+DBXMIlJAmx1lNk73V/
KzpEMDpUeM5W0SAVPF4xEO+6D9l1dh/0K4p4TAsa1yuvwipTHY/GdcP+tMkSp/mg
Xf8/OKpbq9WVpBFBy2nBTU07+Lyje1PqFIZX/B0QT+kiJe/o631/0vUkussg45IF
RjFnldcE4+XnHzX60ByRFxCQLrxJNGlwOt06GlouCAO+cYF3Fkbk7sKj18SZA/Rm
xS8y1jAlPaSh0/oBlW+VLFw2rv2F764qT1doXYeXTdIDEe7GxbLkgRreNQm82sqU
7hffWzIjKIfuP4jgz5XtAayhBMqPay8/5W1o6YZAlEEJoy5DnDTkqHao0P0zof5I
c8JMwSbnpVICrHLzKxsSNBaxERgwW6a/e8pG9GNQRgDcd4akzGjHijdEUSVHz71k
YHFvJlz13rtvsCWYX6iB390UGw3/pHUIQqGzgelaP4cr8iQs3eRj8SgQGaw1l0jz
Ftvgw026yAVCBN+u0de9MEeYh4TqthlZoCh+uk2uznzc6vgr1nhO2KVqQc79/+rE
mjHCzP/HJ7D7HQ0Dgp0KraxpcJwdEVtqhQ85YD0J2PFbGKFoGaAo+eUsm7cYqtQA
A7ZgVrconHpAeB44bYKijGWlIqVCUsQle/bXoyYYMdCuDcuta0Hf3l+8aPFWY5Pe
pTvAdi3UPo2Qbmr1mbQmhqO7VZVwbP2FvzYIfreryngAhG1kZNSD0ZvUi5UrUexb
KlzVdjAYpvX8Y10pxhRYX1boGmhe+hldKq8TF2Uk8FxBqrQEUcyseXHuwmUu/ye6
Bqbq6LcKKjVC0ujrtnh/AoWjk5jBE5/Bl7METUcPQLcgsZV5IviOKYM7u/1Bachz
bku6hvE4i/7bN7R7ebURoNYWtyAcAhBCiuiQrimqgmPFhudEW8LICF5ER7CMo8Vh
nu0UE0IEWbqTDKrxywX8jtX2tjh7q2DeR+/8wog8Lc0Rr6kQgP8DKb2MQcKLWb3j
MftXxyNkS1/op0C36glRA5B9GkE52+suSIgGNqc8ASk8z0xOe3N6lVllDZkFftan
QQvxFmXZNNb2dsr+4JAXL8Ep4W+U6UecOWISM5qwxXI+5ysptpnlVaWR4mfhJ24O
urhGEqD93UiFOcFtPz/lYmY/IkQFtKheYxIyYEkVShz7nNx1GQgwtoi8h8x8rqy6
TbG4fThiJQkNcD1JbByqJTuSzHbIHnGsgTET5qZe/IOcRccYWwSdn0fOGfKyOlYo
4eqn3SegEibIRHeE11HE+UItlgxxSliRL0VC8lYX0FBbUsOs42Xkl88SJqMljyLs
iSdOINxSKc6FYyPt4I2JhP0n7wir8L1jQOq03gCoLVPtAMUo44z1r88YmkCvtBtM
itj5igxcX5bxv6iTY1KRKOjZlMzBYrrG8gY5WwtOmsfTlKt0bk8cXorKIv3XANS3
BlBmB+rOmMR8oFllFbb1utX6WdJKuGkWHXTtFN8jSunddzX25OpCtfFNhDiZoqTS
DiSRQqgs3jhGm3KB2GyKSTJPCOLvsqrN/S1oTyFmGiQMWr088zEedKMgIYeQMDAs
RcjV7wz4HdsoC1o5qlMlJK+B4hO8xwLJXTihmbBGUuqqy+XxY6I9MOX4UPEl3r/I
A/5KtU5gGrhdxl4gBFX7yDZkGhfTHD3FfV8ThWHT0Un8YEYUGaVdyloZliYtF1lV
CKKksOq/dVACFcfgzItBI9NWdUkqiuwkwUHw9Vu7Em8w35RKvW1+4PpfZG9s1GAr
5M7e0d/TCCgYcYxDo2minW5Co+o1qNue3NC5saqtVnmQi/y0m89kcnTVonkotqVp
sSQZaULeAKL28Mo5B3CiMiKhhv5x0LIqdNF2+mtGfVvkFJXwkbpgnUwCyuMF0rcn
4ckjkPN4gIv0HAO0Z5xGOxHLV3T1t6e0rblKQZ8H/KB5c+0G1ZHS/uJbi76UTjrI
15XZ3y6r08qYsBhpgN4q+UwemIwlPx565z3hRH3C3egkRf9qRdnnU14Pu78Syuzn
VES4HtgDgFcybTx0D/HpJ3M6alkCiWiTSaz59RR14n4YGAZ8xcyKSYLKL4WOLm5j
qb5X0WDcbhUOIEwYZAy79RpaX31+cfQGS1Hrc5FcGaZAepIRx6CN5YNIDRjwsbNf
ZMRYLgt8kCOBcuV8my5u6P5Pql+EaHE5Bzx1URpM2mfsZUV7G6glubU3XX5QvqEZ
aJiqRgK6Il0lPMut4OK9p0sMiocI3ACY2AlVN8pN/9wr9y5p0ezlNzCUGAKtw6TE
/Fl83KhRVsMIqkNLmv3ZITwSmjR9hfRZvOQf8JHtFBn1VMPrCNgybOGhx1xF0I/a
VB8h35QAPxqot7+KdAGIqmD9+kCM9CSKwjOPwFRAkR4X9lwb8VOH+1z2wAbADWGQ
auKJXHtMZdmdVeKeTG7cZVisy8yk4SQq6wW8rlSKYgeGgI1UHhDJmpYTAuqXw0Bv
i7k9kQWSlF9fhaMC1iQ86nRotKl4WiKFfQJsdqw3L32Oi2JvqoZAdi2h1uO2uqGc
TS8WbzPCT/chDS6ryHO/ZosrOlFGtN0zhMWPcQuZGEb7aaS8/zioggmOzoTrriTP
qmbf4z4NiIb/v5OS/xOupFi+MrcyyHr7r9cwyR8B3O3qSbzbR5hO8/Vl397pY14D
dhr7uALlQNwFCfeU+So/QkaFj/Zp4bqcmw8YbplLOtbQWRZs6++enGkNaTQWPgnE
/mxwrw2JfIN2SAzSxDHkrJkrddTJHbl2MB+JIPX8dLOpJwazw3jkpJkGlO2+g9zE
XoGbMnQrjIS2tS2HS3C1Q5wo+M8IWsoW5eHeMVwI698btGZfdOOkW5OXB2fLBZKX
LCLSuW9raK0uM4nSzK7ox38VwDWrfpCxcyqjzDmDDwasvdlqxKeUJY6M0UCkkgZp
VjO4iLLp4Kk+ElzpHvv6BzbPKBNOkh/DxeCRaM7BeCkhRy97eih+leIayD3VMQTh
DEIsY/+0IIit1VL+xFfcueLi2QJe6vHTSqmuo+n046XrmblQseQq5R1QcFIUSURu
SV8bAYwGRDGgqYGdvwOeJzfrinHwBYn2HCcI2dDepeCNEiyJ2STj8dcfc53ewtbk
gMMJmGMcNGl7b70Zix4s89NpXoQa2JVCveqLiMlNpKaaEUPQTZPiWsXmQaqr0jhL
Vf9+wjewlpBNrcUYePZgkCust4Nau49fN9Gv8S0NQTn/oiJgeu1+s+VmK38X4Pd/
aNEMgEjbqb62abNQXb8K7nZxlBWHQ9fm5IiNtDDfM02idrQ07IgpD0ZxnsmJrGb7
1GlazKBSkpnIhAdpwf+YGZESyBUAjmGHGzwftHIFeQoBM9n5SbQGMSOLRGdi8vqh
LA58P0N9lJoSOvlbSSHvxQI+CMHv/6ca+UvWQXkPeY5DTxrwEBcnpzWOXiN6GHGx
FRjMT8SuSTJF+nS2VweQ2VTkIhuFnOwAvufsV8FSZ4ZoxJX5d2DSjH355/BnSgiR
xWNa3pC1yL1Otb3OgDUpveZTOsUBlCyIMhmlGmgpslcNHqA9ehZ8hWg7W+bT1h2K
OCb45elQz9aZ0GXOxH12rcMOg3qqw3zysoEmLBpE9VSfavl5UPv0hFNlkaVLUM4q
y04IXePyouArbdPVCVKYfImX4ajFTT0S03BawBVwAwMlaclpZ7bucU1kO0WXceQK
CoRKaF05ZASz5lSK8eDpunJhWz8D8hJDts6RqAczHRrG0DrACVqvHuc55+XHBGs+
fmCjQOrKosvvGXWjFZ/sXdWx5p9H59r07MrfJ4h7mFa/duaujBVPZg//uB2Qdzqt
ro6DisAt5M1FH4zkKlcYkqlsic4foqbgf94bt7Evxsm8rxkW7lp6baMDbtZClR2D
wAKt8v17QlLD+Opp2hYquC5qou5TNsWpmPIKLLEvOJtatsNZH8+CGNgvgnO2rrhz
cjKHMlFF6emq48ApJOo2IIlamCSFD44ty1rupu7Ec5Ebn+sdB45xutBVutdmXGSg
x5Ic4GZay3RiVk0hmQ58JUZidgAKMforQDCi6KIvH55zbSXigGDbbCGZ8yqY63yb
SppqfGdfOin38Kzkbw6bB9cU6NEthfz+U3SW+Ol44M97M6aret5p84v87XyQDzj+
HP7Who7ottF/3pONXi4/eLlJcHiS6ZpxZA1JCWpJTGc96wh61Fc8pFw2KJVp5R78
IlWQA0dBYn9C+scmM9FfpA062YeY6nFmGjJErWvZo29DBhEeRSByGqtetqwNCBPi
S6vImCd5V3l3NwUve/CcP01AXUq9zuTTjEMCcE3DIE+VUMTdTqo6YMFMUB2wDLdb
t73vOTSX0ho6W7TgdcIZDU8ecZmR3bVVGw6AAo/RRVEHmkBx14qZGF6fBnaiRx6F
DkazlVxAvk2dNdgzhBvnrI1cfU8/KTeKRPAY+w6tXgFEVRyqf//4Q97I993Lxqy9
cfhLCuwlrWjEc2zAJ1kgkRKa4/KdIExaub7VLFe7HkN88ub/N/YW1l5CGyKjWgPL
KdZjlNnp8Bej4LNnLovZqcjBw/pd3mPAdwIJW8IHQYa+0bC7jnf4kAMGT7BlLeWZ
QFAQI3INFGb38/u0UYCGHi0Bie8OcmZjCz2WL9Q2VEA++E0llsHVoWcSZDgjjOWe
g/TwJaCs1SElnseDWdJ7b3oTGIQ2aSUxeH6TQHtym/H11HnuLWUajhKtQLEhi7T5
dsk3Bl7nZ27xo1sPVZQe+dYTJbjaj/UzFqxGyH/E52t1vOkYL6iVz6T1di9uVGud
zCrQUoqR5fIScgs6jXfK1lQyrb4RdiJUm47EY3S5UO6XxXelYuSMiZuGuGHynQGu
zVdGpYGHqfMQ0/cXvga0gHLSnjO3ZEDX62xHqdb8gcDBBZYzS0rbweN4h4SFNz5+
8iMrJxeD8RHCUUMPR5WWJYCLKyaSjEePGqgOMbxI70WtgZjM1PiCTGB8EJcef/eD
aIr+bgau6j50G/ThO8CjnakXjX0Flse+Wj04AMu/NcR9Fzqp0buE3d5xVE9QOGAx
9dDVcldnVhuzMKQi/0Ctu+JVWV0MjrDAvn8WwcKi9Z0HqLCqhMrjHjCHKPLgZ6GU
aLgG5AT6Tjp5Ekac32+vUiQUzRkMs85BQ2VA6ly9iZxLPUFJQ0C0n+cp5Yfm2+oe
Ltq7A7BDz6RzS+hSjCZJ/UqBcwr0VIdYP28/ZUDVSBih6xYrW0WXNrdJLWKWWg/3
oZZV28ZU/REr7NzxV+w1Tzn5glddCw6AFgUWiRBCv/uQRq72oTJUG1t5mW7VtVk5
cV1Uxsgeg0Gb12+1IjKPQEw11QN/PMNi+IATcFvhS3yhlggqb9DDr4YDn91yh+zP
KD/k2gzrQf7+0ryS4Z0Z9qx2SpA7zH/vdD04Ra/tAUjcTWLbYN5r1/a8q3aeVinY
GhdQ31Tsok5+52pJV4wVj+IT0Fia2l17JS3G8kQTvJU01g7dn4HzDcIZrWWfhY3o
oHeg+RyPo6RZ2gfe2KytFhYYFyI/NErTG5PqgLHkq1x+lWhaphXTsfDoR7UOPQBr
qcfqOWAadJLm3iEJBLwsKkUL8yrZCQpEktcuyg/4SQA96rgGHE+zIoCIoJ0XAjoH
s43A+kHdRPIupHwEQFx+JiDuSepbXs1PbflL3pL0LTrcZ5fejhVlzX2nzRnS2Tr5
OlCGY6LpZJNhwKH/vv8sboCE/tmM4jOk5C+gVr/WqFyH+uIrPec8YIvfLzAOjPlo
bdSyoTg+8tf+ZgJwE0WBc/VanhGSHS4W0IDrBn3oxuahBtR8KLZUyQB0V3g8ZAyp
KU4kEmzh9BvYtgsokag/b82Ibd6tVyxlZTEDzC+ax81YRe7XoDHW91rjdm23b7mF
KQN2IOpdiywsSoR1K35dZ6zYBSZ1hjLd9AuTAOZ8UD1MAy7QjZ+JaRegzHZCrX8O
xGMgWyxLoFe7rpWQQV5sBxar3D48eassC05tQGbxatsGhdycc7tWPBOpbfv1lNrO
fxk9RywWb7DBmVL1CluE5bM+vdJ/zbpLYO2bv7TDElrfqz4jg5oWsaqarCG/19wB
eGqS2gGVPjnfak1yvfDEord5iaAJXpGBhNHUTGvXKi8ck8+8TEzxmngz+4r37k21
I5GROoX/2WnxN1/ICmQ9WKiIJFU9+c7stAPOdlm0TRq2mKhN5vBf5bzxJlH+tcIF
nJTmUH0zPpdQF2d3+LlF2fxigQpf2YUY0+jX8jU+hf00SVtttdlMcC6YwnDdFOzE
sfnn3XtoYlXhWOc2l8qfpzyk7STQmZaXt0ryUhaEqK9OtOMFI/Ken6SKWm7xCGOu
R8tZprPof5s9vbwjzeAXAphg3COYyju/OSvG7j59tDCrRRjQhTw8Ub9+DfmArneo
aQyiht8His8iEP4rKNOqgRZNEqzktH5YfKdh4R98PePdP/P+Gv8EBvWZmlWK54yc
paecRz0YGtnMj1H5kO4VCWl40xBF0yAmHuHsQk6ULpfsR08pB/BcaFjxgZY/dGVD
Mn9V0blBfQ8F9qZmmaoXb27/pdx/g/zuwPe2H1ZcCWTuVUqVMEeJDbzKXQ+zcWph
ZMua+xQ/4dwMQPB+CBTyQ942PPtOz/FqyAvKF0bMitwD3hYxx0UTkKOkSh9dpqMB
CmHLJgnrh8+I9VdfTjLa28wTBErsMTduM0z/tB16vtHZHu8DUJthn222gxaX2EVI
6fPr5xD3TuamlV1Cac8gLQoSaQllrwPFYHfpKSCLsrnHybkvkiOpIG/e0a/NniS8
OXuB1+WaFpwVSTW8/9m/isD8laZ8XBztY+A6SKoQjUuMT4oP4AbobFCH5U+8u6pu
eEENCJnBI8eBdWfrkT1hyDxp5+ZMgIUFqh4qrXukj/pTJT9OrK1twEB4O9kScemL
Qn61iaizL+Gq8KUwKx/y0OAcUFL6lcfpCTITnGlM7fiMPVRYIbmkO64SOIQmIYX7
8/WbpGVvQf/pkxY3qclzh83ar9DcqjXzo+dlNoN5suFgWxBepncBM0PnoHmRsqP3
5aMLamQH8W2+RTXdPa5fJ6LnIurZM7Mfa4z8RSS2QEkCnWqicW78EXTvBfmvdPfN
ZC/d0sjzNoBIbX/Vc0kbgnJ3DLajcQhTibCvcgQoyPmVhGSejlZpCE6gWEqvL0jP
yz5lIey1p3oRI3vNULAnLt1O7T8TwdGJbCYQzZZkO1lm5G0gJRUEa4Wg9ujcXD+E
3Pb0yqUk4lFRVBAu2p4cWY8nQ2tL5ZbkuwDOQvxJ074zwHxvp0KcoGB7MiMLQhB9
o/OyszaA7vz43lq2nQuXulYGP8kZA1JxZPVroEPmMguOYHM2h60eYqbaJ6TTMnGH
yUdc8x61fBBfokGA+z6scsodpFqWBCAGhfNg8F+6dXhQjDGGrUcp0AvXJcfUVYW3
MDmfeB9zEqhBc1AUtLUw7j7ZTk9ykbJlMlMEKAwFRb+I/S3j1oU2eAtdf5Br0Jdr
27yVHGry0qn0CDmB8WL75QwDuWu9ADJ0SSb/wzdyPyU96dDAy2vEmXODp02YNEuw
NlLlAjDJxGl2jr4frbxnSGYQmhpagMzumbh5SCaHQbyCpPl9azMHGhmcBq8Y89OP
F5Am283d4x2GNTT5IiP3L+JPUbsuOMx3w5GrpbhZWWAM9ICrRfUA0x8L/p1e0HAN
OfCQqle5cPUiOchFndapO323j3P8GazsL8gNOX9m2Sazum5KyOvi0+iy+rvjbc0r
9M86De3NaOKUtbi97dTY2U6I48IwfJT7CUwEIXrW1ASpKDmPKgvG+P1rIK7JGFRm
+gxYa31sy4cmtbxhp5InRa9oORWDFo1qTPkCqrOuL1FBRXyH9iBVezQf4bliyh1K
HJVyU1vdxAAiyJ8cieKAyCt76QGjCn3ZwfiZjUekWxVHun1viiq6EZBAWQuETgSb
MhRX6DkHFVJr+kHP9HGaSW72RuZxjcANsMm03bsojQSdTJHa/uAH9wU0SPGeT8ZE
OFwZsitsxdckNJLGL9mPkdaN/Hr1txdEHvnyCCvpMCiUXXzAIeA1cVvLCa8MRtPH
HiPZHAluW6KaTnBp2bsAnPQwvG/uVi38Ub888RPy0T0GzF4AAEBw+SZArHoBnGeV
sScYcM22SPVfylNTDRyyZ2b+hn+yTARA5TNe9eCpabPhIdOY62eJwFSu/vejqZUY
OEPf/BRmapxl/kMrbLohpmRBUfz9QQNxqg/bkOY5rUHlf3VwNfyDCuCyzSAlHJf9
7RqKTs8PBT1uSesHSvWBaN2tzEUpWpRGNVxgh6U600F3sTycQRyKrDpRyG+q2lkN
cMAZvxqH+g9DHZVN0U9cxIE8CL9nbG4heQ0HhQeWfikxTzfH+RxQylwLxDEF7/76
zo1pvIunfIA7o5PwYyGPl5Q35FNGKxlcQGUlMxjGWVWWo8Xv+QdjoyK1H2MXv0el
zR3xJ5Juqt3XZZIDO7wgCD3Y65SEp78P+dJrxtlslkmNb94YWsdLA09xUyfspaQ9
+AfFxccuNgayhYbu5hKYuCYZlE/RKK2yuKzkFPfvPtVlOQOP42GJnYW0n345U7WO
yGITk4KmvjP09YvOlbTTqrtiVfsbPJEA0WvEYGlWIkovNpXUEEqQwej5xNkFb2ux
I2jWGw+LI+P28JIBjcYb0Eio0laNqwEIRgKExDj2jefxUDlYcFJ8sfqH29abKk/w
iSBWjjaRYYuxwFxQdSRpLH8KVx1Bo255cIBYIE2RYeSqwAoYA3Jdle8Lvqo8oFs0
0QYepvCj8bjUHLWX+rLzVGdOIes2YgoSBSnhrOeUycc4TvztZtieAyKqBjhDbNPl
IiIwU5mCmWLyJro+YqRGMLkGyo+2tp+Qab5pxIeHnypE5WnpqGzjT3uqD+dBwDtr
rnuXd7NnQi0HegR2ZPNFk4w0PjN/cYaZ6PaZ300NdE2u1iD+9j4Ew+vDOgvHtFtw
PSDt5UOtpYZ1FG0tAlR9ULpag/lWWFeIR3IyV+OFYlnYxuh49OxhWl3nD4rI2m5n
qBn4rVqq85P5p1gQ3AZSzn9Vq2dWUBW1pDQC0eJxVHUAZ9/XA1FMyKcw7gf5bpW9
xnS3oVMQDaZysXnVLFdxjop3Z/P4hbBy+BGG09hh6Xa3VbrC0BHaGeG3JYKaIj6H
ICMqvMCgJfN4VOyZAzDvuZSFjJEpKZaw3rsNSLn19wWAgGDJsFP0IeVi4DBIo37g
0qQevdN0TebcBeZaGWo5AjKprV2BuG3Iumk9QneGv9JzjITJFa0iQTe2tImvgHJv
ZcpCVTKGmsDnukXSI53pgzjTM8e6Ku3/fn2yhGCg82HbKWCLmswlrIfGQKGV7E9v
xpc7jVJ0RysICFaBimIxG9lLCRJdzLw04WQ/qUo3PG79OU7A+6HwNU+ZO6DiYBzb
JQwWOVsRpEDzAxllgAKmB2+5hAG4tnpZEu/t3dDhXMB6tDb6BZJTTX6PR3zbKJ7N
Ps/Op0HW0yAuU95yZFvLPUwbck501roUn+l40VAqC+h9UaKt0m7ByLYXjCSzEDbP
PLYw9/3tIaYMuJKzNBvEJvszQY0Xpc4dbZnlQlqPMFaHXQEnMKv2FYbPfwLqsu/C
C9UWXwZwpAuBQUs3TkunCXvK15StePfyiomJvYaU40LwupQsz1if3pNDKctjmQli
xWST/jil5cGEWcJbZhZg6+TBR4c1N8sE3Cm37xtMxnqEi8YHF1+lksNVboACe/GB
fwrRO2PYjOdWOYx5q7nPcLCM5i8nsvlBYbicGRRCbp+7VRzAaYl9jTiBZFbeCWE/
Dp5rVbOhMBod/stzQ4IhdiQw8SNrLT03kE+05TlurwmjjGaaYjA1iITgKTB/ig4B
3VpdBwXtd+JAHhQJJYBfRHzjWy5xIlmofeB0pUL80s0xJ7Cay6+0tIcYBEMyRN3n
wQNPES9U4t6rgbUzjtoyqBWhRaqw2eydqi55/lbuU2jovV6lCpMMecdWYL6FZPN+
gLiES3NaqCNs0aQ/RJBvWQ8PjvBclvCXOOae7YyzDgfpYzV9i1bVFDt1raVdw4jE
rVw0tdNEYE9nLrJQ5PCw+pjmKWArgwkLjHunHV3NX3XzY5JMWM+V3dguLh0X9BEA
TGOw431qLuK5HNZ4v1BsJkcAnCVB+wY4Ygdqz0YnE37rbxQPIT6Q6D05g7PVp3Ib
dI0ROfPEs8Yh3cy0Do7c+yPTaEo1wVvwjKHmxOvJRplDMqbrDhSc87yAyiTYr/Ld
/zjBcqNbH0aypGRuiwFsi7HhWqs2YnMPkaQNImqcKTAj+JptbiV+rlAEB7K6XFXM
2FJZS20/CTn0kJ5sFeFNIV521rgok+Z3SgzqIrk2O/qj/iibw505sGnt0/oRmj7a
gs5zWnf/3KGNwnktbz2vHizrT6q9fdrdokFDK3bayNhL363SoR40UzWAhz79DAKe
ssvTWEWO0A2uygABYJOOIOIb0oHfmnrRFjH5T7hJ3uInH48r2InuRscaEWd5NSOm
MNKULJMDiCr4mn7eFjaEXyyROleWpLba2frZyO+7lPFoofycJev8SMbJftFtOyp1
v6Xbyb2BqMbtoqY9WQV43WXyx7lUQbElYoO4PGnR090QrpoO2fCc9fbkoAAQSEgc
KDd0UrC7dYJJfVB8iknqa/jg0DfnLCHGyRZlYOWLnmPWKbMAFJ2sswL57l46tYhB
Fp5RWhNGKZrY32Rvo1qxjW/z64FsO19WyulDfwpo/3hytgq2JGCyWjBbTdRpZf3h
DTQ9E1HNL3VnDHBkfVdhPBYpP7TGGZ12eyw+vf4bg7ZX4KJ0cNsgs/B/mP0PPX9V
hwNOyIvCgBmkK6Sh+XhtAcVIxfUVsxHIcy7LvDXLxOkT8y4egd2xWRmk0qkXu0XP
uerwhgGk4+FZG2pBpEhagtL3khXpMezEj3ryyu/xA3QNMMyxEJu7ewsMPTeb419/
d9kce6jGxGdrY1YIb/oMguGLNr7DZ4DiMnr1cXMUPUWKnt6kn7Nw8BKYvuYQz+ck
uNV3B3Q/xZwx2QDMLHXRpw9emtgcOHUeKAm5hgkNAOy1R7sTclwyaf+/IhUG8HEd
LNWtYavDPtdYCMzAPjHsKwdCuSmcNIVn5UcJmv7HEEyIMV2aOLOAabvJP8VWJXsF
ZbIwspUswMxzjV3fRxYDoUq4Pc/43b3rvU8fgC0X/sAZ3wdZizpcmpg+UaEktpA/
gPez6l1tn2M7uFvX6OglyOXqB1JUwrlg6ojJFSKjQNltW53/qMlPDFn/sp6EEYbk
uAfF/hiQTmE9HJXoa5ablpNfzB3NoTTNeCketWLDKoLpmeqMexNHCTbdWu+WhoQy
naPbl9Y6daQb26czEP/Tb6vflyeoGBuEgpayMDTU2yO4DeKReCdg+4kpU1kb9ood
R+OYHEG97ti5VW9ilEqxs6oO+XJoYA8VyrKi73rWOZOujowL/xIo+6GIDO1jN9q7
xpvNWx9dM3h/KN80sxLJG92GF5LWA2K/OXNnOnLKmgrcIeWEvaWZUvKjTmGuFqBw
0gtS80T3BtVmBqpAE17cZfmmtS8aOnALolayWreo5VPtq44zt4it7J1zkwZN89wm
lN8WUU4iwF8XfgxgVes72wkBRw0JpVPUaXZVIlA6rPTmZq1Sb0bBkLuOOV1Sxb7A
gmTtYOqRALd7dZjXo1ucUHiuyj3FYkrfIZrdeYUEE6M2bHSa7iNonPtJbSXf0EKI
qoTW1GQNMzxBEdjad2jAesqcJ3VGT8OE3IJtcfYKDARA071aOinPl8OIdmyxtFS9
GviigVtpKfQIIZvTBeEOBg1ZwhlJVsLYdtnJKr1o1GjCbxUz+G1u4mnVAK+aIfGo
PFuLyo+nfxhj0AWJ+28YpzQytbWFbP0YBqdWFxq2IFAQEjrOHXquW4Ekn+0NoeiU
5OHmrwp+XLWN0gdlSCVjOBoDJnrTeifNO2jEu5C1SRGKSXqKt9OtJGY907ZTb4XZ
jFhIgiQ/Sb7LiSMtVyM7zwC2QZ7aMJ/S7yIRo4B1SqGXF+QNGU5/xB1wA1XlYVf0
+FIN+tcOQDsIAevrgyI0S+SBl6uyHojnmmj9coGv90T8JEibcCjlAqmHhpw5nWEH
5c38y8Y8Wb6zhsWz2z93/2imm2ES+fgJJuBxX0N4xDMOE5No+mPqXVTTvrTdPFTy
Y24GxDzfCc5DDqVj1YJbAbVIC0VeR43+5UdISzil1XdMX+2VuPsQxE+4MJqVosXt
Uamhi+wcATAe7jlk8ArbVAhqvEzI7qQ+1q/qVmy8j6n8rcffFo45DXh7dDcxX+ff
h421KvNZcd8IYIDzJPrbsGXuQ0t3iPSozmHs6RP3NCLYECuk0VSpMaLufGUj5zUK
HHDbOrDZ4FQc7t6s0KJPzVj2nR+PJqQoqkNvyynmfLEGRrzQIsiww5D9H6TgbFc6
f//J8i/xUrHy7/qnhMdNYmcbRoWT6rF5ik29431EJz2wQmG1q1d9pnr6VeEl8qiG
FtTQmWt1vFijr5OmLjXVlvuKFWeBHtdP8KnNJKROLcj1dygqrajP1JOI3ESmRGN9
DnYFfqKlnsLUjxBgZX7mhBZ0tkNNTtpgcPYQPe+BpdwI8hILAT/cm/G46IkVnTor
O2l+rkZNUublOAZPbQhJ0BfvvrAQrfs/URg+nhr7bsrRyT61Mpo+FjU/t6wMGRpe
PMAKy3YwcAlICYK8fuT6lWrUUV8/NjP47yAE/VL1GYfilMeMzKCxPsJxTj5UKRGP
izFDlIUT9K71WLrnCGw6k6JVSQUXDCA8WS2tczfY1YEcroaNbg5+hcPzOA89OQcE
27kbd6Nr8LxB24wHKoe8jGaA4HNuLpbY7I0VArv5CUBGET+aw/hG7V++Afvum2Uh
iv5Bgi/ICb33G+x8PaoYjQO0/EdjsgInVdfgKbd+Nu8I4ASBj70Q8TNYyeKC0xwM
Qw6VF/OIK5piu/edsptJWRKEhv0g3Eq/sFJiPTblSTODprBBT2F/pPH86m2sILGv
xqA91OPl+SuzJTfwem4xWYEDpdCtbaJKZvjLARoCLWQNAj1qdJYVMjqVJMz03ALa
0ItrMeQMZFArUhCeyozylnauObHIzhemxfzxMVuj4YTQwPmeq9Gny3nHx3Cs8/YG
yGVEV0IDYigm9zco5mDJ51K6dbQ9tUlP+Np/u67UUToVnpNlHsy1gg772wWHIMvs
d9L3kjhDEtVtqxvEdOZ6282e+wk8QSzqJ1VzsxePvRaqa220ZeEFYFuORItT/C5w
heiPtTkFpNcuWhI5sIsMms42YBfWop2GIOQg25hRDlCLTiwAE8Ligmumd3zT+4Rp
f4oseeZVCqp9homtA+wDFTEt+qnLa/HNF77Uo6z6CxPXaTA2qY1+KfAFwmJLUeQP
iS7H0nopbNQ3T3do9LTS5VAE0xsYOUhuWY4JbPHRhL7Zu8V7bZT2SFfZaJQTBLhA
mxx3pRoQgXxTqmhVL+Myd6y9XmNTj61W2rboHAlpaTSub71l5vxREseK9PcG1aEV
SoychyuLGLvYB3wxOTfxkWF5Sx56XkRnZpo2nFuXNAkq2G+7VLJOwAJY0wpOAVop
5yyZyDoZHBx0wf//nuKXF9m4kWNawLyOa+isIjKDwNJnd6vsuUASvQAFgcNcmO30
A6QQlv+mcSG03P40QHz51HranEOoKxVjryYabyIpBuiw7cG9GjxtVYRgSNe7+9tT
rRS2gayYf+dM3bes5BooHndfMnHlTOVNEf016OAriDo0BMUTWNl7kPouTSOzPgmw
8NznUpuobQob14xALTCFgOJTb2tIFhCACd/9MAziQfLP9jTQ3DzMFTIt5qVr6BtQ
V3eeSBDF9g1NucJFy4u5A75/dFndc2HRvGcc8N0bBcK6P+dfhXYGxUBWiMBoEYEs
UzNtt5hPfqaV2Xzli7dyLLH8sSyzMu6MsFEySLmmA4RNd84JmJfy9aXb6I2Znzeb
adfn7W2CctRAqgYq17c9hSqAxBdWn0vlLHpe2f/6JGOyNIRqPG3+o9p8Pa1GDBki
Be7L9NG4SPhXfxx82rnOw1OBc66EpFsZQhCrVGciWYkFXfiZbu0i1+DlZx4xZ0yo
YxAL/qGGfQiK3vHyqoSp9jvDSprRiNtIiKuX8pdcoWOF6YA+JrLOO1msvbWrIxWl
uviMI9P9XRP/SFwnUlOVawE5SeQeBZQ03Ie2mwJLVlE5HJU1EpXNQ6shfs5kEbF3
oH9Ak9qXhUwQpjkk9ed/alFZ/8lRrgCCEzP4QH6aZMHI419xJlO1WpF8bc9G6K0k
gUQIIhWQPn8XF+tYJ45uivZoXLtelfbncyj3CiOXSc8fPzPnqJFsNVp3FHBporF+
od3Eu1EkjAPU+zDpIEM7oGPFkRu4DzO1g8lPZCFumN6ROov46sAmehWPTnbXL6tg
iv11Hog3bhHD0SoaNwEaY45CPgRgSuszesQhFpCL9Q16FZujQDDsA2dpH3/1A0TN
Rf+gLGAqrKwCjnoqgPuNmYzK1MhpiFiS+UqTH6K8AeQlWDVejHjEIA598vdN86r3
C9j9wnaBcKhh2lgANAiaj/Dtwx/12d3wN7mwf8zWtK5kx+hJ8joN29/wKCn1SJJp
kSelgXgEaWZSXO/TTE0uyUifPEULbEgNEsTY/OtYPp7pZBUTgi3T4lYQfXpPmSKL
oK8u9BLKywNUKWiifeCYoX8zu84x1IRDdAPgnzCySlJMqzZ4jMVdSNrNoWQlAivt
vxMYxx7qJ+stx+qdzY9LEFmWvDsmtVCuJ3kez0FQil7R1Yis1ZswHo+04cY7qzRX
cqaFZcRv0FHFULEKzPtY9rnTxtYu5WnYi0eXbM4FpyyUslmP3bsRHpVppAfhN1lQ
TRC5e2PHPcxQC3TCjd0P0nFpncpUNckfRmcZ5PiWd/Y/1ZFEqB6tcq5RqOn5dGof
b8sra+yXKTfdrZJm4igiYHmKQQOoUXTe37+WE0c1DW9uIdqTHbJCQEpJtWUYr0Rz
2OmK5FIpHBfUaAuVlsR2W6X0m7J6zQh6zKuSWIWeMPKutJMHvAJqpKnB4qdaTLhk
+QDKiZAJIryIQjqRzErPVSYy5rKibGr399Lwe5mudyulbqlfLZNoKUT2jigJNeC8
c6jWHM38FrtgPKWNeXmBH9d7DtScD5UbxlU1cA/0VKB/Cho18MQWNeL/vrFu3Mv/
SOPFtB+UHulg3f7XS3PnFPfvnjQWLpplsehSaW9HPHa8ufS9yiXy3XJpZ7QnxXPu
Hpnk0bffVAo4JZZ3KGagxmmlf3q03IkIQba5eaDmAV2xzfuxaxGssRvoPUmgWBZ7
EpNLLFD38yoDTddh1e3x+AI2V/sxsQcphbLNcTUshKFSLCwh0PB/IVtpjxPWp8pt
/5T7daDdlYFVtujix54QAOa/urdqDeKw4VMmsGTgqSlA97NAcYHnPz+Lxg+TqxYb
kY56wFGb0GueklBMkZOrlA7/bBBBxk42mCyidV8EqF/YcLyYtgGwp9fPAaSDTVRJ
ZfCHcn9zaKXWvj2k1d0W4ZTk2C391WF2+0JSkyV/FUF1avIZvz8hbg/QJczmloIr
wCiOqb/gtT89Byb20px8WX/cRR8fmzhz6MzUIFGBDkD1XtaPGmazkaljn4IJdVK0
+Qf3perEy9MKls7nXCRA2eIf0baIDE0elDX3jwHmXNfXDnY6+sx25km1Z+cEs+Q/
p6HZNpK0Nw0/mv6YCRrPqioyYO+XYOM7vHX4pNB+IpiHCsYOZP9C1FKP4v5Kbfvq
RMg5wICx6/sfLQjwtUgL/3UIa3KBo78a3b6LCIhm6ZlDQocndQVD82vgpPukHh25
KKKFK06fMyVHZlWEZ5j780/1LR7jtlKoQHO3EuM++yS1yUMAUvmoKgQ0Q77awLwf
P6FoureuW3nNF2wvTOhwIb41Tn32wNOKayeGPJWo4eysuns5C2W8ym65yZ2028lq
P4aq3GPW4qiQLfN3GSxYAcmHkwGPX82TNwKEZr+6UXWtncVmqFnwb0Z4k+Ur45Rx
OOep4tXZJxDqyHhQTaBZu1g05Q/TnPt/QF6a5ap52HUWd+WrVbEka9BVZQbYUXiG
kK/v9A6Sfsf7LC1CdsWo2b6TOhlMmpiXXG3ylGW7SBO5zJ9ZOgjZJ/49EZie/KK3
Gu0qtgQbHGXOuOj9uGGqdZ6p/2vwFPODxuZs0G3yvtyt69mscqxuVUkiUpN1Rd5b
d04+4/S1ruAnk8QT81QXVTbVjZkGpniRiC8SbI4mwRJhR4DG2VYHAynuUC2lyMhh
s3ViVKMkozxFPvU7+H4DJSoYoLahacGAApD/iYFPGbVaeNyGw7NnWxLFehTgmOJB
e09xXkbc8xAT7+xlKcxdPusLoZFEA7yE1I2ZOYQ+ajknIO+uGay2XpFtX+S25OAP
laDVnEh0b7QRFgBTYxYlOU7LOTrB8UXwfWuN1b8ziVmDGKYk9jCTywHNRB1eITPo
ZDwc/wy5bvOwukvrqiDxy6TdThi7GN9a2MSTJCbfXHSmuSmevqG/w/taoassLxPD
E9uBi3KGuTrHT2CLy7B8RskkJdNJ4ep9WItfYqbBnrK6a+j69t8kVjlebnMfBMok
5/kZHLMcuZHtuHNTn+6srxgc+x/qZnUs4tVB2H+udMOiZVLDrm56NNF69X6fvucU
sV0BgDapMoDNlHIwbUSuFm7/RwQW/2lidPsADp1w+YMaDgnDdXWOQDZI2TDC47PE
cruzUfqa2Bp5Qr1IP6RKdowOgpBiMzqNSh+2drv8WL8SHHlWMhLMyU57jTWBe9UP
U6DPQDALtdj4R1a3ggDHxG6aVfl6pkgnHprbRTtoUBbZnKGJUYISLCex5ohB4exc
A7ZPSHf80eyLfV29kNC5YJtf07bZuQU3vIZhoR8GQmVP2tQFSLrxNwzzjCB8B4mB
cuMIDqKVGHraw1kybGmWYu1bMq4EiFOG1iZWteaGe1CKXoXC8bMIzgnqQzAieD6y
hSWqI2ijqoxLTPfH4K9zoku+yMcjUWJH1weredQl7C5GI8cB35fN1zKvQPDaXIXr
8lxWM1N0QHDa4GpM+LmpCtywbu3n5I8krdZEUfphG0WkoJRIT+n+f/LbF61pwarQ
9UPvnls2mezWh7aQvWrhtiPAw9FGY2PceP44YeoHQkJXLYcb7C4wzWOYSQMVAI7p
kSOB6ffjcyVPti3TLyFtEywCi0Kv9VAMEBBJ1sz7U9n5w5I43asEiJ4+OzuhbYaL
/tWoe0jGSVldU1t7qpAAhR0bo1bKHnfd0I/x8RE4JBgX3FZ+l5ao27swgAFM9yBQ
ZS7dWjgNU0mdQomb6VyxHrgXh0uuocjgIJ2eUmkRZf1yTopQM3DBHzkIx9uM/6Uh
uxiFarryX2BWNILqBoussaeK9fp74kQXEPnnn7VwZMpryDgilI/Ewsyjogq6Iche
zj8lQINvfKWesgSn9xwMFcxmNUOgKZFp6GbzpRd7S2IHwZJr+5skghWMrgjp8qYu
nNEkn2XoSHxOoMaoFQ3jK4mJdfYGFQqzoW1m4usLd+Hb0OssOUws/8uRszr/sgQS
ZRA7wXUZWWC1FAyNplfGJQX7w4/KchPUZtzYkMTMg9abVBk2rMJxDrU10LfBUzrK
jeQXpBg2ftpU/stJsu6QMapqrpwQjPaC3+7I4rO/qCY+RfN6URJHvw1OImuRp8/d
0JFDYwxX9+5C6xJC1bQBXQosck+z55FhS//8g+hrCwbGH1pyRpZXupAQlnfhUf/F
DYPRbkI6tAUt5oYsLDHGjF21S8Wwika/chWMyao6YhPUTcQQcU+3Ka7/mgENS/Fq
Htm3wkRYyIKdDcYY/dJY84atAIabMRhqci4kL2YXxH+3WTZ5LKyu0oDLAW5EXFJw
y2EjrsrQqr+Gpz1AzmmqkIqHi+Jxa7GR6UbnKqN5gwvxr4OwHJh4LnxXXiN8NViU
sU4JBv+/AdJaA0EAFhyfm1P2N2wTwkBCFbWUQ2edqpnxqrsNxyT8QMsmdKl602h1
NQK1VXD/+pXXWlNO0XEA9yT01H0RyTnrMPk5x4nWjSQPsvzH/cjtHUKcxqQGzqqi
/AShnUgK27vmhik/nlek4GlMuGyrJuWO5pkDo3FvwA0eAlSXfkCKO1k1Wne6KHQH
4IaFx7dN5paC5V4pAGxa0UVCxSkL5YKgUIeUVBWsqOsfvaHSiA6B83eN2KGPPgXE
R6YoN8sRkrUXINWhBkVsBkJbfxoEr12sg75bPH2WH1+tKTIT9NfemIUb5LcJbzdK
rCoC9KWMpAddZJNWPdQJSIzn9p9oF3KbYXBhohCRz2kAoJ53xLWGQvTX/J+zp3VN
DBiVjtPYp7cawi1/YU53c06cYuEwU9/KCQGx0HufSAk8PLwEQBcHNXrw2EoycuA6
0laMyS3wp8n/eonDwI6h+aR+4sGbwKPRv8JRgzHho1ay85YNnOk8rzqy5MuLEe0H
UCHIcWK3jtPC6aSGxbcisGoWG5GzWQ7nG3fMIkHjCVAv+lP/iHWHDT9qzMqaXfUF
bxkQuCqAQuCTuCGOAdnga9S/DgFGCRVa65+2HdUXt8+uYdcx1waE7phkyii6v/Ua
1DTYfD/ifgDwEWbQm0aF4mc+ShR9Omn4Ap+9UVdn6zYf/zED/oPOK1fYd3Mgr1tV
aRWQrIciS7TPLLPotTaP9BGdkqkLBzHbyELwXN22DeuzbRAwtGClRr4AWhJ8ZV7h
nqvuLTZ0+683TNp1EhFc1UL1DcE6aWnWj2v/EctCq9sw/eJgaxW9rGkg2JAjZkMg
ILZ1+UaRgWmggEqw804PK+KNISPnOmAdoyF8nNuiGEuZcRueYkJ2FnxtxwgbIAYK
/gSc5Od4vaAPK4hj1X0CnYiu5WqJpoRzyrhG++27aRCWTH/mxwOs+dID4iCaEcpJ
9IAzzjdUBnpXBJTOk9v36h7NeidrA5UOzYHOPbqeSuWBbtXEC6IhDymo9aH8vDTq
cv7wEbup6LJJ6BDXup08IATwh+F0JAywyfjc83JfBxev4Dt0RB8SL9sjqRzww81/
Eo5IOCzek19IBvg+ebcKcpa25Q+oDqKmmComXtqnfk03n5vv52ctUWlqAhmybOCl
nyXjOE+PFX5Ps1FAdR4uR+bblWsLFAPAl0+mSw6aJgfuCp5Yc+OaSfL5AV5K/9S5
IIVTr+Yj/VLU2lCPF4YMOXv1/ARB2jqiUaxCg5rUFb6ImQ4Ls33ecBlrrJkGsL4D
/Cg4pJ4q7xtoIzCEWgkCmvUhUD/49F7vu/f8xLUtLo9llMmq71uPo/xykYMOn/Iu
ni0EgGE57kA512y1FmtyoML8HOKqeX0ETmyb08l8YU5HYiEZ2xgdjgtQ2RtHv9ml
GJCReboRZNR1wXzUUUmDegCKaCotMDUaxBKP9CQdVzjxXfKttL2Upe0kV/gqfwul
WS45z2KsoHREWM1wcPa+6AHdjKC1s6MpI3nCvBze1aInDxf5mNGxOfyFnJc3mbk5
3XaQAFGGJUAknJOb83jXXHPgKvLct6BHX7YIP8H+TgyO5rMS6DtJy4LiWkBzW43P
1orRxjqjI/XPwG/HKoiwVAXPj11AUDhqIjOKb3CZuOlV13dP1lWb8c9L7GZYO9pU
skmVNiv81vgz+oGyGpamj76jEH89DQE8EcuKrIGPpcubV0B9cFaTQLA65ZwtC3+b
dMHHqynqlX03aRO2kMF9jV4HCLOMA2JQStSindb4TLHOV/e4u7BhO8KrM+MKVsjB
WzxmsVF2eanmypb/xxqH9YsJR3Wy9wBhfKWh54YgtTA+BPa+HMFCObMMswXt7WO8
j9ywjN0BGnIDNWXXsF5fyrnMQE1Uw704rwJrX5eHvh7WCVwfe4R/qYSAVC5ADUSS
xAJMZsKYK2UGEILljdvuZGK3mwudSDA2hphPA/Z9HU0TINPdC+mBq7QTFMIJ+a2z
4+RqO1tYkRYEUU40Q7W9lQtAeJduFTknYhRp77Lb+2u1196gtT5rB8dsNCKOwgrU
3kvrkY+Y3xh24pnExVyT/XFqB2t+7qPM4yrwoml3v2IUJtILCYOB+3w2VO8IDsi8
S/c5GATocb3T/cyCEfZMrHHey4SHKoezMQ4iDJb/mzEY6wRQ9meamrK9QChWaC3n
JMAAS32gp8jOgLqYH0ZDoO8RgxTnzWZ112GjeGXq3Ik8j+O88wKB7QumgiXcXMv2
/IOfITEr0MRWQ/SbYVrd4w7m4EyxFlXILlnqpPYVhpSVVrrxGiDTP60Ig1JtAFtL
V8lp48NfIPj5/E86egRyxFZbEKOCNUqpEmvd+757aHRShnhg7GVinfQftJ6xKMxe
PgtM1UFTcIQWSZt65QEHSZtYG7BIpi/K70mc/xZKeDXadqzPZl3DbxawBnF/mLfE
6G2gvXjr8HwOKbE4LzZax/ZJOYA+jqGDbc18CSOor39oKlp+rzVPGg56+FHw+D4f
tAPcQ4GRVk1WiaaBmomO730qzMyX020z/Xg/nmOXlRSyQyWu0J2tS6gHEvXAJ6MD
9Nr1Rh+KimjGJTvyCGGLf25HiMJoywBLP3qeebquyScAHn/QMKwmtBhwX4ulgGhG
A8nWRDqIf+CvPwe4ZW2+WGZhVCNVPMOi5qNRiTbaZcgD5a+b5HqjqaEPRs4jWwTG
wJ0sEqrWY/9pm2u8Yv/24tZ9cvaRBu/zf703eHp+9ldZTDZ8XzFZmKOCObh5OMZd
pkQ6IcSAFmv5fMzob7Jm7GBtS/VWYwsvhDvcY6gIY/04kglCj76Xu/eQi/VE5bts
e6nO7iY08tSmlDsWeExn/g7Xr9a2cfwswVtfRlnX6LnGXpvxiqbXd+NtszNF6ny1
VBXUZbbL+D1EndPKqcEM51Oim3SyBieAQn6xWm5UVybWxJq+k1aDymG6Z5oYa1lK
fEe5AfDu7RaKsgJr27E0w2CZjkLNkJrmpz2s6W1vXFF6VHy2jPzUthQGSuLO4U1d
9c/9O18CIdVhjzTCIIM3xbMOgoei8k+7hCRK9gMlshkTMXQ/idYpZz6bYgGFakDP
M36pyLrij//VhnPKiJ8wdBdZC8gQ2GxSj3hkMA6NM/fklhIV2e7dfAFqJgz2HJos
jCMoXl7wjO9dJDLEkZwBzZOIilMhUYHiQMf8BEaZ2fL5NJ/FtWCdfo47YuftzUFs
PmCZSVrmluFliL/aZHakNiOtXWhJV16d75iHWTW8/JNl6cloQ1wTRm/YBoiblowh
w+ktUFc/NAkOwsE4UZZvRsokB/q0F9fH7hz862MG+3g1MXNtfvMg18m3xj10m8y6
0H7eW4DevgnQoO7Nr4fDZ+JR6vhZKv9GyVtdjzfTWysWKrMavOkxvx5vAixbsGGC
eYJ2jvA/b5tJVy+XEHOr8iCmBjQaBfir267llJMlP+l5zEd8Z3iw7OXsrZQL1jjc
QYJyvyI6+xWb/cmtClf2p13Gt37jlpyfJo6k9quaOgo8YpYPLzbDj+nKjEpIZ1cj
oIZD7rw2q95wGeq1Tbt/CSws+SvoM8DY/bGMmKa3cCISeqGXEAdO/Tpv5Z4lXwYC
Nw9a4lMwePfBTVS/pRlCiNh+HLDWMuAmrfXXkHL1dEJ7udlhqJl3dwVUrj13pqWN
tALZw1J5rb94NwW5NTFF2rDWUzwTqOzKMMHUz+Aq1oFHZP9rvtiN8VQyI0fTAO9A
pXZrmUyO6S7H4pMHrYT56snvy7g9b76gmTv2d2sOsol91CMTvhCxOzavvSc9df3Z
DCLiPSgiF3mEwKrPD8pZRC1fozbPdYH7HczEoApTLgQKv1zE/ONYa6kBFcOtG2Ib
0Y375kutLE02Sk3uIORhSDW4b4Kxqn3No4QOdN08abnvT+ED9BVttAL0/SDjiV3c
lVJPgZGRHNY5pbTUOHQgd06O0PuYCSJx0c0B9enh3jE9fnpIn7t7aKEMB1gNdPye
PlPvja5ulk36QkH5tfvyb6lPJJulReuRBtNLepn42lGSf1sDuNcn46XdQEZw4TkH
dgF6lRlUXyLvWD1nkr/CaEcV8k8D21BOUYtuEeY0L4R0xZkBwW+rwiKKZMFwRpJt
49XINxazZ8HlvqpYE1Q/U3sG5fG8WOVJURO+pOs2btfKBKREAMdOXK2FCqop5N5a
DoyUDMk6J2uAYGA6E8RJc8bJXCgKjLGnS3ps3LIVMFP8jdpXgKY9D482F4JNEsHf
kaM6jJU7Dx8ISoBV+O3jjiFvc6t7JNUAsIpbfU6c+M5FXAMh3P6I3P0EWw+CT6eL
PPriWqpI04rjRqEy2qUDUErbuVi0zrqaIZ4IKDELhrNs/ZaSBc3gmpVHNn1deQZA
4/c8VUPgUn48tmgBbUawZ9GmbqPBeBsU6BAmMEKdRpqVbrdsoflAA0dpi7gbOaNE
rC+kygGT7zR1LmVXFmVP673+7o3xB+T6P4FAPLVCZE9wI/HE2MfdODT2aAtx5ipC
l3W/ZBHMs2G12nzCeJVOt09q9OjLGVHIXx/z0QQckvQDL/4l2HrM/4p7YssJU5ln
yNAAo+V/KWkouuJqGMG5O+E++jPPC8I0huiOI6v9AfasANUQcEKBZQv0ugXeP4K4
ybPWjrYey4n01rOTT+8kCgtyaYlYjeR9R+FcYa3onQuybm0xiVnc6yi4ETQAshoI
CFVfpoLFFwUx48s1XqMjpkmiBngkRm+KgUQkc7SRBuQrM8dsohcNSFJrNL9Ith/P
4MftQAy5RAM98eqEDeeUPPPkX17WJfxxCWVI/sfn05TzdkqRi2fYTxud34l2hDer
qT4XUDGz8SiJjPRT2tHzYcF7UaZvWtbSVTwSTGiq1V14xciqc+sS1kiMLD7FgcLX
l6iM4k29drkfyH7+kzEOt0pBulX275UnyD5OB9wZFGqv8cJBJtT++MVm3LVGDoET
Ce1PV2DajxOkMYcnsQ2HOxn2D+6tEB32Q9bgbqG98Cy8xrF+6kfZWcWJRCPGbkOs
/AfZAkrRV19YKV5cYp8WeinPvO96ITjOLzfSvZAi95kv6+L6skiMITBvpqZng2Ou
VeT0ricv4xfGCM9SUUwMmOJKQdOsSXc2AvaZ+Rf6QwZuc/yxZ72kQomFqLFtQmUU
tl09qOamClKnyQRZI3FQP6GI4bE4OhQjdoWfYT/K3Bsx9a0lk7Gh5f+mD+Yf2za0
jcmFYnVeFTtVWbSIbGERaQHOZRw7OONSApWj5VhtSpUqpdMdSA9lsek859xbkj9K
YRi6krAIDL3IcZWqgKt5fC8IEFUS0Dq81lOfF2tbpZRnc0/ggoJH/p06wH1iwWvq
84M3G9yjkOwaqkYVXFvNltHInyjsUs8pj8bvSJbaWrVJkPC/lFVros5BZ8k6RD3Y
d9B4cP1DiVfB4N2n+qRIixSbN9wWiVzfRXVbTiXdvKPr9jmweuYKzj4THLzTPp4a
AqLR7WKP5too5Lz+q0rJIEtxGOk2ayaD98wiCatvjeWTSUB7YvxMXDAHjDXBHnqS
ZbZTXek7hO7s8K/3t6z2gfHeeeLa4TfcRKYUkm5G5nOnXxfbLD7pS+ApCh7vx9wl
0hbG/k6xXoccF0vgwRwzP2OB8IggavBc/AQQ4DAJjw/ySoN9rdXdn7kYjL2HYLNO
COdC+ZI9OrSBUbvZAlbf6rjMeEKv4oUuHGqP0MasMwK4uIcLsJdDHXSxF0RsFSR5
l3/z19/W1IymTmlIVB0K5LICCQn13thxGjjZomNW/QKxQkDrCqSNJyLKhdSxYjwf
7kJFYseUE+zeyAQ99/Ip/+5OAVcmD0DXoF40627xp/jZkmb8FPA7lpE4ofqovGm/
CitOzwB+SIK8xn43GIYyZkPREuJSnXH2QCaeszFgtPbzbd5HxilADPaa1IKKBHsL
PgHpOhdHo0uJ+JtHYqsOufIvAXqcBuhZd5W5j/1jMP0dF6jOAf/lvLIfgvk4Hii3
IMZZTJPs0vK4slxoEanehGLRGmzLJLsniW1PGmvON3qSvbWbBGgsMiIUkxu7knQ8
uZOBGQJ9qsAyRet+D5h3zS0tpftxkWTwBXuAeAUrHHboFZuncQvRN523Y4I4dEui
z1duF1FRM1OkdqWOrCO7uEdybUTbF7EVn8XS+woAd07a4wjsqkNSJfIgY/lvleMB
g41P+fBaL/0u3sDf9ZviNF6XWO1Cw1r2VhOgVPsn5oxR0xD6pLlUPC90D0EmEDqq
pH80VExqeQIcbURVDrDjFZlGpNpXfHlJ353vtKnUF8yArs/9XoTr7lVUluPS/Wld
kjEKdPOJa15nBBdRCN4/o8a70SDrCiMJpiRIkR5jA8j7l/Rx7Pp6Qn3b89pZwSCn
qVt3TndLNhW7TvZTZOd4iQfsU6DM3j/OqQZkTYFkSUrLv54N70rUjHxaamyd5blR
BlHQDolnG6x9KxQpwKqKZNxMIWppLb4CNW5YxYvkr1yFb3o1Xm7yztEbfNgDVzGu
iGST4wx2V9+Ie0yy9OP2cso87cvJmKKaDtINj8ECt7vWReLap5+AngvO1liLRTje
6+u5o6/Pe6dCQ6HX8aAHqZusVqJmZ4AyeWTQQPQwJKCp106mMQ0ynD/Sheey65gN
7kTJtnM6l1YPMU35+qg1AzXfeZTQzjvJtGpez8YsABVMBGcaF88jnO+AYSjytlbu
zOH/3vfBVj749XLwue1lMqn4FFEtT1HwRXjuYmKNfinMkAS6K9XwvAZf7WXGykOj
gLQ8HbtlNg3aRb+mXswb7ee37KVtJB5ztTjM0ZLCrq1MOCN4J8uqbF6EYneJ6uPw
qOelJ1je+6dzrJ/bLJT2tDQiQNoHUqLTm2bNIhyFeuBtSsXrXvOiGerPahhOYgjZ
TMpQNU+sOTNg73y/3s0KgldolWEluDcL/maR0we1o2NYV3FhgFC8GP/aI7upbHj7
jp5lvE/8/cXLhHFdt/yfsnFMYYjjM4zDC+SWwyROd86zo3iJ5Z4Ak31t1sNVkD8B
LuAE7CEPjyuIQyeiuanVmWBw5niIZaMFb9o8tiLYVidW5b4BLMd/oYGt6mU66jxv
0LhKBX/14n7n4tTPOLhgxCQYkcbejUzkekuXELYxkXxn9GgrPRqakRkRXh0VwJNy
5mlgF3GAWBvQHe20Nc/ZJmzdDzaAgmnTdaqt7zG0C94SxmVHwV2VnKmRFZflrv/V
/HX0oXYzrTdDZ03qjfMerxNOlnTBM4r7dvT+1GpNN83A0tD7mllc+z6GgGL/zovZ
hYJBal0ojkWA63Ci8YEOdfLWRp1ZkF7Jq4tbwdBQ4Mis7OUBernxsgQo1K1Yt5LN
RRHN4ch6TxUmFPTGNJ9iHRHDAI6TPlYT1/LIOZo+9ATOqcnu386ZwTdW/+KIzJ90
GtpQ+6A/OWoXNkbIVX0bL3gwYwMxXbxfABQ7bWqixXoDdViqXU/i83SZ/3M7UrnN
kQsKgUdoAnSbSSQrefgfKSPhMIp+LJhbni1tB1cSmTKJMOtUh0TcdaFPSEXeSrKM
pyO/+YHoCoPvSEuNUbLR6yvf0iwEOj/rKRTqrn035bRhGXfknMlq695w/lXnVTaE
eFK6XFnfDMoKIYLouMWqDWKp72hpvktemZlPq+lf+OU1ZXEQlgsPen9vKMd+xWyL
Ka/SRwsgDDCJ5S6FFk03Vw0jiVnUW4GViOyVdpxX9gdL5hGc0bIdK3wKYzBUsnZM
aDHRiTqxrrXdATpDDOi9V47bzrNbzmAjeENwTSMXxfsRXCbJPXvgd/sDdITDvr69
EABGdlDCbSb6BRzISflAk3j+/T97+rVbTv2d4H2hq3RAu+8xlPe0+L4SE9wA/+9o
fuloLASpRGz/CQU13v+cA7/N/DxBPJSzLM4YSTVEwyrzxtn06y3V9j80nYwa35Ai
kel0e3dIuEEdHdB5DagOCr3+AZhcBQ+ZeJ3TUgQ5lk+prp3LsvjqgQ5CKn4KiyJu
JFTdQaylWAAX9Yi/y3wqtVPoFa9skI8YSfVep89vteuMnqFoquWMds+5EOEw57B4
2nSvBM+MMYcPByBTdeAGqDWoGQU8hlIhL2nilllNfBEnI4edeadQ4ExeyvPE1lrY
yWd1pAKgNtRf7aOfjhbTUhkDFs489tTGATE3Hc/4wNCB2XNjk6s5JJM4rwxkBAWi
kSAsGKZPPuP5+jaLNej+b9GThep5ushZp/E4rFWPFSaYtMlwNDkfWWdtjmCCUHyA
cjQSxjheX9xPExrVBAZg2WWYQQeu/5ZyAxQzApEFo1HsgE3/KZ3YvqAuKo5chXLF
3zT8N2Ff6l0CGhfswPgqS3mqmTGuxdty0kijrQXoIazF48et3Jwtqi0KCobA/Q2q
ADVDbEzSIZyAJm1bwiqCYro/chFcVTLI6pFxIxrJ4tZv4pmtvBZ18karWA+F5HU8
8Vq+EAh8Iokaj0fEDV846Bf1I/AtRxEt9E4682Dn4DtJPbo7vIDXNpq5dXhRZAtk
RflI0pFb/tITov0cRUvJbiiXiaXs4Kss/dR4JPUoIPYLusb9NIA0p3AsLRUGBjgh
tihR515600Dw1YDwJ7v5dwJtEtoHLiJAepE4JuMBkDzoztWvW3RkNh2JXLtRoaKO
NVFSP9XqYQohiHhtDj5cFiN1pbnf+M8F3+CUnUxDG4wj/9vay50Etc3GufoJ42/u
LlfirQpyeBasrEK1H+D3IqaiHEngrgGpxLUTIVD0WBubYwsnSfKYtl6JlNwECfaY
ubffrPMzx5M1RDg6zQFcR/9IZpbhtg7vTbaBQyM1XNm0PjFLrx3Ykty07FoVXdT+
yraCUOABbB5lNYWj8j/FraPbMKopN1Wjf9jCzjjFMX410bRtavqIxGfK4m8P1TEJ
Ci0z6dEIsnX1/Hs928byAbxPnJHUkDsW1hFA3sW6sXuVBEzeKjD6/4cZFxQwEXq2
0t37fXd3qLZ4+xx7bPcrwCUxbUBiFItzddjUwlYJguudi6mCNqRf3gy+ruFIdMyR
v0irwVu3T0n1azACU5id//2T75NTTTAbMN1DcJhPZTqXwXXLimsdKRe3dPKQWBQm
sfteythnG+hylnTRYwHiFkxsWREN4QaXWpnGadT0J6PaC+UteUWtKyGBocV9Qfbd
xhe+xTM/V7dDr0DQxQzNIE89wlAINrpCxGa5Hv06q4SHlrDV5DShkS8aKhByOs6E
QAjg9QogAwiVkVO0D5zfc1z9smn0j1CQS8Bi7VQG2oZGIn5g3+Y2R4fhzF1nGQbx
JRWUW4PJV1kzI73EJVD3b3RcXA+btHu9RSt7fz8WA9jGW2JztLpYmsdJwpGUeTSH
CK+kfzbrS2frDW7iAkprtF2Kjl2js1qH8LX8AfzquKLpe3eyf7pGTVnBXezgkpcf
cx8mU7L3yCMIU0F+DYpYIj3j2SkWCdMPHwy7imMrnIG6oAIP9SO1AQn/c7JXdbB+
wQrNT4oOXxh9epRwquZjBtMUs7K39t+5aCpaxM7A+40Y+n3IPSD8DpbHLFrfJkXe
EVbresEquDvlocHeCF4xPB+XyHwQ17ygVjF6hWMg/xXl++xtPPWN715kJYtUVjdL
353ZtAcsyf8v2C/caHYSe8zLGvPxs8maarVNdhJLd78PRGSMoAFbUu98rHOwiE3s
QQzZ5dWl2Yo7vBAAtIgvGZ/EDpBOPPaeMGRNzv4OFV5fF64llXSM4vsmgi8vmtZx
KssiiRhgg9IfWv0S84O6A0V6r2W4K4a/decL6xbLbHBlQUBm9hFdDtbgGa4iDTFR
9avJgaW2FkZPsMn0ohID+FdyNHwsI1t+5XXrYlEvJAiIR5knq6geY1RMq6Cs+X61
lDX5NYgqPizLabcovMp1dtbCab3qK486fg2a40LdGCczZmbpoC15+qP51t0u6AeN
zdv+4ltloWAzoEQHeMLupXGGh7fayfcJyolsXUL152Tp09qubpWrHJEYwsDwZK4c
0ipBNgFtRc85652thdaqcL3ggASnSZtsdLsYb/gKWotGRD50GsZq7fWj+ImYe76T
vShqpxscWvXj2yi9ksG3TMgD6zAw9gatS6F0EnrodjyHJzLdmz7IDs7PEyLuzoMa
ooHg0j4Lqb8FSQvy5fbaU6TfOFD8C70GtFHeJ5UNqLv8IpKu/kLWXj9lJC7V/rh9
ATRPbmuABrjw7kTfEPzD0Rpa0okrkr2AJZzthIpjSSyGW72eVj4ojy6xY7mKgSRe
yLassoFtoKkhSNfokrQEBZPgpjocuehQKMTKm9Xe/iAEkgNoy/z2uuLvXIC8Gv/I
ogK89d07Vv9RL3zW2E2BSGO9w0WkD/BCTzr5uLobGh4lmjDqUcoZ1MZVyL7OsWzd
wIZlAWTreHyLLfnHnHvhAwTM6pNARRAHmpOhvhGT9mMYFTgyGnB0yG+WGaks0MhV
eJXtxYE2p34LSxflLTOc3/pOcTdUTNN/RoRGlyjXJz79E0/RaWdF+Td8JUPlwfm4
8570HbcxHBBqNRo/VE1LQ2zpVIuXl60g0mHTk79QLPXPP0fJ1h9cwraHejHhnNhZ
6ovyiXN1uqdUS2KpyuG6ifEI+hvih8bwYFX9+gwGH+3xHdobaAs8sbNo/6KF+/YT
ylu5jydOjTgMziuw8jFNazJEm2NfK9qgc8wdzxzmF7c3Woh3xp2ixSb8ogRqTpwk
y5wt8LIOxZdZiZvIYBPUVDd7gxYP4S9mXWEZTmzJNR+i8dYpTYdfUbXqekXNcQ60
NylYtCWu1OcTS29/bdhOpE5dTnRIqzqeWazJ+2Lr3//f+gumQEUZNJKyjx1Nr6Z4
br9f+WXB+9+10m/pskXZLGOU51fENOcc20+ZdbovNzaWUucrGdrfsnn+/Ts9rbI2
5GT62J5fL7YmvdbyVuup+0y25q58xxckVH9coqo6GXKJsDvbQdYAfXUzZkrlftH2
v4tOJgYqPQwkQJxV11Eqljp12fCQZCLeEDRvJpa6/O197svEpafqPgOQv9+AfaSy
vfcCZWNC1bhRhzgOtD0Ba/8euZMm3xaBzgJa+ri2vmjBZsg0rRHu6m/KJKCY5Dal
MUTO5eXAkd3BoP/xhr94nmgGQoqLCXfAsF5n1OcUszP4FCWyrrc4d8mqs0jXsK12
oUItUEo3A8vM94K4A3VG3u/5Jqg8lgvTIIjKOamjQt7VDvsdqP/E8QTN+K24VEei
ictP3Lto67HPX2mJzJqFRXjpB89RfmHFurdL8bkl0fGn4RxprA5rK9OPwpTmp4m8
1LvjQ6+N2DCQtYXsh0a3NhcfJyGflZnqWOM+2u0jsxZDePYEI+dNzQu8/mjpaZer
+WAKii9CEvYNS0QwwPKDv26mrXBWI6N3c/wzmtoQEvIHB/rLNn0zDcrEuSJYjkWn
ZBbWpDQaN7q4Vtuvdd7zROOaBw1VeuPZzt3YaNSVe5XdEcnSlu4/d1i/iPCD2SHI
tJdWyur22BfgQMQ+pzM01CkcGyftQAYpOtpNFWb1b1xIi+VWi+BtSe1lC4vK5xH7
VJati9tgTs/w/9942cTJT6F4sq7n5UafzEBUdBOVO5tNoYOcxIy+CK3SDr4ane05
zz3rHzzxjVp1Hj/kX5c65Q+rKQp2kWM7q/HXjYbX+CC8AtJseAbf7e/8uRyGIrcW
9UIpx9c374DZ6arFhVZ44tcRDQEymWX1RGVAA020R1rCedbI3N8YU7xlr7wm2n19
LK2aeEbCpZBxiy1KarbOXyYwlF0OR6tX8MbwEkhC4HAn7nd1C96ouTOSHvdLwEJY
0ToZCZaQLybG4x/IU1YAyg9DXRinmjzUIAZ3FTlhWHDlxkgKOj4eDESk+3LV7jbM
LfVGCpo3Ot2nNb8/mo7Imfk2RfnWI2Jp04duvKoLFRWQXLIcqpjFbZptTAf2Fjcq
q+87G6eho7TIMdeCGpBkmqPGjsbiVEvabFOb6zIaFZHJZOuhq0jvtUDXw93yOZl5
v+gN/mstGEf+gBDYH3/JuveYMUvn8Pro2mAYrzQSv//zFL9+W9qTjBO33xq/ltv8
D2nGgh5brUZdCaX3e6tmXsdIKHgXlxQmkp6BYrZRrqS42QW9gXuj9LsOV1SwnHsK
hwQLcpF2olK+Lpp3mZ8UiSgEyj+S6Z6Sk5R6xvL4ELYUk7qmOlHBS1aN6ilNO8cg
sl8l8Tfw+s4jt5q2TxlCy9quUgYe8dzmiYgPLYqVy3OUmfNp88F6AmmL3mZO8n6A
Cws+zsl9ylQ0Xm1BDMxO+WWYqcup7+NfSPSH+ui3uMc4VcAYn43NTqLmH8KxbxkO
QcuRvt1kV+gODtxvnsL4ZjDbKECi959S7m0wic+dMFsakCpUEkd3kvKoG+ICmvSk
ytCrAiSVlViGnBbNnfPDMqX2mPGWGr92l8+OiRjd/jTNUc7BVDCB24vkA5W7Sui5
PUGnSj3rjByRhaillRlwIrAhsGNI90CP4XlnBshjvIvDE0/CS8KXfkUP4OexSYKA
mIUt3AWQUeX7/2kJBv2yOt9mtfeaceIw0cx6dDvOcIRi4eiSt0JC6WEV8qxkFReV
w9WmsEP7aT4CrmKiDjEt7RDtf49sTZHPSVx3yBYddpf8oy1jDjHKAxGl3rx5Zalh
OthZ5T0iw4P6yxUO7CnkRk9CbMqq1tlf7uLVrZSD6d2LRoSN8dYt6Q5fCJb92+Wz
TSlWC99AaRvYWm2Lh215MPcMfgk8axQrbCGWm7owFnRRMn4Agegs92sb3WHmbrNK
WokrJwH5ON0K045KVdH9K+3GmjU9rSnfcZR00ww9k3uIIHOU+kQuBI8ULTA+kSII
h4xroOApZlLFjwQ0iDF52cBTguavxupTZmtHYXq+5fQUYdUC5CDJx9qNG6id5UTO
0+AkuLKhvB9w2XTWtNo2qpR6+V43F18aVkqg/P0+1e1cXFBwGT2p0vNdQwjBB87I
M4RgxnLbheO/6FE9/tjYpozm8dm3gFfSKRVvKxYWhUNVmkN7Tx2U6JX5FwhZ2vs7
28sYU5r6HWi/6SiqqqMDJbbAegRPkcab9KgvYklkrezdLppsJm/MRxNoKp9YCm8u
I1s32cj6uA4B37O4nbBN0SntmSA9tKo4g238ZrOF2HGUN5WXLdN1+LwM6VPK0YAe
iUZXFikto8tBKtKhvgNrW/Uk3bVYN8j8WpRFSlJLAdWp+dcMxHq3TtBWNLutaBrK
Pr761eodph6ELoHN4lpBVHuCHlNuqPfx2VM37wILtbHNqRyMNcD6tCeAALhavTWH
nTDcFB37g+tWuDlaPVBObIT6uBrm7WDH+82nTAeG8B2184L0RJOQxU/FYPx0plgJ
1cI6285JYqIS/56mjIa2RtZUo3x1/YgbUVWdhGfCsmMFElkBYx3Kh/uMpMQVBgzq
hF1soyJr53aglN0cki0JHF40K9U41s5P7c9+LT8jxBh3xKQjppB2PmBOVP+Fs5r3
YtNHAh4UKQEkjigQRBvwSHUzUpuNJgBU2YEFgGY5mXahualQqlaLs6wKUo01WiOS
DrFb32r86NqfiD/fL9QxtDNafIz0UdEyFlfgGTOuBPBAmyH+/5pRAnA7hIOQ94hO
cyVWEVSocxffCvQgjqiSfio6orKhuul6bSDH7Pk199ldsrc1o6jwOqDKRbqjZ5OL
H2hrwI/6CToX/l2nnmRVg4hOEo1Gv5tgZN7U89e0CuzhUuV+OuGmaHXSkhBVOafd
PDPt3Eh7UhxX52Tj5GZw0hsrArnhb9iaokX4K3gZs9eUsy5uEMY1TmmW4ZVeaRz3
1sZMdQEVmONyfGIi7qWyuTKGC46mjQMVOaIayw+FCGFtbBctZe1i/lqbPbPoDVR8
cH8tt4+Bj9BgSSHDGoLT1SNf9PJeMVrmMQxD5AbhElmh1cK+ZAjcf86cSMkeXUJ9
yF0/1tV6hD+Q+qxFArfB3c5uGVMOVB5ps8t3HezqToQrKx4ydmXt7NRksED6pTEa
RsNUluzv9MzhxC1foTCX8VgB5asM1Y2EmsdJlqiUiTYmDT2D2OMR5hNa1/DjFClv
xJWIBD6neicka7uV0X+pQUqZ9K+X2ONaXVuLw32U7IgxsvOUqSoRx8mWmvdfXvVV
E/tFO/xOt6s9mne3LfQYdOJxRbr8J9FurMKTRXqT89hNfkONiEaw6o06KnW81AZd
+YvhfIJbJl7IHvijobYozzUcQ91t/s05318KBBb3fFCWbNRXaC37ts4SMbNRbn6W
lo85zE3vHc1CL4xThSgVbjmJ1H6qMp+j3tTxhkg6tYEBh7ViFCOw+QyoOcLz9Ww1
sZ8UTbb8Nk5HqxiMFAkb2XZYI/yEJJUu51v5/M9mYwG0G3PEzkjm53lQYHwidAYO
hZGmdqhY06nwPs/YN7QUzo3mDX5ELKN/JLGNKGb7/fWZEcYPOtHC9TGZwajE4MNB
v2ba0ey8etdA5To233VS1dIvJpCcB/k7CepoLsg2dKpbkuirPYHt9djserfsc6qW
ca69pcjE7eL1kTyY2wFLQf/nouRZe8NI1kN/Yr5fybf89lUMaFa0ZtrXZnzlwMtT
qdc+Io1wZV2MyYPHd0c5i7/APhed1yf+V7jJ4qLxzeA9dWLadSETEUUMs7k6glib
3IQAf9WFLItOsEGeNb+/MmUIZEYbBeMLFyCKiHauyviHEeLvjmA6l3FZFay/UMBc
Cty1O2/FQW8Oep6mCiBrC0lYS1xE/8mu+DSafHMtRyq/TBFyTCDXuAU47OCSqela
+GvsJu0L6fwXghRSQlevcvOwTkwqbJOXlIrWgXC7J0ZMeFjBWR4mLGMQ367iehmQ
PLBnu/luE6nORD2rGKwsXFGFmNfiBjYDST115s/nCum3LX33O2CbNUoqf/TGcTk8
9AAxh519yVN2UEkPw2JJT7dqxyTZpM6YP8s3s4cHdh4w5C6La2CwurXEh7H6WKSe
o873nzHl3WNb+MRVA7fQJD8Ak9fN+L0RIQpDJ1iGvpqghyFBjsCU5VZPlVcOEuII
f83clFohEa+WFyVrbUIAUwQawsVhobV+W7mKz9t6Ef8IwSmzQ2X25+8he/zGtnd7
qHZwbsvvAuMshC0onLPMyPv6TTtdefFhK19gEyOG9FsD9nOyklCFnLUwwXqjIIlQ
t8QHELTwn5SxiEuAHNfxSYVpmZqD/xLtZMq2YTZNpbLk+acsp+gfb+LQf9p429Iq
tLoeD/EqXoXfMbnxzvAFHBSIs6cxM3U8bH6y5I50OdeiXrxYlaL5/DGsE8+feh9B
dhAenx14F2uerhV0MQqstSFNjyLG63O2JmaHUn20RB2iXGgRX+GczHJQwFvJRvDN
p5AT5jWAu6d3INqc2NKlsR/YGGstsFS6Mvwh6RhqkeK2H/1fcpOkw28BrZ632D9o
MPiKAYCU/a6CYAdVgndyQ8y9ms3z43EuH449RT1nUvsxLp+IR5XdJQvPhJdm1FUv
7OaZgiIGtGLs4vAi4F5dtoQu/VEMhOHxLCHGb81AVOxJJAnFOaFM+7cFcmtlr8qw
yhMRXz+2HdjI3zxLmRqjmhh6zIjr/CEL3saPjHj7iRBpHovtRLJFa7p2wHobkXBp
n1twU4/mTUyCiPz6VMlC0ObNqn2sxi/H+Uu4mrNLC7asi1h4OHMO37x26IAZGYzS
D5HjwQHIWeLv/n728L1rucS2LRAJWi69MglcJCJIjs8eAWoeXofsdOrvpoRBSclv
seY7HbMaSLiGDDHYffLlUL6GRH5lNROLF/nEVwTv2AlLiiYmLIzKNgzvBAjB3W5I
5jN67V1EN+7PXRuWDe/UwOR9tNBbdT9TYNgXmrzNz4sJtxZLBQ90t3wQ29dXtkcP
N49JmjFgi1AhXprkNsRzwShbEg+GCJfjYe4Ay7IBUbNvQr9AzyJhBsKdzjsxWSOg
8oudkXc66RfNdMckcUMrt9w/GT4dghCJcvTlAk6E61rgmXsORpQ2ZjcQ4epVUWa6
h+WhjbNbAKKUIBVFoWcWWuK++vEUIHlvvr66HSBGF9NU5f6apsSGAbql0fwyApeI
2QpaCzu3U9GHSKaTVY4XwQMAUOtaFHqgO2NKOy+MvW6wNOxUvHeUbfvdznmS16wP
FhSH+os15t9imb7dSPfo5OUDzmJR6MIhTBTivwlBw+YHE6zrBhpKJZsVXY+5rGf3
gFQ1h4X0o0xWSS8hYK3Zzts9K5GKKdkG3MQ6iNVPVULH04itUE5eUYNp9XNK1yNQ
t3njsd8IGrYFGrGy8cNoKKjpOC9nH2B/6lcQQS/8ZmingcDBFqyxnklB6NbI4Ybv
FmAFhk2aM/YPqSVGwJ5aj8seuHzUn+A4YbGq00UTibnfyvB10vsEVQDDQ0kSnUE5
oQcJnLT8tuVaqanI/1I/rC8PobZeP9xVtlPLRnze0nKOyidUNBL5unPJmeVi3jbg
NSiTKLlPUqpkUEW812ACY2vV0zx/V3o4CMm0Dkaj/ie0vjBG2XvuabvbuXYzOn91
k+lkmh2HwcBbaelZaarqsrm1lANj1QsC0/KIWV7jHXQ/bDhMb2aiHHs8Kf1pl2cw
zRjjdw+OROWM/viQaIpogSReqpVPoEph3DQ8Jge/N2AOWb6j79W47zOAmDRjc3ZM
AdSYipXgbD+EzyR5pg/MiIrAv5H6EZhh/BmpudZdJ4TrWP05e5YA5WTbhrB/uFFc
HfO9AcCdWR3UvpRgKHR3rh1GdUCCpM2QD6lJwMy676JzCkpU5PrgqJTzvk+7w65n
+qXsf661y3dj2RpZ++YCXZLe5T4NqHrBb9efupsh3mlPUDkKA/JNbG8Dvn+DmukD
GvEUDujx/QfUHqo0ifEMtSn28F0VyglAJ+2MGjVPCttWCi0HzpF7JZREIas110tx
kOj8iQbJpBPlAAy+XuVPgRaTavdlmC0vbpA+w3yrCAx8VcoVbVWoeCIKXXhQP45s
ignJNRd9YxV9b3s6IPT7JBDmeV4Xc8NnYdqIy5l+0b9gLpsRU3v154+ygeW1CuGI
f5W6HAeyksid1Vdbx4EGc0WGEYmliymB6BJgT7Oug/bngMN64MUtkXNZImpnW/ci
SNw+Mu7ksNRAuyp5OkASeLv385wG5CASlM01V8zd7tCvsnPah42S8XgEak++pZFr
0Su9CFE4SF1wZy86/wurZPY3P3Lai1mDHJBJJIgWOarB1+q4ukdu4dHbYAA98z43
InJC42eNHErvI/uAM6VX1Wz3JQl75is0EPMuAhTzWqU9U3T53DZZ5sKBqGpVOC5B
inqiKmFUCTsxwpmuUSTTHHJuZt2H5zG/C0LtHZTWE9QFWtFKQOQhD7l0jtNXdXZ8
ZN9vZM8YxWSwcFcX7QbsYomPYpQk5r7Bc8KSlDzMmJXRr9/HXo91lw8bvhMRsHAh
JA/kRtViyRn2zMTzzPrA/T6UJ8RKv6KOi9SYQ1eY0kGpDBcUBsKniBq4cGd8gjzi
0KPn3UCmiNrXNomposrgjtawtOz82dssxtq6jAQJ54qLeOBWGVaP7SmT1reILoJR
OSridK6f+nuQZoeq1tXy7/WBz3BnDnLRcEdb6/0oUvbqA5edtLdr+INlLGVojm/I
2mMUtNdxEMRWvP26TTjuzZ9Ige+dBOL83b7m2GGRY6mkm+R1HNIbn/h9LEwy1Cue
uXAu0UAqdITZjt2T4lWLmqgo+/MSR9/Hsc3RFZ+W7iCTxHOwVXjCj3yZpUQYRbrh
aE0iKdPJ376uJfheZjbR5VwexG5v6cKyOAHxRlfF3A69WOXn1ntib5h66JsfJ5P/
Z5YAivthp17C+qH94pG7CUQvgXX9FXJply0KKkfh86VD/GVjqB+UXdD72US7SO/H
544dOzM/GYUyCR87AMQNp93YXMqsZEb3zXpLQF/iCt8DPVHaqAwDy0g+W3UJEzZ7
iukJ0/Gt2DyMJoRsfIlI7iqNHeR7/Tuh1XPYq7azJbAxOl8ggCGiOPTQBaDTusj3
Fp8WOH/0HocVrpbSFxICyU3H3IHZyKXC99LPsIwLj8EqTSmF+pLrUrjTnrYpf5Rc
kNHYK+Y/YXxFZcdSuvm0Cuk1v6P2Av02Lkm3UMWZJ8DsFIbCx4Nc9aPQ96Qs2pcy
DOXi3BSmIVw87Dn+fFUnXMEl63F1MjgJ2ZdzU7J2AaMnz5P48bA7hRRJhg9X7hAo
LoLOCPW0m2TrC4yZ0C+hH3fze0uWy0Qs5arULuBpkuOBHGym4SeWg9Fa/2Pv9K8r
R7sxvcNOycdPhn+7C1SRJtC3lZc6z2n/y9FUhxJviAzjo9t/5/2byLwMO3l1P0te
BYZh4C1H8fzOjJucFIn1zGIRdUSYU9c3xJpnokHPQ68JP4GNH4w2mkjmeukGrMXv
sqzQi5YkKExtTWriFk4MGNfagxmZdyNUkU4zIuzAf59/Z1DQDvCBXXV5w3F/uXEw
5R9sl+BCTlf1CRwXokG0D6XBjKCvMzaOYIwPRbhp9GqNgqVVERQddsYWjRV5336w
zvBq4Yz8g1diPRMS2qTwBsgQ4V6bwjujTpqjZoxH6yuweW0dXc/YsimKlOIwaNO8
k8fEariPLFIt/y9J+zvQGcKmrmh2jfAu8n0S9dHM8DWZrI/ZASsfDLadelLFdrCi
DZFCfIwnbnQWBk8F839n3faYkDbsMbRKUiG70AO20FIGP2+DnJZQxqBmbPukKb3J
bjN7S+JegNnUTNxQx/YkgXmHaiQKzRe5c6pM1InrWBJqE37PEbrKUwk6oWVXL3uV
CD2y4hUfKx0uiygMKAtfme1HRFJ+c4DnnAL0yWfRo10MYFcZUcjbG51HuP/2L5ks
DIMFvI/OnaoHYFJkX5lIThVZ8lwfYVjJic0kAhh/emZZBiwnsfG3+pzFRUl0N4Ym
ADiB5bvED0y49S8Ty618Y5bpXONy3MLkX0ZyFy2jssPVfZReRLz9Eh4YZs6FSSBD
n8ijsltrZ0Qfg/X50Udq1OVHuVr6tfibXAsSV/rTwryZ2W5n6n6O6lOA9wfO/ilV
VMBS1ZGWdaMvH/Z//edbUUeANhaOGIwx08hH7pxiPNpx6K6M0X2mSLIwyK1pmlaE
mf0a3+udN96xo4I3oVX3gGuxx+W4o5CjPBlCkJxzQHvC5BE/wlcrBzgQ32KDh4E/
LpbWNjQ7eAJZdXSAawGWpNAeDD4V94MGaZUT1tkDFfRNpmEpm7KrQHek5RMx48YO
jIEw3RoxdEykt2GYONUB6wnr2iMST1R/HK2MPiA3OLsTBOPW6eY9NP0vHDiB5R3K
qA0OVjqpuXmZHJNlFTzqAOGd5VegSK/4FSw/sJeoXWp3+po8vRHnDnMD++RujX4G
R76FhbehyAxyzsaRI8TfN1edRaAKWjumIpBTPO8UEq9rzcHMqqg2IbpThW5Dd/ij
96ANdPPhnB1EaWYbqmpUA/F+FudaarariU2vEiN60SfLrMGx7ANEf+ST2aWwCCI5
r5r0tFMyyjWajYph6t73NJx0Yu2Caqixvnno51ZMfuxayRn/3HXas3sESVMn8279
jFZCC860U+OiZeVghPLXhrOjEdEcaLC2Tg0ZwDC7J4HMtAVXXgMrshlaVFeVPeFy
3ja1QblTYgTkUIYJy0kVVSWJ8Y/pz2QHhdaBzN+AH5GzGT05xEOQLEmrcofRyvcL
5JJVOY27P8LVBL9a++8KxdLZ7GSTujGJS/C2EFi3JKNiwv6qTLeX4M37CW79Uw+9
VXIq4DhVXH+Sesxbm5ka9lADaJ/tPJwhkOIM7HBS4jKJZFng4BIVwQBy6DQaW3Pl
jXmrC8Iqr70ieqm3lNL/SUsw3h0ibRM1kQ5BJdSAJFjjTGhVJBJfPH8Doiv7ojdD
nH8SbP2MEjRcZHFGiSx+GFU3jKgCMikT7Y7lp55bVscVWQU3TYFH42+2qqfJ5oDL
RgkF7Vn0LKTiwCg/csR2TwKH6D7+mtBrKWdbeG5UDiKqp+cV37u12x4CeMf5izn4
D57Kb5Kr1SEQ8Gdx3ppGmVAsHugB1wH8YOIIAITL1i16WZ6umoQ7rIhVFk4hMu1c
u6VlLzOq3AAmLCAfFAqnRAp6j3Shx+AJ9yXAQQzKQApx7XxiXI7TfqEIcq6UDw0M
8rdfflKEZXqhS7sxQzRFNi+XGQaf5ETzErMUwGwiOoMm/nBsC/n4Kfaer7kD5gno
XSA4wAgkIljIRDVtv4nM2VOiH6klUipLJX6lgrAjmA6cH+cTbohCQoqX/ikkUBP6
Pi9LOkcmYqmmI3tkC8TzlrhEnM6EZAB8L567x9mklLJP4jwk+SOT7X3KRW6r90e8
Qzg7MXRR+Snex3nxzH6luNyNM0Q/0DNj5YyuRJZfUPL/9QWx/W6wSq/DS0lNYNTC
ANRLTSaO6byUzUxYEzP+2VDm5p2BW+Bk1odE1p1H/ZMpYvjDz4TnsG9WsoloPvbM
3XGclixC3hktO/N6DmM4wmCK+dnOq9mlRyFvWJellap3dS1bqcWfVH7JTsp7aUSQ
ZoNxWTR7uwVXRDmmmbQ/gMrzYhf0O5GMbwi0JsWt7NBxz4WNN+ljQS/a94qQyfTO
4/fH400U6642CQ33mKPYl/g+U8zzfEIss6D7OuG9eQhXNhSzLLL55xT0KgkzsGk1
UvM9wll85twGjdFAy2dUj+zH8h/ZEWIBcJlwW8s+A/KM8n1hxlVWNwRAn+eU++Xk
x0wWdaeJ4BS1Z5H2TMIOSfnDeBn0O5HsOcJqbMpnC9IhesKGBZ0E2HuXrzC4Z87p
eL7iQoVReoHTEJaGbd+pX41sQJExlAtPl6T4Sw29sTeVHaBBNekiOBJjgZ6UdID6
hvQh5y9XKJ98voKfOHSsk768/xNme6zX2UrcdkZzAeTLRazXxbqcVgaid6TEe1CL
M84lbh4JAaAUCtZlNo050am7DrOmoWk26G5qECWrCgZtyq3dQw3jVyXhDkQv9fiF
pYfYDbVr6h3DselNl+5VuhdAuuI1IVU1kPneZ8fA1D8uFVC/RAmczKHESVThvr1d
i9jWXONlnlthz1CINS2ZsqSMjinGp6wnn+HIjCjPnl+JMO6fSIMkMYaGJ+Wco64X
vliRoYZy28zcUK1wfi2ojkE7HDl+uHC6dsgfM8bnVUYkzzO8y386r9IBdO5gOy7/
xdfLo8/KqkK17lVrdexRe3UkGk+UgyfQC5ohpRYd1Pvz4F/5ORrVr6ir5cT0O2mi
EzMOWpybQXGjDcd67i5ZTAPQC9sW3PuQ1XAm0P+U0Er06FVYWTncPm83jBv05IWX
aasV7yQAhqZVZv8C+ofp207CDutZPiSPiwgOdUgzK5g9jU1Hx4dY+rg9CERPIri9
vBJkfgOueJWTg+ktXEDyxrGO0gRs00Lk2l/b4hRu+1iN87DDsWwAHqofZ5gV18kv
seMlhE66Okvm7aH0BSBQGTv0KVZKNltdpEqbhNiqqZbbKdC00UOofjzBTR5Yue4L
NWARoX1vLFPjFXCq3AuEvFNQB9z4h51F0W+papCLaQq6HNZgbWIn4PQLBse+IHoe
ex+nPa1VXK3ApGTDxY3ibgaRQCIbYFsMFrpPdLLesU5vKmXWTuoBH/NGCcinCJ5a
tNcY4dWDXL+tCVyYOXIw4Gw3XzYip6sC15PdiVRPEQXfBY9fH22EUwlsGRJK178b
AUmLvHz9x4slHuTP641odBYwlzhhdyZU4CGQ66zYiar4Z5x2nkQBKBULIxYskvSg
b+SJqHIEvC5YhN0ACn1qZ+OeZWL5U/7joAuDs8JpN2UBqYi0wTGn+rTE/MLQf4mF
Ub1zpquQoVNW+V2LRllKbYQWoL5Su9G39AkMhdXS0+MAyFf21Tnq6LvSDpp4GMsB
Gnrx45Ay+OfbWNv75k+psIFPtKLCyh3M7MayjRj/jMFi2O/yeSVf5Z/KkUcxoUem
RQUGlU/+/7CIYJU1kUxtBRnM0Phk3TnIbFOyTk3XRyHluQOuitCrgi/TvyazwwnG
1nTmXVJiawAVPNdQRXOAIp9+ESNGXQ7go3QrM6sKaP4jwsO2Jpfpkv6tjDgNOQH9
aHi4Dyyftwz2543z9EyLNaLI6Btb2l5ZWz+irKgft4673BLaQmPM+DMO3jhlLbqw
fILPwym9HAoYExfX/Vt2Vii2odwW8lKZ54AVdzVxtTYcyTp6hg2rKemeZgwy/IQg
5Ko9CoIEN+b5kRaA2ZNTdCKhqNQJRtx81CbYupytaNj/6FmStlek2lhKCPUOUVG6
qvTPRRwSP2vFNnkBbeLahJWX4n4Ajcc12uxf9mkO5b4N/8+d22CjwCl8kNd6aeqn
1cJZs6wevOj+cQnKll7AOR8q5OxIJx/u4gAmxFE4SXRXWhVCg1oLe7SQMW9WiGq1
1YmPI4OvVQs58PxuhpdQBNjnPerK1fLFYpqSs93w/WGKXtT3K//qQNL9TjSDZSC5
rH4p/A6ELFnieW5N1bLE/VO+Mo83hKyFUJLkiQfIc8jdvBTsajoKC2FCfoV0Ev7h
flAHYfBfOrR9pSffjckY3OxlpiR5gQ4f5AyuHNj7lWbtle9MO2sT/M0lNii/yZgd
UI+s/nZAPWegNF9/49ybec0dBkP4skulh/+xQ1LpTF1ym7W/NncrdvDhA0vgJu41
WeX/+G4qeoZZC6jl4DKGvM1CKe/H/U5eqVSbe2GucuIP9gQBZ9aXgrhZKAGhGN3G
YIGoAGPSeYmDvVvqitmFtI53Q+teCDy/HElXs6jhvVy/ql37DSWKjF5M6l2BYkIb
ooH4KEq7gXTciyHR1FlTAcV4TCwMLjCsKbQziDzsFr90BDmsMSPdcXDXvpJVtf8o
4NJqo6w9USuv9jfUMGqIcu6topiTZjgHgDv1lWQhogxepN8s3nCkgzMx+9kNI2x6
b5kK11RVYlOFy77HuFboYH90HCXZW7G9FweR5nFArJh7MXbe2bAshYVgUbNzGjNl
CcZgF5XaU9M6cjBBnoq1LaaAuzNfDbVPB+2aKdPOPyHqJxykk2eLQck7HxD4Z1Hi
eQef42L5mWJ8+cfc8CmYLjgM1xLDXMvHzwQDuyG8idO8tOq7Byq9ibNqdzvU8ZZ+
V0khz2g2WsWORBHoNZVYQDzqYTR3+MkhL5HR4aUN1l9FYqia8rTvJN8vwPNrIpWX
Fct6dnLhhbRcPDLvjJEf6JrcThI+vGFtZR4HGKI6uv/nltRFQXCLebZmRyheuMLj
YXG8lxXbPpfypXh82S1aEodObSRBcP+sb/JclrdTOxZk0ztI31o/8JFi2gZYgYwI
1RNvk6BfH7/SBYWK8hZWb+MBrUQYKKecOisO8djrpOSnPUV7C4MZ/Iy73eNBXPJ2
4S5bLZSpBdOPG3v/66pEpTzIkUDzgXAs9N1iIi+wyejfIbg/ZIXFmlaWjrQLmPz8
HHE2xZ5DHUI82+/TkmNmpkaZ0c7KET5kQVO7Yc2qsvIBuEACUjkagPE/de5erhIb
AEHqQ0kwvMWp3Hg37GpTH556f7/UMSzeHYIupEKEC95raHd1E182XidU6eF9eiTG
n7PvTto0zZcENdiLoV6gb+gXCglkk21WaiCj5gNUsl1k6qtmfCQM6mZGYoYJK3Lj
0M1waB/PBXfRZEH3oNfCSp90T0RnjiqkEoYrf0A9LRJKMuV3d1d47GHLyFckh3MK
evL+befbG19Cuol+iGxjC75q6S1Mm/f3zIIlZcPYwA1F1oWRc8yEx/m4mUA6IA/8
gsCi6T0oCj25ccJSBRT82XPoxi2kX1RGrYmadGOXqAN/c5SSn0EFuSO8NClZUmXv
RCMpn8dO2JDRInPasTxKK0KFGUQCDrzjM4RllJKE2CYLZLw73dttUlMBeg0iLfJP
UQSd4uR/TVFUSPswpzLmlBqPLR8il/qwhqCFqJKTMl51WCDl0+VljpKQfjub6++k
gQW6LaHTpYgfnK+Qvzk7rX6hyfQFfSvJvC/hDN0RP0WHiwOhRbNbC20QadJEM2fC
weWeT0Xtv9TwINnVLwGm9UKGR3H+ov+EX92K4K6Xxi5DSwNU+spjamkbJpjooHbj
Xx1X1Px6ydW2KhDwguwCFuIFrk1gNh8wN+mF8B4AYoWWYdbrDdmZzi+jcHRf2uOz
9qN0Et/hxX/d1xagtXyBgKBM0vsTDHEEPXmX/YuOK8an+dxjxashG02mt09YzcBM
+FEPfbC9u8xm3CfObnyPRSNmbK9zWxSnwHkgId9Y96Ui1uRwLHbXOA1PCVyIMvRf
P38gbPR7vCaRffHVAk1FPuRV9a6JA25CUN4BYhYND8k9sQPLZjhuRW8qzeKGdJKv
Xw0bjvG27bJ2eFe5Zq3hgPstYI0YNf2RKp49v0JM8JAU/fMGxI31kYTbISwHEj/R
IUUxuxGBkuFmQmuIl6/w45Ug+es7Tnj7h5DyUxMyJqE0X2Et9dyzxrWPLEgMvAbl
oc4vAzUF2JC7IpCe8glWXNIRB171Jd4VXJikaaWzX1/sKO7ejOOxp5JeivB16yZP
en0OwbqTM15z76y+NkSOJtedWF0VLIt6N/bvf6mp33F7bm1X3PQhHLBkakemdFwk
bxcGldjoRb+tKvhFCWkNPA6NoX95adLQbrCRJv+gpMQCgT61aAoZY/RHbT7jBi+1
XWW2uDat/ZjOQzUKh77ilGG8kKqoXIk/8dwjZ0Qci5w5CLSynQjhRcVJAf690sfl
O2kZk4Z8keUb2WX2L40LMarCpIrtWJBJt7q3B0LZzI0hf+whZ2mkPZsyvfunIWZJ
HVkULJmmycYkOn0zsELOJwq+mmtovNuyvRR+xgh8oTp8KtNg89sBX9CBmVMjZBfO
F4PloGiXo2sEA/tdpt0K8jyIIdtfhNNfYuZ8L/OZUnsK3Pr3QZW1ZFHntNJskiS9
UcymL6jlxGDasQbGkWSpse1/OIGAr6SB2RVXOODLnQLsazeDgCF3kmCw5yKfDyGO
77l/oENuNsrGP7lAWWuA/oRS2c1TM77v5PySEgCJVPJ+y2sNCswR99nQMT/Di4t3
Lb36GMHn5fNf+ccpO1WFKgGVI5RRNa1bxhnhMmhKEFG48HEQKFQBZFN4rUyKVF54
slDZ1c0eOkPE4PA5V06R8nD9z8iPKCqEasl4OCrF5OTK4lc8olb2ycO6wclajZFA
4pOqbfyD/1DujTtTqgVBMq0Y3qlg354QXKzPPSf4quXUyF0iMtSNvkjv+3HPMMsk
INhN0N0JDMQF0wJh429/lQAbsT+HLzcjSqaLWOg1Ib62k8fApHKzxFkUkKIBODku
YiAmYiFvWjGLc2B7qxd/FzJs8EL6DqFgWpBWHv1F6NI1XSISH8mMXaG89R11d/S/
sYB7GxVEcgip1iyBbtRLT7aF9bLP/cUQ3sUprj0BcYs21vbjUOz2eQFlDlcx3ZlU
BzERTNml60pbZzibk/ZSjGWiRrSKw37EULHWTFkFyNcHZQJwAMp9csm/VaxSCyw6
38nuMrghDEW3VYky4xhRzQJ9Jn+cZKHWXPDePyzFmfJAiIxGEMXhSzvWxnCSg7TN
iZ4k8y0gLiC1ZvvCVqjFfSy7Alq9wi9eongi34aLDeeKldG6R+Mhauyvw4XHnl5g
A7PhBdloiR9jXmxcEueljmgXdk2FMJw9nr9hoeawhkQwnuWMXHDPAzwkmLKSinBB
HYkFIZs3Dde6qmejhxQrJQi+ooi4+uSn+beKAuiLiY58qqmr1fBuXbZ3M/ywWoH7
JjkN7Nr97Fi/7njnCSm4jojQGM4M4+NizDq0xY7DYoYmlZBpA/PP8AwJREaauafA
BJzeUJAcLxFRlrDkSKjsh/lDEsecSLv11Vcon44HwjfvQpChuAGcwY/4t3BLO0he
qWluu/bPHIfg9OBKaI5Y2vCiOQsIG/3fHqBtjo9t3EGmnudnrd0Te6suszfvGIud
rEoKeZuJm9FuiFdV2LBj+x23lWYTxZuzKts4iqst/wUXawc7Qi5N6nUux/EgM+ry
9zWRv2rgJKzArabzItbug7CLtxSFkYY/c1TQsDbiofavhe89aRb8DpmjpR8qeo7s
ydql8eqkvwnLv2zfz1MUWgJkp/7rAN5ZBv7m23PlZ648NipiaPal6B77kB7l138R
jqtJBjTIPSJCPTtnHtGB17rF/IFi0N+lBaNDpl+5rgAQV+a4BpWbEar1t2cKSBu3
l6ZR7nVUvVwU84CtHmxqeK89LcxBRlRhmzL4WE3uWTWFL0tnJyuu8AHkMWl9fpra
QNPeAcGDvFoHN16fVld+ifM/DrZSVfrFUl8PEfT03ki992XQ0vRuzdJdFzC8GMU1
SwZV9AwqkWsns+AqYOeTVUKp+N9gAuWVqih5gNvTvJWWenEWKJDuNY+nEWQQomDu
2nO15rlJyJdj7IJxOwCO2Q5uOt+T7wYxRb4MSnkVAF5279vbz+f4gJ3gIdvrA1tY
woOwgJtPzfwu2lhgCRnEOZa3k6LiFBodOOfhNEdco3OxGOsJ8JiRkRwS1BL3f6rJ
USTbo+7LMzx+wyPaUTSEsapl4waR4HDpC6oqs+y3rsD6iX9sG8QGw6BLdJPkYvx/
P5pwK1OUoYrKltI67E/o7YVZJPmECemPPnWLUZwD1MaQH4V07BH0a6IaqeinAs9+
L4eUKhBMQ3oTvXaP7yymrhv39gOPg1IGUtl+p7TMm2mriqtd0a0nfOLmmnQSYqZ8
D+Cv4fdcfwceTgPjP5xVGvPnLrqxGzGHN7JrROq4uRR/rbPRAx23KyesP16wlps9
5TcAtiaUJd6ViArqGx6WCVPQeDSGXRqv1aG3HR6bCHo/PGRI3IjssSeUMtTv2HP4
8PvHkjdaIHYiX5ORfFfxNxCiDHRKATyiuRAUgXxkuIZR6/FldYGx0gGWguYUu3xm
NNWdZAW3wZInGZWBZsx8Fn3V1m9QadqtwGKoZ5T/t5fKTTPYjSSNKIJ+TlsToJqN
4A/1XwrzeyECIH6XZBA3SDsbS3OWSiik+hGoyWt1evb6iws4Gy+KpipXpy5wTAJq
cWfBPzLsDlxMZYTaFtMBLyXmqG/NhsYYgw2gVhV/Wyf15mI13X4VjOuwzlGroger
BCSnuJWe6PQMdhlo16MUHSPhGyUGM60drgzc3f0OfNjdLwN/XGZn1xZtxO5Lqjc6
5ZJu1NEH+f2sqiZtot8Fv7FGvO8TmcXFkVQMLnIJAk536F8/SQ56992jlmO39UFo
ObCsCRbPZzwv8aEWSWnRt+zp3Bt7kWpwSZyVyL+6DGYqREeVsjJJhIVIvGiZAixD
hvioN3BF8gZ+C394oWZmujg3tVdXlZDLtFv7LdGuxpMXgVOtgihv6pE0DLYTui7D
ZxxYyorqCMp/Nk04/0Mt/tbCSZT0uxD4CkwEMa0eeFJZniU945kHVpg/1FyX78j6
NTXuGTbCPLwTpvvljwl7VVkslx/phdwHaK8DDenrfIEvIL62dtIX3YfvZi5iXPPx
x4qn6l3EAhs9hJZV3lj6jznpSWSGLg3RXLwldyNnrFNaQQEHLl7YZ2i4GI3TjE42
Qf/VIF8V+ZnlQBvUEYW8VYbVrupRHyEgOWyE2qfd5UYgMF+aw0WlIVRvNZTX66Fb
tZgmaxovYFHdzxydNXuEBevcuo1e2juC02ymxAaUZJCbb8eLH5EgOB3LxHzqH3Li
JZK73mMQTYuEn/hyteT+ptcG5Y8LWQtQzQ+ylKyV/w24v8xFtUqdjkQKspkbmzNs
AW+5bQMRR+7ATBuciEXoSo6DWuvRrwkd1quiOZYTUgKymW3fM494+Gfu3oT8XqAJ
Vz2M7xfr8IZY5Xrim0nniGAm6AfWBieeEntkETLcT+n54rd4xL7LZExYi2FpdeVl
Lj61DqlXdSYrbfsWnGhDDrROfD7VqaTGDXIZJ0ehv7vb+STH8Q0iEI/jQ5e/vUPt
bjkyHtLJQ6zHUmpRS9I3yB8Pqo+4N3MXT+gT7KYfxvruckl5rK/zXMuJrWEWBsVY
HzLENREtNfZwMmP70P4+sJowWCDMhVlcknqdVczPl4/sXvYJxvwQh7xthHgC+VYw
ayPRZJqKM5tZhPUXaWbu1/a8w9LEHj8dPk4BMe1mKTxQMfFY0U8Ee9+2Yo+WakL1
dtG89wzt8L6rWUt9af5KAZLg1ZiZZt4SDNZCMCTXuDsLgs2RNmKBaBnD18nbkmdV
nh6065qmia328fvDnN5Rt2c8IOVpDuQPmDdWacxIqKsgn0CnZmcER59XSFSLQDWN
lG8zoJ41YhX+QhNbngB0LzRrIuSeSFaBJVRntAp7iz82EpFylJ9GDCTti/k8NP7b
oH1skwkq8fIWeY/As84vyhBDTVCvjbHLq+duH2SopXCzxxI31nR/bME+U55kWWfR
7bvowwdQPMjor5MOG+9xlPm07vM54yrdETy9pr5UYaVZI3rUpH3hb1JCJ9K5rElN
RoHdHWOv367NxXGSFZfkcCH6NPTxhHd2+Fkt0tICyMoZNjDh9Ma24uX7EH7h4+Qn
FUC8enWWhdS2dVkhBhIlxz+K2c+ZiDZ5NpzbBlSBDjSYjoH5nzSmC9O5+NEwFgd+
siRf92e7iQXPkQSwP4uaTrtozneuzzg4rIrG+TFx2TVvM9FC30MV7dhGzCcs/Z2p
IeZBY7XJrGIqN/I6FpeIdUm6V9wNXjv8MlZnw+fvjKrrEU5IKuPFyRO+haQiXM2J
euKjxP0Jqeh31GzUc9sBRcbLt8VKHanOSHk53ioaJc3JycUHdA2J7l1pYQUd6iRj
oSQ4abZ673xiv78geU+X+1OfDyNblBjkAqqq14BHPOgoWyNq+1IgboSyZYvbxTOj
6dXzhCJjndoIj6u3+bD+dLvYgoka+EdwPejuJNjf57EsK1jhvObcyNR3/o9Yn807
UTWDScxHhg+m5PEnFILBNIcxsu/f79MTASeengNOXRIFL0pauGD36EcQlhkYRsY0
gB6YF6e5KcMxykYM7RO2iWJ6WbVn4MDYm8th2xv8ghCzEAEcDBI0ZAU+vAF99nH9
l04TknMbKbSmFc+Tsek8pY0qU1iBBQdzavC/VWcHDCrQRDr58T0cX+ZGvi+w+Lhw
byYQFVYWX+MF7DlfLuVVMWLYGM5R+eS9gPkKiVZiNrbNCM0LH/xBoQm+obW3yneI
M5e1gQT5SLvOuAmCebblVBbfQw5pCXj+u2/CuCDGA2CisGRakc80ga0EhXcs3pto
vMZQBpaSzfb7nHVMBh9SzktJjl7DCjb7szYcAGchxkTWZd3/08mRV8C1SMF/yEX6
axK+7hG1Zn8APGpMY8dVVKnBjgqtF29/W2kDEiPKxNeYZnoUMsVzdJ0c17AMgURF
2Uw+uCz3d7n2iaumKwZVgcbsKttx1CNUwWGw9Vlg4S/1toQCXAEM0uPl5ituegmu
f3X7s/jQxAebViW3bIQuI308ASy4q26hmygZGVtZ7O0JdepDXxkesX07BvBkiSN0
DzPQRkkxCU9kFaYClSEGkQpzePl1nwTnQC8AMJ0bASMEh2zZVoRyW2XtGOT5ym0x
4Xbq35xlhGDJ5oTSlPG6XHU/yU1iWlzQlwN6JrBzcs1kBhvywQD5TKhShmObKgg3
eQq1EDjVrpn2LY/iKI7ZkmmJPiSDdhAftWGNLVLvMrGhusHHUAWsdhDFXp1UwDzV
MQMWEDBHyT3x/R9sVLAT9jqfr3zOQOqdo5jdJtXpK0SpC2nDT1lKLmtbgWVw8mgb
3h3fkWY5epc89DNSpfp0yh2iE3OTUUgGluapmMfvq90hWaAyh3bPvx/I7pCRiq2d
dWbyiEItC4NxG1Km18/GEyWChla7Xjq+TYOWtqELKQuJ26NfrBg/8rQ8+A4veSRA
esGTKSEysuLQHCiXeAkNjTSXQq1BovQ2iHdEFJM3sDUNQuBO+SxD6pYXyux0Z+O+
5g0RJBkJ3+zxX/eV87+C1Dr4PKPPKDEACd56PXldRJpYFrHnFLc8qeYzMAL4Wdy7
osl56rsUeoxjleUXGt6nIuWq7HbwRstCwybDDL3cSuGVTxZn4cjs+94YkFSTGD9b
RMGtG1wQdGSJs12zcS54FbOM0OIWhzg27cdWvDzMWFLLFwp73eCHTEetGULsVK/P
W1e5h75lMIgbUxQILbWNVfCqsvQMGyAd8WbaSjyPcofRwfw/ACEoptro5DOU+ga3
6EsUKppXhb+o0+UKjNmbly35tK4ttDc9wdaUWD7dKfG5nquVh8olDAafN1t/qIpr
m+3qeCVWTwnu6rR3I+rgaUaigBbiM+tN3O3+k+YK41b4zx7PCfQQgTqhZu/MTeRq
y8XqsNhMOfpl7iyBWC7VlGrrEFb5Rdb/jJWHOFl1braXHZdK650xPnb3q+NRoFNK
7d8i88PGfh0oOnzMtiDxFqu1sBtFpMu4mNctHp75HwGWUoTAAlkxoz+5Il/My/Aw
btAuRyCHAcUJH55iamME+5+QbEsHKh+i2podPasSEsufv7wEvQuCJ2p8PW1mXX6j
mKw3qGFjU6m3obvZY0M3pXmKYKLku8Phz946BNGeXI1A6krJx2QQfLmXIIX13zw4
R8vUnfszeXnlE+JDlqNuRUt0MoCxxgIa1LH0cpwWOGmejjhuFVI/awhPvQahIS0N
7dDWIqGQT8Z/LxPWgBg7isk44RMSAGRrhHsqG0cwSEDmWYNDEs3rCS1QTejWDUsL
vOug5JaW5mty4Dd8Fsj0aJlqo+Nv3LTx3IbhuwT+UVgCIgYKSKjokMm2UkCysQ8d
uZJYcrP6pJWIWYk0lb2STB0vDmVgitj2vdt7t8ejfhBv2uCxlLf3vIEOrddN1Yxs
eDOPiVXbAYFY+6p70FiVxJciTcVMESUnTniqo6QIzZFiUKCkpmL4FDxU0n8iNBJw
hvyFMGzK8+iPUA7N3dtZITNWVN42dK2aJvo3G+hjOo5A6OFJdRyGWyAFNEcpwbM2
6KIihiafQ0S3soMelJ06SQ6cus25EH5sOig8HNPLvdsBz0d0Nzgiij+lj+sdByRg
2AnAB3hmiw7WkelDJ4cNZFoq/EvMUduLo2F8hrfxm95SnV3hffYpW/jgQGezZ9lS
An4BuHh31mbJHvOTcW5PR1ekBpXvqfWrH5RoQPVnyPkhmUtHvC/k7TsiCF1hVFxO
wrEvcLUKBuBjS9LmFSbMIqLnWZFCdBo+yJgY1hA1UHMxmDBeNWDIR/EqN8O/9dqD
XPuHD7rxgugnLsPpMTDg7OkLWr+wtOO99H0xMdic/Zu94xG0ZJubU5GDYykkQNg5
2whbVoMrxVqMg40wifvI7cNHz1fE4sRCJ+dfnYZFWPQ+YxU/2xY09zPMGj0zIrJT
YtKjwg7AbIDKR0He9yraXUi+48OzI4QfVazi1MBiZ0Mc2bjim1bckpqCw4/wWPY/
gGLTO2irGGEiXuUQuC4HGLulHPL1ZIwbKjxZsOksEkHOeOmJjtvXGrethfAxZKF4
5HrheyNBTocoeZAMFNIWYI0iZskfu7CwVwAXzP3u34XP3+BxQL1njfjYRKvw3WRr
OxfeRbsbhWN8JK8zXBKx1kPce9A2P2zsq294pN1LMdx1NdnfM00Mz4I5NYmF1uzo
eAUpaqDFNtn+EguNX9e1PEXTln4vZOan+eKmpvMD/3AjfjQ4r4DQkqBvUelP96oH
ujuaRgQZYcAI/YSTbbxCz7RjJepIIrLiWlvsLIFVdf1g29yhADf7lKxGzcID89VU
bxE+NscvXGq0OW7ewxfcNA2BlczaoqcqHcgZoqbNazPaT21C00rbmb/3ci3FBQVT
r7YbeuKQFd3CWLCyZkEZPBXAVRWvD7icEfYf7I1H9sdVXBlkhYsk8C/JjGU7vIcY
y9xEzritlqfcXKdU6OdgpUSyJBKKIzmQDkH6Dg666o7E88255ebrJMYI+oQuTlCR
mAlHMuog/MG6HX6ukHmQYQNTEdEniJIswgBlVyvBBYz2jIC2esxzHEbN8QzUK6L7
lgEvotdtcdoXdhw2/JYfJ/O3OfQdlce2sLl2VM1pDm0F0wc9gzYhEUs6hhegcxYa
NHmYJTmbahpwCUaeovAhQg/oIOmwQQ24Buaopcq/U8X2fFtGYHDPwWuQ0kotEpT7
DUzB4bYOaJx3niu9XHxI4Y6lPd4pBXOZnVYkJZb1Rtu9YICgWmtwt51pzAJ/Na1s
z5+LzhhIR4b649FO2BcpSSKF0xN4rLyJTZz+028HeHXkCoMSPiO8wA1iOttVDj/g
CS3R5yfOBRqV7QCC+OmibSDkWXnDve8N+FRgQvTg2frED7lJXmQeUlnLYbxG20yi
02eVYga0nVtylZ5XtiXg0F3L79vgTBbu5Fa2RPgPp5H6WM9f3tRVdlkyH2Ui9mSE
XCHToyQNGQkkxvhQa64/EG25JCqBrheHpsdH//n//Vod9ZrMC8WUK7vR8CdZbbB6
T++SNX8ZtCOgK/1fXpTUN2Nzxj4hK8KDL98VBsrNr7I6gr7UI6m7BgtqME3pSrNT
Ogn/sy8h3tqLRwtNmMMZqkAFFARmPw/D36fc6VAUuzmWyWs2178G3IOa1CIRkgU4
FNQtnB40VvmNguRmxZeTgj90cwH+UDtA8N9ZtATB/MZqQLcrhSbGTjiA8AxsKJBq
dcBMqOwPNlI/CaGSO9/SomhDKJ+7M3HPmlfHSM1miJOKJt67oPBzFcmVAySnDIlM
RGwT/x+YeFb5OeA9aCwlcgHr8+wA/0vg8Ut+A93cwSxmxpF+k3oBvDud1jQrnWya
zYhMGaksl+gfIqrkIPOi3z8zFX/ywCufYzFMis3Q++wIhmC7Pz6COYnKu8+RDR21
yBMbttMZ+2Bttk8JzqcjM+lB46sMAIIHGeWhkyvd5baiQBqR18h44ffzkXAiokqH
ttrttNuoWqVH+NUNdUKKwPhEttaR53fAQvaWy40a65LayO4rdMWvmgyYJ5FydBCj
/swXFXGt8DkIpUx4LD+Sj6IWIOOmfK5BxOnyd9kawxDSgN1w62TBTpEuBuOq8egy
lGtRAFIkPGvYuH94hzr9gVQauEBvDEU0wRhkaJPtCd6+4UKbEDv11XtfOKKbgCXc
ks9POyQKXvhgvqH4j8sM8asSCiSSpgrgWA05dCz0BWC5eqq8IaCcyoKiBWttzSBn
fxPRfr2HDxAJwEg282IJ0dFcgQVVqVXEtKvkQGUF1tJXrvePIY6wh+f8My/uvYkp
JOhodDhaPbTmJqxFxGvBH87DPkRwx032SJb5qUUhOZla1bRCrHzegFNrT3IOg5vh
4wyWzUG2SU2kLCO3FyWUUiz7k2ph1MrakQKq2p8QTe6Qu+UKdD3+8pmguh0NEUHs
Q52MDiOj9Zxjv92EEtdmuVxybh0zWRGdmINd34j3/bilMsZCnd+2iaBnxqHimfPr
YulUNxs42sQxT7ZeAVCLbMtNpi4M3t/KVxDaXvDpF0oUeRIVnJO2Ug154YIidedS
BIjkhtJoR2pUCQoQTBb37DpNsFtNzxgSOwSEYFMBU9cen0T6kp6STy06f5aLV7o9
N4RLLyTSDfI8+pBz6x6PLzebyzO6l4v7xz2sMiExW/E8pnmoSIjH3rRdHT4imDEy
mF1poEOYFfVW1lqPyYwug8u+xe0hbTL+wrITJ/Y94W6LwgKV4YgNF2OGi2fJpJ3N
cKOZWD72wIGenZTT0J3rIImDPlx2VckCYchGl6BsZTaxGjh/8vowa9wjpJMeRaRT
i+t1LJPMZWVccDMkML50wrU/N9+qV29FcyMMTBRrj/aM42sbmvf1HQNEORYOjdWb
OgFi0O6yjxBR146sKIf/uDH6ygw/x9sEYAh4CpGskxRMD9l196RsnclX2d45mdZa
XbZbxGq4Z1amxvqmWjTYIwoW/zb910bb3dK4HiDb5KRkdEE2Vi9cyZALDUgccGyW
5V5hTj5it8EKP4hFsckNr/9glYICMWjK6f1Ip5Roe5IEqSh+6XGvxihnTuSbVjGj
TtMJre7Ply6+Q2C/ESuu8hihkhsjIkthi0aXiNg3DE7vVMWtF7ABAbrajO0HG8fv
Wkk12IGFmjf8czQh/FUYCwzNLaTj0OgMjbr+1ra0LVTn2Q0TvSeu9x998a4hYlmK
K1ahKKhPERl/SlgEO3kOXMU24uSu0nBwM3dYMNb7PDLbwjDpr20AdCw0ldbtXolL
bdVHBIK6GMyjjyv6qH+n7Ky2OGrKG6t8qk3uV2LaCNpL4Cylb828/4sm76i0kH8p
9pFsD8snlD0oeSvnIU0XChBwzqHi5Lpcg2AFeZvRwgrUaUrHcNJidqCndNW5VhSP
AuARp2Wc1Zyj2fUndHAEnuOlEEZwoAa0ih+Cp1DdXcMNDZDk7wePZMYgahSJBQP/
enxN7EnHIzzS1rkyPu1RsDHXTpEyeKEGbvYNlIj4z48yPrcGnIOng4TbEuUEQopm
u80mhvzhpA4h3sqGeqwI9YwODRJtsSU710Kd0Q+PutOs8EOI9KqDCVEcDYVYul5e
dOJPh8e0jDJTmiD1Mf8yjYs0ptOZzDsd0Gn2C3jbTvMfb3aKoR5lIhMEFeaA1ZIl
zzDr/dLAFvbc7k3yFF3+Bj+g5f3zNgdS56xGVLCd68A4x1vel3FGDdzj2rZLlNuG
/fPl4ngk4J30GB3EhF6RS8QrUYyoOes5Tk7462NGqP1GrrTs/24eaUXa5YA4JLz9
N0jyP0VDNepkhr7rGfGfOgf8mnvqOQkjtR7TUOajzqcp5UxGB+dwF6cL0BWT+MBD
uJfhwQPHRIvOmlt3Y4j8udlxZpUG/BJLY7dFPj5nzw89PQ38/J6W0eJ5hZTrCyay
dTZxYmZLoB0ub1tvtuE3r3KaJal0ecPnjh9j41E9T9v0kn6mUcLwy6CUslHcMXFV
8I8SzP3qjATCeu1kmEc6GAQmo2QLiQTsWD+xkdwx38b3r5BZfCWXvTfZfVTff/zH
u34mc2rln+qdUoeyrayfhkT61id9xeBtRyhBk+8zQDFIQDuuBZMlWfrL6SwXV0hW
sERhyb/qHIK5ogldQMZQKj/Pbcewefpd+XskYbHHO/NY16zkdNMJklp8kZzx74If
+wkoMOTD4ldtplota2qla3ovvWQG/AIvwH6N3uQbTwAmUlVSqaF8eYl+f9nNLfNY
2VhXdNuv9ll894WSytLlXCtSCxqlvJeqcCaD/lP0kltGhtHDahGGkUhNQxmknshR
zlGJQnq+c4UqvFKYffgosS3Wi8LnYwWEJDkF09ryJuE2BWJJFygi5QTjNQhcZJ98
Rr75sZWAqmporZBmjriBs3zZOBOP1DL+TdeYSHtKGDE3ndfFGLq077y2L8wd9VDq
4zuahvRP6fy6fIUYi8wxbH2ZPsRVZcKHxAlyLmwnJW0pnueZC8JXerU3+i3ovbKs
MwaS3anc4mX+6t/2PShcnVFGxJLIpktuc5vhv2fbsWO4+OYh1WR6MtiB01d8mScS
+bSGeJ2jPrCRleBLoOKI6cSL+2M6M++tX0mEQ0+Fc6+Jx8A/l2DNC/Rn4b4W8Uj8
VcZDwaIt8/NuuNAg5+yNF89Mm5GaUhUReqsJrDxyy28qNMh1SaN/S0bhQgW12BVX
FUBuuTAZ7ZR+TyxNoEcwQhvnpBkuZHQEeb/uVEih5Y6wGUktM9tsoVxE4o7+4xSl
fceRKBxfyRhi8cWAPTaHpM/zX1XgBlH3SMo2ikfwvmCNH4QQfjVZs/mc010it3G5
glUnYo6WLmvlhXBUU5JIqsX+l/nWvh4up0CgY5jTxk+GdYe3u0QIn6hE0teKRoid
0ZQvhwfThTOE/1ZMXI8mtuAe2LOYE9gaB5MmAGfwz2/i3RTn8hREC33uNAPv6nl7
4hm6b9HV2V00K54QWHMPeU6+ddNbqoTgdy4ihZs/YwI8iEQ12qNlqxs+4uCpKLUY
4WOF+OljETrTTgbFraESBKkuui5i7SMcLiFKQTSvXDsmAZxSyiup89CJV+pMgO6H
BHsWnOCRk+2Ow+Fk3ds4ylrCQXj9YDHUEiiSyH4SkuKOeRw7H6BkurlOwx6iUu0V
sSdMgwLseEz27K2z0aeQ3hVU+5ZQ/gr7W797e7JsQMdMgBjFO88ax0B6qGjPPpiS
C8ny7/0dCS5ciHb/sqIMCuWJJBSOfTWxiqi+CjhiMmhb/BS6GfKe8fBc0R03vrcd
JW3oFQu2Evg9JQP5aoIstULMk8ai2z1KkxlFDMaea2XohfdcSI60499YqlxnKFib
6jJEaOjjoY9C0/oI1/qqmrVrK1IkWh/B5qbhq93ZW/yF5DZ6SuT0S1OoHzX5KzUk
w/tVsLVvi15C3pt9gaBC8Xl7SvErFRtQG/IVx8quTSsqeyJNRP6Z0x6wGKve20Lk
oHxqYfgG492tuc0pIZOmQ8EDg479x2TFfceMsaeY6o1T5GLqozIVG0piminPWYsg
P2bz+fr2kH8FHN4PgPY8kJrypYDbqfA4TlXzC+4BMKIoJX1Ty7L1h0kqiCjkXOsE
vZmooMH6UxPvY6uTqAtuoJxZLX1C+3ZblSWOWy9+zfDdtMw0fr99XPtQsQrSJIcq
vQr73H5DAb7UGLahhSEytyZT9LpfHcHVlStpCaMh+yy9Fqs3JNhAbX5SrI2aG1t2
UrqO/PPEbtZDNFqcPRj9La6KV0a7VMuhN8mnS5Ak2+r7ppBYNlzcfwGKxn8pfqnJ
jdGTD523j6uOcuDEN6qaISOh2y0fdMPaKIGB8eTZkofoihWdfbWE2u9FrjlRw+v3
UHCEYrXTLn9kI87k/rDJ5PRrFq53txaDV1TTzm6dt+wIgzU1yFGODX4KCxBM02jI
qb2xn5aaMtTGtZfyjycLs6YQu8V20K+fyW4k6ftWLFixWfHuxEy2fLM/HYreKjJW
n9+4cvPVWB2xmIXN5fntxG7GnB/AV2I5Xq1oGikHIriyrp865P9T+mNYStLL2UxW
3f51JXhIAzzY+nxpFzgMGNwrikyZuuSlNnnMofX73r7oh9qIB1xoBQYTb9YGGRmR
kIGj7pmZgm0eMutsfbuapB4e8sKZ/B4hi953uov8FmwA2Uso8IwFWDB6HnEtMZVV
fp4I3NJVjsa3WjNCSb3gnjXqagCkVEQV0xgFmJMZLeb1zbOockZOnDGgfRkr/By/
iZZaTeQb7MVFbG/pf2XvNSdfurgKMBVuFxjF7D/sHzYeMaV+hzkupF21QMPjAuck
VbM1LsGW0npLUtEw7NwLc8jfUDau0k6gmgKDfGYCJ1GTf57/kfdkE1PnJ6cq4VIj
Jm//B9DpmP7dR/1TMKastssnEkZbaWTsT8rLawas/Tacjqmud+uQhuYPNpEYlo8C
UPdy2Sy2F7NVZSe0pBA6vS44ql3Al5McZ//+zXbdjdYZkwYZ+gGGq1u90d+pr9Xf
UAj9lfNbEIRyFszFVIkc4vOkVcIDqUqcPBkH28wnPmIJxczGGCwLO3ymeheFzjRo
8I/J3fGGnBFQ8YaX16exRjqK/HpGrhtPzINyG5JRqxE9hF+m6kMYrSGWGQPieohI
IRWWnP9Gy6qfx7n+qALMYpo/1UGaIvKkJGW+XMecOXpM8xXmXjhTwfmtmwa+617l
vtqzvIinXrO5NO4GSmPl/unImICjd/wkpfGLTafp4+M1l3aHELrQIPrMZ4aJ7+L3
FiZ6qWNiKSiT6f3u48uCcUtmjOn/l2+7i+buxFGL7wyG1vVMGT2TzreC6AFNai/c
QuVz+nxaR+ssCPkCsBT+u5Os68RgdKw7U4IRRzTnueKScxS/bhiyoUoA+GhSH8dX
DDGdThZN37GAW6vFv/OaW1C8Liml8ew7OC1VA5YDpCkOHkQ6XljqfOC+N0Xg8RmY
OQ1Rh7o0G3pbmH6hN6+VXfDu1qiWOq/6kd6BQjuGZbizmr4BF4OdDM7sex7IsOtR
H0vXi4H59+xrmNin3kcRtw9VcPcVYt4CeFB0ZBnyrMchvpy5NUSKUgwktfP6TU/X
HPWiKpp4f+eRafqUM782b1ZAoSMrtobo3M7vqqrJBOb8A/rA2NAPQIu84O2/e/11
MkO0M0qNgTupVZllqFwaOPqx0vb32hd1In/Ek5RYkkHFOueTS12r1Babn5Yeo3nh
ikdzGe1FF97aLs4dob/7LHZeYafW7QGYt0k+JCQvozQOkWgmzDD1sIWJ1atHzAyc
DQuWNWyLrkGA+MHF794vSG24+/l5WcT2Jh8tgdgWWqjxe7f3WWknERZmVzwyBpyn
Ad2fCHWH0ykBuQC1/Nt9WA8Bu1AwjB51/dtuHlEyelvoMbIDAlgRxK1xhJy6cucS
2QJGWmj+CmwOp/t6bj1LjvynzaHXKTp2QpJvY02BCfT3kmpgqTY5rImMC4bm2Z/6
4VZVJv3bkFt6Qqrk30TuVU9TJOnj7dFv+1pHbb4LjwiY3a6IMi0fNOKFGK0H+Sfo
jBg45Ao+TEJxzIo3nD03cacDixs+7CTs8hLehxX/I3tWTghjnGXHiLWRQHquzac8
ZLF484GBb/CH7/vl4xBq2Gp99yXqMhgyN3Bq1exe+L9w9SQwdXKtaVnuoyeRBfSI
1eqisUMb07ZDY175fit54ay7bx+5v1OJ4RFzSMRnRBVA462B7ijhD0A/ZtUF4/hX
9pNDbuoS62JQs1hqMENA4qZqn0b3uVrIpC3IYQ/V39DoJGhd/GXQ8MN2lf1J48vQ
JG/akGxu5fypY0C69ACvSbG05/l+3WVm4yOipabWDvx+WNW066js3B8leSXpoRah
Z5VmtVJmYdx6xfW4iUzwlOBhCRsHLfR7Swq9qTnAJPfLWVeZnQfdJ8nlMg7ygB19
42Gef63SfUXPra0XEDLNhKd4qGSv2dv3dISIgRxVOkRhTYKPoJKI8REw6G6pHQr/
IXZrzDj3VEGrtXp1vgdlO3nD9F2P3Cj+jC+aJlsCdXHfDT/vHdzX7gTBqKhP22Vc
LguPBH7m4ShCSw28JXsQtRBS+CRfoMUVlepuvgESyeeOhLNhhltPBo0kN9rk9SkS
AaRkQUOyXUMsftt0wuvzxjGb98o4lgWhCuzWvufVweqxu8ZFmeZHxpZ0WDAVIiF3
9EZ7MLuEIaEE3ShfxyQ+ZaDC/q49XAyBTwBdEw/yPQQsZZzDoaCeyrp5NPynZ2dT
e6A6Oy+oLnXrWiC30E3lRb4mXOqnnQ8Bpc5H2Syuaiz93BGu8JAz7KhOondoiOxL
Uge4GoNxcENqWgTeTZcBaYaho4UyE83q76yjbJJ9hORqzdgORjSz5oEgFRmYatok
+2F1GTBjrJlSGMPxak8/maPRftmfWHt/Oe/jkmEfbcfi5SG8mXfbZKj1QGwna8Lx
7X56F7gYk1xwwTyFlN3T3zBn0U/I/wRXprv+ejq77dwemAs23obcl8hgx1e6p3zn
p+IL6KggaRSOyg5SmY0VIr6nvlYsXxzJzzk7fw0roCewfakbo8ja62xXoperXH4j
mMRtaSpuWg4qqXbwnwzFvGtaHWXZDYAp6E4MFGL8yVuZfaaUikS4gkIusRsgWL2Z
TIMCKgdsBf9XMMCUY9rJlcO3BFgZK6Ek35VRQ+bHww1ONckcWxg4RjosU+rTHjXu
QQ4saosJmeMhApWHXM2CNAwzvQ/Yq5sPwhSx7vxCS50IFUmu9jHAwoqCl9xd5xH7
0I9e4Jt/DlGACyEpkHij8ByhrOKjUaGv8jnZG8kGAkAiQVCDR8EAayxjSJhFZ5EH
i+b5hMjA5+0jsUJIIlpvQ26MVeXETywKEdTD0zbu/lzpuij+cmxQLdm51ZLXlhGD
pX6QR03QAbCy0SPMDFprjjs3L5O28qIW5wcYiapi5H9qzu630wjZBsLtwmeWzo/3
G9lcMAkZlEBlkhPrLIO0poywLBLI2u8+m0Dwy/B4sZcHcqvU60nmGVuCbpKtpq3b
HshjNnmuNjwKplMC/hKxyT2CpHefLHExXK8NkoagfbQp+ZdkKTWl3SzH3o7MEA2c
dL0Rpw+7UsUhM+C7jb9nhfxfpQAQ+0Kq0KuWXWWeUSpR/GQvyaJ8veZ0TUjktzjB
WI4YvGXxuUGMWxKnvb+f9CH2J5LbHtpgHuGxHYZno45MuwwDqifyVKNstirZR8O9
u1EpW38DeafCrfdIjSGWVCQNaKA1Vhl1wQpT3a5XD4cO5s7lTRwOCRyIpkN/Bo7k
vnHHNDmSDohKZ1mpTH9nvjzcoP+/EasboQfH5Lc33whm7lBn6Br7E41cXO74ooBh
Xl+oxm+NG4iBYMfovvDUYXCSDH60k+b7jALuuzr4OGWfes4Gpar4kRmajT0MJKjR
vHBEXIyFSTs9FIVELysabGEfk/Uyf9qVJ+tIBXrCDSaHsijlNfdNts2MqS1fu8gb
jeB0UwDxfCUeE2B/mOXAc+t0kbgZTDIstqTyawQGhhLgKVQxW9UDUc6pGb+SANph
oz/PghkeG7kZ0VJ+pEzGodcB6w24n3zi7Yv9bUYGy2jYfcLtVxQ/wGMuNPKzFXZ1
SiS9uONInyL4Njf5ff8kt8TbG+2ZifAA0tnxYC98TQfH8VnpCW3wRgmi+NeRJKJM
Daxdpc95h5vywzxOcKfNLxXOMX9xSecBVOM86qzAznxF8wgB3nVeV4vdNZ8a2bDB
NMZhNjsRzP+1Pdeh5QruG15Yz+lfBv8NszzL90Y4YxlXplICjL+Dvf6bQyEgMS6s
S4Y4wde/ydbwgRBheklLBSN7hg9IBMjV4UTkWpZYj4hMPbif0mxxadGvRanXG7C2
biD0pF43cgoF3x/h8GwOzWwRKE+eiGrhdcBQ7AKm4t7FbU7R2qUxmiWdGfUZoGY0
BcxuzsKkjHp1Guqo4wOtNl0H+gNJMwOtYXlj3xkZjMCRc1F/D17aCZtiJa61MUlL
755YYp8A8rXsXQs2ymJ2dpECwVRrWbpsBTKRRcJtYGGwhbUkX7S48z/C8ebnkZfH
FVzdhN18wLKnvIqDRxyWDmZXjhAMmnnciIaZ0VTufw9eUJA4dFuH5KNnmZ91NqiB
VbZr6DHkzrDcRHer5FiAewRDmIWt6zPjZ415I8pc/JvTjimvmNmKKlbPifg6HyxS
YCSOdRRDO8XyQMU0+X+7QACknk6O6XFVi6UP4kpr/Gg+GFP7zctaQpZ7oNp05Yiw
hcrdfI7uULGwXUljhu4cjDHsP7W4bpLeEJlHDaftRWX1VFV14FgnCZA+V6gh7fAd
p8WWRKYXb6iJh7gBI8hVoAuppy21BIaPf9IL0F6CuqILoDDbYsBuIyDmiO0xE07I
gKjkFKbPedGvvJBELKMnTFYoLmhqmDLV10o5oPCzp2asEU5+GcwKfqSQGbRqvpAF
ETxMjgxSyw0XEuSp6BFQrejDBYbZreqJiLuljoytsW03oQOibkEsctnT0cFWXG/d
kcYEqX3qXf2jC7l50Fvl/YgGHWdF62jretYMrqV/0OvYtEMWvmmkVuPsT+2q8m+o
d5Br8nMcs2pIWouwI30tF0bJ5Mm894uLfHAwX4Hpcs+Zy0RW6p4aI9Yrfx52PIby
/7VEjmvXGVQNl3zz2tBKKmBvna+4GzGEQwXO1OdGYwOjsiykO1lGgWuGbEIu/o3b
tKo7VPNJlmcQSTBkJDd7nGvTycdhyLw7m0UMXt5HMPpQ+NpwP+QDoqp4ogIZzQaH
Y1cYe8SdY2XuQi2gECXxig/v7S3q457w97DpIq5jITNvMu/KiALSk/bzy32TI6YZ
/bxKHx65/ZHA/DLW3BPy0wiZSRtM/+ZIruIbUR4zzyhTn48hwaAfKexe+FhTniE7
/OjtzLUyb4IQdMADgzqwuM2slusXc8H6DO73wa/WlCtppg0g27Cn0CwBtolI5QM8
P9P2ONj0+oWJawPMv2spJc72GZUnZppGlRicc8BwX9g24UEd0S2q/0SIibG9UvWG
F3IwKUklfcB6rK72FkuZGDRjmD4kgTrT8CSh/xlF3l+PCONpucohc9wT8ReObt0o
1zdqCPXJA/7POCKaOXCa3l9LUQSdWPT5ZsTsnvhWhki6PSspeRshYROMFbFdEEr6
Wed4C0F7xCpPkJE1qo5R4G67oqkbSeK5vBL169iIdXXMfp6lzKBDEJc39oWub0nj
XMFctnkUqmRNbvnHidlrHwNIaqPJ87gYnUhp/lmG8fGfWK/aMu87ZW1XJTZizw0a
xLqmV8psS0VCv+csb30N6zGsJVvODigD6QTOzr0dUhSyCviCDM8h7Bjw3Pcv69Zg
dbFTZpdE7Ig8AgiDHO7QzPy2BuvyQbGo4G1WG/5e0++2XhjyZI72qgfozmRJyiNE
LUPOLCzOHX/5fP2MBZ7YsgWqXqRvc+6oUBglA84JGPwWQ+7p9mpmSokN7BVrqzkM
9jKN7B9+d7hIzJC+Q6s4teepWYBXof7hV4KBRMgszdRuf09FemTezQdtn9pdWU9h
4ifG9xg5eschbndGv04mUdw7nvJ7372tahfPTV6DOdvJDtosS5hwf7JENTbTx63i
fD/0EuHNzqVw3tT/wmRGZy9WYfqXaWr+O6s6R0IYWWvp2nybtTQT/9ec+oRP4gew
Up7Ykkt2eGCWo8bsvv+3poxLoWrcYTIJ39vdSTFaCByEcDCrPQCq1y1CUVzxxqPv
1GabT8CsUKfXUU2BNjHXUWpzVANT42FNl2UgfsIdqLWniGtJhjdHuNbUZZb49lyv
Q8tFuD6DV5E8bY4x1GLHTKy1kJhnzZF8EXepLNUmU25Xekkw2bQcqPsfA+6K8dbt
HoRjwyUnG+wMnMZwJrYw2/llKkKnhaYxts2QcXqB5mPkkk9qPRSlwwexGpEIdOLm
Mb9fwvifEfrqIDnbATwuEal4tqjsKLeLAz0KwI/AlWX+T5LdFDaG5lTtEU2kXCDr
/5OQKTjXmtR9tSn13yGTFUhI0GKMnPeRfiDpw9NdxrsjgShFh6l9CReciRJYE3PI
6xuuJyI7WaFYheTr1jyBhMv2K3Ig2YY87qlIDSp7TaIaB6MpQ6LNYvZURmsu4bHS
NCCbk0X1LGV0AsJTVqnWe0tjWBax1Dlsh3SU56hCKyq4ddgk8By5DVtTbsQ4U0D+
eTdQV8t4Zt+x/ZF6Pg2iZWJ9W2q0Kz9Ng60Gmcc5IW9MYM3JOaAGVNkCc3UEG/+v
GkHKZWjDEF7AzY9lE95PrNA/0+ov5e1Y0Q2vAuptjilUe1qTKb64/kqgqFuZDI3x
mSez8/JQ/5BsBiLvZTVX5oPRd8bVEMGdvaZc6ecP869fzTPRSQ+w+T9b0vvbaEW+
EqmWIxMGyAPMlzySvYb1OZ9reDBI2LMeSM1E9RgNrj72bmWfHabGguIUK9mhx1IG
n2GBgEBoU6jdg+aXMD7i9NHE5Zb53dW0OQ0ZVqkj1lYODitBO9nShK7zvpeiueAR
KTK4YhlVev9kRjOv1PsAt8Ak8GXkxn64wQKmGrflO5BAkx9n0h1HzGrCNq1zq5MC
xEA0Geqd7Undptax7tnIjsBakWzeyIFyzIt46GfcL1ZXOOE74ohJdG4d8UXnrRKu
RX+NmRWtJtj7KegPwGp0Cd4dmE17aO7e5ACSfNpXf7+Np3g836rZ9k9eIR3L/6vg
7LVr3yfRsDPcKZtEoOmvFSiWXMSwyDpC9r0KRc1uc7SpkmwTGXrOFHONm46gQmNE
kDXkMAJISeZR6lidHlIoO73i0d1tK7q6GZMCg7cTy7xrZjscFd8wEgoCOHppq9vq
HAqSeqHoU+951NS+3krfEXoRps2CWMbxLmEqlZ2QURXL9olVJzv6GK/yYKi2LrPM
z/tUnvP8UBrrh7vYkFNqvDIGKL0CjqmmR2JhZJurSaCUaXVcWheyZFWNBEhPS3yp
vXQACGyF8NBYYtpUvxNJnbbKVf72Ltd7ZsKJzd+K8xCJdgIZJ7gdy0aEiAyWUXOF
w8HfC7pXShCCTdUF2DfilX3DEW+pwvexiOgRaJvPBk4iIgnOE9PIA8k9/eTYKLIE
vPgguVhYWW5gEKOHN5wwf3YHFRdTYklV/9OBcvd49Y0gb5rhsQJQDr700quturIk
oTO4O1xa2YRKYa3GiJbq9H5kzxGKqIYqRYUeqlhiyqrSdy4bJlAxdct/zMZ4bdUf
njhQHpTlAjJchihmI7cTRPWi2Z81ybA0/uWRIB56XC6vJ5u6fIql5F/aldPNQWh2
nUotvtzC9otDI7T1kX+C11U4SjRCeWUvuJnDgqwzL5GEeYFQfIWDLL7mtk3B9eZ4
VClqX/7ToXjzAhabPmid1eKIrPj1rPCiX6XY9TVdDVYtqSPHRgoD5WiqYOEgMKZy
DYHYf9wwcamffNc8DpMRdulJ64WZrf/KAVAeGE5dL2+2ypy4ABXxG3G2gm655E1k
wxgVA1dh9Iiw+0vrigfzimrnQNpCe7YW1H7PE0O0l5BTs3TFuR2Nw3XVUTCuMoo/
tTapH7ExxXgnRCbJ2oXvZQhGE/hoXzmoSL62YKc8EjlvwbiDIML2mwftZusIy3SS
7YdUanRTfbtnWBtWC7/6Zli63YRjE2mO46eAwSE+8BP58G4V45Gn7q+v7RN3uiEP
nSwntALzl1qkR/kStyCyLDQ9SRKsl/LwcFL5FCgEy9v3GFd5TPMsvn6lgEwkz+Lb
MBeX23OyCzUEZzMG7984JeX0pmQGlEcz926FbVqAHOTuicqeuelqFgu7jZxCU9Tw
t97S45ffH6yz4g88LRFfWGaGqCzXhQgQolIgDboQDvaT4ltSGu8YiVK9Rt9ZibzA
p3+lBeCEwGI1eiOI64cXBxF3C/gVSgPzP3R3muAxHiNWfgarMUbyca1TCedtZRTM
sXWd73irpp/xl7CnlAXNOasRPH2DMXQJNUwNbeFGxU8ZmpRz4AytYHYpkH0FJslC
krW/+knuemMOpBIKFyCOCSTsiylqDoFd0kqoJr/LOogfzWnPns8vuWtckgBPmHLx
oemvFRV3cyp9qJjyinS0eXNJtMk+BdOZKFyA79NyP0MK+OMdCUWkAlOWo1rmmKi6
aJ+EoMp5gh+juB02jqaj3BnJlsB70U5lNqWkXzzOi9y7Mkoi0fiEAcDRKRPs8Zfg
x4li2C8N+purLbsNP7KECNVXWF9Q9ekvWng/JoMJNrbe3YOsGFrIgsENzP6vPgsG
jBO0Wfvu4Z/LK25RN1Kbz7pd+SMwuUd37WWMLasrYOPXNnWI4w1MfRe4r/LZimJ1
QngPajqw3KieQ/x5gKTp53JKp+tuaQgUiW6ndIXc5+/s9hrj0aHaBFlU8VI8Ydci
q9qDENd5xjy18I35k+9kA1eeyjF1cIrjSaqmUIYKq1NsjbDhFWpdAEWCpfoJ6Mz6
PnrezRvm0g5QHxuZS4N2tRen48AddTdiJF9Kkx5LERUySr3iz/eUiXi1Y7FsJ50P
PaNZlsloaTVvDJeCeHIUA9QAXWXVl4f4WFxQ86l7dyiHPhMK2blnwZhobV3J9bf7
N8WRsj0+lhi2OjuwoxIem1jG8SfPy4OVoLaUHs3wn0FjrfdF+UCoN/F0hCjMT1VV
vf+y53BLmj/ZGW/l2Gd9ZHPXEiGUL6Oeu6imlXa2v3dFrNXYHbG2LjgNa9yU8zIR
8FDrbuu2ZhmGylx51vLGfPlx03HqxxyfFDNbi+QNYOp8IXAiEd5zdb8QI00+K5c/
ixkwmSTJ5L4KkrZXfyEP4kZmaILpjua+0iGgl4jbAvNz1Ody4QvOEEEzu67Wr23Z
r0Z9g9M3uZFnHhtZiK/VYg5Q7Dn4GfuHm4rXFcosSj8aY8NdYsTJvQUpHNHZc3bq
eh6IZNQt9nh4LCPv869LXkYGdQsEtBlYcBClWgKKa9NQqeHhgRXa0FxioJJ1raZC
2KqxM8Z3Yl21NFLs4BdptcInu8Wj85IwTe/YXxIQNstKwXZyzacrJULsbm5VYQh7
1kKGHbJBRiu1+C14cJ2vwmG/mDrFuRH+wV9zNSsOTfBAaBMUvi0URKfMqCJeRJyh
dd7/ne7QRkqyAYsy2K69xgCDLZrL+P5K+LyHqa5CJnDfYHlqfAMuRm93Sql233py
YhyC8BkmJS4HeTbgBmBq1gBnGnMpXe6QadFBzpL7BOtPDk2oEox1mUMFuPsRrMyv
BZJ/sTdvyLkZu+jdNcCz1ClQlePon2I5KN6fSPasFU7TV6KMGURkRO6cr3XyCaBk
j5FJqcbqsDOKvgCF7LTJ9Wt7fMzElgeML2DqyY3ZD7Evyi2CylPuJgC733a0AV7a
JqUywCagh4UD6VlK+qDIIFbLio8HOqHz+SKnPWxLwqCl4R7mAU8w7dQrdO0exj6K
BULnaz5C5tA4xPtmLKXeGtqLB8ojNbNyxJaL63/y6Rpb5hyg0n7Y4HuWr840321J
pAp8QeHr4klHj1CxxEA/34NUJeIq0S7rqcXg08J8sWTyedBKzzJU0LCN1QWanZHa
ZRklcbXz1N1B0Df+m6Wwy9pl2j/oYvtdQy85uCgvceC4i/UY4nnKKPkoPH3KDuz/
++D3GNBatRSCgj9Ysu+XrBHpsAIf48l0s96lVfK2l3RWwfjPPrJzOtGYyR4091bH
G02d90JNWKUwgM1OS69eLuQdSPiS5n2Z5bEB+ao0KUXCfurh1nVbXMoRsrCydAqT
fijeJzyad/Np2UPP+gR1QoWxWW6KyHCrOvEvhEzM44uLenHgzoW2K3prVfgCwty3
4hzTLxzbB0xSLJmXaboR6S4Iy1Qx41a3zNx7kopRFh5rnM6xRPX5BR9xu0E4sHcP
u20QwG/EffskaSAmnLQmZBkTI5dc3zfetwvqD3p+cxCOFMK8r9XqdGUOHgEv85ok
1latIlauKZPXUe+kltdDrmzaBKGlYcLxNfy8D+GpaXeksync1Z/0m5aGZHttSb2K
c9RNyCIGkMaxfdoSZvfxDpKiz8V3NuUtrCY4UlmY6wRqigq78ZxwhZriS1uU0Uw6
6HefLruiJ2D1SCBsVF0RSKs7iqeD9LZb8S8vtB8Mk2ZPTuhiqAHjmyJN26sm8SUu
PzAmB76IVKbkm6PYO/sXz8qa6pRYT9oMU6CfCKPnJdP6IWomz07wJb1l6OKkaK1t
dkcbxJTVk6mkfHZ5PC5GEcfWmpxe6PGZ38MkNKaQlvrWEi7uvpNcnWsTBZ+qEBvm
mmsNonCrimyBede21tIhvCRQ4h72bZjYUh8fnWTKSEJlLFWXghU6bT/xzVP/0THZ
C9Pbnkqsp6U5eHu08USRJN9KQEhJ/lnKV3/OUJYxr+gN1uGF7kNIdFQd9nymqAVA
IqBELKpMh6vQ3wD+0+a60CSZelEzYpdP4ijA1k7YUuRraHqIdotTs1Ea/SdxJ5sk
dS9RJkfHxq+6WsbvVStrVAVKH0rsKbeMXrgSmS34CoVBYCzPHlrEqO3+FZ9CSyKd
9eMQJRxkZyjNfF6jnqQtzJKhPqB2y9Ud5har5aBnE4hYpmzLOXbMXb3D82qGyn8S
bqv1syk2NEJ8lTGqPirRfMUcdec0JvKRoLtx2qn3afI9EkBYxr//cZ/XMzXLWp6d
pCnZXkvwc7R0TIB7Qtedrdrvdzq0Wzl5NQ/uLKXMDbchfQ10auIeZAzwb6sYc+ik
/ExRAQ4CWMvUctXesOWgMJPWSsd9HT2gDlI+Q8s3eGemwy8DfRK0Zhe6fSVBvZrE
rHROXA3BVuEQ20VFjqOuKfIZMcCbRWI0yPEn7+GMA80p5Ku+pr+86fYAy9X+rsSW
HjFdlwMFc8C/dumliD9EltJ+M9fbMtr19XH4KMCFGdDDkYIOhY/fUl1doJ66MAy8
DVSR9jtzqp/2xS1Joj1ogOXxeUnRATDuiG+P4jGirtK801unDSka3n+gj4lrCtsO
MJ5iwr3ZrHnKQWFX7wIzLF2vkc7M6AKJOvzYBPu4+sdMq1DEqNiTEls24IW3qzMb
u6v66dJQmnzv++zdtPseLMjwfWNQM3HAbKbDYLPlI2gjc3w5l98TBefk6bAy1aqt
1unDNKdw9gG4c9tz6pOO/yLHW69qNKnjoyUSOeHXfz3x0AiEybklO6me/ZQYjQ4m
dYMtG5FwhR0Q8ImrBIN+mFlpkRrqBD/4mvzng9m5cBEGqD/jMnAFGR3lAV1NQPVH
FweZSxnMCx39l13V/rod9XuT2gbZGqYIYTXXtiivRE9jlC3gjQJLxjN1zCBRS47w
BFMcbURAHgYkGgt/pJ8IvrRsOuLKdbrUuioqiiYg1jaSwNONIUTXXTE7/3riMORa
cQYvj/6oW/0tjtbC1mWIt5Wnx/xVYBtwNfcjwMfgvkKEQGl8Ue5l45zAgL7+AH6T
BwMdWXkk4hZ92lXqhH2rUeFMSl1OgPVdyrlcR2FoY88N/u4z/7bPKaaZ+ttYKS3/
H3fFGShq6jUtFtJzEqD5GGM6x0K/f8ZPdTDK3p9YHpsreOz7ZwAv2UfCIa7i5PI4
7pj95VVZdk7DXb+aK+baB/TreHTUA77IhtQ9H4VvGlIXJVlOPbIWz7jIply3tJ3n
MkqSIaxw9aS9En1NcGnd18YL5zW6jpaxLerNMIe99dp3rlvCQRcXWUslJJhTalS+
CDkHZspANh7fC0Ba5njqcZjphv/0m3+MSgqeRpdw7pQTy+m645FHqUpt8dCwwbH2
OPP5xP1eA6WDpgy8OD2K4qZDLNDLj+g+BkvcISqT6OPSXZmbmoS/Kod9DElP8Uhm
eoRZd0kbrZvdYbs1vbXTSTBeTJLYlTsTcgTwdsqVvOomTuh7AfFV87qQa/E1w73N
QrkVton3VE7MtfR4KTuVIMvK8rUx3GN+0VpIxsHICa8pZZBzbtcGjt6SENJzLPgf
9DaeGnu0IYWduwIRG+N+B1illfIsgB2V6NqD3y8E65LqSQzMVe1tWjL4ZmMJoNFB
/tv3/x4a167i5x7nDLGUpmBUHKXORYrkTw6H6kq8P3I359tySJCubTk1QDi21g9/
gR6SWD+++UOxNOUynK21tUnCHUVsHqf4r16q8FK4oBjA43urEG4DxIpK9zrk4k7N
z2aZ9w41ry3w0pYVa8xDkKA2moS0RHgdxhomLtbT+oP2JoTeRziqcM70OFMgJq5S
KDFHrPTOTTyRvEhKg9gaHeQFVhht/UiqRrCbnx6iuxl+lqxjN6BzFH7GU5Q+LAwA
yGUgEQklaNn3Mu+T4gbVTZY5YkNiugqkaynRiUtr1S/EZ2dZh+gx6bC3FaTCHGHp
td+7NTN1q757NOWwG2MFTK5rhGt62dU50KRnO/fOKl99LByS/YNu2B/MdupJ99sA
GF/oqOD4+KrQlYwXjK+LNE7Foh8fgtRakMVag62GtIlk2DwQ/+wsqyChOLTqC4g5
7r4iWO4U3OjEdyFU2E3aEJMumiZXB7dRHi7ESLCGu+UNo/epc9ezUsaxSfizAgZM
HXn4D6kbryPftMPjT+ro3ddCUngmX7rmcdR9xTswmJFxUKsjdoQohL4wsWOyKI0H
1ulV5P/GW0PxT4FO7sJeoPOqa3UZ9zqKPe/hkNjdoZv0vQvP9dWtrhDk9qHVzQi+
Cj5dPw1g0LE28PHbpBrqTMA7JKgnVCtVxGzJbelguk3Ac9l+OfAMATpn4vztKTa2
EBwiEgNeYRO8njlpUoAm5RaceXYqrETKEWudxJOBrt5ifhBkGXnJCUGKqEvrWGlv
Ma9RSq28pvP7rjDBuXbUolGZnrOIsbo+FmDMDNf7oscg56B5ofxgP0fegI5sX8SZ
cgHDl8jqExxKud66ewpLeYO9KJHt27FUt5vKO72OHhnFgnt2L4xolMGZNgB8lJfn
VPtTmGWunL5M3Z2Bb0JTyeceHqaLIbdGgBUc//0oTfARG+8WC93KWKNh3HuGwzyD
GEo5uNhWwmMTx1UPkp/+ZMb1yXkxb9t9+f3DfcaErcMLGdaju1SYzH6wcDPl6tMw
vGARJtSwH+d+gwX1rLqtgqdteH9Ie+wpxugyHFAJTaJQLJOK75/h+EQ4PCEq2v0M
rMX0vu/84o8Ucqf4lrhMD8uL+2a+5aettUnebLDlOzP5xwPHoX4yO/eYtSGRaEyj
+ujyjdPqr4un0k72IDGfFTI0lij6Rmch0tqls+FGQGZLAELJjoGuJIsjdCY4ZdxD
73np7XkOG2+uJ/TNU0iffn/oNXKPRcqwOo8E0UCDPQawAMxW9/Dueo3IY5gziAko
iW2YAeHehGA7yG9nagzSdrTfzA5v4ahokHESJCzPVa2A2Ft7l+ydgxKLWBTUceGs
t74t76rtpIVqObbix6wnTmYtt+G2g8JuszkfUhmmF5TWXbYC09F925STes/u7NtG
L/JhxdsswXUlRusSXv5aqrdXBrzQULuFKlV6yXGI4qMdxBymGnkWxQhvoRGejVa7
Hu+7K7f59NjV892soeiHCmyJratNiSrioofdcbbe18bXjTAG5G087EnQDCvHntj6
EcZqkJU0Ghaco36Kv6HDqwTkq8Wd86aoqlDmN+gOame2kJsYS3mTvCDw6SJL5HEH
zZBzPMHkbHNaxn0PALRXrDzvj7bSp23jh6kIjbnP4RkXe3doyK9ErEjX6yAtxy1/
s1MLN9NxBkk1Gm2tMejpMikfccrt6hwkv4+hx88SMjOarJzA0HnfiOzx4+X1mxZH
MQFl1OLpukHQSQ81LydU0ywr3mSLs/MBnUlZcjVwo9bhLWgm5rle46S0/3+SRd2e
Bz/tgXTl7W4ZrzHoM05lxYzNF7Z3xVkqYp1OerrvWBBHrZqahsFPed0d1hwWDddc
vyzA0MAjCY4Tb45CrhI7Is69ad6v+6c8NEPYvQP/JLDovdPWZfIQYH+KHKMmwADy
aKzS+0+1FpxtWopBnPuw4b37OMG7FsE+6P4gseOnmvHvjyF6OX2mtwj4cYoUcpRn
NzmI61gyT7/Yd5RrJzpwuGYV7VMczkLinVqllcUWUoo9OBzXTm6BJeN4Eqevmzss
oTXrewugSSQ+BjzmJ9vKKYcpybSvmk/WT/mdvcOBg/K9JQ4cewv12nxKMua+LzOt
/DE7x2aDJbE2dEHgER0MBH+e76KvSiTP/G/OFW+oTQ8GGOxzAj04rrjWb5HI8jjp
rYeXDoHRqvbv4wUgpb88zVVIdLV+tTlowYbH3fa4Hn4L9AgJOzEcex3yOnmr8bRg
ZNAo2eWhU0/zRZR+0mtS2N0mQ8AGfknVU4TogxsUiK++BDnXbl8FDolf6/1NQt4N
kSmdxZNQhihGQ1SwRUUjqmtZzM8O/m+cW5IJmQi+x+ea/uLsEVL63y1ro5P8A3Mi
hyZdyYiPmLlHgjBnpH2Lwcy5/xN3KbEOgxu5tFXDjsuK+9Hn2OcqbI3O4Wt8ffLd
lObGG582xUAMxDiuILFoQkbd22G2IGbHfqT6XpnLjG4qJigU+csDsq+N56muRFmK
S0R/WWI6TjlNYm4qFnb/T+9pKK9OHXmlTMXamI4SqO4yVAGrD3jbScmzRes/6WV4
O9YMIDYS4mlHcbChxNBGaZMRFEw2Dvtw6Z465ka67IYMVbEi1S7UelKv5Hd//SgM
eeLX8DhMcIymNsqyWY26DkQfuupJoQd6whiYR/bFFfaqS4drDMGtiqKGw5qrC6ky
iakYR9/oHsQsZ7KJiy4VSEsFe+Q0mPktZ+ongUiDm/Zswl/SHNj1Lg2VLneuHEiy
OpjlZ+w47yiqGsSlaCaI+2qAkkvPDvlVbwLZiX3BjsVPFneCgBA2U3kOR1U4NI1c
5Ns5c+lD7x+7TXxDEtdQc/yt+5ETrltNfNJ8a3MziNdN6lUrLyCDP75KrN2fMej3
Nw4+ICQe6C+kQwJDoCesht3o5qyTkR4MnQ0S/koAyR6Vo6SCAk9qmUbxax0S4Dg1
JFejRfgoVx2+ihrmqKSUI9Wu0zUGnVMF5yWqIw7Dk9v7Bvx16WFX+HiCUAy+Zkv2
12+ZqITUQ5hPy6byDXuGish7+GViRijfk7JyVPmDvuAUbV0iEwhPIBpFdeu2Nrbm
bpvPZc3qKhjZrILW6o1Wf7NOqXsDz5JOCGh7IqLdaQOSidQbsEIl5BEQHxfNvhgy
x+Nvqg+LiL9UABDbuMcT+9WZRwhIrkVFUCsvrtiQpOgsOr6fDU6jFRbjEowVFPe5
vdyBQjlBEVgYgCvQPE3ZA1hMjHJjXk09Qs2qLjdfPl7aJMbtnBMNmbYuKBUliUBA
hktAPWbb5UAEKa3RbaaE38Cubin4MTfGQmLvJYv1/Is9v1Y2+pm58ScAOW6wCgVV
u4OO7sQ5Qua3TrEN8MoVe9TEQAzVTpnWPww7H3llAsZ7bunV9g/liyQGj1EYAu+/
0Ym2Cje+fotdpAPDIQW4UulyINUe6byzw+VeW+t+Zti+dbkEhBgpssZ4kMvyCkjf
PfjA22HPfXNboQxJ5bUk/MrV6rEqjaPuN/fByg55YYaxbMWeP66TTNTzgyvdLZha
I4wj+k8PHbYBzPAgjAH1MaSKBdFMAYfKsYdYlsNTKlur4atY3jS4VBNTkzJsi9u8
3j/QiARNCMTi99mD7BW8qztL2MmWXXv0ueD02Y4NeicnRYEVwN8K3aHaUEDVdQG6
9Bp76QJky7Y4KKI69N0IlFaxLhJAy2mEsG2cCgJYl0BBwPspxUwG9/3+pVK0/KcR
2PMt1bTFyPqHscA/Y+FGpGADOKOefyGR/SNz7isLYYzd7Rv3g0dZbb1acQJ/hPNG
Cerm8i/YWUhGvfWUSPuZTOQZQp/0oQCbQSSGPEzij3l5sSX5/WFiiN3UP+BeouSy
8r529oLiCx9QOxRUkWPgiZSo0ufAUUDakisNAO8SmxklSqr5jXT0yrsDHPXYKE5x
MvmafxKGP1wZA+Wp8LcT8r0YAH0w94Gys0hOoGvS9hXSOFAkUczXZQqJEqK8eeAP
xjafYy/B+SzfcV0ooSQMAtbIYyQHXHpZTi5hu22P/iTqcQdj/RujZpdo62LzwXIf
HHwPsYhrhzXThcCCC3d1RDMUsHb0ErHAA/6YzyAgKJFJjkdbdvYyozW+hrrToZ9Z
RMeuzk8dggA2PRWbIzu67NbvH3OgcFJObztvIQIdOmUCeKbRQo4hULFEgwkNMRy9
mdLeCvgaWjmEXNXBPdrP6/0e9+xk1YcyC5Qs90vJWhAg5fRUb5eMR5Ys6KF53FtH
KqAB1ubDoiV5VkLPamxWs8R6C4pD4Pa8Kmtgs8FZRO/r6Vi1ZNXOwIAg1RrzYxQS
ZiJgThfYNWfc8qFy37RVlxXlD6mVRxnoYHahDTjlewyctkc75AFbsPr7axLrzFUA
uJo8wYjirAj881dD0VJPKNP5NTX7/IWyFoSA4/JS6iQPE5kEiO0TJn2+qQgJorwU
zu4r6kxZVhtGqY2Jhtp1WdZrvEVv/WSOwz1k6EBU+90s4VcVqJbqUU9FJFwBjhU8
pTczOPMFxQq423nlrOu/f2erp3stD34nxhvaNUq9wtZk3kxA/iyVEXV83hRhxHyA
BZeAk4QWJrz9JmNfHeughMVsA7Cg5gOTaW2NhgQF0P7+irG2xR89HctBwxOIJhPb
0fjrNmWPjendyhN8l/UomWc235IMLSf5oMNvRiZ+IdOwvi3BT6LOjLAAgTeI+gFM
6KrLh5nf/FBGe7rifA/vDL5xQV7Ug/a2hl07l+gtjOekmcJe/OKnPTEv7dRKiy9D
E5/yzPUNBRM7U7hYAwbVSqVyAApl7en2X9v7b4QPaSRAEzlQwPZiY4WyelU5rR1m
YpDdXSbzTsZA1U+Czm264lXVzuTAB4jAXGs3QBDyn+2NM1BZ1jhlbLCcronp6U6p
M2mWkeLOS5FBAuwY/l0tgAzOBPGxKSG8xUpZ3RKZTxsaTR6rS6m2F+kGmh+fRdRo
SxQCu3uyhHzdZN/5zeoATUl3gdxWg1GnZP3gOrR0Yb3RKcLitSX6LpNkPJhB7FqW
N25tsSRQ5fn9WeqdQhzXRiLA2nJ8H7AFaqIXnEswEIrHdjQp6thWfLWPAWXQth8/
JwjeR7z4fNDDoRrdctILXK0D30rH998+2op1mdK2CP9SXAH3kVh3pJTvkC2esXfU
li5U2YERS0kfyZEPWT0giDPqpH4Nbm5b9g/m7UmVTpH6ZOIBT2opafRtGJ2Aa2a3
Te+O09p2knTbp+D9HS5H/Bys33GUtFokIpZf2LyV9mwN8F62GRCKiyFLwvS8uJm8
mFhzRUT9x6wTbeP7EsOHHtRPaOti9glW/wRDaC7L2RhDU9Oyu30iqLS8B7aXySxH
So+7xKEYUw7vKo0O5I5gE7LTM9oGBB2zZ4XWjBjoq+obT7koVeo8+F1hZSyb7hJL
SFz5KRz0myc2xZl1PysjBPs4OkNujRzQCuggEWkM2pr9KWtxqe71gYVid2d2hEij
hBqejKrguuILd2WVGK3jk5nyppQPgmbIJs7Ww9wQJiw+m9tZwRIfzY4x+YpalSpb
CVXNv9w9nzbMCRX8dPB/q0W2ZXE2ylxZ8sM/YqawOsEAhejvsgnteNJ8qpxlc9CE
lGZ5CeFJOdufyxJhbxv+dTSy82Yc0DREnsG4OnyGdbkcmp0+CX01dfaa06uHlcjM
R0Xwetk9ATcFBNS9H6f1RyGqKEQij9tTdc0Mk9P5wHZzmM4XUklnfdGHtVz1oNNy
b5bIw3mCmp1S4e7kgPNyn4xg2VDachDdtLXHnvhfqcqEPLqHIZuXvf8Lo0+BE9im
RGwCnly6g4nc6sxM6Xuk7QoW7So16FumGB34NEkykrhwIhP7Hus1GomzRzX2SOOU
LaXmuAGM+SWrG3iKO/YLZD4GiUo0lGU7twSJlqxzh+zKc6ySUYGFQKfuBl2JBmeX
iQacD95UdN0RY18+v5HFLciMKCfwq9OwzU9k1q8JPeSd6GUBch8XV6JBP88nuzUj
Bnzs5e9wFRmnZ8eRP62Iln4gcffVQRu6IyBNnc9sXc5HzCGVvv4KWhifoks/tift
MUN7sSyPkeWMcNcZt3K9DGnaIi5H/xKuhOgl32ojTd7xDeQrVTflHjHq2DgTvQqe
vEmWztQImf1RWa0EmnUMTb5CUDjOnPs0hYrxvt9zmCmQO4PhaCx5QqXFNVPTP24i
2hqc8uu3JlaeLFP1mB6TkwmsDvn1OrguGW7CoB0rFtSx6qwmbd/xJT12FN8AI7fm
rQE4S8nbcxGvVOBNBpt9/U6D9VpaDaMfs1dFuI0iwT6Qje3qbVPckf+NW6L/gt1c
mxvyd6/JDSEJbHJPLEdoT1RwkxOlO3Q0VvgnQik6e881w1XrE35khAd1dwO2WJI9
IpceKvrZgC84lWSrZDDTKZyR64sviJvJajNcj7hI5bWJrKX3Ud2u6L3f/6UmZvfx
WaaEgoMaHAqVCe4DYSOvR8qDMmMcuiTJWQPe4ro6pBbYivQuePLtXCBE4EuWP4Y4
knaM+P9Wvmtb43d9HeJK3RooL22JQODF3yuqM9X5zzKAFtEyrydGhNMnbpQtPmxm
gBKLsPrFglGiEJgk4jISfQqCYqwx41uP6vgzdDLrDU3qSbFLkyCYzRFT9fnxWnR/
n8+2rkGqiv+BGhOW+zipnF60C2F07EdlDnD/RalkK5OLklOctdmzg3Hp2psfmpOv
hS/Pv/Yuhkr5PzLqOhAE0O8LEoPBGM0FJRBNbChPXQsIMFLErtVqjsvRgCdaHPxA
zaR3+GbwtS4NU7jNW1ViYE5NB9DWev3Eye7kGZcA1H51Svj5FPO6MDx7Hi3TLmbV
C8e23V5//kYAD3Lh3PmhhzaV6RI4qwHkqbF1GuFoQ3AwN+aC/Gs6rcyAVm3/dP6i
YKN+4hW3t6IwF3sM4hslxk5qDIxHsMSMVbRNscXd3kNW+LZxA5cneRqtiD2q0wiM
l0Zmb3LFBv3hzuw83poId7Eq26fCYuYPtN5JHY2+j7MC4Cah/3QDqSPxuts1Sw1L
WaCG7w+e2xaZOu72KSU6vObdICPcaey0WGuZbQ92AjJzKIvviwbyN28jgQ3qZPcR
wtdgBxrqZlH8Cc75pSKPSDcj8W9U83KDqeyYGua5n/vqkXOvIr57Dgug2wJPY72S
4xvZinR33SJRyKTXH3zp35HGEEblJNy4H85uPixSYhcKbTs/wl6F0LRO4oU163z/
URxvnhGkrK8ukUZHdAwS7jzeSh46kULVCNtX3+oXK81T0koM61Eh8o2LYAj37JmY
ZVPUbsrBV1rUOaCpieLGltzxPrlxUHKBKEsobJfnedudF41aHwQvoFpTxlCipucb
pWIZvC2nkQAiEtiuBNyruh24YkOgpcic7dj04xFZPVLc38bACzwA45X5sDttR+vR
6XMboQYS6BRxZ26qBw3TsysQmgLlnI+ZNOFbIOzxGNFXz8ouiXFN9NYW7NjuSc60
9Nzp8MqfGu6xdlNUdHcp0NZ4rVwz0gaOTM6SZ/RyWAc/mHZxWA4B/BZKgutUY2cW
WK81ZP4GxN85wEuQNJRxpLo9rvWi5vVP/YOb2Yiu08jO872FioW9EJVW7HLOCE4p
j/dFPjyueZcHHp3A5OakzzUqL9BFP4a3Y9Gbhs4Sb77UQw8e9cw/TI9KENnZU+9g
WpMf9haXi21BQdMLIThwjSeUYLq36FO6zbS2rPsdngPcXN6iZdCJgwzL/RufZSM4
bzyDaNDbNx0EM7RcLYoBq+FbvbKZPe1ONe+X87Hp2CGujub0mz9Al0RuusvkvECR
ePZ5BM4TPNJiGDepUiwBoDN/qGKsxYxD0F2mbddOqrso7GhFdhHhR8rHGt/jvnp9
Ay9//KI64sQbL7WvfQFsKIZQnKShGCKhWDi2Qp909JB8Sglr3hHl/pHAXTaK9+Jw
5hIlJxb4VKtPGQSCnKJRqXx5EBaZuagJuBRaAUNWGR41O2h/DLIvSeTVuzmaHIUi
PfzmAYxD/tF7rb7Na3pidlPydeVHXPtslYopglhPJj1nAITRIOeq3bLpWhhNLDlg
I4ADJ8/Ib5H0WatZF66Ja8gs0AGoSSrHWpJ+c4/4b3DyZzignSFFmBytLQ5aNLC3
8u2O7szP7mhXRz/35ADNd4tYGI8wSiqEAiRDWUfZFaTIroQGUrYdql5F9P15IEq8
TpQ5+J4YnEflNNuts3uPN5wSlHgWOzVBWwdMOhDbbcqcWmYQNaiINQKyX7CFr8rw
pkL4ly0q7OVJwo8GkWbSJogDcwln96Dqu91Ppd9kEvdiuc4VEjTqFjjrww3mWWd5
KN5rUJWFVKce9ymJAe4zkENj/kXfM4pwkliFcWpe0voDuSXOw1zs4x5HH8atsjcB
siRyfFgKLNAg39I6hPX7Ias1mEu1z5uhNgFHsOe8hThb0pZUsMYIAbgNp0KX9M8y
A56EUuf0LC3kcqTsMXW0+OEEAEWFqYVuWL1QnXNxv2im5aUsgZqqx/YqGXeqSh2S
lvfU0kZbh7QRPeAQTJzMRdK8Tl0VkZea82v9gao55z46/xO229sLK5ba/15ImJt+
FMCy/LjNGKM+tdZ0R+Vu2WJeRbjVjTQ5D8KKZubvMNQnrE5oC2/bJ4EZPPlkZaj2
AHSwd3tfsdAHhZJNINj+IA48/4HFvIpOBmzgC/ih6BUFhAdrKIzYsxyduzl8M4oJ
3YNX6gLQnVzX2ACbw2i9BLQtYXjZOLaD/VblI9xBk8ODXeae2Sil0SXhZUa9it6P
81D8NInhfDct89y1LPudjLbgAztfbBDON+5gKyPh4v1lxNrYnc3kz5tEHuGWfnBv
XWUjQQFQBxCSPW+CF4tm1oDLEF3n3iY8zsw4Fd24MJtSIWtKYzjGumY9y366zSlV
jRWAbogTtlKhSyYFe8KYGpOPt+QMnCwTquRe4yHKpaiDlh8HhHr9xTQDpXNRfPmE
9U3g8KjgiJkLxcOnTjMb+4FELg1t9tE/GzFQAfaVU5eJ/EGS8nWKKeOuXWWS/cDP
xXQuWwOxAj+oPSx20JmlImrdkEXzdHh3zuf4bhryLIrdziEAuX2HFZB4/7RFBjkj
t9AnHXXy+IJ5T3aTOHUgJ1vcbfJP91hyJIH9YUK62e99yQ9c4hIclBAiifF9q/+j
ywcaflFdsUgCfLSIiOrMLIsj4W8SVu+o8coklw76xAYHUGlaEggo3ZQZ3zlcOqgh
kOQ1RfisBf0tkmbE8mfNBX6/Yytjq2bKl1GPl+oepQLZSsn6O91z546EugEnbS3p
FwM4OUbh/CaIAd8btEKmmAsqPTxbBAXjiin03gxORsHfHGeF7QEu+7IcuFpotBbY
QoASP3E+OzLtE9BXAKG+lfVLhPNFLzwkloorUZHVc4kfK1AhLJdi1TpsSyAfxKSQ
ZbAMqb0doVHcshHX+M2btsEDA75wKAowmQDJUfb2qrayEm6khjy48MYpYbdbzxQj
I3Fts8PKS/pspG1Jqit8sHSTwuej9YYyouCQBP/HGytNK0M03Yz231Rk8t7N0FgA
32yf1jmdQTelVW6FkTe9Aw9jzrGPc5NLetFcGM61KycBWeMf+1EpWGRm4KrAa1R1
ekjzSbZQdrCBTgFRl8FFRbFfff6FFpRckaXycS1l1gEv6y7D7w3+itp4DMlS1J5H
sEEfP3hsy2Uw+ALCRRu1s2cfHzlF9yvoiUcghNztvODABuwHACPVeWQefOrlCUle
nxikAZQLEMJuHROpwLfHeAFj5SF4s470j+krXACuiYwQ7OsQ/uN9WZtEkVGnEQZy
X4J/6gUOloKs62XEna46iRQZcQyvCEzmrYX9gEuVoNVtl2H0lB5+YEPCc/8OgRxu
jVnj8pE33+w/bPC27OlqQ6hvg/Vseo1CzjV6F1RQK4aTq7hLySBDsRszOwF+HEyK
ZowUDvufdJSFmngxxg+ir+f2N/9QnkOmIxm3xbkeWRGfj+lYZOVoSfuE5m0eF5j0
SgqZj5fhy5KbeXsp+QOtj+evfceZANU26jPHCQ29mzqtudTWf25FR5j5M+g7FIkK
HS6HAHMR/UUQ9eTnXPgVAKHZmGh29Tn3an2GZI3Zv/0S136Z2vfd4uAFgjVnX2JG
GmyxyAKSbrLjg9eV7toeRhiPwXr0dZG/zFsZHZGnFMF1d+kDOr4Mpaq7EV+EUKIk
xvzaZlubpGFj0WHDe1MOBnqTiOLZcK1MfQbUf1r3qlGy5nSF3wpH3MUZ8wPJMV1Y
lAV8DRvge7h+xTKLnXgcBXtSl+AixbURtJ702eAxhA64PpdYE/JDfOu0uEsbp0BH
wLIUC5tGZsuPOsDUypAVYR2tcqxcM8Wuj4cT8tbllF7NFJwOj7pmRSCf2QHDN8zl
fli3KXI6nitDNm2QSugC/JbHXuC+205RZxK8qM8igF5osfofMCKPVAbUtmIjcOx+
RknbTnw3pxcm4JA6gksUwCs3a9UiqfjPBGB+IHPndzevjEu6MuGPdm05kLTV0Kff
8iBVsLwmpfMmaC33Yhb107jQYaW/ZURwFAlASIJSepLgTcHzVL9XktTE9heg5ZKO
QoYDKK1ATj5QwPateYJQCv2lAXwHzOXWYKMx2CxyuLdoVdIb4G8s+b16mMWYPmAd
6qFla6xBHZG3b98AdWeOnt36ieUrxHHXa0wD8lYBTxGFZ63WjdwJxeehXFiqLX6z
8kc0Z+7LDpsUHOmFpSdHAIag83VtbcOx9zgtcF/EqoE8rQ+XxHh48/ckboGoo4iA
st3AacOoI83QEb+wZuPG9wYYrKHG/F6hUt5JyAA3Lc9oj2wFPq3uDXuuVip6+0GM
bB1VGWw4DWbq7NjI8XuWEsui5JplU6RTmccoJZOPMLQp1pzN7wrUI3VgZikFBjnS
Ss/b8ZsPmaJb+VeOqy0Q+DT7tZlIedixPCHveKHtoEg5Lr8KEDWjQoIy2uudsTKh
NBngKHj8h3vHtKthyxKjVUENtU5t5XsKnsQEEQABQaSLZzNLD6EjdQ3CiRxaKkAl
5Z/WJBhqziSlfAjhA6E4RYyiBXPdQd1k+F/r+XzC1GWUKD7zkLZfoRfoj7nGZoe7
iKpZqATwzZloBZeUkI27U1xD03iObc/cfMxXNIfTV43HQnKmmnoRYxxed3iHZhqH
HUwA6BMZOO4MKeKQMjb6ba8AQcs0MvoE0/ltZi09fDbAQvzlzCfpZEK8pj+GqoH6
/RVMEljMxDBSVaGWWy6jaEVbQ9FiQuKEQQN5x4iOAQb2eqpIlgToIx9KGdFOIEXG
mB01i8EG+EAG5sAxEBjZlPa8NnybNv51rN6AdzkbX4bCzDGW5SS6C4OqKUNrjRx6
pIaKfP13VK3f0sLkwFeYzbyOhuNKgMPaqXiBKAiDtQ72ajkOe0Mv3qNp0R9Myc8T
aOk77fD2qVgKtXLWzZ67wjRtAoAiL1Kp9CK61pggsWg2CpKOp2iTvZ3NVJAY89E/
bnuGnAETbOABR6YDbwKrREyXD6oXLJuJS4ig9eXKxfO53MM7XvwPtDNjbIZv6gPU
2s6AnOtqGPoIopvLOPuvOA8Ng4GDKSsxe3I4Fl51bPkQbmxUllqAJdvAOb75fHq8
x9D9r2pV7VS9Q8XpWBn1dhkW3OL40RC/N1EBQh/OdqtzVZt5N5y+q0DvgU08WJjp
rZC+6hGtv5ZDpukbHXGJiArJi9OtbzxpnuUtEWSVqJAfXkL5DO2Sb4UteAOvyMuA
GyHmrj0lSxeqFU1GgJIVXHWmt8s+0Kp/FIc5fYL3Wf1DsviXKBR0abW1sRnL/XxE
7nEPdpiCDKwkt4KWztBZSEs7R2h8sLdy7U6fN0FxdyjcNIcakKVCARMSiuzZgrcq
7cIbkv78Qov3XIXyxfGNuVZXjlNoh7wQHcTWZJcARq1QbH0sBzuR+epES1dERF6Z
qPEL4veuppmdtuzjE5eXuXyvsi5RNiQaCmfX5wkJ8xKSH8hz8bATufcsuQDrx9XT
K47Mfg6jrQUH51o2oW+VwGgVs3Qqc34R7QT2qa3jwVhtQk9AP9Q2JDUOr0BotQxM
NkBrctc9g2Pi2cLPfw2hImLnL+V7u6qEZCprqKBk3d6jan6gXFRnznqxqcOENCxm
sMxacO1OGf4sMMHyErjB4mjKRHMrDEnPXG/YoAtgMVW6k5veMxfiILh3JiZc9MDc
Jg7IdGpOvZCNaeVGSCkXPDbs7xFejZK1lQLYTW2gTL0ytN/229NVVkQsn9U3L6qi
2ZF4D2CweitxM5UQc6lB0m6z/66Ze+ymAe+iFIHTwPRIYcwfNL7iMAuScNcBn4M/
ASaTAibHR0vHRstdP6o/iVJg2HHzVux0kuSekfsUd+6RraghaXhkjQDQccPjrN+i
3+QT2ABvR7GTGZLFw1w7r5jjIic61dq+hir7w2QRZ4azixLLAMQq1x0lGlbuHyBs
j7bFVajokVWT4M5BFZgYEXpiak/DQxIRTlkBu6ZMYhJm5e7MhEYIXcEg/Mcwvmy6
p4dauGsepyEiYnIwiDbf1zNCM1yYZAekSZfQRcXHfY/GBeQiSzmxZpGAxVnh/FUl
jaovmdviIU+HHJP6ea3dDz05XwhQ/qb31JOYL32oN9maWqq93Zc1T6H7+9TxCdWP
no+bCzvi0iTYCDhgQYz9nlOt0Kh3+E359OMNQ7eIgbUWt4ruyXcbgPG6xOFhZ535
AJAgnRdOI0oHLJy30EY4n9piWoI1/xIH/4qgoWfSPIIy5qFUiErlc7fyvznyxA/2
pma/obGMoOTfdBwcJ5IdXNSKkeCXzcUEjoVVCP4IV8mahHuUB9so8hXlibmOsmSe
8qauMULKK2m8fPOy5u9ay++v6qOhh+8VsHg5sm4Rb1ukQYYzQa5sf/BhpVmOXpuz
RLr7CN6mgio87PF0rCA1szz2HO/o/Ah3UlLhjypj5XSLKm7IXux79DD+0nsfcMfL
gzxCivHuIZBJj/DfvcS6t9uMXThb3WCgQ24Kuby6O7OXQEj2YBv1p4Yai9yXS6EL
rYuNGPXxOjpbz6sPWGoRD9BBctypJxxzvEi3Q7LeChsMV2qPRcwxDmgwXzvqqhue
dvhO4apATxaqpBFXP0ioC8oOM1QxMneiNDQH1ZxTbH6TBCu/0IgKkNbxA+GOmjjI
9tKzcDHD1ad6+9pyJZFi8Ke7dVs0e1B8CLB/IU/iZwSeuuu4JtCasbPZKUkOFevh
9VO/CYszPAdS8ei57rBxdKuYH35r2rXlP2O/IBEQt4ZGOWYeXOqz9raJhLN3oaD7
kCtUgs4uw9EmQ+lENV9lB2xdX45ZDrz4ekSmoEOg3sggUTSwU2OSkqo1ylPmlflP
Phybf+7XjybIszITVSsUQ2BWXIpcnei12+OIl6vvrIN0F1PCg03gCWOu4/2SOLu3
2W2ZuXpmRg8Vt3m66waotF2QidfQ6YswxaOxoyNHtboQOGmWc7ClJw5psk/6mV+X
fszt4nY1nKMAJ9kuaKLjdwAV/WdVal56j3Ho9DkCqMDugeR/d4JLijMvmZOGSlBZ
bNY6q3Zm51CLOSImDmF1lGj3fk251Dl7X7G02cT0Mlp3T55xw3Miv/p4dCpjIBLn
gXLOnd6Ocy41S8xtWJQfUC0prFWlN7+zxdjI4XHMayQ+xL5p1su0NKaVzWBXOFrv
qz6mUoWtY1LhM3sBnGtpMPYnQawK1fMBOONDruILLlg1KOrrmbJuMKIA//pRCr9+
AgkE8oI9uQ8CEdkMG4crIIEpkNoHvb7VmsVtHG1S34XR1CuSWTaiPebzRRfpp2V2
76s29u7QMVbnbyGgkaripx7KwuMb2zWihkM+m8mBxzPmt1Izjm+slEcWwrAYRFn1
nw/gbJkbUoNIZAm43SAZMalBoRHW9rpJIGje+cvhVg/yFdqO9zJhU1Jq3Xcr2t9E
xH9hxq9Kjh1MA84QBRnj8wortDn/bAhSy4qnveqZSYq9/LB3vTUp49GnQyxTuREA
x9EpMLJj1rGac+XYsS800V80wuZ87L3jTZSO+7Ml5N0CS/Vxl6cqeV9+Zqr1hfVR
r73MXdoPatGVz086a+CrW4E27ObivCcmskWrrwuOUQ0ARnINBBwpHj//da7yE7ZR
7x/1xkyGmvXsH+2O0QRUPm6dg0bM3xJenvQT/cKhEk9vqY4rXyUqbxuQ3cLIGh1W
2x+XiPPhGyqVw7RqI4nlrV6shyceKlw7EXQAR7pGR2CYizMY2d2f3/+ajp7Lh1Ht
mrINS7E7sqXz5ipe/DP0Pp6jjOjvxake4IDxpNba7Rl3EBzfsDHkuOgUiEKmRMbH
Im1dTnPOuS8VP23fheVqqNyPMns2rmeUvihi1oAdDCR9TU5Uu/E3wxOgJ0WrmLTa
IBAIXzbBTYvhK1JWo+W5Q2MePZ/JZQ6FAA+JLAhLqjxdlUSTs7+njrfWr3rzUcT4
km04Docqv6W08Pr6i7iKkrwWCP+Ar12vWaiWfXWPaRrosxPCp3NYWtUpDRICseyT
0TA3sSXEwpJlU/xysqy6eqyaU8NfBuMGNLSarYyy2vVmJLLIuIrhQclAblDLY5Px
G1N2zgU5VxNbhhm2E0HRMoM++fAkhtE/TNZx7d6Q/DrFRdDvgCXEqxdohuK1ObR0
jkJorRnVBZRHvEvki+7fY4VjhHA3r/jb57S0+lws1NksmcM6rSWXxSLKCncw0QYP
V0jvXDkRBd9Ao9kX6xNAnBSjmQjj3OAOY5bS2YLul4966JH3hv0Na9lIlis7+Alr
jW1U19VhFMIl6xJERoDOjV/zDJKxJ4r8vVOqElqa3tjIHw3lAqaW+VnBKeh0us0k
3reaoWWoBKrPh42HYmp86maeUyft7qaRzxX9EzC5JlA992CWYyZS7ozMWufY89t/
twmUze2u7BFKJYIKP5Zt9+lFRV8PFzfiNMT7DIQuvFIc9+6EGxKIS1LMoy6i21MS
3Oe14vvil8tMWGpYzIBWzYoXmfkyvGJUqIO9ocaSV6rrt2q6NUb4et965TlQrtbg
pbgi+JKWwplYMhKJFJw85OLYMVfA2KphCERSVBvfnzpvrbs7T8aSnLdITMER8PpP
M9u3A0cYCVUaGa3wsrG6xtJx1iqwm78XhVXAp0iq6Yc+D0Ixn/MWKLXxNtN8osN5
PhXYhBmWSukigkUbaP5gflC3nQ7JYnTPJ/Wyb33SIGAoGZFb8FspKWqcpeNBnsY5
IVrM8lMi0YzLPHZxJrSTFCPOFQU0EXc13oWMevxFte/QVsWT88X7oc/CB+ASFqNp
+P0g0QUY4X3KmHCfyohCrvcQE6k7oNHROg+wR79OE6jox0ZkvQrCE9/FZOjf+JHM
UjreT0W6ENcTIJmm0VD6VQ4BuqZ4Om48zQ1IgHDCto7C4dVqTzyOmr3gMXrEqYTs
GgWwX2/nm9xja2FA1FM3gSPkGUcTHDJ1Mn11TUGHSlcAkzEtm/FhsGSppPVvYrxK
JLr4/shvgs8NM/u+QsS74oeLFDdxkYGe2UkrgQtHVQNiJfdxcK3+FJP7ux1bK7c/
EZLJK/2yoHYSoTmxiMSQWvGg37i3ummnXNxC+lX/1RUHmayvTYiqvzFX+iqhhCnO
kOcdXG4FoQOFjfDei7W//4HKlw+tyQ6lKMG1QNEYPdhQ5vtuadENeT90fIesj6um
m3MlfduoURGFRqUl9Pj1exa9QQCqWJM1elATF4l2/p73PYqkcGDOja5Rxxtkuefh
BCM4gaNJDJQLqzpYuNuG/cZ9Xd2rypD1WAAj/6d4SPoydhftF8TdaOKjY1ILMBMF
hnufABoYLwX++bGKQXeARgMqGbBAW9phclYZsGffW+uHvhNiGeXT6/kDRjD9hclp
WxZVC+E57d4AcikuEFtBV7kcHJk+ChS5BKx4en//qLX/kCoyGT6fEYG2wOdYUCPw
a+MEWA9f1VetdgHjrWbTYvF2C+o81QVf1GGu7uAwOkLa+li++PEOUfxHRRbFEvne
c6XWxjME+YomR2M0vfMCmQASMqS5b7FxAwwlVC6qOSls1buM9TZtcIWdEHajrXw9
1UvdrjCBhLBcwCrzltBztANZ8sM86K7VIJOSeBs/Hyo6Ia69A3awGDhOsdVX0nIm
5jnYH4o6pK6fSJuR2EFq+Xblq3r6VFbmTu5wamciE/WoAQ3NVZXEZysRMjTev6iz
sxqPHZvRr7Q1Z3bf10Cck/pX6ItjL6NWkWo1iSlg1q8aZRPlIiMGZBWywvY/qydC
vx9AQUDHe944U4V/QMpbQMuFJVZ7GjERuIiiDOQLaeIpS4A1LD4rCpZDCYN/tD1M
QZpPzbqw2oxHAB2ihw0RKm+JYaUvvf8cni0bNLdo6FD2b4z6jYu0J/HxUqKtlksh
/jV+7hoGzXu/WEeFeO+IZ1NpFANuAnwdS1agxX0Ed6XeRuX+Kis6cDkfXR5kDJlE
CkN9kfRiCbAKh7Nw2fkKs/v1gT/rFFLyS9JnBUYFJlRuOuToJZ42rJMVCyIfwTvr
gpz2THLRAnGdZOA51dJUpmJoA2aUHbKu6mMpxBN7e39ZKe3LN9KhIh0MCFGwsccU
7UddgyAjtvvd5pcJZWof5+kqAI+JE5knu7u0DQNj1F9wjqzBazDfC2xGnz65n6Ff
KeSvPESJmtvlW3hjsu0ljD6nSd8aBJz6C+JGAmCqg3c3QyclWjAiF2I2pGbVzEbd
zaksrziSMgCk3lngh5alJ1/ptLdzTTLUxlGLnWgVnLnZjHc7u//GaBlx556mcx1U
D2iUN3Qww1STudaFDdZ4EKpVlyljxJx53oI1iJ3eQYlrPpNaKSkpcyoNPIKJtSdH
7iXiN/DxP4q3jGsCHk460AkEUYyB8octqqb8gRkphpU56i7qIUdyzxT08IAyu+iP
y+e2YrKIToSYCgG48xFgMsJrObmXh2j9xWtJrRPaz7atWQiGkObYRsiVa5iRj6uQ
JPwS76JcLdJffC37gt779hIgJ1uEzoqqqJZmKZGh4lmrekGTrqnLQrlL7OG5y1yn
wD5gw72WfYJy6TjzVZi5va33OgtkZf9Y0XoF8j3Qx0gRU9jt5HLzJhxRDO65mjWA
mLqmryK8Dr6hL7L0Rm84l9o3kSD3iax1rfzekazTX7ewPoFCx7KWKV3RMnYbjDSz
iVqZKCqVIUvm1VhZTPBfS7dsUKW0R/dfpBXPmmNFtVt+LiP1A+rNH1Ok4deeaL49
zulBTzEYOrPnVTM8NmHB0LWhRIwmKYX68Ds2u2HnOfN9cesZ/BeIh/tY/pPzIy42
33jhe4dtstyQi1lbpH7XQKE7T7oUdRXGPl3HNL1PIE8ho1cBBupWIkvsd/G9xeM+
k42uArwUuiB4TkNLX8wGnN3V5FJAzpHqNs6l/fMkBaFclJwp1l26D+alu0PREaUm
9rgJMHhUvQZfokFphhB8hrlr9g0jc5iHhIAPRQbNTqpL1hXb4U+/YX/Uvv1gNbZx
Ce9ke0Q8NeptADR6AX0L3dRC3oCb2MbtEkhiJU1o8LtJ16ajLXogbzSoXpqClaNT
10Aszz4sWMWM6R/veAmUfm0iohn6sgyZjroQhtUP5BNopud9EWxKfP4/a3VKGn9a
Oc6uedMfIVkcwDY/0+P7lasDIDUoZWGhTBPh388x/YEUXCzK27RyFYdYXYbKv9WA
MG4qTIIqmDIqTIafPdrfSJtSs1yJ3tvEuj8iw/k8GbhpQFcl+CdTtADQoTSVkA6M
Ute6OBknoKjN9wED8jb7tetCbPTVYT1KAF7dvWyMIImV9lMC+RAD8OTdeNt7K4jd
QVnhWDGOOPrHL5Mu5JxXBARkRTdkrabNhYA2QMnHeGIiNRcHsNgJUXLZ62o725KR
zZXB8HgZXqr+6gF4cPajMhOD66uKnWAhtNnN9jlHBhllzASGZtLW08aBFGkjQHxt
waqBUK7p0dg8qMRAhdfbGfMzL8EcJ247AlQkFNubHz1k5rQjqm3e4ixXbV/2cdmz
zXhtEnGBarZvzuJEzil03LWBwQmtEEJGDCauVIRrNcwV/UjVHVl2JdS8p2WuhnrN
qWUG12d/AKlQU6hby6BmDAF3DE8XhBtJe8EYJjCWFeIWH1Oy/JLGK7v9QQDWnAKN
fSky8UKxtqzl+sKrICCe/FC+ev7UiNrS1eW4UTa3+ogsKtnBHhc5kE7I16es6kJH
RsNcwlVWAblYjjYUg7PiuRHy4QTPao0h3p4z7Lm8MPPEJfNGdeAwZdvhqw2pDZX7
439AKNX/P3ZPPTAFAhvvhToflf3CMnN0/MPUZXVR/Lgmgn/MbJMldKnjJYRxiM2N
loY1MA1/NW7FCROp7M4c2vvhTwA9W8epF/SZXlZtDLx2az/JXDgZfxJVDGFcXguq
5tZ0oQIlQo0pTEIeaqgNoVNjGJWavYWO3PcD99WHEyUletKc2r3oSasc6xgenImN
q6iH6pN9OLr0al611fo3HgHaHkeCqW3rsUCwwDaFK7XO4LAc+sGNtUIFBDmQIZuy
hvwvdisNfGiHaubpsaVwgmCgdX0xkTNbX1dINZM2AwV2PQJv/IW4JiHLVYeWc2MJ
+fT1wOke5BkvYGGPA5WXn6W+++vYDkby8BtuvSIHukYb8ky7aDhZMmaWnaIsilNK
AQmzyOjNkHF+j5+jtCo7vipAq8aX26VYwJi+Xfbcwz2ekJot9tv7oU8uj/k0fH0c
U8gJtrK4VR29BJ3IZ4cvquw9N/CvdjPjeE36ivNt+zPV5Wn/fKBa+PJU5XbxR78O
znmE4QfyVhLMKCXYyOpk9aCubZhFDG03FShGa4Wx0dvXJ7d3TFUnyF0Jh3xSdaHQ
D0ap5PhKUY4JEf43iq/f06/Drs22pGtVV+jWUMYzqqPyExybftrvkWbi0nt1j+k3
1NRP8yNDqxjyMVNxvCgWBw3ztfCDZZMem/7As3/fxO7ujtX75ZaXo3BxcLvVbLQT
ccidtnc9AGInuXwog+UPzLJyZRXhLOfgPxpA+fJD8v1YcrnJTkEIOF3wT7WWRBJU
vIcEE/LU0mEsv1lYpGrU55F3czVRPMTRHWdCW3JmbwMcO23Xufe349pobeBwp/ji
1urb9Rc4+q7feJE7IhYStfLAr7DPVBu48EFirG5byUFhIaz3GAgUnQ1a684PbGsD
qHUCDGrvTeeotqdxFtdmZh8z8xaKXqFXyk9YOT/shaGuzhQxFUq1nlH+tPkRNwfk
aul+TdIGHu2BDajFIhWhcPmZMIIw5y5y8dPgCVhiiQNG+eHnR05JS6y/sI6PaNLn
/nwnWXWMSEhDdtcqdx6WTF3WPIw3XWpBjSY+oacSBX+CzWHyzA+Go6zj7jgxvS35
QfPKuYveSVmyvG90oInTqzV8MlOuMnTwyfzlACbaJBoDhjh4ycS27qZNazF7t+Ld
5h/S/orjmDnVtd5j36ImJ6hE9YL8evLyS0cNZhEtYs1SiphguovBHaMjQ3Wp8Bkn
pK9VK9915wYbHuZKuCWwpF/6V6mO3Y8oQatGU5GV2OQnlv/LpwCarw3PaG9zqsrw
6A6HuciLEASpjuHyM5I3tj4SCqSbS9aTNs1FS4jcNBzGxGCxE2ktcGMp16HsAtA9
W7TjBjbF7TSWJ5eOjqsjm900RNRvzhz6x2z4O1siUdSmCXOWOFzAv6kNR1Uq9sNC
O7bHmQRfoot/52VNOxVU8vhvoFadZpF2G89v6Vn+UH3HBMBcmvFose+4z0Wbbd8i
UluFkwMNAp/AG2TYheBlFF7k6hw1Y8+q9XuyKXqfG94EusyW6EuOpcgF3pRvfYga
QAQS2gFefxxR4zWdlyodd5ChVdlKbHy/luLPDcqDpHnfMfWR0xJROOOrvQTAU4vA
3CYC1o4apTbj7icL2emxcRPV4aaEf4259uRyRp2x8+AT650zoAoyEsvMKmdRN5bL
ieejGLfS2ndnauOglO7DksqQs/3Ty2gQSiLwteAfAOv1zl5uH63EniEmNgp+bmGA
l8lUxvzN4+sb7ZzG5BqXrrRFKyIAEMzcfidO2C5cCuqfxc42ryjfHSx10i2Tm85P
rmv0AHNRNqSAerAjFUU4r9I2xjt6KqVooIof9cmoyTaAPDMFj4vqI86olj0KIzGq
h8i9KUKTmvUjvMznJzrzEuCib56mVCfGkjY/6UV/qEjvdoKp+n9xHtiD362tRemg
i1q1QkdVYmUyCldlJIU9LK88n7idXX1E8JiMXB+mu70blsfaH93tG60TBZdz8M33
Y17B3o9wrma22cCP3Pcon76PsDbvmO6xP1qk2fHUdlrMCIc/ECk8jmICAgieXJxu
16di70oOMjuQIVNP6IsKgbCVk3Qndea7+py4xUF3cVI+aqrmzT6oKJ9EIkhG3HQu
71BB213oyGaUX8gZQooYQM+3LgH7gKwEv5c7pRRrz9/QqrIa1XzZqx4ELdlUFnOT
7ATZAccs5euu3ULq+tfeytWyC4XZf1+TltCsQTluXsC/FZX3+J6PRk8A2/aS47Qs
3lUpaAvUfUvUtnmMgNn2CnL8LjXTwXv6jwFjDA7hH10uvAy0aXQtJazMDkwfedkb
YG4LGGdvBfDXiZl0LBw5PoLf3JpbwolL6xNLg/pIC0BsUdyOe9fwsoAPiXTvmOpk
dBWhwg7m2xJDezynTPp/JbTVQtntg6jEGfUap5tLKjBJdmNu/EMCWR2knNzYtkP2
N7NZ5p/OD9fFVZhUG9BN3VzP+DvwkHZOrQxVMnomU3jnAnVqPS/VsRkxnBa2v50s
3fGqJBFY9vDlKPWh9hsiilyaVA06/82Z+/E0bf3LBV9lSRZJi8wRq5wCAfCvAiWY
nGTKgin1TdCqC4CdSQOKmuHIguKMmX5eC0FLsC8lCMAmiSrA4J+9qUSKu7faTyJp
tBVXSsxAD0EVOCDREEr2C+HrRYsOmulo2ryocye1Pf3T0ZqBvD2nfvyFWMNsk5eh
oFdzR6bBQ9baOi20JHYEB151fHlmxXOB08m/tp6kLUqo1xn5DMLLI1NCHTM//Zez
1LIq9Ob+buj5bEXWvNx+prl/95jfEu5Eu4Vl53tTYWfet2V37uAE4SgS3zyNbH3S
tene/hk8GtGo67D8QuQS2uLnXZibtkKC10kBuzbQ3Tg5q1sGlkIBZFopZAhRG4PK
h3HTafK5frhCM9+TOEHiFyo+CyYhse713A1n0L4FpknVb+H/+UOZfyRpebRTrhkU
OSGGbg1NYPJikmW+z2Vkbo98hj6+gxwXvbm3vJwOJbLGxwe1FAyUqWMGRYwFvLO/
DFNV13btT2V5xMAofSoIX1kYGsg7I2Bo7/Z7VAoHlOJ2a/RVwcN/r5U8NZFAmTkJ
uOvhghSgmN7uvfrgzOUoB2aIq4kERZumZTxj9rAQd2/bRCm6TN36/W6O+nDkIBBX
HPSEv6qqrZN5mXHDYqbJ5liL9AB+rMRpZA2lWtsbj497bg/MonFgjFAq08plIkQ0
Ggt2l9KKP8PJDsdBlU115xxFK8EBerRUSj9zARGQCUeyqIsI4Amo6a+ywo6z8ZPE
Au6HOyp7A6+EDuwzt7XtV0K8G4y6hQ4MWGi+uZ3mm8IxKnTjcg8h6RS7pX0XKI12
43LyJpGj8V/dZClR9y2KUH/f4pV7wYYFc+rDRjWhvgYub5lMK2hfl48R7rKLlS/E
/YWLakOz4LGbKhq5Fk84ZwcwU/VLpcIJprPb42R+d5vmGNHzpm8ZQQaY/cScAmUg
ejiQJUseqOew3v8qpkyIxQUSinxX2wI+hEp0zwJyVzIBUaOfFLBTBdYDaq6NKcOb
s1wh4wjsSKpcK/3voZoy019FdmJVy0iMLRsmKRMODZ7xZlLsZj/zokoNRPMUQx6k
IOol1lw6rlH/rO7e89ZGFbhgntd4Tam34Qk8reoesb8l7M+boeDDFSZSvSenU+20
JPeZSWIlbLs1DHFqp3sSvZjygWWHUrPdVlBku+hmaAfW7drs92lezrMBr1x7KuGz
ygSSamaR+4LY5rhBGFq56JDgvICm0wDjPedmEofntXS9uDoJyqGAStJuMeJWif/l
IMDk/GAte9c0nRtHA7psAPom4ADN/UYsYISMKB9hxTV5Q5Ke6etyqpJZqRJO64mM
0BQZk+XYC+C34Y0rRmV6Vhhl1uuXr3tWaAojxnPOXHkmaRwli4ae3I7F5PBghH6l
Z9YN/1eQ0IKnGIQtz4SV7W4GzScYeVZarJfCwdvDlpRr7yibu7YL4zJhbHo7kdNh
QCmqqv6NEe/NaK7hehcAMxcgo/ZXUldm+U67Ei+14YkpfdyDHOghnxTRLslwn+Uc
kDcqM6QQ9C2dVlDdMnm2xRdX4Z5qlNkI8Xfww3PUKFtQedR/V3Tah3zw/7NBGc+X
rq1hGiyPk9CKzrOf7oWTDF+X1yL6RH04Wzb6JvnRU9ciLUbleYyIjBz10FsLrv2e
ayYv6m7UuJ1ofcCbNZFVYv7RcBo8x6kZh31OcUA/g3YRZCdEBB5IBTs5BafBfRw5
mcSPKV+YgYAhLCVTJKZ9K9gvc0GT6nLvG9/5z2gICFLg7gMhhD60Is2dq3g+J8Jy
YO25vH3ioHl5ybcsSZ+5MJPM0D2GRmDevoI82H9saKHHZPN/2ruaQJVRe67PNvCy
VtEpsh2lPrUKJb/3A5Orog/3dCTcnf3ppBaiSMC4RhGnkIp2x56FXthS7GgKsTmC
sAgAzkMbAQKMR69lChq8XmhRypEO4ayR7N/SXbbr/dwjqOXZXyVl1HUXxuVgGCi+
/iutwPPcpGq6vMvvJ30BOwjUFGtd+QxeCSL2nBjIzr8O10UroA49k/+npd0hoZn7
w/DW2JD/Xg644bwIG/C+p/+IsC0Z3Bujjq+wpQgIDuD1FmLos07jnPGuqWmSGDAI
qhg6XkeeILg0tNynKwvzORAY54Wl+Im2ZyPzyUpGFh/w51bBBz5Y7jAbyxf2Rm4D
Y1u5mH8o4YywQFOTyCSA39PdpRbiPw1n35+9lS5QF7ua9uSeje4ql4Wdi0MzgSmk
hwS0xIu+e7FxzjxwNUouC2RJ3gNrD1037Co52jifONYTjQm4R0HVGfhEkXykjI87
oPYKgitYONJKuh2UzXBvOTPzJ6uh7lZaKygKw0TQojZpx4vHKcoavJO2pD0R3xJs
pRxwCEtg3OW7HfybXtJmAbpOMWNjTOHiEfq6pgGrvqswPuFXXVkaK9l4dyA4bA1R
aTTfTycuA8WpiNWm44Aww7LN8xh37FzDp/q/YJj+4/PwVErF5r7fzupSKltH4O2r
6gX3b0Hu+E1bAkV0FZ4Uwpe10FSf+1lnxBlr3QCiXPhtsIs52hnORYtLYL1WTcWH
eIa8rIZjkMSDEyWSd8T9WeMBYsVzeIwGJi/Q2oQ/0K+Iq5OhpmXBuccQ4CORdu/Y
26gEK3Rjv93I3N8ZpmKQn5sDq9gz7uygNfhxvwtTXqTcTggnoKgUFoix+HLtrnhE
otxQ4VRPwOvvPCvfc5L6DlJx+X4jEKw5nqPkdghkJaymb//xlOGkWg6VxPpAe9n/
FgnMvinx7vpeED6K2j2D3kIr6QA5HBcOZGqdoMJizDGVWMFvj7oPQrGzMoeOnVIm
Yu+W7okof1emNxI5Bjb/Fi60hU6qk8+d6PqFIJvvkubRAtKtwRStzV8iKa8D2uGL
olJ6kbvviqpWqeH2XQWDfDVtemezO+Gcz7H9dfiggG9Rxp+/hm5pLOBq1LoV8xdF
DQAXVLQ0dwy7Nq1icaGj+vLTGZgqeQdMN7RntRtYUCf5eIfrg+xGFvN5cHsr/6et
+5GUp94GnQJwfiAArEoMS5goKXF4zxXmclqEA6e9ux6KUwjzEKZUDZv2cBqHqeUP
jJNCNiV71pgzWG7ssvdjV3BSwxqS8OkuEvQTpL+8T4T4J1V5DaC+zN5Jy7LZ/6Fv
LBEavyZpWsjv9mx0nyWxFuCb+13oj7IP1FEPkqvVXX2rch5ggBSQVr1ZVb9Da3LP
r3Ba/bGBtEq7TzgAyO5BNxpXZW625Ff3X1Bhs7Ea5ahyqvW4WXhxiNWMmV8mBWsp
ctCrHWw9nx0RdRYFnM11PKq+1EAkTAEp0vef661Ayk7NRAkXbGQ77iIwhmfnrEtp
vU+CVR9Nv0YFAAVlST1ntLESPyTzITbp9Tl8h2i3xQwyVL0Uii22Wgv8cB19shtH
30fIvbRj1t/ISeiQyEgJc0EBKKZ6J3h/QItjfYEPvtAbC56QebteGnCMoOyKEFkV
/iel5RDV+KIUuEr+2u5h4NrFzjl2QXZtALsf7TenkOMJUoTB5pUXn2F+WlB9i1Kd
UHVvodzMgSGcS51wxQKwTdxcBb9G+kcLArjYl5gA8xcEuu3gXIYBWbeI2Lu9V/gI
/AOw1/jn2wUYhQfGAKHyNas1GaJUrLoTpe4+LaqAZjtJoNxKoZ88Q3gJQTHA6XwL
BbwpM5ex/ZZsFSQYVo27Tl5tFkBzdPeg0QLNdGMNrowbPgFs8CzzTcJpjZ5bm201
hCjCM5eAurs0FOEB+0/J7pMrpIQYWHZaPp9h8JqhNLxqy5cMSenQxAtrzJyT2qgV
e/t4zbG9MH/OslbaXUbkNLx92C35o7vWL1MdXOWZ3QkY554aW77bXJU3GgxVbMbz
yyuvvkZJoMGMRyEhYTAlSZmCw8O+NiyMdjSkE5d0diVQAPWvfNRvk3tiUUI30lxF
ClBC8LysTxzJKYtqBBmFrJt8yz8ArwR2y1Wc0FooXC8oDPQn33UwhehKz3HKqC2P
HbnOAHOEQfKA8CUyckvlCXSut0Z+lx+zyRHiUTX6ys2aS8fIlQhpcr7PDljXo/eQ
UC3VkpRFvnVdudkkCbLxy+XWur1qFIDE8H4jPG+lfz48yxdiq+Zz92Nrj+86+/O6
0ZfpQcgHneAqWinEJVYnOZGGiDYAloQwvsLO6s1oL24cZe7X+Y9luz+YZFh0iymE
hCTtRVm3DOu3FZCzKUo5DzhjHXNiAXaUmnvAxTgxHDk6UUnsVRo31kTW7+XMF6xF
QI1EtZXEdhhKanRUTXIs3ijg9zMc5WMOwr9LvJcG9itWYPZ4atHhwqGBI49HCs8+
Fpc6IiSh9VPqkYt6HrGqH+8mWEl/6Ui4/CnRe1p/1UtVlrLoqZ0rtrnWMvepf2T7
d/lyZWcu+bDYE5NStiY/S1bt0TbWfnt5JTQXevycKBumn/t2GpqUdMCSCbOuj8AB
UCEgjjJxrkD8pBKKM3Fyq9F47q+4rIvhA/fYG+aXjErqO6z3buS751xCiQ3sVPKy
+XglM8PfkNd785oSokH1A0fzWCcrMOfUuMbdDMVB8ovzW+qnqjbJ2ZXb+fIa5DsQ
X+NEmHwpNNsZeTLoRa966FXYWhXJAhmiMM+Ak+/ortwo4G0D3gNnD8o6k+1U0TQ1
rWE00XbQdmbdQy5Iu4GFnSdNXzRah+hvaGNLRYZ2XK1ibE1RkB+SgiptjJJrfpIO
9QQgg/gnmAl745ubSrtiErheKt8fkKLCgKBcpj7cz6WE0DtORJyQwAxtZE7Fosmq
JHaTZDUbZ/+G1E/Z/PZ6wHZg1dNdELSigu5y9JYjj6p9piEkxXmh82ekY3sXNPHG
2PQZWf4xpqILcZ6xEEg86p08KQmn/Stc13WG99rhY7sopMMDCxf2zYplpqy2G2Fl
M671NndbQnGgOecXOabPqioAFZfkLuaVriqSmcCR6b3opTzE/5ulPhdLPGEMsR2V
MyciCpsOiYdR9DXVxIPv0PNoF2/9t52cEp1kRGRA/zwWRzA3vjLrcOlpR0tQtqds
CngMflN9QDGw2XY8MP1qsn/NjEk6UXkN+u8PI3xzoB9LXsL1vlMvFpmhx7z9WMQX
IeUzVnAepHiq5sK/q8wqkQxHNVmFskRLN7E15lJWjC2LdnRO7QdBCGaJ1TXK/76+
HaizIyAk97fdATnWH2xdNKgf9THVtE59Wo+cR4+U+OwQkc1wxRsjkhlr6KAWMymh
fg4r+GTgYb8SbqUHgvsL76opu2kXUmsB2m9qtDXDqxOhA20FfauPYsMdhfaXxGmS
SJmWN7lSp2QucFfg4PU1TQzmVRkNvhLTK2qvIZwI8qg6B8WMAIrW3NR0c054zXYA
qdZE8jraMJ6GJJZPaF/ie6DQ6n5uuDPrvpvaYDgANaYhx12Y/vnJD69eGqAY97/j
BxwpJYfa+zexd+dnqslwlwyeh2KrobJ3lm9emthoJvmWiDxDWQF/W9jmetzeHHKJ
ADP+phNlYar4gk+bzWRxd6l/JBOoo+2YEmHbv5R5oifxQKeTgKw66neco4C95No8
kenoUrNWZdHnj9UbTT0A9TqcFzsq+MMUPdsKD3tARoTslJna4qdlF2h/duqYFIIs
5YGBP3S+Zki6Yk8M4stI8xV23j7yMFPoR9WN3JOU00NEoY+g/DN4WA+cNCTtFewC
Jpc3ddlYFMYaIXSMEagNynHA2ZuCLSff906ZrcJihL4+i1AWb3flyS9Qu0y+UsqQ
FF1p8rF2Zm36PzoNvwH5thyuYiga8jZl09hLFPc+3S6KZ8AV9864dHsxweFYHqqS
nN75iSEozSmEmlv0h9w0RN2GBiq5CC/eO3RAY2FkeyHYWZycX4vOYMs2CmQgGDUR
n7HFLbnaVMjKp0qqM6QWVkyqdRA35jjQ8Eeu0lVO/FMgUpucEEPhgadTq+nK6TKp
2TWJIQnDpVDd/Z8q4k2QtZpNJnndK3soki9lGnpCpQZNmCGVHoJdrLLs9KaElhL3
qpCRrqxTcydHfqpU/T6ntzZXDzihfYrPmzbwTzrOH3oaqH0c6ZQWgJQEZET00zTi
0FDZrpx7Xpr45NemPg05ZkeKz7SGijIFQgdurKCy709TkLiLXBuw6hg0LskvLLrb
5dhVE6h3j0Pk+rzYuJxKEryYOU1M987DvfTzb0j6Q/4Ife+YJUto20X4Sv6NDxpL
VV6IQsl2xLXfvuBFubw7qiDqOtHCoBC3NHseItQS2VaXtYeY47R615kRpKCZeJi3
WsRzppihpHsmUVxeQHGxOQqR8CVQUt7Taeibx5gYNZNu1QGT3ztoaln0wmvs1CR0
yzcB20ghxGJ9aAx33d01yy/SzHyI793nBhpoJ+LmoFMBOzlubEx+BmshXJH0S/bU
TKpGJ6sAtsryY4SCjKIvdxvmzo7xI4hbrytwYKK+gdQuz3vbNx3LjaP+cb58aiGa
aD1ZFG74amVxmo/WUFEZNYJFvnlZ6tO+1JPkXSV+cSreUGVgUDbjkCyfA0O4f/cu
1yHdcrcZCQrc75JnVh86SwnIm6GGDUs0LnE77KpltcS7he4K0lZZ4lQWFzzto26Y
VUllvCsjdHqMCoCh3m8GGYhR/hA5Xwvpkqibvsa4NZI6OFZLzoLj/lHRl9JTs76W
E5Orm3Sg1/O3kLumDpOzf1bJFvBXoXzn9gMg8aOMz7TWVcsBAr1sJtZseWN39ovj
lNhrUNdHDX0ZnrgTWjVHKx7Z/lXFI3tJIUxwUQ9sar8drCYSwuubOE3hzO6BA3TJ
2DkxnRGr+9FA5xzjQxy6F+eSEzTQzNumFrwxsSuQHfx1vnXmxrFsgP5tv4QIBiO+
IZYVfzUM7DIzY0LfdKtafD+hQtQhs7bz6gRO3hKtfxRu4Mu6KPSWsQsS+cjHoyuZ
CZXrBD0DV3e8eR+YSyH4cIzP/Gsl3/nAtFwZcPKYtFkURuxqR8vb5BZP7WXB6qul
mG+oJWVWORpUogmoRwYuh+Eqhg/6qUPegC9EXDlPvncjVQH8IpASRYL+aYcL7J4R
oBspcNZIpDBq6VnGJKc6cPaEEL3KZOeqhfYWdkZTXF3Z10j0V2uklWS92NWvTKCB
IB3Z4cZbs60vIIYOw+zuZUJUERfDf38XoB/2JLVi/AyAaEirRwkYxxZHu5o2YCER
U8ROEMWb3nAN+EvOSAwbqmbeE9DkfaGJVGBskSRFdgwz4SwGV01sgRoyYcaEwibt
5dLZVAOTwGLzC3dl9AmS/Q2KWKrNya7bEgCQ4ly/Ix6oQypzsUVY90yHb9f3SQYf
Hzu3vJ+ufD52clHaraLft7P2LThTOU1yxbGdIRd7ngfmTQJjGqxgH26mfBUNH8Ei
mx82Yq/fzSIg1oWM86BUjNty2ULpQpsFGJqF56iBrP0AdbKsteu5DN03+cqy8TvJ
dN7oEAeTzRjQPGBkmUbijOXaL1Um0VlQTnwEDzjyZ0GsClyQ/RN17XBzlI+U/HR2
g0/0vfVLyNK3fKEXp/vRPldU1W9oKRDtNvqajTT8afkJ/eNvKUDi7PYDYuOX7zjB
Bh8M0RaohNd9v2kYL7Qp+oWvXKI7tOZZSRKu4fhuFgCaeRswvQSk8xhQt1M00AxC
jDxlZHbyB+cJtBKMHmaz8Gn0C6SYu2+uCDMLPoXOz1NQU3ZYJrH6QbB4goKlRgqE
EmT/cfCUQ1tSso6gaZQKXqDqd4F6BL8/F4hc0o/kME4KSI3DD7t7WtsES9zbUt/J
nVcunmQWAKYYbrIqmAk9nkhFzYw4uuwtdQSoVCPror82GiUguGvkSUolemW/RkfI
G6XBZMGpUqG3gVi8CHh80UJ5Y4BMgHqLKnamBPmmME121eX7kjNuEtmvX3vcGRlH
v8ukDQK/ANE0BmxP/qFSrOzbuSI1JPnPc5oJft4rX1duT6xwvx1zsEOaLTWG08NS
N0KiPmBZ/vP7xdOVXKh9I4Wl/SZYqvvnV2TfkQ9OwmxSerJskaIMQC9T4BZNRwiF
ECAIobMPiVz1zpkxbuevOSm6JtLcFRCdxXVt15ueAJ30nKsIdBJKOP1ShOOpe4yG
QcrfnZBlHEacKwtgD+D8rLVcEZ4x2UwlPOzVxsH/8CLFObvgIDo+fwZ/xMjx+Ag8
HECqYqc02hWuGfXbgrx9wNheJPD481HALSt9izofCxzrKUdkVY8ymOc2QHp5xUFt
cNpGGXt4AbXvNUtnp2KpoBhZUyQoNenxv9yeYx1JgO0fKrl5yHT4bkge1vNCoCFP
vAONXdXpJDz6rhhR59Fl6LgJKlAnC7n78rLqBJuJV/6ouVh1ZjquPNHd6fViCNvI
dzVLzoLTtKotE5fb3xQzP9J6nBDCcw7zVYpITix7CSJT1A+x6aSlLDFXoHGe5WHv
Tc9FdiQNbDacBzpUzGe4j3mgYITv8/Jkfra7yBf0sNvZq8IbGXqULU6zLEqwhy8u
pCrRjq3mJqLg7Yz8lSSLzi1e34ldP/uVEnfg24uwFdCxqLqrUMO2iq+30u/ixSj+
tAArBiqK7cu5plteiJyMOciSVo0R3u+HSutvHuKXnfwALhZed6IIq7mNM7+1gIkj
pFppPu5g9k+Wbg/JAD7v+8BkNRD8W6rYw+ZxzV0gUzBNe35cF1lozfBDJ3k4ECwG
r1mQ5oQwsh63DmOggsShn4ubfFp2vH5O8+fiDszHGG+jNNDUeoz9mWS5X+mfnSbe
rVouFXMwE1jEkN1bfHUwm2roepyxhZGV0Q3LMuNQPNL68K+FAtMb1johvPSriJKs
oCv0XYka+mSk4CaBwpFjNnwtD1793cKGDs6J0oZsnzzV5Eeed8u3ofV7VscGnCx9
qntKt6IGG1Db95ag8mDZ0dC60d8D6iVwMrnpIaJGohnhFGvxbv16xpp6AE6JmtNh
vutP3pfgEFwl4Icxv4IAP0b9RSJNRSIapaomKcJyaTpYD/GQ7QmxNlWiTqXxFsjs
iHaPnm+kVhfJVK0kmiziR2T89M0sQvMgGR+Ju/1tL50ICi33YLz3WpaylZrfpged
RHt6dbc43FF3cZ8jYErvv1z/JEa1HFaJqQswfi0bhxhKgsBjAeNKYuLBF3HCD+3R
uI1mMlirF8GIYSYgCQUbDJg4tG4clfp2pAlHwQuqO6vbnnyJZbD2csSkQnOgU3q3
u0LuJt9SJj6P0BDTAkFYP6VPr+tzyeVq/jLn/nGrm1rO7Pz3AkqrrpiOAQ/WZqP7
P5q+OpYs/oCDTGTwjDY/JPTIJHfharZiyzhuZ/noJzJgfydXwLZUbaH5A1HQcArR
0QWawSJeLfH1WDX4rwg1B0S6lnRpUGdhQ6buYsirOPydmMKpEEsZisPy55228dEv
Ag/BNfOIivzfbU0Q8ctTaDOmVW7NHAoQtNAqfNrTUja/ANBlmi2fY7vr4YM3kYzz
6H8FSwj05TuSa+zKDNZL1aTr1KUdFLYnILhh660sEOMnas5o7PnzNeCPDCm9TiTY
FH+tgO2IW+xWNJUYcwZDQwzmSWanWWRcLYTdbCaXZNC3JX4I287zhR+6wE8oHQW9
VuBrfjdbF0sJku/cpgkFHshj0q+Y1YRdGrvnp2t8PFhfJwXkziCdJMqSYQLSnEMy
9oX1YC05elw1rboHIwbTpHtGajIlsmQQCrZHDVlnSOjxxcYn83lzD3QvwbYq7MFY
EAruuomdRvQnAHan83VD4/QP44/lY9+5ohfshhM2MY4xrTFoExt1cHBNf7LrF/o5
I5p90hLdTM85aD69fHRMYxNOpZkRI0lKC4dd3daHtM5r8UWvXmWjh4Ok4VGSFSaZ
AMKsZNJ0gCkY56PPVoIpK+ZVC9Ur5yI2i6ep1E/Z4uHHs0LXxLCkkIf7qA+BgNr7
EctsgONReZuapvNsSMLhhW2E3srfIjq9UjIpF2xuqBclF2hebpwNPp7391McqSTe
Yr655WhKQh/U+eO7bmsEJVjn3Y40WNjytgeMmQyjh3bhhJZHGWTlq7T+uPXvEnRB
wxWixvQyE20WXMnJ4eCXg73jQPKpWZRZBxbVJlhAZQvnVY/cppFW84VWbYU+D3G/
W482xJyqBJ5Y+enj5RapMDtzGc2tFq+8FeTmeFitL0Vfs4wrSukFi43Q9bwnNrhy
aGevR5Y9O+n9OFgKldxjyRgoU/GTzUX2xyHZ+mxA0Pr0gv9FspLFCIRK68B6NbhK
dkNWdslptZCvgv2MdeAH4RHKEjaef+lmtX1t39X3QDxlEgnB6C/4/IOAlh2MxFmT
WZKlqaJ90an8Gw9sAWCjahKwpDS6i9ToXREVPuMjR6jasr65gOlFLnDlO5AdidI3
S/BifinMUgtRO3O+HRN038bnokm5HhI/ms/rBUd0TQAjiqmUziEBCUNWSEGCfcwc
6XItS4dkqRm+24JLxh0dxLm/oU02lWUiplPNKWWrOrVZMrDk6QqqrjSZzVIocsmA
O2kK2JjScQh893cS/ouKAUbryQH683IdvelC28mKJiiVVvVd5FyjY7MNzImMJ/y9
aSSpx82pKw+Cu+F7EQpCE5H0ivIewUdEDNnoDI5/la/AjdsiOjD5WdPFjmkiBEnz
PfUIjOnTzZOlCx6mQCgTHp/9fRfo1DoO7qjGG5pE8YUGf4ru1hueLRhMcfqquSZD
zarvjMMyYO1qPAkwaCDeaNQDzZotdA4cQY2nwcJRISWcS3x+RbSdWaW2qR5KyFZW
RXJ2QOUk4WtzMeFdHK9VY9Ij4FrTAnygCbLbJvlUFD58bVHprbH0rvTZGfLwJJKM
E9h16JPEtcB+mXlL9QxqcG+9P7XixxHy+YzxvJlqyUHww5lXAb9JjP/eWrFwHIT2
s+HekRAy4Ju2RywO/PTAEmzBZ8ZFeEfet4LnrIfsVZKc8rZfnbxTLtnhBw7AVDBD
c5b17oa75K4NH6rP/U4U8IJWQez4iZZjlRl4519wl4MEIWSX3SOQznQr1vyFPr04
6LVADE2GT/o0kWAcFASY0soWiAfsvi8SoaatfAkKqkBcMGdcmJKgE3l7/hWPI9ka
vqVa3iY1l1rLNENP2+XKy746CTocw7wpGLPIffQqjgFHSDx7zJGCJEu9hKysOk6Q
7SEchOWDCNGIIybfA82gYWbu82GJtveRakB1p6U8yGxK+GwkCQV8hPAsWhDe36qC
NJaFnkJHTgHmorPWWT+I8y5E/i/xRxjgHI139JuXPEkjYAS5xJ7TBRXaLZmLJizh
IynsPrpclSRCpWcWSGbbMpu+jIzwKgxSrBYXlZxTLUDRUdaxe5tGeIaFGwMFXPBY
8NWxyhgECmARtUpQBt8xOMpbkdN+tfG1ycPA44hqlKuIJasRAFI67daEMKHSpI3q
S1fEEqO6J2uitwXdD/025ovkIf0ow17qYo+on0Y5af2A4BNSdl9GiNddBf+8Mfy0
ez/M5H/gr63aqMCRI3zbFpa+9pwAyhFOX2Ciprab9LQGM479ueH1XBxFZ+rmNJGo
2LElJ/KzjFCRjZ6iTONo6VCklXepWCBc+MZKpOTSJXCbdor5M2USvaXSGGUKX0+o
BasnWrkdkcPJZFT7PIbWwS84Bx9/ni4oIJLCXOLC9yWz34bvxdwTT8fCAF73WAy3
CWpRJFtEYru/c+rybOKNqg88uDgTbniThWQNakrNXLX0/hnEAbYxekdr5OklZH+O
AMQ0Y+tR4F1G7nYs3igAyk/93clEmNqhbv58KswJhz71G4m5BYLE9BJ3ibsXN53x
HiLqL39q2Y3XvUtsIf7150lepLeIBvrFVRji84VWWeo+1eW0Imf2sfLIDpt8JRV+
d5N/GduAUEkFwh+fO0aEX3NrgINZzczDWL8eps2ceVQSGdMUXQyKNS+Adcc/0kBR
6GylV5QQUhOU+TFUohI8v+VmpvxvtmCQ2keB2B72HfM9m3DNgEkZWpBopy6zxyA9
c2DWEyDL3aFJxZuXtD8EARbEYNk1ySyYk0QZUaj+JOh7GYMWIR7TvxRW7VNxrbK0
kXGgV+VUFek2wWZmcOnEZebMKNEI3G9+SVHNv+bmUY0gY+OKoyPwUCiRcn463w+h
l72D6eWqWgpwy860692TDEh0SXze5SICwWDbA+FJoz9c+9LYPfefJRJLRw5L0sxB
9MEsr4Md1j5nfQwS3liGd3AfCXAPHZ3Q9RfxJMij6pLr4mUnZqX/RPYFN+LPJDq8
4KpHRQKlvmLKgHfSleMeXmD6ND90bO029rZIGMt8Cb37UPglUgLYQ5X6QwEZdDC+
xb3SJ3L59gPczDTqltJaN8p+4MUCHGujFkZf2ZFBMiue6dGvCszVJOuFzWyL1nj4
RAaEAIr8WJZI6YA+yoqkRfhUPeA4Aoh4nU4AL7SIUiFQxZsRvSO2O5MZmDdC+QFu
iZGxdIiGYp0IRnncDQU8A7Bpsneq+SCRzUYsVJn6S1zav1+DNrO0n1xQ01lnBLbM
jZrDrD97nvQYVby+/Uv3YUQrlninIs228k+vOOeAqBf2LCgRXq+oWJshGmrXT+qO
n2naTBGupvF2P7G6tofOyRRgxAoNemlw2O4tjJCKjbIdcQt5otE6MWutdm8Pq7OR
pcAAS89zD3cx9iQxH+sEXKB5iTThBWuogo/9XOduplMcO9t7GgtI0f6VFgCuwYqD
eVgRagntw4bx4Ft/ZOHQ29XBPFwVGvZ9r1200D/ZdO/ZXAcSW9R6ZJ6iayijqVhY
kt2N6/KGiDqrAbtUHASRm7BPhHpP1yghLTvF8up6fdpHEn5wFlC5vMWmZst66n0z
eajx8Yq9RqcdtdWa50iGsreWNKodhIWQNfv8l1UnRvDVP2Ko5Ti9PKSTrMWTLyc2
sBxAR5ybMi9vYqgiTgSaqdzKKRHZ3duQaoaKjWamkVbhrSpmARcCAUqLQl0ZBdLM
0zGCJuOwLhpAXU+Q8vdKr0pagG3FW+Y1iZ/X55+p/6WnjyzmP7Ynd7ejgdgOa3kM
Bt6JMhUuk63He8Eb2RRxq8jlYXjaB/XpdvZF9ldAjirg1HeWdtaokyvVR2BnMiJ5
th5MmOiJjeOUwPx8UD4oaYZICy+qvK9qgPgp28vSRx2BzPx2BUHmVjEuD2blgOpB
pTwieQhl9no382cAZxUaf1gC/e3L/5GjpHrlSY8PjqYj+YzJyxXypVbbNoxxyzA8
9e1wovv6WG2o/yb+gHJovo7w3xYwihCEKiOO82gyoNPM5/aZCUFVCah/u2lKkHqx
9PAqNyAYJtow86Gbh0w0MXuPP0BExCJo9kXZvvUEXQQ7yw2eqk/SdOjFHtiNgT5h
7RYTlDvTfIZpI7z0vtph0muq68ZcbKXqjmoHCiu90tzMz6zM1ntPgayTvMAJggAq
RbgWSHAO3uOsvVWWfvXn97CYfZeFAvAbLcomkYLEvN7iG+D+N9PHvO5KxxdW+nIT
qg9e+z7T48Ot/w2LM7faPM1k8eDUO1J/bWyJxgjbyhyZeP0RwKE++p1fpCQsvpQK
HB4z1s+BMUygtzWo9/6L/IwYA+tXcCvAzDkdyXEFCoNhRN4i2tTZn/Cznkl97el8
+RadOkRZhu9PCo6N1+seg3SYhTD19CsprD+zJ1LR7KrmQ1A27si6hdBJHRaBLpyj
FrrMdpwZxHXF93ukVpf+tzAY2V74BZYp0L0BuwWeUUppAyLkQ4GTtlrOyHNl/adm
5XkKFfl4lWi7f4T/tojrpeGKyJiPi7RbGeN49vCGGXzXEo2Tq85/vS3M//sIC0kk
pKKepiZWzIRsnd6i2BOoxXzeMS1N5dPEL7ZGFWDFl+4Wiz2kRtrv5YCyDOm7GJwK
EHe4zfsmGmEfPG86YB1G84slhClC+eelflZ4mOjAkz6j+YJAhoSQ2pDWZp471gFR
Fr8rAjJFfL1+jww23SEqTi52+iGsarSZn4qRGlU8QJBAe72f/UPJhB34zALPRJRM
W2EYiygz+lDvyBgppiN4N7RppISRYP9S74CtV7r7PCPJ5OzQBc0zFklUlQVHOBmx
Yw+3soyp32yTj1pX6nGFFvROogNtkEm0zn2yEIlUnN+ZXoRHVM3oxTSyvIq+J2JP
4YdOF7R4OJER9Lq8Lqq44gFYM95D/KZFb00fxqhIH2iY+TpYT/Bjaz3epbs09AZy
gaR2MDeOvkHM7SVEoRbqRXRRE8N9j6QId8izYZEDbOrDw+kVhEMoombNhSS0O7ro
iWCfRN8IT6u/Cr+SZFl5orKI8xRXye+UPJ4j3ku/h1M3a1rjnPTf4W941CLruNAI
Cvq7sFTkM8n8lT+PR48N2aDx6qzCy5ejWdQJGymMGWmtBpcpv7NXwX2XvPguW0Xa
YG+85z+bNZwQFzK732nYRTZ5JSgUBUOeE12O3iiuRtEOwxh8ncO7EXnBfOkk4TcU
kmcxDcbGPH5dTwv7mc13GG90FusYadWAnc8olYoVOBHdQOYr49enarTkLMLDXMu0
9aeqg8vEyz5Lawr8pP2eq96gJxmLTq0i4gfr7IPYsZ/g2ndehYhN5q/+jjBxKaAO
aXtBwhQvq4FvQgKmccSTJGbB/I0ppWqKHR9Ee86+4rtzDEf59FPsqWXQvyiqH5/2
OzeUGjxteaUX53Y7m9jB+lDr+cYunVph+5KPLSxmHlqNX+qKk676pIJ3ACg02m6C
pxg9G5r0m1CdPFLyQ6rw/frf5HWn/HjVaSACFrBC5n1okenZcOpF/2dEv0cR1I8z
xfg5uP/B5n2Dd/HzTmbs5AuFVDrB6lHZstoBjYswiLTxJsWeWNAFtzszmtnseDKn
vdFBKsz5gDckYWxsWDye6msBlXWILJ0jKtT8ZY3oU2T7UE3K8P9BECjXN+R50SPw
vZHUa8YegsABwag9RVk3R7bSOs6kFe7vtTWSiyqmL0qo5Rh7noXu+SOGqtZvj1hs
RWMArnNY6RhhAlebakG+psJFB6kHJZALOdeEVcLfl6crutqhuygVgvet/I1p1+2y
V/NzsfeEA+sDPbWPALn/VXodMDFtkbGhmO03q4WUk8zjsNtZy4nXFd6y5TDL7iJN
u4h/4VuYNCR/Bf24UphNY9kfkSeX5boO9W8y7zjG7/e3+L98bCAQGD0O4EFlP3Ak
IiRbipt0j9mn2l35W7aDmmI0hfGeg7xE+OmEZDtkyjDlbOaP4ONr+6IPJm+Bdk84
vD+GQUOIiykZ0yHhOWYGcWDUecWVo6eYwpOpXQ11PB4Vg1z++YXPU6H4/4ghtyPs
QNHCuI+JaoGgISw2rEVs2fqXtBoo30UMqtsbZJCj2szbyc9bD8H7hPF3e2YllMzs
Qyk8OyKDtWsGppCqbkh+WJWRld92AMPePTqFAkrkfIrTCm7ysSud9e3MxN/2h9bt
60Z+UHqp/DDD+XcjzSWDE8t0flcD/sI3VkvWgsdWw1oaR7u9IRGA1nr8UOjGKNas
GroLeofLAHPXoO/cn5wWDNl8o/pEMMNr8vOwourZrWdvujYrkDxl3wo+NBpmNVRh
nNsULFPUSm4KoJOZLUTr8rwNnbPspU5cka0KKEbC0Lz5kGQjb4G7e1zqNdXICwxW
v3DS+pQ5wuKwbfNe1ur67yTajqSGL9Dklcni9CXUZli9XlOgG6wumsDrOeCAr86q
eqVWdbYfzK9py9GxIXvTa6w19D0wTx5Qd+IZ7jBASTCmGsSQ0X1olJexRDrfGsZu
bwSu7hxRUyQ5kHY+PCEI/09ByWVqG/B909naMg+40qAR8bmzp9UBNqIdLF/vK2Ji
K+FQ29BLnahmOfvvQtyumd+TCXh8yVXbB6vixLZG7lnNxHJOPq39otTuwWDye0kk
Vi2JRtIQqYyfZXmHxheOx6tsVmCeeuGdO/NOy2njsrCW1x8pPCORQwXIsZohDlsI
wmuMISGr0D3vd4UHrfD+SknkXoL6L7049NPDGvXhO1d3fo2jHbW0fojCDhI6ZjfO
WR1y2vAStTy0F87/6bbGOlKruvn+KAW+56sN4m9g5pMcKJmLMmCTdE7Wi/ridUi1
yep1FzJHl9Omy5LnS6JUtD1Vv4sy9ewXnr8uoAOLsR6Cv/BT1WLtbexOatx9VK8s
fWnQ7bREK7iL53Jq4Yjiap1epsiSgsM6PMp/Io/KxA/JlmCnNsdY4pOUKooU7wFU
NErIs3PmEbFE1ZUIoIqpnUOWm3wv2HSiU+QKcO05uyKlraa1w4/pyUmJ6L46uNJ/
Ow6f4Qn9ryU7WhzK3SQ4Ysi9o1Y+6DmqyO1wIhwrUPPUw3mkHc+5jSNTcHKXjH15
MCeH3ZtofNC6kWk2cbLtfyX0kSWyKpx9blHvo/Sp6EvHUIl1chnp37ETrGYuN8Ow
blOSkjiJ0r9Vats6XPkxZe2kjsHLYGY5aSbtrJ9Lmrlrz8ZKxt1G84yDDMkoeyOq
jRZRSYfXTe/J3TnyCTxEr2Q2BL8AsxrtekWJ21X8kK4UlZ7WvFEADKZ465LS8ZaL
w2dvjbe8+4r/E0dL1kcVh3z+S1OIf6TGITs1n/LBFGZkuPn7ORhtQ1armZ8YrLJF
IhoPdUp/tqrNbXoSHUngHZROyVsANy3mTjmpVBMS/pCCraQYv8tJtCwOXlRe5Lyp
iED3ZRdozeCGljpzc4obxrxsEz4MBsiIxmeYFa85qdoHg1C+g4yFzrM20o8qk5T2
6GtbIEeqIozpVEXYAa03abh/LhSgIhJ+3Z+3rfzcAHaLNv3KC1s/Q8oyOrX0u8D8
Sf6keO1UgU4iKNeuQ7KgZRsOkyNEcvLqTuchHLKqxZJdMKVqccBWO3DuEUtlRJtd
iS4csVZptMLU/b6ZeGERDhipDlOldYd1i3CEBWHOOUzrQnXmE2DLo9Gqb4Mqv40H
zFJcAO1nTjAZpg1kOgdg7VkIeDCMpNbO2BwmShKZg8rgnSl7NKGie3L0zVb2NeCJ
ugVs0T3/JxzggzXkiATYVUdGkTf4xj7NbOyT4W1sP64KAL9/GyQ1TnCyxk5NDe8M
hFMg3lA2ZZM7oHV3QUDj8bdHiGAweKR4BmEGnHR2Y8cwr1k76dZiB7P4M/ghYhnm
tCRHLOeJIJ04/JKc1gnT4RzP6ua4Nw4gdrhKzRQ6lJ6f+czktPYZQI+0u1xgfxxb
BqDg9K7xwM2NihMPOWfA1lCz8AxJMoG+4mirL57EuRGrKDqT4SXPSRSc2EqcTtPG
KlrRCPlrjKINxD4PXjeTAboNMgS3q08qCJQKT3rWLYsxNT5lNxYiDcr7ePelrD3g
GVLEWwPg3WIb9Hw7otFwYm+3hUIqvJcxfAuC7ePoiw/lmqVd1Y7mcT2KsjX9lf0H
HaSeqwwPe29N5QYnMzT5rcgS8+PBoQ0WKoPSrp/crheOOKTbbq8j3pneKLLe9iKv
b29H/yY85khhc6GtFpUqWNU/V17tFEZo0HHiJrmDBNFoTVMRj8P6NZ7uMHjee/z8
CR1OXPYSsT8ewTF3e9fSLz+yMJDtQST91CzJFMoaX0OLsxlohxeeh79AWtP4k8Iy
c/CyKzSzR7aMGOnN3xYis0CDmfR5cMRzbExXtkz0YbT0kVL+8JyYvvQGUWcZO+fn
grnjNY/UAo5euGzBEv8xCjrJhIY9RpN81vDn28Q/6y0dFUUKL7MQ70DB5m8QIaxi
Yxz6xN7WgrDSzKZNFDTk/GlrZGoV4DPqoe8a7udsvbr2cbADoJNx6AknbVNCwX19
aOIb4IsTWOAc9UXeAvVjaS9SDPKfZwyidDQqqp5lAtotlpPRjObfjjL52cLLt56K
yEFTh0wo55dscHH1Oj2WCyUUn60TbsvaTK2cfB2YA5J+dmW+pDY5UlQdqs5G0MMC
nDCxLpgrNX6IywLpHXF0gyKFmNkrEdOf9bQYz8o2kHlHdbqb26ojKRbFnnD0famC
Iq74R1ctcDvf1vjuSzfy/mU5+F7UKVlhMBWnulhB/wV+yUVVVNYqTH+eHbWtKg/x
nheUCEIhd0R3Wf/8XK/E8nbbO9BtxEEi/huGbmYiDnwIrsF9IVOFoKl+YnQQtCG4
UULoPp4kA7CgYS1s8TOkATo6b01jmQEHW0HKsGf3+t2GMETnMzRmZVCfFdrL7Z6C
2xKv563O77olLKgm7mnIGjSgWV810BnIWNIpRzdX1nZuNQo7QRw5aCULJnAGdE/N
lbknVUpNuUZA6wNPoWg3Hn8XjlgNwEI25BVxSz5oW68q+uB5ohBm1r4nlJMARxe3
WWNjh+yQ8Mxo/AhZYuKwrveN3DG+APKPGteOnnxGN1HaUQq3jfeeldKn+m2fOAWp
SMO6vHHzME0bq2AVZnJe98YE1t4NJsE6DgTlsRAbyds8fKv84SWjazdhYQfMSZ3m
KedEsGUWtTKmFg+0cJJa7BdbSGE6J2NK4A/wlMYjlKd7WgTqjVS/+96m3KxImZat
B3rstXorokx49RAHbub2vZlU33qlzSmAttyOz4G8tkUkTN5Aql7eXDDOp3Bkkc9N
tm8fPN9XsL+zUt3JHxVCuBrQ4R+5M2mrQrCMG/hPaLcHQmR05jVFVnVNocwP+LNK
tsZJLsOaVsJpm52NSUXXl1p9V8W2sCm1e2aIgILwimtoTaJdY/KJJQ28b6wlwLfc
3yZJOZXK0rb7/RqCf3N6X0mRmFT9kI5PQpexVdSaFiQaluh0IBm0KaDdlHNZxSZz
9k4Nhyawinerr7NyWwGbcMKeacqEYUidw0W/laF/BSLu9ejMGAayBdSkFCkK2E5a
Hu+Rhexc5MGNrohfGWwOqKQmt3zg3ReZMW4fbpDu2j9+XVxkcE3NQ8afE1/6mDNL
gfeYjOMvQYYhy5/FaaktlDryQ9goxPnWdCPyOs/aUHBbpKbRu69mft417cNsDK4a
S40aAQr9RPQUnaDZ5TrJAF50npkongJi4pyKVxYSJgj2fsRH3ZA/k/hBO3JJx5Q7
rU6buC56K2NC/0m0fivIxA6fgNH2CsWX/aJ+1SOxN7SIkOKkJhrM3cx0dTQQ7FJs
clLMxNQSnPR0rJdIN74KQri5Q4dMn+9r+3ihqYlauM7SUt2CcbeeSy2oHqVosUgS
+tsEBqKvoZXFeF8+QXWULpyNXkZJVg4bDxohCKqLOolcduKqyuQhm43eoW7E0fWh
GqmJyr8Fimkw2MjjDyZ1Kudh7uzG5yjp87CNohrjdb9IBFzBgPr6LS3e0YJ30c7v
o/hljGVICGZNmEcFcrn2/kZ1g2ZfbcwrWCdTO9V83JaJBl0B2A9yTjtCCm6RLGVv
SYTqrnMdP7xo0aXgCZufx2KESkBR133E/zUOx+xJLvNDTyRi46WnWDZrfl27MNIF
+kiBozr/DpRzCNg5qQp5UIUzJ1muRbb/O3xG36rQ2M43ifPb/AOjXMyEi3VLziAD
IrfFgS1b61REaE9tOlgCSkFcxIS1APdSCtNlnF/ZVo70MAFBfFFm+C8wH6JydXIP
L8i+SAFjnwJinyiZJhadMXFEIPJ5k4X6fTqZi69aLS98Lu3c4l8vFl2CrtT2X5XL
F9w8AOOwDdLmcqyQEOZ2GMeVEeb1vEoZ5GAhCH8Q6K5k8+x0+4iqrpbsnauToq3l
JBrpVg267EXmFvnqY+rW1TrdtMcl8f+FGkRgTBmgEYZ9h869RNZhWNN3qUr/QW8V
alk9yh665nf+vS/r8TWuX3adTNGjZjFpNmMAd1qkYSgOGdxsj92IP1mdaNxLV88Q
H/3GVNqt179GAA4dElUvbLPW7xjRKw1NrwwrPFRhyVNM+Xuwi2niG7TrtEMdfw+9
+L6sK+1gWkvVv8s8gOc8YH7KCvSfvUWSVVmOHg7as9Kt82YC0QEBFKMBqgbjRe2C
mC0RZH70J/0HmVn414ZPfJ6AxCjjxAXMcyCG9eAiWXjOfS1JxRhq+OxQn5tpyius
yPcoJ68DVIBJk55KkVOKlS3Byem/cjG7xYJTLe2kqvXfeGuT5XcGWlL7jZIyBJN5
m3khw+Jm5O6byTbp0yfdFj3/pPL3HEBSc+kWz1wXOnBXWzcttS/MZHJtEHAeuzj6
yeaqCwvvIjrZ+7zFErcvcCwWTQ/vfB1KXEeDv5FB+7pUG3XmAEPmU5KBgwLQ+g8U
6UBId/A8wbQDeNLDDiTlA0cABEzhQ0H3VtrPhl4t6zuL/uHjsJudfP89yx3jpyoW
BwApJOnf4fSVa1GxBlv0U2ddOV/eRlzD5d2ETXkB979+I4fpWvky4TrnfZLyCcGe
7C0BjkdqyUvyfc1hx0zTHD++DaUahD191gmbaCOWF5Q7/NY+jNZKjlYMjElOVPsW
1BZbmH5n0zsx1nMXq6ywbtTwKUAZUJKtNnZPkdS4xixkHRzIrU93MPX9LOs9JGTX
Zb8dlovv3zg/Y+u1RrkuV1aFjOB0jkXUw+oEcFCg2GuYjeu3xOJPL1oX89pWUCsR
f33/2jS20P2ajlVP9tWrCrelI9kv8E3Aa+SPq5hTfq+pIdmy1yHwJR1Ig5SGjsJD
5noPiBenwUyxSzcY3hA/5ydOb4KybFeuDrJcsSTVjIAB2/xxaK0s7U5dsgDUiUi4
38fTy+pg76TWh5iQQRzQyOzyLszdbhf7j2482gbCui+N6APyZ12IbB6pmNXDSGX5
9SRD90fosq6TZW+dz8DCPHF4IWsl2/xCxptMSsw6RLRDTC3HFGRto+w9XTQny10U
72Piz1qiE72FhgUozCsPOOrawqQMlYsR5QQGGMAllZjNA7xl1+r9R4r8IbdJXivE
Uh/9fT+ERckK7aMZoG6jL6stz1gofs0VrFqRYi1U4MhEIyYkxevYaJrrD2B/gKk3
PSTNozSzFAh5T+2EKK7echgiMSLxfw/G/qlPVDYrFLElKZO0tH27MaGQZhehRlqy
lw5ftUGseBplYQ8BrItXgLZL1saU+uPP6re0IN50BZGq9scgeDggfQKLU9+yQZQD
gi2hRqeK3rGdHKrdLTlnmxdVLRrX4/PzOh6xVcPDVD8V52TzpnhKixbVY32o/Cfn
xgndIZXsG2QgHQNXEHGtJ/3ioKM3ZonBoMSlezs/D3WbdWO8/WHcbPnpW8jLnJGU
TUhR/PNP2gv5QUikrwueI84oZ6VY9uRFjyksfVkYn1PTDkFIGniqDCzfxvPw1tLP
vSCT47JQPQ0U2Rjr75r/Txv1SEkFMfRaMub+xjHtpmbamIhAs5i02vD6vRy2r04D
gOejHGVwJwiJEcmaVqaUglY1ptqBDDKzivCmrlLl1nXGdExxz/Q0qb7Tl/wLvF9w
9xkHJWrxEijhFT19iHwhcIeVAvK3MpmIOUfPG1b8yUgkd79P4kAVKmoZ3LfNHRNz
HKGeMxsFYKYQGjhaJd5GqyVHU/hweEZ87016aF7iW4VKuxTbgBsIvddp5S3l1RX7
wubT612ShqQ4CSTGLiE6DuE8uzQDfw9QKZGBVTWSJ6hNPvrsH5Kg9Lm7wPIaTqK1
UMQ2rPEm828+jdDRnvbtw8S56fXPSbHdwlyyzXM9M1dNtFpZngw4XlSsNwE4e6PI
yJpVlaqhiMFvy9gnUoBKm43s/p/IGF5IOTvmGV+9IQ49wLRznWyjHqXlqibFhQRp
41VlwnsnwpESqDsuJCc3eE1Qbw5daTZDENcmDnL0b9wZGymW2BW3hQbpZHFh7VY6
OfCQvh8KQQa9NgbL3p0LW5H83Kb6tPmzmXG3b3IL7XS8/nDjKlmllShUpKgaorI6
oaZ6nJ7VMTf0dHRIBINFEHU51aqWJr0jBj9wPGs0OUjUqGL27Bm/xgJMoS6oxlhe
QCrp3Ey92uBPTrImXfp/niWmsCsdUwl7j2IC4o61mlB8+lxIdJx2lzqMFbPYzAdt
wOy/ZYxsd4txiGeuW8TmMg5xYBFsMVSwBVz3rC95F6Kk7Lunfe0HGimjfRxbzqw7
c6U/aNfpKRSUrikTTZrBz8DdppD4n9nZDf7Z9BzyROmxyp6fRZWtBnXeVKVpjaJi
eOH1zLjQ2Qx/05ju+2f3s8ARcob562O3ffwUcq/aHX9e/hibp2L2X1QB/1wkXMO5
TeVzA2RHRUB9Y5AmYmAKqzBu/pRFeLvJvq7iDjLyeYQc/gay9liSYZ0hxQRfplsU
eUC6xMaQhABYtVZRSzeJeIc8FGGD2IhnvqxOYsweeZYlnR70RXsmwcB+zNghad1X
7LdnJgJbJMIkTU+22niTyxho0offh1tbYlVdaRFj7N/97xoqBsYdMFk1hsT6zATU
pMQkwNUUIOqm4SnnoUSd+/xCBFxaQ5uWoE93wICZLpV9MOZtYsus0LKm5dhuxZbh
EnXYFrGu6he7X2HISZPrc0HQSQw2txcUSt9HDu8/iSyXLdS2yb3e+Oa2pDXO5Y8c
pAQdLyBPtniT3zLfcNQHWCrazoOc07uMXdYzp01RnB33Gvmu7HgKGtxDgh3I7Kb9
2mC1h68gKXyx6Pk73EJhsquCFfHTuSw89XJlWKxRZYF3DFpsnwvgL1AYEqN/90OE
a6FeWMCCZCxH48HJdqIfS0s5+Dyr/l8ouB5JiPPPsLcq+gBuDIcNgcf4sUc+rhW0
TMzG2UFjFYPsCEZYFNs8oJhzNVwwpphK9h2P+KU7r5yCVduxAFJ4DnniY6rFU7Dy
u7BqPuQHwT8XpOgaVMDk/N/Sm9abS8J3RAPUrJVaGQYujP4vvcaemuPwIohOUsyB
Fk0fA7mqsp727wyI0xV6y9EThO3v7ZfiJbS/SYUZM6YpEDJ7wSMG+a8fXzOyFNwy
QVkMS8ZnzE0WP79QOsPsp/fhDt9UJ260g5zk5onrDsbc+Tt3r7Fsxzy8EIl5QLk7
BXBIZHeApvLCTTMLjREv8lpeu7eplOqVV0OatJZWsRdEohWxGe1M4xNdem0eEwIs
S4KhpMqfL05yapQaVFtSfQvVkYRnM4A7UXGOJgZOuUDaJ4QnRddSIrshZrVd+SvF
T5lhlJqLrilo+ho0iRm9URA20tmd1r2irKVQh6GnPjZ+gi7rj3Cp+qZg0lFgbCpc
7GPyUWb8xRMz0IaTvJDLl63oD+pC9LDxrLKRN+iKfZvnjyltQjDeSl/W8K9E520z
sJfZqF5cbJAi3ILXqd0KmZ2xgOw/RPJl+SDqNIYiUedS4zgsFp9uIVgeEz8QYLwI
xslaoqlGYzq0Ti9yF3H0a9TT5gKUTQQVsUVWAAt/x7MrbuS+aNm4XAve1H8MM+YU
mrh/kX66CHBW2bHwcuf7KYRX6lwqj283cQjdqTIfpMZ+OHsDT2nkund2eIUtGagE
LiAcOtWoj/RNpT/xSen8RSrJdBp9dtnt65KZ7yECpdGaxdiHbkirDYIwiRPDxMWb
aS710l9z+OVwlHppNaYPO+pFa6Hj0Fk+xK5nDhAVsNyVdEWgX4Xv/vt+OZt11DKw
CkfuEkEy0Av1btOihQw1WDiYlYjsmoxB6WQh9NrGj/oJk56dh6tz+wkliGpuXNpY
GZi6O1S6qaRUsNQ3/Mm2EbkYL0sWwGvPafFHdtIbfR6XcqMgbPZyS1fJQqN0RjFc
/Sjo2/44UEwORInI3bxHL83Gk/MQxSP2FTVBjcCOX0sTTQC25FnZ1OJUVroGW0+U
Fpl+ekr2OTsRmTm5e4Wjx1QqFqF77cyNTS3xr6sIS+rmqO/4GMTkkwCRPoym4V0t
0oA4qGzFtHyyoUwfWrJ5nDtqk5yy6b0D5V2Ld1s2drsLHjBpTHzJ4srU8p1juhy/
WdDR9wD3xLAHEQWMatVBpC7cRkJ7nNGrlzDJ3TFHK5lsWixnruFQUg4+HTq2dKTx
jrJ/qec2Qe2/aoUwYDzcNssZilJcTo2gAkZWJGxxHLeH1+8s2ICrhwbaLmrTT7ga
oGHOu7BY67iOab17HbPorYKV9jiRgO+GqaPcmYBOoTeZQ8WP6J37a2yQ/SwRfRjb
we1dwgjCJDLkuI3ZkDg8qAKdJFSGsRrfqBdt/cOl/CWXisgGggXeKU0DLZEWZxlZ
Yl5WpjA6R6zApizCL/iD0amUCBBOB04CzXzBx75lmkiJZRva1E7X2oZymzYNn224
5Fa2bSwwGY6Fe8yqt2qSE8EvKiR61fJ1gjXIirjjnNFmVuwsnZNRe62693lu09q0
twxL0qZCGuKZTsKcjG92h/6wEuIMnVfm+GVkARoRnf2D8p5+TMpz7SEb51ptfD6D
jV5DCv4OZIPZQkN18FPlai1KHKSXHZPBmDDR3i6Mj3oxE436hYfAtY59+TLIGz45
qTT8HHxrsNPEf7RGU0BtYLKRAIKkkfUcYkcUPuEbStOtWXJ4jnrOewORYBpfefVV
6tdzUPSoJ+htFW4ikKGoLSIogn7b8yV2pkFlTEMBL4mrEbmqdHCNcEdojoKo8c4J
eUzpDm/0B7rrwcsBAfhve8p+1abbPJEUqOlk7NFwdUWc3JyeYvZaajs1z0nMRdl4
qVd9wxxepxyOs/tAwOE2qp5w3szNz/626dIo+ime1nVv8AEz5Fi3QMPp/c1Z05pq
lM34ar95i6MdiYysHfPp4nLWD47K/GLl5tXyRUxf0AS3YdR0lQznBkxopQqVfd7S
rzEM7IiPeXV1gA4KmKznu7HkoIDWywrV5QfmBkb8jGeXTcUb+Xt8qzcupfd3iOFI
BTjdSZENzy5LGz/lM6wwg/+wHbJWJSa9kS5RU+FEObEenFGEWgjwihjqRb2Gcqqd
SS3W/Ak4MdhtZ71VdKhd1GogaKvwk51vfX0Qh9Fb0d0v8b5qzR5tbVL5AjE8pL1N
J1DosivUAt2Ph/RVuYcY/lXDrLffvhxwaRImgIQ9Lf9zZbCJYtf8f2QguuZNZNZC
fhMKZAIJZG28DCOIBodZPLzhLHSjNSmlC9v+OgPi14n8O/TzJvKUKcDBqh2kXpG2
11JRa4XsG6bBcFdxs9Jh3bPMcWSWV6RJOOx/s1plcafeosHG3XtMH1WP2tPobbgU
gzmYHtX5T72fy4woOYyJhlhSy8U3mFtm7ksPEXqKFjhujsUYKyLsDv7d0rAj4PSx
Tbr7gmt9IgnX1DPbHMH/o34RIKcUmTilxj2IHAUP/2uJW2AS5qUsySgqf6E/PVcq
Gr9yNloZyBl3udeY4bNZsBL3UwPOTOk5b1WwsZxmPYOzL4GEp57QyIeR+GglW831
4NmxQevuDE+TXlViIttJ0taI7dazNMyEEcfz7h1YpVCHwCoRGLp32kpMF/vavHXu
wBBurzy3nselW+OCQKZcfhXCbDb0xRJkv048AoTlumA83YCj15OYaN4pGFeIsQ69
pAY8I0pdh48f1MUAJgWd0lt/Ud/bn0gn3LjeKHCaHRG9MgPihqmubzZN0kzi5ynr
lgAxmblgziYwPVGY7zduVklsUdsBGD1jsFesY5eYsJVOae5/tAuinDzADOl7/K6L
FU6I7RHgi8rp26s/nTueWRP8bv5r6GJ1Es1BL5A99qC/MRmIuMdtprWT0QLW9xhG
9G8wRu4nXj9tAdFLz3FoQCRZ7KBFrglGY7tQgaSlmo2eC22/ZqYRJJS2lGgvKWql
hb1pEqmmHxIeCtaYxTcH3lyvCXdUcL+3pO6bAK1NU26LCH0tE9/apR6vMJGjKYu1
tTp92SnRitvUNm2BawfQyTOih0fXLn6VNHgFoJwFCOqtC0T4JIghHpQ8U+wxYT5W
u/eNvBZMuqK4XOFmiAvY3Rc0SFjFfSWZ7HkoO0ZGNryu8+b0dd3qY1aO/tlbfm6+
Lx0D3DOD0DXI+IJNG4g0+GWFW+Jlsr4M1C9vG6KH9iXEh4f3rZGVtDbot00PKhQG
lEGx4AAjqsbOSYFOuPMIrgLoPqCNEhCeuP+xCf79sn3dZUjVLiLrY4Kbt/dNLD90
sQKUeOjzDXBuIVZZNpxIrUNFpWYQeBHh8M82ZcxhJgMJUN6GZmvEfVuD4ht8NCMc
d5h4TljGjH578hexzJIS1H/L3l2dIEGzye5by3eFD7rSPaJDLGWDu0Xk5PvoF2Bz
Mvk4BMduSYLjTavrudNVUqABaNSl5J2/M8WPVgEV6tiVIgqm23icmb+XxGQNBCwq
hYQTxRhFuw617QhHk9I9aXa3F+vAyeNOlp4CxcTGvrVFUgYMCBIznZmQm5MJQ+4J
G99YXc379t4vliz2Fc5nDUr0EYBSXRNTIzFe/yti3FOjMAXbpOX0kbutCucF4WX8
zSfi5FtKpOVkTYTYEiNKgkdoDBlUD8L7XUq30+u7f2e6LUdrRVCMS7021Z7TBcru
ISzb25O37pO/TeW+kvnvpMkFuFUtIweHC/ExntKRiWOll/T8QuBpvZnLLejMIpuM
ntKKaNsxf7GvfmqiYTA2NEruyzzDs4VwOx1zPc745WiF95BDLBJGpLtFxe8jvo+V
Ah/NdveIFbLzwSizhjNGOuJa0uXTh5WePHHgofkNCMc/3bpvFD+z20QGneGKACSv
UTzdi3t8eM6kEQbeA6isBaz+03BGD8vWoeFVU3cHdDR/t+H4ZF43EAiwI4m7CMCk
D0aZMPqten7eZ9YMwa6vUDWyxM9y+1EgO3qkzl9Tyfyiv4sOaWiv9Zj/RvghoVDJ
sfqA3W+w2UI+i41jrKDYXXzUNlGD4f2ciaINaixzV0Gh8/Ke2DRDkKZsZ/5OS+O+
m83vde+vg6QP5wJmt2L6ZKl97nLBqepOm2FL5yIy+7GZcUHykesCwJ2JaSOG2TaD
mW1+M+ZciaAPNDBFc8HsszS0hRHd3mPG5zKnqC5TspiD02HMcl4iLEFuIVbzLvHF
+ttI//qjapXibTBnmBlAOBU8YeEUYDhdk7/fcSfmDKWi1ogps0AJHH/OAAIRgudk
phCNx6W4lD/YRmcv0JK6wFy8x1yjLL/NvyIFypnPDO16ge7AYfN41TzgCNWhNCEv
Fk3GR13cAShVAGCF7phgapGC4i3oEQOQ+aX62nUoWmXE/udxXoLnPuyaGpp7iffb
eVFTyUNjwaGTilOSjw/3vkNHHrtIeAs3okYkCOKeE3qFw9W6XZffOOnxS9EtNUUi
0qSW9qSLJPh1C6JN+e63urvZuhI4a5hPPUCdthUKsmSwXLKj4o8nnjHarqX5LXBG
U4Vzp5L1NnpHj00+i4rrpEAckooczhZ+aqWZc7/9e4SoMRNKWuBL/k5qp3IRBUb6
3V2Dj8kV3/le+2rQ9bCpSYYeqF1itJWWHnNitI4XaXytIMQfKKfUJfPfzuZ4byTc
+ysksUoftYCMYqjferyqs5hh0DAALcCTMvngg84u6dY1nkablfQqCTPv8d5K+2YQ
EtXSD6WoNmRYaEBYn5EUQ0stbZn7VmvyudPAh2cwA79adA0SvajwoYAWq1dmVenJ
ZOSfBakN3HJQH/c8XmuCOti5BeqDiFuD/pFyOXE39gCyXtYwwa8KGvKJZpvRxkod
L2NzjUL0oB4vNMLj17Dc6jbYA2Q0wBtfR1yLYOe+wqDrGDMRwd0cPXGCqkCSto8g
9yQhJze6caOptDJMc9mKtfQcbXHrHGovvzhf2VCF9emG99VjI8W63cPS86EiEOYb
iQAwpULSlk8gnpIpKNV06Cfzu13fPgLDTU8MMIknfFRCSoNhhVoEdQU/urD4AHbO
kLSphwi3a1LwYsnQr4ZGlD/sctLsjNCi/2v0JhJMa6KKNbhmLE+o7qIs+Q2QErcY
R6OKDTlRRG7P4W4WXNN42aT2K8Xj3l1DwY5qkJwuPIy1EvkSheO/NBVDAEI2dFUc
pyhqEwZnj2qGMtQMcir8nJWDDnbVvrGAK4PhJZSAC9iXEO1jcdPEJS5j0MUyDfAA
deCz3SjgcqQpuI3dNBlPhfHMlcpnLkfsxvZ10m4yjdmxUbh292jHkAyHzl/Ts/8t
2tZfA5LIDzXr0lqVU8pS0kQb51rVXO0sUEEZ0MJVO/YGTZ5eHlXZ+MpOP5PRA/RJ
P5bA0cmoALaTOG5QwvDehnbznw6BnMP6emmtplLT8pl1okzzylwFUy+Ldkgc2EUQ
lXNjB3UT0Dp3sE6encsMx2rD3uQmdJfFKmtSMS/TZZqXifL5Bm58PSVF5Ljcclaj
rwH7dk6PK25CRMNl4lS+lTNI4xQz+YU6QGGwTB3YEF/vg2kPiGp51NAFO4qNBEc5
O+EiaBvIIam/5KUKqa/Zg9OzVy1+lyoiWk0+KO+F7LifS3HF9cMXIXHZ0lM4vFoU
XjJTO3V7crTFlEa9x8OK6rWslAtx3lXRFckrq5XAZP0GczFR3bScMmMTU9/rPH2c
e8umuZZvddmP8ZuCWTiajGnrDeq6thxRnj26Ju3/80Y98PZJtCetXNOJ0Cuvll3N
bNyMVRBZBhBgh37tF+ZZKulNPGkCEc1aqi0EZvmdBXhiWFGXER16KkmZTEk2kKyv
Qs1qzQSnlqcWQ4wVQFqlRZ65e0s3/Nb6PzOYPFAYqa4vc8u98LhkD7NOMiWc8AiU
4nfOCYJDblzHuAiWyAnsTdwmbTlxv50NEGcTprB6FlFF9yBOhZZfBuFeZ9ZX0FlL
+9naj5kkwXfiRtILeY3zuvsu8I45phLEQ9PpFplNQreVhvrK36mRlMGwZ4qvnZuw
Ak9Mmqfv1e+8aPIdvbkO7003yb41g89SG0XoYkvirH+vcnnRktjCPz7h8pLb6aaq
8l/hVb4wcJhVWaYlFtFFMDJas2xd/EVMKWuPpVLQ8728mxoNfL6hDOPJ8jL2VWg/
QoeV7E5UNBvkWdDgJs7MufB31bw5wTHlEuv+oUe6utH0TZlHpDRZcM1CUU1o7vOf
zGGHQHbRshray0JkHRniLFZH+DkcdSVSCQ0U/GpypM3j8qBXdzcO5TFKWI3zmfU/
OmL/pXlTK77hWacFi/Z7uASTGtDMqBoYNYB2rVp2/dMxUKTeSbhcdRWDoL9NUwQg
AslINya2HkvbRNt6Gl026hJcWW6zT8s4fj03+Y9jlBFXzc5LLGg4mOZN2o9qLq/n
oxQ7LGsxpwjpbZHF9Y8xJCKWYtfX58oEUy71ig734ZZZ3MEScNoSnfvKSfiOGVqZ
phLGFM4pCzJDVkg11IegRTMex7krPnah2KKePbPWY1GYnteS8/DA3enmDbx+ULHx
aCXsF1V/vKDcGZ+9/O40uaWDrVUGBuD7g64rjVQJx4Ezcde1cB5uKf1ih43aUgAL
7I9aInTyUhjRyU35vjh8PtKvb1E7T7/pcw+lvX+zCZAVFixXkIQTvCwI0GhtNEBJ
nWE2EUooDZM/6/dO/ffO6GI9OkqStEjf26lAVmPP+bg1KNBsLlXPQAwDyTboWf3E
D/7gYx+SQs1hj4r8hEgTptCMsnLd/F/2DLYFttcArerKffLFm21eeR4mw6Y+Dhxq
/whh86p+8Zg2OQ8WKGh3YnBUe6HfYWDFIYIuGyCNmM8LtghGFldkbuHP+fwvxThR
Ku/7z3fsVQOvfC3td6c8mncN1cC/P8i6fM3uL0nspwTqAIbyzS6Azu6PJW7Kmojd
PZkU+JXIjtYXMZJaQW8p3EO8HXtMKVkrcf6d0DKkijID9jm3a7TGfSnZIbO4hHfF
OCD6oPy02q7OIFnP0BP/Xm03rmvL+Xw17hSYMJ1d88kG73JeH9g3R8+lxxXbI9PZ
7KwrnuFy7bBNKiqr0kzy2h2JGGmNOqFUpH83WTRFt/My9YB+jKcH6cfqbLVzxKER
2gc5Qh6bGolsf6PeQpipi8j+bDZ1FAwZO95jRBkecs9qrJv/XoPaw90MZJ5ZghF2
r2MXIC8f7azj1rTjNiXB9O7RNEcuOrMtKGEwt1UZuRVH5KxXbCs/tzxrFq668woR
aLNTOZSB8fvM6kkewV1iDjywUNcrNrDg/hoDu73UIEHKEVa8RfatzwxYX4LZjOg/
L0/Sk98LXkXEeZhiLKAcbQyNqJRs0X+7/PcdIF9fKfwHNOfhuzHyueEHlSVHz9kC
RsObYzm60kr5PqkBK6YYur04aSk6rnl6KCI5MRvxowZqVzFZdlQcdsfh5abZtYUk
F54ARs46yUJi2ZM2qpMMc//2xx2siakCADbnQyKUWILtlNHkahXgf1POlMM62SUL
iEKUlKhXK4Baiw7luVlHpAW2mtXW1wnBzapppqiornVSGXv8Z6BgPdboYp3qE5ec
+vLuW//hTpXhzOYxymTFLUUxZIgDbKH65yOI030ydsKMoTt/G8mMYL+CbkqGThrl
YqH5mX9GGDyC/jeSp3njxbifdDG7grxCuLqMay1sHK3MZWnCNVOuCqltx9o32z2G
8Gb6G3/kGZA5uXkPbnGTUFc+yN50FQWgr5DY92fmy6EtnlYWNbq6oQO87oNT80wK
lSRq3hV5niSRb1lIHD/lGkuEBN6zjO/JmT+u1jT37T4E0cEhJomL802hSHmQyXhc
fJm4CzE2rgqtdVWOZNdaPIRmbO+ORlSyc3w9Awdkljz2iTGI4R4ML/HzDeYC4yAm
z9ooLFGGRBuOki3qXSKdGgzUOl/XdCKBADBc8LOkU4tavVEmv1BiD8IHExYFTDYy
TAc+OyOoc/HafPqHzjJe1w9SUKMcyiik0L662CPhj6xaT3wGsT+cF4fI/zdahx68
cdBUxBLthccMWcovyTMd0THGgZxbQocxyMAv0/Kf9wRm+gGLvUe8KK7TvWcS7q8K
AOHia/lofBqcq3YF94omT25vM07LbayV0dxw5S1qrXv2dtDiXFSs8YyGvveEZXAd
Pg6L/c2v82VCOwzXW2tBWnI8C+DGI+FtFVLgIs7wS+m+zsgEseX3FagxeiPOiTbc
MQRNQCpaji6V5dHxvecuG+YUSuWcLfCT3CdWrbfA9JkumZNlxQkSsvlpzjAIbBMp
wibr/CQmwMPBHRBYG0JK8vtFHd4lp19agQydnPDf+jT2QSRpbMy+8/AHn0xyjA1q
jQqLrfdVi8QBoBLQc5CecGnPMzr7CELkLCQCG/dTwJAbfFaELXECfOl3pBXYr8rf
4rleGeB41CoBUqjRgn5oMQqp6DLD6tZNG1o0h5qKxtyZ0JwLrF3PkPXOm8hCWrQu
B37/W91CLNpNGBey4Bc2PFaPw0M3d13Dn8KnOSut06mZEI5pk1xo+5DFuxL35syq
nJtxs5k99caNJoW/QAoHni8Kpj3AfllvJIgR5GaUGNshj6FTWDyxAsv4qsHBTSnk
zzCu6Y7+Rr3EZCzyXsOBa6l4TqWh99nHBIuCClcF/DxR0KyWM6K8dc4b613fFnxZ
JZuqCNdoYCjyOh1CIcHx4SvtNDosi/8+s9l4ufHFcITJdRaZbDEtADW6NslV0m6U
xZ6ShuRvfa+Z1RyTU7xRVZMFjnLcFxYWAf/9QjSLjqZkdnIIB/9mK7cjvWmS8Zl2
hJhoTMwQcGKKXX40CfHBH+u/HGeKjRbJ7jxlAIdDbequJ6kv7eTIxraBpndpb6px
eXlH5FGIIC06FBleY9rc6CVcgGDtbU+YzvEO6h12DPKXaOyEa35xYG3l6MhxEOmX
hB4LtN9QgnHp91lVzRgJ3b1UBboMXJxjX7scjh4a9FDstG20r0A1JNXYVIibybqE
3DKrp6f34zwXEFxpY6dP0QiisxjY/jnKZl04PiUxgb2a+jCKaPCry3TkXLGaRTUz
tOz5Z7HeGCZl5vKGQUTLLkpAaQao8NnmCckdwLABmHex/UgG646A7eG5diJ5wmpM
F1RIlE1tMI1PzmxO2C059/u8QXtsRTNcavx0U1Wkk9bdw2lt7Uga9h31pTISEjQL
dhGQ/ZBEoFV96UFwGxgF1g0Ieh4nVZ5pWpuqfqNYc/nLDl4gV9b/9c2F2ILArS3r
CgX036j9sJo1JpOv1i0Nz49N9J8GML8hQARywoTkpgr5Jj1cx9DUmlAkBGlmoXFl
efkq7CLceXjrn1BZF88DmwBkoY9Q/WFeSkoCeMK2Gvq+1U32+j67a9DcVAZjtige
k33roQypwLOBO69EDbdVluki6oQ7WJNFw8aOhV9c+9nKfzfghJf0gcWz2TEo5rU0
Sw2SMB1eBRaH8jFvm60OIDeeAXegN0gNs1Hw60aaTsK+UTyctfiyB7BrYp35136J
BRmElCCWQd2/OgGo151mk2zv/ZilkwEiz3FZt/wuwbpfw9fQEhpo8O++DkRArl1D
HmiVXJHwazKCpPgssKU8va3RhSMA9rMF5EXgk7I9qT3TSgSpkL9eJU0BHMYxjaFx
bs9BzvQ+KxRtRfA4i2zDP95QxpbJi/gdzQBgUAEsIsavIQVJi99Hk8Y+rnz0Twu+
uLQ1woapOd6AbJEof0UEyqZsFkkbLLJ7ETRU4ewCcKxCVoHVH/l8krZaw5UT3QDB
YWaaiB0IIUmYubFKLEyePwHKg0C00dXvJfEGWEz+TdIpVqm9c+UOI9WmXviFHxLp
digxtbPb9QyxTWirALAvDyG9e+vKrbQH7N+FaZOu5bpcFS/dlRTf7DLghNaKw2M9
b6MIeoBLXUokoqNPhlHbKqUV6Cgm5aipdh3+X08FnLBuj/CepCp/uFrCM3eaEuRY
BRnPie0BwdriERDH55mJegXY9flgk7KNVWEq8Gdc3RkT9tBigv/YQssjkDfCtoqm
1+Fuv/Kbf2uBrxm6P69EMedo+tje4sJGdix5sIK1QBlumUlU+z57LgFGAYy7vySo
3NUQ45EEg2gI2WuT7uB/60Lyh8notUzfzRk8aP9NEOjgdHiP+Ixgj14XCpi2+KTq
G4ZYMl6vZrRgCLXC1FoI3xU/yW4kGtIwRVvREQgl8Vffd3JOYF2N7lhvoFLINCpu
s0rtKzc1X7yaoCaQz5EdmTnrP+MHgK8jpVNcp1aGhuyEhOJ78swZZLUFxuiXaoVE
xOmgmPAYND2LoM3tTiSgF2hZKzJ5ZEVt4WyIAPXWixGz20hxTZFS/iycZVvjFFtw
rG3DcHzn3Mb7992n09zLcVwOQgIiSNnvN/ECojwtfR6+v7WhPmK2NiNZhjQOzRM8
PwPLbcTtqLZaDUWIqwQHNNS4OjZdKfcDPx2dBsguiPyfeUHJi5FtMqlvaa/IVKYy
Mi/NXkxRMG7U0Alzr7dRTsZZDUkknaHz8N5H0/FviCS+PDpbVH9ae7kX9mBlvU1k
XgBGYGOYDZgrtRoUozZxPNzaUgOQw1wQeWGRfgg4wTBZ2GhdBs3kR08YqZP5ApPS
gSTSGd5jajHuMZYXoPsgylcKdDDDEVpmvnslSx6tpZm6ZRw4YtDAehTL3q26rzYK
kY99B7CftjrcRZzWO2aV94wsv17SDz3qw8KaRJB/40FUjrKpFGU/4YdrTS9AB6Of
bHFF/sQogDB/qn08sJO0mXJTdvOLYya1bpsVmFujFVh/twRJz3lY6gfnF0YC3pPy
QdzHapxy3Lgxm8Wyb0orXadC0NLAv0hUQmQy9PoeyXDGdlVFec40vW7o/RrPvoY/
GKXuOye/thTaFymIEGUT5YFdyxYpT/qcEx9Ry+OuNLRzxiNbWuTFkydd7je4VMyX
JwgZQ92uVrwLfUwmRgD8Nh3qSwB1LaQJAQ/DACzucIm9uHv241tTWvbOe928SN1L
ftgG5/4wuFsHhhjoHf/V4m6BKo4qbBw02lucDBiwLqaqrOaqRtqa1C6c+a7uE/um
HBb7b7AasR7rqyvCAq+BhyPUPnyrPRaTTP0HpYSJowgc62/PcQJJGEla0fw60KIt
YwRKJShXsXY6b6gaugOJkCDFujeylcwxrXH8QYrgBOpwtnNbW+aQkRbIcA9BHcd/
If8AcdSUwlfjALb1UY3twwMAwThmV+Iye+G9lL5puwUcw/aMJaZdv3X6I61wOnbr
KyS232QRuge//ByJLJoJ1jlczcFCm/pIbQrlBSJwZWL7X4iftAsJD7V8nbEg8tHF
bV35d/9gD0Xj+nmt0AwONssmQ8UdeT6+nr2ppBxm54fSiOxWRHLjtVEbunFldwRI
kAQ9XC1VOw47HJwCcfJJhLAW1eqv6/DQvB5slTdht+Lv4FjCbIJLUxQO+u3zpkr3
Vhw/asFqKYBSURxUNYMmRpDdjXkh2ded9io60BwrayGeVvK8jVQZPeHYM2my4zPn
/jPuYos1U6YSb2uPQN0RFGvWx9DLIbtEDD5F0KC14ZObJvyWiwDPpksRg4iZZuyE
Ptz9Hb5clqJWFBd1JIIj1IwzFH40f4of0KONAHGOis4SUNCrrgNwmU1n4FMKBHFu
J2/lzqMy/56loao+rc+aJSi/PWTtDQhhXahKjVSqJvB2VKtt3OEU1ln2hKPYMtra
vyQ47z+440kX+erG61qGZEyPZEu+1LtXiNt69PrMUuxJrYsR/igoD7HRr8FqVyMX
kEz5qKo14GtDakGunSbITCQWIwp/+sZJ2Sy1LBXhEm7CMlKKeHeu/fQGoXoIuCdI
QUnP72OjxsY/SfCON815WuQ9cEifMspG99PaDNvbAg0NxZG84lTPF+t+kbvOajyR
2o56Z5geli+MG349Y/xebmy+dDir3oJWsVf7mRpLjrOgxBZv86O1ODX0PA+1UhAv
HpLmqZvZs4HTZ6gv3/CBrcW4ZMuX3xb9HkVdEBr1tfxCiTwLTnOrVENw8lEx3cDa
+YdP6eSmn/6Fr9MFp08c7FvcImlyR8dXKiZIi3VI4V/bXrluLW3wTzstaF7tgjpJ
UEyDbGvUpFGRyG9yxKU3FMFf32U4XoqSrq/Wq8/PkdLIxqOMB1xvlDvV8I0FTC1o
8XFLKEuvMF1ywpg9O9sz2x3w1Md/Em7nYFSiFkIeUe9GJg3yuqveS9L11v1VHmXa
st8UVK3NEJQDS6HdroLR3bh0IRdqm3oJH+1C9QtvtynMTAu1Hg4+be3ht3xUOXQv
+e2q9peiKsviOq/bGffjnwKUiK+peKXTLu+/7BCMjMqM1NzTLjLigFmBkBPWRhe+
yKD3xHe9KZcUjnroayUN544y++hDLt2O7LvGm8KfGmwQTSjLInx7OMB8pkLMEzRt
+nxv6JummiKPlsCogTuUOXDKgHDI4+ye8+o5ktJtZvB6Cou+h4/eQdoDR5+5qyhT
OcB8kgJOQqJhG1xNh5D53rUoCZZLucqdlg5G240GIsL4sOuBW9da2Pdaq12dm242
eSiQ/0+OHggAATJSHBhM/WVuIORHZMadOQR0P3y3DFxDN8DFu2PIBhKlK308IBJg
xs16QNr9we79y+RyRsjPI3wkMuVwPiAq5pHMpt/nWHKcbeLOv6RgJsot+w9rQP3B
nkvy3acJYRheoDopUc8wSAcDmvkor8UmAUp/hi3ZcoQ4azMrZeOPn7E+GeFxp58b
dF63P3T9HSDQ+OcZjPXerHc8Mk654wc9I2SOdBGJhAN8QyXiC/A28HUZ+4PVYy+U
B8eZ8VZtrDdGm2SdLlZCdpoBx36G2U2p4GmkgnlS+GwYBfSSUDkd6BxJpEYgJyDI
5NulxVW0S6qwbpABYiYWFTe00UfpSEzpgugbAfJyWcyXQ/ywNeL+Mjk6sSjjcawf
cU5lCEYFiF21B28bqV+G7AfejGDK2eECymcFPr5/CSNSnJB7ZZo8tdk8BZy6kh+w
kqHihLzZ32scVNl1KpOgtApoq7H2DJ0jmfec/9fTD/Qi21TiCzUkpNcl8oJ/cpn0
cCibgSmmK10LoKLK7MVz/2zCdlAdT4bAJyU6oGNBtID9ho5xZffQE0iWKIC/G5yY
TgZxYzqZGrb0o13yf6JpSA7dXbZM7jq+M2QvicK6cz/vTk3DfkR4NDXPq7kCimDi
AIovj7V48te3ngf1xeutA/n3RcBL+erY59zMhFK6s54N4irIcXn3siCYcYRk0N4N
WxUbFZ/Xv8xmL96f32hCrmqn1ppbTjpB1hnIdaB55brwbazsGhPldcghmob/PCoU
afQ6BI6FqYLBH8MVfoJ7Zrdyf9x5ozUJhJs7ATCckh/1k4k6ACtWQ8P9PIEHjdQN
maYePcjhpYCUckzUIkIrrj2CADSWbPpgS+ovJqjrUX83NaPiWto7vUWiZOCtE0su
Z1wG660evagHsKtYiRweLen/nCqgCqTDkb8TQitccYqtuyF2VK6irzk5wEdB4q06
11BBzMGzyyT1aw/6iQUpjBl1xzw4mmJkqRd2XFEiQLhrukuFdodnewxI+2gKDqEn
s6TNlaghgiHGzQJT6BTUoMnKb/anUtRaR7Q3V7Eos2s9Ofq3G3yRd80+GX4vzit3
wTOZw84JwUQJyb2IOLGzDFUIwAn/OsbfXwhGTBMgIAbzueAXppQT/7VfCAm7ErsX
RQraURCoGULtdellb47+TunSUswN0Kv5CLJGf0RghAUMnUTWXBVUmZSpJsz3nYVM
khnrDSs5eqTqkrqNz9K+WZ34sPrx5P+fvuYcNSRYTG+ZUqfmtDu3wrKzm9+w3YZv
tfRxXysj1Tgdcz4z2udWNk83iEsrDCIwyV/v3ly6xKktVNtfjw2e18mcB8EOZt+i
KwU+occ9s4JiNtqIvMLpsEhPCRrjSJc3gfpkWccLap2Y4+/If2x5biK1oENqzA5u
9fNIrNKN7RbwdPrZoitAy5BdOnf7nBnKeGo5qIrW2HDRMIb68TIk+Qk0qGb2MigC
LOmJoGvMlXeRXB3zHXT6yqOXZbmBeS+SWy6etytHlC0VQN5S2I2O2EK2U1GNZLCg
4GldXGB3xRYA+LxQa1uMx5fxTMqJtlz/ir5TPrnX3hXpPgxWUnlgq0+IKXu1/EKG
eF/pfoIRYjItRHuHVDObYjuog2/hndI9caTI9Nd/z7w7cgsoOurBpqG82UnnW20z
l8ieeVdIBX1/D0gSsHNzlsyvzHAZUSVVuylgVBj910upozBrs4g0DjbjLAaPVMmj
eikRlg7JZ9J3MN5AotTtiMDYlElhMS+Vj13yWK35WAN/FxkdxzzDq7c3QqIPwMDo
CkLrX+kLWkSsx2nWyM7XmnNPdPsB0xgisV1qJo/XzHjAY6W20fNnsDViz/HqPZ3Z
6HsWqjYHnadjsIMGwZ5TUleYYjQpNqPjRuVg8C+ww2OEUeS4YzAbD1odmOiLRmVu
ZlwdDMpmzKfFsqK/AbTD0AFyfXXy+OaK665zI0Cn04y2p3++uTJs5YsV68HXrC0X
v7NPg7VSdmOc294zbUOJbuTCfgrtHHbSCTQxMuadBXrCEjalIb0ip7+Dnx26j1Pr
0IFfm+TCzqwt84iQflz2QgHsKalWJ09I2bzx1JrGpUL2XLVvr4GZA8DBsYMg6uts
LMHiMM0C6PWTkwYcxA0NhywA6XwZ0tju9aUWTkAMB6of2wdU3F0SMUDyp0ns+C2M
FQH8EQuq6h5VIpNOlEyQZi0z9goOVkGh6l0qgOJjGGczssdjbFMzlW+cX/CrvbPA
VkjNDQuberPj1ev7nGTvYTZsGvfgRq3/tOGpJ8LNJxANL8sSeTyyfyxHRnjAJsRZ
a/5xkoqXUWeKKrzsx+xUR751BbbJ/7OsF1w4Sz2zyLMIw3bcsQQzcvKsgWL6f8PQ
8cCM4VqVWc6nHTBsDvYOf6/qidoTAE0qsp0BzCi5EGBGcThX8WPWkdocfmjHWU0N
upYMX5q+1FFsn7/SIwseyPbxCyFSpH+Vi7/HF5ggU8gZFneVcpEe2AU3IXsk3dBQ
07HYNdkwifEwQSSAomCWbEk13A3BkhAkofP5FwPZ8v72y49yr4mQuPG5Mb9jWqUX
OczJ+CYg9paBTG1qLXCtoCFztLnPuaLIufewsnd0J3YiM7n9p0xngYESHHF4ByIP
PPisiqFL4vDqBH9zTXGzO+LMtAxRuLbmhNHw86D0S6P5zO3VVYzci6sQG7DefMEJ
ZJ6rfyQIhsk9gi0s5KHoK8CvN0WJe5mycfrEOiWmuo6oRyiSqYCklLzprWOITWo0
XA07n0vIWhqtlOqB3kSufgJVhPyqrDeOF33iUmU6zEDHiIKr4iw8dOFwQf0SnoL5
yfa2UXSwoyyWFBimeSJISw5AK0dfCjP4RjetoCFl6F3kipC5Nb0P3bGz6s0zOSVx
/JdSlcyd5kLFN3c9NY2Apmvh/C/LbKUeAdKOKdgOAjk6GQDqj6PItmF7+4v2w91R
H0byPwoerSj0SDh58/lnwRtQM2RgN5cgXTZExLZ7njsV5Xj1fNc85FqeAcFVnx44
Q8ydf1fWfIxTJxUznoCp3Jp7t6XjJIobV8Pz3R4q4MPVVnhwIr4+wsUz382U0GgX
mF9edc5Awbe4zKAwGaG1gvb3NrhOd2P3K/UeBeoY/8UASUSaPMMKM0UT05yYVVxd
5yrnIGoSstNEwDMUdkyzBsXL/WMOSTOujnTx2mYwnyz3lJfDRNwNc6Z/GnFrSUAO
ALC8ECpBPkDydKDM+Ccgkw6vy1Y7bB9g8l5oIboMhqmf/kOj8TQj9Tlu5R7N4SL/
GlzQ0ITHr6sXUGYnbdb9Rkt0H/SchiG4ii/jzk1582VInB5m9IyBKIBY0OdW2HQk
ep+7hPKtczWNwaRnBVrsO94lXRPIbYwAkgk6CdoM21HNn0+Ri5C+Pw3rn2CZc5lF
gUvvRZ8+scmwYaUPSq6tn2jl/7EkEM7uNU5mHbw8xC0Mxb8TEqY1sqUbx+efY9BD
/GzyU2POq6svFxPfPA+rKQ8Jsy8vbpXUHI617Gueww1zC6J3Wg/Wy6gjgQn2jLPV
Acc5EQ6MetN7YcJkJEQbu6rPmSdnqsVbiDKZyEeIZOpzT8afemXrRlvZmAffe7YJ
P34KMC10FMYiJzFVbwJfelh5JXRIL/6sSPpZHUs+hST0hWXHDAcKPVJXOlo6YS1p
wjFlWB+vIni/6YXk6DkpfBQY1XiWFAHVeGMtNoyBbwfHPm1gyq222cMLYuQjDzyv
IkVEm+Byr8wvygWtl3u/GZaLMliA3FtPhzqCcDllDTYmOOvQepyEzlVthWLa1qmT
cZfrhJILflS8wuVuge77mFIkB9rNVal7jlbM1+G05a+vChlsXPaf3DEUis6EEaai
aZ5LlxSE0tcFKu+NL+TGfhs6T2w52vPxAUMs8JGTM2E80/L6++lXKqqXkl4LqUSk
uxcRAEcrThFnFnI+iF9uO3utoJqvQvLL1sD3LlMctirNU1pkInEd6RzRJozuSMOy
AVNg1gZLjIK/6jeiCctsINK3ao8aDL5p9XGdO4oeP9XlzNO+THAX5Nv2+otYT0hv
+VQ7pcKvTeSW869htO+EqT72PSx8EZ2U7MjLM4QnD9GUS1GDbm0xGK/vx6rkB+k2
ZJsCwsLjJXyAPePup0srnBACmHE2jmTBwMOnGAuj8WGuU4QEtbAQzfvE6NCleUio
dZyqm2pmDpH7Jnwq8FYn1jrjOI9H+n6zE2RcMlMxX4BSNCA6Y8WETdzqnMfqewBP
KuVPoAbwTmdJGk1Xm4LW+Wk7VwoaNxZxVQb6KRpy77lBsjYVz8+JSN9x+loUkGqQ
TctgX3qql/kwJhH8IaDBAcrU/RyPEdKRGTr745hHejkwYzdbqF7NaFMIa3afmQzG
Dc8W4E249bpPPkTpTyaIeCQ/QsuuEzUylH8JtVyUGzpt1IY9VX7HzLvWbwG6R1GL
hr2KZynOJOWQIkuOOZJwNG+Ip1j6Cbqr0jAEuOuqrXw1zzExI9JZwTdy4lKV9tjW
oKrmtrq3sPiKPqZJU8KFpU2phXrYW5SF3Uw1yuegBBw0f9Lz7YB3Kb/ym0y/3UlR
GSVHg65jnQflckcD2Pt8GKf3Gge9IHe8HZn77Y3z7zpP/1+LDd16xoR+QCfECG6C
pR3ynMgMGzPu/OPC2hl0HFvK1eC2DcXP+rC8AWM7PyXeO9fbz/+sO6Kauu/zGZ+L
cmrQkb1tIj09HiE0EUxF0DSKcqlIm5CpZe1VakUUUWCt10V7G4tK4nIkdktMOQjN
5OeA9sT4b5KX8eG7CLLydDNm/TdjHgiMcSAHWK0zGmS8xN76d0EXI/yE5ettb6bE
NFONUEFs0mhCIwk+vrSYc8zEFJbqVO18xkSVhb3oCZhScIPbaL6kBd+0W6dROfQC
i6H635w3TyQuG/zuosqUVfuFtYIptpEdLn+fevMPvHx4JSkRzQbfqHQXtsOOYY/r
UZQr3sPai++Z1LaNn8OTC2kReA1msdVK4KZ5a9S4fCC9rGknjNSZlwVqgSbUxr3E
YIm7u83GG/U5TIUaELBCtj9Jz7JOm2tN7+NjSRXA/cDe+f4QerMcSj+T+tnISn8H
QwHlj887bp5jAGboeqKbxcrchhncDJpQNUwjCcEwFKgYZIsAbzQslC4so8X3gpta
q7O2GWThmsH+92zgerrR4IIIr66oVjq2152PmNinLQEQbyVXMletqramEPbvWdZn
36QbPzjg+aWfuEtWMwYV6HAE5Zx/fKJIsFrEvjxuF2+B4kmJMkRhIgfcbb+AyAXE
MhUY/xQ6/zSEsXWeoQOkbCeDz9cMy63xKf2sosduFXNSv3qdoQW79W+wiqk/wjyA
BvMbHiYKQmWq6QlQF7Cn3NDD4UB70+qQ/rvuS3APRnUVrkzU3fnERYzvTvX9jFq4
ETBVu1lCZDX2NCIdQFFZOxs/nvDwLY1r5K5BrfqM5IN8qRF77Mb1q+Q8cw0N9jdv
JIFAQS+7aQZlZ1aDMbPzBlFcFtreR1FlTHn00d79tfl1xmLJbvbfvXpA3j2Ddiuv
uDTp3rlfyXASPWRSUcF16DJ57F9Rpv7l/+ypw5m94POcywFvHPn5uUnrIZ2zxl2E
J/YroK90Dzxu5J9TzCNgfMXFh5Jc51ID8BO9CToJEW34fWa61309EY4V5amj8Pp+
qlB5Q0/vrRDb3N5N42qafe1ZxcOj+Pg3tXKg23ZqeuKWiNS3JwuvG2oLzo+ON+ZQ
tw/NUlfDpwRI494kwhXryo7EZr0Vj4zsm6wrRjojFsl5ic/AYXDdJny655vrrKTn
FmfnD8a1vD3ScNVbl3XtmG9AxpXaF1d12pPC6DK7eLayE8eLfA0DHo6QcFqvA6dx
g9XK8VKjd6tjhDTqJ6nhohGZMA3w9Z2yOxRWmjzZYJ3KDUQJmS0eQZ7NYzfYEKYo
dzQZtgXVA5kpGp8eNB2FSOBE4ceUMQo2Yo99v/OR5aSH6lmOvTuk+PmycL6RNjjJ
P3ZhtSjokaJwExPkQDVGpyCW1xMyovXvc78xMkKCNI7zLPG25RY5o05y3UFx7hur
jmuC6ddVTfRN2iiiB1etOu2MV+2p12BLpYpibrmEqN6BHf7AtiH9SDRtCfmj/4TN
1qYiF61LbwSaAKAPC+WXb86dLln6WMfO0Qej8W6Y52rLaMMRpvf/vHA6W0fE7/5r
HyObqhRrp0QNdEOItUR5dePbUCIGJP/Bz6k+E3fC5Tf2foUXawPd68mI1V08khN/
PWvouWgHdNsv/YHefapgYi5MO7W7GxP8zJnZd56koDdc/6AV9cjBWuJvlJ2rsw81
2PB/InFqmPuj6VrDOjUgqS1VGw1olbnlhzCKVvkYc0uHbgazydehTy7aPHWH95Fc
jCxcFpzna4r+tDlL8zYqD6o6ydZ98IJppKvAnkhhp16AtTbzn6qwhC/hmRUI31O9
geee4CaJTlOyJv6p7JVTck+fEf5M5V8NsjXuxa2GWY7A8eEaFelupjwHxvtMwOMM
ywQw5ogJVGMdlk+hJTxN2zm/kKuedCvUoVv/hahyxX0QM/87FIS6DsQkV/2RT6rv
TcCuYEu8E1PGOaswq8Q35508SEGKt5nAR9XCrKVvDQeoBjwIBG/syQL1Fh12yuxm
Rz5J8Lq9TawqYxawk4resWmqcVNw8C/8+sIURB/hXFQZ8NlEwfYfgW28Kwr4PQu6
IGgsZjL4IRecWJbyKm/Br7gVk97yFnQHXbDREaWJmzksWefTxj8JWwArOLo9/N4h
Nw1G3BjAeDQFR/b9FsPeWVrdog2f6A0F57myriTcCeDAuJHZX8DjCgBA3yaIWNJD
pn257K8USepy4TuN/Jiok9MnWpk4eWr8jKCacjP7tSIM1oZim5z68Ae+ZrNSmS14
0IkOTe6rdVRJScCS2lQS7ZF0E6YwpXzNqNAGzU2HC6KHfE3FLuS58NzCtuiBda9D
VayCo3R65sglktyXeyIin69T/FAbt42JXBq7kOp1H06Z2y7myl1o9F3S6y0PUih8
UHLbjp7jDbxUv5tEpHXBakvW8kGQofdPVAS4VbR8ngRK3jwuJFtiMP3prhrlamxr
dxtqWcLxxdrhKa+QHq+pPIWAGvisAjsFl+xtrxtLRHkcScDM7EZHjmzLxx5OIkV0
25aBpUV4yhdbuOaSwLoCeOHyIxhaXopeWmXjorrEc4AeseWgYc1oijScUX9bn5PG
9kpMvBNzHev8PH/eHSZZGU/sguBR1jNDW9PA2vftjAg3+YItIhG3+H8Xpnj2GIon
Zn77ULsAalLKFWmUZAb3KntNjqfY4m+AvYT+99Q+PaOjyzZcZO79fZTCzlozZsRa
zAHhGMNrVFUfd0rKYZozQynxbWspd4vejXHEzNJVHXTJbjFYAP8e52su3jJ98ZE9
LlypUuX1RScvaeGr4KdTNw+JGB32IQmEaYVatzdScJMOzy276bdULudy9U2mXwjB
N8F201xw9CgzrK1a+SMtr32Z8gTEjsMLsyMKxPj6MWjZ5hEkJ/ZSc8ATILltWeLu
NAqcXz/FGijjO+/UORG6cBExW4UAdXDPlUkgXxDhsx2ZGsRE3YtuQTbhw7HNmYcT
TY5Vd2lh885yuw9/J+jLdY/ZRTfwVFWW6QD6nBBZka6w0usu9EikPm7SfsPaTOWi
69ZnxuUYswhmjn8ypI9Tug18Svz4eE5wckdZvhukDsGgwT6KXFCapXgy/JfMjob7
Yz5Qb0bsmKW9EZGcGdoP6xJtZ6mDS6fosDbfE2iDMrCzQ7UhN6ry9pOkyQS7ANyz
ceGfhx6FHXWYirFWngCTs7lY5je8vhTiMdPZ9grIfmKOwCyjKLMXPf7hptTiaNjR
1DGLoRl6y+/ndAXvC/R5vCYAWRrpHFtWJiYDgRAjJHafCgLh0CB8hLo7DXN4ZCPS
3j2oKeA+B5bidGNZeTgFN6znMdU2bB7/MZBwUHAeoPzAQCcvfsjQQOCjTqZU0y9W
JB9dmjmKDoq9VdCWU4LbBeyksuI6crMao5CpLS+KFFWiUg2CLYcYLldZd4FnFrbF
6MYj9LD5E7zSsNCKwGgi1JMZYNTrNJuqBji6/45WFAmr6o7bx6p4JNJrxLDZClYZ
uUzbhg5/5AEfLgAEJcrKDnkv6WmHNVYyeY0jCQTugEymgkCWQK57ZnybXzlfQj2u
R+GkIVG8dF3ITNxseNp6DBqmcAFxl7VDHuXzA6peJdHfgXk5bL6LzKv91d5SdZ/E
Om1x7hFxqNFLzH7C/YfYqL+W/hNJOBKz8XEaWVGXvEuxgEkf7APjDQ+K9OwS+R7v
dP679rdYrVCguJ0dmvViS+JCJGQtGZ9qZp5Ec4VlGJsABO4RgFTHoVcbVC4nkxC3
kDN62g1ECvhNisXAxz2ZIQY3Y8kx3Ye3kASXSHAa4/DXs4Q4iZz6rN81K6sB8ulR
up7ysoE6Jc7KPiw/kwbOiErkaNT42CupCYt5UjlxnospROu90rFmogQ89o1SamGJ
Y06XUowVh8DHKc+AiwPmKG0eMO2hOBr/28Gq7OV8OMQ0iBxkX6qK7OW5I/tWtiu1
ynZO3nydqW6SnThRmoMcOONBektWqPeP+3gqlUt5xmnRU/KUFQqkcA10ZovZHlJT
dpDg2ch0+XzFdIlybYtec4FNnSPz9nTjBvS8DTHWAGu6Tr3306Bzzwpm2ewUSduw
K7HlwLu84eQCz938Bbp/eIaCenJ4jwauoJEADhG0TQQsOQJCjdmSZ3uZHTcPJ2gj
CG0ZHCo45xVn+yRurjbE2t/vwtXXh3TUJEOF86rEKvffTojAwagLtwq5QQPtmPBk
HKx6bAC7m3uvFmkHlXrtyny0vXm7YiSr3YdMKR20+tvsKKXnRv0hztZ5LO518JcS
J9Ulo69d55dbpgqAH9i3OQqj/6HQSznOovL/8Sv1rE6fPPD4Gex30XVHTGU5ub3C
oLS8jSWFKMQP1gkOS6iqL9FMRbqWt0zrvnN6q6Nm31H438BKh4kW8OqWkZWDnRP1
6b9gcFL0TFCuVPsKfHByTHLa9NJ16oosDt0b8qbIa6ecI1TIqhN9cQ9Lc5HYAy8F
9l+bFqMHtatWaRqFfWS4gCAWKaMzKjVZbnPxwI0g0ughOM9eWiZT+dD+DDvzQPLz
r5Wbom7672o5WXzZBR0UbiGEZ8i2Nf8M0QhpxtNnU84Nvj+I+yn7b2kQom5bOjgJ
zMgCgztP/j54VFCeQ8pPyAArOzuhScqayO4x12as+gTXczVWRt2Ji47uwxc70Y88
EPZsZjgmYcl8sjGHjkPgMwcfCuHX4R+iBQmIHT+laxigi47Wsacev6UgvW/LFIw7
WDfOvp2bHHi9NOVGcKMBrpakCm1BP0j3ulfPNB3DIyYlqKCkAc1Ch/dBnBDta6n5
ZJovozrM11zdRm6juIzTmMpzUUn7T26TdF6W6EEXn7off1AfKH4Tkaa9j2qfHi3d
3qEeq5nE0OoRHDOn+4yeR5sqURL/fhkVx+14Sl8VKKR71Wqz+TvFMFciNPhDEGb0
w6Fyz1EwlVGf6cI+N8yr9xmrdgrXP/ihl1h1HJ/gfAWbukcu15QpaNLbMkwfUiAY
063aPCw3P4VrjxD9DNBnK62+J8tMj9ueK9QtFr0G4vpGErC/w9wjdhzwMtYH+Os8
brlbcqt+odvP2uuDFp7ajjkkVn7k4d3V5D6GJRVliQ7XsVSHqf01S6lsDhE08sdW
3xqhN3hbXWuAz60shK5wOAXkx3gfAwTCqlYmH3ryvtainrZtavpRr+/awiYwNaPm
cgqCckJqwZqHjnG8LUfouTfEa7SvyDHnjc9MzLwZQpTqknkcGt2gw8nAA9WxTJ/f
Dlcc+P+n/4qZ7As0ifKRt2ZODNHPjzhAWukFq+GzYkyLDOHERoLiq5snADifqrJc
spctlAgF+qVBlsGdrdOCxuveouIX9ay7mqTYIuDfWXT8MIWjPVATp9FYehBJV8aw
kg0H8mfWBqaTTwCJ1TzBTaTeKBafynrbgxWjwDzLdRBxAn/k5G3KtrvX25+G3rTe
79FBPSSMpijJdx7Pr9X/iars+CLoAIoNx7YCn3fJA36OqeGe9Vn/WTQc2/uZ3sKp
yzfu/ggD758dWhLu3Cv94HA7wQoAguTqNbZ8uCbSMzXLkYYLOO/NdsjfnAV8pmbt
aR+sVJOvIiSA9oHi/nmMx6fttXkqJfpxkyLGMthFpGMGzRtvDgLFs78SuX0p6vMO
v2CQuvZBLenbe5j2TRMtAU9ubrC1sHPmZQKQX/+5FxXzWeOcqEySWCUFE5Ye64nf
abG5FC/F9BXEeqwNmP3PEpQdrWglr70ZlMi5mnYxkxToz68nx21s4P4WtiNDNLFF
df1g2usM+wEzCVKFKXeUPh2goMeTbTiQY2J0kQLt+bSsaR79BV1zWvvxzhm+lGCp
D7yCNodOLcTSfkxyYKBzl4eG/wUtGos5z1YJCAuK+8GxwQOb57b/FLp3vhHjQEml
Bez+WmdbyCwIgqwhx/fNLzrNIqO/LVWbNy6ztCM9PASUYQD+3peMDRv4RnjuZgFx
c8Z9TSGS3bdex3furOV9gEBTjsF6oGhadwQcnt1/U+KHjdo1z2Wmu5kf2oXO0cWo
ayXjmEuqycC/5Un7Sa/+r1FLG71oBVgOmlvv0xr8sFZ+qZq7GhEEKWtJOpV03wV0
ScjZE4x2dj6+WnhGKxAnsxdSgfg2i6jRpe/8YF0bPAYbTgvLPo8WQCXH7Tvbdavc
MuLie3dY/MSX2FPj/gmml0uMPv6maLEm6AamdEV9QQRB4MqaIHT7HCNK9wV/MAPg
nn/Ft4+OMMjGFRBnOj+AiJRR+PlNN4YRx5uxODy/ogK9PP82sXeeBMKvN9lXUfL7
GNv9G0A84u6Q1yPj7G6rnjE48+UFt5Q8eHSmzTg6G9FDrTbk470d3Afze3parGZw
5Ng7FoG0OdXFFlc7taHlOsMvnBMj5SX0UHhJAEgqa8BA+67zNJvTG+yEvsbJ9hA0
JcRqoGE+FwgWbCCKreSGZGh6pRWQWAleF4R4WrgF0h3bBe06AYfSI8dCneEpQ88r
yn8oEyUfZIHZyJW69aLSsQOW5lZIB/yHaDXhuOHSuaUwkDpSrAGusPoHLdyMlZHc
0ZVARCoZiCnR+6BU/ePw8g8EC6onGAeG7MN4y5Ivay43rKcRbZ0B8aBM3vdSXPlf
o9unyd2InnsEQ4QRhKylmZlJtwQPeeb/WL+ZOerPjt5UNpXf1OYpnlidBAn0T8ER
qbbQnbntZ8rj8+FcLbh44EKQt3OdVKoui1YvqyuAuC23E+EYcDWvKmqdX5F1mCuO
sXZlhrKwxx9j06FYJBo7rJ0Os+0Filp4Z2zX31qC87sCcsQ9Ds4lVjZs8mWWZDwt
01f+KZ5HFTQnKHI9VQaFzXEQq5CA9pqrfubwbuyO4bvsbdM3ncbVi9EHw2KqEzth
qD7qCeuU8FAPucdH0ZZxh1+hdzoNbb/41YlIAtF/mJzhY0dwUPz/w+yCH3G/1IkY
iHztpP5s0ILC3kuNfb612AoyVFjeH93fBxaR15AekhNbF3NT8zS2NzGVKWGRTLpl
lEKo0bVrRMybWE/NDLBo8zXZU2uFSQaNsk4bv870rWpgqrBq2dzJQ5WkFnUZdYMc
MU5tzFGbjAsGUl+aWqJfdDjAVrYJlJPczDQtxFBFQsDR2XfzWX+/Lyb37JsfFJ1+
eMT2EU95jtXQ1nq/YFHAJdX/z+Q2AfGOEe2lIsE7ZuD3t3b2QEc9Js73BeC/ovMd
M4H6GZOVl2wyaZ811gOeZi4csIVbrdvIxWjSVo/zNqO5ZVm9n0Yejgp+d39sdPmQ
8SaNSCx7/H8/ESgcfDyywSI8eyq2xzCiFOYx4lXxcXZBPfdvE0jJERNktPCEtoIt
pcnMI/fm7x+0CJ5GvRIJiyDhfpscxXOF6nRewMh8xYEU4wtmkjLx1BsOnIBsLetE
R8b52LF3EcRYgtQAbP8Zq36oQnAwdwxxcVNBoP1TXvwfKA9b889hbtjFaucxjR11
yV26nMahsQ92bDktpNTz7yBcyRswA5gHTt4IsGacbKHTVYVF95IBaqZPRtp2yuwi
jSS3mvB9Tv64FmhmPIUmfQl91Gta/uthVoTqDNjH2pLgPCJ5lTBlShYlOIzXx+D9
tZw5QRQUlmNCmaj4E7HDwEEitvi+ZtLWWTToXvwPoi/ec7Z5XSWPKIF2GCfAHFTC
CY40uOq5f8TBL2k2NvB7nXvljttkBGGPAg3g+JtIlLnOpXDavegIbZWCyoUweADO
PZGgoCC7kbCMX07jP7CfsnegGXIdCcKF0a0oQ8TtI1D0YPkPiSqY3Aob4AcQIZFB
SwCO8wI45O4C2Fo8g//e0ySCkLUxqdbDc/DFVciNm4NVPR2cqv0F+mItih0rOtrp
QrKSuZD8aqtgGgzEa3N7M3rASqk0vJiJq6Wlowk/WmSZFa61ECRAq5Y4JcS9hX7S
aLXGu0km8IVcRMchNxhIS+pF0EhOGV71+4zwEzU6HBbCa3QVTebHXL02GLU5D+M1
E95dquVeTWTobLYaTQpvDM+lrxKLWzQG65NGUmCIxbiLws5QgAXthxXEzbbQ/pms
MUmfNs6PJLknHJT03xfq2VO7YPekHmvO/F1JbwIqRQWHcjTiYHhDQn/sy6Q3qIp3
hB5tS8ZWCsQqH6S5iUjagHbmwI1MqCDTSQ660ngf5evgwDgEJbqIFheyJVSGaD48
PKVA7opMhmuRqh9Of0nfym+xBntuoZGGgoRQ5j4L+EChsKHPRWpG42fkfN5mfACS
XavQpHvG2OEh+ImIFu7MsIrbrVuRdBsc06NHkTIv9aynoSloVulmb6TyqX8xCPhC
ftm0IfCYoIWOIrRbGnPjbGEaFjy7P/hBAiZuH5CJxEMCiUbD8bv77oxewDaChdQh
oK9B1CJq6AMW4n6Wq5PSpRxY0P+ko5KxsFyNjAV80pQMH97/4sTMv048u7R03wy/
bx9efrwbOYetuz1rR1EkzGue4c5VMrFdnPDij8tn/ESDnZ4Opl80ZJWNOaUnhMa9
rJEwCUh1wmH4RGumwTANZC4f2/gzZmEI1idKKPQhy73sIEZwF7X/RKouynlXYUiN
01MRYfs1zTdejiAaxqGkFGxvnoM7p1/Oazn0NgTUACFKffsGFpFOHalw4JdedbiH
kgkvT1NupL7rKmGs5OSTWjBvggD/4SAug4LiCPJZaEpUBxKV8CsHO7hgULxtmZsM
Qdd1ILQHiPXLHFOf7yMkvau/8r64NJUSJviXrmXUJZzj5uPtnH+GHxtf/gk05e4Z
S77BZVAFJ5DHvcdfLGriLwpoG8ikj2uqmHNV2HR65cOayhqnzGGUypcPDxo2c6cy
xaAWPYW/OMC9fLhTRC2kX5hGfy5Po8zAmaOR5Ai8ihg0HUoDUOQQfpFEkHLmnDJL
GDVdl7wtr4BUXuMvKFmr04rSbP4DUAIq5+1NNBLIbqkLDxq7nhwu7QiTDVfoj4tW
A1sH/ce+/Alth7cB3ActR5u3imGZLMXYAQHjCgDQEeNgqgkcyMrHfHuNoC5w+lQ0
A4JNgaRFLtNgmwuz2dzSu4SbB1bmakuOgzOUYDtti9EfKyoEx9eOoNxM8uojkTCk
52Ohx0U/CWPVHmE2cK9eWdidq+X5uo1pMKz3GtHarEddOpcZbMspR92e+oVuUrXi
zD/ssH2x0wFiYJ8oftot3kPPbqEEMVTudhKrD3YDKcEE+j3PViT8HldL84kxsvQF
E0nsrBtHhAk7HgiIK4R1UtzF801D9PAk3CejbdkmsyuRmz0ktm5n/m0DtPdkpO8f
GV3f+QpBQ2000tZX/i4Y1sd/XDN8Frp1KidK8HhqmRSs6IkGI4pwnCsCN88Vquyv
C8u2+L159Iz7CyqGew632YoP8fdmz/jskvy+yHGowzXUfMzQeHPuaccPbZJ/EwvM
EA0+ru7Di9802j/98Zie6BiPSCkGPnVvbPkW/gjyfxuntdGzw6XWnEgF2RXOoY+D
coHWsqQrAnlKHA5oRdirsD9sP8VFgpCDHnvO9+BrkS76JlR1iZfVrxWnL925Zn00
4NdtCQBQgCpu4FUNj0AUp7WAKCedUCMCfBd1wsuXy7gIKQFyl6vM+ofbj3rxGEa2
6yBbOTwZAcPlvEAcPTL+sgdonyNfLAZ3bT2gh0iYsJO3ptKYxtNEL7YO0Nd6zxIc
cRgXzqfw5c7OtsBdgbxJK+HGrwhT8l0FQzRQDyqnmcm+qC1lAYPkw+hd6Xax7tsx
93iFdDk3OGhkSvr9HQmsKYgDJRViWcMFA3eEbYn0RHmoFx2XDJOv1jEcnBk3uxFT
qfQsSuVxXhgMq0v7JZpaKetbwWw44cBy8QPBZPtzMZLfEvwL/xkA+8ohivVMdi6P
yCZiUtiL18RlBiBkJ4Pv+xANDUp4y+/3+1kQScnkIgH27/9afA2O5kah4PYrPKcU
jha5yb/wJhMibLlBWHREiGFvY/Bi6IhgcurjQjx6NrHAESySfpo3YtbMFN9+hmL+
BtyRY882HJQYjBvVUhPK4mx1+A2AmZwPqygmXdQ/jPJCTlSviGAbSrIXltVhxNbr
IR1cHx3X+uQE7lVUi3bwrFVBTyXeduOnGzB+WYbi+4dc94pgLhYJnyRW+RpZJJY5
yY+0k1VCDGXzYxeYFmSjCK0kWwK3SSZ6gqfJgEy20j3b4RUqzRXg/qtaWqm0dAVD
ogpqFrFi/Qgdv50pxP4l6mihpllWmK5gzDmAV1Y8L1XZ36fpXhHkpow9J6ZyECVj
2tfSURfq1Ztdcx/NyI2Jy1rbC7ji/J3/BOK+s2Bxq1SQVrYmHytPy/wICqgPP12C
LUxQvG+foINVtFdtZ1e7YtbEOpxTOLtltL9/G3K6K9y1NWws28cnIXTvjTqeyCQO
O2Zhz/R2PkBqjoB2orfW3jjiI4zRb8qVcRlbosCPirUtEYM0KsTM4rfR/C5u6Iye
l5MR4Jpmy9RXgwaEjajoYaTGl4IvzaZY9F8fLlKXYxM3rGVBeZjftHlCLK7k2YHi
mdnAYOfgoz/H2TCgYxY+xfdQ4kR6THftZOGVDshZEtO4ia6y8d9ZsyhMqDjG0VCp
RIQi/DDuvzJ/HGfQrGUDEyRFJZhtdkrGKUzSOVgfxev2pDQZNPGqY4BMeAlOO4Ko
RBi3v1Hl58Jtj6bZhTDd+gUZ3sybm+xBGIfWdRYMYEzTTRAuSaTmEIUsZ5Hne63X
SJncZAs9hBdobtsq5NK/o80ZWFQ6abbtdv7+hzpxEKPyU0RVXFrrwV0eSM3TvTDf
zkKlVXaa6e9y5056ng9HuAwkK1o5fH6dB30l9HJd596r6hh1nsyyu2ZbQL8mQDE5
cI8/5KucCD2dShOKprZCaZCZ4V95diAcY2LMd5BEeqIU8Kjwbtndp3Zo9D9RO+kc
EKpy3M9OOOpOAo1wXlROyLduOy9PcXPOa8RcfFsmyATz19viP/O6seesh0BWPccb
ch8f58ocVK6Pi5kZ4ibY52EfKvztvCuWVcW293UHh8ueXeTgkrD8PjWN3BXxj4Il
hrXQ06gox+9+qRVOK2+xMPOFAds5lngqbyjqvLjzpl+zwuUj0BI1+t1YfCqkygf2
02saizNJI6Jg0AaE0PPHyrQGRnrt3uan7gTUa32aGdmWSgo3QeR4TAFgA7lg/Xfl
tP26bC/lNr9DnnHgbtCWcfs1xs+gDU9IOHNSfhs4ZTC0XtXtrY+MFG9F4tAtFA3i
Ye/2SKS2WJbv9RQDAUu/o86bjVuOOUz3eKiACNjDATV8+joMcm05JENX6HqRgfmY
Jv01yoGnPry10WWdAWbGHeESKsmrox8oqtDiIb0wD4hkv8MF4LAnzieahg0GX3wu
n4+MK1qAaN4IX4bpOjpsiOFeodPmnIFyF8GFkUJqY2MFVF1SgXnPloI+PD54Wrds
WigeIbVEHQo90WOgIgfSGX7bPpyCtFRoJR0BtX6Xq13W7lOAEuai3kVlOZvP/+wc
O56eWTE4BaJMcMh7sZM9K/nUgtcl5mV8SSJNF+oYiLVuNHHiT1jZa82ZYq4oHZpE
nGUsNieyisg4lDC0B2Mcziq6wtZWq4YTH09Ds95nUdSBGulqAfekC5Ra7SbZJtf+
dP+WqpWCvkm79ZTFdk4blN4omSFxEYjDHfWoMi77I3JDM9crPa6FlONdMdi/h3my
kYz470xTVD3gbB8RAL1tK1JurNNIBXCfuo1Sep43QNr1xNHnavvrV58OZJjDdGZt
i6BYe+lbdhx44ReRp9uQFrt1xdZOeXPydHAl/YfLjeOBirvbf+pMtZc85XSfMtun
P7oT4kNEay5MO5wgch2DO6f2EHdjTDM8kuRsbgBuAvxDJ9PjwRQPPbLJOinyrYj/
HNHrtT/5Cwpg0AtzZx8VcLfA6sF9GQBpberDtJbWR7RvU1pQjzWttElNDearXG/i
LolKWvEZ1cBPqt916VlgFJ6nXkyCvHtYGg1mJtgdj/mrLJXAmDY6LpaEe/vbYhmF
nQIwYnGryeavbfAZ8KrGxv15V+6ZOSasan85J+nZR4k97/MsObsI3ReP4uIlQ4qG
CfNRxode0IXd69b84s0mFg6F+DOez4ou5vKGZPrhLaJnyHW/ywqcxJ3z9TlmmHgU
cce/C4K9ie7PsoauVq2p8fQwugf6Z2xP2IXUcvLMZsmy8fscdQcUG1Ekh8GVEZqr
3OvcZpueSWezCUPJzsSmRZ7gCNIfU5J+WlqcniJjWG5R37BM/6CHMV4Bq69aLXM6
BFGYaWKvwx20G463AbmyyDukzuKrl7xMtoAfUZsTK8rF+4YZTkaFHHhiJlUVBCnX
TLkVb0xbNYVLYhw3JuC3FhrHVMWoXSkIw/TtAe/LapIQ3zneEwYA8R9xdSNZGPfg
xZh73AvgIgkyB8tFIQ4CpXjt0XFW4MVVqCW6myRhMOxDWpU92OMhFTTLtxN5mkeE
Y+o86ocyXTEsYXw0o5pPUpQaO8gD3KciCaR6WqK0N0F0a8Bw1GycWDfZuGghxKRk
6MsxY9oK0QX8k1R1WvS8ErhsQhnq8IutoYhO01CC3hcASWs60HgAy55kbfDkyll7
3m7VcKM3FNRUrR0Jk4EQIOi0eNYCNQAv9qVjpdN83JnFaxVq2C8tC3q2ltvqHNFC
7PBXPryuUJbJIig+QWmdc5Twscc0NMsVRkEnpLe6WW3HVsN/cW1lgPzBvNq5WULk
BP8Jhn/K/Q+VU8flb6Eqdg2jCDoJfxXbcZxsgt1L2hjFlRIL5cPnYxAyaSCDZUhp
HwojyaCxDhNy8DH61dgey58dq5GKPs39cwP2YxX2/R7pTebEDBHLNRVmQkpm8rBT
nXvYWYE2MFMW9ycsS0Q39a6bEtwL3dL/+8Q2DhvgjcJzZTqTdISXnLgzH9F7hkbh
wSagWisvLTJUc1TdhWNshHlTMdynyrvZ8S18lJeeKDFIQE4b4OAe94CHjKdfvZZR
rEm/zAVe5Yo5yZowgk86Fgmczyy38Aw2+whGbbWTcTufgMYvIpd2b8Q4HJ4jeplb
iV7q+Apycn2ht+/pRKKu8hxVWBOdb2fj3hHKKohyEF+ssqHNf/hphqaNuUC75xE7
0d/FPDZKe7bCE2V7Yfnf/DdmDF7YkB0oytlKKTosAG0ZBKOM64D9Ac2qnj2aKHjl
2pcTSqTJEnllbbTQacnCuOs+WRNJGztnyVSSyOHr7tQJRc9t0rG/WdVQ4ho/RyI1
Oag8BvPonWK6SUenqQrT+UzOjmRiaPO/kvul38ml2+1pdq7cCzxA/+4pClJcWGmg
wCcgbZ0AWcYVWUnJfsUqDy4cQ9YEWTGUD16DwxMaj6LA9ApBhXZKR1VBlnXRpx/A
quJVUGOS7aluwfnuA2bdfVFd7xtCHnnWsKf1JwVgJzW6GRqlBJXtHdeNLABokXPd
Lnn54M/2aGP8xdSEwtFQJcPkgSqRw2cyUHNszdSp2zCFM2VZojqiaQWyvGn7JKOA
MFEKosfd/8CYBl6vLyOWBNRf78O34aeJo+5zJM8Kvf8p4zWmwRFdYYR8duqEWpHi
lXsxyWWvhDJ9cL78fc6/6t/clU8obiMm42D+XrP/XIHF4taMCjItbPxUFEdOpHEu
1E/lXZeWgBeGcg2nhR0IeAuXkipGb3P9uH6E+S7ZhVZbuG1QRp8nR4A3/NOIGlZ6
aZvXdtH8VuRm9yJwynfXDOQuQL1e3BuNvyMNCHszR/nG8AvqM3zUk6G85rQoMYIA
eCJD0PU+ORozNfr5VtcxenH5Dk9Uo6M7LMM7Y3w0sXiuz7ck7ea2tga+IUxdGeLu
ohz1o/Dw8IxlsBaCT06tHabs24Lk34p1Fmt2VfThr1W53Tyh93pdU2gBoh3x9w5a
3+P+H/2GTmfyoP+LeLMuemkhYVR6Tec4UUfbLqGjSd2gOGxP4ZcsmgQ+sOuIOJ2a
7c1yTDPqHIITqNYUG8TlTFzlJtVO2lzlc56YbZcUoyqQOftPYFvUkpTmV5ryuzAf
xLRCvHVSsWvFhAA/8eaZ0yG2xUAJmzKZI8z/xFmmizEmJpxYi//GD5SRkWpJ66Ag
2rosw3Orr6i52qPsDeUrCdbtsjmKB/SDyM0KwWH1R9V1JQ8AkgaSGcfcGrKrMK0V
P8FIlZ8T8FUi9uPP6d9bIyOLh98Ep2qsSf235dmRW2i3dsW9Sk9ahe6PsDerOxhu
+JFy8T3knqpHPL+9Epm5j2vG34xHe7pR5XOBLCPWtT06mYgJRXnrzxMH4KfDC+Os
GWcW/YOou30GzDKyuM+0NBkqdScdAebW13pTeZgNaEBMRRlkyPPhFX8lNIyauwDI
ofdp8G3msUmRwHfqjJ2ln4YOewU78S+cDhztYLIkKhk0kFAL/RdmXsOWzG+2SXqW
bwqmjeY4H1/Mwpzni5oxyGkRMYhOTiWI5aiVu+BQCvWku2LU5xy3ho7U1UVSCXwZ
6RKEJ1E0076ZB44H94hgk630bfDLSpkjazDESE8dWX7Wtt1uZ3Lc1dzdSXBFO+Ia
bhJZZEvuwDekI1PjQiakqACsah8F3daLusxp/R+2Zm2Osb4wYStKlF1rxZollyMB
o7fnDIkvI8oQQ85/r+l8rS4aPNOFIWt1AoPkl700zO9juvj0yT/9bSAnCIk8TW1C
qEGFrWprGuMoZcVdesaqMg0BmK3ckVdoqjkSYWvPZk+hPcdySmmRrm2kYaJxN/mx
X60llgL591H0/bzsH4wo0nMsbYJjaswTpGjtPMkACkP12O44G18F90TBMyN9nBhq
LRBGkmLG3N/3XMj6XwpoHYwDqxEHJZk30O6gHOuI6ajXO36LdeNDD6TauSlajrXQ
eiJXtKumUkJC4/ZQxB2ADgP/qqdWXy3+Th70mm/hDFS6zHXdRrjPcDAZyEjOQ6nT
R9LgJ0OMuk0zWCaDVBpnkowqlYDZIgrR9QprzUiwU2eC+Gxzo3I17ISXZYmskNf3
Vcc9ucpHQdnn1Tvhpxn7vaNSzpgBWeuQ9wbuRbl2qMzcsW3T8/uJPXAE8r6c0EYF
oS6MWLsEs+g/B0ED+5UkKB6mSRI5VLkSkJZ1Byuv6SF6QnV6RVhd1tdf4d9MVJ37
24w8AXhGZwwPsxJJaNyeE6OvfherTeEBnw5mBU35HDugADRZ/Ute4ELF7S7c1mGk
DgpIpzZRX6vJqQC9tw8wEw0letJ/6M0/k2Jo1Ef1aN42YgjI5jiGxjXqwpqWYAo/
/xgcLgeohxPhAh1mrNd7MiyaROB/1bQlDQV9QO6fCbiuZ2tCs+/Rk+LCgP/ezTyI
Hey7pM8Xxzk7KAPxMlz5PKFAqbPcdLn11XGNrVqQqLr9LP805WYTdVdxwP39mBId
F+SWFH3UJm27Nsm5BBg3XgJTjIud1bdY+iVEz9LSnNYUrsxgpSLsWgBhD42cF+fg
Hn6IL8zhbM7EEeYWJvgyb587yDjjhoY8Q3VYRSrKkz1xosyMOX3i8IoFQEpsjpgp
3t0GryqUzYJal5HsXx2z4h+7nQagtjbiFupXRsqkFibkN5RuBUagDH0CFQwH9VZQ
EoRRzrxyf5sgnntKaAr/mXFBGFL0yf6MrgGIF79oLEWpVK1/8+9nUdwrOwJSQsDa
24xv7OiAx5P6gy09J22z1X+t1dSx2OPtUoEoH4JF0i/JJCuI6YjxPOroBiguFMps
5SR8BNUYRiPcFckW3XjWIwronuuZyfpmQ0QaNa12WFbNwNk+ptL+/vJ5qQa4SqFK
7vJiytNt73HDoHVF/uQGcz2bfDj5vqHkXtjjceUCRBjx1xFog6R3gSmut/T0aMTW
iID+s51tl7b+ZTRxNGKVHKs9j3f1Jl9d5bSexMnOosjN7czjq0WGbiSFZNCsbrAS
hapr0DKLqrCcnA4mP0jP3hty0YRiCoa8V/cb1O+RIcPue12q4L9wxwFJCY6B1rAZ
z33cBMiaCKuKHczDKRMWDvdyv8Ju5i3FOsZWqzajS6arU6nt8+14pQH0/PD8HKG+
pVcx76rYBigUUAUz7SZD4u7evWjkH0aHlwQYvjC5f8XAvnOMG38Eb8aVg77Ht+x+
TYLFTCx7XXw/c0ErJNbHSP8CJ6WFqxXpYrTPpqLKrHeEW/mlIlhnZAarAT/2GrDS
7lT6vIOaf3Dg850Zh2/g/8aCHu9gPw3vUFOpN63um+uObphGBHlduu3zegZnQGp8
Lt4YyK5Zi0G1Y+LW5bHlTJ9JA5KpjJ3Vw6V2DPd98wjeFD/KVtnt/DSitMo2e8FB
e/188Hh4v/APLjjagNSmYcECATS3kAWbGGqwGNdgZpRS5Wgt9iNx2i8mY4EsInim
oLvnyynthxUlgrb9cLxyVYHmQn5EVoBTspAjUO9A1LLTGtuElBfptXYZq1xtcdNo
8g5TVIJCLEOAa2HI5c6aXe5fpp5b2bUV/d+McPgZo/nkCFRto6Lhge/lgfG0OT+c
nHXeNl+7wzJd80tQzd8Mt2EqKfp6nsiWbNhHr2YJyaBd9A3nAPXC0s/w8HWWZS3L
cNX9L2KqBNGBwVtMnVvt/+kDTe40by/8esaCiAho7njRdaUK/K/W/EX70wLmWjc6
dULhYqNfl5Tmko5V50Tz5pWG6vkwqzfJF5xrpNB9ZrTZjhioL5TH12EVp1iMZok0
rROysVYcnqrEeOvYEk3NfUThgZ5nxMe4hunJ9dJTiNnl2v53NU1KU8T91mBqY+PY
KZBtdiXfmSaT2DeclpBKkcuONmMdwiJ+R1UwuXqn0mWVdsJEUGdRn2D+hczqakys
paNrp/o8ukqP8XK2VScpgpAjRczTKGCg5m2b4EIRbWu+D1zAWP4PNY8pI2LMa/q9
wYXvhnIiuiW5bYKk/RXMqNCO67ck6nEvy8NQNtdNinzxP336iZG/3E+3+BBrvMET
1LPeVnCmMFYzKKT5+bFZ8orbg+6eGmdOj8zGrWLOkUTQ0/Xf/Wkl+TL2ARrJz/PF
gXI8uJb1njqrQer/Jyh7cx/ODoCLZ2QzgTtJqdPywi4d7nzQbrYbpOCEbSejMDTZ
rQZ8SVE7G61bkYSV54anCqYi+BzdFyYQij6cFDUO9MtbtPzfZDkehZfE81Rcf7qv
HkfFcumoYxLWxI+wUdgiJ2DkaMW85xTmf92L9IUSq/BvsrxmMA55tiKx5kHZiAwM
JNptysggbchrPRgPQCBLRQBjKg0Yt2kZ8O09NGsoa6lfuXx+0RIej3vT27LVltYA
yRGx+YIao8WbPv8ThyvWkWfhF57urLkmXUeitagoqaRnwndtSUC1QPJV3BsqJ+rn
cUXZGQS1z4ab5wqohLM0JrOdOc3nLvd+19wEuMa9yn/gT/vW4103tgVb6qrE31Eq
dqhCU2tcq4CQ1DnSoWPcchJs2DXIZw0+SNW/u/VbXLIgD16QSXmMtYDNdCLA/u3v
zH5GvqpnuR/szxAOCpfG9BoSuQiphBoR1iRlrJ3lVKmD7itSfbXbwyFuewv0YKEh
z0T0eZHuHYwiwEh5oQ2GoGXsTlbC9nU/ciLp7CgCdInsq45NKnGAem8mAoKFKNql
ao+kkoxMVW0aYJ7dnWLy2Yzce5uVxIDJnxnlzd+ClYnZv/CVGg0+9v36orjKEaJR
f5w8Ed6xsRYWu4FYOXYQfOb9S7dMk7aJTByEfu/m9rmVNCe8mPRnhHAbUgK+JWMO
y/KRWKrzMtoK1Az5PbnCtydLwDimiZtcLZIuBZm5eXNg6M7Y6I8t63f0aMi0Yd+n
GpBo8FT6+e2Y2LNpmUPzIu74KFg0y+SScdTbdu1HkuXGTuTeGGBwJ688d+NIYWrX
Ren19Pr9hhSg21m8rJKPlUTd4HaTDNPss+9r6eT4atkGEYKupnbWNfBNu6JmZWQc
uIBP/LNSuI+yAwKOv2xUslV8h4wPFGgR1Ds/S4IyekI4+bPKkfq4hVQbPHG5Gwi/
wf1K7KfHkI72Bl2Xffn/8GJ8q5uEEncOUWFjm4Q+g1MkjJO/Un2c1PflnWPqLh2t
a3G2NC2bLwxPhTLm4f4WsTfvJHeSrWS8xJMe8A5XAAa2TAOU3bhe9C3QMHQGhsc9
0BxjQbIwnHphxsaG+NohB8oqYad24A7juWjsXft04FsJedJEiS+HEAye43iP+ap1
bQGt63WmQWzv4QO/ej3lPQoiQasW4CnvjH8AgRCVvYRViIcxLiw8xoG62fnxY1Bj
jnGODgQXtPG/dvUlAQaR8JA5dgLpgkp+7bOGtCYxwz3ymDN/oCDo2NCode5tMAnC
7gc4FXGPxYWlWBru/qUhLnJPiJ1ZHFXnGgo89dMuILJYNc2ZM7g60oSAiS/VBYy8
NutDmWEcbWxBTYWKqNpn6xjwB18rnujT4d60/YTtejjbNE0fpEFLF8izMe+uogQ1
ScDQjYVONeBfPl32KqYwgP/Jl2rgtbkruvk1iBuWjJYDQ8DclOInRByiPkTacFA4
7XbQoMXG18GydXwHViBUieb8JwUK2gBHm2P3X5nEEsbeWH/rELANRbKSnMzRBERS
Kx5yL7gkbjDV+3An7CJcqa4QDO5fzSU4g2pqJtTUlr/AO+xuWQPjSNAqoKnI0WvG
gruHKLViNCrXUL0zqHNIyy9Aqclqf0RBVUwit1L5yqczuv4EneQOmpYQX9k7BdC6
QmlWqmf8zPSgdvYhkWL7w4Wk0PL2msuTa6kdTSikIhzBh9QvHThSkxLUvkSR6JQa
YOqMAxaSlbyzKgdKz5siaIZ0jVRjb0VH44gqMCqDBD+FFacg8hfz4S4wFWZlghOz
NNdX/PmYcDP6HT556+JHoSgeADdjhP9dPtqt3BGN9eqaSOOM9GisspXc1cYkBobN
blFa5XeE9LB7/JduPYtX4msN6bJ+ReTyT5P2/+3deLiyZgAwQYeal/S9fcwKlTQu
u1+DhjU7UMhZQtbqBc7yXjLr4EHpJ8zhNPAhnvlQoYqHAXcZKCOFzgoZs1RWoTW7
cu61hZRd7W6KAM0emqaNTqThuECUsBV19ooA3cQN8vAMldXGFJ91Yv2qkSHSCD+S
HvfpKzxmvxp4M8y2GK5BXOv2OD66UpkdrVjplotk75ljlgrLvrqMbFbtzcMJ6iFL
J2EEdyd1P4evTJ/FMlSk7ZLCVhJpczIOCoU33RwtM/Q7absR2kjIlQyMzXJzIOPs
nmr6jyqpyGfEC1lpV9WirOMf8ezLwZuKAa8I/N+rx2pzoJiFj+w+VEOIGTauJ/5k
jFkmRZr07Vm9xwHWDkAm+HE0BY5LXp1VxMy2dzzhanow9QJHmyC7ebKQ8oOcUanw
BpXvPuyOUrXuBin3zgoupC7lf5IcuxAnOuU98x9RmAhSeSVQnvqf53YAJ0fuNooq
QB+FcrOpXlA4b4oQ84454nXRqwenjzbGvejtoozLKndGevXBe4piEDvSD4+Vw4a+
jESGjelApwvccs+NM49l9hrbdUPiX9si4NeRdR009qWRMvDv10LDnt8sn6sA2P27
uc3fWn4bBDMgx5+2eXOfpp5CNebGGAzRt2xR89kd56unvfePhpFTF6ixnktuW1g8
MRcXhmmUXu+uI6/Cx5PKK2fT/PgcL/LU96VscMauLjchLGo5BQgGAfHP+2Op16cR
rbgs8X0oBh1bPA3G2wZV53nHxt6DaYD2k4r2nTBh1yudb5Bu510D1oIQYoJlIOe6
AhTSXW/sAsxJ8oXL8mHyXVTq0aENW++3d1jjAyzohnFKuRTFXuLbrO1mMpDWxSIS
ZApIi1F64zXY5PPzjvnb0YEoaeu1iH4AyILiP9lViAtN3TmGkx0yU4bJehVhyZ/e
mpWuNsYt4pxR+iis2iYKi9jPAgyNYSAXPzjzxkjb1c8rMDDv0l2kqvcuD+LS0Ak+
SOGuE3f/aBRZHtX7djHkBrvr3nvdplC3BJFs5VG23BwmhSGIe5UWK4nHv4Hfb09B
9mdQ6TwbMGjEoShbAZAfHw+GFFDHNRACqbV82CnUHw4/+wlcnO4Tk2fcR425nYTr
YNuicmgBDcCm4hH655250iry/nwoQQBO3yPg2hG1TyzpW7EH1lou9oDLHiw6u/RN
uBgyYFOTdav5mIiCr2GgNoLtH48BjyhJ9RQFTg/kfGKMxvAFNnp0veWk6MtAFTB6
zXkmCu9K5wjNha9HJ43KFJxAopvug0TP2/XY9bEimjB95VYZPwPCho0IaQAWjFYx
M1xnqUrSTWRd9BuLefjiRGp4ah2RMpaJbIr25FZuM9NlKrL859B4fBt1Xdxm2+8s
3ps1MU5yQ2Nk7aZazhLIi9cUgudRY2L6jVD3KjtRZqkrtrqLTVvyld/PTxRHfuLG
aUEiDrLxDaWsmjXlNHg/vN4KaaHSxpg6Km06+XCrNwvW+RX0pxnHFhmsD7Dphjqv
Vc9DsnBZ82RIs6J37o8EERDbYSXKido/wiJUnefK+tRJ+sdxN7Dfhc8PFgz6csOE
ft5q+WF5pro0CmeXVQTCox463c+SGyj1aPW1c+HaXFjjKIXMoIj3FeFN0lRnNiAl
A8tcLao6N6NxDd5ratkmBzNmbotUWlW8vYQl/+x+WiAMC0bYgNvo0JSuPlpwCeGz
qp7HyJdCzpnQjUXaYDDmuxrnq/yYE4Q1AV8FZwp8Q02YRdO588cesunpb1+iXWKq
xT5hO4Uy+4xGmAOEJ1R8VLXnIiz9KO1mxkIwqfAFtS0sfzidKt3u8+72E9jVpFmh
RyenMMr6sNs7VI4kvuqUIVbkDHz8ugr+07eczrmmN+HrXgoLN0HNPZe9vd4ozpGc
EXv8XELrbYrTrCYjuXzl3Ed1yARnLi/iJ5B/QhnhMcF/FQ2KDSvdaLshoQtCfGWC
Vdg7HxdIe6rG3wGr/zNoZwUgTQ0ByymceHf9rPVtD2YPlKFq1I7048tiVa679e2h
MftK1wTTz6LlaqnSRAP8dHWGwCkOAEGW6C9wqo6HsTQ9rnXRQZb878lw/eLdYYUC
w08+FyDcRUoiXPo1QOZa8WDTQlkmLtZHf4BU8nLmQZ8JTKWvzJpvx4gSY3232UaC
FN1TOz5rBCH8yUTZEB65cQ0RDP9IVAOT31VJAyBv1SGr0YoJhPFR0O0BfvBnsg9A
MFNlkCFu9jTFaCAqNJ3OjB0OcmYcG+Fd4WBv4cPV1pCPj5aP7QySmUnHJb2BYekd
H9V6kvt9DuYMZfeFTbBbRzMo9EYe8xpnv9L9hc5HjJvRANkm7e7+8bQ9B24Wfdhl
q11vlDphCOG8ldokXXL9P6R70nnoNjn8dFf3t+uqjfBEfXoh4SAeDbc+wJh7pWV1
hIuXl3a81M2zc+FNwT+E0XZT+ywqpkLjsAN7g28XlLOPZfLDcPuF0ysKS6XnaR+8
W2REkHaac/L23bb/964ybB55EX7sQ8AhanRrgkUJsxAQLf93Bx92gyz2JDuzYJOY
P9bucIKohMU3CM1cQULaZ6b6NNn6mDET/7qFTTnWOruRDzsLsDGBr1ak/t/jba1S
acrdMxoP6e1kMeU4zXCvt5yMyrO6qSqT+jfKfMxg2oTmcT7Dne4H8cZZT4auBZyr
ZDG3KBULSQm1+H2iAGPu/tGxMi2ye4mNggSdoReZk2nV/fUq06udKb1O8REvwjz2
HGUp05IJQnmTavjsamV+cxeoJBrmg6A4NBJDwvMs+XH47zIf6BQvFvXoYtxCTsVq
q34SrZt9kXvNX2OGNrEKBd2G7z+78i3des5aKh5uxNgSRiRNw9HMNJzfTvAlzZO8
/sSJCw8cKUpsr+snOlR67/gz5rlYJxpHS1Dcj0c8bHz3pNV4YJMT0CLFGXPeNreW
oQ3MxzTIuy1mtc0dnAnY1JUcVBmLEBOpdvXJkhaxSABepz+y3SLSpQK6ZH0DrM99
rprZPBcB3y79oCArV4QgouZzeapss1oS2851ekzT1LLCFCK5o85FAzAMVKCZc4Uv
dL98BJSqu6TIK/+VevJP+wsAIwkpQtba9dDEmDuryoKZuoh1SlxvkoiF5qJWH5Ak
dTYT/Y/BQyThNjM/dbLLLr2S7noJ1E5W6Q8mTM7cDOrADkEeNULBPG48J0hWuRcA
FLwM85G1CgUSKrICB5UofhWJeSfeyojHeGDdp8KzBfpeDiNzMwlondI1zE4SnhwI
jyyRNZr30Njd+ay3wfav4v0gFNEHx9ygjdLJhcY+RogX1TGMhecZKQbdpCJi5+ka
fSKddQbwxhbW3YUfLcqb+x8DDnw75bHIwjbPETHLyeidkKkCU/eHwMlVkKD5O9Fj
l+F6cE+OKyM1r9+Q0w978O+TDuzBKUfzy3EmkxAn5Ds5GBHeQ+BpBkrwVOUNo1nv
ly6V1opGPyVrRx700rOgSIVKznFDvhkGRCnAdrooSi83J5eexVl40a90U4ZNvPSa
ZFWGL6YcvvBSedOVqHCDsTr+wGDuv2vj18S1blzZ8STFc1tGxfHDlyJ9oCcCyGNs
xEeU0/26j0byAkJIQIrp0NhtGG2e1X2MXUIAKzoUZotqOsv1iaOGLx77L2fhI2xe
TSTrcXfaDJc+aYMTTidWgXBI+81lOnfz1kfUWDmsGXltxHC7Phg/rroUNEEnvys9
JE5m6yi1j0No/MEvYG/IZl9/R+Gv1G7gPLdzmxxmsqjdALflVQdEjlwAGE7wR4fH
SHsPXs1OTADrdbxGDtN8JlhwZQTZeUlWX2FFJKZYN3Iphmdcj2anVc00hbRGVj0x
qbWX1OudeOyvSvDHXhsn64fwRbfbGwBR5v4S4lM1wy5LeItCnPZSmOj/CvuSdCc0
vpDU2bXdnog71vd+L15j4vEDNus261GzmRv+ijkklrDbbaz4XsnofxjLScm6zyoc
6sr0L/EYUyFcS+0oa48ZLJBXxPy2q147tj/LLLSbpVlPEcWxtFyPIfJfHdSarMe2
lBoAU/h8CQ6LZv5c62sWXjOaOVfS5Qj/W9DEJz+pyxqIkX0XbWe57I5EkYfYDzRZ
xg8XCd0bS5qtA1LlMPnHSfSP14T6Q7wfUvL5lYIh0h1VT1SmoStEdrM0aQQQWumb
DSb/7A7MTTVb7ZTOnnpEVuBkDm4y4FKrajQAkTXC2lrUJO+dYSSWDk6fd4w+ox/r
ctuHSyZKTDtFSImPp5Wuu3168iKNj26BV+MxzUMez0XCTeRERxd+2lXrBeeqO7Pq
4S8LVzj1rMUchzubr13HzTMSHUP4/NcDdmRUCMhS4qdNTvFX93NgcVo8N0PtnhB2
gIuP7CM5z8q3HVAZM30qZ8PS7klaqjf8d7jMbb0G8EyT2EAcrU8XzQS8bHPjohnn
EydXbuBH7Hyo/iBurz+YentY32bzCbSHwuHgcEmOgLKKxrkBmp80F+dZxcuQNc2Z
LMWuC4FO/m2RmeqY0QL1/09/+NZMuB2k7TUIUzS7XAlU0bZGcPZQb5QyaKbOHbcH
kN07Ee9rXVT73kuMkUmhaQd+Q3750Zk1/n/gQUZ31qQzpSDVe9tJTHM3B5L/aa3/
H3ufFvhXp5CCNNxmb8B7Oa4tzsPaGwTxGafMOzobzuzuYqyUFe5ZPfVVBscx6CWb
METnF+tKGjidLQwkNzgAu49wPdgoyKb5XAsc6a4EqUPyuDlAQJsVKJ/gHNtY6gLb
bXAgLHOKjjXu8hmeG3FIW/fq+X0PM5ClyVa82wgSaGqBxJgkUUuJCt8oa+9Cvk3M
ngpnQuhyTQKpukDvzLyNrv0uxmb9W2VlR8gI/As5dV79+6GUdo0cqHAumbLwqvG+
er5AS0AGh1JbB2GXH3jXv+5PUwH7Ulio8LFyj8kRPPDLwizcsR8ga2FCnp+YKK95
NYfrqgFcmK7SGxi4FDa0HH4Dx3t2WgaS1APR23mjd6DMiMF+JmXVjsIeI9rnN8sZ
W20PoFOay639/DRgH2W2IzcpxkTfxnKDzDCpSH2v0BZ3pEBETjipYFJvI33waocR
16ZIaeZA47dRdIZvjKxIVt/+V/uI1N/EjAjRcPx0KNWYYEGwQa3k0/eLH0YAjve0
htHBRP2ONB+6v5Bc/CVM6XRNUMOlwl1Hfol2Ol0IxQRyOLEMna4X9MfQ//8kutov
74OoqO7XAT+3RKWQ3Zy9oTkaeQNAKkhhzAK9nW+Ed20yfGM2aTxbSHlZSwOCHDy/
gNQOT6HGc3WDJWm6OzLQou7xDduvbbofroTWqR/ypNQ0+PO+L2Gfxk6RRrekz5RD
fMz7VpFK5Bu5crzqZ1Rxqm7nkAuipeec8+2aWTJULdXtfJ2/yOvMbXJHnwx4Q+Uf
BCItLVzfrVak7T1Rns6uQr37UWdYHNFwZXuEQEoWzbBwIpBt9m1CRO/YufOfoiyy
wNidWZNBwG3VMn31n/L4r6WC0NVELf6pZrNm1mCcAKgnn8CgU6aufwh6H7GzRN3k
WPAlqijil9/JLd1IJOlKt2Wl+24w2sCMR7BGri6MzJtOVJ8NZ439r+moJ3AUuEnJ
Xe2s38HuaaZgYQ/URNECZlJUnRTDMPKNNKt/asxb7AqLvd/JXYgUZQXdL2Vk1rap
8rXeVVkKqhz61e4Po5VEljXnQdDbWEfNwWYLHG48lr/rH4egP5hsZd5DpG6VKT3l
vN92q5NupjQqKzs+MXHsteit2OGTbwY1MNzbPZ6wdhMd4l0GMiWExamoLzUck6ji
bSRNl/89Y2wEXCT1BpUxs17FNGzIK+YAu4CpQFEfFHV/mfx4MdWjKmL0xu+BC24z
15zchpKOqifx5YOrovtQx6Vh6c6akKZqj6hYPv+DeS5TdMZjV6Qc2lvjRuoLUXfo
HNGUr/59g32JziAzaBcG5jf8vSFh9x8c4ro6m6d4UC6q4FDivGp9BJ+3MkaOrnoT
2j3RX/4J0UK+hnRO9jrk+QSOHKvUj9GIEdNTIx17iFDgE3nocVZ9tJeGqhRcWXdK
MYh3CGFnHZmPLQ0QKvUhj4cKmeUUzC1DU8wXqQ2Ua34nslvMhloqhjjq2FXHOVbf
mQgpR1CicmTgASJBxzmYlWrzoz0QX7eEK5fibcOcT4G84sbaVP+/WrLiIPlWg1Vu
HfcBUBd4Y/VSx2kgD7I26Ns5h16zY7Kth3UzOOsYMT4Hs8rochDBMdkrwiqH2OW3
mwcQKCchQ6pMfWpdLv7a1Plwg4mnyp1CoueHszL83TdZflM0zGIfkf6xUUUsrtCd
EriVZJSawCi8zSeIAC4scjR620RU8JAtJEcYokLXap+TfQt2+KIvMkn+LMdfGDbp
x0uBaWQczrqHcGuSf2Xor7W0qWqz8/awmgKF1xA5R8Ss6raaL35QdCHHMtbWMiHg
JgA/npNdksYRzr5ZvJgmcFI7zPPTiMb1JuYlLJIQyRrYTdRguzjfXMGsLKI2u6kW
AmSgsZtESstRinNpXWhfhfgXUepIIeFdiEs3K4GV7Cb/0pZ7RAOlykpFaQrZYVM5
de+zgdumFlw38n2t00mlLc9Rp2LPM6gdFOPrJzeZw1DMvYELLPeGhwrkafQvNEpS
3M6tuDSMYZfr6Ir755sMOadDs9vES7Ank2aaKMykeLftZsTr2OQaH2Wfn5m2+/8y
EB5mEQDGWucLwzsrh3WPNSxeStUMkwFUHF5iD3iJ7RB4J6suXnN4MeQ2OZgh3zdw
A9Hzk+3ZRa3pFBaossbRZ7kIpWpv35QlqgRL30NDRNSEaGeoPRk0GqGJvSXSHLlO
CQBIV7B/NjvOcZ7sWlzeSVlAl/V9H+yb4V6Jx+iFjm4rtq0izSiEcwvphWWWwgxj
jW7iD1ilsof1UY4zjmysdNQ4m8yKHbF6Ms52pmJzCHinZ67gaNnbVJ68vkQG/Ujk
FXu/h6OsNizxQ5696ucYOQSUlHPmHbs6bx4a6ZscimUn486cWZoRDcrREy7n9ygD
R8ZDCtT458u9x1LqH9PBo9Dd4HM6TNMLCsoz/DhGaTnMy1x1e4AQqf8aBVcUGRjz
3fYpbTPEDQRftmtYmIDDQsSrIMkIz28jDKzG8mbcV+zTJbrILKimIneo3ee7F4bp
ECU5tMiCPh+X7WPhb6Hya2Z8cpJZczDqepud1t7VktQtYYUnux6KgtMSTd63urxm
nwTsl1EfWQc1SXazJaluy9omN5rZEJvm2OxgUoKDr3g8GperE84NPTayRsKWz9J7
BYw3Q+kJ7+DXAEdf64jbIdSouKW1dYRB5zTcvF6Rt4J+c5h3JRSuzAlOpRzT/hwW
HIYd6f4RpH7KnBnb4kXDu/AwlcqZkdyLJP77BQVC19GlGSvF/IHAUXFaMdrsje+W
BLJ89176BntrQunxBLS2Rv17OdYh5GIdg4N8621uFHmNBIMImrik/PThhXEC6Re+
GIOwvJME/HdSIbZ53n0ohPUWeSdUNza8gNsqFjnzRMdbKgPIxm++isLhf5ODXWH3
+b8d2zk/E+83sIqW/hdUJn45SqfRxCizF83rby8KpeeWHs9Ic7fQxqgn2kCqeUZb
r6C1P60SxdwnpnqirjeBUp+ckvAObl+IPPSq6sltni+rtYdhjVdy2OXwgFUhPIpU
wSAP66FiDjcZqJCiy3dRHziz42ZpIAsgThVm72swmtvv5uKjPSnr6jb81iNaIS6W
v1Z2KK1Ml19odhUqr458gKG7QhWl1/0OPIT7MLIoFfPpYKAF06IUq5chXYznZvtY
bf1I3/m7Kf/wQbWnhwOsW7ubFs0VymVHv3cdrUZ8YgnCt4Q0u+V4VY1H4I0TKqne
ZKO0YQbwZUfelaTHYjoB5LcwYNXPlBcs7Lw3AO1RqRK012ZqAGbiGsWT+hZcI90l
llbcoRs1zVB4vr8urV1kEqjZYiu/nvbYJSkVZX6LIRzYKI4KeVcrPrToj5OD5Rlc
72ihyaf8JemXPnB10KOu92VaXix0JrC+fAxYuib4GLTJGZLmXiNJ7zB8Wh5ITFsS
fUqdTqdJs1bTR4Ejk/glvrjBnsdnRUjHrnssiz4LIGK5erC0KjGXRMktrX17pFJd
/7kLjD01VYt3kuITja0NtFtT9v2e9494iYI6vA/iYPQCJoiG+3cnc/YZulFSkmil
dyOb5+U5qN5VHG/K8dyfq6Joz7fbP1qsbtZLIe4JbXOaPyGzga+rzbXuT542K/XE
Y84aPfblbvQJtz6C1GcDoweZA6/2mKf8+YMvLZqiltC1H3RGLefjAIJTh9th6zzr
LpB8unBOrXhE+5Cn023XBPd6SqBu2ymkGZwAmAxuvuOvd7tDpmGHk4n5UlZiYpjb
tFmDAKrQVfg9NAOm/tdSO4VRa1px7dlRpuz5Z2THbLuMmuzAeIQIk/PK2fgUJ3mz
Ql0roIIZ+3yavFW7sQpRqdojlkYagOR0fS5PKBHf36Vzo4Lk1lchGCWYAzfzIa9d
3b4Ub2YU6WUJqvGdjiZJtrM8CCmxA/6PB9ugR3eL84X2R+1BeLkK+bA+DUfq4rLB
rQwgSUULXo8jZKvhZevq2VzwIe+6YUZWm/vs2B3mmbePqeEEUaypDPffWA7O7eUe
r2T2thhMWAm87Qv9IC2rjhI8Xf5G5ma8E35PkmdiN6q3Ctf1zji5g5v5sQZD2Ldt
H8ORj7L08SWcddypYpQeybIZj1Kmglov41OoieNAAJLDNo75ZV3TP9gZbYEJQq9B
mhqCK0Toye8QmVtAlcH2/LwrpiY+WSlaC8kjAiAplGQSJ4az8Bx69oG3U65XLYjN
Yj/6/K2VEIws1Q27aLlJes/Ke1SkJ4byTydBNJ80GC1HfSbMnkYSlBQszPQatG3J
hZNjXNBg+8WFqyR+RjMMdGKp7843HR+ZK5b2uzgxItiUoUmDgDzTenXJ3WhXoz2R
TFa1xTfFk64xnTbDxxy3F2MCMW08qdjsRL6dOc0zqk1P7CGqt6BNdVNiqq08yRRN
DGw/PTbhvRDpKcR6i5tYCkqO+KJWsz4YvRLq/aGeUrwUGQ2UzEe70dR4PeJl/nhd
wbXOvgt3l+Y0brvL/v3v1+fBB9kWJDoCucqQJTPAKutqnNYgmj3BhuRyX8H83iWd
OkPmPW/zyk+sFHhTFZk+n/q90Ei/QfZ2kIH0/Ht9zECI0BQ4ezxRoFIdpys8xgax
oKZGNlP6Sqpsq3rD1inyI+EgG/B1CgpUF8aKS2TMmb8yInQfA2+cFKf7NVtsLYcz
B+CW3HzO9PfXg+rclMzl6UYs837Qma5BF/1UUPAFvQg+3U14NHFVXHAP0IGTngbv
EIEByqVvBARr7IUqCeZOZwaOJZSuqQE99M8bxyANVj4zmFQNeCYxPU7LWODYEEdq
oPv42iDDlaKJiJa1abV7nQ2fWWeF/ZcY84iZIoSS++VbVmZj2o84u1WUcXyObrBR
RfPct30wca6j/K5xdgT2m/TyT/94LieOmuUYjBtJnTdM0yBIQtYSSNjWhXLPiCL/
TCCdw1S1nI8AfE5Fch1VzVrTu0mc99X1JbG1ss/S0V/nM/j9RCO7Oi8Av9yG843r
AkraEfT77TAamc6Yq1DCaKvDpR1f5l/hs35rAxxbRcym/RPP43zfz7rX5NuaucIn
MAkCAggU7aLQoGs9AdWIHLZHuZXnnG/qt+r3+C83PjvRgB+5GRDFvIGI8v4boMYX
wtj0JM76pNUnC+UGf1xwVBCi/398gK56XeO19oczuErS3sX4zx7oIsTeJPS+d2xy
CfEAqcci7Tfbvft7Sx7TV+VxhI/japTJNN+quv/xAWdlMinqWRcVQOAPGDXVKtqX
Zk2gFCkvyxvMAgTznU8aDf6+/UcOIr1CSs+AyzCY8HdQ+AwZHYy+Q3Ru48XqPYd+
J9EH3zHCtI2FaZ0aClORKFnWjquJlFB3y8fPosejSCvKVaT2WPVS+3YNw0++WtT+
AdzXHS2LGRD8AR3E6rQ7kbZUeUEWhisGrf5iLr+7S+bIgVhqWDd0ksjYkt8ykaKC
c0px1U+GD3mfJI5qEqMoVkEiL2j1TT2/Y2GL2tiN5QWiaVi9j9SYjaPKdOIZF4e1
1qCbLGiigW6x5dh93FdAQgxyNOwshHShaGINmxOo65BfOf3VRswX3ioT/5nhxTly
k8+BB3961AEB7jokOqCWZfNWLOMnHjs82OIUqQ+4W0d3LYsIr4tQFmVknHujpF+X
i2rI1lHd/8MycYmIHzxqTEIXYfnPKzqHL5GqMkuBt3QQAd9CPNo4v0c2ackgOT9q
3IsZHjc/pOHvdxZlWe37ddHdx0hOl6FnnabWaVL7aiAIcCSI5Mv7EBeHHsRA9qrO
THrGzI4DWTSAOtimAy1G745jX2Z+VArsDm1oaOqA+iK3YFErrqRN4zZu/fEa12nm
Zdd0F7EVshnNrsw6Rrz/vcuOThYu1Uo43IGqxHvPj5rqoiLyTKPlWGgpWh3ta+dl
HEA2slX17qjzf14bWDUni6wgAvHIC+0U9aq5goyRAcg5l8yqAC9e034QE4qPso8W
d+GBrWGKGTcgonkj6OeRUcPnaPPJGpdXJl3Mc4AvZk7HXUyRIAEr2wcoxnU7q3IQ
0d6edTvWD/HgMt9Pw3bJaw8FkMQuGQinQdTXee5eH1D+xYe3MFatbGrZuPBYLNpw
MgqVTiJlHoUnjnfhiorfLL97lRNG3Duwq1AOtwgodYGy5zg7AOVKBK6F0ycSyT7p
I/AeZQVVSBGjV8sQ5nN2emMF5yuu3tWNatU8xoOZA06p6D51heoY1FnUXYT8j1+b
hTQGK945je8x3HNhSSPfz+tH5jyArNlIixibjtR+IjnGa4RON0iwQCpMU675otGm
TP1qtJvKmDTD+oWxXNYfbNrERIaOuViPexjwp2re/3fZ1UU+cbdQvsPBnmRzq0SW
YiQKPKNThZMtxk0bWImG04pTFHv0E/tLhCdfxOflRjsRKGCrtKXOrwcI7QFSz5BY
cH1bj+V/4dnK6ZkQpgtYdrl/Uh/oQ0G9MNb/2xMiUEBUgaxuvpMPlGXLdcmqe5cL
f6IP6FrFsXzmcjlmIt/CFiMs7whszFx6zmrLqoNjQjP5ReL0cErd4MUUPmAIXiFw
B6ToCn6mnVcZ5q8hSGpW6yGDntqAFIpOn/Oxdyqifx31B3B+bkaxq71OjtDZqsuw
cyk7mn19kwdRGtUjA8DfJylAC7gwYhWfjf1W+t9eX3qSzWLoLzOS5hPdnw59OAkW
aXlzihADZeBqJTBa/u7wtC/xjMuZpiaulmsH+xD8OVzmDzCEu/fCbIz7XmuDHd4T
fUxP4kt28rr8ws/lsUESmhj96xVbK0kEiom6w6x4RERY7/r+D+pFqYEqKzZmxBBo
JCjopt3UDDiQM3XqtmEpzjkeNSsyzCh9spZknfMULtEWs1qHMFZMm4N/5BU1qfPz
SI99g8fW7h7d1glOOmlhGGCIZYnLUZaYrmR8ca2oppz21Nj02Rj+bCP0U1vqb5Gy
qIUD1id05y0Fs0e0ksXifcfIXbFUmt8g6DMkZulPZa55TknPC+vCK/tanJdMZUQl
OIEx7YMAb0xyLg3fScO5E1g5RoAqFtB++ynqUCEMEts1KpabTPd/FSv1r2xf3/HY
N1F/9+dUP9fcFnOaSbbV0UuQkblg43h0WRmJ7JDaYQv1+El98C/CuNpMk792pAB7
lLt1vAKJmvuxDWV/F1wy7qyvOBlXeeD/RJmcL8CWsWJ8zPRhDj2LlXYmP+UxJ8hn
BrwIMs/+TDYjmJNwSSDPsD0IJd4BH67Qsqa6uo0eOZtAcZW8WzrVHKmpBS7Zvf6H
Qei3Hqj6d7juaLb0j0M4dGow249gCaRotjA2gmVS6BgI5nMvN0oadEV5g0pio8O/
pBUdZMvFLZJdGxDdkW5bH/I+Hg93BTh4ERWaacWQJWCBkHI0l/3veg5mwiVc9I09
Jjm8NEEBVrpBVl+lnwW9NClwcC1pxg/qSpKUX+6yx2rGUevodtTsBOGpmXqP4zUd
1FJ4G57yhgG28HrntJbQaFsdUlN3kyJ4w2Ryqa74ngXXWL7WPYXiWnKPvO8bW0/d
HwE1aJ7yoKJYEPCehEwQPqwAMptsuI0jZZ08wnmVYrNpqXl32xgysXRM1vM1x95W
Uyaop1J/mu6NBC8RUDmtxZ+n+3EfiDk1eDXZYNrfwoREYA/oHhVsMfexLiMwJ4C1
RGGk/GQSWMZQw0bQWFc/HyNOo/dyEQcXNys0BKdb7QbSlz0PX1GrcCRr+wcKuT1i
PL8iSmDweHC4h2VRKrLPorMyqDtBwvYEiBzv57lqqTRm8UcEboxNWrRheCvMCsIB
aAS9DPuEfO3yATPYyr0/PA6X/HLTHb6JUvkRKpkJujbBqYrrJsOe/f++G+SCLctV
lweX1a1gJnrISGjUg9BltbbsRFvncc1UTrFk8XleyiPr6AuVmvKS6AMTUlWc9lED
6bowr4Qb/5kYQVs4DK9rfkT4m9prK8Tng77ATjT0NyulQ68zSB7Z+nf8nVLu3QyJ
1rCc2hDTHzYk0JJkLq2PN/MGosIbn2+Ch8XItdReKo6YVyrWJv5Vl+ZaZFidefPU
F+A1onzexo4HoC51r0i2IUqmaEfQ34ZZhqYq+ro88kgUyZOy+yiBk+bDj82ODU9N
zH8ziqplZ8gnkPW781fR6n6DKjaiijfpFPEAcLnFtat8/N+zFgIrhiOYvSsJqQRc
VIVgVP2fRZ88SBoxHLnJZTtM4tZZ9DdGJZ39z4iVr75sNcYJoJgxO3Izwa8bXQIl
NIxCwUVBnHz4wD1nhplVA+MNNx7/v0b/qIzbDRiTOllkb5KFcL5Y/Z2w5/6TagVL
Zdc4cx0ra6IwZ7XRWxx8IMliJtOTB3hkpPDynbTtJwOs7NLdhDYNp245y4ZGXGrk
y17UyJNJ/IVS+lh6NbQ3tjI2XV/6TCjqwgDkM236fBSJgeMz5WYipM3XzxUaC2Lj
41RNrJp93lGf5b4Vo5/374T2edCfZm9xjfxdAK1INayU8O2vmnWtewBF5oXyzvJ6
/Kq1R3S6ADi/EnMWMlYj1kuNPXC4SGbjzp0B3opsa3ZbUiXgQVz/jZCinrbkW1hI
BbHaaTLPwraahLZm0b59htcKYhamknpw52p4p+5Jaa9Oj/k1jSEVOIu2WHrS7bub
m5CWVnNFrf+tBQTccUNNxyu8H6dr7NAmA6VONzXD9Hm1SqYT4M143Ji0Zn6OVtpf
hGPsgWeUXi+WEel8uepecAC3mfXCEDhkeUpKpqZISt0i3E8HygieySR9R7+nq03+
zQ/ueLZIOwescn7pgFYYOThMyIIgR4+MelDElLy2Xrw5D/mthqUADhJW/uJ0SLiq
snunqqevmYLOc5pVMxCue//AV23/RJUPVpahErEGgkoujmMgWhFBlhCmtHvcS0Bf
o4ReBO2ZecqBpe4QDuzAFLHc5wrvtKb2izQQL9LPUC4nc3MEXY51wtI06sRYjnek
VYGwn4bHtwVrLoBNyfr9LeNYluGXuzB0SZPNMGYbtJC5UpzWYJsOBV5uVc6oQGb8
a2q/M07pNER5zBoJlGuNmvR32kPSiOvVNto473ZOY4h4LzmNmwm70kMA76YUzSjv
hhpOAZpv0S487DBoBkdoMge8waroC+YjPrTQ4tRc5Yzhm70CojniV6HdeChOI2J8
ekiC1dt6FwqKiSMBwB/LyzPiVfHASIbES7oVcMh8GcE/sHmLMmTUCt/84LQtApFM
5CV5U3zd5CZW71G/xiFv/Qg3bWxaXozo36tGRXzPAl7FfQlwW9kdYeUxsqYABk9G
9AivNKi2jOaRQkvDRqHv4W8bFAzlCeqVaGYUXSWI9BPth5GHw2mou/2znotIHZfY
hEq0nA1Mji5wrVdTS3LZoia7S+woUzhLrbiAtF7xJ9O23Y3mcYhGmykf/kf8RVEZ
EuiwEaBomA2jwGJ1MezFH7TrXhUR1A5AIWiV2J/SWZLfxeZPHKqfq2wI8/z6+FWG
kkVpfUEugbFieuG0GbY5jALqfm9KcnryZFcNbLLewyB1wqYI+oFEVpGtM86Mj4qm
FOeMD1RVBofC6d1Kw3KVapON3iegMimTJ3VwQ4pKhATnpKyye/ME8u670xc+P5bb
/OfKWpw0kM5Bswe6cK9l8/eErBwtXi8pX8+GIxn/YPgqsGxpmPPG0ihkmKgWxVT4
3PEPcS+Gl1heX+IuC4OTbUYvY5D1K9g8ZFlffddsUQIquFNAqm/rsXfuYGrCPu/D
++kkbqfQY+BLaJhB+0jMvT/32OwWxNsjnRsveUBCU8Jhtwqvu0BJxZvFDv3IDlM+
aeKpbGasG7x7F0owuqFaYydip8gEjD1jCUOEmmcqDiOS1FIM54dgKieUnpvQpH6J
cjtPv/ezYyjR189iIwPsGIJFzSK6je2IStlM7PSxxhJZAtfQKvKo6BnJEJ+MkK4s
guC3DNWv7JpLOogSkIbLoQd9pNRbZWN6+x3CKbSJa3MSvFLcih3Oc72QMb/y0kOu
cXOxMKN8adsXPl6GPgx+5lMLuiI/1wZLExAiBt6+WgRYupvptFzitQzEQKJxN3c3
/aKChR/y3NjsNjFeGPwgg/s83ff5mJkXYsMumlXJc+7eE9gGjk04NPWjqGBYIKur
JXMET5o5zVtHWH8w1MhYTtiDOknQr+EVFRrYb+xmaHuME50VhFd+SSqs8TahRBvo
UbTiVHxV+MlIAJ3TC0ZmlM+20ivEfV4xqVDxK6DFi+zyNb8az/MmrmOJHNNdQaH3
m02cB4iJedvZ+y3oTV3TZrgrqcH8QXrGNCwF/KXcMUZmwAGaDJ4g1kwZ/8Kvn3El
vDuceVNe3OepIB5FGRraksDFHSw1/B4rF5SNaeQCzOz/B8YiyMfPcJ8ltZ2QUMB6
kmBLEi2J1pmKxqXSYVDPF5BQ9RghRhNP/Af1xXQNe9GBfu47w3p0bigrUZwrsIFq
rkmEd8r0v6QdkOk7AZTAi/2Es1z1S2Xj6OtD4Ar6MhbbSQU40N806+RwFjGTiAws
qsgklyl4qi2BIyCK4Tyz3svSulc0h2UFvxn9OU+DmrBzFPbanTha9e7xJTbgb6d+
HzBZ6L0Qd22OR4TD+LVKdoSFBNGAfbtjogkbvxU7HOd4eAFNplsoFBrXJfL/q6j3
HP2dowZEcQWZ0HFB7787nyz2liCz39L+tXuY1fkuCjj5mB1Mx2HdGWBdapmzfftd
C3mHT1YnfzDXxwQI3aLQKH4TNIYhvKrf1DlAmBkxo/pNzGm6hjEVxtbraoWq74n7
NiLG/LerqyCCxWMkJ5xl3hJti2wyDUIbdXuCAf3EJ2AnM5lawde6s/zPKcRP1FtP
plI1Tk9w1RaMsfNIeLlz3U2Tk42XIRlYJfZYxc5UNtxniB/2c7XICRbbamWY/Aun
xKIMgAJocMpJaI1Jo6VQAAziFOgjtcSqbhFU+UqGKaVEKMZ3U2OkxfSCi6YdkOH1
U0CGNLqI4/tWvOFCyucTJ5epeR2eo4WZA0cy6/0VM34Byl2jFmSyMOj/Gl0Yd4u0
In8ZPPDEc1o/9Yb2NQmmwxrXiX4Ht6brC56pPb2XnmYCi0W4sFo8MJgzurCHLgaq
u1z3Q+B4QCS+NwF42buTNcSvrNVz1DGXxdiBn8wOXF2B0WfOvL7QIVQdmdmoUwog
WLhx7nD98xKL5B+RCptKi/FAnhHJz6VmSr84l1tD50hS/aDnuTMlHYjCo9QHmFpF
ZB9x9NpL6/G/sfVN1p/wkT3r9n9iR4GDMFaDsl1lHXvqLWiyjQONgJ53kVvYQllo
sEyf0SWxFT4T1E19WqE5KkPnSHUCsM18cjk8vZkUNPdY20+wvNTiPxjvGqvh0Fgz
k3//u5h4Eh9tHNs4DgEo13QXo3dBaKJCbJ+geFVTyMBxMru1TUF/Rkt4EKmy0uXq
n4WfdDuBhfJUhrqGy1UCh1ikJjTSb7izNaYBB71bqwAEIgSKVWccnLL/8KdCiJFz
5uRwcLA7tLgO+JkfiPlg+P4J8P/hQpUqM9vp7kZnofq1uJxCZnbMQ0szv7+/NmkB
guYTaOSraBA41eYwGUFs2zxneEQnXA9SV9fghpHrjI9qUxWz9PMm7XxD0VfwdJKB
0mIiaOF+DPUFrthvhd/Fa4imKyOlTcg8ru9m+yrwmx2ELBxMLM5riNbW+rz8tskh
8Ou9RQYt0q1jODE2D6Xqvy373vG6ZMVQj+YMFCMMprugy67qwd5u9r0uK8ZFtu5t
igdf7Xc5yxjRzMRJ2uHy/bPlgLeER7pqOKFDHENqtB1i9/10irU3OoACwZJmqNiH
1QGETjhhIb6kozplCfPh7uNmcfeXyNbCxRvR3zsml90DEO3JCtvYi2yPKgm9gFVH
Cs59lewnhQsn/2R3MO3rcZbhxecYJXcBn/47OpplkHBEpUX27Vvo76ZUwXgFJa46
RNj66/ko/wgb5CIFb24vZVBvzCAXcLVJY2VeLDLPCZyHA4+tOhJYmsOy4FQmhqht
jcYW2fE7Pe5NxWLFe2e4j4eisgWvHdaHIL08UQ7cdy2phdS7qL/wJwMoVvWtWLze
Ts/tj9RGNeBQxl0FyN5mT56v/hoB7Dpeke1+sHDkk3iluZ29pmCyDrCWItgui+z1
Ss4G//vynhjZMgSXZbQOP5byijoSXRN8EQfsiwQRqAf+M8dnuWpZME5UglvYuEuZ
Q36NdgjtftrQn8xxzRbFHo4IV6zGHn8KrCwKfVD0zQiNUnEGYR8pzdn5e2aIDKmI
6Nq1hofruQZEnleYq8M3psjY0cHHCiZUjhup8KsBfGFyr0so6C2zPaGs3FDPQMxP
KM9HsTKE4Jc+aKwcD3zdouxpZUsAlUuX2Foua5nhz0nBBvzOP7C9/nZ8mAhiXuV9
Gra3pEz3Wr58+ALM3KUMPeA4r7KBNxerYXRy5xOiYU6vW6tOiVMbC0E36Nv1WqpU
EaVXuGtbSVoDZYGuJTS69nW2XKYoj4mW+wD2hs7CyserJCahqCmj+jAUjBwk3cyO
a4DergBn01EkDDFL41wpgZ6yZ3F9Qm+yLMvNoqJj05v/3Ngqdcy1yDMGYWv3Yy3N
c0WD7v8LdYsOtFk4subf7sx6n0GlpxnqYp2D1lalJDAce/lzLHzRDYJrQmIZ+S4W
bnCiH184Hih2Bb8CvTKQeL125PqYsrne8Fji9VXa/tIn2Sb14h4YXWd7j7F9IxaQ
fRUVAWEkLIfKTvPJbY+Gqy5RnLe4gtqqAc4TVgcwEr0R4s1pr3s8UNvqgtSxdUe3
MmVfydv3PuFhPHWKiKM06cRz9H5aBiarOQjSSUQ/Nfi5YcMRZoJGKzaurwnr8hRF
jZjYEX8YxiIlV20hKUyaw7FYxuwDyN3Wc2PlhG+kqoOzEzvUOAZwWbWEI81WEz84
5XHMfD2dtOY7o5jnWis/G/fhrTsiegGSZAqQEx7jap3LGYywANGYXw1kXw9f6so+
hSO2v/2FGOkVRbw3JrM3SM9HqKzZpy28WmpmX+KjyWE5xrKw6lsuCdYj9zDNzMEn
JTDSZTUjUGPKDKapcQ0AI6Ll33bG9fyRk83pmEJUyF1f0nbBvQGC+uMEbYeLPkgY
UCjV2PJ6bgkEdMjCgH/cRAgRmhGWBOmHUVRlQEYnhBU3IPHH8TdyUkC1h/LR5sSX
99Qkum1mEdWiaqyui+srzXmBvdvLleO4hzXnKBBJ+BjBWhuwzxTSc+lTQssMAl0y
FCmNG4LsZb6XmWZtDb4n5R614MWCxlrQM/PiCk0VoX+LL0xRiyf3iyU6d7e5TVrE
8dr0fabbXS+wRyzEWwows+uwF4Fbtm8dqSxXiHBaRhxhW7oBlEsSbbsKPsHwNbhH
fvt3ebUShjVthbOQJhB8b1OsgmmtZUcMzF+qcIVblkecn/fBtXt/Y1HV/N7OOYED
Gx1WsUKIPRJuDL/Sj6ieQLxyuAonuIh7bcjIC/1U0a0ntMdwrqcVMIYN/+AesVrh
tVyDgsT8KIStCk6O7dD7VRRnasH+mrMQxUJR82mXw6RRa0/R4r3eY6C5Ex6WpfQ8
TvfTSPTYzYGetGWFCYXMJc9/zNOtNFe/YMU3lNlJKM1xXVrj3ti0TcDsfr+tyygP
Yww7SK69qaxIO00cxc3Y7Cj/umMbdfcPWD3InyCfRM9Ey6vVqhVnPBUAoG8LsCwL
Xh98+fLcTY0sh6AoDOTVnzCIweZD2BJ6w8gGrLkyanezXa9FuQsFspJxL/QR9sk3
8zBm8oTGbGT8hyseBWq8q/TfNfgBYc4FQiZODEwRJ5DpOXnfzL6d5lHwEu1UtlvX
t6zQ5E/OAS1fmsZ5QU9HiXDXOjY6l2ex2RwA6wGa/cs7LnGu5jxemC3vI3jx2OgW
oneRM2ROSeyRt9h2vZgBITSpdF0RipE58BgVIGCjKn8r8G/kLF3UhIJkaiIMUSda
DMPpTnzkslxIEkB2y6vl4VI39NVqqaxTSedfH2JgIY/XieXNaXWAneHCdGES9zQH
Yq2aL6CYSZxWJX5c8C4/SM92Z0nURAoEXc672RP2dREWqiocL0bk7Vxs8SvLq1g+
YUIfTljKgJBRENAOOEWZExgISqBlaHQfpDpLn2fM5atdhBCZRSOqAvJCratbFzOT
vMTAEeXSXNR8UqKHGk5jbnmAXMCtP+u85kks5Xyuxwx5mtyC2nkuNjBadg6Ew9QO
dcOrQqKcHVbSTl69hHnfM+QIdPyZbR91HA28mdOS2zqWJmma8v2/vWhNV0BtDK8W
Xks9FazF6MpoDePm2gdxMB4lIFnAPhlclTYpHOjOix4ufjNgWSvDQafeQ7ZtX9rz
i35jr239EbBsAwrEJgYesbraDNe+PIFIOCIf6VFJ4lvtmS5z9q9NGBw5L5RAIB+5
Cd5oN4CIAd51ydRJQQUDHv8WmYISjiqZaWM8lpZKxCJi630I728Tyh77IXe3Lw2f
H3g4xpST6+/SCSdmV4578vWDzfC6oh70V9F2YSklYXfIdd57NQ3zxpOG+o1IXTtN
JVD9lTgw8zt7nqrt6mvGA/miAZvhlDVKLu+Mt3PPcYZZwSE94l94yFVr1MWW31En
kI3uYsd+AijJa8LjkIWlUhqn3wuaPLCF7jbJw4uPK8kWSBQsDY6o9xvveDXeVula
wnItnZHJp75sFJITYBC9k/lqZ8OtvPY1Lq5bn0TjAgq0FXVC2wElVuzoyKtFGfJ2
zuvfP+Vwa7lDdwCBTAA8QHXsl1AJ2eU3bBP9tvNxbadiiXeHEE/fPtMLH9aB/9AQ
Gj2W+CpjbcjAN/zEhw8x2gJJPeZRlhtRvYNndZrE16k6BfdJHiA2BoPOSRhsICNY
cnkZbl2Xc+6V15ulS4W8mSBINaDI834MQGBOewseDQtLS9tJe8+1EhrJZTneHDUz
s9TPWxUiFXF54DXRPMxAmDixwWFcn/r5i+xyGHba3Pn28ZG4NdqOLD3//vqpfs57
kfygnoDH3L9nDO/MtAGy7NaF51Wn7eLkcHJCX/gVKrZ9PlgR6l86gNkWp5skcEhs
xnMJThfXcorb09lRHoNStN+DjanHurOgPk/t5AaNa6QWly+XCWFs7CXKKJ/m7SYf
L3Ri9mqZBRYwOnNuXusN+x65KaC+11+4HOJDGhis3n5ZcIkjE1q84mrhgMwTLTgq
bdh/K0MQcJ/zIbhn7qcZy3/ii3SgS7pbGJ+pnE2pzISVCcDUXlAgfklZbmoPIpaB
MMJTJM1KIOrl/r7xDCvA31FCkHarf+NHimZ1WnLr9UZrdhpKORwWvEis79zXiiNH
Uf1DkSeJMPeqlwGQ9Gi6oGXTf/Ymm5L6Ct83f5e12i+S0CRuWO0SM1S2wRUz3V88
f8r1FP+XLs7UBD/nLY9Q7pFTBd/VE1a9UrHT4xPWqRC0s96iTwKxVdxfLpErs/jN
nV4RXmcA5wpO9U4AJ2gEGhLxUW+KMPb/rja1+GTTp8W5LWsS2tsu6jqC5+3c71D6
L5rXY2IYhPCcNkd7ns/nMDvqh/7/AgYEEc4gDcPbdDRWyGodXIif+ss5ZtNyXYB9
S0RrZaNuVRkBxus+A1E2/Ac34sI6MH+e1M2o2Ymb4nC68bumeZ+9f4nWBKcr6Zs3
rPSa7M1dx5Ow8JuSY4JhcckIfXis7J/HHIwHQARUg9bd6/db8rRrJPqbP7Qs/znQ
gB8B8XoJ/i8Z/cQuwL0rvJvynbCl1GcIvgbsd1UHBq2uGUQkiHPx6XZTlxV0oiYC
UkwURhpgLBULgMcDSpy9qqo983icifh5koCoVbzdXmuyOgnBFur/QyNKHZj4OmSD
BwBiJ5Ek1dEOVjutHc/h1pJ9pqOLkUGAEzcfWsfV51j6EFTA/gUmePTPgUVgW6nQ
m/I7MgJkRZkGluWfcJJz8yt2/xnIwYFA4Uk9x4Vov8+TzrH5bc/vAoXaxkJme4ZE
Ueh+14/NoOm3lqIjNHgw2CLtnEfUOeVmRhuneSAH6H+lMA1cLLXlb2Ttw1O8Tdcu
QLUc9hudyzkXMbMazJQAV4/1Pmu8ZiZLpo24HZm4f7om0UdpJu+1yi/833RliVQH
g1CZCRuTqUwYigyiEUvUFOEtihAflyciecT2aZ9xHKI8fWX3RssNYTC1GhtwYpuy
PHdm0ujRF3M3QsOzN2NsKWxslqRO3kvkS0V7R9+HhKoXq/NekXKEIYOvJomKkduv
bgFguEf/u6Z9PzLRsd0XI13eK8vxMQBbFlSrFcDEssfWADr1kR3KhPmQdGcTtw/3
bGTY0Myv/hDXso07E2k6IK0HPicKdQyKm7V9lz1fQLFVQlfoP7jpmH+MUX3aYevh
M+nON5uqoSEmAIdDjBQ+jHY56BA07D8gZhgxobsQKBu10Ok+C84hEHVKH46o3yxW
j858I4TpFPq/wK5InxwdMWHBTAv5xrDlBKl3zxAeg6gmS9HhZujJ9QlizHQxBeHX
Lanyn/dp+NUpXMxFWluDw6cOfomFSBqX9j246MdukVsol264nr7POawfKa4mvAtW
cefexbTQNUiV7ZEloceRiLDZtPETvo+aBsWw4hhgfvrFU3/NVNkHaLQJTFdWx4k7
TZxOl3o3wWhIaJqhPSciVnU9E8+mGDxB/WoKOQlNDf5ZjJkTURADGaV3L36Yfk1b
ymAdpi9BxOcySooMcgKexuSozHwscQu3BVaUfx+osVGeW7rcqTTRdrpVTazh51re
Cdjv30eUI8MV4VGFVi2be8bSx/ylxjUqrpub8p7BY7FxS2NmmAuQaAdAd3VKQMH3
JCC87lBwDlgnZvfTUWtMPG2LgK2hoyN/lQ6n4CayQLUKFud2wia4Ra8tezWplEbf
vsxMEOItG8N3+VGA0qZYeJ+nyWGT1dDdND7NIBpkSzbqV1WxeraymWlf4C8hEGIz
NK0P/QqpUUXx6/9+Rdj2QXNaAswY1lBrkKYMDj69TqOih6SMiPstvkIyCrHUZbXn
K2dhmo8Ku2v07JNZemqygVsFzMs2W4WESUhHKmZabLP63MOzk9dYA8eC8PJTeCmo
dtykHIbRTu1IhCdR68prEIz5OsmXZi5DUaqXp0ls/UDZVgLFGy/1+6N3/xZcBMTp
Uf3L1IJbVjdvv6Spmp6HOZ4SSbO1FH/NHVtQ+jMM9Qlwun3MR8J7p+UME6/rb56Q
/nPZUuSkHQydRzPki1utQBkCk2a/FTo4LOyJNxkQc9n5xybH+ycFAWxVfaPVDVUy
ZfqsjNNJOnc3IRUVr4w1CrubzThFmc3wdwFV8TAn1LZb+1qzzREFRutgN1Ht8k8K
ZMnMozX+FOEYO4uUrjn4NudxnB0OvzTAz4OzPh/0JNpBlpk23CMYQGoZ1zrAMwYQ
0FArICh05XBoVqvhSYPbSWlOhLh3tIqczMciZEvxfF45cvaMJN0tm791Eljk+RCj
quwTDMQ3DiJRQqMBLE5mvaHGVSrLW8rAYWfwXEKLyyH0BtOsbxswgFVKlmXo3gz6
nh2gd8s4pLBoAufjKTGEAc9qOIMg0D4Xpe3JqgGAMyWFA1j546CdpSdPhTgwV1Et
0JE64b+tkKFmTZM+SaxTQI9l7KGCTWqMKIk4BUpJ5sdgoX0W0ahX+IMBSNIRaNBJ
5laZ9YG6KRAx1ncC4DorfQc9neTVw5zbuX9GBWdcXD5NJN3M12veUfkn+X8UAPle
3yI9sZHgaIewG2elyRpvfN98GZjJ+q/wNdvN0JdYPHWHOFgo9SXDQK1MU5qmt+R/
jfSvLT4fk6yN3YGLMU04d3jeyj2ad+jlzL71f86FU3P2+kKGQ6Wb/kBcMsFmZHex
+T297DhaoFU9jXGZApLK1UHX07TlFRw6OQqsgj4WElPvnlyvszx4lEEtnEveXip+
EgaCJtILhls4E4C6v8BCGJm/OzimOuuy2oXowZif+l5uC6xByjF5pAqRimxrSb0K
ljlU8olVdSXfU1DMmmP2ANugcJYPCYwElqdmkf3skSAQVzJWWq26/4JAVs4MaSnF
uZCaQjLSFvHuo+sb/0OFQ/VQmcSHMc3YM/FuSwAvWgfwFaNy7RgQLleEwzhvGJPj
mezdZjOatPVXrZQFEX/47m2AubvK1AAXNqi/YJ0EDiFh2jzx2ZK08IPQWZB1Rjw3
PMFmLmTnpsazLDKj1JaHbc1CmTIExFV6Y1JlulKvC2HAHrJUsIxZp/bnVjPY6BES
Mg0vP3uaMxtzYeDaauOy4GummYiqNMg6/SfamK6pgvpqBoHW/IpQllVSAowYKZac
ynf36aSCE6aMFX/ujKQVGaBBij4sgVkUJlbKTOn1GjXtoYJq//NaQOTiipGmZjOt
oK4V6B1wtZI/BwBneJUO6O+jaV/37JjsndK1Lnt9OKz/aRrY/pYL0WgfbrkC+bYz
3pWWzi1PVTbr543xVPlCZnnpofkuQkalPvIFFmg5aeGM7aUDgjQwq6AP6qNVvnIW
xpUlly3ZZ3QyMOGWRNHbyVYk+6bu1KBm8sZ8sFt6m8zbsrcIEqGhW2AW1Son9S5l
foVlSDul2Rujs8ZIAy33dWYSakjVlEgNBonwro9xZfzJlhWtNZ3yuUQycDItnYYi
AloUMrS+v5zWhEWANKQF3jAEFG0eNLi3CZ4oUdetYchN8GyPxyKrX5JfherYFIER
pbsuXhOgx3xI5rM2d8D8iaGlUsihn0hc70loEVBs7VHSQ1Y9A3bFKw/Db3XqvYAn
IfnCpH4DHiYe5kUgzfN0EtrwiZRDId4Kz/jrMNAGt7MNUe2AMdGFeHofjXdVjqvB
egLZqw4916zaNgRDZwxGjTYWiVaMhwT8slfmmxTcTTru6oxxpEmB7zn15qkl8WfF
xmAmGgUYmRRfYFjYsajJcZnZhfLSyGEad+O9m8M3RCsvqI1MfsVp8AB1Goof6gQk
kxvXhAWgcQ2ObF11g7DycdYKQVdhSyfu9H/Os36gDmj/j57vv5bbSOGGlT+elrBU
ZPR8AVVqHQPP+n5BmoC+0kIVT506KuguidC2smE32LQ8+vwIPmEVufZmVQCauQKw
Iv+rfOXWM1YulKM78Fe55sKiNdWG69YVroK8f4cgGMhSIcrGSEiVnAf1i219Q3er
2vDxrelfFJ6oFIAJ6z7kPBkEkJcd/9FDyrX184LDVdkxsTAL2A9uqwrTz6UPiqjS
WTz8WQ6UwrgMYFvVt9mTQOPSymhcoCVFqrpbBpF4VZegb5jIVm5wANq4hYYm6JWn
jj/dD1fxMSzSgGoe7pdc/O3MadUnhZEbZkYQ97nwxhMHSmfJbTlLJfskpGFIjTXy
QYqCHnODf2gJ0IM+bUGuO7BzGKEhN4Fgh56CD0Og5eoncdAcy3xbTFEIPlqzMxhP
47GTP6pmKJ8uC10sOUdREV/6znn35CUk/xRXtxG+wCXSN9Mb4CiSzEx++qL5b4Ly
D2UAeQisd2P6UN7dfEes1YWtaqR5Apn8tlt4//nDFaf5pYsrMbiysAWaAIGHt7Az
gJz703l2dyFF+u20QQPQd8i9yaZeOzNuhNNUhp2uQ9JVB9u+MMaLszhlyckA3sNR
89otcuQAdekEUV/QL/vQTFtyHddfFhzm0xZS4rvgQ8uJjpgLecT5nk+q8MjAijjn
kNGHx4UoQwh8ZxodGbO7uQseNs2YlR9GKZ7EQpfgOhJcWNhoj4FlBxSqXGbDqhn+
g6TvCd/h/+NVmTZfabQhr9O5YiT01EaTy7iPe7wCaxDgaQjMbMRHEbfDY0hYQX8i
ipQZJZLA004jPHJS2QD2cgI9TdAZZFW8AqSLGsjAk75WE1Eca7NZeW6IwBbvrBfg
18Je50b1Ev5DYFbsItsPFyIRHl4YLNd0RrSDFtUHaUTulSmITLVdncLThYkUvqLa
XutxFHGgJTrsq4YOonhOps+2+Y9uKVwGVprOVwuetBtF5mNfk0VdX2NL7W3Mmcqt
SB9kvSHKmQsKqzdgaVqpu4z3nWWxxr60dITBO0FjM3CzK7RyRrLRWVHlH213LuQJ
xqAnTceEy3RkYsPafzFHE9qyXrtPDBywCgyI8kpFwJWOTieN1K86ql3i0VPiRz3y
AQAxJVl7y9j+OyoyOoE4l+gsRqQS7R/Z+xMuDS/C9aHqa+U//Qjg5Q/imaehAN/Q
VysQ/eOHeYbltCFxu2LK1+vcGMQu3O1ab/Vkw4seBsNA7iPPa2M36B2d/eFrpJi9
27TuD1NWK5QWDZpDvWJPhjg7sbexAa3Ibe/KaqlGJSIcjjbsdFLLEIa/BXNi1wKc
JnRhiCEP6Bp5crCd9kKeqZ5eSjMyPkZk9xsDhy3kmgsSR8RXi+h7AeApdYYVxdKo
UNlBpouxEm1Xf+foQf0zdH8hI+K0aG6F6SZfaGx7kJ5u9mPx1+qJ9kt4UXDmeKBa
Q7CzAU/RTjOXzoRLT43Y/ZTVF3Zj0B964n7Mfp+60G52SfCQUFUdaTHt5BFsuZdZ
zxAHiYLPW08Hukux3od3FCmFYUznIBTONn1bE3Wka2+jxSy/ahYbFlgYy6ptJVJE
91+K7dtTDmuOMcmZUBlFo8BgyzV6LA5PZZQSVb9WLkJ2AUUqeQDPzbvVDGzzda2x
PRRlozPWlcQG7IQcWP+neiJqrSf4timZbpMJunBh5jSC43eQ3NgA4Ni7KxfyE5jI
PqdqRnCyx5gCxqvDLcFjBVqmll2isIKaeAipJtdv9bosg/D0GhT3i/M7DEUswP2u
pg5mgZ72/3iGPIkw2+aSGhRlMJfFpdr+duk8MuKeG+3VICIBW2yST5JZZpaLKSXt
iAFbn2+Prcm0Iplpb9mzPqpyk98x0aH98WairTKc4vf4IDCGMShsG4sHcMjDt0W+
CI8KOX5g7POqW49zXe+QYc5VTBSKIIh6BLZGJKMqO4r8Kzy6HgIREE/axEzRYxVw
1oJDaM9mOZVLVnCQef7YxloblJEw/kaA95hkzRk8rO1e9M27ga/nr+9znTBhfMls
tMjF2dn655SzCv0uHdjigWR9Mzq5KPW4Z/IlrRKkGGRBqsWGBMT+idgN6gMCKWkQ
BgiF4tUF6xySHVVwqMrxGai84FM0izmMK3mfwUcfWZohMrRmclI005UUtUi3H92M
MepBc/kGSMVd9WSWPPcwyD8XnBB5mYI9ynNtGOGtjA+YKbOHLlXB90KJCLAeVayz
X3zsCla98ir4eGDoFG+k2UBBNIomZUxL91CNY19stwGj4aVVDdeAnkOiwwowaMfo
K2NmBu+iRCM3v73Zz+IEiiZz2RK24KuM1k9p+0vrn6tpU0638+2WJh0IU1g5dtBW
xRAm4LcTJaoyJD+6ZsrfTOLGbR3BWDWLJCj6xwmAfLOOQknfZz5w+U8nIB1MPQXz
7GjMGT+wYzxN7HiCs4Q36n5CGvGFvZOx1dBUUyIIaQW5UePzmAfHoQ7tMrRYD4c1
0+eYyH292cks08h/tlBAN6LhKq10+QtbJtx8f+zIed2NoR5oexSbHc5A8YwZY6G0
l/qiwQL/jWvWc8LAvSV0ZgbQo5xY0u+/gpA5zDZ0r9HNDmT/Mlx1aSIwmqeCsyLm
qg65xywSZlIs1veq4jeCwg5wMG2vQAN8LPKsch/mnHF3Rs4TjP1fQxGd/hG1BmJE
R1+6kmuDQArPc1gRyXxs0s9LiFM86ceUIelm14tfzVTiDJde+IOEPabrCt99bxO7
i/p5Lo6hdfB7Md8vhqBNerl4XVC3aWyWoRn4bpppwzxy78rijHyQY02/F6N+wyLK
aAK1zcrd0+3EA0uceDohO48vXO0AhXeQl/O6HV7gPHoj82MaCfnQ56F8NEMnZXYZ
xVXTf5D+yxP7oGGCcS6PP99usKG3/1fKwLO7B1MV0Ops2Kq5Odl/pBEw/GeS0STI
2234iGJeujrofDYxXEffyQsSTAJYgnQXKjqyrwBo7q/JWnxXszZ3DiMsxc2uDF6V
eGApDg2Urg3fblsr6es5HuLtos7t2qgdGpDPQiUXUfuiVMOeqSjNSMI9cl8A4q47
lPcbV5i71RLwGC8FOCeFdMSM9LBOE9x8WYax/8E1/OHF3HvfvaWTWQjTD/obVyIt
gjYXmBjXVlZ8ZKvGUQw521gLI1Kku6GfWSqEsHmY0fVVNNVWfohUsvf61d48F9hK
WAuYeTT19LGd8ThkYr6mzJYvrB2Gs+iffrMQZtJAfkfVVDiBDp3+XVOJOzSIT3jk
8BXnbTZjGJ4OJIyMbHx1c/EBiF+GIXAv7rwF2V5ePHrD/OrbSAFjlsdxNNIysHsO
CVuHiG2WH60yblKb3hndFJ7xKqMe8rQ7cV5A6D98X54z3HsQcd5iNXbp0/6Ya+Ic
NkHDWuE/49Vab9is4NltjYaVD6xcym/BZZijMcSw93l01p7gPRVa8igft974rq9M
EX5D8QLENVLYyQOvFtutk9jgbWxvhQUFWa4PT/uwwdkCI0JBfQnGb25J9/qyew89
UyCNeC6aFD7q32W7ECYMIM88sdHZzEbRy3r2dVxj3EMvLjmn/ra2gE25lua2Sovg
BkXgbKIIu4T385piamyPVuYqFjIh87DmFYYuY+108TFBy/OtdbihLVPjW+oSDc6/
Uxertkurm8/x53E+WtLoKRVmHTzL5vsnM/aShKNxFeCnjH3S54ilP7UTzhG5JqRE
uuiaVxMwpY9hA61mwf3grZiOJXEaDjSXcWL0uzvS8c71R4CtHSShici7qSqQ1AEI
SlscjWTNfaRn/bzoqbsBF7Xzvrqbzm6SHsIMA1HNpb+tkBRoQN8edbWePngYQQnW
2REYQWJhL6b8cKF4oBo+CZ+zq+AtUCRXd4PSyjexOiGdeaTJwE/E0w91mNzaEUFQ
KdTPi/deFmjYq0R0hTK4ZZ1SkVBASfBJR+07+U6nWeOR87pnINYcMmMVNtEBidVl
UenK0W3bLevAQnLICccNJQc6oLvrFc+3b2ddCSkjHcBDZr1i95TqpvL5l+vWM6TV
JfPwDkmVbi/3wTslnV71HJYLLJfmRcfjbg7qusbbtzJIMcn8yfqAMvuOPc1eFQ8y
wxBscGkSK0mlqdGWiU0cayh4yllLGtPh1rvPqqoOW7RTQo6T7LjlVhNmVLBk58qS
kxisa9nsyHTm5DesJeLbaAN7SXjhdjE4bGyw1l+4aZxRx0TguXbyfdDStB7muyY6
xqzrFKHUVRD4vZdeOPZIWbvlPCq+ZxLa/d5WVenRlpXow2id4yhAZBr60+O99woW
zbRW1GpI3BuB2AYBRRJ5hcjZkP3mo4kK6/9wri3BubxNimd62c9AAU4op5sr/xnT
iRnTGTUgKipkhNk8Bu3WTrZCoFL5656s74zRMIPt8C+DJm5NWGnqP7eMBOkP8v6s
hVjcuXMIK4L30GyFCbckoe3C6WyNrekOIhpoLXLVhAQiAO0QGM6xNSvuXVj17tqN
9GZ4+NXODUIS8NeU4MDM1KSQpBGmJgebheqmLtIT1fyHXA0NGMeL0TOHgi36yMsu
+sZUoAERHgZbpKt/mlYwLrgAWWK+SdjtW+DsKOsNph/o3TraSLbMd2AIVdWbWsOZ
98zzmO0EVENEJfCQt8vqUudpAD9DYC2CjE1WNRXzs8DpU/xWgSx4+wdRhKfCN9MR
iZ0HnAEEvQI4z5VBNzEfFoE9NYZ/ntsrEYPdjk4KcQmZinxCuroNElOtKBi+S6Ij
BKBOHj7ZxXsfgfbh/eHpxGi4MBqgXi9Q78LjD8mwAYkZnOHjlYu0ABZM9UmGZ8vD
/H8UuqIjwxjtOFHB5hPzXU9F9UUz4d+m1Az4cpduF0QdMjvb5U++1i3XHJDBSHo4
f+ankdW0SKQ/yR+cChEjLadBn+un1QWC6+YypVAq1UOZcA8Tivn3CqHrLoj5tLDd
i7ymW0cK/DzLsfxfILv+hGLrI8C7b6qRYpNP22aeXe9x08wRrqRdLnFoQtRXTlH4
ezmxWO4yGIRiaBNr4PX6uAqji0LU9J2tThFQHHUfDDbyDkoVzUk6kXFhzksJQAJe
Piz4pqiwjjBY4EgD9uxbM0v3KZqyu5W7j53rOEefrYplaRPdQi4N9LwJLZCKRWiC
QZ/dicny9V5LQtzumCMi7J89naSHXk+D3sh6mQIjURDH0maZqkq6eLAtus5GeriT
YPoDiMQ27qMOzD5Oj4VQXX7DnjWmx8q6TbUEn295bBhciEccV/R25wfhj2PKj0p3
FBA4qozZGl1QAM0r/rCWLCfG5JVoK1YanfXrvERL0JJaPUcklXmidvUjPxZoPBMC
VGAh725j9z69BFwDljs6lj2Dh+hXKT/2Ola36WxHyOxsAiu9OnOL/nEu8AONkQHf
x76aZ7efZy7BIOHQD09n8V4LtTE7WjT0t4cirKYGsKjc0YaF0yMluujsvrbYzDre
nU2GbzSZCDL0YsIY4RZrnuKc/NeOR9W616BxlpxkTpGDPpps+7Hx4LGyYLNcfXoD
5m9QYGvhIGCkZxmJP88I9/QSGn2GHwbheTNw++YLrFU6WFqjdVjMbKjF1KARKAQV
pXt5jmlCxVdHohSmismSs+z5wWF9IgvkOQ7A/zTXQHWtdHmBiEScWkRwRy9kvNUF
NLWyNe6u5pZ2xa0DV/US0iGVCW5trqongQY7oqlP+lQUeMNTkLpOOsFX2+8FJQR2
6Vuk4aT5x7qJlauH31nvc3KOhrHLOmonqJkCG+SgXUreVH0t7qXZ5UlrRYgUwQnH
WEkydR80IxM5zYh+HfzCDRhoyON6qGYKXuuvbPlmdDDdXhVaOnNJH3Qz3ayC8LhA
6IHPyAo55PNCqd+3BHDbCkTXHyvEM/sZAzgZcbYWzoGMhHEV1mB3aVQ4xDntctQT
6pz7YIUCKmtsvHF5Dn5CQibO4fl+qHh/bb1Ft5aRc92208FNjABjSSAQXE9K1RuZ
mzTzRGOhyNEJy/jxu66Hck66Q6dLp9OrD3RECAEryG/hHaZfLPFScqeAf/r9Z0LH
YY/xYjt4ChDXlM7Cjtt2i4qfgnmNQ0e0FYIYClctNb62+otVi4FlHtTd5tF7/KDZ
p322rUNHUZP2cf2FcPBQ+cmuzEYUPlCkhfQunnV6pSMxUFLCMvwV5bLlhNrClCjb
9DOrMZ9m+DDkmHBJDt0GiauhuFlDYV+IpLNMgpmjob9kyVFAB0e/FtvDAZvyTLMl
SshDDdXkryU0wQKHYPyuSPUl2TnsHXdr2cNnO9HPe7hSGKH2EVdQ+YQBAxaAYvWt
dF242yAfus9cMgHHJUG4X6DrJ0qLp1iaOD/f8T9l61YJZGaaMaeEYNxcEEyWzlqV
Vxbz5KSDZSZ5OSlAjfAWOB4foTbcY3HGo1ATlNKz4E32DuzQogVDI1f6MYHq083d
XJNKsUEdXoj+poAm3jEvsrnMawO9h6RwNXu0PuUgsnT+twKg69Kgyftnnd+WrmhY
6ViR2X+ixm+ojpAvSPSu+5RioUu62YTxzGloMZkx0ahKkWdaj/cpkuQEaeBb/Gzm
LoSrV6ls48FR5asDP+cjdflMtFS8awu3j2GcRmlFHSxWZIdpQNO9LaETBabJ0rBF
6yefZ5Fonqn+qTwdYQyDJOOt2OeZApQ65KNNQePtNHRicwrsRRBJSTpQNWbU7o6h
9bRt5HV7BQ4ORN6FY3V00o8HjrYdl8/Yfc6NVER+xE7j1+PLTVNFFwr3oi6D25Ws
aoiJ11urXLnp/lCKkHFpQuUJ7KVw27/wSEWbNLKfiugtf48fcdfJ0jdpU3HwxHnP
cT+CcHUIeqdGqxrU3EcC+yp1J+4LJRlwxQIcCJcgvaPo0q/kvxTTUAXlCfzLXu/k
x43lBMxC1zBU4MzoopJoAtdRFeeD7vAPtWNmipg0pXgHpu7D1Knzy4G1J32dfrlL
IcSgAG70kp9WtfMKo9REYtFjmkDQ1wp8W87sIWosj5/aPEnbNu9tbIKN4tmP6XL/
RfeX3Ft8gNCC8vJyDwBiZtpypiC10qre1DAdtDrIoo4rZf0f0F0Gzx1g/5Q9x3Pq
4Y2hRLun/+iJ0dnhCJVx6CKXrAmUEgqFElvuJsqLMMRpxohsg60nUJAGUWy9U5sn
M44RT7VE1DVJbYHxshtzY2V9JULNqKJcnzssJTxl5TmBDIlVn3SRySBUjgk/SCSv
Au5BQpkjikEe2ZvGi37RgJSVknCGgJHV32dIToQWeMX09Kz0rqAtrePYZohs3YDR
8zcSIt5KrSjuizAnbNQCdTyFJm1wmzrMGZEaB1XMzkYXwQqoDLMiPRJ7aqxCH7zG
VXvUyEShOU60vEng/lhMiBTCT3h2gYWZ5ypaVLVfFDQKwwYi9Bwv0cSafyzTzY3P
DYRhi6/Mx/FAbrj7L3Jm5GyXk8RYCfAWp5UaNAaRxd2r9n3D4SLVtiVPaYIrHbHL
IM3fDQUgRayXD9CZxtyEYbN/F8a1WVGy46+LwoMvxSqZRsgjom3IFrw8bO7ZqY4l
WthDt0O8Es2JwR+iMTDEoNqM5A3bq9wqMQ6UszaF8yj2nSfqfCfvaYSq5Bued623
exzJYk5c7TNyN+PaLzBkSoeWmdFmhvpbveb5XnvfqAWE1Ro0Pi8oD6i1xeCGGKcx
nUMbz6SYU2xe57gGAqGYgxDZIZvr1+SLx8ATA4QkTkwtdGH/tevz9EGtUBZdrHB8
Vzg1oyKB4MHVm9YNoqBnKN3Heiu6KkapTRXzwKxNxdUR+VUR+uxsvVEb2WKPNmya
Zt9esVx4VatJjin/ivrrwdhdfqsA7o8Zj9pVT5chYfmknFs+Lw0S9UTSymtlsWit
swurLE1sKAH+kM0pk3BbF+78pYHIngy1WBOg7+3FDWoYCVFUIyVSaLPkjGWRGic5
Wk9zEw4K2AdiZmv7M4YFYfZeaINVrz55vPFIPvF+yR5RM9iTLIhb2XA5Qjs9QVOh
znIJs/+TEutF2hTc7CkQEja1ZSiu2ZiwigusHuXbYf/1wE4XkF0uLwaecWYysWQv
6m7Ay9cL8NBIURumU7M80Bh4eoV1MzjGkOEVGNCRFyMzOn8fTJtaCkcoH4lZq32X
7CsfLfCNiq4jOtgRHuKy/eDayW7QUZXlMcNICOGl85NqLGxOk8Uxu5flHzZUp8O9
VHAgt72cugUc4nkA1c1jTWvi8Z/gfxwFaaiYENwCTsQqXGDKI+x9tX710DuzXVxN
9G7zcueRebHGQudkGjhsQa1i9IsNlHoEiMutTH7eHsF/pvEYxlbh16DFKcY+LaBy
D/KeJb+OurLkw2MACdr+00EY44DQdYMz+S93ydiw3nbCZ6GIPdsnqaGQG+LcI/RA
VFq6LoEvS5X6rIAnLuwJ0RMnhWDAlE//wiyY3MYYjzoo+s+G6vOWfUUxUxlmEo/J
EDSibl/Zu5MkLc4ChF9uGoLiSE7XC/2z5DJ/Q09Em5pxyUTPXzqe/4lCHA/0k+KC
ENtVuDMS7IFMqAV1PiuEaykLG9OzMcYcaK+l+ySWeDQ9/tiScjVdlLCQHgyYVH+w
OY1g+F128WWUoWTW09zliDLm8k0I+77hzdSxU2qpnQQdEij0Lp7Iu/SxQavKFfVQ
8Xi0jmUG9YmxFjg/YXsXHta75fk3WJAzv0UyCFFssJi9yVaO8pN+wDxg7q96/eRP
hmm6xQmPufRLk2FSMwE0mE9Rxti5j0avSwc7TecwW5D1u22HuJjtUkJrCYxwGY80
i+N5d6uSq5l/3FvpAMTg+u9wwYrkJV/m/qRoQHzPC/94ILME333D2rAOqOF3paD0
E4XlogOlgfoNaV2hWpXe06zRCHsIhg4hwlEuwLJ0ZWoozjDzhep3lFV0a0y1Ds13
JRccwgIVQpCJJgfcTwD1gX9frttwXAcbdMrrQB3LN1U+PuOmNbhQQOIj6cry6yFq
jahFJMvNegt0dIUvZp4/FTYY1cT639TZY+ae4THAtAn2VaCyXt3EK1D5UlP4XvSa
qsiTc8v3XYqx2/UXxaNVuMo8t2OMcWAUIDkzab6hdlKvl6yxSD9mdAl6It+vMyt+
+Qzq2PWr7PIjc2nMW8Nd2D6UzTv8NMrECYy+FT/ypl6V+a5zvEzT8J2uU9ANK+nl
98V8lXO/DdQWUol7lhDfGs4EWBuB3YnrhoJNBmgewn8zoQx/Ytee72xEVkRMjkIP
73Ev3IPTNs+xYuOaetLLuvHQrPOzJH41edIVOaldgNBqQZ3sahFk2F4GawZxepbZ
V5Rqg/OxOEeIsVUwL3H+A9VI+usvowIIJ8TSDGJPtpE/CUSeLATlFCXKIEnmN6TW
IL7C5PBXz1ynocLay6ih56cCihpHM6ZJdADFCYLZnizw852ztJFyLhdvT4wg9G8j
ES/k4KqYZUASsoUJqNHoF/PvzcbO6KQY69JRVEp81/eYzdTXY4TQDwAp+8gcChEG
PKGPgMQOZkXEFeZRY6KNKL6j+VB3fuNyr8unxYm9O6NFnVXOkrbbuXwGw4iqR9qA
H7pVu8dOmAd8Vxc82Ru30rCAREazqTon75pLkt+RbIEOYHnH03k30tENC1pgmnaJ
DOqJ+pPojqcfgzM23YxyOJ8MgCyAUWqACiOO710hZuS92BUKMV68SVmLsweJvDGu
5W8p8Wpu1xaWAKNja7U7QDHPFyPehqSmCgGXSrbyhIkjp85Z7AIm6Q4bzypcuu+O
WURZ9LWTpz18WgZ0rOAZ3ySwpL7eKhS95Eqz2Hm1OgYtps57g0E6KbsCDfKBcnqP
AAJC4Fusb4Lk7xPDbJ2quGgNdL48yhU3L3u+m8EjWzNXI/GLborur0VeO++BPsDq
3SWJ8o8yUNehzvLB0+jqCDj4wNzprw2DxzACB6OVxgYHqD24TFTsjSFLneYRWHS5
IBkFCwBlYTzhL896R/snO2vDU1dEnaKoT1yhJtT731O+oLmSgrd3NhwITeGAh826
TpTxp7KwXtPfTqU2KFqE5aIGE5hkZACI4X2oe7NDkkTBLcAt9+LrUHe9/GCbR2Jp
yI0YqA3aCzv+2kinOvWuXAVegTLmD8SFMDYbUah1whXUbg1a9CfpmYxImum4/j5q
kRzv8jTol7liHhgolL8FDYtWCiNK6+FmVJkZnWC76vd2IRzjvyIjmVadREuimpoB
87JxC0qB0yTzI8kJnSmP8MRt6I8MHVJN9kA+47cRIMQwE7SqMHJZ1SSUnvNh91/u
bJLENPPyo/u76lmEFF17g1DSIY7tclMjMh76MMJoVSFi2BMGlLNDUzmZi7WXaS1n
EunmW2sfZ2EN3O4wM8IfPUy0UKi8FfooOZa7vd31+8/tETngtEkENwD/jhrbwOxb
/qNuC3uCrKDO+5shT0vyy5iG+PBoGpaSoal6x9ZjQNHwJmF7fV6d3+eDiuP+C2s5
rLoHBJV+IUQVoNgJ/Hxw+xzEwg5hU+T9BmMtM6bG32XqS5MzY+6jjg1FnljltjnR
S4Nf3kyFMAwD9obbPjW0FeNoPHSHoMB1MQoloZFS+CcvjdsVzuOvhyNRAApd15n9
NsJ+V1aWWPOMfQ5FyDDk1+ebtPKMh4ybKNI8FK1N801SkKhI3hbIT9J0Jndz5WRO
hbzXAJkT0NahTH14jIg6VhANcgb1PpFvTqwUfw40EiDR+vDg3KluBZTugA1X2BBK
e4nTKF4bcllvht+OQRfmpBmnRfLINH6oKMGoaHoSZChKLQtWhOqOxjxKOP/hIgMC
8iJcqWT4hcJmeb68G7jNAAPLuzH2gSzWq/aswof4bVDC7tX6cRJnLlJ3QgZ+HnpE
iLZbGWOhoyxO9Hx1c6DRaa4nFqLFcZKEmEpxOyNHzN9AtJZ9EAMma03JTw0tcoj7
J9rlUPRrjPjIIZN3Wfnj/7xHyXvDPiUauDVmhQaAneBpUz0oQpfxD+ErPoA2j5AW
OEbGanH4HZsn1/9qMRiRAXzAr8QoWHvGJD7R/coOSCKDT5kLX/PPDrv/BH7GvBEs
AowotqneWHieKn4VureYa4YZlbm1L5eHacrPpmneBKXVRHUGBnenRThu4f/8wQ3c
Im3ra8rYaXD2Oy+qI85PZlQYNwIBqI3Itb/UrEHBoNeew4Flfdh/T0lOJcqIjFqd
LOkf5De6UIm8U8i61Kfol982UEd0m5hLqoefAPR3f8OncWaqSSJ4MQ9wLXFX6XBT
VorzB+W4/FzHZtiL+QX956nvbhw/j7zLfcSUaXvRnmuOEO2yDgWjLaJliwNIE1JU
tQU4A7a3Mro9c8GomOiurt870+rmv8sD/03RMamIExYLHpjcAqpoH2+RH0D3PwHV
S8vkKkWHQqEAqzkYeDG5aeKBTiIUmHPd5Fr6rKqx3d4LSqbCQ11QTuPtOn2ct9eS
NjMfBYbyRQRoZvUF4tRqH02du8dLutLayE5787fe2rLLjb16J/GFYRkg+WnuBA9Y
mbVwgrsbdidbBqVcQNx1gi9bFgA/4dVzB6LUAWh8pWe6HrlzA2ZfjtGH6o6sOAvT
TovQGjl4TTmPi7hycxeC62NY5eQUpqBtCABVKM7ZiQH7uNNIOojBXP3G+u1nm5Az
G3WzpuhWUdXhB8J/cYj4K/Zqi+FckUA+Q85DkUVmCVBrcSQiNpCY+8Zkv8IzciPu
lMqggER2yvYmiA8/DJe4IrzSPKEs7FW8oOy/XmDjlS2dElRN10+XLeWJn2CT3PdJ
YnU0y7daHZn0i+4x/IYgo1nCz7ce3rU2j+JMvd81T/FL9Uha4Gwu1N9O40gmyAmD
NPC0O9REuN1E5BL1ws8XGpYWxkvSxOe6BSJYoe3xwrBNgPmZaoLwdO5KnejkGs+k
vRhznwnEmlFWQx9NRTM021WZU5oYa0ZLgU4oNtT1iCKxBfmgdyUjbrWxURKqsMKW
rRxQnCZPAPM9EcwYXbvNp3Cq94bO11NTsn9c5HEHds9JOIMKPjJHHE2UqGrab5gc
WsSvhlxtrYevO4qbtBr8UC3QTK4YjWzeFPFMYN+WJZ9osAGwLEk+IwaNIXlCQDRK
kAGNvYgXNe0wF3YPYlOlNGbq5bQIVgAFuipKhBs+UTrUIhHxHlp6S2aZ4Uvgzhgf
4aT9eZc46fu+RonpC7zz+llhpuBOSqx3l8LhNNEwIbwVf2xYIok2iC8Sg8TvxITj
pWBL3i3k2Eyzgz4yZyM2VwFO0pS2LTmfu2MmNWEoTV8sbSpVEOfPdFaG6p9+Uyf+
xfT8OBIdEsw+CHt93JPpDWedoQdeYRTNtRvwb6Qv2zPjEeEVBjtJLrxEziv2R9i/
SBN4bnhr5jQ5asdFRVq5Yju7PJCfNj6jLw1DK6VfVF5n/W/aie8hx+qxHUUELS2o
Ah3DXgBRNJ2IGRP2vRV5mKp7bpP7wtqoJ2Fqrb74ZP6Oy2z9hKk3rg93QLCeZ+Wv
6rOV2M0WmyQOteHwc9U+2kx8oT6DjWgTV5/Pw3DDFlCvziNE0PsAQ7sPePA5qrYA
d1fp+VSm2eEEDvskQIrMcC9nbxHD6PXiWEnmEJvxT1Nm7eLw8xTCJtlcKUIR9A5v
kV5z56vriml9yswKpPQWT+ErwTMU8gSqEyV4gLOsLJ6wjXTqkqWIQZFdfDRLzps2
Tz7enrt9rgzf3Bzm2SGXB4bq7pOQ0jE43XuUlPSDLBil7jIbExybym035WSRrwQ6
iz8TRIJWg9uYSXGAw2EMqOq0BqPd5eaXn4ORU/+MqZ8ABMYF2SZrxDg140Uso59+
JnB2kmakCc+H7bHliGSpFyIeYekp6EPh+0kqV7eab9vSOzvOybHzgp2G8iRZAl6E
8gKPewc2/r9hJFRIXtA9eaVrFxnrh4IXc8H1+K0eU/qVdEKb988BZYnDZbDd7UTh
kYPIERsJ5+jVsus/OipfNriz66XaQTWl/ZJDQKW+zeFu85owL01Fvb4tkC4IfaFN
B3P9XAICXV+osK2EeZoLp83PkWSysWfuFOiOgWuGq885gfgELmOyHIFk6F2zBlQ+
S1VdwjLLm+dE4C9SJfGJtOIHL7ba25iu4zjfY72tKL1PtrwdPtX2EQ/jhXaIWQZ8
A78eacGGj+4R8rZtdXqAbbJm9II8T9veHlcc8WPmNyZI0dQja6h+6XQ16X68uY9e
6Czl228L/fs7zdaybvibWuwabJKM4a5pdX7/5doqXMEDQw3FqplzQoztT9emd5cH
3vzCyQI45Ao4M1y8NxLbNPKaJh9SjQYtFo6vgsir/WEKZehlwJNHJcjT/KyZQ/wl
0Dz3tXQI9+ldLc0UbUk1yu6htzZxD+0Xx25uGy577H59dCpNdZ9KKdwV3pqq2Jt8
t+QXHXJlS4pNGA01q04xYHwjVaEw0AjbRdZ8F45snzoPS6pkJ3O99Wet4s4hgC/U
ErJ8OQaswqfjfA4LuINugwQxVYsTtuoW7CzgWQ1NS9HALZvWlUrlK+Asg1U+uhLK
HRor/xrRY+d26O5c5dlgqV3Lmnd/7/BC2DqdYz6095/hsZw1KYkRIL+asZ9N/UdE
84XfwCCUpf71GzxLkNEjQXbfqM70ihyJjphp/xmJnzti5gS4NbHLsskNsWvjK1RR
WFIn9er9oWKrWqYgGx9PZzwFiZvZdg49MZ5FDAaGsBx5jCpjnS6P9L4J9DB04lUu
X0tjWB18hcj2mye11KnXM2tMWrj5exFKGWt7KOhpC74kWVFLjD4vsrYYDwMzMkV7
r25IjIIk5YCDqAqIjiQ0vLhkyEYy6f3dTMhe9LLWgWnB4J7Ki6zJNpAC5Muzy6z8
c4OkuEWo59YVhmERYJ+eEx7Sb1cxvK21jwfuXyOmoskeTYG3GDrgpH4htkOVfZiy
Cdmm93XeWMdG6BHo2uVMdCbClUDsop7nfbV8TMByvG32SsdjTugk/JGOaA6gRWCR
AZL3EI9qHNUDK0P9BK85cFuYGkazE4jc/xMlQcrsjNUydQ+XualFHykpWU9cuND3
lSOvKoqhrkx5bkrl+7fnGcxhEHS8nWxwS77gpisYwrQrTXAMKN8iq308nrcVCm8f
b4+4NU/jA6JmuUkAPCbiLQs3blBGncwm+Gu7rC3XiF7/7Ra4XBwx0BXO+25F616/
5HJQibDTx4Qg6XhZgDw8BwsZQBiUULD3jYRI5qhbMuKN1hvXuCbQkDB4+7PMsojp
0kMsT2GaF7469ecPn1I5Mo4wERQFRJ06TySaThzuIYBH3xbQNsRd4rqJchI+hfA1
ZX4ccXdkvLEof9gKElmCfxAM23TA+cRZGN7gAhgMTJ3RpvYFXNkYjFaRa24vnO+m
t34iS5v3G3Hj8YXY69SDI3UI5g0QveGnf7RLkGjgrnYF1kL9P013fxBz/MdHx5dR
YFdstnbDO8ZHtbIwSEMdY0D3k5q5uNwtloDOgmmUlXt1r2ZsFbWMRkjSNgvR43H0
SCRHq3qfxyqeOq5zf5HxFeazlJYcT2DFwv++TNgo7kZVtDDekK5ArhKjMQCRt3CK
2BcCv/FAOxFxL1qSNNSc5DvVd96HwS6/psnEQQCROuHhqFOj544mO5CbEyuNTAe4
czHKCQwaND5EdXOIntwdB+qztxJwPbYgtJvMyOZvuGvs9wAYEPGJ3OOz8A+Azn7s
PY1V2BttmDw7BVQxCFBp9ppNZpsZ9r0bNcsED36jBWXoq2ZPOeEfqwUOt29RQwu0
77i/eCqVJIMu12qLEplsBsMGQgT0CAqYDHN5mUzopHuLwGDLD07J20l+CwMLYKuU
RWrcrHf8Mb1MSBR12d/MDo+6gc7XbsUv0jTMFgf/4rT0EQ7G1aP+XaUEbj3XEIwD
bJ/viZVWy3nuQyu/3VoVSGE07vqVZpU9fB1EjcR24DZWAeobzKgdearXB8XwigpJ
jYvqJzHqzOqVp8YBuUD4Uuo+mPJFGmjR1qqKcosJUbQv/r6ZOUJiGzKrvY+1i0QZ
v2wGpZR2y2DQdau/OFg2Bi+rOhA4bFsPVAKomFgvAijwHcS+hlqwgTBNzvipU5ly
OOLOynwkhFWIJjN44Z5IOt4viWPSZN1G6jP51pwoDgbdOvhlM3qI7a4IkxemWY5P
Z678MXjSMqvc/Oxl2qeDXmjgI2PERciNAl7qHk48SPeFanxxzoaM61Jot/cY4Jxf
cN2ftV1OaqlaBUawgGRrW8tUQJR48Md5x+TroK7HK8TpDFS7f9lm/ZFj4n+qWnmx
mNXc9do/+XRXhmYPdGxkdxcNrWUaHI/HOXlWmqER/plIN5H0xd4qNf7Q+3cE2gns
uDXvresj96kVzOpAe3anx7TegQRACPMCrJ44KcBeSbIbAPHdcVkQ6aj4GmsppHaf
Df4r8A3tr8mCXZt5Oz2mz2J8t1fGJtkE1xx+PlQU5cau1QULofhhaUaNrM8vtDeR
2LvcG4LDymcPeRrfClWISndLvzMvDEOY5VuhvVDm1BOEHNZK6VHvc8q5wMZ1tQOJ
j7APQU2SoJvQ9F6QrfmOCtHgIMtkPyoX6MmS73wti9HMliknB1VU71HizjfDaba6
EpCzsQxlCVKqpxDg1rN16nshphMzCyXQSfw2zgINld3utnYzgs/5a2MeR3dLmWqZ
4obBzhsk7o1Lh52XV6LOqRR1fhPC6StyjslfFBv85hA8FJIbFUsH4yi7t6OvoBxU
QrkuazVChEwRbi8Y7pR6tQqZx0h68SoBFFWfqyJzNf4R7dun1/ndHkzTnoYukNy4
GYS+6vWClRNMM8Beh5jSnPgzacazJRLsTHHQCvNKPFzohZZcI0aD42pWhTEEL/6L
IATyDywH9bwCNI7Gnu8CqVXKONohNpILCmyeuU3ZYfV7ZHy8ZeN7DGb9NK+ca0pQ
F1QdeOPbX+/24RobqFUOgGp486KSyHDO6Ik3aqGiqYQ9d3TfbTrj3PM1FCyku2IY
W/5PMaOAxqL6jFZ3lXOtk5c4Y7Azgw7EohQNobUOXrxCgMzsBajbsmfzh4ixNE48
ilyMHVrdC9yZ9gn6NODpUsP/IHNTSXQ3YQj9JTp+lIVl1TbUtJPspYjU04Vierhc
3spV6OFCYIhGykuGcu8MosWwalovD0UADa2AYbdIyx0fgpXMSZI2eywZhuUlMxsC
Al8E8FRfgFBAHwiALFFg/bQ+iBv4prg9ONNVfYqFJ9uZ1YMng+n4s6t/cA4wyKQo
NqXg65UlAsyrKorIvWuu5bc5HMGEouy/QEn7L8BB+KWIO9QK9VTlmJQ7xTduKhYS
seHmMZj3W4YxFivLBPdUGhzKGMzp3XeZaWRnHjBERyy5hKcHy+r+R+i0o3HKJe0L
f7bm5nWPzJ2bTBJ2B6QzIk/R2LTKoN0nhI3EizHX5OSgv/rfqCR2i535Oc2abQvn
tk8bovWwwMYUSGFcdARFtPuCJ88Pmmg06o14hIa+dGpuXk6mqj7RB/ZgsnDJEXlm
024BNUlqO3Mb9ADXgqBLf18zwKFLMDFiuNAji3kgwMLW41vsm/Tb4tZyghZrZafd
RSeUhYmJIdHg+K1Npbrrz+I8IjsB8NoJjeUYwMSpHtQCl2kUpcfgRv7cW8iCy2sg
1prCZRaUPh6LvRCw4HP1mq+/bIlIP01/UQgL+vLBMrBAPN7h28QX7Mgf32ffNCLr
WNAIvxOn1q0rnSeMNGjxzdDVhj1cJ4BLgZhgVBi8VjOeaZq6+0hAAUYrTYVYAt9x
4GuSzVx7usZO7qETTR1BKMPFUeoUDY1zlqSLtNhF0yTOc/tZc5kSggewDcWOTQ/H
eQvfKLlrsdiipFi9FaI0K4ulmvf80IcT0hm/m/2JVBBGHoP5h8D8j0+Kp7uVj8OL
GsEsKUE1t06obXr3YGQO86eNERXuuurJbkMsVZF8aFY9KVJ8Pg6KZmHqwG8OuVMe
YlXdu2Wbi37xusX8oamaVeSw3fhi7mCy7g2Pel2KVZqhuJE1Cfd4VeSLrzO9sJvz
XeNIyhVsMUkAZ1gVXCVbuxulqZRQXBJ4VpfaCtzD+AfT6gkUM6gvU6CkN7UpX4WU
IlbzXXBjxrGgMAgZ4nqSBkhFFIlofGZHfJAAzy8OEUhNc/QdviccGBsG3P4rP5Ty
xMV8i4WVnT50tlr1tZc3DiKW6CxU3cCeu3ruSXVRh3qQhvto09m/X0q8nuuRYTbD
xkQpEwoYvI853DIc+S7bn/biNa9VezcdtzaAR2RISxzwWTOFNiDJ+GsqY8V/v2UZ
43zK7vr97vQDKCubQDhPvdm12A8PBznNdMUx5b9GYRLpbhVuTHtbezvjSN+XNvS8
v9G3wDyVdG1KUcUOCPdAI/x8WdzM/O0GxXR3PE86mYlWFZXQa9nP344FN4q0wU2E
Ar6wtkBkIVaHrz6nvVqIGrUqUrKX0wXZblv5jllZisL2lWsyneExIuyWWS7lJTpX
yo4BH18HCoujuL4vW+HW2GctOSe+tklXAvFUhJgHmQtRhAzTSPUYw1WvyUF7UAAl
8r62sZW7NBFLnxNN1FOuwdLvtkNpu6aGql55PmYcKX+yvcptsdqiJQ5zn0aYmQEA
EV8RBvgCvr+exBo5xtTPXd3IpNBHMkmcaVjTD2HWftK8hc7caJ5PfESRNit1ZlCY
5x7yy343tjHoTZl8beKgZzyERvu+uchNzfFgz2+z/qrHVbbGpOhZg1BQVNqGgxZL
GE4XhE6M7XG7RK29YISx0FxMDMeaz//RK/e6vDBv67KL2ho2DiUU06ijrzAOGkap
4ej+3tfAO90XCfsvTDzbrcapZ2mau+MF/1OsrTxQTHlUR0KRfjpveIK4ZzfnlpEz
WChFYvPRZ4e75IR91IfBpDF/Ks74PlGaap3YkXj2H+gtaW9gsS1ODgwZwJOv2BWU
ceSyqPgr5H2i5SCw1Xb6F4zlnycu7VXRfmlCpb1s6bKaxefMtgeT+SSR5UeBKUE9
lNAuilDBdCwUqE/cYGSK2mz3azSmvHFIRszo9OL6yP6BdRXOdE71Rrxcwxc69hxx
erBOMxw3OCXUaFqcHtTH0E5dLQ83klA/OenZABgzndMSfGA0s+EY4hUFBcqxyCTF
5U0KQPTcGL1YIAvq4Jw0BpjC8IXwOcdVloKrtQhoYUITGKlJb4OrgSHRB8jm88l6
nc2sQLSnXTjY68j1eRozcf+ufVOQJ9AVJZ1Rbc2ib3ie7KjJiOTcoADiXPjEn2mr
pMS0tOFNYOKcGBDVJrVz9OVefXnPrMfC4dbau/7YywfPh4TDRqCAUujAz9K02EbN
SV+jwHKEITfRxPFXGSu/bL4QFhtPXq6pQNL56T0+Lu7UvmcZ4TbE0Y93WdAeb2ZW
XTDD7WqSQ2bvzSgVHuzI5EP3aWEdTejAvWBqYgbqlG/LwvYaD3DJwcCsN5Qm26Yv
6FdzWofIzG93tmV0wwWo6vvr7lkg/efzjYhdRlI18wZN9SWWclBi6X5J3WbDsbka
EltvbW+qZ+WzeqxqhmcaQ0kyFsyeKLSPK6p5JFNhtlqsHGyO50Ok3ApOaNAMi6iC
eXtkQf9Bfra4D/M5N3MVS0j9PAhFVYfuFfti5A3jig31JyagGdg+Nar5XT7wQsEO
19XQXbQyGIWpLYDcplfHFGOl+OhxiEMcKuJnaFTB9ELIAbUfQxN4c/VXtcGeCKqt
zbrFQTQy4qpW91WhxHQjwTdUCdLTq+1nGQHV7AI6Gng9vWCz+VpGAPijcCz5QUeM
fMQU92K3l+eG8z+MhUqhkyNObThPJW0gDBRJS2Ss9GxVlT11QKMS99WxH52l+CKx
7Fj9T2eZSfT0xNgfYWByKg1v4oPMA0EBtq8OzaFb3PdfykDduy0JwrX/7hp200EY
kbPdbl1TgSNTigt0elxei2NzJESgTHoHnh7KMWOwaPsAe3W5jG4UbGVv04Aakzpt
4aDr+1SIz4IFGxewN3V6JrPTKQ7BtGKqCYyd1PRMQE8VhJZCmfx6Q1olS9AZ+L5t
QBP/yafWJ4GOUwjlMKQMdhCS8uX1zM6RJUsMa/l2jaQZ8TsvKDzgHwLtwNcK7KuC
k0PUrR5e8EsHYQ0H2N2gzKGJayrfGaK4f9UEKxQ02F7OPmqc46WHa9p8dB3LVjTm
VbR0gxO9+/y4uwd5rvFpanHPOtda38o7sOOehGdfmzB11NuQSEFRJse4XhQ9d6W0
VfsYFb6GSnQvJWKYRj1m4ZUTxK+R6Poz16a2exqvogqqUtnLdC9Uc43GSz2mNvVO
pCbcUElHruqkcXGVARa92ghOh8vvzgtWmUhnE/5RYrR/ONXIcm6WEdgsHHHj91dc
Z+JetiVIENV4ZNTwkACppQHFtxR1UnbaHcra/TG8NrTEsSAt/85CnGWt6T65qZIr
N/AHibIW6A8lFYGKRnvOtoI7m4WOPOKch/zoP4ZbkRisshUjf2wAveU9o5ypPVzN
aazpR4uCyBT2jS4Vt7ZGr/tx5ZCob4ZR5W9AvJG+BnOWjee+7lFbgb7FUxSM0/2O
8M50hQKbWJ8FoPLFPZ339LX7sMG6pDro9QJeo8AD5MQwfdHAJKaulhkxtcRZ4/lo
ILIbb5MQjj7TBmI8ileWNPyUGhQKbbpaavUq2XN4CQrR3jXnWcFSfXuEmvNp4TyD
pEN+yR6iLdJYRzNFt9SQedm5yPdYsvVvTOS/ZyZmRnE7Zv4XXA93x9p7r2OlaZ+e
lL296VzVauzUnzV3ZKXQn8ISfw+/FUBxac5VLSJzocN2FaA3M2p6Y4WpswuG3Fp0
cQ51pzUD1J9fx7z5OBtamBDkG9x0lb1kdxLB17tmC0Ks+L2vj/byRHtxlv3KTo6j
GU5vxn/OqzFlAdgoCdBFzzTCmoTvkrAnCKxVAuipo0DIQeGSmTJKVTHlynafYURP
luOAQFnwvaHM4LBMZAE/euA//sgUNLA9jORS+FH88BygHLhCa6A3FlzLEzGE5k2j
ASEYd//MBU7B5j9GIteH306SlOIJzZq4sYaK2JJDd/vjnWEdAx1UGKBwG+FGYlxT
+eSaOGWTKwtLdiCGlRoPuVcPg9+eY2lRwB1rTnhNCHrlhTo2i93LWtC+T6aQpGAC
nfRM44q7PEBngErAlY4Qzqu+pn6JKeCah0+WCb51F0BQi966S9VksCowbXqvc1Ju
rqF7ohYSZwwMpQoJXJvhCWToemx1w9YVsXN2DaVP9q1ZKJ5pmEeY5jhfoI1wW58C
MPvub2RN9ppCORcIctsH5rSIdapU5/gEY7IplvTye6p+tH1fBP2Fjl9O/g7jDfSN
PsxMZ0YMLKVH89rxCcju6Zc3UUmKa57OY3EuagV1zkUpgbL4poks1Tx3L4W7w+g7
vUUnNWkmpfOvXSIXRxT9nMgbEIH6o4w5RnZQFggZFiM2DLBD29s/dOjtNc2/ekXr
zEhnmsQ8vilO7DAGaNuOD3VnC5E8W4L4LcPsAv7lK6IQWGuHHSNSfoLJAckKgc1I
eDIeJ7wzQGWP2rPf3NDI/vo6+MjGMq46hoWZ2i+DYpNIi3RIZqJJDS0h0Cfrc2uM
UCrqSmTf3MQ8XVrBesySRNdi4pDKVMrcbM1LQMtcRDkLwFMHgvLZHFnQLNDGoz6q
iu/LSPkfnPGuF00pVV2ICMAMXb2QXYkYOgdDHSW/gNc/XpIfi/0+BPXFFFalFkBZ
aLlJ0BRayWZ8Nq8upnGo3eUNVPvP5jTl7jKxfhHTAl86/tAluEiTB9u2CV3aWXSO
IJ7PJJFRSkj2nUp6afOOrGTB/cYOAAW/u8dNN18YAQuTpubtSmC5MW4CsNTOOwQ7
cpXC3pRK37xa5ca4yERALMT0bWha47AaPBBldgwivnqzR3yV50oS3nXB04gKjXbp
6iatXepqhaCr1EmfDvnTb5FFA5hWLzN31LL8p+FKBjfHuU60Eb9x3O2QEX9E3w1f
xrREpPX9BgbffZ3LPDaz67VKofyalZS8UlXIgcwqJMgNO7R9noWdsl2JWUSKGJIY
JFyOx0mnaA1OmNtRLwaR+EExmwL8asRL2cL4nLatE+P5LyAF4tT8l4R7oXta1VtS
b9QzS0cJYtl5RiXCreMyMJJnRHWRiWlmZBJCCjqxTyYI72wmr0C3OrBQgCu0KmyH
IxkHdKRdrC+J5w7Pr8ctbpxIRrCtgyUFvssSSDL5QK79mw7NI4pJV1Ko3iU64tpQ
9TVHc9fedQo3ZhuvICvL3hkLivkTJQoDd8SA0CMWFIn6HIXgFnqNwjwYd9h23MuG
uUZ5NzwoEUC+sYsHXhGYXvlxETJPNbnrVH39mZsUF+o16/dtvxwMm4Ri19HrP5Xa
OXa8RZ0Spe3SJGR/IxiI0/pMCWQIgiIwuqKjpFC9TznZnItHeOmpjRYr9/PvbZEN
yoaE9OJCLW0nTiyiWidfUazSL2JFQG7RYZNS5pPtTRVvXj7UJZ6X8l0rl+H7+i1E
U50UplWBETM4TX3spEPCuG7+CsoGJtZaX7cREUPBnxiPPYnHXjLAqyV/WHKKmOZI
71vxeExxuInf9DhL6v/gGdQfhOnT9qorzWyawcW9Bc8nZPcF6lZOWUSzuRvipYIv
DOsqyn2YeZGkBhWQlBVY6gJ1oBXb7Lls6Ff8MuSc+V3K6gIfaqhJO/ZCy7pa4zT6
Cf4bARCns0Nxz0ysxBRxkUiNHsGHmxw9F8j74uSnxOoQRSRzl0TWsi4KVOnKHT3u
R7taQpej6U9p53LVgTH1KgQ1b2CShTOgpxyByeHT7L8P/zgy5J2Qt9IZKy7AIBoY
KOk7KIO9a2Tis+FoxoVQJR4tl9zZj2Ru5JBRholZljZhRjHSHvCn0q0EHAyCz3Jc
NQhaNqfwAsmhxP0MdvbfJ2QQUyPAWqxUBkkUPyPCIeHtDkSWVkvwkX/mEaBAQo9/
O5sR8Jg4m8ikN/ITMwio2BhhVp1ajR8+ucyb6FBt3d84oOyNaDQRRTPkfDSLKAHi
9ThN/NA4PWJRSMo+Hb1BuXOqOa1jBepfZ82y3yCIydVI07eYm4KUI7uAMMj4MFG+
DDBm459t3Zew6WY1Zz/qFp6Q0Lv6FqLkNXnAs7M+ZuKJYMgwBlx7WMCR3UNmjzPS
/9pHwi0JMvqR3I8z8/6gadt5efMWfWRDuyuA2FUiH5xeLFijrt9bLQTNO8o1CovI
TqeYxT2agFXyWWYhmI5xKRzLIebGjvWls4MeVI0LFPVL2FQOXfJKCIG63tymz8ci
O4Zp1Z38O6DH7V6IncpbDVN149gxKfuiJc+EZ12yrKaPYwWG9YjAMHKuV2k5ngVP
m6syB6ibEMBhMsVFu0EEF93XHcfMH/IisztuRmgvYWXh/77k2kbvtomOL6MsFUCy
YO0liIQhO+zpsu33w/ItrAYIBtD8HbvZkImwT4/gZjKCpqfi7uOuX8Bxeyf6r0zV
e9wZOHdyt5KIEkw2AUcpgDAn6QqW2EJhOkHyL/CFQUz1ErTNY6jqb1m01DgvjZm8
qWtjDt+KMci5aNspCv7Rf6LwpvBhgCGyPThOuhxDqFveSyJsXJx/qFPKHThO2bUY
gC2Fjw/xOB4ylzgd33FEXIG4Pvxi8+eQbzgSiyFEUHyldljlOIhrLkpKQ26572Of
xXd8iMZPh9dSsrhoCD84cz6MwI39dOiRvl1jG9oAy/Uyzcs3aq501qYTHkoosZ3V
/+7CTLa1TAhosfkDjV14qHWYmFI+/S67L+L+0j2Ul8q0+QvJu0RqcOdkzBSjvzWm
NNpU3gcvVPIYT+XevPiNz35LCatea0+TYyuPPjgQWjaM6zTJwvesERfpXIawUKI0
8xms2mqixCQdpMdzdVuLvbWOUw3hekNCE//2b3JT0bHSv27E4ZeFbpGCm4BUigpW
4rshP+FBgSUYTa3KlhakXoUPabWoXNEiOoOltbbahKtcFXuoMWsLb21ebairJc22
qKBxrYMeRS4H6Wt29eWlORhs1Bpuyh2L4nPjvC9ttm5oujJrQz8um1SHzc5fgvG4
tXjz48aQ0Gbr6PAWHWjg6/J5aWNUIMKwUW7WARhB/5MTVCSdLQb3Swfl2qKOMSrv
iwVTFeWYGaM+adiKWuJ2Nbi1CE1obPQYJDBbvub8J/ZUMMzp8UkhZfQla37NTSKv
zAW9WPI3cRjMcn+HVbZJ4cURCmZw2Bxn7TJ6myG5GOoVFK4vFEgJNbpUYDES1u7W
kelAqJxpyhx/uNml8Y+equ5jJlLyaFZ6SwV0vgX3rFnDzW/GBeUOCZxMPvOueL39
Qdeaq7p71Gn1rbQBNIqAaXJU4Whnw4MMbBZ74jdsjfETy/I+b6AcWpdI9h6jbuRw
PVRvnqIOY91enIqLA3flVpy+EJbkIflmeJTR1qXskun5Rn1+VXf/J4+PApsWuYKc
eIbFd+WlymCV1i9FRZBkgwpLmyot17+RWb5kOrJb3IK0FJ7IRW1qXgK/zA+Q3OHY
12wQfpenEade6Ae34x9Qp0D4OMB7+FCRt2wYPhZPYH+mPPjEMwQdYQDZJqEr5IbR
p66NN4sc/qhQV0Oy8qrnvbrVUCMnCrXCPsTij1/kPO1pvUBUCddXUHDsG3IuuiUK
xTHqt3Fjt+vkwXYkRlC34ZdlNi+tItHW1w1ATFV5h+b2lJkIniYpvS5jBYO3OBzJ
E0YoX+rrYXBdpiZpmNbDVA9Q6eeiYElb9uSRLMcdLgQ52iMOBKe4xn75xo/1s43q
c46FuuhxBxUPR68mNEg8/NCVtonLZuEKf5kuCcutfu54DiG0qdnyH0veSmGgJC2g
HonigcNCJu8aH+CrpURV0Dl1l07KMnt+XcMomiddeIBrv9kDKUfEigU3x9kELEsp
z0Kv/82ine3I8TGdY7yeKDODsjkHk+dLsThzOuv6igZ2RwY7N8NGIA6uBJz+7yfm
DcgvSd3/AUlSff0glvtP3WSwXWQAGj3k9KZXBdZ6WXVsfLokPo2OwiSkZEkifU8H
zq2sS8PlqEIZLz8xW6t0TTLduictgekxFBmf9Wb3woHVEOz6TCteKHVNIIyNt1rV
Y19p9FXihC743nj+dE67SmuFkhCkCrHcgFk2LG1E6/I4K9bIcxwOX4RZU0bBfP1f
JKZA+D04X8x+T4LZ6zdacRxp1NT1R8T9YWanpCxPqGO0RdoBsy2WU1pRu2I4Ucu1
xfF1gitYRoMiNm6MCs+llifvnoYAeReaGxE1LCuwespNxaqQZl2FGzwqymchblqu
goyzvIzoP65ekUP+ElXWFztILUZ8e4cW50LdG8qqAkLuTXxUu2OMTGSbHzQc2BjR
/IxSN1op+JIV2PhW3FyDL6dIQ/IuTJ2yJblibvA7MuKI0KBuij64657WISdTUX1e
t+/JMoEcdsXQdhNXHmFqPkoKOtU1oG9JiP6CFlpRv26iE6UdcN6yegq6vBROqT1A
uOUNaX+IZ/V/0lMOVw4NnnRS7+1f3u5j9BpeuwS/4o+zOUz+XBwTiCNJdhda69VO
GqhwiXvuyPtYIKwfoKjdkMA97kZv0nXAekFnvaANKoLfdBcKlCUKVZriDX/6sotN
ICnsuIPOT36Z57vFCSXjuM9uHWebX8ASPuKF7THP5qHlXTPE5Mv7qa8YOgwbcEG9
BHip5gKo6TQGhvsJffd+EydRvyRTFsMlUof25UAu+sK+s0PE7ts6ldXpyA2640R/
AXYKsjkgsgigHeoqfoWIRGNQURHKmQk8XF+1Sf8Q7vjsrkCs/2HEBK+btRHnTBlA
lEzuMov0o71+LCrsdIA9TnxocKEKGRyvrpL/cI4C1D+zADtPq6sV1TyBjGK/ksP7
5uODvD/WXEQxE9X6tdVmqUsb+SWpi3dVfGAUeRzlCQ2zqw5gI41i+BaXgcywRE/g
dEU36q0Mf+DnxRnKZzZxZ+2lMinfpKvThrzNhzzSeRwKDoOPNYGKPQ3EMlj1rbtr
Omj3i/rYzGZov8eDiLbsWR3fDnY5IKNb2YmRDVhwAqEp0J/7SpE+De25iC0LcJIn
pEmA1ij6RbuK0/r3QtEd+2xCusAxvqEakp8KkeY7fQQiQfyHzkgzh0RtMQMl0VL1
thgNCaqYwWuT0FgH/PCoTcdF+nKk5sHsK9FipvZht4Forf/iM/9fR7OV6yyksYLA
guEwE6dSiwL4YBs7G3csn4wX58rbjzBTgGkEqR7afz70nRY5sX8a/lZ3UW103iF1
hiCoesnjHJ8Ms61kpKortIMa7xX+oIub6biKRAQmaBFQIx8GieUShY0EHLp/kasS
G84+ZraHrKsB5OOi+ofk61sLnf9RIDk459eaq8UhEpryISBYPn8exERZj/MFY4Pn
484QZhs1J30lxXUAfEFyf5DmQ3YAJoKbGIXg5Fq4RuKbTqjZCJkwGmrJD+EnRrsm
ciercdivYj1R2XsgCbrl4vdAZ/tdGdPPBVIPb1ZDYorcjFrFzB3KQCuQZ6H9PWfh
6v6prxTcyq1OBYdDCsd8zvDuw+/rsIgyk+XkBVZEi4E4tawQ8a9fwTg29kJlnL1U
7/XVJX3huau434b/Bdap4ofnjfQPKEL8AxQunAcmtSRZ852ixxqAcMX+txJMvYh7
6itaPwdUbAv4TudccDarldElPVkujnpVh3l3WLGnrnPAqSIPIMeJRkit0wOnE4Vc
kfMizXzkbuByIHKd8BM4HNWWZ4PxdMRq1Ep6U4ECpJuKlNBUEj4KqoWo2FoBpqdf
fE3RMr2gZPDRFa3GXhG/wLk8vfPpl+ZaZS7Csn9YyVQhZTeYKrffRtS/h7qs6FTX
fz+yzVoSrIoN9Bx/ALULf9ES/EO46KaQnrTAdrE2Ph7XwfJ/LloSgPhuyB8CLHwZ
/pqGcEgHGkOmCeN+lFOqNQPioMbR2fK8Q45QaQgmKsSPx4o3Q/Tv+cQS9SM7tFRY
pLX9Vp4Q2VfO2HCpTDnqpRkit9IsUwBB7LGAXjQce7/Fb4kmFLbjE9Tn6IoVZ49h
TkfFJr3o7VibQJdqzAfk3WGtF84u4VPdgk8xs5Xjbq6EaqG2Ddw6EguR6l1YmdSY
znbXS8xqh6rnzxPzb9JrYcLXKifxTffjsGybQTbEQ76V6jQZ7mBANPzRGEPxxA8g
FxOXTHNNEd994R0M0Igkx39nXVIsZV0j9YkAipVRMSJKCmGwNCCgc3P/V+LQTIpC
M4CN6jDzxee118McSRX2Mk2r8K3BLJmTsB6BluOpRO5lCXG9xuf0cDWsNnImjJqL
rx/FsyJPT/5R48d+vx1dYI7BCq0rH4HZS349Oaqn21SOFLpkeQFXWtkeCyaNXAWm
nmse0Zxuf3/wME+UeFJINbiB8l82YWlTkJ8t1LGhEan3XjI6CPvErc/yi9TTFYWM
I7GbzYMiRRMvAFMIiTWfrkqbgLW+/lOYSo6Q5NlJL6lGB6gYmT/0yqIJ6SyvxQjZ
qTB6JwvinkxkekEY/AZNCp29u7C5xS4rt8eb84+BrWWGz0dbBYBa9ZVLcwDf+qLQ
mQ0MxBlIm5AfAxXm9N0JX8o1igyDEtqgfJa9+Pr4spD4sXUuXW3I8Zm9NmCOFkao
WDeTT6nwLnnnsIzqEvH39uERS7yebcARyUcIqjuM4WHbxH6qo/n3UmDm91rH5rQo
UwKAL/FcHhSWwT1rZjjbMbMZQyqdVvpWsd8NHJkklc+FDcjH4sn0w2KcVlLkpyRG
fLEsaURAMG2mS9zBm0x9gJxty92sXSmTB8p1dov/jGKE220eVHx14AHWwJvA1uwe
1qa2yvFrLqehtL/WVUHQH8jX6wMx8C8UDEWTF7V6zNhDudOUZqH4nnXJ+3lLDp3M
E8HUtfzEO+/1R05z/KJ2uPsKsmIkVI7Vyc2aGSIaY4J35WS7/doI8uz08fWGaN2r
qPseo0R0Nd6iq3tsSyOoakplZi1X9nouXCSh/3K0DpGiWccePDrSrvYdHtTeV4gK
kYA1k/ZQ+fV1d/fbsjupuCKMoM7C/WGiaRgVGpXiv1XRVl6sLxYDCMt56+X1fxDE
9cG7rehYw5wu0PN6NmT2kGLeBu1anuYxDXieZEn7FBfKrX0Rsnxi2EPnKcLwIvm6
MAr5P8KF4ksGlSblRaHDHf23TmLv29VxEnGq9PzLuhST+QWyxp8L4712ufjtzL4j
ebLA+MxHpBmtCUQZNtvv4yJzRMieX5QBJHaVZ0WwfWao8QJ64bP8uB4iiCUsNUnB
Ub+dYwAtogDCiTI+aoy33l0Gu/GmYGBwBKSdoGzjQxUFyG7Loq1WZ83Bv346uc1W
QUZy9VWHDyyZymQybUxBwlu8il5z/yLEa16ixFOGJe/7SY3BQGmch56JMsYRTRmp
nkUte+f+7XLg9NLe67shKh7s4R8Id+og1XBi10NXPiM6tWL+MSaUvzWzursE2dYK
q6osIX+pBhzYLniLWiGCUmbpAerYm+514GnYE/DmBUWmHtocnN1Ftoo8UlB5jNZh
0Y+LGGTcyl8fPJFsjNMEh/sVXzCzqcdGJ1g0CRqeZCHwei/Crkz45v90NewFZ532
6DtJPbsn/IhWmKmqrcYl0TQD+pJasgto5BvTRrtenZ+WWAiMmEZew/Ora02riLvo
aU8MhpRYVPLapn8QH9lDEX3Glm6py1GRnVzjOAuNZjnB6CEFbRgECVxE/KKcTQAc
/K5Ctq8kzutfECk6WCPIcgMQZfjMjLe0PIxdEcIixN8LJzAfeNHJjwIqnay2anLA
L+NrG6mzqtgbsNv3FYb6ltiugAtJBVOFaZg+PHFjqHppZv4Rv1LcY/7c2kKvtB3o
cYWvxNSLEb0k++VVFYDEP1qeQd8OEsDJeTS5355Foqy7yTOK4+X/LkHpu7CildC0
1zdx5jB9vg0lzQ9MkCdQPUaN4s3VxHkprCT7NPG+StWDZtPm7h2sPQoxx6QJOKW9
+I5z8TIncgFZA4lzBjHwsPHcy4GtenvFvtgzXVX4TH/zfZiDyUylieQ/y+MShZKV
lpSF6EJFWkKaI4scFZlz+pIS/KhgaF7bkLY2eBGaVnnergyZwy3shl5mD4QS4+f6
5LqbXefzvo/221JqtYlrdVUbTz56jlgI9p/JHEDkWHIGKIp+I+RymWoK8CRnR+Ej
U33dm4elXmUbB5dGoy0mHS1NOTeum+5NWFzQMn6tYqYgPgDGyECcgjeB7tQSfpk0
Zfyq/epo4bYJp4otPspcClDflNZpsBxZt62CiWKeyUwcsVlkS4RjHxBlfqMwT7Dx
AbCuKYFZSJ81OMNH9JuWbV8WrrttZeDg+SYYDM5UIGfMlY2+6s7uCBHRSIDzH2TJ
om5OIUdTOxTwh5Pv6/YLF86xY75Bf8+WdZmc73VVcjGEkHkpt0GsfJ6DkjoSO+/b
6idXontMisruJr0daQzpss8BB/a6RxBayLrZS6JuEFjgUmFkyrSOkiikTgq9cE7/
oIve4R1g+oFedpGdzESNtE2yBmuGdXUe7axXLocPThIwZnygj3pnlTSxl7tJ1+NX
nuS67nVhj8h8BPby3Euaua+FihoruFrsYwrXwewNqxKwDrgdmaN7cC3VJFsghZRn
pYQUAi4Y8n3lEHX+4WcQ32ljIJfB7ZlX1w7c8LxPFnXa1SIhZ+qrUsWTwv3dOY/h
008zBeVdfzCwokMq0yjA6QrlAa3pLW++qi4tcBMUjWqS22bPPQLoIL5NOhlGn7gA
Mlax04HRxs4cVU3wvZ7cD73TJCb35aAZ1pQHTGZuLBTST7AgBraTaVE5Kovo0Rcd
TyVoi5vsevV8tviJLI14phhs0cMA42vaJKtlP0/zrVydMdDCHUXOMxvqhLLz4Wke
aBegWdeVZ8NGI59REtBSR28BqcyllCtY5itXmJ44ToAB2okQPbGAPqTHo9FTxcJF
J2szjGdcl4unSoYHykHcjXmivqbZGCXAsrZ7Jx6BKj4mmDBn+OEgbjoq/gVvRhNt
oZ64zutfc9ZzuAn7ELVhomDWOUxR+wA+v5r4m6l+UeEHPcaJx0eFFsQJHL+iSFCH
EFqBRqtAIeUYBwTMnIJ1yO2ynmsmACAG/sucKmTLzcfO64Y1LjfxHOnoAKtIuQrv
2uejqiz6kGFvYTJO4kM1QP3TuZwmHuwubarKrq6p5Js3L76i09Vqyi7RuM75q3+/
lgtKqZKRj190FNowVSxLPYGKlsbsVefv8o94IF1PjCBG871uFgJxMW7y3qT4+XVA
haYwcMMyN0myibwpG3eYYX2hIcQ329vPw66SUJVzugN9rj5xsVSXOzUmiRpyidC3
zAiIrpCY24Av6wr/chOUZpxKbt8zfn5/xdEh3fJtjovnvBjM1c/LcbcRIbOYtB7Y
XkdYFAHtfEATpZZ2O+802de3Uk+YiUs56tg9wZmiBJU8a63iNy6XzvQV/buKtv1l
3Po+SrLj+Zb5m2hQo8olbfU3je7wCZpn2sqOoRoFy+sUnKj/droPLVinRESSvP9M
zq29lTdTT57+QZRd/ot/uMUkHnteexVLKQgASfc8sbUyntocfbNWblup6PZM959Z
NjUNvWa+sigKlklnHCWxJ3Iepr5fQyp5oHfqAMM/J8u1WcPt3vrBEwA5SiOGQ6Bc
1b94L7AhdbcVoaOp1KYfOvkYArzQ90AczjkKeHZ0USky3QQXYXj96FCnAN34fWqg
iwApRP2k2J4Feq1i5jkptRZoCGN/fkZ3yvrGfRP8WuFjgc2NIUi6CRNnRlK6RHxR
R15LfKRFgcBeM2zferqYjOZpnLUFMewEMLQGTIU0gGwnsff+RLcMTTQ/bKT/RuWe
14AtiNfeNvqTOJf8n7KwwQKrhADuVz/zxgR53Sov+QeMeVc5h6vvsknEzP74A93C
9PAK5eXqxTakpaqXVBjC7HxjGKpTszJRuUxB7XmtT9kx6Zd/jLubX6mB3NkW0tS6
yimG1BSs4wMBO/PnvgtrJitAJHoTjrwsGgGu9Lojm+AIuN4p4IZ6wsFLUNuByLfG
D9l4aMdKDHzLi6adoWLEiwAr6G3i3YMln3iIFJ2DWCE01vVvGacA8OofNqPYJIRe
omeML1krY8FwwH4xuiPwUTcxNe0TNqHx03iwy9IXUwG9ZQEcSxaSJ24DADMEK4wV
Vf8q7Q6R7CmvC40BxeslWe4jc4fyDSfUysXfW/brhuFz63U0JjtIfnIYJarwy5hv
kCYyd1b5VWN83g/kHETieQm7TZwXgCiDxr+Y4qPiXikqOzAfaUq5lZraPqCdKvjI
wQGBE5+XScvxPaxA8OPgsQKz69NUAfS66tMfSEdkonwDxGnpS61nELXX0QVIj32C
l438HCZGpHNYqESVpo8DHos+QNgZ74clESUj1cv9dmjz5nWmWqPWWq7UNV8Q2azi
kwcuEPrgaaNRNqrOcIywAEELIYtjS5s1W2G8jWWcgsTSwEQ+GrZJ0giBhz6JSftB
lN/HiaL7YuZ8pMzgR1+IjMytGH3DUrVO2izB8RiNBvuPEtbMy0H5MmimPRhgWjMQ
YfmYOmr80XB/JNmbNEQfSoNV7NraQ1wAositXGWYHeueoFndP9LoDJLKfs8RdErm
akgsP++QvcGgV6K4P7/tN9mqplifn+29TG3NSm/ICpz55rlIK9fh86GOs9b1rU6W
9sT+kEFVQRp+hdzaEYJ1j6BlJupfuS2sLWzdMDoCCbD8gmUPnErvvG4r4mmGJCZh
q5bQhuYAQ+w621wa2PiwXEksvNpOyD73OyABhlxECE/lWTGafOqTcgjFKfs5lr55
tjcLinpapiEl4Fn0HNPfBCiZ7SUqDFVKRINR23KkNpLyQagVs+NhFp7OLoymlVI3
9WDnaRwV/A3raCZxk3aojzWlqeNniua9fdpx1QUpKgRoG1PUZW8mgZY/IbO8l+DI
2Z3hqNHkSezedGTwO46I6oDRoxjxo4jNrNTiico27uGuuZAdcypkT6p9bVShxeKF
Wr47TZww8lvuzR07Q8FvfHmLTBFe1vyJB0VE1bPGCD0YpXbvNuM9khnxuRg8Ikk9
tz1SVo7xjk76f0IBNMWSkteN60/oMLmqG8L21HoMImnQDWaoQDYAt/4HlDtUVH/3
dCkz+64eryQ+h+qlUuUJsnLZXpyRAmDyYjmAl1gjqn9ebjMHDyCAKvppdk8TwEmQ
P7zCtStxDS/9h0kLtH7wG3yz7TmthX1nTDq77HIpMxo4x9LpDgzWCd+sw44lXHKh
ss+s7Ne4QxlLbE2XxKYQEduvfLvbg7gWE7O8B4hIEYXgkBMeFtxCMVJyuFKr/WBP
2G73sAXKpCG55h4w515y/K1p4hDxuanfzRtO9i5HwGaFUO4pglLv/4Sb6KC245zL
HpMhYhaEL8XoiT7SbuwkG1w4bqOEmpm32boq7EmFhq4+je/+kl7tXekQ1rEB6FlE
xhWBWTJWWGnd7gwVIEBjRkA/QDDGAfKHBEmXUtqiE0+Hnubwyv4GflEsydNKMdiQ
e+Ejg97PCpHtG6KejmK1zkSBLsLtQolsuC0/Y+OzAM2le3AVsoaf7gmD37RhUaHw
ZUb5SsnsPzPEe/w86XwsQXkvauI96kKDxzRun01UwpCG6wGobj0vCVmSuGiT+HQX
fqqCrZVI0D92ypFdvPnTMh6phJ6FnTCxWQYfzf+yr1Lel4gbYsaZt/vaQSewxWPM
ybewL7i52ooH0quyHBor33rSKGog3TPO0sXL9EJnp4wiUa5e0u4Zt+nI07fSFhbJ
XxTXZHuO2jkY8akOakg9HkzwxIuxtfsSxQOPsd3gDNltTnQP2VxuJZDO/eHbzhxY
UvU3TsjdR/a8Hk7UIPqNpEYHdMmS1xV7CvBgyCbt8+kcPBEQzsLvx9rhvTGI/3rN
f+pPYSLFCddIa+ZRNr/WAJct4nw9Xo5GBcl56yJFePZF0Dp/+mgjgh1ik80dxNCy
ReqdCZJ4+TUmP3Ml1o/j8JOhasvuDLeu+0fSlEjorI5ZGzINqsDwH3xICa0Qhr6a
IVV+gIEdScIjWGv3VnMnKFfXMEXnxjaATuuZvRmnROTIpsJJ6DV+8qXKpnl42n4S
ex/JlFmG3ikSYk+qD7Npedxil4etwk3WFca8rn2KT/5ilbq6ULQs2MBHO/WmrDE0
+ANOxIz42LeDkyNt7j7G1f27Gx75hzrUMU3CMlreJwP2Q/bTOXv0IMXRGTJezdpR
30DjlnlU9jyfXNzvpwSfs2g7IoGFOQutCaEN/waxlryRA/Vec++ELzMTzKxaoWFb
O1GLzsm2nLWHpHq+x5ECr4ca0Ew+vlCBsGiiTJ3JbXEP3VGki3kMsks3CJyUrGPx
mlox4/nrUNHVfe+W63H2yru2MIkQZCm2MKm6GdW75Pes+MWY0Gs8kuvuTa1EwKd3
kQPW0w2oLxtlVlCcmn1Ejhk6pBzM+C6LhsPwgmdKsI0QRBymLMP0G+H++2J8fnov
C9LzUM54HgmCBmEoiCnbTuX8bR1wR7f2W38bjNTgrcxOgNI5hk34RQ/qseENrVoM
E6MpVR/diCwPx3pkHRqOTPb3PEa50zRe20e5mIBx5ataMyFLicJzNqU9q8EXYjv8
xq7HzKwBPsPoHgEhpN7IDEF+cf7rKW1YORGHmkmQffzBIwJT9V7nkfMVZVlQiPoi
eUaN/Mt4QqJ0pXam5cWFvWn4DucmXBGdQyJsZaPMiLDZJqxEUj499jQtxevtm/KL
YHYN6ZF6ETNpNzHKu2Fji0sHy1Y1jzCmJJHYPlRTmvWKUjpT+jh4oGeMXJfZ9MNa
FUMDlM2eVn2JcfTwPffo7LSFm/ImvGSWhJEN+8vkRjXa6T7xCqq84UeKu4ki1uuv
FGKa3qr1WU/S6JK+wkbb2bU3luPSa40xZsP1MEJb9/vUsSSxF6ghBFALe/5izU0P
jCybGI+KJ53jQUa5TuFiseQRUMTLckunGRYAGYFq5FUQbtDb/g3eHGhSpEzGfm2j
up169o6ANAo8TJAr7sK4drWycwObBiZOjX8kBmC423i3wZF/cRMdRHT48R1pX7Ww
6FSxgWe8o7+TC3M3rt9YORRHwJ5w+ALVpAmaxaGy8A5lG2w7hWWHzd58oSyid59B
vbWgclO6RHy/Jc+jr5JRjRc57YHjhubhBoVvcmfZNG3flGfdO3iJzQLinn1SRKWU
P+eG2zLA/nSND9xovZuoAYqfjL5fRqK3GmDUQhyoa4IHAB1GXNfux3LPW3KSA9hR
nPiIKcdSnSFF6X1fNQRZJ+lIruzwWOr0+558O1NEeBTXVZP/5a5QXREBAw4+b2V6
2ss/Vq1UthdAH3JpWvh13+8M7bToBXcdCTb3jPv/iy5raeVODn9hbb1+LLW1XNj6
JwbvQWbjOZY7A3L/gf9cf3vd8oPlsf/QIWEJOUQWV9AgVvAWBASbdfDKYjbfl5dU
L5LV3cl4PaDnnHMwa2j0YTl+hXoKQmnztkziBTirmW99D4MR5/GUKTz6c3rMqV0J
hwPbQM/bIhKVUb8TXsUzSjYa6aMPKeRbwJ4PdHNey9ueUlmCoo6nXZLTVurhJ5gy
bG38811kFk39cuYuzFrnDchfXnGgvW2MZAkx2swSnPs5Hm1xbflMQjgtFKVYRRM7
qzPk14Vjv56LZhGKEh3or30rTpIXF8g/n5hc+1QowBOSAqBd/IEmOAbtn4WoZFox
50GzEwbeh0wSJT6IXDbbefuW3YRGx0yXSs9ritQyKP4Hfm9bWtqcIg5FdCv1EpUy
7CwgnbhcuymwSPoAxJ94wWyMiqm9H0zogCYjKFJaLZGYwkqdQjOZI2ZrSQmqlMQb
JN3cALYZDVq/hQs7B3eN9NmvUaZ1t04JOOa9DC+63/h+aYG6WeNdyPUlU8QBOJfO
q1rzURbWmW6sRsS0wBXOhGU/FwAcXuIGhWhiykG8DC13R86m9xGT0cKYqLif5Yto
wE3kwIPRh12ijDjvF9rT8hNPih6bh/HAjGNlZWvRs8aaRvr3wR/E99obxd6Fh6Ba
Rizx/j/oUB1g4heDUhUg/KNcAstzkw7sL609maccMsIfl/TixIz8J66jVEgrThLd
wEZ3NSDeOI5J6reWQ8eyiOzg4q5zzqqtX72xy4dr1GrRCzqIEaPzo8c38qEBJCQX
O9jd+QRje3iygX2bPgi5dBoTf6PmxLDQO13He1bkZrcwteDNilO3iG60v6oyjA3L
bB5tRGF1/+yvhUFHddMOyNZxZ5EfycYzPmP5Eayh73o4l5sC9HlWstOghKQx4zsu
t3+SA55OtT7QRb2edhWDKkjlxz4OzNIKURZ4GQ4GVwMCWX4qTTU7OgMpkTbHmKAw
hEZdQzegZKmEhEhB519UganveQ88dnGy+L2C0TTkUU/kExU2f1eeEQNceusbITZC
QM9xyqPgD0+yodRE2boVWf2t9u+lk0ryqEXjytMaxO3eQNaYDiWQE8xpVJKKEtLM
biHmLI3VlTHJcdA7aoI/wVoeYjjqKxtwmOrAsT6EQqsXIDmj4g9AStlJW0DCErZc
eqmP1jmPznmRXnVI+WOw7Z4RkQPnqMhCuuFlpFpOLo6oTqyg+6sXq0jQ7lko9mlt
srdXWpOdR/rziXj6dD18nDYql+HYjPP6yMbIEFmWAKA+gb6P0UsDkitUxhsMbsG7
qM6DQ1qp+aq9VuJ+C5MY66MujZk1ocOCPFVBqr+6/OAUyNKFML9/wiDBCPY9votE
PP/w+3d/Ej/4v1Vp/wf5yNMcR5jlBIlv1awj5tnPFlRAJA8+xqIKLm4/ycq5RJr4
TkQl1H4SNupATSYtmwYuaBPxo6aYr90JCXbyEXnwDj+RidCNnqs6MbcL42zh7tV6
j91nFD9RPIEQD5t/7/ZSxE4GiiEfhvidwg1USG1u1qty3eBD+QmCdCbQL+ezEWz5
L/88cbfGUucgooOVmdag1N637p1f7+3aCdjAF+L9IfXMjHRz5cuLtPTcimygdQvA
9tJnm//VdozgxSd0mllSCiDzRp5Z8anUEuHhdErd3FvysaFcZj30rq9eg9t4PB/O
8oUG9jcr9rMjGhbfQ4m8EnxQDRadF6V8CZ0ubliB5RtxoaOIgz+Be+2+Zl4hRLN+
gxb3UquIXoM1WfCHbKjctLzrg/WTGRbKQTmF3izXYi5IZDO5T4P04sJ/TdfCSXf8
4ZlmhDHEWDvt22WCs/9Edsb2UgzwAsrbTCTZj3dNOWsu4hj4zkA+D7Je6zz3Rji3
ZlcSGhNkn1tX0RniDjE1gM5BlG4szBLJE4qmzhOAnCxBht5hjfl+eip1PhgWXkhh
Syi1xpLhGyVPgHMXwoPWww0BKaqhJfcYEbA7Z5jxQHreGoLTjK1vontwUuQVbyTH
0jQbt6dGRrUfnzZ8SpCOFvFcU98MmDMaxkWq6XhXkCEomkOtOU7RBm2uAdD3xKXa
lY9Nse5503GmO0zeuBDY3ftTseeiv/xzegwIRtGbu1aDN1f0HYAzlFtI0xLU5eM6
XzOoA+v1Xf88MW3xgCVzp89d/MQyjxgY6FWHLX7koWy3tw9Tok04BjCZgnN+GSxp
H3ZaQWJXQxB5WnO0SgJSeOAPG5NCpAkw76PRNheR5fSXOyRwwbSv8TUTg6HZ9S79
rJhY2LKH4+BW/xFX2HWXnHGyjmELNr9Hctf5eOH1ntfG1wKHFG9H5GpJDXspOC9B
tMP/RY8F/SbfLOeeZ2eep+7vmeLcU/NYUEA0fCMgApSGbOLU9/twnvdtd3zqg7zm
z+8axJvXc/K1IQr3c262pQJ+PasnjYcOYN2GPQrdr6C4eggroXO41qUwTAXvgC4l
diQFmp10QVRj07g97BjvZApk0O9NOg5wz2Nfs4H0SQhhJe2u4kdXCJ+/NuptryKP
ijh5jPMFqshRKNSZZNCFSb+aw7kZP3hIfV5ButfroJ/emEcmtx6NKEaFNTuVM0OI
VCqlN+psDFM4IbC7JZ+mX5U55n6O+UziIgUs7GNCMrN0GrmtYbxil1PumdtmKulr
c2K3BB+2v2pbxdVWnJRWtpD5V4GM7T5Vu93KIGuhVw1iQhW4BeucmmP2Be7/iqm5
IM8KHkwcAolV2n6IjlDYEeHYDabBuW9xFF6w8owhJSa3EUMcUUOy4yhX7bhJdWM7
ABdT5hySqQZ9xmqs4bf7jpICw+JArd6DttXw9ypcD+EPuc74ilkD6k68qk2rKLmf
HhcUWRlZqsx2IzQuKcm0tgbpmL37GUzys6OgMmuVkCB1/CHZnwusKx45/G+4hl8A
NuQUQ84FaDV3rBi4jlFk6+1YmTlwG3H1Y52QptFxsLYWQeRncd5OgGjH5giTjjaY
9B/+chhQCPV9D2O9tQktQeQhMUzvUa8s0rl/vhiGh1jcAEiPnq2IueXpL2qdsUFT
eeR/PlGHc0oM8p5P6rMw0zztyyt4JwVuBD7YtMFlA0sufoVjYtJJKjD3kgW67unV
PYOyotmm9yPxnuPwly94hXnIhA+aPUFni6Y+1gBu7zAcvu30bf47tQL3uir7Jh9m
R6myMEIaUSM2RPGKiqKE8CvXZ6BZGBfOJGDiniwxzfkQkvdUrW6jh6EaMOaI7o2D
zy2Efhw9pZkd1CjXF3stHdTnRWKzudrbNF58SVNe+jp8Tfy9pBSn4RrfmHx5lEZR
limpBy5O4vUOIBuMbPdassl7R7+Orm0regHTf2bg4OJPEVniR2a8rG0TOlWiIfd4
2herBW2VxHk9PFHButpgXTA/FXt3b0F/zM+RxhOKUFF3ZW2q1lIws9UFHruTeJmd
egJdgPGwaMTvycH6AVAPWN8/fIuyMSeyV+U1twpk62qdT8fiIpetSgJRNvZdbyUm
wkTjyfO/0DrSwFRnAmCfHzkr/ybu6Hi0ND7Ya/O0XlpZsIiiScQBHZHvKqGrPfqo
26mFwPB+92iTjgWuzal2pau2MCUdhxKOAM1YETp1JhNJSgDAunqHCo5+NP6jDEYq
a91cGXMpVbRUQ/Ov+G1no9V5Er+HWDZ/FCdu75wB1noXa71cgmnvq/U+pRjAhKSJ
eBqzU9+2KgShH3mzcTc3ezU9XgMjpGHeawOU8UuVC5bW5mMQEA947m1PC7NhtAmN
kthm5muzzz/z9RcCf0i6KzxdkXecH732q1B7bIJnfczeX9wvq9AzXUq0PnsadBOV
D7Hf64Jwu6kK6QjIQwGlpSygxwbjjlmpSVBnvpB6dCwDhUctTzD9myXGo+afRodf
9JCdtx5uh5lj7K+rix2KqZDLPyX6kD1a9YOF9Fr6C4dF3vxXvp9nTQ+seLoEJ3dw
v+MLcZ0V5h9UvYvP60SOp63Yef8wIS6XYR2ppSOceyT65l1VLYGID/bewMGBxVBu
PgF045AV8ufovH3NGuI4eJzF09l73UNEeAAXMgTw53K0y2ARTZICXtslhZVVSQb1
0cHFqU5+8Zm9HPicegzInCZbPyi6LJlHjlKrdkHwVpSTFXaXDtgJOkKTkhpapPrV
NxqwR5zVbg5WFzc2tmo0gYL6i2CeKeEgzaYnwYYoNnwNjqe9VFuVmxF+Qiaf2wZy
uW+MJIcd2/08oGEo6GmZzZGcyytWODAZcmDDgxOCcybbFX93QX+UFIoZLbKMRjbU
qjuskDXvV671KmrPY2ycI6mKV5vWXjFCgaUhC3UXUhOS3T0IqWoAKVZE8t1UeHOI
pFtr9IqgZvf4eMNyt9Q0ekXtwyOeFxB1imjnkz8mDn/I4SbbDjD1vTGS145995Pd
XdWGJFaVg+S933mqT79hOnYLwcquzLpuFmnJwm/2ILQBtrB2Z5zdvGEmL/xLiSqU
rm23+uuPFF5uSL3OePAEto7NKWOFFE30Ll27R82DBfA6y555t+TeVS9alE6L3u0d
czu1KXaXg8ZrFIIFJZQoy1CvFIai8tFzC4d3Dz3zRrS4T6ysIat598Jqn+Zc5xEz
t1EtNO/r7onW1or0IGWHgkew12/XBZWipJkR4cQBKM6ECqbEHAPWvuGq4tqJGDwr
Bc3GVcl6YRbG932UaMcAoeEWfokalV35VvuHNS0qKpjhQU4/4rhfCj+VtGVOb6Hk
JyXtGCOOshv3f/ZHylhsV4g73YJ2C2tebCbNbtd2vWuMK+D5gfYaPHEJJsx2IMeE
ruVgE0foNNo2TdLcmn8hxUZ2ALHabOShjXkX55hg6IfaC/dJZA3yfuIeJnDqQRnn
Hf/BHjIFiyDrlg/pG5/8MIIPzYB7+bLJZlgrD07UZ+kU93MigrSaTzqlf3oTJKGH
BY2aRo06wv06KOZon2kjCRkwzWpOS3/3eJfevH+55wWFf4JB39tzFmLWEE4HgGlm
AwTDzD304Vn0k42rODWSn/NC0z44Ek7qTumphADCuSM02P7ID6Je8hEFKK1vDUPs
TyPU2luc5TYNEYZ6/FAlp8cd2dZ9Iyb9E63GQPr61Wg/ibBzZQe9p+ke6owJsd07
4pHvzdCh2/FvYqJ8AxQ1hnIZ74H/G7zFbxMg0zTjLiIg78evoopJbFGmf9mHptUZ
FvmYRl4YdIyOonayV2RDrOpGvKJtjOQXQPiJ02ZsEionF8DatKxHiG54N49GtSY2
+UVYIO00XQr8t5ytEXFx3yDa9IpmpcAl254skin0wffwOEspR9QOuvCwK0Kvqph6
jGVGWefD/SOk6ZA6Lm+5Znr9UxLMkqTJOa0RwM3xJPFm0uFUsjsebgyUnfjD7X+J
naBRwHlYg3/swMaheq8I7/bQOY289JsJSN/vrqaFeDRSTB8m3q0CsdAoq5+m1fOd
Buxb+FBkfKWv+qN41C/HqtyMoD5JGHjLju/u5hYkTFHdomCA5HaRasHkZ0SENtjA
cBxyP8mnHIdQ0F873AO9/lme8f5gdDJig6cXclBfZofNbUFBmGbYElzXzxJJq3Z5
O7n4o6FD5edWO8uoBwmrccUiB8EMj+oPWZDpzmmLkjiXkLvgm+4bwGyUsdNnhYGq
KjJqcUE0xVTMXYALkvRqcB9z1cKCCabKyFbITf+e2TB6U03xU/TEihrAralyq58z
ROZhQ5Zia23CyYbmWd79cmRaeUnL5bMKJELmCrKFuZH5+TndhlhD5zAHmdwa+q53
0sLCSKxRD6xkjMJRW+iCWPrix1udTiKcMpPRHqjJsa0cxV+69Qpa8d/TNCbAajkE
1P9qdK0GASkKJtxmI8Q+f18DhYOIACrC7L3pVviisV0Yg0gSEzANZdtcqFFImrrQ
qNWPNSsaIolOW2uF6J27ukN0+a1MOvXV9rDa/tTREe/CikPWIx/koS9do3PNyeiq
ziTgRO0WevA01sb1ZU8R2PXv2rN2tcwPFn0rW9tealqe0rD8+pyKKPNrsZg4BcE6
yfkGdcA8QROsw9fwQCNMS2ijeb7erDQ8OsFEyhHRNMrtbVG0+Oe+3NnejS62s/W6
qIq0UHP37BE06MsUmuNqsfpMPqnZbwJnOs2mvB7l3iy5LNMoLKZAFt9tT6bswbQ/
hHDUkEDoibFFncBIazX56idYoVryZCpllZzU9hQInBOTi1ib9OKhEI+zI1a/f5/b
Jz4faj63yfL6/5xzIv31vX1de+fEhFUSnBGBsL8p1jhhglrlz+o7WjSZOWNJD6fS
w6SFPriamK2ehnNlSKvw31RvU2heAN/A/RDjMfMbhnWxsfplPceEdmP+JjI7cKhr
m0QXTrXwxZYN7VZYcwGN6ZY7/Yr74dqWlB7G7+tJMtDrtp8jfIbAdTeYRRSPLQ2C
BIRveUzqQML+BOo7sTv6/Q7PCw0Bf56lgHlBODgfFExTPzi346iDby89bAm8xJZW
Dc3yJQVjfekmaMvw/GpoVpElGPsFOrqjxc1CM8YVCF6QoO+hW7HpEAnac2HQ7NjV
L6M8TU65qsOqE7oI9nAQMt6Efj42PH0SzBAfKaXicWJK/ff10MsZ9b7FlMC38dd6
XuvMce82ldP6O2uLacXG3kU6zDep52c9m3htKjTuiJ9QlA+Z9P2Dq19RLrQ/wXc1
UqxTBCi7SuyT+4rEygq5zTIboCPwx5UseEDh9nXgrdjCg1HL99Vn04+ckXb4dIgY
QsZOWK82RQ8lRDg2ou+c9Qc0ukpTtMLpxbqxq3rcNfiaz674p7l1ko8mHZcGQhcK
oHsV5o1JpE0BhzFfbKGlSqzB/sVixOUlvX59Bgru11wwnPnDvpUqlrAwqGdT6Mc7
A7G0iSOPvsUKlCU5h1wcA/UjOgaVqj1j1YTAGh/uTIUvRgLn6zQIzKxgDlL3lhz9
tvLLJi0POd2KsEVmcg1gRpLVn3xtUXR1eTFb72vMpk/huRHkpb5j88eLMFWpXsQR
BSd+m1zo133SqYG5wK5rabah+OJV/LoVHeW3lOf1E1C00GiobO0NYl8zJf0jY/xV
pqd1o1SBhjsqXY8Bl6LT4L3SIcEwZy7uq7ytQDbPl+xdcqQvh1fTPRxcBoxJ1oU+
y7r7SCdcRZeOkI1rUCyQHghQlQ9dklWVbnz5W2T0hTCJP5vF3w/TjyGPEfhEZoiN
E6LTstUDe0TEkRiOR3ZoOut6pb2Zh10A7q3aLSl58eFZl5NFLsUBFkJRC1xrql78
6190evcMmSVYY2xHy4ehK84mDx313oUKmgkW1zaiMa6/dARJV2Z8kj8zxw+qR0lY
6KcKEuptKt/RpEq9IN8rJykNHmyTFoSL7R0maJIOmsYmEmw7dkPtGDU9FvoP4SyG
yDFQVQYnHOzAYg2m9liD+ZLDTvKhVoutxc3PMpfYIXRpKxty6cJ7O3IZs7a5B5eu
HwqhgWf4ipIofc0LnQqaWUGdiLzaDH0buSwefzLtUzhOizdmpsfh2wR1HL6BDc1I
hsjTbxUIqS2CPJ/XJz6C9UbVNLR6AaEzMn4pTrtIdyHidmIQtW6UTRW32ghFg2gm
7veiD9oiGqJsYfY7sRvLDItyWQinAgadaCxMGL6tF3skqVOatJZvH0N49WpFrpoX
V+LeWgYD0Qk6+PWEDJHjgrzI5q2ZQopL8jockxc3M0YRkRVL53SF7H+gjgW/rcCP
GQK6Ubx8h4mbzLYJS9+nhIvDaBKAZI8AKcCRpEPr1+AZDw1JXfrNOEIBRzdDcfAJ
c1+ZO8a03aj4Hwh5ZcZ5bkPIvF8ohIJJ7SnlkqJD7+Xo2sOWvU5POsUDc486xl0X
sNGozGT+HJlI36G3CJlqzEjiDvODsQj6LXWdvk5y99SuQruQHZEFboiJ5l77ng4L
wNhItEybplQPaFUmZzzu3cY2r1/UdP+VDdopQ1k1kWedQ4et4lSxV23imTscDKsJ
PDneRcHf5Pt77CpSisAmLMEgPQ3gAQ/vZbmSKRa3QsYCdUU6YGtrHCfR7zFTUXiz
6o2XxRtSK7g6aAdH4Br7SaTjr7mQ4ZcXrCYw4SXsDNcGJ0DRMJZ7Qv5HXY8NYPNk
6PrehqjW211C/8MMQldvonXS06eebI5cu+HzX7vTFhQDp/8E6Uwp/JAFxhg7jHR8
cL9C250lMKZ/mgGXjQCFM4KJTLEdUwtNbEQpNd5nhtovN1/XUYjI0aXGhvSc8us6
1qkTe3qzASjNMpP2Ml1l3M2Y8vpJlRKwy/URl0jUtBko/yclCjWr8UVOU/aQF8cv
AXHTWaPha1/ZDijwJtA0smpLMwM7SjhVSiz6VzwqV9dYSaPI//WqT8KJz07/HSMR
r3Ze23nPXWiin60y5bHVxmdFN4sAfoVxK7UVmjxhaJp//PVF8ViBmaaYxWz7vtJz
i93szfWwWO7LHJcZPDcdqlx/oxDrR241ZT6VRA0dTDD2Gnu2QZLfAwUmS27FvBMC
NypxHuEHwi0MaHRux6rnt8HNSEQzlK7HLgnJbkKG8jHXHD9gtyM8WpAX+UtgdOWg
68vqwrZa1kW5N5SE37duQlU09HN/6kUv4tRSB+tqqZszCv0ty7S2B0QnI+hiH0U0
lZgVFWh3+Btd0EyIHwTfJLDYXzJsPyrjHaOkCfdA7K8KkzXGFx1LdVdoZ549Rsso
vkK/hBzb9LM2ri8UvOCD8ulIBwN7+8EIfBS2nstbf4DNiL1VF6xTG1SKY6lJi71Z
9gq++gNInlpd2xSHadglBE5ijghh4kGVxvk4knXervhW+CJgP/ksjP2cTvjC8SOT
igJmslb5VavLc14coKFFHFrmDzPlWWm36F8KfXFU+sNT9yzHNj/wJN/eD9jh7s29
L4eOmH2tonViX/lVZXEjNTTwx5HA8MIcZ0pnTv8Jtpw2WldKnggYyvzhW2L4rY1A
UA9W8Wnp52XawEo6jCzusd4KCJ7BeU9b7L9bMsAVPYfQykRxj9roOc2qnGhcmET7
9vEsCNLGKVVTzyXcN9jox7w6r/fe1FBThk72qJOvHrVMuW1by9/pDq8aLBgEh9US
y4HQzsXVLkK8VsKiEOUBQrN4pJORuNHAK2KiAyoHiowbttF0vAFwXxj7PQ96K9ll
A1M8S7VOI0F0OK1xDrE1JZ0yZ/SoUqb3vnerUYfcNCqvFRHJXOVftpl0Q4kPHvS4
9CyUkffztqTTyfZfUqqAZLACMlwSSasmgj1MBucXstEbwUI76TKG9e4IdxgnN0x6
TqAtuaa91PWDlPQAZRYf6jTAvBz745zwtCm9i++c+YMOVv3NoXlsj6El5gsVnjrp
HXEe49gxiQ86YIcjihwtyvpNFOQgtw1ksBU8z2S0YkbQ/amy5DGFTgBiCX9nR/fX
CoiblnbSpYZXe/pDpu7iOTm5ZNlGVMBalDdb5+TV7WhO86mm3Hc850YxsCTpEyOU
PT46dAT5IAm6YQkr5YJmwB8jeoF5e6LRWsEHqsky9d8y/2aSQneYNKwETCwpSoOP
XIYjQnU21JosxaDy8oIGSty2wLvVbpIK0BTGdUG0nWlOha6WR96fJ1fIW/xMyc3M
LQcVcril9ms5eceDrDf7tmiCPamYnwG/oOSctbODijnFVTRBOxgg27DWiPOg2MJI
ykZggACKjTOoO4fkS79eJFElQUK+BQ+Z4+GDEyQZv/BnIWLYrxczeOuIO//JlS0g
tkImGv32pymmkyg8nd825T8va6lFMqFtLbJoGmIMr1sW5WVvJKV0ReZjVykzGhCp
NnWDqWSGhW3q4n8SgHr+uklfp5a67tDKmXl8OYY3vzjUdbGFp3JCE4kPCiQCBN5f
kGgLrY2NJEmRw+pcXswtP983az3cyjP1rNvxxgEvoL149V89eADUnKwPc4qy15N6
3nWOJa5cuYDXoHUnX8OTh58aAmTG1+ZbJIwn6kh8T3GFXi0yJlJ6YOHfX4h7ztJU
Vyuy9rmebX7lM6K4X+4+OLi+tDQG93PJbAh21SR80jxQtDPFLQs5lCtVfB/RLjQo
jgcA3joiJk7J/kbZD2RVS+/A+9XH9FuaZ5SiIwEs+htW8+pJY8+9VZjt9UWrPY8q
LYjGRdFn7xZZMIcSilsQ7UjDjCyIaja0/R0SCc5GFAK9V8sbAax98xWHNGM3qceD
oZq9QQ6lyo81uP7zqgMD5lVmQcUqRSIsvzLDu6oHHli+zzoeKKat0u7/LsrKqL9S
Vmxe8OfmS1nCRTA6NG4Ytc5erd57PsaridCqpMxn0taQUbNA1IFm8PgIHQjHbGNb
+znKU16bMotvWLSkz5WD/xl+kwYTD1wUrCN8aXhRz2f8PlIafksDDs2ispPCsZ24
EJwLstZZkcuU8iMwaSKOxPsCPTPVELFO/WVwQKjnm9ElUn3Su5PGDTOXkSSmvV+L
XKeapvEwk9NCz48R3E+R/V04iTrbyf4uhaL8S1mmu7azV9PqPhgHY19mBxv1e2mo
i/ykj5qGBtsEptzVzBBPzEKD2JdxmKpS5h3UUNEHKtqOaUEknkb8j0G9zFQRAvER
/M2ecHym4c5efWfSDoqRZk9Ry+qcCvqQXk5UmtYFKxSeDjUpEh+uRS6AkOTuj5HG
RNw5lftUfV8ivgG5s5cWG0sFtkwpps/hIaXWMrqL6H5LufgK81fiLDA1dIJmrKOx
SHbWbr2VJWO/7/6vq0Gi5e04ATCwpMtLoq8eyNTE1+qlQC3e3G+nvQ521MH8c8EW
pd2nyR3vJZljWda0FpY75doYmhOkPtxI6wEL86W1fnSFYvQU3o/f9oTbFwAyK8Od
kIy9OUuZvw+l3a0+i4s5iCMHXmAbUe3K+RlBheRiJu4nW/Oq2k1Emm8IeYIqBtp7
z0Wxrkb6ALWaasLzGgfCYOvNKzGzG2OKUTTYEHmJALa1kjjHa1F1njBze/tqVrfp
I2iaG41NJhdEh56XTPEJkvN6o/cJcXWtC6xvwABnyXbzK58s1a3zRNpoLrGnJVfT
O6e7PcaufWcM8StoLlGOw1ERgg3p0tKFgE0fgdP5ZSevgarcfDMYFM1XcX66wwCF
QWVHi+P3o7+Cqrz1p/sgYotkHq3j+nKYYObykjHgaqJFz+LQp/WqBoYNnFZ2kGFu
NXj6iiVtcv9Q1xVXnS3EfW/taBGxcl/MJA7hXrh00UuRi8I9EErWSoAXp+T5loIO
ZPKZ9Oyais1VHfuFGAg6ElPasXY9KBchSumX06Kh2oGbBn8TpcfNGPodKbzXDRn1
oDfOOpZTITjXf0OVJpkEFQouArujXjdrk2R/ig9XR3ccSAsW8UwiiDwg8HVPG/4K
B12c9rWnSJD/D0NG4jM129AQy5umsPmrsi+UXcIIKTJADsMjQmsAzi+GYKMB8s3l
sO95whdqeUBTCQ1J5mHiuiCam/EO15ip6OPFHesc6ivoKDY8OoLwi/RQjTk7MCdq
Ogs7cOcJLzuR5pUNLsKws4z4Gz0Pq+m/YBSK1qDz2NBQSqz3D/GSm5NWNKHVjEAb
dU7BajK9J18HQ1Z8VZ0uApDPc6OoEkWm9zVEmhVqyQIAFQml2N5fwHsos1JmrCbP
+sy8adurkW8brXzt8sVBpA2xeFOdPn95mrcAaQ28xBppz6SE5PBkyOu/Xkx1mk9X
PMuNlsB9xeJqjHrLvENm4QA1aVtnpDHCdcLHMg6qIRtq5uQh9LxJKJehmheRNMhl
bGAz5LMDMtCB8iCCAG4OKcCSq2EyoSrDVHtSww9BTpzl7vVrnoEEclMifA165ZNy
wgNjRJycsuy+ft0lYi+nQLIqdFaIyhLjX0cfFMQ0nLZYiO0SuhomuVO5UNDGsn+w
/OQAoLKBQZFGxBbbXpA75EUgzJFCYEwIAEdzAbwLeznUrdH0JiGfx7QTAJYAt7MU
97mVy08+2cNJLECpzFxXBHLLOuIo7wnrpvBmDwn+vNpyk5bVr7H4Len3thgqk0sB
zxoYjrWdfPKaeFOtkqGcUxYp/kDMZ8999SLx9QfVhzsp7CYeaWVbKwUbfennsCM9
hVC+phf8obHmfGq4dD6na8bpG7CIfBEhKQ+HzyIKC4UF7pg0xecvyVWWqhQdGVMQ
R7f+WPpY4Xaom8gmz/TQopoQLYQtjZSHLKvilGcehvq2DdCf8ek6VDkwbQJ/0daq
15GOQ2fYWrbBhEvpIiQ3ZmOu4gOTTlc7oO42J0x4oHrCOwowfirqT48ZssACqL7U
bdiH0baQO8rpgm4EJBqSxDytD78B2BPVjTK9tXCSTXwEpp4Jqwbzqz6NVbJXVth/
2D65nmbsbSpZrAlrf0CPCVqVZkXZZjI7Sf47MJPnWRpsC6P4t2A3w7k5MtuYOsli
160UqwlLpuqOOUJjQy7arquR7hP/V9CNaUUkIJsrB5o0uVqgs/PUrCzFtF4uBsWK
2vHJcll7UHGEaN7mPh+t2y1GecVQne1/LO3KmRiCQ3vysv5shVo6zzdJ9SHpjpp0
oAi6eAAwjsX7wgG96NiuiptXBZnWyDvMTGYxhqSIqpT6QMWa3BjcSWMw3b4aGJvQ
ookm3PB8Im5qyNJIc0SV+lb/xH2JdIEr1A6jL6pyIqeRB9dXLQz8sdFj0ELbWcB0
XuwW5TX+5Y7QyCg7g2j9sV0bJCV2y7k19549fJG81Ww1aCp3lSW4coxGuj0w8FXX
BPZkq/VF0DxEsnHxaqyLnSOZn0wrerwHB8rD+jhNwx3h6Z/3zdQwwBLNX4aAKGRT
4VBMCUi5d8wQWIB4Wx7B7DW9Wj5v+sqLfeS2RqE+uOVQa+tHx0OZl6F+eI/+QjCu
4LeF6A27DLE2mKGQ+pMDbyQ96ohIPCLdnc7vD58qt5bvOMFy43bA1/WgkP3cs6Lj
UfbHe7ADgtctPZFJzkNZKCxvlW1Y/HOoezvuwZ4Mj/5ZUmrTbpmG4yfkeLS3+iIq
RnH1q6kzfVLm3rfEI5vT5sPLR/d7wi2c9ou5I2ZFWiDJFIRxZpMhN4f8gR4bgPNC
NWJ8v1vH0rABMzdLSrXSdo7ec0NbGWNTkSPz070iuOJkmvE1FRq0Xpf7uqerhbgq
0wMNSosKGUDVGcfdfSLKogQ7IXN9R5G0ejY+Mq3u4NgogeDMbqX0STAhz+obe8ak
HkdKQPaOtB4rIwn6KsDhLmJKFoEA+jZ8rkmzItJUNZ0Kzcj/B+XohTuIeya2+8Xm
nV5E6Ns6JJf4mqB4pBEaoTo6bq0/4FSnZ4k215turc7djGYKDnAJLfkhjiw4Cccb
MfIf+vjwvbOpMYvmw5/pKsRF3sZ70Ffi3mgZrjtFpyMO9ggG9qsDZTe32YkjUelr
J/iUYn5bJLKTqUI8OKsZyNk4kSDw5MXBvgTNjjb5NPKxsMKiWNi0Z27iw4g7eLyd
o5iHuNpgeqU9kPxCyv1fE7hUwZZtVfwNO3XUpkOLIA7PznHdXn0uCU3PYpT4qBE7
7QeO2kn2uWjzqUiLPfm3MB8xYgsNJypcZRNsRy4bp2ymbX1Hl4As2K+AxoBYeqkP
TeyI6f0AHcdpPaur/mTQY6LylAHKSrO8HRvjg/RixIcSFMB3B25nWr2fcPs/PP6s
w6eCpR28hBhDL3QhPwpo7+rQDEAKoyipwuDQA0ISmYKoXGh8KXtesp2NHn2HvMut
HHOa06kJp68Z1OnRfZTsV1X05jyYGfo9kp3+e8glNRy/79vaL3griqzfQp+VcPo+
nxfymYEUYAmK8K/7KbH316TAFSQUCXWFA1Vpu5KNZgT7aGUPEmoclf21KuQOi8cw
Dd8Db4kLM38/JcsNLbEIAwh5f/ed9nwhluvOHfyiHwwypgplBrjqlVp+j3Aj5QiM
5ZmNZqaq+Ks7/X2HEKjR5TSrZqOwI1AupKVY6AaH85rCUsQ7RBo3bagqPtMviziy
uFIVSXiKn3rpuf3CM/7oGTnS1KXNuASRiA/Nm+wJKBtJZa2/t/o/J3dRQq+rJjjw
d88m/90igEpEh0sFqWNnZ+zTZRzBYyC0pm7eT8fu1VBLtWJkQYwzXewZNwl882uZ
z92t2A0GGu2CXi5siVMJfRN9Il+U6JTrvHCAPGoUNEr83e2xseYkcjL9hn9bEo3w
5iT+TWfoF5YJGAIUdmew9w8wH5he27MSfXX3EaFJY1p0Jcgy5BrY6kB74otFXb5v
aBqGmNNw/nA7I8hEapL0ixaHECMSxV5AIRFwTWE1KrDzsKKDZSRk8fK6gGHDw2m9
KWjHNDiEuio2iSAIeXzZVWfPmAMHmt6j1A88Cql5OjsKLSpxgXj4PICR63BriuGn
9zcR/+OiJzU29INppRANYnKA3rKPlWGasH4ykm8NcCA/3bsgfuAR8Ei2prLJAXbU
Rtw4tieEre5UwA8X7CtkVktSmzPhn9HvXUBa/D5zocR+ZItG6E/JReBBqjI8zw8Z
4B9lij87nN5JPRShKjbxWiMY9pQYT1BBGnuLIHr1yl6+QE+DQJ2is/G40aIWStMJ
9QsCR4Q9cZ555I1cbNYou0kTsbhDwsWH15Uy7oNuBSJjTrSjcig7/IoTKhWMoGbh
y9Pd6lV9RaphrkQ0ZEmdESB1EFRjPJzPqyRPeNgjDgaHgw9tCJHmZcA4OM73nxaF
Bget7TzjeVG+4JQR98+8FCzyvmPR8GPC2oIbm0L2QFB8zI4PNz8E9yDsGar1Alz9
ySc42Cnni0iGvZ1l8aXZJhLkrZq3WWn3wsXqUO/BgOSKO57ilWnxC27zzYsHbPBs
JKVuy2FD1VOXx9JlyDv9I1cor/i9Pq4kVa48G+xt8BN6piHfIypsxfVq6+W3W6q/
gdfRXP/628MgESGQgRgl+dUUYIcn0MwqwLbXwpj5MRcaLxwSTQyICI4tmZVIr1N1
pR7kUlk/r2Ha33YDyuLlv5g52zJC9Qeq203hSJStsnzdP6DxgzJOT4okWnOscqZg
11bDRSsDkjgCEE2/VpMp5B4jjUcoWt4CTq27mp1H+/9DxqbSGDWiCHjgl/F0kIkB
+cEKHvJ1wBzY3tdX9p65VswE2e9fcp54GYx5ETk7RN66yU4OmYU3TyTqqFLM9BIX
E8PLVsHGWNPGyJocRsfUcFUZoSlF10bIl5bvCG97+dj17SRtBWvfqyIVbNOwdOIe
AMetmS9AfPMPPodJlTGPgftKuAmweRqkEPwVEHYEpRoUFg4D9ZrCnbmQezBnmTMH
86fwhakcv9Cu0S/BKL9sR6pFNkyW76aJoYFaPKVlNb9G4d+m3gqryB300NKBwAMc
YUg3FuYGbsHi4P+xiWGEuNs61Y6H21q4v/033DP2xhCQChnAljufo2Q239Mp2kv7
kmqI3iKLPb9H+W+lMZbGhR31Agf/G7Et/7r0U0vC2mDP5tm6ECX5iosvK96WcjGV
dR4wfmy9xf8g/g1AXGk8FIl6VvTcv/W6k3CAw1hQ+wUzD9zvoGMq7kpOuRKd+ZKN
Z2Hq7XnoTrO7XyQneC2/G4SKLTgTA0BIEXctVphGEM6r4yMeS8WzDRSzkUOHICiv
v33B7zwWg8Bxl5JtrlyfHdrp7nhX576rbNxVTBK9nQskkYiU0RaTl6GFg8gjo1FF
ZE8Mc/b6DeZ72nd09jW1Huv/ESovIsY4OamBGosvNcnODe+M/I70xmsbHW9OubrH
s6rjpQ7H2uaXTV4W4Gywg9jB3/X2v+XFJHbodV9NPgXL5hGI+TFgYcUZFDp3eoHt
xgd9ysbbB4Gi9HPwxAjVYM43+mZ/L+9dIQviIL4gF+RHVKlp9+kpTZT4Y4WcT6BM
vMbniv2yHgUGcTh/wcNvwZzn/X7CrWq6veaUqJETS842EKvg00+zweLxmFATEzHv
F1UypLZL/NciTAN4D9aVgwI3RMLGXj9VO8X4GeWt4EAVfrBMyRRvgvGDV8jQtO/e
2VdRyO6M4kposatccjM53Wy1KZr+5v2X/RmzflPYdB2iE+xGV+L2JLJCfFGwNhOO
D0rgpTBqzNw4R1cCIoMlHQYM//Vev5gYKnX27Xewukyap1i0MkHLxguDM9G8Syr4
te3J7lzhcBUdS2XmmfM+Afh8g5NQ8Uk+XWonedwxQZFs+qFjTBx3NiwVdkbhSX+O
5kAg4A3i5I/5N6eNqd76QNAEZXx/Jzg7bjOOoRgV5ZYcH6b1S91RGIQSyB0jomQM
9FfgwLBCg+SJC80o+32O+PLCkA6CWnNoIJrU2NZndfUsENz5VhDnLb2tLNOqGGC9
zO5ulngMCFEQKBYezEFe5w30VCjo3mnvhUhR1uhWClzNq40iSv/5EypTczoZVika
EohIVIsvPNo1OzSGorsOf6ObwPfSnmw4+vgXx8q/wHLGVGbGsbrTsfl4kYfh0pfP
HWiRj/zWq0K0It/PP+ChriJxoibl6t1k3Q+F8xLRp+aK5zZppBEFNWvj6WjdExi+
f9uYZnpJzQh3yrdwgpKRN8qIneKLnagLprg7h80L7SvjrSj5LfoaLw9vSWeGrYzu
DPTl/U1ZiMf8MN+xhpcw0Iusyps+F24Khkc27YOeijciyAwhD7IGEcHgca4Ql8Vd
VoBd2548/BOf+747zluT0ZXT8DlquCyRD552O+7L333jaF37JLbNxfnJK+ZvX2Gu
wH0E4nZN8FZ1VlGgHpuGcnSHOEmttdMBNNka+65/TiV1TVUc97yOrNcBNSrEseM1
/pGiy6JY2vDOKuStPCIfxjNgYSfcP25/X6RlWeMlLzwc/1a1NdEzTIfxmR9RGQN1
3NmP/Ot5hEiz8KqJe5NSqx6XgyGefzMePC65avpOPzzyULrASXOhQ5Ol68AGSrfZ
hu7TAx2mQRQ8V5rny8IuYSYhxuskcB+gxyh7rLuWrnfwFn3Hc9heOMI+qN977jGY
1NkwiVDTM6HEGhe+wWi7zhvrEdYnMBdxqsdzismdPbeJJJmr6+5t3BFbm1kIIsle
m2i9mwiHUwaoyYyaQrzL/IinPeTIBVPUjmDS0odvgIC2moWlYCj4NPQEo4yrEj/W
HfIpWRz/iAldF+W2GNRIozcQCsx9Htq7C6PHFdRRplHH1+CERkzQPqG7sPcw9jzs
3uz2c+Kuu8jqVddWdU9awkBj4xkr51DkKHUmjYpSQVKgu9+4T6GSu/+5j/zA2S2i
uR/shut5vScngazhaRlgp9jBQU2/hVCRtEZpNWs44lhnpFEydxiNJfu1eQLBa4pl
ffu9Q1MSJa8tmuUWJLQw9IzTzEwUY0Q9hvAtR/LsuAKVxTXtLQ6kOcGpNphR0eUv
E5IqIZoCIc00RsGJ4foX+fEvqJ34Etm9FBiN9amOWb72dmoAg7Po0nMRIJ8yrykR
EDuL0o+VIZBZvZGMsc+5/ND+FFgu1ZOavZ6MyYxWDnCR7wBu9v9o5A6V9n/rlvMZ
DBWCd0eegMonAZ50sHwRmHgK9C835MZXE78yjc8f8qhzV7a1BV1sOJSoHvAmDz2z
BOKbKP9Cb8Obq+8ehsERA4XJ+xyyZ9FzDeuoL7I8ECLOP6NSBdapGI2uBsPwS6Q4
AwB9TMOGPFgVQ/HiPLAl4Tqd2emfolANfZ7AK7LuGQoWl3rkVNO7FjDpMHEx1mWH
kcIEq5E44CIFLwBqxLbMClFYoC3BoOF+LU63vkmr9EneSxn8/YQTI6mreN/FikD7
E6KJwKM+NzJ98fQQCUNnQDO13w258NuREGruL+2S5ShmIpljn7Zx4JhjTau24DNl
YKtBeV/4azBI9+ZbOkjT9LGwDALb/C7ieFNUgWAo3EP0qz1IXsisrpq5NT2MpsoP
Y4HCQEITBRJTjkXYqnV7uFjTuQGSyf/dhTv+bhdiHQIrMoiilvnlrglSNiUKHu+Q
G7u3DKnaKHnmbaUtLfdDe+5/0rB84aSCpuLtCq0j85TU05ijpzY/pHzq0y06qtYg
XF68DpwtEmSBdCtzgDB8kinRy3EA1EzBYmu8kk4AU6I0maBUoWRbHo7UNQJGzrnM
dzUs5ByMwHUj6h0eKAMvPlu7svkzo3Ncg3ucaey5pl0yvIw1xDbkRMQvFIXVLbdi
E4+lrwRNRbaGwp4wfuLRjpz9oivmCSBe60hVWNRUUL6FEV6sNXYuVqfKeTOWm8O7
qAus9jbigYR7msueUqIf6JlJ4WkhMvGmgzpeRCYMwLchqqyNko3Jm8dy3N2E59N4
Dq/AbQGH1Pb6O6tdjqdr1jC2EZd2ycokHl6sxZR+WO50hbGOEsJcPbOYy0AmO8db
YQ38wImu5YznW7wbgsNgMOB60yrSKZoOuxOZL5goEyB55yYA/ySizqXnzF+Akz9T
iQJhv3uw6ahZasYsWAiFDS0P9iUsippVD+CAeQEJ194q9uq6BZ2rlQfJNPcPH3ts
HF70qeUjykYZJupsVOsQypby+jaecpd/BncGoNcX5ociI8t0IReJjt5c4+Gxrdi0
BIoKZjhktqVGm/pmY7v2X73ek80zk4Fo3dHpMuNLciVsJPBC56ATp7cObRk3BNle
GZ/l0iS7qNw/pLVQPtOaZxdfchUEYuEjTfuG5S6xOi1qMj4DA5oKaR8fCQFGS+RC
wIVfp/nSZWQMOsDiyi8uTh33pQmAdSJKVR8ASZIjSb5UXg1vNNsE7JSB4+C1Auyr
wIE2Bdu7YVqD7Ss+saCi2Gngewx3q3BtlCrORvsT0bViQER8kwphjqmp3W/9bx9P
kX5o6wynTRmGUPHuh+ks63sBE+vd/jgY9r8ikIZwOq9q774ZbhHn+lVKZtkV2VKV
crv3kUlqbYc/WTZ4W4OV1asbmE/vtaWHVaZdXN1hT9eP9MvrXaB6M0knJ1wJYFZF
2NouRKd5w77rXjK9UKq1RQbcIiuF4MyJms1PHfJR4YypK3et7cQuW/MpShVXL/BF
M+bMzsOaKQj3CNruWfiK0YKos0kxzn+/ptcM4PF1feUXSftmj/wT+qmXZk+QR+KT
SxEAyAJnP/DfdUeFg8VEZcYW6iHsmAc2R3LRokgRVs3f3ThIG9kiOSt98GdhrDxN
TK6/b2u99YMYfMa47ddTsB2sG+y4TzaTovOxqg1z3N4J5JEP9JIbJ/hsuAzA2tPt
PMvh83mfDhyJ8ProobdP0nxpAc3ay2qRLynTNuhN0zYRL9fdsfD9TePTErvcq24r
pGOGiDhIw67HC4wfzuvVTLfr/mD2+hcIZEGHXk+0EFTp/qcLNOHAZ2WQy8NXupe5
G+PaTsH7QlFGK9gHQbj9ee2hYB8Ulh1tVl/TVCnUClDphlztAvFdp3u53cIm7cEU
G5uG4mIm8J/7neCJxeQ7p+THqES71irOp+6/rWU/zqrzzdczk6H8iQpmUuMzF0ia
CjLVZpJgZAz4yau1SDbwB43DZoOd28hKud/a4xfMyOW6IvJ9YuW/iwVn11QtPOQ+
jir/8VHjMjkCI5pGbbBlvYlmEEaKYYgKuoF2ZDeD9Kq+QC5bBnk0DR0OrSFzk/9D
V6TX0qGb74IcR2OwWq75XR6P4ahEIVnY9CxUPYTvgLLK1lAW2+c12L/GnkM3g2HF
WRy4QUMl67qTo3zMISET4J+lhff5rE+6fMVhqgmRWoYx618VIVNMRR2BZzPNxCFp
3SZ1iKA/1YnZzLK7omcmfM9yILQxdyX4GpYJ/9+jUEByCl2UckxTkrBNPyZembL8
Lq/7ZpUXM7/v8ljCpei1oTRbhZZ2VPr4k6mYXkgWt0F+UXhIezCOq48QNaJblv5i
HflDN58ZHfu9cUGxDUgk6vlXnqHvK52/hyfBHtiIb6Rx2+04FocF9iS9rGnPXC2J
3ZRIvbc26QrJibtsgtPBkz66d/urDtHqIIdIyE9DTHKy/BuehNS32uMZZAa5FZXu
wq3uQRFNYL2Ch49MNvt93d5LTvX0ARf3mQe5WTJnYXEY4QmyK5b6p9eMpnckxd51
2mA2dHgIFUs7WJi4l+gCYClKVB68wbGrxnnOVLLCEy4hiUOnbyCtdqR2tL8v3o+L
PxGdODJDBtMRYgsAs/VmXVQlITg5G6ZUOqpWyT670teqpKjzV7i3Tk0YdhBx6V5M
7gQsvc/IliexHLsBVpDmKOo9uldugiwAqpX4WSi5g6dNtWVpGaAh09fHvx3QDlJS
HZZZQ/OEbw1KWLPkJ6KmgG7t4Sl/uwzryJLGLu5lCnWwim8KaHtNxeKErrfkjlfP
rFWjNEuFtYRGG6Gq7acLhqrOKAe43epFOoDGRVykmJd1XmfcS3Um2bJ11X7ZvXKw
BcOFvt2tpjzsw9PPcUAW7jb2H6GN/Q6XxoeCY4GEDgjbjXW7ojuAJW8pOZFni+ez
ZjbA1io3d+O0PhLv6u7TckpO+9DaMG7p2FRnpqzO1U/76J7x4kzBwcmtqIjjC3j1
YD2dfm0suYJf5Oy8qmPHLdm+k/b4MKYN5zHUNmMcLqSzS6M5yo+pXGZ9IicRip7Y
/I4dLHg9OU5kJBrHYzRM++mDa0e1ilXe/7LCrJNeCC3wrbXmV/5QpXGQ3a1NpMWA
6rAXlB7NK3O8DCetp2QOXYO4dQjoDUEBCENJ6wnO/7zW45VHtGq8wVArEeKKgjNX
HTtOHa5HjezoWhfPFDFzV1HuHcHG7aO4DxCo2rmgXehnw+m4NFPjkMpWbOVZNUTI
EeCH+6N7bzv99zB1VPLqp31wqY1Y5SuxgAQskrpEf2pzmQ5XoZr179AG96oA/7RU
RKioGdxockKeEsCUmqU1jo635MOcZmkK+wcH2IyhcLcNUDJdlg12QNzFQJFdOqiY
TXjIBjTEsoBq9bW5m/Z2Pov8tcFxQRnK5nw+biKx0XmyX+exWnkuGZCB8QAlJqCv
d7nKc8ZM65rTD2mnyWz8zX6bz7VqBl72iPhemz9oeZm2dt2ddgYmAiTk5o7iiczP
JIKLi+Viuc7lcZsS/NRiIamRZUlKC0RRq/6QoTmS+rkYRz9WTPml62nZNiTlXEhO
kAIskXciIVHHrThCyCc+J/kPrV3OaQJbRAyd63se7b2U7iWgDkcy7nOeMjvAuJn+
vQ0qBoLz36WQCCYZbFiaSYz7brP9RlDXn+9bEiyOd9rpVZ2ea0Zl/uqOlBczh624
Koa0WQqhd/s7Q2OdBRR4AabAvFNkbBI/Xlrn2bAX0NmloOo2X/wmNhe26cShxdAb
7c21O6P2UlNWdbK5V+RbM7IUZ5R9ciLfUwmwt3TLkJm3uvXxgX1FkyXE3uATh3ZO
MYg7QUIsrrm01WCFwbINfwpjzqGwUx4JwslYw9RjuKlvBmKkYj2rT6XfL3t/2QQV
YP87q+TAOFxnjjRCR39GBj63z8wUyjjPx1djaSMaph4anR5XPjeHQWEuAmsOcaFg
K9SVr0ybCVQlrzzWhQhMwemGq4L53jibH5ZjXFJMiPsGjMmOzuWWA9bdgNkNmDQh
aGdofE9jIChTNdCr/Aqk33GkU7ml4KlwIm0zuNHZzi2W0BZMrau/PmhrDJZpmSjR
rbIhWMfSchY1pGtQ+/Fr2qOD61PaxVTEbL5lNCmmgIQRGw8LP+WbrnKCsz9kelYu
3AVCsxNbLVM58rL3SBQ2dk6AWSSrjn0JzzfgywfK/xd13vqLtuw/4TQAeVn1mJcY
YIBwD2RDSfa8Qy6mkcZ/zkAW3D/syCXG8BdCayFutLH/JUbk+0Wz7dDqXLU6td4s
0vWHU64axyCm8zl0cazoEUH08QCRqe1B+aUEMLj/Khte2qsDmDG3VoVb4OTydI9c
DKa1JPpdN7KawTPPSZwn8cKy2GuYDEYQ7rjwWrvenkhLBzvgzn+rU+bZGYDieKlM
I5nVF9p2W3dIGx3UdEo3BIsPUBM8a83L0D/4rPvVABpSPGfQ1G8V5jQJ8eACTls6
ul05bttJDzBJYTIzthLj+uvTvdWEVUh2Fpw+04dRkCN6SWQreAlPc9oPEt7HNBEq
bsFMGyXhfJ9wQaXGSmYXwtbKMQq9mirx5xIWt8NX7Nn+N0E2GLwrvTLtX5O8khs8
vMes6nzBSpGS0O/MMnvY0op3ib6BsCvHJO80XzvRKXaynY7cUvGSDBQpERAKOuWU
+zZABLX87iNDQenPvl7qrCxZZfJ2/DaXBZKgcGjyLvoBk/T5x8ugWl81HDqWaYk+
LZUEfdtEHZlWK56Qad9Nf0aPdg5vDHy27ZkuCNJvSAduzgpzjG66RyCYobReI5NV
AWFv281Ehc4G78rZamKif9hYv+VKxfJLN3DChIYIxxl6kyE13Gd3CpZKIpToQT8h
54yL5ZWa6ytfuz5AI7+2VKfP8O3jxBbgENDrok9q/zwMQf8oYzBlcL7EOd/zdAj8
NZj07z5O1to4NqCkhzTXKyL8toONLguKi5ns0MKjoL/yFhJaxXhTNJFTCYN1+KJ8
4rWQ/pxOo+RpmJbu1ZWaGCQ2kqmkm/DYPdFnwbDIWCjzoheCvK9jLIcj1VjmgN1c
LlHX8o7fn/j8wPrk5vOYWsddTVEqlvvM4/8mTan6aqViZx2V+PWkk5jWf8ZFgH3x
TMwWmH4JQO/vZMAx47sCpvF/7TYksxQBJlom6ixszvnJ2za8BuUDL0x1O6YL9Mpk
8y2EhGeWv8yE1MVn/VWY9iv2BDmvT5CRakx1ISF2RVprycaqsPeQ1rOaM7mHJbZ2
ir2tChIPOzycjFjRmt6kpRrlsCj9ZjcxQejL50O6OtBssZLqvwGi8yJG7rPj21Rb
q15yW9tCiS/JY/Orif4Qv4/z169fvvya8D6Hany8xs+jVNxGwL78TsSWxST1ide/
OQSRsunxmnfDSW26Wz5shDDoyay/YxxeIwNpATtF6jCZDaLSlEoAOya4LL4LSP7g
cgoLfSjCHVl546v24CfaIfSfnpk46iPxWpgtbTyCyhufL5qbJZseZONY5TjPtd2A
jD63A2VYzaqkoRTTW56iKvm1BFIogHOzoAPJ+WRykC5oh5DJG4R1v2NfF7QC9Yig
SvJB3Lk+bDrVBfeH2u9N9v0SbzEf+DRTK7IFnLLdjvZmGjmwK/3/QFTd1oSl+1XU
ZoWGn+rs/Cq41gmGd+yMzIEl0qgZ9N3fg0Lz1/8ZXiiftKs+84KnPchhiz6SCSqO
qTIOtCuNnmQH5jw+W1P+xZo7Z8I8mN3lrnvQlhkeX2kM13OpvP2VYHINNLDl2i7T
NBX45jtXeeubBF8Y6UWS31SHnctiN7VMdxS2Lfi0PF/YlK0PHueCXYXCHMrCVNR3
nlqvQidZcJR6TnCq5GHjm0WisqmhgqJ1ZKlfH/IrPL7Un8B9QB1iPpYiXzj+fuzI
GXTGAUN7JGi3d/DRld/BYS2z1OrblzlqBHoKXYnwVTPb+V0GcindxFil+PYqPImY
FPJ/kHnvkeKqtE2hAWXoIbbRGPYh5Hi2A94ZJ/k2sm7keg5GYVvbTfniCYQJ7n3o
oYOwFHcUtBvrQG6Bk5GxJ8Pkcnt6n4v+8R/4ZI8B+piiacMR4fIn2xXj7e96Lgb2
7tgv+2rpnt+DYur7mG4E0+9rLlMxyYjorBRbHlsZmbZUOyRZYrmDSwdk0sUSifcv
M8cn3ssIrA25X+0K1b3GIez4ycRAC3yfmy0YaG02m0711J2lfSmZvHZlbw6WaY/x
aBMN+b0whTId+pEZkMhl0xb5HkJJDKMDLO7HXXTo9YpoJVSrEVGt+aZCnGZdgBvb
rou3U8CYelGEfXJuaZFH/wXGpOYa6O47VmAz4fA7Y1WBwE4CZR5w5YCyalf7XIkQ
dIh8VMHvxnXpnMdVZjDwO81IB9oMdHXslVo5y7geyQ0azbK9XJRxuVNd8GccgDLt
Qe8oK8l4rhhHi16BqbGPHVGa2foc2Jlu2b5287hEfCXNG5xXblAXLAThm7hI9Ikz
RhQNlkzBncoNpoIFYzNZ+yfZGc22l2KwyOzm/F2Obyxz2xQCVwrI9U8QUbaCFPJj
oheIIXmj9+vdi1V4MXV/1ic2jUjWEF38X9i3S5D6j7BHmf5gZyjVdpYHAyUYC8UU
eXkTws11X6C/InFWpCZBvkIog9u49WTaFBJh4rRwsBEdKJDlmRYgOZADmVJz7W33
12MyJUsTKGlqmSzJgvkFp7Didkye3NRj6O7MSW1BeK3TRMIMXxuRCY0slPQErUlO
7YOVzYiDjalZY9ahl94up9TMisRCxMHOfLKIlihveTCdZyLS9B3FiqrTUpHaac5H
3tlm/n5Ty11P4mAlHzYNf7+a5o+0NFNDD3VdCXPRHfo1bDl5wSwxrxTVeo85MrSh
ROna0DI++6c1VKhZlPfSSKJwypNWd1s3D9izMf+kLw8Xl2DYGCRPdJfKg3XZUs/4
X+wm3W4M3zUCziUZIY3gYC6/4uREIo6BTuWvlhgO02gumQd6EpMlYrVdvPyvs2Vj
Oq57JMCc+IYvlxQuqiiSEF2eRFyDqOqDbmLIe0jbIB+O9bVkRbqDE4Q1qwRT1OEK
xxrgBfprgDX4QZvmv9ezyGiGGe5loLK8waXh1ZdaM9bJKWTNYGKZqebcv9dDuXXW
NrGJaG6WGbaMEU4iCPtT9I3KY+ASqZdTDfj6JCRxTYSijge0apzt+oZTqHeQs6bL
GQAuR6F2Ba4+bsZxu3O2PnmRmKbin396sKr7Zv+T7GjA50F6Aqm+/z50+dzQZuhi
9gQDoI/21NdRG45yeYJjCG0EQGvZcRy/jKbzx0Dw+pp0wmkT8o/epzEhq7g7/HOv
GMkBUvO8KLfw5EnHACoaCkUmrKs9SnXvs/Z5VV2IfN0SjZuL5P9u2C4ORfnlz+ug
hUFxx1CBb3BB6O1LhlocIF78OX8wgMc5E+kQE2RswAK/q1+4qipxKtwUIXfwszyj
esU7m8kvI/VwcL3la+u666RzsQ7htbinY51rbENdGQWwX1wCm8q2u2z8TWB/NNVj
Y+WFtlv02H3qaxclp1ENVnswGU3iTvlgi4kskCzfHo9h2Wea7arlpI2K75E4f61t
mrmwZ9/nUXp/7PyhjFRWgVq5j/B9+bZJf7v0yH+TBqZokPT3tVF1pz9ypY/3GI5c
azjQeQ7ydBa2N8Cua65L5m1AagXGI/YefH3zTpxJLEEAR6c/LP1AJarhkAYYPUmF
XxrkuArkfs2olXUDZM3NMcUW5kLKX6eG5TKjiXJEl9fL31csvkU5cbBO1jX/lIeZ
aHo1XjTgQeKv1M1FhPlrlDrJToUJuOq212e0IPJEbwqmToUxf913gWw9NSGwu8xC
/ei6YR6Oe5GosHI+xPoabOMxtdCxHQTIMuGC3VZygjJEPoP0ZDIHzMuAyjcORcW2
m21sBIKJtfj3VjVuSnckj5lZ5aBqizDX0qOwelIjhBKjsUsYExfq/qLXXlkmPaSl
DjB7be2wBCpIuMvjIZhumI5R3RMmloa1nGw/8Q3xHAZBISmsy3liqSmNsAo4WV53
7FgvfgymJnONyboGNtccgOtWkagYdqBrv7TUK9iFfsT8RwIzywE6JwdeTsoP0aUr
QGn+BbgRw7kJp6dpOJkf+uNzF90QcA6mvKH8q7I0MC+KG0uxyLHHKS8QgHddr60e
CuY12IemK6SH+v1ULlcIFZfDnbpZib+rWJhK2UDYaTUqm7FHdxiHAoVHnCq5YiRT
I1raP3Gd5Fm+FYnO5BeprHh2G8Q3dUlef/cgwPYUCi5RSfDVCCTKGIr9veUgCAos
YNTuTDwMljJcr3io+Z3btPL7Ei0P5KpwESIchgOlwwviNkBbM/HlY2Ue3synggSX
FjZHdJBbDqCzO+xoTIen0Wg6d+zA6f3hhl1Dd3ibVdL6BCBIFaBhDN/UluY+D+3p
fLU3et3cPHiI6AWmKU8cwOfpy9j/+hzFQNa6LlRMZIwwBB9tTh+PDZieTv+OPqsB
/bjqU+t4hUG/K2U9Z3XudmhGr+Wxk4shr0XHchnR/zQaJj1IE1iuasn7B4G4dmC0
6oYzC6DBMpX6B4WY3gz8Ppu2LPP93BjvbC+9+2k2II5fWVoyk6/s/NL83dy9RS9y
9evgQc+x+Z3Gb0qrLu5/2udVshswupd+6mJIGcdo3Fu0ArMl0QMg+XeOvz50HY58
/GInqjCwNY2fXBei55OE15eUVlv1b1KDU9JHwpq2rIjSey0TSTi09SHgRrN2uLEf
e/Ev2MckJm1JET8fDK6h1V8QWcSFoyQvBsjM/1ar3ZfYgxiN+WdQesXFoUwUl/mJ
y+UIKBPmt+qb5vVzL4jSG4m2G/fBZavJ4hqfmENIL0G41eEF721fI/pAvYVZnWkw
lgogsM/gXXJ17iym0YPDSPFllhN2oowj0jvV4rtwF2TR5z5KgkYz51xOprTOJhi+
nOS9VdHkO/rjv1ZjA8L7PUQfxYxDLzllBkQC0jU0EL3uGh0alcW/y+HlYJR4Uvj0
2K9sNQ+a8PLSUZLkAkJXuP3pWQNC4Q6EmwuK7Q9dI/FfMe9t7k6ZeaeB5kFT48th
6H7unHXedL37NoQl87+eFX6nTtMfmJvzlWdLm46Dhm8/2qtRl9UH1TJorcyXms86
kMmMfJJAOTAUKIDH7VHQ8lTURfkcKBUMYeE2QFmCdA5Jjz9LHatD3IhGZ3n8eoba
VQIVGKn4nvSyB/pBUnVisNw896CROLdmbATMdiuTPXWJpuBeCqB0afHLTlx1fm9t
LWPIYo+/VAdBjZAInhCbxMZMOKIh+9vi0IXnIF3LhsioGhCU52xdosDsI89SJSza
qlNFIiHVKAj0epBbTATPBYwjhIOQrHm4XZ1YGlaTyzomq5/QKK0aj/ayAVaGCslL
k075qfJAeycL+QNyb8ZZiZO+t4tihUWx/9sX4OFl8QsmlF5IEHNfOw/hA84EszTj
nHf9dvpG5InFdXz5OevK1VJzJh5hJDQ/WPeREcb5PM83v4Np3pr6Ub4U9nKBnKpr
qzGI1f9Xl/6sAH0KnFTJojfZ1I+ao7ube5QtRo3so+AjzOFN/clEmDnlcMmVheQD
j8zJgk8w8ez/G8Mkt7kvdwbVpze5lKVjLEXyRdRZQVXlbs2+zMJA8SurNkUbVfBh
mscTOG1sFztOvdF6en6bdJJo8OvukelXGXhQZiDtncIkG0gN4L8ZY9lwsa4kKsTR
g6KIEwIzVGXz7/UWca5yfBRUvkUDVTi/1S0rEFe9tSExQ0eLB5HCiE6mVmGWIZCR
t6l0mRkGXlb0LekF2V6u31Lpw8Y4SVSuBM+He/QLBjevRl7UKnuyIqz4/8V8EfLP
YLC8Z8bXSOwMasWbtAC0ba+53RDYOETpMGDe9gyWf6cZev56Bl6LnCbj/Who7Iz/
2QhM5dcQdaAD9sJfJljBJ0/ST5sEKlZiQYQtmTC3mPk+7UmiosVLv7h2xLm/+4Kj
eU1F2idEHd4KwcpasykugTNRh0oIIMKNu4JnXa9YWzgQqOUgjLqOyyq/UkoL+toU
ZfDK4CVzI9dg9NskL+EjKVxqUhpaMGJwJLT0mT1lIlW0FWaSOgGioopOPjx6S0ma
4PnVBIFH203i5HmXzyvWXxB6nLknKsPEuIVjR1BvCh32o+k/F0pCDORSkKIpi8Vd
te1mwbi1aZsqZNqyaNyM6WwAgG9qci6/Jvbjo/r2cFYj7596m5yG9zsMRQXGvShB
UbhFfFsUR8f3J7gPL4YEw6OPlDKTaNIxw0ZbEq+tbQr/jkn8xT6xD2cgXJZwahIg
oxT74njuqiwA3G/2EAxHwM+YBqX4mCQ8wUxbFC+fe5T5Oc5iqslkEo5fCfuES0nd
SJpbSaY4kPiUdr7tPkBIQwxIO66box7yGASNwh+ohYScRHR+cVEzkbyUCZdhku3q
0JuJ7rRx6MMgMFQYc+9IuL9Al1iiktY87U01UnkW+/6KCCu2pd+gXdpTYWo6ryT9
+nH1R6kHyIJbwJdaMTzycmhzZaBqJbL7WqCrsyCpFSXnfBiRLdQiyApRMiR478b4
PzI3wlPJ6jbJCl6H5zuE671n2OcfnNtzBA3LduEtiuRuVLRLowNK4ZTWJYJ+dMw7
8ftJHRozv16oGQlWqABUV4+h5E8Td81WNUNFLHKV2gBzG/3ErT2hqJoWlXG1HVrx
ygfbKiLpnc/lt5IyRDTMM+GHGELow/QDTTGtYg2ZyZFcX+jp6pA7HS86gQWJWVqH
vvaqzQyzfi5eEw8j8a2QdCaeqbOcCuP6wfoSDszWq1F3LLsogsayga7GcYq4RCZH
q0hNSrdpPCQNZXWKGOqTdcv1JstCiffn2vE4yvp7b4KpnUuDY4f3x2KWVzmmtxQN
SrKlbIqoAu0y+YeoIEulSezry137ZUPMKZzIfsfbAB4MFNi97ysELWfjzFVezbtv
HD15NIShpj1v9TEgaMYEhr4CowYTOXuugwMqvuly5e/maKsKYuEfdGhRTDY3CXx+
OV47Sh5zUdLkV0uK2yB7wHlCEIU3Og47uYK69Iq5uQT2bXgNxrLUcksQDI6u1whO
t/gy6U+hd//ChUzourmrzDDCfFvPxPBiTvLPbHRDtOR9aoZn0qTFh3IUrVntU99H
YoXpAhaNCXre3nTr3nGS1Jx+mLS2vjlDsn49l6eD411m03RnzZizjbIkQgfzLM7f
g+oP9VWRS3e7VkYbfU8VFgKecqBJbysooDnvPffJJ6NSusnAFNkbkcYCwNHOIRpW
sIn2NIGge/aFJdRw/wSKvxJNoB7jJu7u3aKH5UWb4cARD+HRnVlBO/CQU+gviyfs
5YsJccGS5KKSYF2uWvoGRT1WdR/o9t5Oya990ZYKBlUKOzoWchqQR0WS/yqnkgpJ
nRe+05CjYBARsc/c438xYz4ZQbITsE0Z+Lg3JfRYhewK/3BCOzEFVXtZbm0EqRGB
+J35OxKmd3A98G5lvATCDs8444oXxQykKVd0F559xNByZJx2LmdHM3Rf83KKVb//
0I45frPe/oT6Jbh7TRqTROae61/PVUIABK7ICGuriM7rWCH/bt1XEMmlkWVIRcBq
iSBypR5QH6Jrgre0SAKnzCPHPyK+WbljSu1VWvRbwMlPJ53X13fy0ZJmYBdbddAY
CSUTChlpjH2YszQFI7g5POTLqfDHBvonPueBt4OGDS2PROjrILZUDxsdmqRZTqpx
aqgTPx3470KOCs0RQHVmZ9Ia0wQvc6lG4aK+hpB938g8oi2IHAH0xkVVDMlzoXis
BLfxEbbUerVoTR6ZLXwj4gZiYWobiKz/5JwjADAClWmnWhqvJavyRn4ivyqDgyXS
YovmjQ78GKFY/gFRASNvMKB9N2mqgFaJnT/7tGPDempfrQkPX8kRcebKMhfPuT0D
DKY8TV6USynPOvtmjVQc/Ok0S1YIQ1OYc4bNizhrxUThSd+OtairduZgcEBb88fw
+nRWScVOxdx5gMbtMCoV6fxIkbFC4NM1J965XAPXa+r/Sc9jDWZoDsVKT8UGsfqY
g1jqShSa2By56V9vkcTV7CTT1xxjeF1aFzfFqRiDDiLjsF1NBCAr5ZwlHFQi53x9
Qv0K7xu/KkU9PS/fzw+BDHtOdJvkuuVaKLny3YMLX424cwAueiD4gPklaNw3CAK1
WJDyMkwQky18Q2idxV53TA+S+ZRXmzZOa5izjsoVzgOaXf8CLszVyT4rJszhYDZW
f1junpl3b5pWZL/zFRS5snYcrrrX4SZRIGbOdYr+V69dPJt4hTmkWrM459F8j/iA
JxhVGu1tema2fN1szueLvFZ2PBtBSszfyqpT7Bf5qP1hC9ErS7TLl1hLRhcTrA0Q
rvDXsp6nb9A7IFOBbimugBlW2za9bw6EZpp4k/Mwt+Am8H1NVd1IMweUktBcIu24
Fc6P4LHikqyk0/tA+M5ouj1WPx8/9uG2FL9QyCjyLB64dHBHWExUM+7+xUDqrQe1
av2tb/XUElpH3aZT0nm9/01HWf1FXKNfi7tAqEEm7dtxfzdZ2IvVLr3SGbSCSNCG
PwzDCoSCpTfKm3bDikDQiIp/cQvk1mGMxxO9w2D2LNnudpI1wvqATWQRdLzH4WiI
2D8fzoCiEg/n4nY79WNpNRFh7FBVxU5avTon/lgi4+PfDMUBHmVw5rq3KoeJOvwT
/jHGsRnTiuCJ3HHgdgQOZPa2qpQJ07HdUkIgdYRRArhj+t7n1IS0Vu4KmteovHVk
6c7bU8KeZg+XEavuUAfr07XSVLDWB8QDN5qC7IV6l0MEWwSDxo8G0rfmE51P2n5Z
ITIMKuCPAjmk7x3rzti4QYVQiau43uAypW/USfxKYsYdwB8o4nyn+lfztH0bGs5s
iGO+crktGH4VQ0gffU3tImB5ESc0dP8w4K5e15wRzm4tXFVcC81VOoxCe4RB1bGN
AYqO0JTjpuNGpfIzqwFK0AQxqVcsshtnIjxMSzjMediALV+Wst//zkEyR6OKPTho
K4XZsVcw+HnEteTtVF7SXt0nqB8mzinjO7BfPauCTxGkdqyBR+WRTokuXzicOOWd
MsHZPsjlRpO1tweDzq1VaHobjkQbtnNx/HZP1ZmHOcXQ6Y5BRGifn5IQl3GQkr99
Y0lt+wKV3bqpgHomfwY9RxtKP7lhFcBMJyG6yJSguj48ZD4dCScP1SfepCd+TA/H
hobnZPJKx563tL/mTnA0s7YBebolonFVRoQc9HO0hBskbR0hAIsVl6ltu2GM4WiP
mQ3OvxZg6jYj9vcKFC0DnaC9z/PDrDmDnGzzBwRSZJxm6IostmkEuQQASSKJywo/
cxwrvY++XvBvDryAdNStNx269LL+/TJepnMzRxSfYeR8JeiEUQwrxPCnPW9fQPbS
lzLWJiwJiA0UpfMOHDJYtupEHByzLgIAB+Ge1aveWdVkCp9f7V80rGBj/DyIOJRV
BTAXsG24Dmn5lnidSQRjRcSoOTLdXQzCOZHn2kFWvnrOGaWFsJ1VGNYR2Q1JoG6I
w4lOlFoUUjcPBhLvA0LGDYxROI3Ure1AcCtvIV/N0gvIgMYJVyFOCtZIcMs/d0YT
k6L9o4NeBGzYFJwwj/CEVgTTs85fSggzN/6eFr1ff/+doyiqNrezyq0WROmXOK1w
0GjWtWKUDqvWlV7Jb0DBn8tQjkb7/3FfubZbfxvFkTQZm/lKHFiMEIrLTxvNCPtO
WJ0PQsK9OiD44hlMTPs0JBQm5kHixtXvPrABT7qiNZH2EhIUCUl6CF/KQ8fpJ1mf
WpG+/e86uLRis3M21vO6yNPFfX1PiBY7brx9juSNQalWwFaO4Rt8z2PUvuBJi5um
j2z2Xhat0dv+vdGQu8KDaHXtZwiGpJIciHveCRr1Vz3JkUuR7hmkqaJr4o2xZXeF
6dmO3e9ACr14C79RzFONtUiCzQEo8dw+T1RZ7bUNuEh9zRWfjoOaf2Qmxi5EdjmI
uEN1m0qCjFlLkDc+/QKDEclxoP98m2WbU1q1SuQNzVVyyRFt61vhseEryHHeTbSx
8O3uh21Fpb3xLUpJHIA6Dl/Ab6asdbiivg07q0bHs5KiWKipMSC21YrdCNw9xHjQ
pCpA33/L99buERqrkmpCsDNCKz1S7tA+jH87bE0MdsHhlYFT979A7IRucMoB8M9e
OWwsWvUG7QbYXKKECkjxui2ARHVmupPXOKHcKD0svuJWdtGy3MfyUPAtZMiyX6J5
UepXyXJUiZ0CKtamlLzxXQh1ZA6pXEUiuB40ezIcTX8V2DihXuj02IBpXKXwSj+C
dWYAnNUkMs1rh4xmx6N4pcpUfWkPq1HsiojEE7RnlErwhNPwHuKxbxWXFd9tB02m
usyLtRNFZUUc3gjbQSI++NZfXiIM/Ew9SaTZBAphLDcwLTz+JHk/nPA4IE+ANhFS
kMNue6LfQnak1ZwFGAbVOwFscwfJ9FxI5jvM7bFQDwXciWDpq07FRlaOgCM+0C+n
yS83piJLXlo86Ps9ARnrGYNZ/Oo700TlM9++Zkz7pqClo1VEc1em1WooPDbT9AoO
rPm1z0TpM/DdfBjaa1XawU9q/UHByJSTSFhDbLXXRkSs30XUq3hz2vF8QQEIab5M
JfNYcVUO2yK5N8V3CpSaGEuwHX22ItPM5eRcuw3VTB71b0Nqd1gjom1aJXOkEliH
i1zNxZ2Q1rwvNLjp0TxfzVIjR79z0vptRaYk+q/h4VWYYc89GhAMWWoH4XLaSFdb
LfQSX9zIXJ6F6FEEPqdb7L2NGhSOYAJ23u+TEVvSwxhnhOjs9nOVUkwFRQsErBwo
YHygYdZqX+8jTkXk2/gAiwenrlzW4nvkZD546XeVEV+pYUciJYotlzhMPDxUXKEq
SyyFqzHzxl+184DeIptPqvL38vR3MWIp1f5oTM/gXGkmZxZBOcvTeTAyn3gugSNx
SoJB3CzDtHQX35Ji/je7cBsGPzYACcga0JAwEqNBnrQKDHgiBeYOyfkOpTx8Zugs
eA+JnXjEmS7xurhv866su0KuexeIxImHBKGYsr3MmPYDplG4wCYQbTL1pPe5VcR9
O+Fn4gqBAGuUzY6+fxsOCW1HU4RLUo46U6LO4i2hUtt/JCbQKMJVq1CCQ+6ct6MF
o1YPrfRvzwe13pyrGdDBAalprIzgGWRMuQCZUK/wjEGcpCqmNxFRMnGMjDWDPXDy
OqKCBNiWRT+/799UUPj5Q6NYvlfSyiHAocHtH5UIPvaLGerLIEtmOYVMabxU6e0i
vgy0ftAtKNNJL91MUuCcGLXj+gPJ7oCKroMXB8l0CjsPl58TwBBjYDiyfSLQq9L5
kcXMWX9vTW8LJONDZ5/0nXiGN6Y5uIMmUkTlSox7z2t7/TuPKExy9Obag+lAGRAQ
vrwPnmadjwXVLe3htmCDzQnnsaKjH8yykGvDZYlML0NaUrzICSTmgeL+mdoPcNOx
HrBLd3sx58jW3ItRsyExgjbCkwl6g0r+XPuoZYJuwoSpG6lIkNeDyBFpKchFeUOQ
AQWNqQX915iqUu2IQPLgU099On4emLNuTfv3PgXd2JYv2x1yTofNvcURogShQ+kZ
1peB3Ddd0acPQwON0XQVHLC54361pisiryp1n5IsfJs0JbPTR4IpuvIFGyWBV4Ey
9tSQewnd6xITdKvkcz3zJYu/rByb0hiIGURHCnmvCKXicEFQt6gvVnbH1N/2n9Og
I43o0cz9DZvRSUoKgQ4PXOAPBpRG3aX0MG/aqZ5aCdAauC0bwh7uRm7LEbj/1/vS
nTNB0FTEEFfWheuPkrVFECHZYO4HhibHzspG/cImC4/caRf3fWa/9BErEXzaf1F+
OSr0I0xitLugtWZENqGKJ69bWt8wSgLU83LPVZGoIiyU3PA2GA/oxyZgP+JSnYZY
4qlwziuWeletqt7RrKe3Q3colTK0b7j8D8Sjr/kZhlytIp0VfSx3rBlsAuV8NVKB
P2Yi8bTzpQe077+SBdjF8naKveAsa6V4FshqnyTTUGQ0TRVg/Pwi0EEg4z5ZsCCd
i2K5yUi++pN0gpMy/BZCMAVBfQk+AhXVe5McwKxPsqNeuVSwHjry8dnJHjwTLht0
diYn+dVWg1Qb0jKwl5Z/CUdZnqjvaXzhTQzYBG3FEWO7JdCPumO9nsrO5IfNeI7n
y90dcjIWzGQxo3UwWtMzeRM2UzpNC1/lT8iMPYYyKG0awYj9fiJFB6FWDc1lJEty
4yarMrZNfM6sFoTy8qjP+wIxb2Q10+1ItfFRyILw+rM/4XC86Klg7KDQqtabORPC
iwLUDg8y8JHl/GHNHgWNvA0z7j9qSsVe7JlJUlUqwcs5Wepc66f38PdrvLZ64dqP
FExQPhQ6eh4cijAr/hEIfx+ceImuTKyYajBGyHN2pPy92D4EFd+FsmjdCGO7gZqS
hPeeM1jj+YTu8LqhDyoTo4Y4rVNoARk0Si2DltD1y7SboKrf/9fknW3APY9ccGnG
B+bvj8XVMoocYTgxrxawErP2SfSlpnelp60sTGv7YaXpV3l81MM8f7EjwG/RztA5
4HlUhCrmyWgO2MgDEk/24AUdlYOMMULUCc0MAYKAXSbAmpz/MAHsTxf5/XapsGNR
mdJKAL6CzPEQ2HxzxVS/mITkLFblM35aQMJzeDbqC1qGw3CdNhUEI5ScLM/gMu8n
nwXEIoc01bXac7Ksnvx1EveNkxk3lN1ZF4oJk5HG59FgkX1+MCcOu+hPx4oczBc0
v4moKd0j4ZFrsdNFybqD3N+oXowK5MGA2+AL8CoYkr0rcXJudpMvReBqYXqWYYhY
0IkSGLC20xtUegkmxzSPnftQa/qqEM2kFmRXCsWL0PxXr2WNLsBmwCr74neloRbv
Vlk6KyFwaEGn7cCDn/OSjYiavmaIfyjgJvgY46xkbjDQ+hIhSLGxVlOCh3vlBzh+
9SegBwDFoYncykuzAhnnDv4uCS1GJVuOcIgKxQooz9r0fD9DlU4mSIitqcxC5vWx
ILlR2A794sxxuwGqnEW1DFqENxE4KVGj4Z7xjAXiUobHDIhNsVezQZYmbXOYFZ2y
JewibVh8WyyMk66E+nZswADHzPdIagDMCGWZqDF90NN9guQGtHz0q/eAveOyTE4G
T5B7VFvj9LOnd/DzXjg7TC6nvFjFQivUzoOOt+ZzhkmklLn6AUXYQHa0w0ewNKJq
qfhcLboy/QRjy89yUYQgJld+am9NrY3cUnMvtC6KeDnvRAMob7dPLSzKncY+Ykte
e/lA8GzZi/w+6xp0073JcihSFjb46hW4cmpa23EoqYD5/d+3Nn6+I46xSpUGyY0a
LTy2Ce0umR9LJ4Gkdka/H29Szk0CYFHID3t+67QlNFyHCBsaIRWPgKJbF2uG2V3b
uVKkgsHwpt9LIzZhKmUipjwWBGDmMmqNXFvwF1c4FO8LScmNMvOJBZBKEhOOn3e1
FjxwRJpNsgddSkYDPJEmRz8PlIBAxbMedBMIrwOo+zX7vHylf+ok1I/ElunhJ2lV
uRqo6Ej6C75toQaGpe40G/DAuhfnV3H7kvPBjzwpDyIkPZ/01RIcN5pwJaVAYC2k
l3BPS7m8EDfcYD47NGPcmLpU3bIhVhwVv5YcWhBeg+RDjWL3pStiWwYL8b1vl8Hs
zAtaAio+R+TcaWERB8RSuM1sGDK8keUL9qV/TK/PwReYUuGi4DTqQcd5SrMGHaXV
WE9whlpdAKhbvGlOP7Nxe7ZuEOmDx9jfK1apu/NVNTnmcdmtt3xZpVd8rNDoJCgt
hUHOuv7WQ+t+EePiIzlI5UisRVUl3W7nJ7AiJx2DvgFwnba/1kxOFBK5ePb1IAod
fsbqc/sf0NPiSDcovRhvthABydKl6zC0+yMLjipyPgTvwdvV8mIlxgpzf7u9BP0p
DSzST1AVovWgExEtTamOybDg/j/ybeRtHWcyBaCSZgYyZRI5Nbe4PEcANIkbVbca
acgrjTnjaeJhSyE6kCaQmjD/y43/kwWaa8t2zEBGxUNZYkVW33R8h1xyeOUewcoR
B8utEJmuQXUAbW3YC9exkPzYYe7ubyFAqe0A4PaolUozzWN9adNehc6m5kMZACtN
tvC2raM25USoQ+Y8bpn1aw6DhC6khHwmRtF55ucaobJ1qELKMjuaQA4zixjQQDYh
ea62NekPZnvTUbnvyv7yD1XH5kkh2PyzpXU7GQ6L/QkItMJjGW6lZqzpVvFb32cq
VRbE6Af89aZ4xT5aSFM7qohKBx7Gd6CN8/1yZIPyEf5aimFYtkybDFdQ/iDlObbY
QwDlhPMkgYj0k2FNmQREW+W0t0PeVhDYhhrkA+3sf68u+8QWOv52iBP+5o4ACTu3
n0s2dRnmVqYjFfWy7qeY9CDrdsfh36AEcI9lgKYVFdePIhAX6VhijTRFSOqFtSbx
mmvX9RbKJLwZToAXMowuRL8S/0Oq1mTeCKNClIwAzI+Icfok1rULP9ikyck43+B0
/CkSh2+reeeOknYBOmGmJUf3xqbl8+lucgOv/YuPVB6Qx4NndBHHBYU5xibZsH4X
iBGoiZkaKO2eAjRHhh9hAato9XSePzI65nAmbbIY3PD0Z10hY2L5k/dO9rL70WRr
2YtpKXRfRWyp4MWmvKYqwcKZBsV//nfM914ONkv4ZEi5LdBGt0oSQHjY6C3zdxE8
NptAuKtwUpCxSIp0xeVDi3UgSlvclNv5p0DbtbaAycQL5sXd8WyapUy6WUesr+L+
PaARUgYWt6tDPZKR3GyHme8ncAIXT8GmaO7lJKCeNAYLC9aqnvOkPdRAoXjIOfyL
4Mmemx9oTvL48kMHwPjw2JaemRxCG9fnz5q3fOuugPAn2AtKlsxWFK11BONLrZiE
gKOvMCZ03OCLiXRtNEaIZ/oaXVEqeFpcleW93VT/fTooUY9MfFKRApt/KXL5OTaX
pSS1AceteiVwddlkqk7IS3f0lrIF7PZgZn3CKxwMQgTYC9uIbmbzgk8YkfIYSl4K
6rEN496bxfxLK+wabg6LxNian/n227JTXxmurKfu9HueEKpjl1Rvtan0axV1VETi
5PT11g1NhooBZTAE+7Q5LlthZ+f5BhkwNGkqgAzNASs9o+sj1TcF3AqaLc9Eusmk
zpKAjacmRoR4g0wpBSB95uWVFXFCsTWRWQQpeSqmFvu+x8XJWJBHHEUVHCBP/rDO
PDLfYrQBUOOpF6F+rennPJfJvH4YrVunHUTFiLt5dqy7tRYPcSCF0atlUkoROSpT
bgVd1bFTIc/jHLqBpy6Y0cXMS6474QoqQXbX3fmzrhOCo8cSVTr14uKNeLmKBGY0
89z3ktvXMfMuRWnCtCAEYM/s7nO/Y5n1MljlX/ROhqsNEnJbny5JQOyd7e03NemM
uZQ7RorPV/s1cWUEzLq0l6DYnW+KtPxy/C+CNfphXldsMKSTY07j3iXO6CGGAkFM
y+3rN4Nhvw25ZwNXE+K+tq2bGBoXUVuVw7OmJGv/gFQcVm53t6u4orUKBUob0+cI
baayzQ2hUVgBoOaNWfaQRZIqKFhC5keqmtPMXNL2w61hQeHijC2L5ULCp9afT21X
/pRMRG6g1+ylORTXbbLUM3j6eWU8Lvalg1iu3lYXF5Lad3sk7YyCtUioB/Xo66ao
sHRIO2cX4WKKGMHJ81dZvMmpw0GYNowKwuA441xbxSM5YYdvFfp2hQL9Nx92ftN/
T+aBDTmr8YRhQyF7jHSv2cAf9Esdkm47wXrJZSPr1MSgi5QZUZPXZo2/skK9YIoR
S50pDGUYFKE8O/PwIFq6kW8DNYUrItMGxmLZxVikJ137KhyvWgw/uJ7Yjtdasljg
LIxahsuHso3VLLpFb/OS/3tPp9LeqFfD48CxjrI81o96utBL6cwYZiLwvYTskgiP
wWe6kYpMImpgBq5BqtRZpgxJP97H+QTT4YhM/RFHPZ/h3tnwyWxwPfwGduVaaMwq
l93VIRaBXLgQoJAHH+93E76OzJ0YiWHK2VD997kd4p9HfNfZQt53D2AwQDi0JVRh
hx5urx2wo7B8ru1q8QFzcWweucjLyHwF8YZQWTVr5JgIhKrvZb7SGRAtj3zqN/w1
J2VWrmBK9LWbKHSQXKJvL5KzpETWvn7UoNEHvgnlL7QdMZwBacxcZLG2/0crsyg0
d0z5udSxaQd8bUQ+I0y55a+z8FS/wuFfPzRAeQbMxbfQEjSQxhK4DZL21iIJCXe0
FxsjCqcMshTjDBumrzsF++BU0uOQ/q6QUx8PhkZ7jmMxT33FWhZCeJmuX/bSgJqg
kjsWeRa+IN0+YO0cQZSZGAB/ZN24Yvomu7RPZI6Ty+Ssnyv2whT4LR4lSdlVU7WJ
+qoXCVsnzhzy0ERnMS3o/SzHOh2qy9lr49W0/x9cnCc9Br3mExOHqLk87L4XQ6Pr
zvMhoChExHooZ4uRb/XOpOHlmaIJyQsCVA7UEQa0m5RFZU/uMI4LDRwlJCxwmxkD
ZWJRTzG7KaLepaIlADPybpgbNPqYcIKRsHXfNXrjMk0isEIYu9rcmyuEAsf7IBEI
LEVsyLqTeHqN03rLuBpvmqZ02m4dOb585EmgvFCmTU7vsE1EGg8y7LHGai5Tll+r
ZubRKjY4eNJHvkH1WJw3x0nKO9osyNjVSDJW1M8tEV/HIEjX+RZeJpi4NPSn3BHh
IYap/K7l/cY3pOq62zWCrl0QPHQFsCGx/2j8hhtN2mEAa/JCvjeJ2DNDnY3OL2r5
5NQxjjhm5qKbjun345OVqIP7CM//LM5YFpeQ4gqrL7GeqMIV4ZSLSDetmLfiWxy6
w/z65XQ8ndk8oriAUY2oSAkaGSmJHFwcg85uNdjhBuoZEi/uE5udR29f43JsR5gS
I4aip+6BnRcNVpimG71yZdltUW/bmysowMz9f2IGvJvm/trSwQK1nGaPRfQfh0no
SLQmI0u12AOj9lKytgL+Htx1/ojOdRDUFBBVhttJiX9GqFC0hi/rSBscziwgy4Rd
yqbzd97QZMbuHQ9OGehMI/dZ3SUiuIHhuehsZcNlhD+q8adv1WFD23/78EdZIvz/
4smZD73gNGDT0cJiQ2cC2w/qOu7B7feIFs5oh1Hzz0NNwOh10YzqiPhajIT1cUQh
Gfh1/bWFtdE8dc+JmkozoaFWoWwefDRBvnzBlsmkuACUTWBzwYqDlr9JI+DHX8uN
t0AzWZO0+nWevhAr4uTXfxSAsdtaVJdDLh3rJJelftrfYvFrOtY5kmq5/RtZ8fes
ctz9+j7LXW08JNnCt7iXsAZnoORNglSszlw+6oBCo3YEOBzJxuwakpTTAYEx2G1t
zSj3G7IVDwh5EJV4CH1V2T9Gs72Cj6YXVvpgAxgRtGrEUKx0PLuXBvjTEFYzZuxg
fhp9Fp+q0xZ9+dkA6L/EmjPHe3a1j1TceSC8KavwH+FHsDLYZcOlJlYeuh65d2Tm
nQvY7d3QLZTtLKenqhhiIGEaBYg6ktx5mLFhZ02x1bD3fL34Vi12GfNBP8BPmINc
Q6xbgLSSO+XAmyxpGIxHK1EIKjMJMkncP7v1gWA7XgGcM3/lI9tG0KZyyl208eXF
9EfQK2u2KLaofB3nujVUByZ/scFNzlz4QWRXp/HvQVFxQGYRLmxBzSY0QR9YVFx4
eZT1H+RuomAGAvASJBlTG0rRR/G5FHvYwfstFQ9sGBoSCj/ITSV2UiMZO0P6bUQ9
tWMqcd02fGUpuuvw3jLfiTRWi2+Q8wp4+kuIhiHp3QvdsK8e4x7WHtuD3a5t2fz/
EnKy/Fc9r6S+I8zZsLiBMIKjlcgRrb2vsGapRpyOfS7owO3eQjB+Wo4v5bnHKC9R
gqh2TWVJACKTKr/afRs0cQOnEPAvxDp4MW/zvc53lExSjvlp23plcllSnDqflhb4
MRIM1OPStsOTjwuP+txiPIw0RjluzF6kEGLENXoxI68pRK2ynftMGU8H9EAARoBC
jYLjwpqANCLMTVu8ZmZT/ZWXqpwwKM5Y7Fi6AS3T0IJJEmkKVWT4IPc3GZmcs5qT
Mbz/PTWoCPq9/19I9lav3JwnyTzkNtv7qXl698UC7aaPLtEeUCVXbKMwCgebjOPR
7fAsB07Nmv2yl98YWpAZew1G5L0C4VBY6/ECwcLSScMATsLuE/88jYz1Oz7xHeiv
IiQtx60EbOHJ/zPfsuJKaTYIU1wT6LxN6jm09BP7RFwKMxRHyOFYSGapGnKqy7Sn
XGopJX3RRWdQ395TcLHQPQkH4oCnupwfK3vcvhRmjLv9Qf+g3uem87ZVyWmN+5v8
dEmSHlN8JJOZAJ7sUm0D9IgPOdr/m4brxf70rGmAgDsO26974tznI10LkJyVvb3i
DoCEvbJAPVxe5BmGLdGsIEAm5E1WcKTeeLyWloAPQDj9vQZFx0dx/ttugcSGVBJc
SO0DpI73H+m1xs9hbcG7xOwWwkOAjZ+wzQqWtUGBF55NdNDDYzcx/CjS0vv0Qczg
RfaEFYdhSOCdyHy1GFXqa7SoOpbSJLx94TfmclQGxkUOEgsQ9T98qYOV9v7uRNze
qyrfhELkLVL/jUR3X5duCVdcXu6sm5LYQfZC8LPQ/6MT/AXtD/eQqyDMpK65+61O
/erTISAZibVB4RvpqzVUhfoh1FzmL5GdRnCVwQ3v5drBNtMV6QixSML2/bpucub6
m0OEDl7oB7LM4PzNZztGTSnCsFHvQC73Qm5v8wIBxsxswCNMIvzmGdY8qD2DP7BK
OBKbbts9caefGjCze4Wwn7bke8wFZ7sIdmneBsOyuPBiAyAUymjvbKhCZ+7WqQth
hyl1aKTlh0K9aL+WTkiNXdJsgAbTd8DKhK+4YLJU8Voi8Pcd+ynl89vKdGG/QPm9
NCDbOdT3iZeSg9oIRCMWEslliRnBnvpmvQYeZfcFBjxQdn54XIWyBFl/AEferCmi
hgX3yWny9J/kcnt9uNIcR0AmjwINhZb+NwVOs2Pz1S1QUhW0+Nqpitd5ONVRSFOT
zquq4Fcbw7Z8ZNWxRmrYnkzQaP3ecNg7CxDKC8TUxjKlAYewsXT4Ox8QQOlSnWuK
Jp+l4Of3nspG1G91VOC/rryMgL9hXTW8ObeXHZ/C/J+o5Ey2n9gyD6kndZfH+N4D
WJ3YeKAVACqx3ij6WoMhEVY11SNcA00jej4MuZOjhF6EorVxGRVq8obQN8Nf4s+a
FCyq9FVNKcLH97/PGLtghl7EhKnYmxvmJoKz4tPjbQIB0aFpMRkz0HcjMavZJQXW
mfJ1LgCvAlE/jNm5CO71wsZGmtw+0JJ7ilZF5qi+ezetShwCEh6OVezmaj73LByZ
b3nAXW279U6nFMfYQARtV2222LRHo87g5XBE3zQGkxgTFw8gJnPHgaugJYquekeS
3BAwZtACNF1a2rksDfYEwVyKCoidPj8+HV4nsQkNZGmPbBKbQmqPtm2au/Bucp1u
mC1Ra5neAbwtMmZBIyTHMWFxHNp3OTa3j9fvwJtSA4Fiz4Vy+sIJ54Rt3JxHatq5
Sl1ktPXtXKvADwzP3maYWXoTbpW1cS3104lw1885swm2BdVhtt5RtqZmxL9xq+4V
qk03yMwECLffm95iCDsm8T8nACaQHhKzR308k279/C3ZSJgqXKmEFgyHlIQkf7Ji
iU5YjEFyqAiH6nOq5a/FsKmdBWYV8Adq40GRu8+12LAkVezMPrLthjLQL0lQI2Ad
TGERxPFBL05oegu+rv/hP3OS+euHZHMOMLJeNU2rg6IKhJRj9245eF9kpYLTcNbS
Fkvw3W6MAtkj40lzI42AgpGRvgxzY+M+pGiaf5ies+V1XQz9+9WzfbHOFaV27JT0
0vZLEBiz6+xvl2tnTh8BJ20b9mUHclyINxk3mI7NTtOkOWDD62+n27ztJGyPd8Nk
SYZlGKyTyyn/dBlep4sv2fiVyHWlKmns45plm4QR+0lbnNWEzvC90wQQ4KhZpCO/
lg+vP7FFBiI7UcqQSWM3JM9caWeNRnHyWGdIPyAWIz3nVhUQPD+O5cHHj4XU3skO
MtaUby7N03oCshTKKuZsbhxaPdU5JXM3Y4rzE9iJ58eV4itzLs3A1OLWYfb7XaT1
4/r4toKYH0ESnVWUaWnwyxBEinwMkYgNeJyqs1xInPy5K/qQ7E9vsUEXelAj8W39
F80vnYwfQCO9JMA1r8Axn3az0nCzI78jtXUAtfsZVBX3emQaUYthx2uTdTpvDsTV
KeP9OvgFjXV5PND4REzrTPzX3KJAHsVLKxNLMTO0HhhHAg9SXyC1VPsQjbU4foba
HvTwGvj/5Mffh0Uo6fkER2R09VLP/wyqBpgq8ffSgbXzGUgjcOL/9Lh4NYII+ZRk
+PLyoO1SpPpFT/rv+4h3+4k4TV3+fZDDYyzo5qtUCjY8Nsu7PV/zqHyiRWEdgjly
JmVU+tUWrmPlmUgkQ2eNi6nWgpuorkdPEcVUaI3SK+ORqgdWwJ49yj025aowxSvv
pbi1VCnoZJXrbFAJXO13/norOQAIHFAz8xMkvCyPaphmN5a7HHYkzmbYHjTG8BQt
FN+gfc1/77IP2TZEW+tNIng1rBNREkVJ60Zn15hZsHaxy0dmJTWewl2la8bI1lE0
3f8UnrNrEfFTMYQxUBtFcsUAYaIqY6jkwppJWCkcTF9a9U6LhTlGDVR83OSFMUxl
AJw5yXYQIM4LtlxUTayL6PbyHvRqJkEz6X1dz8nEfDi3MIP26Si6AgiAta9D/DzD
n8n6ZI5zkyyfeMRqx/EqFFe1a47IivX31Qg5Z9mS6kksljOa0s/6eo1HfAG/8Glj
GWfEsOgBMVtXfvBHjaaB+SleWThEZx5wCdnaUhSP8fCPPWLE/OtUlmm1BfSmUuR2
xZSbUUAxRf2bDlOgP+l5yWwMT/jgE9X3OgZIFQdJKWt2YXH2o3L/VPiBVeYv3Sye
+zFUWddJj9AIR+DDcMT9++pHT0zBFcMvw5cBG9PXIHT/pxZuOEZTVwQZxiNYxxOA
iHAjvArB3YdAbOsxzyUoWx4Ua3WXtG0/gkz0Xq+o4BN2azTm8frY4fvvMv+AOVrH
yLMmGQo1+R4DUnjBXtLbKaeirP2cV1vchIhMY7wSI3jS0XykF/ocWy+eqfyy7XXO
uf63myY/ZIXMW+3tyiUB1dW65cn/5CNuWXZVqL/HYpYgtdpkMvTm1BDS0HaXo5OX
sSsckiwTlB6E0IuHeV/slTGWWdpTMx6QLlJhjQ5JeWufOOwol3+3YoK45Ct2A4EC
zp0EG0dtBi96yTnjZBNu1X+b0AhNV+lvgRPhDO0dDccy3G+qAqU7VJZzexZrGP11
PgyZkKHRQj88vrA6/5zTeQzcS68cd9edh03MqKkausumKcdEj7uuOa7krhxHuIj1
f8hfqAe1GhHNASV4x4iKerkIuzynB9rHKDrHUXSI2eFzM3vP9JCciWMRqz/o1Azq
4GA277clMnxhPSl+H/TUL0vWf2zlyI/HqbdRIgp3Cuoe/CzKHE5ljm5CzEFSNW9R
uN/cCzABMuT7kZ4JLIpyB1IST0MvAz5hjILbsZzwA+b1OZKI0GgbDpXOcYaTiZRP
X2oeTfkdzmvbCyGHj9UNix1TOOfrhB2E7ElSuN7AItvChkmYcU7DGzfAhG7fJi3p
mPtfiBSnYGyvhE6d7h+DzhzgvMZga6MXyEIgfaa/k7iIgNPRcBb9IGOnHdGYRZxW
XmLCJ8v7v7io6ThG3KMeT5o6sX5yARlv8l3d0y5CFn9kPScPFCpA83VwZkXZx8j3
xGE/He533dxF4+OQnmLIdKETdlZPUHj7WUCQ6OUf3vU+Ht1eoMs0vDMaCYq6rIAc
Bnze66jpNVWPrOKGslknGk3M8yPG+OKY2WkBo8mZHbEHSBgAexICy2jtwlO9KguO
r15vgMXi4+j8hE1+kGDJlIj88Fs0zCp2oYL8fZIsRn2tULG0HicrV5SJWw+ktmNR
rLaFncs14XYJy9/NJ0oasrTizONUsJIGZJCegSeKGCgCnF9sAFiSIVnTcibddxsp
vaPiqZI16zgQbkG2ljNy1AvFwdIG8+dZJN9YNKOBK4kmZMI0M2v7r2q7h5oY2TRR
Me+YH4fY2mcuFjL0AEe2WD7++NFMm2LR+PJrLT4SP8Y59v43pm+r4ALstBY9m8iX
wDfkpPF+Iq6WwNKFmeWhgbdptySBilpj6kBPMeasqwjaj5E1dKr7WCXVSvkqR4jn
3ZaV3rXfJmbLh6QRNlLgQUwtfREnoXJnI4Pbj8HABW/k8so+pgNkDbIZiidohntj
9ShNmxmDL7oYczl0Xubp4HasShCw0RZIzPPTRxT7chcKRccQdwACtzB5zx0bWzaJ
3EeI9vEOWx2tBLzN/boWYGJsbybcHUCJvgi5UlhLteXmkchdfc514ZDN6/fZ0HP7
bw2lhdfsIm6kqC0RTlcNA5x1hPuOksW/iV6RnV/PSWIu91hKs3z187sfNAOfqZnG
PPQ8ljqF437LMbSZ8mvoxzD7TLQ3VbAKbfAoAhRDHywyv+TfO1ljvJIq8Hf4VmDR
behMg3pYxOkpE/dhRi0Gp7UNz1Hzp36e+YkCHF+fSFtbmqI76OQeNbN3Av4SLV8t
b2GgYtamZe9k3Ohsf6l3aBrDv/0gdYFlixxRhRzjpRd1jNYWH4QgriQY3+NT9Zn1
FF5xXaJ6X6dlP1l7qhFYgxZuSZ3mOV4FRV8JQDu3dJ4tF2SeWSTVibERTuFqxv7F
06M1dkYIZYA0CY/u08bW5xSqKZqw69wSXH3XH+RL1TazNjJuBfQ7VGdGBxMu7fzD
U1dGyJn0u561RRN69Y/2A63dnue/1AHanlVLmi/koz55parjwPHcUQIN800cg52j
JXIJOA9LN6COdiSu0jOuyQVuIOoAOCkW/6JDyeOIPeRRe4V1HmqD7a2MLzvOImRk
BJXKdRF8xDEuhbEmW99aoE1B2Q572jlSX6CFVjj65MNwfBU7jhX3gjSQ4cAkcTkx
zZpReKg1x22XxfpNGw2iFwUDk25sfXwFulaVTjuAobNcKSc2LjYBSvKxinINyurR
qR67sCJurUFwUhEkjNOkE6EBl/z5iex0AOtkTj6AyEVGtFu1+1JwoemCAbOkbBX3
GpDR2EqjSJkY4gnikkhX6oJEusV4NC+IO3PvSKPcIFUWFb16UVmDV1mwMSrCOqZ4
LKuiokMCh+Ko+aB1x4e1Ga/UutNgvttmYYt0FEsvclkK/inPCU8seeJU6mjFSPp8
VaL20GuV0OHJMtC3WXMRwg0DiBRJGavZMeFRd/ABM9zY4ef/eoPJMImNWWZmkBMF
7UGFcrCHX9gzKKSm2RTNGo0BWh6u67URJ9jN/SYzw5ZzMjryzbA+BVJsEyrmgpyh
Xax4NqIq3sYCl3N1hOyuxUEnlK4hq+Xo2FxONP9oI07PM7EoCvVym35DBMcZ4WPH
iRMTc/Ay5kl1krPljgipvwrtsbAT5Y0Po5Ar7PFyR3denxpvam3QyVemP0BjFo8i
MHT9d7n9k5xTqglkWc7AFv+VZ0aRgPjjD4+PSl1sg89J8yxqQeDj+uJzawaMlQfO
59jJaVsqGsjv+oc8BmkWPvu81pODXVjlURwPxEe1RiMQb/G7wM5W8zG6coQLs/5u
PWjK3pDFckwMXgPkStcZ5BY6UdUwjKOc6pqaAphv/svr/PMqR2KXzJoNRMjXf7K/
vrIuXV8Ip2FmR+D3naYvkjK+ZGU610pS7d/M6zVgDYHP4eoPqjZJqBDq6iqoQCKY
D91gV1L0yQn1n5Sh8+4wpqxlGZm5WxKJcsG4Gv2ZUDEloPBQL/eZzCALNW8xEUw+
/1qxhexfiZAi9j5yh6EP948yIfFs20JmFJd0mw6VrNPm9bDPMB0/vaHMCmEU92hm
rFLdAXo0rtK7/ZUXkVLhDOmQnLb/pXCmYojwy2Th9+FmkOMyp4WtExif++PHYWRN
9CatjcHx6MdnIjaJgFAF8SuBgbRTO6F27f/e6rRpT73Orshs659Ak7DmZsAmkKH/
jj1EWWa4OYYT67sBvnRTzwef6Hqt6zjVYeRsfTxwkg6DSG6BmjUGC3tvU/elUHSh
Hapz2LCiEAwjjv0NE7UUUq8yxcZdP0L2sBHUtQMX7M3iFV+7/OO8BqZatPtW3/Jd
D5topOCIooiK7FsvuxH11HleJ3eSwpY205aEAgBdkppR48hPBR6MlPYH5e1F0eJj
IqDFENiulHQ7naX+DQVNW03Ika0ofVhVTdKV76brhvGFLIS1UZETNx8ekKF7uvG/
7zxVwQaN7XHG19qdByMjkmfqxlt7oote4WQmAgraez/kjIbmcD4Gp1BAS/OqxnXQ
ml7zJGxLeHf2uh16UeGeeJjAoUes3W6hXfNPh6foeacU97FR5/skfq73S71tH6Or
LLSnOSBk/JWxhEsiyPhep6HvQuBkSgX3tva8A58k0i6cVRyYSjWkNXJW8Xlnizdc
hEoxx9z0QXc7rUUU4Vde/5OY7Y+wg/SzWoMVdaEllN6tE9q23CYTeQWGtsDZC/FA
zswGk1xRi0ctUCsRcn/pbd1F9imuD6AQZDsIPiWeWq849p5H3+PSijDbNBgcrqDw
a7sapgyhzOLFrN8Yy2eETZl+BheMywhZDj6B2JNAsIqm8XQJYhTclEtRNhZDWMJI
BvhoBfTEei0AIcTnNsqrKGT4hvcgtX/L9AjotcHH2SuAxCfbQ6ms9chSp96FhBR7
uyfCT/tKiaNolbfNJ+i9ugATfZS2uHwVr110mmssPRC/pFeE1OPRL8sKUX2ktdUV
dBZW+G9PEfnbMjmn1xbb2dH6wLfLtksBqcSRVJdoqJOdI5VGwR6X3zLqwVs0Iwf+
URvnDDep0SIL35Z20GbfK46I9vtL30T9A7h6GULrzeg3Lm1MBzSIa/C58jUEOR0u
V2isGuYalW7rbO1gsHg92PWfs6ifjUATg5obh6McWjmmK1kTi1cV4cf3TIa7TS28
DcsXbE+9/uK6h9fjbhqdXPJaM9uLJZKbpZ5NM5dRLvjCx9TH43VjpGAp7eW2o/gx
lgGu9rMSsMelx4ZRojSGaIQoN0M9Na5O5Fk4WqjA8Ku//MIl4w7ZMaxfClOvnUsu
B/InJK1MZEAwPc10tla7QKTR9VGa/ZOExahYE8KPBpQlsirZ2lg193xoyvjtZ8Hq
7Rgian9m99EJ1FBuKEsJFlovL7B0vkRX66zgvE3KIjspqA4doIongq5kTtaS6jXy
T4HbN7sKqpCGOuIBWCHuNw9Upa4B/FOS921fd5TPapITQ2LPcj0+KVSQnHfGDz2t
m41vv/XrmJnto06IfmIcEc7VMAZfjyi2OmNEUq0mikFG8EQ+DTWcGMMN4XfaBBji
Fnh8VDxlBT64gPF3GmbOwqMvgAaH3CLtVDXySEARLxbpRVK/efxLy7QQErF8Ax+3
ZblgldZDhA9Z725g4Zt9OO5Ry/wVQQK5F7mho1+KZU1TSUnCL9HpHdMXmla+NtOn
7NAhzg0uFJv94UtNwByTbm2u/zDgPnBM+Ha6UcpV8kBvAHuyGsW9kKI6XgikX4QI
ks5n1XgOZsUuQ8eJzj7TeDZyud05sdjSCZDHfD5TWQxKHdxhRQYwnmi/nta3nsRp
2NWGxr1EdY96eUXId9TpNE1zj9LNjirx5EH+ajt3eEnzOlzo75xgEiiY0tZTcG8p
uOWs7xe3GLPsCZ+kLwOpqiI5Ksfk6q6gIbToPMboga7wlfnV/sLPHBMAhlBb3nQk
vt4GGGWXOWsYkW5Ur9ApmNa96C3Kcjh+22eoDK/m5718QL2F6GeJ1vtRUg5Q7z1b
gBGrXpZmY5bgh++CQz4ELZxT0ssUohNuyW0e1C0avQp/IrShwfTaqxI+qsNWePgU
9pokCOkKZqZytLvycBEzQ8Sq1ITmN6RLWjx9vygfYxifkACYthdrAeAqbF9/QZoJ
yyxHINqQX2wbYr/vO8ZbuH9mpJiRKZzSa/T4zzSr/QbMSyzQngdQpUz6BllUgjUz
hh2k9XOmY8lsn39oZtsBnQLn/bjXFLmiG3QZXKbvaBd1EGUIx2Es6zBeYFpTyw01
AaG9W2pAw99r3MN6OAFZEZJT8J+K/dPiImnJe/LUrkeGv5ACOiJ9XwLbCWJLfhwY
Lkb0HXN15kRAiJWrNcf/DXetkwTIS0WGrIEJ1okL6AGEPUC7Kc7hEPbyPU3gc23V
5sMGIdgMD6JOYHlRHxTYvcWxY4tNN1Dsl00/QxFq1HJEuEPL5RhFcYHxARs4DNyV
chv9F12W8FEwSA8t4Iq9KUYgG6TXTVibwJCNUwTuTwgyR4wzA77Yce/qR7qXQo9E
iyUMwEa9FvE4VOxwPbbtvFADUUwebzwVwMLBqTH4X5uj5cMxEKC7PGhKRzX7Y9gY
GaSV26bsmm8zLjADITdlE10uRi4H+9h/+/ngzEBgvJvYHqzrbo3/ZLQDoOnpdPaL
0jFLVDsoh/Mg+vvxsvKzrQCWgRozZCHR25cdjTUc88Lhb/NcszEYcBawKOuSvf3+
L9K+5jjz55TlI+Thfi+rf1BGjJAtdKY3UjiuL/RijxupLR+gwO7Pidr9iMHUAig1
aY3KnlrPdIi+xufn0mu4yWYp0S4OQ47bj7hANLUmF1Mbq2nE/go6EV93Q5ARFFAk
tHchWpeUwyKO72Fho+qYLYXLu6JHsVPh01eRmjyCexaRsTNxk5xVqFWERlE/1BxT
SGqXFABLQdTZiEE8p4zjw/IHUWfUW1h3V6z4/knar8sIRVeBpoggEYrk33ie4GbR
a8LV83y/cJfS2vCk8zE0VXlpJrXnVOGz/k/ZFmshU6H1Mk9xF8kcBsg5wXQHM2uo
wnLhrr6wAi/MPyAOIeDKWc5UEBDA5BQJSztOqn1PrjzbDBbXTVXiZxXNKe35eJRn
H+r8KPh/wRbvENCpJUuEkRqHjTFY9U0qzZLJKA2A8isokRrPE0OnD4XLZ3EIyAxM
EupY6WZnwruf06Bd0gME6VSz5lr50SJq7C5mI/+b1IfkjpiNSHaBY/fGSMQxkF3t
1+ko6AArtf9lwneh9t643gJKsgu7T45h+qRss0u7Tz40Qz2JZtjVn6eOuQNDejnU
/8o41uCOjSnKhbBB0M8Pks2L0GXL7nYX2Ffk1m04+bD6k0d84qPNlmpFOqDo25zP
1jqXa8NHyYLTwJfVwRf0WyRxfFIHV6ksp5kDTNfqVp735CEG8KLM2hMShOtB5BQ9
EU0uTQqPrMdjZCpNcVRRQTxCzj8TkzAZl9/wzTvnLEPOZh9dfzjn6T8qsuFNRFRb
GdLRnPRDw2DImyU5yKMzxZHXiVBAsUfrl9ssI0G0OLOe4DtuAycqbaLk4l4AWwm9
3cs/Cv87wTKWplENv/HGy0gzUdCwS2+Gv96Uw0PEMqDuws6AL6YEcVaJL4J1HEJ9
Lo5x/K5yyHmVlzKY15z3g1oRgxZw9uFQhkc4a60lH415ZkIToD22E4gbQU2CgpXi
qH6h+XCjqt1boOd+xO8sbEEDNZshScBpJUcrXWnhqN6R78ERP5nNc4EDHNefJK0E
RnJ/FBvQLqDWAMWjZG0gmRBEXbsi+7oVX3TKg5+kebhb8lOupXpFoi+oT9bt/Oxa
a9yYGMEJGEY7f/Q3p1lDJ2tK5RSbnfnfnabO23OJn/QXzU+TbVfMzyizHxzLaxaT
hsa9YBNGdMUTnC9jf3T03NuIytEz+AxpW5WhtTd4TKNFNTQHFhHLXjwuEb1Db9FL
MqbcwvDIi78ELsoNuZY4mMY3ie0aw2KAWBzxxL3N/x9/e5gCS10HVtZI9wnRyVrT
SDbOrLuBDxWx2857w/hrrKHDWKj3zaOaESW3q6zeJroxi+oKkLepF13pj8BhAL31
489SK/UUdaK6yqjM8BurFs7hkgBhCC6cN6k/FEAb9Nwkd+xVIpHr0oWk7lMKM45h
p2bPxVgq6x9mkgY//Ex8+F96u+qWjyL8nvfk7VYBha7BoncoJvSIr2LnhgvbbrGe
wpO+sN3b3V0BUYzJ7Y3U1mQ80CpxSg4E0NMOW4o78gqJWDMRydyAfEc5/91L5PAB
9vcycG8VWVIvwDDOOFf3DL/mtmbRnZKHgn7hkQrZi+LKDGSWea6zzOAcXM/aKoRW
Oiv3yn+xOrrwlO7uKDMcs0dlvl5DR+b/Ingl4ySP73iCUyRgmAdwvVaBc1w4DdBJ
EEMin27/vqR73MWXemCopZojJWgNFqI4mZDpSF3b+PMrB711DWf8Qmb68K32mcw+
UUMpluuZuCEyT0Wv4KwsCg2s61SzBThcq9G8NHBMHZ4WS0YWuRO2cGIU96xyqvwl
2HLk+swKMF4FGYw3gwk//8P0q9e7OQOMlqAIIwYm80o87QaeZKmWG3zc5BN3wy8F
mhhg8zLj7RVGyOyMEVQD+V+Tns9207dTitqCRRMOnAfrvzcpf2suCAVaNwhBNydx
TgxnDRp7hvWOJxq2pK1ycaOeXe5GXpSW+yb0BPCmPyFvCYgt68XaRELgdtLxIrnk
uWJt/tSBHBrdfLKhxi/V2XudomBI8Cp+4LnLbg+MfBUVVe6G+3DugTI0L4Gec3zS
Go7o77E7IfWAThH6004s0xvOKgC1D782n1jMCn+uuN3k2RKBp/ex67kRuDYS7rx7
23+SXZeLHhvc/XSEfw/lF0kTAH+HupzLWuh3cF3az0Lf+L95zN2Fp3SYx2VWZvIa
FMP2Fxv7qjOFEPl6it8SxRZofnPtEKKpQsGAaWU8Oz961AI+Z+sRQrFyPx0720e1
t5+7N49azvOwEhIEYmAq1tnAayKtQ2UFpffyIW7DqznRu0/77O98wWr1uZXmSLxj
IFNE62SZV22e6XPMcJFIEVEs+CtXZB7bLX6W20gj3y784m/ZI5dSgdN09HXcq+sv
rul5oC0u7uEvWTQnVar2O5gAlbmPFh1r1f8xfll16RfX/AzuNh0MzQSWXUf2dLxU
d2+I8upsPYrNRs9K9HApcAaLiuMesTddaHdS6mNiT6kkTXQTd/rx7kpgp0gT31bj
Tg4wHYjsgxmx+uXgiA7I7QgKJNjkdwOYsgWDz4KtWhLMrdQh4PmmKPmPU24X21j1
MQDNRsD3yZFVr/HE6Rq7wyqgJIy94jk/5XemXu0fYniV6ff/rn0Moh8KVCVTSHcf
hagwX+S/x3Vz92WAJyfZukJUkRDQMw7s1O/EYWJE7CFQwTESk7l6v6v/WYaq8Fix
flMbqAbm3ovY0ff56pLO8CJcGHeuIWj7VnypfyqM6t9cbVI7zzAivTDSt+yxeP7Y
jkU1g05+OOLwCaDrWcoVwElWdXsf5EUbMph0knPrTeI1JqNAAURpiW6M65d09d5P
UkDdutYzQFwvaxdTvmvhq5VLFrmeAK6WiPlc1Ble1hsmMS/Qxg3OFZiMd3cpl3jl
OFGbxy4FoCu5+mdnrcqO+NRH8PNZOGSeevz9qdIFc1Ugstgydp2GcyiU78NvWG5T
+gLRdLX3NbJDNV9aBfeMUQi0T0dHLz7RI3t8J7GQj4mPGyCNJDQro6KzLxVTlMBZ
wEfHp9vSGtk1pJ6DUjJzuOjRokUZZWY//UHyRFMdxln3zKX00S1od96uKsHi6fC/
q1EzBMJZk4Ubk0vfGO4BedPODwhzEt/kujkZRCbLN1nwJHVjq+PcMxoI8pcM2OFI
VtOnj2pjy3No5JA3tmfnNS972dWULZhEYTGtWvfkkI4CvI4qQOBGGK9zqgaKmIEB
+NhTRHRdRWtqs7x8ieMB/WZELd0TCyShzs+8znfs3MXX/YjoAGgE7JB0XjV+klcs
0U1HpUGEmOsygM7gQ/K9j0eHRi6c/g/h4Fen2THhSA1yMefl4dHNMIJIfRfJxCth
KfkXoEsWX1ftHWTwDkUukLw9W7IdmBQ7PqtkXVUb83fkvgLiKMaPLaZRu6sgryAW
aed8AXjcbFQ5ltxTd3FIoyQvpTYLjVRtLtpAL8b4RU31E+HZmicWtOv8uQl2dRzE
KZotsjQFEe1VoJIhKL/Uc7zokHnLrNzxHEmAr7VUPp6D4OhHt9rtfyFOng9VJJZ9
zsGvpzh99V2PFDsQrjdbNndE3bEZwOLMqR5Enlp300sUtlqFT0QMpNo8xhRw0SBh
I1dIxYwU8BkSPtey0QjkVIP4Nktm1NFqv6iGuxFufmYW7//iYH1AbGHaXteZFXMd
a1FOmFWSGhMKb7blb1uAhzN/cDwquefyP0aDfFCw1McKQZCPqxpmk3jrQKBARSm5
m+bwfdBkjR9sZZNBGvyOf+LYLSZBXqV0RPg1e7RHGF8+qzLlpUCEzOruwwEuNXTX
Va8lHE+5Rn6LbvxEOxp5o7PMPwQMpHVHXa7Tpt48Pm5B8rbo+KeSzPD8DyWAmjxV
/5CNhb+ebzSVxA0WzBU7PdJinSKkCrYbUXZ7oy+CGpKMvh2tQnRiddXuzmCuGzfF
VmsQ4TQQplEVIMwDexg0WyONqyDLqFXV2B9ew8M5bC54VsgIS73f631E1wlec2Wk
lDcicZef646D0XC7VyggMbI+GJaVdF8qz/zDY54QGfqn3qRruCtiYjbBb2Hshq52
h7CLmbR59gjJeknjKBaCN78Ab00j6npQJxL0+gGWHVuocmCZUw/NXb+lBuSuVyBA
TEAyM5N4WlGNzSe2QUMhcl7/gLVdOXG7EPlKyW7xuQ4hKCbP0HDyzQpitQ1D29R/
rAPQlAWr70UbT+bvFShKhHr4yLpXl7mdGAI7Uo+pDINop8+p2QKXR7aTKcVSZYxn
U6e3uaf4cJv8bY/aBHlQSWkAoVXQito8K24RHekE9eFb1JDpapCfgS0DhMjTwCCZ
n4xQzOmjneW77Q3f76BfLVpi2JHsWvKh9wFtCFmJadMngYRC0IwNNE0CSiZblyu6
Exf3+j8vxb2Jruu4HbVUTcmPRpVFu8WMGLaFQbfGcwLzHGV2r2wMZrC8bvEKqP7o
jzZ/p1S8kIOQ1juLMZtmhSRYkcYdnDK5hhJ8pZebxOUBoL3hZzCX5a1pNQeZO6KO
ljstiNMJR5qFKUV8zHWhzm8+vmbQcVw0aHOrtynuhRtrcXlxwUuwt0m3a2Fno84S
9Ds1esncpa2pEHq/bYj9NHSRg7oidf8hr0IAAy7S4WBsgl7bpF8q9JTzmMxQkLrm
W6wYaODcZk0sRz5vsDYLkIERqYnz5XIBf0N+Tx5kkz0g5jkvXSW8LPEyzOKJEccJ
ZBgsJqpUakW42cbe64SnnSASuQXm61eZ8SFuG0MVJ0ZIA75VaJ9T14Wwd/0vTVzd
82CCddRATFlqU1JztpvscMP+HlUzKyStVnpcnSmMyohRnKmkrj9TmTNlVGjo/8Ho
YGBZ+agoCVOZlQnyxLWYflpcg0IFxCBlzWzmSQBvt5lO4cgU8ee7Y8xGTuCBl4fj
jTjSD/O1KV3yfGkT2sYCy65JKQvJTzFdJ7tmh++0KiNRgAvS1asmHyV24UfVWeMn
H8ztH4ndvq8UmYXcO2wcC5MHdPVPMSAHEZKC947bSC09DJhFlvzNWz9WnmL+IoGq
7/DwhKOXvcxyrX+b/E6VzvCEYCLLcsVnmVzrRsn2bp8JkHQfinY9m6c99uBLFkin
OgJwV2pocnn6EUcxDODHTiRqHPxt4pz+ZnFP4lbFb07YqlmsjizVo3jjgRjb66bQ
xA4arJ3masP5QjZ/g9ME+ws2AesC3FaTiN831g+EeRtGuJU0QSkPYiTxoTZi+sMD
+ZRf1dnocf2aMESZdpZfMMEf9FztzijCSICrdiyOm6OYvjaNv5nlOOu4BUOLH7EY
JQunx1hmbOH26L5vNGCTQVJpKQ+vufyr+OFEELIvnxcVnlePl3UC6rwP4q8DjYam
vB1ZZ411vw9GgWnRcTcZ8eUhr27XIMzF8V5AxI4t5IrIQpAthcSM/pmBIHR1N8QF
MpnNpdpf/us+IndboQSn/Msd6QlRfrTP0eRGEWrqdBp8ca1tT9pY8wVQ2d1rIja2
4WDcX9pdEnOUB09oqpPKvD5NzX9woccMtyogDq3uMzV9Eokh2mtM8EaqoU9y58yO
7FX+H1RZapwQ0GBVF2/pDgDkCUTYmF9sTVUq7cKtC8OF403Ync5s7AvYT0A36Ay+
fkE/0xS9WmxIQhQdsx02gANfxkq3ZgN66lZ0AHb3Ks+9lFhRtOVKHSFUTwQqnRGa
y8HGPB9x473sf73Nk82WVOlpFIAyIcdY+mRBJArn7qtzueVrlm+3To8p+sjneNk+
JX7bk8dLdeHMVMh1Yuo2/LyWGBswSb6O+kMmVbW93bvdf3Pqq8tqkKWoMFba7Iw6
/qR4azY+Jmz3V/syeZrdrVC+kFUYkLtIO4SwJfQvVOINpvKlG1TJKOsH1B2M/pTG
4E70Mo09l8C5gN4gsHDBGDBCQlTf779qVC/WAnDCbVapUae7uR9dpISiQSPw+tf8
/PcHuILPz8w7AgcZq7VJx+r8vALKdq/VpqUsizr1daFDhGRYntQN6KEUwQI/Q9cB
7zWY1/Y4vbpHlMFFjQ2Yn9sIPE4TataAf7QytfM3yD/TktWjcUTU6+vO8qGNVQL4
LyLUjBlmy5JFHpIhw/3AMbxT0tuCwP3BfuDedVkJXqzLcKYG5T3AfdQpB1lhPvQ7
M04Qt0FQth9xy7dS80ADiVdzh8NC2LH5YTltz3gciVZgnw0dB2tyPih9Hpfwcz6C
jtYqHIzG/xToDVvyk7oksxziKzp5hXmXFztmfSfDnRXCInlf9KWu2IpaDOoCvu9z
SUr5lOVytveNnmnyXJEyIXOGeXv42z2dDVItFMEKPcVQEvPMEl4aUcTQbzJJp9ES
4jaao3tcF9jubLNoo2/HrOBgQJ9SIdnkKDy9JP/lLNZzlBRFIAKG5sdbMH8KKttP
3GAKYa4rjHt+GwbvlmOoKKE2K+txtOaF9tsg1GrAGfZN/m+sQOmYjlxAVwu7N4zx
euTRrKxK6GJ2Vq60bmQMq630KMFFLhEQmXHQwnTuIF7MzjOrzSSvgQuT70Id6Jci
AJfKdlUcdQ5PAYSo/Z+1Hb/5tRxu1+Usdiy3DdVt8vKe9r3cJ3U0cUYdGEqrytJM
60UADAUJ7M9zQtV+onCa1H7R5tnH6VYpahp/MfJAzHyTuCq3P/+QCUVycIKGiIa/
86vT7TfdQX3qlaTSrJum8iygjm9yknxr4pYh1t62F7eqZsOsB8ydVABuUPAo/Qbd
RM801iqn0T5putDrdWhAySgkcQPrU24MIe7J+EjA5ApR1gas5XnP6Dm/WlPxI3tK
03QBsU7Etn6DLRsVbFx0h43LudlqBY2gad+5/Rjz8vGuMOH45AjfO4WYce8nbfLm
rAaYVf5Im/wXsfH2Og0jB0ClUoBae9sTd8lTAif3iNvbv+i0siucvq7SV3405S4U
kEOE6ZaS+PeUD0XMVgXv8rVQEj/yolt8+phj9BHtny8+fNJb3GEyGIyk+41McacX
4vGKa92v1uoSpVMTBrTTz9q/f1UJ+JhSagQQ85nEZcC5dE3mGBRHA3fdFRlUTTe3
H0G0Pbyb6FnxZ2o/i+y3MDCFqJUtcoRiyRssALTUkQZAKiQVrwchHyc7DDT3g+dI
Igjm9H+1VI1gTJslVc61d+kZNhqrt5wnfT2eVgksGiZSFXsTMql4eP2H3xwUHW/0
NZ7a2fg57JIrwHg/zvk9oFWvgwjUYD8CcG/NhPOh0iYLNFtGhKe6fNO+shQtet1L
+SkrMkMJT73wNmTkrFaandnvAqCbV79350FrbMcZYPEne9S1DNzrZkf+BBut8yGM
HGyzTOsFVvuXKD7ToRO/lct2isDP/rRDa10FWkdpWBuSU87FNWBeNJkozfDx1OlI
yEFUQgJw9HUUFYMvr/XcKzjNBGTPm4Id+lcrWYX8rDZRsqanbh/Yao+sdLWrqgoZ
v2QO72XlcpODyz5coxc9jwWl4Ev9S3Mk4WHNsZFgXnVYW2PgG4eT6a/Pg9PAVgmM
1HH/fi/cc/moMwqzpCp+lIAaIuu1v3cYYXIXUsz9iKhdtt7sjuEdG+fF8KIEA1l/
ZPfjDarivSaL9IjZBWGFwAVJaieLND8u3dakZj1kgv9ySYAXU1owDp+MCh7bdUkS
cEmmg3xY7BxzPV9Ol9ai2DpeJ4xcdRF0QRlEa+qJK2cREiq6IpKpc6afLrU4u+Vp
ZP28si1eoN+OecPYHJP0LrU4sXGUnRAJKnubagKtv7AiVBG2dlAgl6nGOBI8XIvL
iZpMNf3FX6hqaLY/GH0geDB5S13N0TtxzVPDiCrecnd4Ar8uObMTxutr8MBArSYD
csP4uPGhNRoTi8i2ElODdTTBb/Es8upPMsNPaG2W3yczqimBxOQm+1Dt13wtdt2M
IoG56nbW7SrY3IzZQwTb8vyJacYvklWoVZWy6rwC6PSqOeb05PerVQZLdWI1m4dP
OuhLyLIOS0reifaTFKypf4RlB/bgfEpULOMMrZkU+0dF/VFrftbDOZKkptyqxBeq
ZphoXCbIc/Aq+HN7c6KaqRcRbd0mVzB0a85CO25Lw/Nf3zou/v8xJO0rDXh22Kuj
E0jq9DcbnVTp3CTZwmJkfMR0+DY8nvLq7OCzZWdnMuoKSwvrS6iV75QwPSIc4h4c
+VH29n0wKEUpKy+xpyaQ2MYm9CFpH4BvmQBpwIQag75DnA69KkslFC+NvnRvADIL
zxdViwYvDib0IU8j/v5De1cuoK54WvkceMCFe7teAxnuxw1mpUCRe8hiwMjTiQDB
WIUH3pGwuDMtipz6Cenig553zUkRULFOvWzjQNDpTd7Sj1HI2z5QecC3AA5RllUt
0HoxYZ0G1poB7HAjyiOXB7W50reN6oo4l5hoc8rg1k+Vg8cXiVxJWpsShU/cm4Z9
k0TJTZBbyalN1EuZDIb6x1Z3HfPnt9ZkEwI2erBLM5U1mXPzg0R/iy5/RXwjpD9b
Gu6gK98GBUtKqfB3Qkg2raQhBsDL1qrAUTIvC1oXYnvUqXQZEsIzIEPFc0Q4/eyU
q2VNHqYnI0pXHwklBLP9G41wLb2EWH3IlP70ptnfhgEGL2643Qoxe6/BI9mgTs4z
SVXYNatU5CneHeXhe1K0AHwlRhRSJ5/eHCQ0lXChRQS2B9YQs8LOGT9JeN3r3AWO
QypceCP5yqRVHmB4H5F1nCPa269SiwETMjgca6XM4BFGRgIOS/nDWnIl+w/Wa9Ox
dqTNexfTlbxwM+Z659/fL+GJ6ncRQ8l0ycHLtXCoM9tm68YWKucDoBRfDwrYX26O
qa0m9iKjCagQPgHgxoRGRX1eUH1i7uDCP5LaELKhRNpB13rOUHA/VpHSZh4dl5Oa
DRJTvMpYvcX9Z0I0Y1pIMD/hSeB5vcdB6G5AtftXIjy4OtXPzrg78UZ5ubP9E0xo
widBlUJIwj8Og+XEmIlPeMNPjDRUVkI/W04Z8+XKJ+Qs3kJfNHADUo2kgA1F1w6f
9tC9gSgkCDTcO0OstRFLXN1aSdPxscqnAIH/mCQPHFKMa51sZDjnY+m/5l2czPW0
loWuya69P0jG48SnkBbyHywN0nUKEvwggKKaJSUpwaHzIqZKR4O4Wfnrq7q8JAkQ
Q1Q4fc2AQC7v1eYsQ2s3VWS8cls5UVBnRO06akfxwpBhGNWc1BW4WvUW81IXHsMQ
zK5ygqdjVqijYOEgOKsrA2FJzDvdXwIkwlnvbnDNxGhkKSLurgwV7bk8/pOaZ2qX
qbYpfaoRV1sr77PFJOftYEqrP5r5eO7DyfkDp9ru1OHoZk6Cim5tHJb9HL0iCJHa
xeFse9H8s1DC7tbxsJcUDWyYq+zHMW1E4q5fWGszOQYnWuHxSSCFV9XCL+qrZNlO
4WITa5GENcGS23c4Cc+hjlPO4WEWxWUv/O5cPWVWDZzrlkKV7Mo9/s6svlwKIBWo
7V3EsOwFL/h0oYNzj9CICPn/KYrCH+7QSCyN8lH1+QBh4x4dlJRRr7qXAUgvrFUl
KmsKZD0yMEfJU1mI9VUIhYJKtzFbDgQZBaPThLzhxKAHg3vGoGMXtBMdllxQxViI
7klDyD2j1cyATlZwnHELgeT4QAg8KY7MYGxBJYhR70sffcJvfotD+afn4Hv9uvTj
8lQ4HMEV54fYSdGIw2tPCtTpVhA7MH2vPD4QRtLmCShDAQLSiMvoUsCLY94EKJ1G
M/dUntZAbHivAaBK40bxw8N2JzrNJ6UOEhFoSPD95UKX0vHiUQeMUXGAXRcrZUhu
jXQbGnILxfZoj32ca5oMftPBt5cSz5CA6dEdvXVOIXp/RvaB7jm3mMNRe31WKkno
/5V7o+I7z+z3oIfTUfDGkgLuHIQzClTTSPxFBUqwf2AMrNrnR+ULuijoCi07KL8i
Wyqi8LXR/RqSyoeWBt5FIVdK3KuN1a2H38tIXV5h64UWj1Kf82CtanAX7HVd2srV
4KLYbAbR462+OgF4W+UuAt4TPKoqykqfLhGXeGsbPyoVEV7vJPOrOXbxZtOxYd3e
KB75Li/pJ/R9twhIZ5DO0lr2AtRWxHXasysMbYDwarpOZ7uIpnbBK+HS4b3NNtxv
O9syX8Z+r9b/n/PdpshTgbI3aTM9CKruGdz+NFf2yKnqj/sObqPmncI0xKEqCTke
fO0o+JlFytdsmGRT/gqiNBD4ydHSQKiKyYb9iTnQkChMRmRqvu6dp5i2y0IEFWRP
mryaI/nEnh5/p6WtOyjJf/y3v+YfaQPVTL1ox/zZ/QR7JSxjFhCzUmGhXk4JmUej
EEYsimH6WuazZTWF/+R7zzP4t73NyrZRBkBaSG+7oWENPsI431GIkNbvrBPfnnc1
z2F6twU/xIRd7SPOJ+Zdy8O/akLEos7LBd1E8CgaIPIDuRHkO33pk8PJXwq6UmKy
s2onuLTFFoIsFpHdbRSDYbUqfzwrnMDH48H1G3Yw1Dbt96OxE+UPXuf9hayJSeyu
VZruQWaUXvBaF8iuxQjyH0bx5CxocbbLN4js2oxOduKKTSd8Cx9K9Ry64G4HYUky
aPOk0BwjmtGzzyl6ewt5TJKNwF4XSOyP97OF00DNBRA9/pL0jTyWraMzZUKV2StA
5rASZhtHmjjo04lKfrrAdNerkAyn9ADry1kFiqTwn9kmMgCF9JnNoDsSz09GMM9L
KfsiW0i6gh3jUi+J/Qsz4pumW+JtlIQjDvltLvphIfgXczZ0X6BE5O9sZ4izY8Rw
P+aJjQmDcjNH4BN6MAP8thZ0wsWRz95HW+UUKagNZD7mRWyelIkROD5ef3K8ILSA
nyfIookXifA2K0JkLmjG7v7V3abQ51VAlWA7gf+Cfr/xWMCSQx9G0zr8g4NXW94O
IXUMfiD7dKwjsDT6/3lQSE5bmGeILKID29m7s1OxfKpIwjWmFG76CJdP78cKU78l
R5tsuPpPltrG8Mds75OUX9oQo8YOJEnJ+81DV5CvQMj08kGYnH05x2OsDJkgfLYu
tCRL7UEvXlLPKFqzfEK9KGsW8lTU7E/V8ENB4WBvLnTiHxHWqJBXdwqD64Pr/BxS
RElmyyhd5etCnwgKjnJ3Nt170vGVi5FwyKkZysvQf9hD09gKDUYy1lSBVd2/Hfj/
qgpQCuMw5RPN+6ZP5u979FkMrNEy2/kNvm+PLO43ozldR0Ndq8KK31eI6094f5l4
h/Pc2tAWIeQTm7e/hbMDew/h/ScCl9nmSr4ZsFMOYo3SHZld5af3uulw9ljVKYeo
NsM2APH7zKeyWeldFHYbFpfwN4aEu7DqKd2Q8YF05BcPwC5hl24Uw2vsLS9T+7On
5jCCKXV89uGCvYq4xxwMV+A0Yvrpp7DYAoto/YyU4HOZdGgcr17w4dNotnOSruZR
AQvShMEkEDLAc31WxeKbVVwRQCb5W22i1EcAipZUgnJdpPk4HypUXFfyccb19Fs4
6/uEmYj7AK5OZ5CnpSRv50owMuVLCQzqndD+ICTbDwtcGwcBiZ37rTjVc1vbWBg+
k/31fg0RPJkWvkEhxrobr8pknUDsFEJ3YebfkGlXdAl3IDH7dR0R47haWT5M80yy
p2N5DSvgO6mL+ZEc8Zuc+exVG5gkUQLIIGdVC2uNCeMJuEvqsrqcsECpOqgYQ8ND
/qWRwP1MRIvbjHSnJuUI3YkRk48aOSaSJcOoVeGrEpdNJ+Xc47/P2z7d9FmpbUmc
PkzwDhpLix8isTCkk49i6IiLbA4LrB6mLcuavcMoE30DvXJHJQPNOyKx8NC7soKq
OwrkG5iS+GGFs8RpualhxILvtohzm/AryXUHt51YWM9DgB9juSbuXnUpsAbniXWn
h7TV1yWfHYkLv0vtCx+D9ly2xLKGB6OX6L5P9TX3L/2Qg1p/cVMDkRJKtUH9iGud
M6o7TDdMo+YqLQqo8gi7xA+z2QLFbWUwvBtZ4B+aDAM7+/5U8NhBw4crxl1PHDbU
6KWU21FD8TQFzaRHbx8x4dWQbFUiV7dw8ckERjIBPFw2O5ndveVZIjBvjWVUlRAG
Yo9H+K0+72nF3JLWqLoaBNZ2/lK77bxMam5AOkKVeAEPNPmzBIFmZoToDHM2TpFW
E3CSpXz0J4HwZGf36YTEqJybBndMkFPto0QMLtdCx6K/nMky5YVWQezegOenw3fT
asTJPuPIW0hFLB+1pAGRGR0jFhT9T2sPkev8RI0JnimeD2EAZp5zxO89LHvjK7dA
nzvlq4U+D2P1a8f8LQI5VGRoFsEhzM4DqfURn/OhSvWcBRaW1GNgFves+8aXSWvq
xUCVW4QGDtkDHKo1zWmF8ZR0ldekWdjvudZtUL/kR3CoC8KfADGQsNegtUsogbvc
8BiYwJ8QUDvzv4jAWfFnOJV1h4/SALtr/LFLe/JtD6sRQWHI0qjt0LVXbyMVEu/X
eD/D1lwlIQncXlbMYVrBbbRcWmMROowY2U7vV69xYYFW3hFveilTr/jXKktwmXsr
TB+xIXs2T6GyxjozQuNg/3nUbr98/jvOC/xWc1qoxWkEEM8Wn5emoit2cxJ0jGbL
eAQy+ib1llvEJO+0cNxzeEF8llAuZvc0FTlXdlAWlIT22SqVaKGD/Jtt7uYAsM1y
tTR+fNb9k6bsJN2MxsBoMSTXpTQQfs73Mcysw7cgyMt04fnIPJtwEdWyjPi+Zi1K
LFF8X7FE7smSiM1tFgYTu5cVguDZGJ9qVDXU2MAy3givG+FkGNAlfmFBqHJzekk3
SxokjOo7jhCCunAdhZwCxgsim36yPqjTnirlfJd6lKWzWjlPLNwtCQOB0nSRupIO
Jjj7c1DLbyVIrtVv63M00e9ibz78RYklSRAAhHHvPxTJGzXVzgey8+XlZk7T6/dg
ifuTTVkvqjiZybI04o/eJx4NyNkaJRzOR95OpGEpFrZqHpD/e/xH01H1olcortj9
qOsxUy05HXgWjS+7zK5cmAbUZDrTphDMvSLV1dWb17WjtABc0jsVE0cSWQVpv7Qh
aX6YB9WvH7qz1V+FRqklBOtB4BHuZk4t03kp7rZ4HZvjxm2zFFvx5fspmUjaTql3
/3+xVqfK7dWOUdkbS9sf1VpuJgZH/KUViUcZ4otnocXWq/bca4hbvEwie8SFWnKb
B6+yEYaIDk264BjSukES3fuHmj7GhnGZQ9v6SLGSiKNQSvp4LanjPdeQ2rfWl6y7
VuZqYZNr1UOsfB812tmAhf4VIedBexUnu+SFLLWY8FVEt8jdQWab0bKkwT7YX8hT
6FOuVbrb9VIjThxH1HYNLuNuqR324N6+Dpa8B2JzMFQ2FIOAkyeoNf/FHE2OKelx
SmZsZUAnVCZ0Cg4JKqESkLKoiYx6eaTleReKyW8ha9ombCBKBAF/k9HmGGZBXsMT
Vs0GO9F03M9j9nFaNEYyC6V1NxuLIbzHp5CPXnhUhv64bWWpfPm7w9ykrTKJsH5h
RVWvhWMw7vz78eDkRntPksAWIRF+b7oA07zldDW1LO+85kch8xLCpQv94LCUh+TZ
B0PcNAn3M8jRdCSuJ4tpljtOPDS7/GkQ3aHvaGBFmMyq3M9YXkyd4G9fN4V8Cvjh
71Uazgksz68eDmJMPbmZJvc4vgzQvS4pUspOnNxPcBwgN4MkmJ7FHjfzZ647vV94
Cr1YHEoR1rLQMy8J8EsrcEpv75ay0PTZC+ZglrPfYZMe8kinhA51aF9KmPyCYDDH
mBbP+TQk+Y5Ce9lqicJsx0DgijAZH9SJWTsQAmk3Bp9INqJGEXsddbwbT3l0mUlX
BQzToMy77OG1V6jsclMfMaq4x5x1jGTWL6n92/ausFu1FSMK+kdDREEg4ocqHDSY
5KHopPsvH3BzugY9LUGwfaGn0cmhBwYyAwYmS5bZmHI1F8thjVLFiGSvTpJ7AGp6
dyefMksWKO2jvAalPX+WrWNn0NS7qVM8Th5oTXDgiwCLqlTdFCfZsylUspLZtz6f
HtgIeyWPYqjCLAW+bNod2QWVbMBTFrZLnHFG0tPIDNO4YuB3DYrw3sXlii18mUzL
jFUCURZkUlaCCYdiu01kuEKtwe5eOIvv71QWxcvT5S+hR1ybSwxqwn8Ss8E16YXm
7LzSA5PknXgo9AbHbEjIs4EfoqZ5mTkG8jXKhh0efVEZ2PJtsK0OPlviXMYyxAWl
K7kASK6UhcYfLXhIMva90UwdWkceR9wWwlEdBaBL2dNh24q33uVO9KN65S/ERk+X
Pcj1Zcc5XFQkze9ON4NvfNJaVE9HqKpFM2w3Ha0yzLcrkm2CDE3e/H7gGMVhI0Ks
J0TQNkT6M1/WKQg7emxHRN3fwsP63eqb9e3jvgDxlD+d5dv24tEGbV7LOs2vgs5t
VV/enYwy54u82T2TaMb5I53QwL/A6ivi1+wC/P6PhKWLeAOkLxL5S9ziLlsqAcpe
0yzFYSC2nFXrCBDuP7zSw4FTV0VWnZyi2sJHenZ/1k8wP87eP001MLa113rZmYGR
bqiEpa8yksJxdRDThzzrxlJv+WS2PFj/3d4JzpipxDV1+OloaJON1USrICn44x/Q
AzyHmluKMbgU4FQg3mJxeOSv1JdjgbWTYx/LSkzT7ITO+fEOVhCTrpfgeBHFKgqs
8JDXvQ3BdUJO3R+9+ImAWVUA1i5ayLK13ipq6TEzAVv3z4lXzcYEV2qNvBedBwdH
2jGTaO4Ci8oLfaH0d+BU12cWATQAsELIjMRNoNA2WzfiPz7CavIQYXSxLMd0dIW6
Jtr10DxE//7RNjYguslmDEbxm9RqToYB07uaXHdlj6kqsSS5cRxFksQdvY0wpDw6
VMkiGTi4Vi6n+cRyDWdAvmB0Am/ZBIfRo9POcLoDyzaVWGoKlVTne7qRU1KOM6UV
4F+gnQHyQ91ovFHaPdU9pFq0sGm3NJ0WoI599DvkKZ00e3EF5lFS5wU6o+lwrphs
yFQf5BgqTx2BakHW14DR2tMrqAHE0TKnkPFguAK+Go3YgrhlyIpAP1HM9bqe/jfK
RdfvfYGKvtQMRnQo+Huj6UUfxIMjvBVB19np6nne9M0j26VcoHNDBUg9cJMbXpDq
z5SFe1t9OzsgXyCSnoLTa5O8r52ZlBIbVNd+8TstXCQkHfpbHTt8vVOea7GThG6D
GBvRiqxNDzGRel5dJh7mfTnBHvXX53T0C08kWRr2mAaA5zJxm+EMfILwiuQf+uf8
g19MK1Ahpv+lhtQGqh2rzLfiTK9sS4PzJGZ07KG+ElDieiNjM1Z1CqsSAyxqwzCl
c9WjeCjksBAOQyL63TIBjz55YaXQU7yuH1+/9gOQPqZETgCu70o/Peamklm8Gs9G
v+RHqdMzMQ+bX96wLkApAfE39Vcm2y5sZtLvDpduSavyJfD6ZIQMBWFkAHJDoiCk
BWu7P+2VRJ/1T+y1lq8sDMR2dbt5vbuTK2PONUS/uRLWh56SkP79UBrOg78o4M69
dKC3ru7YZ5OGDvGZ1J+epfo1B41RUVnpA+kRYcTg7QVlD/UbLcof2UN5vMQku9Fu
SNUV7pi3hRbmQroUy99igvJVhpxACXe0820haDRyHHrYCKn33nvO9bhx7si/A9Bu
Nmh9/DN09qwPBUkkfmCQ4PtjY2ThB6nZO1QRV3XmVfM2NaLIm9cFp8uH8C/uzBxj
amb6szTPJJ0p58X9ObcW6mNnzJkhIQ84wBc6EDiw011BqbRSxL5tbXmrqro3PJQf
EA/Otk4r0HfVNbrDIWr64baEJmNypk0XKQ99svlHM3ZKvVaBihxXIOCSVyvwTfFS
Os5m2qos8IlMgReBP8iamlUdg7FleqZq7GjljBzK8lh75p5LMMxdoUqkjXvplfp5
DWPV6bXE5ZAheV0PMquxEHi7bB8rbswbeLAfy9tnrauTf/pjwUwHSCo/9Yz7e99t
M23gweDc7fm+Xm7KoqYyc5Vx7g+yKwmPctcERIXIMhocbJ+XaNR0AF4/3+L7xBPb
mJZFzGfk7GK9/ld7sTekJShxpkFJThZ3aHjQSLwqs5XniRNfzrjBszo3sHCsggPc
lyq5OuaeixUssatNjtOBH7e+fDg+KPjabNBN50q+hF3Cf9fI39pBrXrM0syE4WMf
1GlG3xGTxmFcdqzm0R/LLbNOilhA+cCEvfhxfsHR8qakDmf1yuKGnEwpnLqzi5sK
Zh0RPbb0L3wBRUJEa5Ps56fMW59zo/I1zfaZVO71t6zN7XVpHLOMhtPpecxAdeVT
iIVjyhYjlcXum7Y4NJct2hsre+OwgH2BixspGw3D/TdrtgP8J3cXlzwFwfwizhoX
h3WNTpk3HbVihWOY1l18GktXfSYPyXlPuWAL+pHLxaXZ3VCZXmBEHr+jPlSJXZS0
0MjqN/eq3rAD06wjdcJ23RlNjWO6tVuCSjtlpdJX7Z78XfG7op8P5QbfF5f4fWY2
4tMCKyagWFx/ALUOHILeeAIB1F5LQtE518m1QK2SH3T3esicvxahaNjSk+vEUB2M
q+/cRDJVTpt/HyTkeUNENXjFsHl4IE/3r7E7fe2Mp64o94FEgFltIj6ClG6vAPyN
nIAX+wmz3Y5eoXnAVD3LbSItyZ/5ncmck6pmfXAdnjwAOikuRNaNOgkgj3igrCZ7
zFo3Nv5c+PtjuSztBcrT/69jCNj64FWsOOITRa9Ko9ibmEq5UCxDXAteqC0Rup+Q
Uff9oDeFP25m+UYbJJIC9+Xgeb70gk9l9PJHeHBb4Evoag+bFxxWqcph9p+I+jJM
gMXPFLEhaFTzw9PdOVt1JRPXFsLwqnz9y0lIOBZEV9Be9MXEIuNpB0VULIp0NuOy
jwQBPVDyBkkKT5uJcNoTZqFQtSJgPfAzcnI+49bpTK6JFfC43W3/r+KPsY1k5rds
5RQMptnZlHkz2/lDfv2rRgYWXxb+xarSCeoqiXfYSfs8MwZS1CBwwKX7/WOWOyg3
ZUMYqyCgpyZLFzmurCblR/ANFsK+14HKugBuJRQQrOBbxABfbZih7BBvSZ4HWrgW
V2VKBgsLtUpYDKMz9Dco5xtzc66ENFuYHPSjT0/36F+j67QAept4GdUyfIl42Pqq
UGu3krhYRa1KHIEKo0PV/L+eXCO/ruYhY8PqBCQwrpdWCKfKIFcFnQT6TsL864VF
tHeOw6mnBST9xDxYNo4r+3wAb0u7wZYyO/U2e4NZKpGazDi09mq49xcu0vTT1n+k
6Y7gW02rsbWmLi41lsdiFPxdrL/dft8D5AkqyaIgfAdXiw0ZFiaBgUM9vLh6EeY1
Ltbw5s2OKZ4g/hHiIk6pv/j5aiL4A+wtUlvKZiZdBdfET2QXpYQ6Uq8oNb2C1tbN
+eBqO/fOHq3V3e55jKh/6Y/DRhGY8hjx129spy1367+gMo7xlCnbo0y4Z4X5PmVf
pxYAiKTJgeHlW783sTih7r00aSQXTRfzLdHdR22fqnYdx8xWA6wcjyyXZunbSaX5
b9veCDZf3ZmjJe7C17Z6nVxGJKqQtjRmspn7CRL4uZzPyoODfmEjLP7U2dNzVy9R
/t2WRsng6Zw3KN0WYUEfEUn3RFVB/4O+9chENRaMlzfnqE4YAk5fAFFNMM+yrNeE
/prMjI+sus8Qer3tOOwGFGRt2pIxedYkTZRkYhunya0miwtgh8Wz6tVjrZe5SvsC
p2Xy0XuiC5NAmEF6PT9gn7jvmvu4/H+LDV72am73ppvINdgopPspHGzXnIQ9Cgag
PopBJ75p244isM01rwkp12CqSXGN/wem6dY5rUEm42DqwOo1eUZvubiv3UvH/mck
BNRFzwjl/jME4B4iDai2Ga+fY6eyefMYyqDZGyqVXHMSqWqKfJbWBFiV8vxIfm/x
sXTNqKxz473/QfXUjV73xNTv4nHFdNEJjxGI7Bn706NbtSCaFrfEPzbofEQke6sA
sOT2zQtKy+VcQYkC1FdQceWNoVE5AWfsAuFb9sHs1i87JXpF3RmB5DmI8TxkpCb1
BwjIAK5SDpTjjbgibg8C/YQnoNdr7eWXA4fQjr7bIwBF19IG7b5XFhLxhqQeN/qc
RZa+2NCDfi0ZsdauqCVd8jJCtZ58utKwrVxgcVsFQpuH9Gi7sd37ZL0kjzo0lz/A
iFqVbkYG+pPFwIynPmDDUdcw2K1Xj14kB9JAChSNe9Rjnh1CXCMFn++OhpHSvDKd
RfIyMs89o/C+YgQJjPOIOBY3Njx7JHIxGk/CmFYHZgT1IIyvcMxXZp5YNut/zWLZ
9fTtBrnTkS59gqXv8V8vQHmDtB6jQfSLOoxzgh1a3DJ/ZIqMe44FQ0chE5gzr5c3
lftTaaQixLl6dzZMq2mqTBrLFe8H3aMAfAFcQNwtyzde73zGVVeSxReFwRmL1Odi
7uzm4XRMszJA460UbwYdOU1rn0jLFhs4U03iTvwPnL+xu/Ub9zF8CL4D2Uq97QZI
7DyayTFiKBzX/ngSfTPE1K43s9I7I8s2viu3DAjoABEECzItBDifXGppFvBPKJEz
yZADuyrLJDfX9uDPHf41XUmx6d+Y3u1UnsnrCylPLXMXfczoILAWe6yY9vn137Qn
5vOQQezCw0Y6LcP4fEik8BYVfJqOayN3ZbRF4WDjLZ1AWpNTOAXlEXMrUrQKlvmE
sqW1pOfsHxaiucnS4i7sRc1/fs4L2vYB+B0qUoiL+zja1GRJBxyxrWi2YjLvR403
A6td5RBKJBQqUGfWQJmslKOg//tNi0YRFoOwJImA0k4LUHz4ZSHvf+dUV+QDCrq0
iYRZmeA2LE1l7a/d0xRhmN7OM8XotyK3EfcBCzzHpQxodv+0Qk/2vfkyByyRu5E9
D7eWqZUSizopSpQTZ6fKHz8YK50vbadAxPAce8kTC5Bh6Qd/z9AMjhfRpDzZ7Anw
HE1DAb9X+cpCE6phBuzBns5FTt4dOXeHrMdQrr00tADutU9GRHdqIbJX7++/fkTG
LM9d64o8bbtEDqORst+rptMxk1l1l3ToBAYww8+AyP9y88LQ71HLW2cIVc+Jrd3c
g6D6BOGlF3cgHb5K/DUtDBue4tXfc2QOMphj7SzLJAphe/f5YiOCkSkdesjWZU+q
VNe2Y+3DogXDJalbRf2TKzu5WxB2uaWnpi7j65JKA0r2taW6WOTbKJ+KTRDVsCxA
BF1OwuA8Wg2k/31kwisfu+806lyAEKiPPC1sx05E+vTOOrJYs/74mGG6dfuCpaIr
UknRNkSW5cUA+//R64tqqNq79A9rNWcxIJfkD+4lWwVoVjz+gN8P3FjYuNmRtOUj
GLu/QDVqF75bOyAP6AlrygtJ1qSgdEx9+jkPhIzOt31M5nEev4n/cJuyKfaYZbDc
IagBQX0ScDBPWi20hsjvQbSzX1A6uPmGGjL6xsvn8H+J/T07EbqB+d0nBDPmsEgS
5Ey7CNO2Z/HlqIKkKwvmJBpj4OpADg2fFps4qIbxpxgvoPWhhhqoA/Q803nQkwV4
+EWa3Dg3bJxR3NzLlVNlHBjJnumQ4qAdCzcmKL3/hsVHBvS0jYN1sOTXC6YOO4q2
rKuXAn3Ktp76g0t20dcqV1KLjW6siEHYC2GfyMReLNz3kDsRRaJtoM26O9Y0XKvq
pPgwz4T4BTa/AUBBzLyfAbgpIJCf2WeEFQD2ZttOrmKfFZ72GAZacP+HKd60Gmgl
hgQDmsazgz9omU7tRTXzOq/+D+wynjllRgHmEe5NHXw9yI6U6Vu+1aTeCk3fBFux
2I5UrrvT2opRN4m/6inYl8zMw0vYzYsV+6nrV4AkltT658Yuv6FywUi4fP5nYFZH
lZ2Q7kHLre2t99a4Y986zSkM8r7x3rs6+stDg1oEVvHcDH6gVBmuzcwa46z5CJaL
v1CkMkBLHJfvFo8XicCMh9t6oivbI8KOUMbTOyhx8gg6co1dPInpIn4ZV8OqGTI2
Sp+jz9q50Vn/dMQ3lq0Y4O3frGhwnPSoF0As71rHCZsodTYFKdx+/peyW9buIxAN
X3O1/TfQ/caI+Dwcf2QlBlY+iV6/r1juNBk65/YM4zCga+5C+Xdh4Bs3W6jJb4S/
TeRJP/Nz4WoJboIIie//63UXcy9g0u4NBvPU7r5BTNTjmSr5EZjZk3Y8nH/Fjbjn
3hLubfPa/+itnZF9lU9S865QkwfCa4i4MzwLkf9CXJpejyACDczIzusqDSbR4yx3
YeO3Nym+Mk6MyKMrjrBwUiiil8ogSnSmNPPgw14U3WeWR36R0TWQUCKmFk6RVQ6j
8NciW25Cc1SjqTQe47h7+y7/1uYy+7+JZT95cBQ9btMApzh76rOGYWUUSah8Roj6
YJ218g6p/A6xsM8ugBhPOroxevuB50uCP4sEnkE1JRxwq0Cem8Pqr146PmN98iLQ
WNa9keFpFEXnaOvx90p6B8GhgkWdcsnEw+OVAKd+/9ZTkFXLEao643b4xfI/sZ3J
9wmmCHn9Gri2I1vm3QMmPyU+d+kjLzFcEhIOQGPqiumYK/GwJTgE8l3u8rdHHSee
K/tPSOUqs6ltn8xVUQliGKtW1KbYjejH1IfyheLFrCN6Fd/k/ZW390S0F3z6AqEi
atwod85cVujaOwiE+ZBQErCLWtUny02Pml62FyHNnxCDLO3dJSGG7FJQcnZjbFIR
tPngZEoiMAXeFmloQqPb4viN8xwA1r9uYfpOTuVTlpZrFsjSoXw8uREuH/54s1Xn
DJt0hU72m4T/rPV1CAritEYcXmEYbADJDeSAgIZ1qoxMhfLmSoNWMOlnVINO4TJG
wBc4l3O3Kdd0TRRAblT3m1LhymVDdPWJ5EZF4YHHqR1j3R+sI4LlWHyS6kAwoJlN
iO+htOe0QaAwvbQov8gmX9hu6nBE1Eb2Tg0UqIZRkMcPNx4tWJ30mVWws3Yh59Tc
U8eOKPx8XtgTxk7ewCyNgZJtHkihxm4FSX8u7ga5zBsy3o3BgtsCuAfm99MZVC30
lhqHXEMCISFK7yuO0TQvIhD2E65kV9g/gIecgEL0VK0XH/dIToTadMCqd7Xc5EGT
cYyAN+ZENlXGK4uMZnsPBTLi9CJPF20bxPNFf6NFbgeblIMZBXgAG4M4BHPWEK0q
v0MMHz5RDmDO5w4DM4aL/7pBW+iqbL9QVIBNWMkKU/oMhWL0qhmC16B0QRK7IS6E
ixk2A1xaYbgKITo5SHtZjVQlCM9ZcuNsxx7ebV5MaLNn2902D8FOiQvRC/TuQCHa
lTohe+cfmTKcZ/ShGymK0XnpD1IYExZYfCka+M4Xvmj8WcZHWXfQKfZlfCh2vJzv
22qEmg2Qi3XJAdar+IqU+0GIKF5g2Rizk+TyNwMAOxDN1SJho2SHcfql+pTpeILT
bTO6/36J+Ligr9pa3wBxjrH1RsJFDgkB5i2dS1fxFHmBQgCl763KnUADmlrM3xts
KX4EN4uKsJxCHwQGr9d+ABWRftGxcwYJnddWnpsBDq7tf9mIyqD5G6YFSRCQJ6lo
/7hC39fjwo7crw72R5KK+WhuFG14s1UO2macaUzT1QSHELSKXVEXNbq40maIRGM4
FcsvNkaZjjcLp2vmKhvmE6YFRPWqdrKmYGrFh8M07nfymMwICkMLgaPWp7e82C/j
ESSXdccffiXLxylAhH5hDmn36gDDLXFtwgEbjx6R+fW6XK8vp0e6FU1mvf18Q+sE
pfhSJ1GGeFexh7dWzt8tCU7cLdj9wFVKjTqpkypBygONpZ464HVt4SsxhPp9mN9o
TK0YohkRpREGPexIiam+Sz5jSQa5ebrL7Zf5gFhJAxs8EUEBDXta9VabTP6ox/2v
DSm/7BqxIuWmxddu5HYPmf0wHUYvTfOx1W2BlH/857Ps/eM6y/LTcloS9e0eh7HQ
i57VbUXSw6E3wTfY6rgj0UM/Co+5EyOhH2Nd2n4656KBRdbRRFQ6JyrQgmlhJTso
PKqQb/bacVnUk32Rboq+3jH6S2Om93FkycTAwF/UOg+AHT1fooM7kcVQ+6enTA/I
8CS0kfArnJqwFcUmVtjZStEZsQyYg/RY1bUV5o4khjElM+3pchRLZYSzUDV7N8Xv
V8MvLPUZXuMYKSAafQqdsZMS10nKn+Xe6sswVc93z38uD5FTh2xVCs3DqQoFg3P1
vvy6UNGYa4MaEwgbChTk0D5r53Mx8rHzgYr4JnLj9v8HsFEag8yvC1lsGzwGJJeI
m/IeTbyLylplLkCW8Yhk+jlGn4XrUmZpltOmZ8Q8ZSd8lCP0uz+tZKGkP4+x19Ht
QHBl4dfjiMZL90sNeW1AkyYA1NhchjP5XUUeePNsh+SZsVVZadV7CWYTII3AGsy+
nrhKqxzYztWdDvnDHm77WeAARorL456OudcKTRowWvfi7EbpwrCpbnlzWnfPtnVS
DHpx8NzrwHFV3Aubz6cf18dlOq5z2Q1EvP+5/Y61So/aF0cxtm7paj2P2RvlwJBb
Jces6I1X2fN5bpvX7omifAy4SOGp72ZzdZ3d3Q8fcFOxP0/UHkHTAuFgydu9ZO/C
yDpAs61wtzgjFHM9xOSM7Syzdg5YxJW8Pdt0XWELrx2LwJdiMtYjxnplDaCnx/mO
luMitZMghsgLe/OPSza8U94QuVIXZFppXyPdZhO885y4eAmNZ5KvTyrwmkpHRz9M
CYa0DpR5mOkaJsQlkjNNn1z9d62JAoclL2l5mDvS1pFAjUvYnnUmY9r2ryUAgsMC
4YYw75DrlFopTX/6cwNzDb6Fv6nplt47SaNbJPN+r38Y4bdN6pIIZ6GQV7GogUbv
JzN7GU1HYHUwex08PixRCXBuz149tkUG6jrn3H41git54sKeNgn+8tjYjtdMp4dZ
vNPYvjM8ZXtKWDpCsLrP8M8Az1xSci4TvSwAPO6WPNPNK01tNd5q67PGeBLaX9Co
222zsPnKpe/KsWKcDoroyybdF43mWBJ6WnyH6ka7kQ/o5a+fKGA9/UW+bcY1ZKB3
MNk0EcD5CcfpBIUbfaT7/Ek/lxsfXo9COuTZhwGL3EdGT0cVVorVPrAOrAy0l0DP
HMjV2RoaCiSNhNrOupBpOKn2qVRiIynf1yEOIdi6NoK+93bQpS4YjRnxpbLyK/XA
vpHJ6cpthWwbJW07jbBoVFbj2VFx/4MrDhBaJ5T0BSj3gI/ipq9TlbWt4YzYzeAy
HicPYcLFyQq9kWywRqT7Olrga19fcXQVwaZQI/tl9ULUnCCBL0Rlee9AGxB/sRQc
OUCGJz2CKd9e6BwMMbMxk/2RiBLxPOQHPQN34yj+lbfWoSLvmwHBL1scNAH16pAm
Cakw/euvX6osB0rP2FyYWpcx7RxTCzXVjEN8FHpZ/ZyaIARfBEaCnj+g2hKo37U2
U5OcDnts8s3uAlOdL8eNVonV70JRvUobn9pIB9qnzoayvbysKpgDyjx1oB7cj5qO
ifkfQO6304SQJTD2r1h4wGRQNR29tZspXfzAvgY00cdXZsICncU6LVn3v7gEiERj
Lv23zdVEKuSieA2Kkfyb0fTspYr+hXYxYybFOSOnGX59Y6nligeuSYtVDDMhDaZJ
JsBArZDlBLUpDJ2XSUXxiCPq5YsYmSCoLKjWqlSFc+UvppXYJWDJZs5sKQL8F2hr
N7k2ijPR6umrQMNFe/tXIxJRHobn59xJ84hP8JVA66ZtmqMV3x0BGNsMYR9gsK7E
RiOw+0+0r1TstmuqkR3kN9X/zk3k8TyR+J1iOzRfxlfbF8PwUNavNrcHN6jQ5oqV
Ip0v+kUEbQVpVTFZ/+9LwDcOvoEGSBzgi8KtdP4skUzmSMVEWEcGVuZ11Q+3h/B0
uIAOKiwJqomm2P2o3nKkZ/TpbBiRFj08WBu9suAr9zYxvKYUvc/+JUn2uX8LsqFb
uuyCY+ZmMKBdSHLCYBwa4udlhCZZBQq1/MFyIK+DBKftnIJ3qSgS7EFfEKYajJLN
EQrhskGcMeiTFaeJ9Ro0NiYdsPyP5gYWEK+hF2dyu1Bk89Xpns9KSlHR1h08RV/z
8VBMhY7qPNLnZ56Aw/25e6Xtw8hiBkaKzFoKEMhl4Q2/S0Lr9klesyohB11dStRC
uwqh9yJ/TTVXlpIo6BohL/UOV9Al2SUHR0ict7dNjrfOdWooB1bzUBN2/YLb1i77
a+a375Ek+JPtZSAk4vpMknt9NB9Qy1FISv2qPZGKAGFAQSEEjzCih6rLZKZXNZzw
81/xU6fASdqmRQh0y8c2b/bkPRck4WNratSoWPuUTH61v7MExqOSypikUfaZafGV
vrW7CAEVLHKG9t5kduueJvIPSgSgtiLV6RaFtY/+UdTUrJKzJu068vo8zuPrFQzv
ITl8FNHGOppIxLpLNlj2Znoj+vLqIaD/ppwkjCS0EtLhG8xeNg7k/HzjN1R8VoPx
5l5QmY+itdGlqGHRxGepxfek5ls1AVVVSsviEzBiNtwQctNwAVrRW76xtXeu8UcH
4Ta2vc7Axl5COdWDufVAFnhW98xqqwPq6OHmpvgMDncMkhvmqBjPi1KL5MZ1Wjdp
thQJIy7VifRAxCh35IvB/HXk1nAyhYwI0/TK2f5kTxJNrNfcKNF2Zcdpn2VdBuA7
EivQUMx0uggk6LYDmjBBVw8qWeYq3axPJBtYg5BHj5TG4L7EBx/wRVePhgBHO06F
uTa7019JAqwVLy2985K5deCR74vWlHk+eW0HGh50VtIHB9NRAVtKrMHjpmbxWizT
Ej0PcAMauf8VekEJ1+WMSEKE7IH9Ysssj0jCpIlMOY3jiXLojv0HbCiVFr/AbrB9
G+t55Ha15WYUAUI7UuMc2DhOauf2Eic5fAPQwo8TbsxjPAKcQtGsRDCJt55Fh2sJ
eze2XWtVuc6RwOjNSlKyi74paMMr3YC1619DQsC9ca14+nYrxhsrR/CqM53WaLkQ
dnwi51igbqpNqUaZKUuuf4V9rApx7eZY1HmG4YYkTK9oXkjogPxbLG7VR6TyOgyF
7LtxBeQ0/1assXH9jtXHIXi8NpkBHW64w1nIn1owx6Ci0HmYrRJbsroWTgL0h8TQ
2pUbXraINPk8ZouWEeZDsKxOHyiSd9EMmCVseQmnmmqK58PDnMRWb/IcLCqmsiza
aFuNyazQGapOUcEugPQM3GkdsfXklmSeFt3qp+oRNi+9w4O7Isdb6G921R1cZZMu
sMd5pIQ4oVl3wMAeWF5DKWWSHz/5AnppbkYQkrayP0YB9gzvMxAVR1dguy7UBNre
TqTWY6V3Ct6N71idCxRcpHHZW/A7IEXFVXduLUN/yA1Vx8dGnxbscwo8yvMFLQCr
GIuxu/TWxL4gsYROzLxjCGY1BIxStycQAbZujUO7OIO6cHTUd66u+Ue49uwqY9a4
V65xiLTRoDWLpOUm7Mt0k3cdoOaKwxXufVo0ja1fqPTdzQQ3I2N2HT1UI/ggRy6u
v4ghb8yYzWumMevyLNp5g44iauuiQx1b+hOhZELUISM8QGd6PeZOL1ha9RK/X8qn
MFnJo+zOgUcTQejhhUcIunU/D0A8w3/Jd20hDlUJqJb4wDNxIxTJx1ujTH39u4+0
DantmHSurdQdH9mFuPGTw+TJsxh2XC9EjAY+9wFsUh09P86RMa11MgK2EzAw07M9
CNmMPmZzb6FG4u7icJMrwF7p82SgTjweoUIlKFBEGshpcMNRQ6Lj58IACKhn2AAB
1PYO0bhkFeuEuolhO96hyddb0wQNjuzUbwW3flpH7gXW0jbcax0mlw6GwTX9VwR/
+qBIBxPvs6Gt2F3R3ORk8vpjC/rL1q7Eb9+thTTNVUT2swU2i1VttRKhEq0ySKwP
7u4HLMjzsx51a7c6oBqjhK2WgZCCQhz0rdXKHrr28gGIb4CCITg4OD97h+jCq0Gg
eiqzZ0x7eqXY2fTDAZYPY9Yg7fRlIEy3d3hkFXMGJTB/kCikmhQxrv1uXnYf74yZ
HcsrTJnS+3tdpdpqzvSYKz9TA3m9hYvvuUkBh9HRWhQTqn4UkWDMd+4AP/dkx5Yq
5EcMv9Hopqxc9OGzDrO6TUIjPzWctfuBwphEHWcL2NkSqp7jmlyQ+fgP5p19/9wt
1t+/ghd+wsnCRwEMSSKTaTR8k2jIWR4UY8uOgN+wsx+GqEuqh/WJVz1IN4XYX97u
o0ITn5zbgQInwsOAWySWLjjYRvhclua/nGEPX/CVJCifh+iJCNb6gm/9j9+/E+86
0KiFj7VMtHQXe588hBeyAWr8XS/7ED4yp4Mo+LU87GSFRnLxuY9q5ADL0FF+83/8
CI0MnbP6e7Y5KHYqfWgNiw838XC5Yk1FTrpOTCWUihsCxRl8jWFp05I5c3dfvN/j
DexZuzlTPvku0uIugXzkeWVrCSE8SglwNn1iSQ7g+1QOtewsSvl287PcWXjLGPDs
ngRLiBJiR2Wp8udkyWieUTsgLcyddseuONaHB0h+lfGqu28FiNKAyHUs18j9jT8o
CVlpZjlOX4AxDLmT8/G/2vhdBtNUtNjUcdX+X2g1xegxP3iwoaptP6gaB1TlngPk
s/nn7+NNtnVTI/m8/VCsLQ3Segj2maVtuS3AIkwfVtTqrC0SEWoFJo/ANkRhPLkc
HYsBKZEqdM8b3tk+nfWAbOgfCc4HwCGP1AjiSghp68fvaqiNDWr9FkaUXkHLozXs
FguqNzOiSXXVmNGZ8Kf+3JY0qp0KXkWh37dNfx3CCtPk9BW9l+IZhaJTcLUG7H5h
Q9bWd+WqHt/BS6FLVIhwXP4Pykk2a/Dq/D266nS4qYuYeD5+La3+RKYxOnA5w81q
EyTGgOjLt2Z+CDrc5uPi7LFRKVndl6rUTAqvG64kLfPf4YShQ6dCPm4lxV63AVkq
icfT4bWr6KwArtykCpAW7sNtrt1EsHAt3B57f/Vu7f+pOdSv4eMw7YLH/O9VqFWW
71WgLOM848ZYWsmaVPtDSm2TTuPOU5pD7eEYNOvGWMH8vB0ORxEoeLRx2Wbm29XC
d0O9LbmDGntpHU7PeK+Zoa4sQAHxgDUEjeDF2D0lUrqS0eBQ1V+HNKGT87c2bWlq
JvbxE34Bq/GVvlnwZifxv6zzycZgbIGA+M3YA/2U1eYh1d8c3vovJOBS8Djh/kEX
YkVsz8iCNODUQpaIxnaIQauO4oRQedjqfP5+ks7ZuFv5qcDPF+KLaxRdGztrBNI4
DqF6V8bOVvTNb0246NCI3MQr5uetu+IaM2rLx/cMZNCWxN9vg6G2mg6H33T6CkFB
EbjrxQCV4QR5XsrVFEYL0So8rWKSCkfDv1QJAD2M5x2oo3OqjKQ8i3qkwXyh5e8F
54v3R3Gi4vl8E28FwdiMwvUBCD9dcfsPkXhJgsn3gwKYw88RYRJ3rA9DUXjpySWq
7SkHAawnrLSYr+dP/0+XVZSQes5Yhpu5GtpIM77XXJ5YjQVStzvlKLlx7UUcowxc
IwCutyvo4eLx04E58T0JUytOE+5k2OxgAy2Xqxt2HjEkkpz+5wd9r2b1ozYkLXgp
jiFGaOgxQOfKteFScTaUR5wwjxxkNkfSsVn3ZjwXiihGXi9Sg8lDjaUS42ZCLvUX
j4gQqimc9Qx26Hdozh/fj+kC5SKwfrCwIbVT4Xk37Dhq2pVUWvIiphCJWfU5X893
+EEKN8bWf0cVqtycGFzC3y5QoQzSCBEgnDTpWIZc5RCDcY5fO+bIdGIo6UigCFDy
gKThrBLzDXw4h3ZC1yFa06C5H5WBqefKjNkRHBU4M5+rjYWsPycKPNXnUoSOcK5r
SHVfUMMoSWCfNVYR0a9/xEb4P2IIpGBE7VkxXoEZ145shwl8H4oyUHFvNzh4ABLw
REiAP2DJ3LkykdMyj6j1qshEKxQH/ONbqfz5fzrGctw1sY6BsB0f/j2cAUO7iBHP
R03iHOjWNd/tNo0kCUuyN8zgRQDOdDc1hnL1rRcNOeiHW9SUR8slZ7VrbcbhOyir
096neD6CbEYKLYXX1qpJ3Qhh9vr8rHCJJYgRHihVf5v66Szh8nsWcgw6fceBeWoy
Zo/4Uxl69fMqi+/F93ZHvrjrk00CepTeDgs59Y69Ts9D9ovnsZPDgfUZ1jaPotrK
reQQcIrS0YMqZFtVPgTN19A66nhM7K6i8RgzGHjXUldSVZnDGoxfVbP/9erx2RTR
mBjWnn7Imvy2rSF9bsUT1rkwYgFsj0JADRfkVLxkvKtwfnhNCNoqQa2yBuX2WW2w
BfzQISEO/O9sEKNT7cUNppJ10SZ6Gv+jNU3do3ZAouo7i0PmoZjjgk7h5FWb8zDW
AHA9CNt6Ow7Jdve38F4NYUzdzo5c/MuSFRMb/XlFkVnS6OG8pw5Bahv5+3eQ0jPW
t1wddyV3YzORNM0QbBUwhZ60zjExcCgtJ1F/yElK6uG8eV5kgwEPBO/ufRUxPeir
3v5MybnAIs2wl2mO/ot9AeMfw0RFK+DsFTdWso3Jbj2n7i2d47psPJsj5K7QVi/m
RsGRAqKTLIXdUhgykky2pq8coP677OEKtxJdD4e9g+zYEhBotQZwhBVfcBN3joSl
XBZ9Ov7yVa2Lg9FI540gMp0+YFGp2GPnXmzNiwryeSuJLzXTtEtyLdfQ7nqjMLwL
AeN+pkXPsqyiIk2cTcmDd5EqXn9qlmkZnwu5Q2ut3mhZeO74SoYDYmxoz56dDyWn
XMbcd0Z7t7nwCEC2W0IL+gueohEY9wlCPmW2R5ArmyGxYQQfKqn1tqB3SfSlrLsN
3gpxj9cpauXJV3SVp/vwwtISA9dGRIiH/RRcTekMB+BOOiJv8wxnO2Z8uTaGPndJ
K7TFidXEe9tuIETO6ho+s8SjK+yMfE/94Ulo7ZpU6CKwOPZC4lxUBDWa8FyU+0q8
82D++1X7idQlhHT2Og4g7E5g/Qtolwjo5dQ/Ii4aldFi8j6OwKBnciTUaAwVzTW0
glTzPvMA6gMfBCPLn24Ztb0rAFQjDSItSpmt11Qeh3ZKnE0Xng+hXZcjZmkexawq
5v0PfXJrlnmrZyAUVGTX4xnVG7k20k3YnD5Ovct4kepqrJ19CoBbxzMG1mo/oViw
xQ7Rlkz4wRO5Ef41I2rREd/I9I/3ggST0i5oAT2uaKJEk8TsY8EyomPIuWyw21bJ
sP7njZ1CJhu2SNYkdQln0j0F8c5es8mQI1wB/YXtv9ufSQ2ByVhUIe/OpGnQPI1n
55s4gtmrNKztGFgikQ0JkEJ65caKpRbRFKu8tdLBpAtIdzmwFBNKx0IzV4WxXc9b
FRd7jIbSjPwSr3LpcbD47XtPp51MjsTYOxe9sjh9M535SDn2XAHV3dVQzUjELOn0
9FNRyRRKLy7AeVmXJHvJB0yAb9RYzdx0n5IziqAV0z4VM5XPNG//lcOlRok+AWRI
MX+/gYT8OCWhEAiKwUfJ6PO9itfGcvH87AGyPFzA9l0pQ8d0kwRChyDwSOBxJr4D
5uPMDCYSCcHpeP0c6DEOuKvYL4wMZ2eVsBC7opbuPCj+Nn2uk92YqPXwATPPNNjF
eqU62EZ5ae+o2m9mvXBtnMU52234C6ysZBOteSUCIEmObItQec0zsucyiJPx/fNs
Bj5CDiCSKaqr9ChHihLmSM6SIxAGyl6MOwFj9B5QNs2hvfzd9fTkU9SAvutmCpk0
ZliUH7NzkAKzfKmOWQGv8vWbpZn2G+l4akSDqUyMF4O6GW+DGO1o806ev4jH3xlk
VO6QylNqun7X6RYPYPyjf8CcHki8725QZLLK88iEbV+wJ6K/+kQCGgDKDVoSw+lT
Stvq5/2Ns9ThQJm5BNvbbCWePuXhiAOjYfrTBHReHX6aSc4VsMbsl+Vhv8bVwvbh
4rYl/UZPFHVuR0pxee1Z3k8T2dB4AQ/uR44Q9SmzBGXTlbaky1LCiGJ51tDPXX0n
isHOId4mN19K0c52KciKLkVTDrrx86ScFpPT2uDtv4oI7HLUnrWRc2IVlStr7mNW
x9yCZsIbu/Y5aVp3P33zWJOrRZNsjVIhkycMdrIpzBiN/ihR+HR74rpGnrqPgth/
ppoCfNSZM0PhzcvlbOUABeJ540im3QklnLXTOCx6yAXaJHFcTcx175DN37K4tkY4
GARFH+Ll1L4pB40w5i6aqRRDj26RTIgSoQWNCvVtOxg3vTsDQMnJtICrigTjK8dP
EbrKKbxtscCWcW3GZEiPOouRPUX1GC3N8Yx9EWHFEoGGXNbLomarb4my3/OnWyOs
fa0X2mui/740mM04UyyxXdowQpyIjlmphMHeUFtAOvD8OtK4BDylNMexHC9/hBYC
7+TPTkXvzCR/IzdcfxaeLlTYyZVmMJQH41rLBs6zPql9G+Vg5BOhzA6r/L8RbaTC
seK2v0DtgXL25EHQCHVgFvVENBZNMo/vsYXreHd4DkwxnBZhAopicui3y/g2Tu0V
gn+NMxnpXjL+WXOWKwZJ51CA01DuQQ4bpPaUMLk8bIgQNguGgMlJSnLaCQ2/HJ6t
J+1M/dt3b3Bes+N9D3lvQt6LK1w1UMcnL13UIihAN+tXaUcXLf06GaehIdZWHh8K
2N24rjy0b6Sj1zPjOnVQRLaAi+oDtMlSMsh+v4NQ//hBb+B3MQMoY3iI+trxsZDJ
W7X3u0tCFHxsl/LaVk9T2Q6V3Hlopq9KzimrpICnF7YieklgS3cHMgp5HCaKbcf4
x5sB5jA/rtUvonn+Mxkq0qEJkHZbSIwLRsj5DbWVybOkErzmMLX3zedk3cQrJvKV
/IvvEYJSTwnW4QHvcD9zRQW4pfvTQCE2iGeB4VNc8X+Pz7xAr3tsbeqjIA8WJSKO
onTvexJEMw7UM/rjOPKGUYKJ9w6y/PCIK5pEJWk4xmUKlCmAtf9icO77OMF6VCNP
/WfcZfIesiFxez6doyEz7uajc6FyJItWmFxbQaOXKrS8RAd/RZC9qX1coH4e0Jbx
BVLblUoLGyrr717BCDrVPRubW6u1ghClRBkrdDNLZyDJd+o+zIrc6QGVnAMKdEet
THq6Aa0L+job2jjLmbqOdB57FkqN74dEFOgl9A+Uwicc4GSVutyB6cuNIDaLSO6H
lzi01sBQJGd0Ert1HpVmrKDzzKpcM4cqvGsXHEDSRdNYQpZuv26oGZgIMOaHimAC
EOqXV1bfGrP4XbLX6oPtNN4Kpe2ojqHTrzTwp8cpUFrq+VrJYfk8qfZtYEyb/uVu
CU4tvLXYLzX3OyIUzT3E2Z5td/WxPR+5fuRHprs8kS8JqIRzat8LJyUlH+CqddSe
njxlT+tpBorgLfWgo+9HXV4BU2c7qOyl68UqCLLEtLnggL9+jrknaLWlrMW0IeZf
+zGD4/cbHnyMpALRvpyLrXpEQI8vHK9dom6sUo02PljzuGmkTJMZiHdey6JOGYlB
MKTqWineelurDc6FFHLBrMevGatDR4ff/Iy29opLVxftKJO8EUUVOb4Qx+qY+KSG
iqcC+kmnV2K5vmDFk2ZCpLwFVuhd9fL27aHLWD0gqdfZkXFqmP9+L84nql1JI9i8
yNWEPt4k9X6Bh8xX+zhiUjUWdkMBsZqYOqi769B6LvhoGgIw2Dhe3OT9XctXVmXV
88LRwScIo9TStUh5xLn2oi588wWOxCyvlB4X56XFrf569SEb9+JyKtywAhPQ1w6J
pnS1b7LLRhWLEEm7c4NAbP/5e+Xlz2lV8MrzF+ieMRhas7G3xlJUJxKGJz+V/ZOm
U8e2wDV3tS1F9Cn+tcUeyzNaC1baOGI4K6IuPYhtC13x6mxEVT03hZSTPmcWG3M0
0gG5JjRqHBu9AOO22bXTaDTZYSkACqiyDTsfQy9vDFHGgAodnmIHuptAxq8E1x53
ccdabItfOnbO03FIGmgQG3sQcYOcdL5jfAuLuumXjyVR0vAjUtzN95NRVK1uPd3V
wrf8k3wf3Rsna1slg+Gy5P1X/FgxeBh4LHKVizvm4yW1O20pCPsEVG124WuxE9ln
G0L/Y4BqPD8nWgW+E5W72C+LwP2DeDOCI8HlJc3wiQVso6C0CurqMPJs7EK3doaZ
W8+QtJ7g4nsC2yIpG7Z33IX7CLdau2VWuJPSgNOh/5056Sv0ZDRojAoVcPgM2zRi
KM2dP04OTU5LBqktkAzEf+ULfVfUESIHAEhMLKfwjoe/rd30chFoAAIXtKuWyClf
ZNjPVwFWW7oSVr5ENz8dEC+QC4fEzOAq5wdquGgY4GoumJsXPvAsxbIRu7qF+RJK
sBLtnJD3jR34aHUB3M5KEtGGhOzoh8qd4ZUAc/AgpCWebn//QFfNAnncX28h0sgk
UDlXYl2NtY4M+IVVsCZIudlq1SW22FcWAPirRfg+eXYpGpXB5dldTAk/SrZJaiaB
Ix0Xl6AI1GxiHTCFtsl7N3ucltvlfRA8B+f3+Ve45hSihek8hf6fd74n1c0TacfJ
551+PT02fHf/auW4LXt7LC2Zv7cSE/JnotXBPb9bEZmL+KcboObHofirY3l62elt
ko73gOUUb0WY/yVp7qkuS0uKXrWVhV5l1gOgX4ZttTgddiQIcFOr7FD72kZeWgh9
WXmsbqgVuBO0tWzgI6wUdLG9+g29S/GqS6Xm6JlxYIxuVMDxT3vaoOy6asnChXwC
GL+VkOnK2IZWudEzYBhhbjQN7cAYjtxcZt2i0ThWXdmFJL5Ec6narE2WrLzELwbb
ofONEoWBMMPVJP8LFTTrgqXInFqjKEsAmqWbAvPCXQXLJHjUwgYW7Bq7RTte8Za9
2fRtrbSts8os6CqkHwUYuV2iyNcWziiXu9iO9m7mIRkuonLx9JpOCMVhhl6f514A
YQLRvlbtRAJAuNSluPXkgGFGPCARjgZBiajuWc1lCQ6i2HYOjstFzfhYe2aJJ2ig
K+GdPRIYQiO/CVtNq39fG6AJ4EHoSVxYLle2NBrgH+HL1sNZxTb5BKLNprrPax+/
2vfZLVkq8YEGNsHl9PhsjUJVztcdkzMnoIIV9flWLyxy9B/H6RHxPEk5WJ1HP48A
SMenq5GppYbpi7xByFbyAwOTWlqBbISfpbZG/wIsaiNbNrg3e7xj6GUsBvxatn7Z
QTHWNYB7Ybqm6/18gPfRQyAGW1vEILGAMrt8iOwnFLoel9Hmk151usl7E7sbMcLn
yAMXPUifsvlIdsgCKBehkx1uI7qoaLFLhHb0Wb9K28SRGA+tShqYAFSnGO/a6jMc
AMeNQUnnHvNb9wrO+uKZspNoW1IQGgMXCF36IfjItBoNTlICtAwqWxt/qEyLjHLA
fSs0NOrVvkVdYsIf+l4uKLogvuB4TMJGYfLTzhySZE3uzkkyGm4G3UAB0PhqPjh0
Uih5msAX5Osh8kHQxdqYRbEzD28F8gc61puSi+HbQgL/oHD2r49qXHZ0gKTzyvVW
5smAt3dKv4O53DDE+KWx8CgcRZlJeXTcdFTjEijiBnTfX1avGoF5XpJ2ZBTZ1caB
3ECeNjpHxgCRMQ7kAOXjBxWv14doTHKyO6rhX7WuCMo+UdDrQbk/Yu9AeGTjfZ4F
icWh3FMxc61EMxkk6JEEeCOBpOpq/LEH55e6nEsR/8c1i+yKS0NCL0XZOlkwGR1Y
aqJk0ZbSZSJ1G9+0MMygzcJtJaN/EKwjPem8IQY+RIAk5FV8hewX++OgKTfolTsM
CZZAsZ9jLjoh6PiyqNLYF/2FdpypCDhsIcvheXEHorTK1BgC0PiU6SIwMrDMq4IN
kj2SqCQqCyFThx7mlT9IivGxb0h5uckKktnXUO8zNPoJbdv7LHeDKFGAPszk1qqs
GCmHKKQdGbKoB0XfSUXlD6yMwig/jfN7irw7Rcb4zRwrm9JeDes/UPma0o2SieKP
kBwZB+Ijck4brz9NBEgf4WJikaVZx4P0VkSy5AiBOL4GDHSQ4klfyjQp1c3uZfPV
OOqK2FMLNhPj77qh4U+FO7z94o/ooGRpb9SNO6jSw1xjLs8mOQBtrwHvRs+XPs+7
YTVUNb3avtm1FgNKORtYbbTquT5/kq3O7lL6d0aXDd/PJwarFcJj5oyxs7O/nhFz
HO/l13MrnuMxhE/JxiOAlMyMU4MaeUK1JG77gbODb+VzifL9TPBU1UuasBCpejxU
e9WF18radKyNhuIgFe0olqTTHmRtLlZkMhf/UzlvirzJVrdwmBSbS7YuLejIRMv4
J73pEaQBQB6fFodZc8k6tMrvy0kAPYBYRLJ6CS/epbdmaBPvNrZ+OC+eGl8a0DFv
OHD+XQoOIIB45z7dUqtlZGYRKmfMjZ8RXtMraMQUWkowkV3fFeK00eBXN+RVI7uK
DX6XSWPkzfUqo/erH91pUZdWGScW9htsqVXaI8iO+lnuN8wze7FpTvumveI+XuOb
7gE7oDl0I09wUp30ve6hn31H0huVeaBtG2nl//uCDL0z5KAXyLqfCn8T+2PZ1w8v
pfjCZhhWYL51Ghi2ozJBvxDeYdykQKgtwe89nuT3JtwYCwwtJyGjLkTJ08I7wa0S
ngZpEmpDGi1WTIkjjAqNlIJeRO8dS2R1eMZ2B2jnlQKxSEKy9GogjpiJmCRpyWEw
jK163C8bChZ8oKEMNe7MgMr3PqWWQeeXWokMogqGKSOwSL70vn8ln/6NTlBt7jum
umRUBd30/W4X/qQPoE3gf6ScU9Cr8XMPR+BUA4hwOUlk79mxMR52Y/IfYg9xGUMN
Wgc7cNYHQpNHsPAaMX8i0We9j1cDQBdP8ojLHuooA78YdQO3gne6fvdXGBUfOuYp
zm5BGwF/O47QplTWpaZJJC5LcpMkMJ2xAzVGqGqvGzAqD+WTKVfLQVLub9mXKEj5
uk1B+g7N4bKJYiWrZHy4XJ+XkrPd2agsOD1ZtSnSJf5JD3pJHPJQQ+hLJI7Nh5Io
UN7o6iQ523UoGAVBmJCTbt8/DDIRR46j9gl0+dC1zo5Dbjkoz8MnhZ/lgAJwyZAR
bEADxAtev+6GKFkPz8Rd4zMrWTj067NJnX8CLMxCbAVouo/6C/uEXMq7/ff+ynjX
mtvWBTy9eWJ1nKzzpgan6N8701sJ1j70HIOuU+bqyK+GiyC0bEYgU54IRZFRPkUn
9tACKOzxqy63E/dTnJA8tGcBqWfsUOdXZepQGuWDMJR89FtpLQxXD5FLsOQRZ4EO
8TecmaRn2tAJSs2V6ZmhGcq1f1FKLmhklOYGetBnhFWYp40wyal6FYeaBzLLx6FN
ZbWoetxLjgGlcAKJ92QRc1rFmjg8qxKqwXQy4LjLHpnN7IXtttXgtIOvl5zWnZPS
0CSvmbNE2vrJ9U/m+O4NnnrCS3ScdmR2reJgN9LOUjDG0rJDu1Djh0sZokc90dY7
VXSXAcxUIp2J5BO/NNw68h2PBN22m3uVHVi1uSwXpb+YAKEtTGv3qLCtAVkpiv/L
C+fMJ/vYPAkP34KVxAohHUYzew2tOt3z26FAw8hRcjSHxvPpicnO0xElfNHxSUwp
d14z9E7LSE5uBOSW2FWosInCSAbsbxzFYefzMnc4Tkzb8eVT7q0hn91bpQS4MfTD
Ybrt9abakci8zwqBfeNlLa+XTvLKFZNiGdn+VLwLcshxg3J9bF+vda6yeuGVhpzb
ijPx1lEIQ0PwjCCKGeIO35gXlML/Txqow4rcjtB2oITFScLl33oYjmu262YLHgI5
vxVkjgKVdzJ+Tgp0MZmuUJxhNKD/liV7qeKpsHwiB3pgm0AZloYW2gFmoytVAj5w
r6QVHhOs0muG9mfARmeT4zzemLhtpK9/4C/OCaA5Szgceol8zLRD6Ddg6lJCh4tm
MxciyEmMTOTHQJIOtAPpnFWoBhXH7zsBOCOd9bEa9jfJXNC0oStWCHpIiqYSisQX
aj6SLK6XBWkkm4DqDhE65uuxL+zBpaCvJcYgHw7W8S8/0cDLNpkj8djgTjZfvhZC
iHBipevUgwYazEXNqC2u21oJO1IgVTdJxXe0F5bIzquN512Q4VI3L0yeHyiSyVdO
yQ05DuUO3Vm2utM1IdxDy5/28BlsJ7qIGbUxkQWf7y568aey5rN4EDZ7OH2UZKCV
EKma7V8b0y0sg9IRfcBLsZVn6R8Z6GEznwbO6Cf633toS/BLbDz63KHTe2EyxCtd
bogD/EAKvzFIHtfw9RYj1104pY0YqVKfoEefLksMN3FcuaiEsChLh0MkRAzo/iNl
E0vD4/LGs4b67muW4O9NIkIM4vzruPnTzCTLkRiCVThDvJ4GsZPXeIlCATSdtY0M
lDhr4MzA2Ama88lztS21qBmGHhPcmkS3+W7puJ1gEd7K8bI8kJuX5hR5x+YMeV+I
VeIIJcnVMahCWm6FV2eT9tB6Nu52YlhvBLf0iUn1HCB6xG06toWdQFiIFsKXECwx
hL4GcGLGyBfS6ifxV4uGe58bZjuq7SnQaO0/WDVrJ/dQRm+tLpWRk777pJZvgixC
bLtnYHxnclCI3z/wnyAHGoYhu2hVmktFJCjZez6SIuWYA5qBvk+FbOSlImped/th
QJF9bSJ6P+3NQ92XzGdT5rlFEhxhASGv1uaNtEElmaP8iGuiBP29WZs7Q8WqQwql
psldYvFQ/OzQcEwrunNHILo90Pg/ZsxsHyQk/v3AzWWqhby/LZl6Vk18+70BbpKA
VzQl/HYvKPMgC/0LuRbAJXfCeSxKXITFu+owvkOKEiBCqVvWXlQVGRoEJmwbS6ml
t4yv4lE6/ZY6hfnNee56SAoWdkPknlxHmiQO5/udsBe/ztVAjWAkazxGL+4VJEir
Ii83JDFpEkRvoR/5+m0P2wGjsb5r2ZuG/ZiP0iZq2J/3HGeCCtVuwuaexyeAuFxz
sDRANCqwB2JvBYhuDsb6sZM/Xa+/+LVFEPTYsd0kyaFAa9z3GK8qysRIMZgmAW/8
ePIXVm9tgajSikbXA+hFyty6XiRzqJFwaRZSL48cVxrWVn4nRD9VrqDT+wk9bmQG
MzPfT0rc04k+18EdHWX0Zg6/f6BFZoDDEZWLSpfBXDxpBoBR4pWr60J6y2aKIEgJ
xNjI1+1UNYrEP4CdEBnKnlDTAqw8QDk0d1B59+qCFXFGfOhyus2Adq+9FTK6e2UY
ZCBEPWniUVmraH3mb5hxYPmC68qrcuciFwRaR/8X6MuTYgtdFrgKEM7jkQKoSOZM
EIQgdGcWsL+5RtBren+wSvYPN6J2jGaFyfGQrTL25cwJm3ibnGbclSc43DDVIfRv
WqceKfg/v0c/imm50Wodg7x3CiQnlGoZ5xRKqcU6s20ZrLOIge8ySFN7NNBWOsN5
XFvDp5Z6aPaCNqvMyXpjI8bKqsYjTO6dOCAAGgwtd7FnDsmHJZfFgfa1N+6FIsUl
aUsaJtnTb1BPd5FP+rrwKfOodaIh3Q4fHHf5tO39YL4cLDB9TrIFC5/xqf2nu4Gz
gy1yXNv6xgodBiHU/qMxLxRQ+LzHC3NZZ17f2D/9FG3/ISJvFd5HcSd3oTFXeEpX
exQovcfRCbd0G6ElMkD7H0fnUepDH60KHiCwqsZiEd2v/L1IgkllLPkbywFiAZEy
hMrCZaEJWovODjN7193J74hWpgiivWjb04+baZJF64PvYci3ClbKB3fQtqBFd6Fd
v8MLWTRFrXv8jeiaWp1FxgtbRKeGdNV39xLZOWQvO9zke3UH1+xjPRtzjNca+wVw
hPjCoyoPmlWX76wuger1Ll5JMRsWrYx+r3oaFG7+Vs8p1FuSJ3dXTGCXspmxmcMW
4igPYhfVDYoJFyS8s1tDqnsoWu6mkLioaTIfwUz+Vv3iKOUtQQBCifH30/rDmV2y
u3k/Z0bs2rKIhU/ZCKq/glayhBC0TTDrgdsi21r2MX/nMJQa+PfOhDh4e/+y0NX2
eY/JyjF1QJG8z3+axfHcpUzRKM79B0fndvAM0xa5e4kJBUDs5pFQrFiLM8MEFAx5
sVJXL+yeh/IEh53a/8axta/cMqfRYLuZWDcKOe2QHkFrRRHfZpHZRm3Pm040geO2
ZnUlwBMnHKNRt30VzF4nJyhE1ijw5PwW1CcvXkS99dS9M6cjidlgD1WuUig/W/jZ
ugJ1kaSc8eEXTrBOuekQEGzjJi5hvVbV3NsSyoWInQr8jbJRSe/R2Hj03GCPz5Q6
+6yZWLY2CZQUVfqxVHvxqh3U1KbZSZNaSvgWxiAlpyoJI56RGS2JA9eUiSuJo2Cy
8p7W8CuHpZbmvF/R+M4aLpM2mFl8bX1a/FMORrq1pUK9XIFQtB4u57NeuD4v8t2x
8hB1V5YP2ahfJMvrZnNhiYLvyvIwSHx6JuoFXXlnl6TdjZd/wnnDZfstqYixh84x
d5p74ATyA8gaPMan5TTqCYNvvWxHvkrCNlhlK4ny2FlFmZkYD0f+f09a+7bBu7EO
R1iOsq1AjzSYSs00HCwFHTBrNrfBIKBi00ngMMCvZBhRRj1T9E96al5cySDfT8qf
lw1X77G9FuGVZ1IqGX3FZHWIATzYZRsLhBnHzU5QzsW5bIh7pBnXACQiY8JBlu0I
QX1O3W2d9MCisamERTw2Q6IkPYF8OcHxFslwfcE1ZGRKUzGhY85JZcdJJrw9wpNh
a5l7HgDHFvwyImIH36qBbJ6QU28lk7fOrCwpHyLNqpbdrZQCTzA+J6kRlj/vx3XG
IAdaxMxExJiVvqBCV9z83BH2htVk4sOoAAdushawJDJl890J2o37WO3W8Yyx8+7k
P4XnMUuJHaXpw/+wOseuiwNAXfJAlqPboojexsBSnGAWKHMy1TbGRu1Ttad70Juc
rlLgyXTo1gAZs1bWHnNlVb2iwki4HrM4h6jUPSmcTtswG70/3J8avMwIsuRRH0iw
Au0GHQwqC9m8l7k/GvAMgdbPHpotYMNqclkKofzXw9wlqI4GLxFjPxzrFd0LTg45
btZyax9qW7URIp4/W5pzwVvo22xzns1VCIj4UN8a2MHKKCg0aRE7st+PB9sO6k5+
hvn4nu22GX/SrxbZDkWRfFjHdUTl8ovLuBFNI2cjWCCTbXQ9a7ykws/NFeEii5l7
uYkD4LyJerZaHIjblxXHU6DzLsgyyjOfdG1MTVPcuSp/Xzth0L8fSHiGYzcSzBBE
L1AB2y5lYIlJeTU5oznB5AzvOTsH0S8lWlkwizzXfy6rZypK7Q7Oa6lEtZZAKSor
cIEwusDjoZMMJGgVlBguwlhCjf48mqzprNWzBuaICy+iJo8jqQYFMQ12818F6x7M
Wa3JbUf9x1uBJ94d1A+UHE/D7LtsESshf2QXPG0TPTpWnCtTTq0n3X0sPXG4p5av
FLGxIdAY6q22Oi7ahDOmT3S4GgubOdTio/xTHZgVkAq0rWK1/Aotg3pVEkL9NFvs
L8JxmG+aTqvnzko9SOf8COcU/FEYVby3iY3MdW40hH4XsSJU2DgxCGmIkRMlQ4ss
+v1C4eCVONuUrYU5NWbDz2HUcF29oVUtH27QnprjTvoY1se3eTm/DK7YXbEzzzjK
KWNjurXhK4Q+n5UIWEJKPmcvsZwh1aotaoxU6Wi39roSu7o17I3sGvxvNSPRMCc8
vOiFwFm7n3GgkcqH4iGTEKtHrxCkmD7kS4vjTL1/1tcnRpLH457HOj4gFIfyyObi
XV3gCFdXgK4/KIXz9S2dFFYJJuUTI/TtT95hvAGYCLZJGUmbCZLMkEUNd9o8HbWN
ubPwV+TJBlDbuMA0HFqUO48HWN2wugYYLJZsMNaBZCvhMX6ySgMf7ZeYGbsSENb2
nkZNGoOreVgPiL9a1WJD4KImGB/jJ6qS5zmYSZ0vdFMnE3LuEryNZ0d9Q6Of72b2
B6hPpoanw/wGVKcXNiIXqphV4NABJxkaTEp6yjreMuCLCnVWJjXApzS5nb4E/yZi
6PBHK39N/d/gPAucpmCA1Q9LuisP9MstOaiyl7R8j7pSleoliCLSHmzdacUJT90N
1AeDi5TJE3rPXO3J+b20yeHBZJKoCOgUV1lBBVCDTK76dmV+IVF5dqG8gVwtq4Ov
FRmjVhpTJNgfutlSbXeWwWn3Gp5frIBW61vgYIa/ogurToThYV/b4skQZ1oafJHu
y+Jwk6fHbpUyHjEIK6chxr7KOoZZIp0fNNSuPK9PyJALXS3D9L5oiMwa6Bnu3alp
JZHgio2jbeu7UxRorsy8fj1JYkf7WI/zddj6sOLgPnYbk0kYiVhOZOa2/oyMQDAT
rQ4oyLntMs50vmP4D+9TGoG3pvE10H3AvHMBkjYh2c6mMsWGBkUj3a/hnCf0zAv9
D+a8z/pJJKeE7u4p/0M6I7qLv4pKYfIqkMeKo3wuNedPzi+fe3e6qSZrm2EQLdn7
+Lj/czdNw2JJM8Q4khp2URcRLSyKAdIbKfgb9P9GQnOobWKzXNgkMyXpjRnKEBAj
ry9399QuXCcfYb0JwrkXlze6Y4gF7N+hrqznuuZkFixNWwBxGf0x8vtONPQc6gdU
MYFd1CuXCpcbQ/ICULNlBBAzzmws0LEovjl9pulEwqKr3yiDO8wvYTYnK0/Bj1E9
htuq07p4S4v8bY7wyjkyJUFZbi/cenW0DnfBDKqCi3GhsfqM0BiO+NTdTdedkx48
vvmxVhBSYqHcdsy0Jono5oo92Didct9+pLRpbNBcOCuEmEf5GnGiwJLvKn3RPYTF
XDs7mBMqnB0n2FdrjGs82pO7JRge/4Zx8RNRRw65R+Fz2il9M7HMRNVIRSQFD8Sg
Xdw0bBirVP0U2eWARq9fCj7HoEDeZem2LSG+F0SgDrHGUK881zcacCon9XEjDmBi
XSnbWwRd2loZivKluQy9uZ91jRRoHfw3ivChZ3G5iXDiHgXakE5yUO6j6tp2lXHq
p+f2KjA/HAyO2DVlzVfWccM6ESKsPGESvhV/FwvlDlakh6QTn9MJ4+L4noHIfUMQ
EqDiJT3oTLSU4mc14MFyKCaJm430Ea2G7zzIwQBUyXctRkPy6oDOMcI8CxQ8KgM2
uFSs0VeBQNCOAPBwBMympapYmOFO6d5dlZ78Mh81r0j5aFHkedKcTNUnc61qykQG
VLA1OyitCUBM1IEAYBsI8FgFFIUn0kXRA4tvpYkIuVpmmGu9pxDeySf6uGbSgQtK
HowMHpAzs/bm4N8dOYiRF8J/NYBiHOYQA/bLrYbFWdQulHXUh/dOrKDGQ7VlG+4H
NxRMd/fkXBc+RHueyyIG7omI1LHt/wst4vNYMgay/V3uB3bFnE5V4nW+/modah/T
iuCOCXtjQnxBDibgvbo3RfDD3Ge2j55p5htgCg0f+CsqgQ23unkP3C1plWgpne/j
yXxPIaeU3yW6lbYYZ6MOaqm/datCWVzs+6YtisKUgurpnomuiNaR6Bvmu8mQTA/a
oJkCjpZFL8AN69zdbLAJ+KEhUZ0MuCMtesl+SDpHKVDMkAI9Kh/LNXvkQQ+VhGuj
7SbGjEND8zUymd6jLQrORy4Raz19fbBQo9qd5Vzhjjak5PVe5UcJyYM8rZIe1xwu
y/Gw/rtYkA8KSsqiLRc7CHstUcj5fDlZMspM3MJnfCHkM3n1FvasqJq/iajv5gQj
2gVZLPxJI2X51JAp2uYYEdRZ3OPJWwm8ByvCz0i/PyP1D98VlDB/FOHvrUHWl3bZ
CISuY9ue29HAYQ9/b9f3ibPSEtj5psIW7PScUJ6epjMMVpQj0eDQeGpbf7CyD+h7
gD6T7fM3h/A3oLc+qqYJpz6Xyi9UeiRuG6cQnLIXMrHEinFW9fhbCwgdEjM0Aljx
5RY651QFAhqicsDz0hsFOY3vkvIc+BwISPdIuF67HhKewOUWPxFlqIELCO21n080
XbPT0YEyhjOyhVnXn+J7hRqKeec6kyd+Wd5Nq9aL54kGGFaj/Q6Z3YHnXZ/kWIbN
Ci7/YSdAxn4G6eCDZhjuN6HmDSScQTQlNd6NMCUKyDnQ04O20Lmcd8C771z41eNO
wTDOie8LejBBJ0d6V/x8X+9pqdMdBadIpS3bwhK09KJgzTKGvs78BNik6VAOx09w
lQl6ahxG2NSvnT436ssRLOiQgB2DU6HOr4UcitWVjjf8RbRdAd9Hkv2RQX2P8XfK
i5l3sM9zBhr1J/Cee8E9l5LEVD4+Q9kJxanPtdjsG8uHQRlGeaXUxauA1ndWxJ+K
IgrEJeLc/1u673Duvf8hke8VwGXWKwA9WOvC2EEYUuyX4RltUSCm6Wtgjxq5cuSL
jV9adNMiRhrPASX/byW+MzjvsOsuDOvjXiGfh4NndhoGxv7v74VPi88GPrI1v4v7
qnBmHY4sCLzWb4dzgJMz7acbpRDPrNNp7Cukb++Y6Ow1uqYDuHuiT8awZZ36HZpq
XU7oSXI7bEVzNxdm7VJEKrtz0tLvurI3t441CCvZ/5Qi0xs0S6g9zr4bi5hyyRCC
dj6O6HUQXVgscXTR65Ccj57uvY2wmgUdm5TPOtIsp3MG318Gld/iIVzq6mQBy2dk
gRol0VD+XXX7dj1LYuGbEbXH9SFBc4cWx7jq3vm3XModLogPnpkDxBDCuQ9BB359
f/ygaLWKoMoz4h4rKJV4b6bxXGMxgz3wMxe+Xi1b9hnB3XB9rQ7PL1lqD/D2vVKy
z7wr31hi612dAYRBCisDqNFajKs8LZyKXNzpYdAG+SbG48EOl5Qm0UdU6FXQ+9Gt
Xh/vf30imlvwvRb85hOzifdtvOBGdraJmssYKx/k6EWf6Y1QCJvs8MUVUN7IBOqu
Wif7ojZDsD+k75xqx5wMVW+WgnGLraBNjOg81fEPZ+PK8mwS1lFx2+/cGqHrcztO
IxS5bPR27jSKU/h10F8DSFdTEdzplemVbCe8I9bDkebae0Ct6ETNJyphdPZgRVHA
oY0z3jpAKXFrH7yhneU2Jpt1V8j2ruXpaX7qJ4Dd1osLsdBTqVLSSdGWfOrYhxiv
DfNpWitfcevx55drdt0G7nVS8o9Xk2iDomxWfMYEdvFmcquFfVK7yfvf15VLZX6x
1N4IY2Mpm0lRE8EQ7FvroXCWJ5DyiCR30OKZLsb9o6FT96p5c6Aty6dgka4MOnjP
eaWNl6YbxeevyXNM+E/KODPPm1p2/n1+YMla09pTANcd+anE1VWa30eU+lSZDDMB
aPe4rUi9YeK4O5fcba4e0z3oEVm0Qt84HCaKonzNPDLDNjnR+tGtP3HgfxsI2M7A
VfB0uEEDcSHdLmjHrMwiek9BV6GWQtP0kzk/vOVrL3m5tyzWbl8o6iAfOUsIBdqG
gDKfZGRFcXymVBAqlOXOo8FlSrnzpWeeT+o+QrUDg9bvsnLNfTBauDAZoIPYEiIF
3s6xDArjW/+xiFbZKHYYtBFyQ8S+psAG/bmdOCxdOm6yZtCicpXXexSEWw0dm6/m
GPKpzsQLqfoTiNkxN7yC/s4szelWUXiTiISRPpdR4jlNzhKCEcI0ZMLaBXLINsoO
+ngg02e5DTisgwfBT9PhpANjhsRT0u1kMSTsQozIm7zWsUk2jTqH/u7Ntw55hVBb
5725IQv6OUW6pVZuz3dD4jNkv8m+ZoGTA/4398L8Idc2UeYk9rW8Z+nbL/eSYmmV
pec7Kf6XqVj/ngHOgkrhPL+XG0ynFcqLxq4BBcRCqeILQr6EMaVJbD3QJTrZDOzP
vbF/2RwbjNrWsByj2ooNPFn2ixJpJG9Gfw70NlprdZ+SfkO3WketXYERunlWe67e
+sgL+ddeXYoXXhI2Tlg/REIefqOM8zes4N4e2/PD0UN8EJ6XK9+nu4xYBz2hfF0N
m85CIGX+rvE4YYTJ7bicVz65VkTE243b4mQ4T9HbZ5DzFcuiJ1EHB7cJ4fwwuX5h
V6RnHsWPYHCyjcCdzAQ1sF/QLVMeEwXpL+JHvXGYkFL8rdEj7alEgWqLxZ+uNtYX
EaOMBRbod9/vURrZoCnsSkf7Sxm6sm4swRj/h7qi2EubQBr8kzTNw0CvwF2GYjBx
sa2h856fwPAyEetn3KGVaywSmjwntkQaVRVT7neQwbRa93noZF42Kw9Eg1g8BDnh
urD/Qer+z8Rje1lnTAljihgLM9tMElKC7nGYdldOqS6utJT42SXlsWDt/VY1bFp6
D4t3ER+Vw/WbJfz46jVPAlCSw/ivsIaRBS5FBLFo+CRXuNMhBWLjyVuBO0G19hUq
3IBOomwV9atCaLj7zzAPqibwtrZAEYt8HK08FUYqdB4R5bzftnMWDToFoKQ0BOFV
9BnCNPeMJDFNF7ha+8NnrQk/djFjmodaOZhIaMrCnqe9bV2klmD/eSKv4+iDO07O
vEYEf5w8u907hwO45KeJvLh5++dIsr4XPECJTl5oa2XM91DYskJHNvp2prjJo/Lf
TNWNrg6F+MiFDlA+/ZNAht8YhRavLcdvOIUJGUFmjqWzcLFKlhvucrnMcgPLMZL9
ojDyxd+1TJW6lcyR5C+e93t+GxJYoUgnm+rmbSHRAWCM90vTjNvJJb3RjKuyn30N
pVodSjZP/u2M2LAX3aDmVQnj9W83fo5/dfYTkpwJgKDnJ8pl4XsS2snM0wmQEh0e
181Kny3KNuO/0lgKuzurGOrGZiF2cUC1iveOVxPC3Lhal2hQmDq7OwlVH6lNolq+
fHo3ULbPwF6Q/GmhACZgg/mFeaBnwuhIeWRbeVkITQ6hjFcSWbM880VTSIkOn+p6
o/mxKM7/TfBO2jTiDt6fM4eBAYHzZFB7BDW7Wakca5VgkX1+K/5Y3yKGQ8Caskjm
CTCQgsqpVdq3nKy/DFGrF1mGIGquaEWN+47HkugHgDdxpnmn7rZtMzOJ8hg5UqlP
i+c21tFKYIRlxH1JLFI9LdrCq0ijwFbt970Mhsg3l84ACTLaSQnazkRucLbkqkLM
3BDQbLocv5mXG9G5s5hG3ugkNX3pcprrAmL+t2qpIV0ISQ8dePDR+0FuNDv0Uaa2
c2SZ5F6nHFBcp5zj3l7CDf9z7iXM0hL7x7fp62lB9nD0Oga7dIa5SjGCRTA46nhZ
yZdOD/gplTQl+rBnsLt/75SRQYN46HhbsdVPIFEotnoOFeMUhvPOF2OyPi5jnQG9
5or2RIWjGTboSwzkWl5YuavHSVUi8mkV8v9O0jKNKcMvuiCNjSLl0qmXXP3nEIvP
ni4jFcUY5GQSIy9Zh7g7oMvQ9XLvrJDuIf8aucfP+0HBcASfLUPA/BiKSrlXBJw2
VkUmYS9iAlBfGwiRSl+O6XwGYKwM7F4M3Eab8qZzvD66An00zUmUR7dcfqERj64W
sOKrj+8Y+bB/J2LUecfsxxfq8EYEySNEJZYQw0qjOJ/6nE1UbwwAeUMTuZV96ULI
LITSUX3he9TYrDTKaTn1NBom7VS6rHYs7c2K1O42QNAsD1DkQtiaih/XFotLpfzi
uWgKTMwWo35nZ6tYOstrFchiMear6qJne5Dvnqu7OFbs31z/aPApoZwQgQwLNcSF
WgKlOYm1fp4gDuaTFRWr/dF7SHaL1BfHopyWpJunH63PAiZl96BwxLl5sOEVUr4g
Q6JVyo1UNLh3WOAaHBROVlaBd61jyFhC+4tpmtqUAQuHOdHyiKIOk1cAO2azKa/0
O1luPb+FBlcqVPOSK7TNgMaPBvHhk8VzBr1O1P1qeoDHbLmKNTYQkll1O3mV0B5I
njm2nRAkEBbGgwx0+aWoh85IGtgJRnNaYjRczVUex1epRA2JobRSnraXZwKEP8CG
K+dQtYYiOP0HCzd+zmyNWXQNt8XnTKIavNUWEP1rnKvEMePVg2krOIEjJaCuj3Da
VMYkuNow+7FnyhlFeI63eCJp43LVlizq9U+uEK/rF9zIcHOx5Samft19aUWKyDlz
IvFyiKSuayI9rCdiKPYGz1N/uUR7xsrXqxrJXXvTO2T88Mr3oAH4UJ2wG1HvikBA
E5QS9X9hWLX8hYZdCPDFMlwi3la0//+5VM5ky7ouvSA0xlnP5SCqB0yP8Exl/oqy
9PuzA/cxzkEsFB9ite22WLYSOhTjWd8EPFbQqUa1VJXpP6FPfk4WxiQMi9QBqzIu
jaP3NR0/tH5nWR5nAiUDl3ezzbVv9qhfQdg612oHSM18VDzmwFI72hmekr2KTgnk
n+MQl00/UhoicXp/ZBQP81/Hhrn2geDz0JvVqFG8AtD8vbW46z7Smjy05eA6go4S
TglKMxKYLlGzGSfE3U71dqn7P689Hpu1PqLG4Z5o/d3oFdDGKZwhqeD+sVsyXLhv
g7aLowR+Ivce2xcmFaRdPL0Ce3CNnZ28gKVoc9iZs30GqjCevz3th6aXFa0g4u0n
lIhKI7ymVMWHV2qS8PThP74F6Oh6x76GowzCyn0svml47gx99HBAAsgiVNKh8kuw
412gg4KGMf8TAouFqEzbI3hLp5yCh0g7nwvYxYrDF2Hg0Kh4CxRbeCnuvhKYQfG/
uCaFQ4kyl5+IX9GJMoq6wa1x6z6AWQh5BkbObCpZxoHPF08Nc0qYf3eSDK76cBr2
Df4j0/2BDBxW6McGxHAOoLqgl44LSrzP5qIgXDPa7n0+06c8Hx12pG/PCLSo1LrT
Toj6gMxCmJgJbnE7yAWQDFc3T4wThT05n4iTekISvSRC93mVUZlg8gAfFePVQx9J
FV0h+/7iGSYP5OKBwCfN0JSZfnDgNfPDN8Q/4YD7/1POWRHWnmAc7DebMDuQ4tGk
gk7980wNNAQb6KjK+hDGKI3tsDh9KkDt4qBZYatqdKrfIgvN3n/dSxuPbMI1gzaF
Kf/B2Ssul1pIm2UsgontaKXeKwfbXhDhLpokzLl31urjZMPmChCa+3fAPH+3yPsc
kog/6+g0CrBAYlQj443zQCA5IdGZ7q6CkLFQAXyAQqZ9H+sgsStX8p87ug9zkMnC
glb9XNqBfs1y5hqZbntZeNw/UbW5bEtOMudZP6agOoPI+a3U5kZQk7k6nsuOxbx+
N8bZb5gGyY4YXE+p6IO7kppWoocQCX5KlXPAMUCenQXf/St1jBZO2KJDgC5CNGM2
v4ApNUGniE7e+DcGLOc/+1RZfXt6Dy3g6fen2lkwLhy3NYrEqRmzaPwagm63BwWC
2qqdD18orAe/ROIm4Og4syDu4Z8zbynYiTgE8jD3UD0cta0fv1BCZp8ny61C8niD
aCWcuJo+Poz46VziuQnR0vWFK2q29U6BGyatE42FDJGpOliqlbFpMEVFUkWXliDC
RQAB+nOBC39pH4ApGDIumoepWrzC6zrph1F3MzS8T/xXdmgus1gQ0IFWMtMi5Gpm
4uGqsH8xnenq4u624q/AKlg8bNlYkv1hNnvT49SwlsH6OLJyF9k9r+mH4S+7rxTo
VD3ZOlrK3CpjZV3hjD/IYy8iE8yLIhOkjM9NgaX4GsBW54+g2aD3CiogNWXHVd5M
eGHqaexeQdCLcXEMxlWN5QLSfYBZs8OeYONTaE9ZgLi80Wb5f8p4nxVS2cFtTadK
fUJLM5VECFIqF9TwjbO9G3vuJk0FHtCTK7tZk21IWGBcN+PLvLHGB2jXskZzsbIQ
QywYXI7LlwbH7D25mogCT603Ssh3/JpMh7O9Ijb6m9bMgibaIGfBhfXiZmh0eNzm
ecfXVacgIaLVpCoi9f0PaQDqmzkR0Ch4Uxl3FPdUq+Yy2QPs3yhu6yG4KsYjAXXf
qc1LwLMmSXNmDdxLkdeu5/twraqWYOAaELLVsicpJH4rOuNdWw4hBNdRsWxSJcUK
pgCqEJz1t3KwEN+5Ly6nUa5L7T77BMOPZzn6LKirpYxnBLpmPjz0xvPbh29BGUTI
hMDdLwKAKr6xG2vELdS1Y2CTP8rKjPzOpLtvVkFmFq2iZ6fkk67MSZF+PUr933dh
UxCRMPojVFMMi3lZwQxPuNlum9LtBo7Chk5+QusGfwuzhULvAKv3bgy6dvyhoZyP
greOL9qaPGEVTAz5vrUQBha1DVKgYxNnSzl6ptFMjcnBVmI1dl8IVO2IXS1qPXZl
1dKiZWBHIpGzYQ4Kv3gCSWCeCEge0bVWsRqC3epEt1H/h3qYo/8xQw6xNQQ1iLD1
SgvD5+ePi2w8QpJoOyapXGtj2MggWQVWs0ZLGWRgEe7rH71KA9SIIPuGpoq0CBAH
QsQAJo39Xq8AWRvTmUwmbGubBMwt4MUSsXQSJWZkSi6z17S/svXw7nKD68Q7rEzz
p24qkE72UHRs9jaTkB50dO2Uaf/vnFbi2UGv15KE2Ne9tFiUeqC7eWiHBMaiSKrU
4nQRuq8BrQmZt8o4gQh2PzPv9InE0Mmf8NkQcnyzcsPvuAZpHjcT6niyuVEmsNq8
nvZHdrzqd+7pHM5gcOfpcl1+NBXU9aR9b55XkWxFre3P3RndABSD+Ib1AdsBfP8r
PyiRet1ROPoqwPRD1aoTE0Oa9NsiaqD+mkXHn2uJJcXSNpDsU0GyR6LUxLte0daH
Zq1Cam9O1cyZbDq4071rQGfBey8fa/Dfdt9BNIMgmueLBbaK6bTYn0i60I/plY9r
uBZNuXxWzVRFuEbC7/aR02MNtakOLkPuoHXYG7B4Q0scGdbioYWU81TDSwJ8tF9r
eOV8QvDth9gN4VpjXjhsXZd2gegIiuVTnRBbh+LkcjJX+S/ixKPcW8jfXPYx4Hn9
3uwIGgrBHp4s+7TRE+JPf24o1WwnO1U4Rl+H0geJtetqZ8GeyBb9Ef9tVlMyQDR5
SIUQc6qghTl4LKcLIJO7itlKtMxjQ0tFCVyYIEHbJnnMJvP2rAzR26mGc36l5ArN
xDMhidarKPfwEBMO1sKe+Th3QJuTtc0ZOaGsygdROCvKDlDOz0yP217BalHr1N/j
s4Gf3KTxr81voQlBGOJd264n6vUYPZOdKK9iMgadethQyjjkI8yklehF/Of9lbpB
H20lS6/zxYEriy55Y0+VrjLOlEMWv2NUkiPB0VBA5pJxKGiJJpmD7z3843vONSoN
ha433+NIWMUMDmkYcat+R5QCDykJXEs3cPBy3GwXclikHP7p+XbRhUJWlD+Edl+3
/oglEXk8WFQNEMK8iOWbZRRSAHdiJAypqXpv/l1+YluPvec9NQW0wo5gbmOb26kh
1Zr5ediVhu1ZNlEY55EOObbbdrv5PAo6fIIBMq63PtvuX23kmbzwJEuKEBOyFAeI
DwyGcgIWI3ofT2sDkeU8tZ7dJcL7JuJFJVSyIVQyVmFtVwM3KTUtU2uIXNFE2u4K
xq/6gVzWT1k6Lh2VDhhcgzPsZBCHIa/qt2vAEQhrxeYqCsAXGb/bjHtiJnLc5za2
m67LoLSCOrqnpF2Jfv28I7nzd17FELoOBJUMuIGLAFMAC5PwK80C9nJl1b558DL4
sIFkjIIEMDNRmCUBuPi8gvh3bJGtGJEoUJ3ov1JNKLe0LBKfqjVkSxGURBabEcb3
7b/TH/Br7REJwoShZkvCGtLcZNR5uNTsPR2bqf150Jkj8m1SYGtpA4U07GaBtFHw
5BAozS5IPbWTl/g1vBCAdC2UavtfpRJPD+aIN7eua40sPBFCU73/SdJjUN+Yrkhr
ilWh9AxJ7ef/2CaYkByAiARojwXEfKvJ+psgMWa9TBSkRk6lEhSIoJvWttJSeqR2
mP7fKteS92tsqemzzJuxxynRRWktcTzyc1fuw03lW5XGdv/RpM476zMwCsTZKptF
ft+LL19MNYJOxqrqcbGwWNX4k2zt21TQf+vOYQdZh3+cj9FHgqzieW1PDRhFK+Bh
zLKPu+hl02a96tDGrC/SR1zuI/TEAwODapCoY8nMgTBLlmJKaTLYaigrYdR8wxuD
hW450ZTOcpv3UPswbhdJydWP5zUXE6hfndUGH6t/qVFD5F116iPD3SXzgR2SYe9E
dGT5t+3n/U0kn9cUzhVJSYuxsv1Y8Jgy4rPNoudlDGZdwaiqYv3D4hUzmIfap7St
HmFkFj0e/X5Vk0L7fZUg0PzR6tNLuIO541TmKQP+t7xOcJz2Ch9ASEXKTqP2IICu
j7THXw0jLSyCAwwGA6m1Vcp4dYrvqm5Yl89wiMNHcz6LJ6rlBwvfaL870oHYdmz7
SMlCNqAU3cxrAT+3EqB+Gnq1IzKy+MQ0gewnHvnU86bhmqacSnZl6zL4ZXzsnCYD
ylPDMEYbIICnEnu17o6YjniM04oT38JTUrVt+Wyg2h0xdkY/wCWYGfqxAA1rJgMB
/vVFLfdFDbkd+9Yts/ZhNJvWhMXA1HixYxWdKJhm0uzyVYuplmM7IdrZ4Jvyx6TJ
qiI0cbvkWHJlYdXx5c3tLZtRMGlAvpIsOg4H1H6ESi7/pcSBPI4EmEs6U3eLA/vr
hKFy7fEOtWqRdJKBiJwKbNQn55oeWBIkC9OPtd+krS/Ia4gppBK4RLfRbimSE7lS
wCV3sty73Q9Lb/Hd8+XHjUMocquO+8V7oZ8oTS21JVkR2fH4nTRWhyuoYfxsq84N
Mv5XcMT068DnM0ZH6oVEG+OSnmyUSdqOvu1kd1sFYjLcpgYsg4Sp0fy/ELOxp9IK
Cc1qetdGapnLxCxLdTkqBZhwLZRKbP8ouPYOKEp0xFLX95dafzMRIBewLesaDphR
a9PQdcDko3W0rDsQYmTWW9yNqVrKzSi0lHcoeeWSSIS/F1vhNTD1W1g3EoG9rFgr
X1ZR8SUJ/iVmzSpC83S6hFCZNob4Ypq5X/7gh9Ybq7pcUCqxYhE/h6xUPUpxUMB0
DFTis+phfZwlhmY3eOOlNOpIuMBDjrS5Xi4xVonqAu04HCQjNeOx/8C7kLXJy31u
g86u8paPqG7m4L1dJvTaH/FpV3hUqpC/dVrUUYjfR+87sqDxSqdqZAikg1SO3Naa
8O4Nh+ScxZ++aBujP2AXSew3BmiP05BDK+T92SyFRL1Pyjxi/Jr2hVNStEgw12dY
WwB6cnBfKNmfEQ1uQN/WIIyrz+bpqc7dz0iYP0O6TebE4lBoIAbS7Vk2t6ZF0Wqn
jiBFu3lNcf4bV3zu6kcloDONObPivsJ/buqomLsQ9f4UwT2wzyDbDCBgm/gB4Zj0
JWZsBlncK0dWffPVQL1fgZ87Jva1Dq/vJtG2fHMZP95YmvDxLJqO8At7m1cWQMK6
d0mgWZ5gqNUazQmGM3u9HACG4dxilorraKUGwYEPfsQ+9+8XG6el19s87tyvhzzy
KzMdhx3MdAcF9gCM6S4R8TtuIP1RTYFQRrCFMRBdgJKkxPr9c2FpWxKjHfadUc52
x2u4xOdE44HTXBeZarmu+yYHF6VODdywvuswva4BdelKBfdiuo1NsKyR8ErNC18O
2WGn99xipOzd61gh3hTiHbPCwzpvDDvgyQQ5g2TWW2gywnO/ldmzQQkLsVpJp3aZ
P/elQwJprPgQ00dX+6rl/GTcEWWBvBTNyS+zqNL0C7m2lWVhAgh4A88VXLrfgPjA
zxy47Qx6QdwfWG0S9QOH8/gAikKUY/0clrQMSnPgEZ69171Z1f4vqhtJHXyd11YI
p70NnYUzLnWafWOHRj6WEVDgHr4lIlVAZGOTs5BdKf0gdSQm220eyrfz1Vw+8IZw
jFXQbOfdP0kqYma11dZA9Sfr3PpCa1Hy95FvjsKzVTckC52XFe/ALwV4ajdcPhnl
9nTKhLBj8HMxKsiEeuBRWHsq15Y7pk+G9yeliK65feORwEN8Cd2nI9QfrZfIC7SB
rjJZIWh5IehzYO7wv/+nC3z4zkeCnm2p75hqx3Yvx3zjIy3Trkg5IvLUua5/XKCY
Is9EfAhLea27WaClCDe1qJ98l3NLlhGD+kindT1rfiaIIweDlxiGBMtcUuLT/Y3t
tGolBudzEdldutw3aH4sUZdzEvg1RCMhUmdlqowYuMquOo8+homnhswsAqftkkge
Zg+5emmTXX925WdL1dxZR/DCbmSLUPEFXPrmscbgZYq/hxNtyUOe00hgyFrERUQo
/a2QbmliShYlG7eJzb+LAz11yNCN+mURXuVYwBokMQ+N63pnSBoctKMCcOO7dx1d
hO3i9DM4XVH1+Uf9ztdLvKZLkFZhJRhKwIYER2dbjHYSYiUG3uGgHtvHVGUuSA3J
0b9ps26JQyB9zFO/q1uErK0jBAvKQNZzMdfJjxek9vZ07ozVg2IJmrglDALyslKI
c1gqUP/S3Xop60gnc49XkEaQlXcu2B4dgwXlZU+VZTzSW9MQpht7z4aeFVAyw5EP
zbX0TO1DcYUXbshlz3i2/rLGbqEKs+9XeSYA9Q5fnQT95ixOeb8i+Obr1XTdfIsG
k8CP2Y9CPFO+7E4YDQfuM+8X3FvgT7CKSxqOyR3S4zvr3RJOoGhMojIA9GLeRozy
T4yF5Ce8UW8lzBLTaeqjcbVzFvDHFajXoQJYACn0QzXoueiArf83ozAf3b2pzcK7
fY/X5S015x1zVBou8B2/W5oKpoZgWDxpQ89RnVUxXeaEYG75EaiTdkW8CX/d7VFr
DX0Z6blwdEpjZd6jwTVraepvum1oeN7AQchZS4ZMwLNRGRH9TV8N+Eg8BwBcaULN
vGjz1JjU5HMWTfoQv8qq2DsJ+lHiNLafynbbBdyV3ldFhtcHykCJUuVm2ajMqKgp
rU/9o7+CQoUmxL1NN75iUgjQAkxo6sqFUH/u+tBGRT+gdGgDciMs1z/kdqJB4e+8
eoJfgA36upUlzcEdiEY8LjGVmTUWqgtatPh3gkL85UpCCMjlb3EI6y5E3i7+VZyc
QyN0IWRhNVPD/LNuKilEK6vnKcYUQtT9o0Pr8qIEmQeOLPARY1Ancu/mWCbSWmmD
S+WIf5doIg4+5SDYnBqLyJkQTNuU34PGKI7WOP37Lyz7fyuzawYtp6R9shCp6q33
diE2FyRu/CTp3jvZi/Pyaz5WHQ9YCMOeArnShY0dfFZ2P+H7gh9n8LOtcKhe0ULP
CY/hC1ge0zsC0ycGnYCrm5Cx3krFy7NdbH8QOjDxW9lVmyOIXqQ22g2t2zCt/4Lj
q2igwUCP9lfNCdxndQbstg2Z8MKRA4Mb/51CfcCoan47crNSlHWtyEJaKaAEPtKM
yuaH6hSKB5mnNmyL9AoeVY3K+goxyMBTtAeSbhtbO1puOtOkBMzhIr2PRHKQezpR
35ehiC3GFmFTUjzgJncCUJuioW9hstrHlcmIAz9mBD9P6Ga5ItNQ/x53TFm33s6n
iTmMc1YduF3AvLExjWW4Uz5+oB8gjvtH7UggwYgwxl5ft223is/2Ozl8beb2iEsQ
Ms1Z6RR5TgeUL3JwJ5zuZ9OFfQBXBvEiJsp8rloq81tyMQ9C61xZvXsic051ybYX
k40zv0VzmALYRql6p8kXhfh9DhLomqmNdMNeMP3totJ6tIGfFNy9NLPQFaUucLOP
6wgj8YZaIWyKDw5Y/3vOOp1pyJYPrSre5U/5+WbegtECun70WzPVS2bA3RgjpZVF
ncqb3HVJ53sPNmtpxYvRHktLaYr72dPhEVtxMkpsfLCzYDoTRi7JRUb1AZCillx9
1zgqqRW1CXavvVgAQNBZm1lI3J7Lw1YcZqPFpe5eJ2zjPFk4lE0yFkWJVwg77mfp
B5wg507TDiB3ZlmoMEYopIWXAbnAv2voVwhLdjXZrnnRn/o0g3jDaufyS2yR2x08
fUKIoKl56EzhhUi7vbXq86Bn/zs1yNg7EcISMEuL2TQd6GNMWfJnXuEQ2n4/LX2R
Xctim3GABfnqb0iCB4LHlycQkZytCR8i9oOMkNhCNgMXVVuUiwmP1mWM1eUWbylk
Gmit3s+Rmg1EGhkEFpD50OfAVEsZ+8+1geZY3awTZzUf3umKtxB8Vk2kAvmTBjTV
6okbB2VIEnAfZuSbbqK7rbxJO/5RUFLQyZf9T5tt7mWPJgq66S+pdcgl1JOmRIH/
u7rlyRizCiEsfcf8DAqjPtnFJ5IaLJcb6W7axXnyXD9qiET8ipsgoTzCqV+UtECa
6Ec0Y30ZOYhNVD/l9s/QsMuGNa1fhziDckGzZlOM+SJaWVftyAnICxLVePuW05vS
fi9kWQlNKP98GA4U3TL6JO8fJ0Ox0VOo7ML5Ww+bd7aeo3OyZ4UvYo0BJQNt8DOC
CbevDCqfTg6gEEheGymHKjMT2nNtazD9106r/vGqiqSph9k0peCaqlKAKg+MhuMr
1OjCQsQkCcCj6aHuK/Yu/Aki+OyveVWWUM83usfVvTfog0MmCTBqnf2f/jSRHkCn
PFqBxI9Yu+X3lxwsCjtnYleLJ12N1jLmYpBLBNs2WlJseB+FVIXo27qrWiY7Pfnd
UdmZhsW7HsUr7gxrv8TDNPiVlue8JAxHiJrDqapu8+IGTX6rCOWoXBOUqpHTXTlP
n9bXbbrho5ym3baEhFDdqjc0tP5zHkJ1p5aqP5SjhwKJZqBShGgs1pYoAmihTl48
ynLmRDpq1kPzVx+6eNVsWo8Dj3NsKiQoZwu0OS21O+3RsLjGvVwhHqKHquS23J72
+KdWUIii5z+IQC5JQrvAR3H08Y3yWS3zaO5PHseMsl68jrW2Kusivh6ZYTv1zwTH
cqNwJQdjbyV4HtGLwa5nyq87K36kxGwZtSFvnOLN/9ue+Nfv+4q677Ri4S+KLzfv
qRG32WBnm2cBjZsMsnbcKE48SQZ2gHoJlVwtRa0bEklHqHFVlSaquLf8Au5/6IC/
vIpAVNUHeRUanyatMt3PLhbIaM9k9fEf4mZFkdd5W/AHI9AKSU9iPogjDpbl0NTP
WvniRCDeHVtpVA3Im+7YUh5i6JlBtw8omqY1txkSlgaiwe4L4faB1Lym+WFlUGyG
l222oInEN7/NeYtRPA8c5vWrlle+bf2en7LZztbIGBT2LVaaKNMK8TU3owfyFba0
V1/2isWIqXYIaPSrldq30Iya6JMBIHGxt156eXXwHXbKDniSiRcab5P5rt2l8y+9
PdQllqJAjEuFJKh7uSRdPCzn1HVRvK6u4uxdqaBSybLYS3OpfD0NfVk0n0ISqcQD
ItaDoMn0GkS76O5C+uev7HB2z0F0DMVegWRdBBjOz2O5CBS6k2VpY3ryMH15NVBi
KOPgnc3FYPAx12IEDbIVRzWaDv0xHa2HD6wu243OMTtWHE/6qfcKxcuxpHszw4hI
2d1TONUTIsHaV1zedCyhriJIGnJy+IQe6fsDiTK7gC5kHGZbgzfh767Ldqc+/Aky
9zuJjGevMwXc4JjwTVNkxCIP4V0P/Nunw7K6OYPmj/7PKTm/y6Am/kSYJQS130+9
lNOPnEeZ9xghOwm3CiPhfh1gN2QdrHLV4GdV44bwajhjen754tO1KbuhZmt63RB1
zzRWZIIU4czgmfy/jjGFsJ4PSdzB8GFXew77MuiPy5fAeQVSsY83dFaL2mOrvYk+
rrB2N7/YM1sZq6SDunrWFVsAPjaUArZG4Z92h1kNOP9MpEu4WnJ82fn4B5F2h2uZ
yN/kdyxVdIgJ2qGpW+baxKw0YSmn5SjI4VVo26CsRj0sFV5iSzG8gNQQ59q37Vek
4D4WswyIowA3RZgu+YaDO5sJ/7NbdLp2/thxJ1bni2gTLGYHlLATwfeqFpW2ul8F
sE7dpRTw3TUw0OvuLR7zlQRogV5wZ1yd8nNtM7E1TgCoh0qtq+f5wI98MPpDpR/J
entntwUtrp6PK3Any11cqwtClmFh8rPxmyFrITiSrUOGIsuqN8egLxMUEfir1mZz
nY7S7GC5Vf+c2LJVbzbdo0K0iBuLISm8A8f+A9ntON2ke2jnoUGOo9V7AW01blxe
f4X0zQ2Ky1D2z+KU4WXOf83xdan5acsVmCMpujIQkEeEUnZuaLTTfU1UCCnL9HDh
c6PPnvqlJsBwrxtm3WiErqJ+592cucbuzxoivODlBgK3N4+ZBuU9fRffkGDaRydU
lGtBShMmkUWG5JCAUT6IMKZJSgtwLJsRoR34VV/7byWWgMTYWqdSiSlbp0MVfd+K
BlaP2W3YXpHeQHa9lH7AZz8ZnXLZcWvC9M3owzLy5yLJzckTg6LLnATLaezqvvNr
G/csGYAn8ezorgVqnKF/Mp80X7cjgT7jaxvUwlw6JLdRiidIMFwj0dWtegxn+BU5
gseWewlVIM2/uir5HxY1ZtyAK6WSYcGUJ8vjb1KvlzCpu3ZW6huoxcbkQEFbgTxk
VAc22u9xnYvAVfj3FiPZ2OGbr6QqfFeusdJcXg44YHb29QchxhpjtFu0bmwC3Ez7
FqG8dR2FIhPQTkUGQuyGVE4dIlYi1gmBohXjjSZOVgui95cOQPpVFyHJFW5ortxh
fvDbmsG+HI8yLjsHQIDwSbNEM3nXVFDmVo+RzqNKwnLFzWaVXBffAHS2QI6FOUq/
jh0zNpmB8dGHnHGqppIUeqS8w7if1WeRRRmMSUXWMtt2cHN2Jpkot3ncRtrZ56Wn
eXE0mBSShJMN8T+Nqg4BlZokgOOSE8zKLYe4mjJkr2hAASFagxnXRb/QHfHQ2H6l
ZCe2Sz6FAyAJwy64RjeGQ7e+WkTfZAS6ckAH+aFYkyEp3aNR+mGuWbteVrgk3HMK
JE4Ins0LEySStsPTCE+dnlIHOu/1TesL1e0Peb15DMbJDkEPEGvyqiso73FzRByo
NNrMVfxZ1qCGEKSAKtisLh7j6UMzXbS4F/G3oo++/dqfta8EInecqtRLrkwwNj9T
2ecIFVbN5Do2qxJkIUy6xIzEkTWuoqv4l3XAPZgvpeEQwQ89E1iEh71sG1g4tKsU
uKJ7sKcNaHt8JcHZRgoSPMJUILGdiRnpyB5brJu/GEXecul0Kvjs76l4XDrVXBQG
62JS68WrtFQinijlp/UCM7Ql0SU3ejggftIZpv+XFHDRbIxLUaGUGHhfrp+N363S
/7H2GzW7IIQK37uxRkTPnj0atHCmFiqbedxvs4KxK7iMwlRG1ZqTIm6GFMFt4EWT
avoB0JzwzoUOHKB9uOCt1k/a/b/bmDeFTBPb4RhEdSQQzdRTfrT8/d3DstCBcwAj
IBvUxMEhjGykdDMXxL9zP0wDI6Eb8dNrED3UtBUPzWqMUwZcdGSBx5BJIkDwcdJ0
lCLefNVuwxH0rT/SUX1LH7VMDE9szG3Tctly5tDtIe5j3aAivJmc1yNQuQOIxmbm
+SoCwF4TWKhY6qxomIHktDHIHCCRcEGA4zMzDZGQI4q6k4F8W0aeLjNdgtBb9sdD
uy+myyZ3QSV4s5kYNovDbx40DdE81nRe1zb4BhOt+Iw+mxrCrhOyBEcPZAHA4Im0
2XhmXXWBQnEckGWoJxOsvc0JdQyu7TQ2bD+sboOnqv0GdICfa2aQcsU8Izu09xS4
aXjLEUjKzxe3a310DLnecVTFE9FaGstOgLY5Jz4T3dRCz4zohNGgnMBhHE0B4dME
1vQxaYVnAy0jpiRmrDtMJSbjeOr1vLPaxQJH2YQpl3uJ5yW0KYNwRSyzmJS7AI5/
3qRVppxBpW7DUHvxHo5Td8i/CiLBcZvXf2cD6Kazsi+G+v8pH+V8oz35dNtKio0Z
W89gcLzyysc6vjHRTWb/0aM1JqSZhvfjMfPhPOXkPou9RwSh3KfJo/NQVsjHXZ2R
pWnM/GfG4Fvexfwrofgfog0sZVySyu6UsJSysVJGeP03sz3GHgzfZ4DT3y3iHibG
/gnU7PC0dJgdQRe9tGFjOdZKRKFde3XqazBd2IRMljpn37ZYF5ku2ntDl8VLl8hb
yfzTe6iev6pHo1O+bwfigcxJUPGCirtFPdTdbWMXP0bmQoo0i0isewRXVoLCvRj+
N9trGPKN6lYZ1sBn2coWgJM3XQvt3laDPdal4c2xdIDYQMtH6/3m+2Ck2YqNWtrk
ZI2W8jZf576S/MOiMwkhiLyGd+KnsglYVcbz7rJCf6Z9OTeCl+4BbNj31gVSLu5J
9Gy8eSrAgwO04OEofyN9Hc0IoV/Gc6vUK03yREQhERH8eAX/TeM5WZkEn4pDc+wU
Q6dFqul5dFWvwvIu9CHd+CC1Gute+ilu+X89NfuSOonFz6mIhY0ZNNCGE0FZD+kM
veo9BAY2JMA1T979+7XDuu15+VrOGb3wpezgkh5RpS4pAY5QC9E4TsMBY79jT8U6
x6Lv6tfXs0z76wIrSieVmrBVyxavti2gM/q6lMCrFJlcEHQZJUlXhe7gmyHoALpa
CC4xdQUKSLmye8mXUzda/wmjUyH/UjaFDck9axz7O5kJ1BB30Q/5svYXwGU9cg0v
TAt3HBjFIw8yzE9KysrYZWcz6RntcOBhq1kLoD3XsjWnlNVH/iKpNnj1/aObbV61
H2+/gjmyBPTEXPoTqyQZ6dqIdfETkXnjaVinGy8kCStTNY7ndScjc1UXePMhgv/n
2EAmNuOMxcL+DL+U8PTOdLSXkdqBYvc8TSo0koRK2rloC/GrEPclGjaN+nCTsbmZ
lvsJf3xxResixb4ymuIOBhtSAPcY84FIMqvi8nyTrXiIM2bhY+l5w9Gh0ggsPqNB
kGjBAUO75yS8eOH/Dkw6Hy22cWvmWe9rEdjG3XeSUH0pVlSku25YC+0FOTxdLMiI
aGDRWc6lqrKjdk7srUQV+j49rh+7+nOWpiqovyALxLvNhHW2cZU8WvUC2w+HZ3hs
UJOksf4h1ZQvVFVVxSm1RF8TuoDclz9KpiFEKcdA2KLKuuEF/TQR4G4znayZZAe0
9QuzxYVhV9NXVqYmt3fP6MYiSr+8bEWUy9qwijzAVCDLR2kxYeGFAzg4hA6oaZgV
X9sjztPPGMHfmQ+dZnC7Y61SiDhHK49SagLC6yug0+85QcoKNkwLp8ewhK2RZsva
3zSbcEhTkEBIp1Y4Q0ectqy10MJQ+l2W7J1SqF0upAgs3hwF20QIedyxhJmG5frm
BkAdK+1q5cffabwtKzbZqakH9YIpDPwT0pzAQ5hXWwUMDOpd6LftLCOqiv5VZ21J
w0bzre0yC+vzc0GQs/Rdypr7upsEoblGl2dVlhHHc2M5YTpAD4yjqDKESsyv8wnc
Di/ZFZEgJH1Rake6IJUWI5D4YZekrFaAw1M89MQbsnOs+R3l7lMOJ0XMhK1ssWuj
2irEsa9PN5tg9eM7jA++f6anlktZzAWKerkXITys2yl/Xn0YqnTMToV3dF8exHhI
omzxZpQLBKkiyyMYqWDOvDsRINu3cHv2rW5iisv09wjwn87c36bmXayDP83EiGGY
dct1coRCwPOaCVxL7Pagp4Q2mM3omr5qWtPvg9xOQOcBgrX27WemibCIfvhj6kJS
Xzr0REbL2UdX4PqG7KYr3/NXodCMlQc1eU8szA5h+Vs9STgmpfxFkE9nmYKewxWk
naG0ntBuiAAY71oEgQoK8Ab2xUjJDkOpyTrOPve7Nq4PvIo60rYzJvesHPJdx45L
ae2p+tACkAh0jQ4HvCUlL+7YpxkuwXxDrrnBIHPM+km5rBrfHJcldY0iv7qo3ehf
ktZJ3sdfuE811/8fiGCfJo0kQFa61AdEietb3tx4xOe0yZ2sY2foDztWA09wPPIz
UK223X8Eew0VXhBJ911jBPuSzahz9UPvP0e3uxkZKSYWWL/zCC8LPSZ6t183GJyB
uhafPcb24yvYaLB4fBimzDqx3vOcpB3bFuj/ZezlNcoHQo+57i7rRQDJjfevA0RN
/nd3yNUhk597tfAUXxIbPczPrRY0clvSlYqWCvIB9C5b68ijB9dhUYRfP9Qj6YFX
kDa5LOCPH0Xqy95zUyyt+VTHDKgkdSt1Pnpi6S4g6xCMMz42vp6IzXiSrjh5H/7n
yZMqIr3IXIJC5BVC6jT4yICcqJP4cdXAEpADQUivAZbAQlWoPFiooW726wzu5D8F
Q7yaJ9lycz2xigcwgneAlhp6bc2v5mGmpwrPM1HVQXCsbrmiNQvhfEmnQ5DCuGIZ
9JS0BS7ei4TUt95Ff1fDiKR1eg8Ied4hZw5c+jL7Z9ccrpC97+tnSeVJ4t1ZKW6S
/fsXoyORFqVPb47mAleqzL3PGzoRK8euja1qIzCOQue616Cl6FI49GJPxIPlinUy
eorcJ2VJpZDSWCkvoPsediUHROmjX6Np4Z3G2O/JzsynMDvWkOQjI7SyZR/hq3LU
OGSushdgklDgWBqDWahcNtgdkiugsiLS0vUAR1Rbnpx7zpW4rlqxI9mpyEWiTIqu
g/sY8/e0pvmqhdmmNLnYfnz2Hil4ELKcoQWW+C2466KFrLczstEQZd6rr9qelK9Y
78IVVzRIhjQDu3f58EWB2Gc35deJuH2orJYGFQ9i1hvs70CG5F2J8W/Q11VDs1FU
uVKY68KI1QWRfVOBzVbOFdJ5oWKhofkyzyuP68JuNOB9IT1h5rX8vD9MYMs6d2KN
HCaAgzxpqeiZvHFkEcY/5dPpx2EG0VLX17r4wEuadqd1WEvgKBMXXC8u6AXvJ4Zb
aCf00tavVk0L0I+gc6OIgJoji1955Gg6OOXPpxRmMSvHvI/j4LX+Lj66Qd83qvXd
CoeFBQndn4I6zxolR7D2URZzMITtztQnipZdbXO5Op4JEFYk14VfIUPWMjPgiLDW
x4tVbzT3n9dnRDPlHje77T6Ia2dzecEPwi5EFtMdGkiJ6360V8oLrXTOBg1JSO6t
rxAuIn2KW1+mm6DEVH/QA+FuzrRRSIjWecLpRuSnfl4vSGwaX9owd3xUyyoKraKH
zFHjjg/1V1Go2/A+AgsaKGDA020/julto8DE6U4pKdoktQ33hZuzVvwFsXqwUB6B
VgaN5sGMxvXHD6XFGf/UZBPxjaCQrZiwY3kd4wDeXGGQx2N6TAiaqeLbkNPvBHgI
OPrqXDS28X2n8xkIpS4g1Tl9pOmIZ2Px5uXJz/bpJ/f+qDet7ikdOGH/qHjaL9ut
lqbT9/iWltH/ofMhB7zTfaljxaasZr8ecdKUZ+7IZR6DAVL1lxC6id51wG8gTjeu
JkJ29GP1pxH/DrBzLnluhstR3tEEQNKjw2YljcpkTZc5fj7kU7Py1OI2QV1ANxU1
ETreqPaqSzvm/owdGceFXtaobDcaEaGIwIWMKC+8mkgN3JVpNUaYbK5YtOUGFybx
+HbBTsXcce9UuxXFKC2xAe4hEsoPcQ2nVsnzomP5nKecC5rmLra9eQaDpkxCC60P
IUx/8JJuvBIGw5enEekco2NBZc0uohJt5cxL149QgGrJsx0V+k7fEt4tkWACoh9a
pKEszWgliqKZQ6cXXfqdMfBbv6NDaqItMHZtXtdrB0l/Nw4cxZRTGumcsY429mg8
pvyvsp0n4Jj3h9vEzglB25PukHjYPrOb5tgfcMNTq0f1Nljm1qAp+BVGeGxhsECw
KY1NwZNHKmmnA/uIgcM7X4K7QOMjKRen6rikCbb7JAo+z77pUh6cUCyBriS6Vmha
Ak+c2PjVXX47LnO2KMD7oKDXC1MxoL1L2TTV7Crm4r4leboQzNTa9QX++ZcIKCJe
ioXeY2ZQpysXuA2Pet4l9/tI14CyCy7vGzYutyCPQWbrLujv4y3MUYJBBPvf5Qzy
vE9DjETFUu0vFfmRBl0vnjR6OpcXs2EEQN2e/kTkR7C+RFN7Fsq/mNpbfKOlFrT2
d6+pVTLOO36/wGyDDcFWdivW7OednNxJ3TdxR1dddBLihRN0OfwbIj/lnUnNSFHd
1zRq/gqQwnm+02n/bMyKtd8iXs12OYLuYGiavstai/9DA/39oHvuPmKIVoE1GfIm
iuc+LIg1tpCXpdDYMJvJ+RyFjmkGHZSVCbHBvuxZRM9AIAoo2M0BtY0gfvhznGjz
2ARL44Z1QUHJleWzB3N9rzRg18YlLLodl47XxN2zuvq8vkbQG1qWx41wDv+eV4Iy
4aqYsxJaisxepC7TbuL9TpHV9HeiQeABm2Y/nyUbfXKB0cIPZDT/dHs/wPKBC4Na
cn6QGgIVANeEunegNRvhsOplO1PZQqNxVMgJAOs/R1L2ZtFYyk3THucSqBZ61Evl
YARhKFSAOlv51sMZgjsQF5GAtluMROntvdlUM1xackADSxdnVqgtrM/2N/mLmZKe
Yzap9K+dw6jA6zDwhKMSuaqvWiSGeG+3Izc6Kmj0mR8KN4cbOPnqDkoC2PxN+eEK
M44cNM6E99D8O3Q9TCM94l+lC1OzSxxSD8RSxndHYop4M10C+dINGoftRkfyZTJf
zyGZ8h1RWBK6pZ3ACg9gdl8FB7WOO0XX75Wa0LvffXzojy3D+JngrpvGVMEzvnbR
eDqGYPO427Ctdg7DfGvPnRPZUBT943MggCutUbcP1kvEzecXdi0+P2WtRgf6AXCC
EB8hrnsRQQf8r5zSQ4dk726j/LrfI67EU8mCtcxAM8tTjr3nPsKZDPJpmMXv5ovM
53wa0XLPMSPnx1UjiWjFQYUiQ5MlEfdHHxwmkKH07uQVjNzZt3nA20FpmNrfEXy+
KPW4mHvu9Iqqyq6nnr3Qp0LY+pK5gSwYj5MngmBpmumU7RFYCcxVJzpRMuRgMJp2
Dqp+ONeCU+JOP8vo2E00gM1PExAPbaNCf6PrF2bSluI/UrVbMTqBr83URz/b2kJN
CsEUheH8JYpj5hAKrEbB8lljZDp/soqsVb+C+U/m7kKEUvXIcHMIngvXQ5hYXRfh
Rz41Hmf7i7C9224As8C/Z7VxvSELrpYeEyd8ChPI2Yhts0tbE+tWZay+MMM+tBFd
NMyuceE7Eqs27YmJUgJFs95Sx0PTy6JeMIzzCz4eoW0YeWzkIDt8NThVCfprmYs2
a5PFaeredNzEdZ2bl1r8wS0IDGEF1okyuuI/O+1Phpjmcpt0GeOxtHkIyrYzPf5v
kSBMKIaepttAGraKlXrhoJGP95lp1+L+7ELoJZ9MIz2zVwT5R8kY81VT4ji5oaSE
zbR9e9jqy9Wmr8lj9w0lUieqp8sWZNJwzuNFNVrbZJHPlzZuWqTdVPAqPhLNkH93
1T0pRtZ5fNsELSwKAEz5TCJfqH1cFcceFzgkixqgkn0UUqgWCHa+0kB/nHl8tJuv
0u9mDYLDu3ZqoWmHiKDbKaW+1gBFprZojw7d1vHK1eBEff3I7UX+AwzDM0ooVR5I
qXOgbQTKlMTgoi2kzhVKsfy4wAG2kRO9/hwBfGVj73zzAmHOBLI2y6ax+7A1G7/3
mLNvyLhHLQAw+X7kOUCdcaPzqahKh4SFZIF6VgnCnl6/rzlyQog9jWq6nRYEZtAJ
tbeUjVDuV1D+0/VuR8TBV6OEkAZxtm2VALqEoyb2zYDHoBpyEDV2+DGGn7ek1HpJ
xW/l3omiL2IGZc+wUSS9emjmwXd9nmxsde92uzsdyLGip9lBAvxpVgcHo46OoSmZ
rRwcFTeHt5bMaVhZbLhO2BICU0jVSIB57kokcfV7Ci0+pQ223jcMwICPXFH0k6/U
jRaMlN+nKvlXeTycUscFGCpsw/8H7M+CewwS/kkd8LZ3OloHR+wtlzqoeDeoq+Rl
Bi+uDYV0EtdiqlHqyeGQKjSIg7uuPusO870T7bIEkNCsC8qKoobMcHYnL5nMzgDR
sDc4eduhBdD6nO2nLuZCPX1M1isEZlDZZFFCzSbFw4ws3BwvA6tSqsN0LMGib6A+
cAiyN5s9a5iPaJsTh3xy0XE/wGt4hqMOx89aNoZXO0FeOsoZgtdzkIsUyHTHRTMc
zNKDgX8Q2ymZkZiofZ24BNkeGYDgeMlMRNJuocK4Bs2ixvpdRwN065ynsNv/oCqB
0WURJ7wOvtTVccZcotg0owPESokXLNLSef9mbuxEjKUkwqCdTvFPD4iNCWlH7vdN
gfWq+y1JQmrzOeJdRbrcceZjCPE+BBVQDO1aGK4b2Yqyh9hm8llMhzt4UKTeeEid
ppe7Yj+FNzvKD4moviuKayBEKvH5Axp424khPNjsvAFjps9+D+eBqLFJ6CrHStA1
8d2GbVD0k1mMt77QJzOfwwGuEtD/tqzoA7B0U7hhxi+pujcjWihs3pezQr/Uq+mF
qeXOdP2MnYo89h0RnUpSIt1AAHz09WV9DCYTWHZCRODKQUTbKpvffX3EA+lL74ZD
GlUgPJqgMqtCxnLkSJNNAC0GR4za329+7RUCZvMrLNSGkn3nsWwpW4cjhz6WR7p6
Z1cVcSVz3TavokEcmzS4CEQvrCorcbof+vTugwGgGZcS82LrGSGRpkwm7Q7W/WwA
ZhoIYHOBmPqKd4K61v9KgkZuZewfVlXkljrOsButZVUiIwa2hB73yJHKskoycYgY
b/Wjsd/SuX+7Bh+8mof0MXF0DZzb5bCVvSRulVhbnwEBdXLLWJg8sVe8ZsNQuJot
4RzuFSxm2rpLbmBkDQEOqewTRDh7r3S73ZD61iCMSb/3nu00bevCy8lp/TIjvnu/
EsHvoGYBHaiMSO7DLj3kUTpaDRtZkrJ1jGssEAkMaRQsOIvQGQ9YR2qkxUYCJNBe
eAVgHncLm+PDFLpzTQW/Pt5oEsLzT0Hh8XmR+C5xa1yvjx3pw/r5CzJ8ne4xX7zP
rxBcci5y6T6JNiWq8Ho2TR24aGPmG+Tn3OtoxAzd+omBAkddmAlx6xxSmMJgbC1f
iKIBx3QiesbW6AlZAyFlXZ7CvqcDLsEReLk8LFMfjPrQ6liwdCdtecamzfoJ7Zly
G7+nwxaZyfotgx8ro3X7vI93wgpjTETJgrIzY+NZvaafQjIKGoPw0t2CVjI3xNYY
WHnSkx75IUTsl75Ju60jeZPUCgoFFZH4Xa6ew6+Y5Rs0zJPVscFAXX79SvDno8ro
Sy2yP+C9Rk8NseDZk8o2azZHU8nXrWbwAwEG5gVd1WXB7Yq2UZa6tPiGqySZLt+X
mipQxQTnAhgX70L76/LSoIo0A7vTJbu8wqopirXS/VH6nnWlGW3ec4R0xo81fNTC
wo7jRleB0DNagu5bRQev53NoF5ardBiF64kXQzcxJ3N1Do32/Q5f0ynhhicefp4c
BPbtqhCvW0J+gGmk3Hmw0Mkxb5lj+si1cH5Pcltzo4CnmL/o5+GTKSW3f96M5LIC
Qt5wIVZ9f0vq+SUN9w9WPJmWRy6S80+0lcb9uZQ1DINVzxWqsVcLytn7FjcITITp
V8UYLK+Sve54kvUKRFyhOg1hK94ov4/UyR/ITi8k0f2hmuUef5joXIpML4xUWntH
G1CBILEeZQHdKmpq5m0JmUqMj+8RpWWPX/93TTfPl+0kCePiJhVdo1I6gWtTFJm7
9ho9JChmJGoYw1XdME5KpjuK9t30QRCnFdAxqtYAemNe07fX1EFS5rFoLNpyTR9H
aO58X1lPwuWbOFf1cS60S0Foeu+S/8ZMUp3/ly2m/CEdXiM1haUY9Z44oT7HKRwB
czFeBRUJkj6nd8ha0nXX6YkB31Q9d5t/xMYXqZOdbro/2d8hOygoAmbF1ZLlvELJ
C9kGZFpyOqwSS8PVvjxCWUkrfhqh/SRNsGCZL8/Krd6hNTb46vSgek+Ch8+YOG2u
vz94sBJPy8BDHRUCs4Px31ut4sgoWucC4xu5lAdDpVxQJIGGp4KsWE8uDlq8E3+T
nxzaD7bNQFwfnUYKb/WXItBHjsjn1E+Qrl8PAVomJZldUIhmc4te9toK+eIQ6NmI
eOYZS80eoSs3BVYdS6+OrTl6ZqejugzpD4G9hq0JB5TvROZucxzZfiLmY0aXnRvQ
YIE20jl6ubr4P86A1/JqqDFoFl3S8mMZr6WEiYTiWjJdTwF4xtJtqdHpPnVrugjd
4IP2bAajKDCD5AyK2RSKRZ+d+ZfpBEW6hCNJXsziJ22PSER1T5xkjb0EznzyXR4c
O4+yQ2J2Y4FA8fpjAfPnnyJduzFo4Jp6T0bXjJbU4TcSsG37CVU6Y40zrQlqcE4r
d6ZnNjjn/4wHgkNDQAM1OiiaYr5b1zyaHtaofxndsAtAllReeRXege9DAZ1TO46x
H2L6jPMsWhA0bi+p84ZaUhAEkUrNZPI+4oShjMK5kX7tInV6yhMeiRs3dB/zsQ3v
ApmimI0Mvo1fIkV68Me9WMY03ZjcPsXtqxfV4W1nPYMqCnBVvIDKRWtWFgSwEuHA
T3JOi3sO19tX0A1rfUWS0WqteEcLwPp+F2y6wUk34eIdRfM8mjpzcGxnfbhEMxh4
21N/38kB/ksVxC+2Pd0aLurlg/m36zx4JLAqhL3ANH29jCdnD4voM9q9kjg4oHVt
4HXe5pSK4xwJVcWKfuGahSDFUDU44f/4S98Bl4iTc58UVACrZ4oe2Ty7gLSvpUa5
BetYFbOqIe1Km+zVyi2DjGc0SXJH1gSuwDAy8mHGuUV0lhHEn0X1WcwutBg5mBBX
/BhYIbYbEjLuYIevXcXmD6uy4BWfgNr63kgDCLr9QkM32dYnK8F5nSCixjnSAaFG
qhyWxvYQ9OneL1zdqeJcN/mIqEX70jc5pDxmhDuDzXQNG+G8Wrdw+gmCtGFhdruU
JIKvvc+gRy6oMv8zfJIp4ef70DneYmDj2XTI7jqzSXZjaTuDwv0exp3mufjhkCsN
pz88RxZ3OtJ8WvIIUT+bJ+8HEWhyBVj+VwyZ3FxiKGub3nAvEE0EUGXFBi94B7eg
HUxdpSk2NJfU+gzKKi/grzEPAq/GNVOjbExfyoeqstZ94fD04IoLXi9XuzSfpMat
0a9R1tCbkvpt0yq8f/VCB/h2C3PCHEgPMUBT6MnjU0aNJ/pbO4XkFr1KWBuB8/EP
QoFHz81B/CFr407wJuEny+SYEsScaEjh0EOSOXKgLMLmRi5aKA2LF/DjHZLSI3/V
Yjg+ziEWKH7HZxN55y7oBcrLtl403NW/DHiNgOj3zBkUIasFRryQf1Xp4ek47UZ+
HJujYb2P30h0T7RCmczLZXaBmO//M0n5+5p5kxQx9QNopnBDB+i/DtaS/oew+Wxt
G5fGXYcyBcZWIhbBV46DE5vvfeY1X5+w5lkQRTcHxRlR6pMeq+h3qBerXirB9yvt
yP78sy2fjcypykO7M1as1EZK3ing0ZApsObHkZbeFX8URisG5lt2J65WeyTTh+Cp
JItwbWHRT8lxJRtyBnlzVePsyPEvukYm7y7SeTCoYb0bRF0oPBMOf7SohSyjNh7E
+5chdTwHiU4JPHjLNYMx75Q6nkrJaFZiebhFALcdgSc3j1PCFOOQGXE2TsJf0Wh7
W7o7PyfflJp1JKz5R5g0A5xjGR1fOGx9L+KYFZYv/1ZJ1FmkEXbuw49dfvoRaod4
vY4vXQbqgzr8DAwe8Ln5RnGlgXA64p/aKLUzInQwx2neTFqzShq9NTegLz9LlIQT
88iv690yVkwRxZGX3OmcJvCGo4Hy6R7yX9Jq0Sty7iwKdyQMoNIUxsh6ZoWY1+1+
X0HTDVZ3wyBCipXmCcfWd4TwmjUHkPhpUSS3LnTj0VZXGuyRMv+ziL4u8osnpVWU
j7eQpuxG2TzRRJdqWtE0WGy8rp8d4KrIXl/hA2/aUHzTyVs8iyHQKlrrtlNeNAXx
Q26F20Rr9FjpeDD40gA5vZcLmYia3eaFhHL6AZOmUJYI84y6GAMsBGCJ/lWxM4OO
0Jqhd3IVKqe3La6yRJXwfG6/hvtx/2HRWlxpEiauco28QNlehMMJ/2gvWxWlSdb7
p/b/vl1mHkZHlLype8xreHOZpJTaxb11Yb42sTFByoaENvaXceKuForck3HDV/2o
dU0dR8EbH6RptFllN8UmyB79xgiATCx+B+kk7g1MzQeYVIrWrZuritAhqd9M6Suq
AF6jAu8UnNxBGI2VHaXLK2BN8F7EWIW6EMhhn/IQeane7942xk0nh0Dgz/PZs+KL
jGtpAbZlcShVaGC71k1tiEMF2tgc7KiCm1BrxAPT4QJbIKU73JnEn7J9DmAv2kSu
pFpKtXC+O0qmD44DZcDk8rkAmevFe65jxy7uYodm+Dl6u+xEC1I6xmYwSdScwRxf
MyEidpDtqvGZt5QvKEPfUx2WuzCmUehH9hSCctBoxOTC015CgrWZGvjTey8hJwLZ
CGJWRFxzm10HW8DW1Wd2CfgNCXFwfTr62uplsfHEVx7cf10cuULCFDtHCB9rLjEP
ibwYj8mF6M53AIaAscnxBRTHRI7B3Oq4awVt4ILTtpRdKC5mdc9FqyP9v4Tn1pgo
QDP9nne1PMilL/0qWGxT0Zod6l9pXv7bGDnYue+k/ieAGiidXeheXuNXuc3q77Ri
ye7LQbzSqIyMTiCnV8/lg4d4QCVC2tgnRJeR60Wygkw8lTBKozFUoC5r1lK6+sA3
1y4qrdhatvXkixSdv9rEwQ3gED0nvTuyz/BXaDkG9c5QlGeppmNtN3JLjWvGQD4h
doGvuhc2jEwBI85FD+7GkJw2xsbJfD3fxRagWvPI7lD7hW1kGeYveHx105lyi3Xg
ATsaveMLBdbg5GLLNVZc5GseTdGlsBghdZ4Qo7r/cu/A6tYQc15EpA2hzyIEc8F8
E5384ezXJoWmd4NvdJ3PjPsgmRyP141auklvKjuabsf2G568lWRIKucdkYwjzcVy
1QiWBrT2E0aDynS2O0ySQEKIj/KhaFWComIy9cKz7Bc794J9KPl6hZKiXf6X0jWZ
RLD2+axK6hbcbA+oTRvfDdO8QhGk1IMbUWQKmatGqqsjZr6tUTQeog2OpQ2UG/Jc
nFE8TQYF54bwzI00Lc4BjU2eChQqdiwiIFRoYZelA4noOwP0fD4iM74cq13YcNBM
Mx4r/FiTfynzqt9BeifcPmOyYHgC9cOtMfTl1PrPOA6xBGGPyxNgtLKfFzgYBYXK
M5liuuHyGAQ+BrvCM/vQtFtwWH2FV2eUg0f+7KiXjWkXnYIUwtYp8yM6mD2ox8nV
Yg8dR3pzcSUiltSA8GZ8Goz1oBHR0Y1jMVQLN356/zs6V+FPyErdyR82VXXEPee1
k8QfBZRvAf5GV0j1JqEQDzAGVDhUD7YlCcRtNKLueEmqfvTYt+OMhsx9xwTtQR1J
Wplfjh4oCxhhlE2tDYCgynTBUzv/GaJ0DzYWFNC2z0kGWm2myGBQQmHMluOajpeg
grT8MC9+KrrU76zvcQXZ6x41tdlylvy+O1/Qk0j942dc5ns3nI9wsI1fzDV8YwwQ
1Sb703vMwNfSMObI8+kyqPtIWuyGyYiZkPzXh1216hT3FHSWYe6nhRZJeJrYMr+i
oyXCORwgfiffHsjG0S0AC4NuhsFa6CtYqvExcjkqgIfuhMDNyKBsagLS2NDhmLra
dqYBr/ac91jBs+LVAETLzWBWnpTq2LdXID7BMv5hcYZR8sErbGbEtnlYalvorQt5
jrk285T6IlQeZRkVuA115pSZQ9x2qcWXYxct1t4URtpODL99OsOubmcOAtXDhxSK
6sHHzaSuC+Mnq/zz9lHbhHNhVlxT34Sj/ox0YZDR8KI+0QXd7jeYGkz7IplU+OUB
VJL6x+4drZx4HmYQwGC/1h99sAvp90YSpS8uAOf0Mra2jbsxwplR0Cjz7yWb61+E
lOZ27bE9XE1w+unXtiUP1Zb49fw26a4j4MOiJQSsrGbuCNHAPFjHmQDDcWoUWyp7
3cYRK+4K0LruOrq7eAFdKEjX3uZWedhnYOE7slNnlBA3r9uKzBIaHK6WzDLMJ7bS
CUOI3A2U0k7AYhdahkB6EjKhcV5oaaV4RoMyftTCJW1yiLBBAe5D4ec8ewvR+ok2
4+vSi8jDsQo6zxFvVkg3bG1O/wUfuk4hZAY37i4SFHzFK1J4D7+OGeZs/wfKFni8
m+EeohquoH/OFerj5LJryjXPrH02ASepVcUaBnMz6GJlzZmYJ4of/AIpkGV6Q5vq
oyXJxx3bkGElnBapdNAyq7/JgsWU6W56noqYhJll3CRE5lWf7Dj4i/YbMn3oHUqC
Gr9uC7GxL9XCAiadlQGSMbY62fcx/r7F4VAeQ7R2ig/HMP7FP3MNjbekXifIRNFt
JZuKivTHfYzMJFUrnUgN8pQ7qdVhIg5oCwiVit1V7ZohLgFL8rvuCcWG6vHFCNj9
Jxg4325EMyf3xfmg9RIJn42Xhh+08XdHF41ZHJe+92ozGYF1HCqBsgxQ+RPBEgko
zcKbc9PyjYWHiH1l7Z8nd9iyKjvL5nXDxJHku8pt/DSxJEHio1C47OSJ76JedCH5
Hsq6RcU4lHxpZv+xz3y5ZmH90/+f/H/s503UWoeIcItCrQ1IDjRR/X3zWFwXqu4e
1xn7aEiB1zj2SoNS2N7DEx94scCZng2gbKEuI4t9DsNmf1PaDhU46B57OUgpSkUh
JeTxq4aI6//ehrwUNYi3ncu8diEp4d4Wa725jOr0jJcZD6KQ4SC/WjbpDJ3VP2f1
zkR6Z8AyEIpukXfQAmJCjGpQELVpGON1fb7Athlj7YFDf5ip68XKlLYfBRKW2c/u
j8mdvFzzfoj7M48ZpMXlIcW8xNxjMFYwjkGlh0/yWNd1xp+Hs43yWvPF3cOB7s5c
JAGwvOdTqi0JGIvu2lxNqluoHPeE3Vsf0qTQU3TjhDHHEBNbgndN4FxAi6rpzydA
phID9Yk+oBASqnAV+SF6mA2Z6YQfRErJirSqzDNfNEo1AsJZpHGqgCBBZ6Kvsbrz
Jz+Lpz7m8uqgWd9TWcJFMal8tnTymInQJSfLDUAS/hh/s4R7W8XEcIOCO+PjWISa
oIli1PFIraNcLMXc7MAjHzsaBdozE+cfBn4MrBUpv33lWl0Yl7lM0uX7C7SqJXgJ
5YnZFPuugW7JpttX/usH2P8mAuwntKRrHQP4HDh6cyuCRlWCpXPS47gPzI82e86y
e9rTQog4gBQRDMu7vgyIU45hjHUyS3ZV0kG2ZZbcjHKi+pjxRTzsuvzbRwyudRaP
kxVRPKjY6wxWjbT0l5kiR/zven9tODRHbH0q2BoE1GaaJonywGFsCki3gisNqWLb
E/ecalK/OlfhIyA0ySF/d3mEJvUvr5IvlP4tUOCNrYOOBc2/R4h9rv6ux2otCWW9
eUKfbbxvMH31x3iIbTmeANvQwGhI8N90UM/KANRHPqfIxEjnaddPYnUeyX7vBFrd
9XAthsD0mVEGL8/FQa84J54mQS15E4oSWIfAWO9BYnLO5AcHtcjhGMlVtS94NufT
L0y364XcCwEt92djzzH6DYB2gn2JIdeNLfo6NgcTMunvTkseC7RErFj18FfzDvUQ
caIqvXPlK9AzAjxq9bFZesvkWYSAGHFeMRieFl484/PVZKSbmHFZXQK8UaesiI7H
pf60Rboq4q4BMej+cpitZnXjcqszqHfNZF13nXwHSUDYBOQyFOrnqQrveEJye/64
XUiOH8dso5kd8m4SzQEOZk/LoXQEPG5bkgSXCAKp7oPpymKm6T9oQcmW//ICMVfp
9pdiUqcHcTZnPck0/S091H7oHYkSSJzsdz/DjlD7VQo9MYPUYKG97ZVm5gJ2bFZq
zsdj7BDKmneMgBund/LviRCtL1y/ppn0RDCXz6XmwL+6/O8yQ6IHBG8ZOdMslBHU
9Duo37S3439ZSer6mqkiyfO6gyxMCQ/yje2OffcC8PlgDAL80WhfFes4MIZJsUcY
xaCREXrgaEpgjeZ28XwgnUUuNYHGDvRDbx0XoEGrLmHXgUluHUYjOIcPc4LpbSw0
quEHu2tBhHkjcy8Td3wSuSU2dN+NIHdYodiHOHHEJtnbmy6VPF5/CydGE2utncA+
mxGt5QSUkQVJbxE1bdyftkLPLsuR3mK6z9rhzxYVzkju3CmwDiU3Rzpb8OofnkHd
CpamWihKvZq7hIfySg8bxcoXqvQiLylsxSanYe9IvQ83ZyAQOU9TL32UzWgcOtuA
WoGF+Y2PJGpAqBJ7wzYYicyFaQNfwAVsrn8U97gyXXMLu2gsXIaPAfdKwAHU/x3x
AnwE0ONCivBNzZus6CxQuF3hxI4cOyMUzre8xrfllq13NKMy8RXSlz+148LkxscZ
9RwUpdCb6o3yYL7srDhpHwrIl/aqlUTnYon3gWMm51LBQW2y+wslIw+9MTpcrGhH
pfHSmv3h2/qhNgt4zkoLhOZDiffDjjU4ipOWxJ1Dt2eDafa7jwt7QWPwv/w5QLAA
KimzbUHL+y1HXuw4KxUS2JYjAtn2l53cKu3DOniZqI6wWlzOhEpYmnXBdMyByDlr
IkeTU6/CTFKAGM16bbr+enAcZASB5RoiCqjEI6yi/bbZSd+F47ewAcQmBKgEZosh
8L+6+MQL9spUdApt9my7CFHTo+MynsvyCLn/fWhUfaL4Oe91K1+JJhyFBw4+ARw0
Aln1eSPm5BrElylyp7sbYV5dj+W8ytwcC/JibNB8LK0QbqpPC302eZykt31b2eMV
PaItd3rw0QeBVtFVu67KvyBPOFi2ZhcDdpZRrIt+ZGaeVyeZgdBjWWJrhOD4VX3W
CZFq4LRFnSGCEQ8ktiDrH/NR9OB3tuYUw6I+qftFDrzBaGAbYmeBkXN48dYfVe5M
9i+3uVrZhppHA9+dXK7f2HOyL9jCF92c9sfgmjJbJ1q5mP5eaPLqm58q5zmy/wLq
uAg0WLVBZfpV5xyv/89j+CEmgIuveF0mUNyOlqRAGk7w1pj//lPM9vFhLwMoJNGP
pNCi+dxuXFtOxNG0foAQB3dw/uIjX85J77BGqckDDBLmf3XUthVfSHuDPQORGAz4
YsoWk2V/0id+a4CKb5AkqozJoF89QbKhKrB+hr0bxad/zsl2rn83v4nzUYz/G9B/
/6vqj5SfsCaNdxN81HhlGK9H+rVXkx1GEhZ65Z4EEx4W947HA8OjNDgwIDf7yzTb
IiEXgvuC58sfrocYwpcjV6FoBZ5P+7XHBAbv4s/BNaNu1c6/hNOdKgHo/y0LgDXI
0q+2e5GibjLsLpo2KYC1kva/0CAkl0dpQ+oPKnLdxv7UUujv3RTD1R8iQA+GNBcw
+TPdHALPni/NX/94hT7ul+gzcilSpAVmqp+ZPSBApkP+Si2wHSxwftRuxmX5yorL
gKx99kjd6xPO1PKW18jrz7PA28cwNcAPCcpoVl78rDCyzEX5YsizU6jy3UjFaLEk
FS+LXMUQ/MH4u5V9vZkbk4cY7IrgKT0bDi9SSdkK21XvlSPo++eQSzoR7Cpm2XOp
f/Wf8dHHkWk62lhB3/bKScXH50J08ST+ACNpbDykxZ0gEFi0suFzk3h8AJXI53w/
L4uVqbknMXaguCRkP8tNMxj7Lsll2kWQ3b/0A0qlZ57cOZeRnH3MOx+/pgt0WrCj
gf5+tl0MuGfPuZ6FJMyfTvTizjKgycz+/9F1Dslunpku0t9mfKgzXAB2nn9vp44q
dFYrZlnEyTYBmkpuAkcmBYcUKSG8oG/ji/jssFtfZtQl9KSEXcc6JmPFTra2cgt1
PUFVy/hwn11C9/eAj2PnwCsXxJoQgIa2eJnxG+jeSh6IBV4VEY7CN1Hgfd2a23Gy
S/jsd0ORtnOhnsp3c7vZdaWNB6rbIvpu+bieKfcfS9xvFEAYhKxV5UpkdNdYi6Nm
46OEV1oKJoXEZN4ZFjnyvQDkSZKX12rTDLK0YVNqokqTLsLSVuBACByXKD4+pK8X
0sLGxJTPIqHSd4XGKTXRTdUhu55PDWrsV9DDtPUoZLqBNrAEObaF029zrWO9DUVd
GT0tYaNO4QMUWUmlCxHM4lHKehaKRKjbP8izpm/erG30y+bK32YRMSQQsvEBkd0R
Q+fHcwIBjBXQgtJ/IMipKRDTSpZnqwtMZj3rxXTfrgLLC4u6FEBe22e3/C2+qDP+
qwxI8+FkmbZmAhWU3NE8ra0WIOaZFMfh31pRhO6m9FVwoIEscByJIoOApWzYxiF3
JDj/n8+tOk39/C7hj+vISN96VAXJtajE3wMqm6QaNsp4krC7WbD6pQQ/3r9uDf9M
+5zLRK4lH/SB0Py3zElHZ3Ple2kv4xmzWthyK4rqMl2aRarzdwTqRQR6DEKsjtls
xcgNSzbOLxRC8VcrSttMJUeDZkEJIcMFrIhI3ectZoBKTAzbtvEPRLZTyNnjaYQv
NUjp+P8BX4xfFAPus9PnGffjxpJ6sDV49f30TapUOjUTqXtCVBAj3fIfpJbsWSWQ
qu9MHB1xJ4SlsmP4VoPhoN3DK0srFded8hyGS2ZxsueO3CRIB36nlweZWdvPjcrG
3B+KY+AIyKA8JlcfQzTOUzzr8RKorHoJ6kB6KgjaN6d0cQqM65uWs+H35mFK8xI3
8zE/Z9P4oMqn6Dtryn7utZcwMOpxe92O8VT5O6hWPXi4W7RfgLd65J0JZvMspNu9
ldtpsg6WXuiznSLyuJ3L5H30MzPVGnHEoImeo77wToqtlxBzzn8vXT6WoB/++HC/
zFBfNfRsFxg3D2bfy0epxVq7HJVln+SyDzi4mzswAjGXB0YYzz+auK/FxXFT4yXp
iHBucM+pS++dn77g/8WXpU+1qGytG+3yU17XrYfV2uxWWIWSpi4Qeyllv89nE+3Z
Fs+vbukkosuzfivdR+eV5NSyXzzHMdXCVvF5/IhmT47z/yxh/Wri2GKsQScijxAX
Q7k53qB2LIt1+fyvEB3juswc6jQlYPvaICGOLa8W2m6omy/LtoLHerM9h/CV77jY
n5yNg9zYR17YVpCIgiPdKqSLofszE602nOtg3jXAGWylVGAiOHGVo1nICs769U/z
ORl7mvQehyFhcEtbaGa0xHys47Ze8Orlx9Bl/SJyppzpVObBHI3imw23pqupvcJq
SkIP6ZPAK+tJOyh+ieh4HL14Fj9cOh1p8PfR2kUZQTfaSTQ9tekrro3N7Tvp0CYp
tiO/YcY+VuWMOPXYivdXxHg6gaDzOShkK6BmJm0n24RTlMnqSkdGo/X5YMS7odZo
9ip5U5km+h+/KSLU/qNo8jJiBBxa8q30QuusfpCSFFF+6DMsUUCEL4xrTDjTRHk4
Ao+MNksz2A+rxN9XukjLFdZ0Re9ggZog5gVb3/mpwQcfEsh7wnjaeVNCLPM8wMSx
pxKLv97Hv8T6oz/sfmw8/wGfUqIUdQom8DhYy9HejCMmB+yYGuSwrRF3Oaw//YnE
Ya8K3ZvOWZCJwWnEuCZbHW9HrN0HO+pYQ+wgFForpryJJBl1sbChhFcKRFChzeBg
rXFXml9A+McaR8ppZxEqf58m0HZWvRGJ70yF5Jc6dI20xpXoUzT0MymoS5od6jzo
lwpmFwU28i+az3MG9lL+jIIM9TSspqaSc1r6XNFm1dX6DUAQDCD/C50Ttmpp6H23
1fBECOlo+ncubjdy9jA+Oq2wD5QT29FxpO2VIU0Bbe81Tv/9A/IOE1myPxeObRIh
abDUCebKa3NXuAJsWtQbg0NOQ+fitUvnSzgR1t575NMlsS6v5BzuGMMdd2pLGCGx
jsmJKEdOG3T2MewTWM0mnv4JaYx4sNlVd8ka2HsnCo6Uw5iaGkN8szNv9Y0u3z8k
uPuLsT1AiB3FgVsWr6RcfrIOJpnTEMj7azt4zNGzdL92mf2ct4Hy7YyVwtZaanpj
hw79nxAO2t5VwZnu56j5KSm2PVOBQUOCZz36w3Utb1tQ56f5PlVmTyTt1qF21oZv
obbLZOBKxyMAxV2r7Qk6Q0uMj9xNNrAuyXfBWMbQBMtFAHj9Ng3QnW7KDAVdsjEo
SpFNDwb4dylE/bz7Y3mg/+PsQ2O4Pb9+C+pme61+fnCiOi61rQJTLBF6iRG9rZXt
aBQQMNDU3gtCiSCM4fAC4lrRYpUk9q7jwVInbnBO9ycXo5nOODaPSr4mwd9nU2ZG
OU/9L8ETXAJbMeCNrvOAiPyvOfqWHcrmYzXHQZzPg3akE9HtMHJtPZCOjZX5b6Wg
Tj3oyi5vLh4/RmuQ6Ve3/r8Ql5q05yFNk7ufBg652IpIj+snzldZbP0Fvtn9P3I8
pEFNpPjwY50HovM/HpXBWHycBbnKm3IkVU4mv75jSKL/UfvgKMFkE2jWU0fw76Rm
z7lVmHXXzOfeHmhAX30tUUvsiMeqrnlnNzUsTgt3mihUpdyvuywDNYGKGzQTK5GX
oj0TMvjxeV7IBT8QApUChPVd5JKD0NYo+p8NBHFAweOdW/vXNmb7r6NTy8ZkeaVs
c9yyLk8OG0T/jY2ZWnU8yi4KiCfReShCcHOiehd5Jkmc3BFYKLjidA+HTMheYxfC
5UslGxiI1A1R6DsUB1b9R2qUNP0BR3trQUMi/wpYzSuBF/JoWxcOIzmmTVDWkQax
2asxGMZGcQH+AOMSP9IBk4iRZ5XjWnHulz5c+VcQj86cWlCFA/n+O2ycPIDqtVWU
m6S0eIjYQYVcDTn5iYurdkMFp08c4501SGflBEqFR6GMOu7RbX/IGPDWw8TsHxjZ
yU4VxBbGGjG1vqNHzuhxXyjsV2eR3G1z+tPq5p+cBMQYqsRmv/sFgfZkBwouBJjd
5VKAit1CFQktY5AzoCNennc/jdXDrP0gN7LN3EUHDdQUkg08U2Vug1eveS4eNQTy
3OTMTSEN7qa2tUevV0Lj+Fol4PIDbJW7RdRYm3BkYjL6dpJPSqj5HKA5n3YToPPw
Ly9JuVjsClSGQ8tVmG5gUujcoeyojVIp75MXWuCP/1GnGUhJLQvxzGASL5P0+oD7
xbZ9CIR3peOdlAEkl2cLYOEN/oMrfqKnAJgB+TMgr4bQd1/IzhXbzKScyrOOnaUU
G13OyxDOazohIcetAcTLx/XBiZIH8I3R4JNNLoHqafXF3WdRHAOjFo5YJJ38cFWF
7ZFxhKAlTdVr5wYgsgEdoPUKscYGq+p9+RikIAZrc9W0aH2d8Ykn7HM86KG2RP/y
jqAwKRa6TFCgOU4DhNrrN0Ywh7mNWVoAcA2E7qVZFd2X9kAHFwdPV5vO8ZnDmwLu
ozdYh+qjYFXkbAd3TRf+nHut3AW+YggPQwuS+P/yY4ivhihXbF4AaTaKlyDewrS1
gbPbVu/YOv+Lpu/rvt2VT32qezDiv9/77M5Izp3SZwW5LPpHD7aZA13al5OVeAJf
ciVzv9Jl2Oq/gU9rrfJg4cpYL42yEWty+y0nxKg7azhhckxgXk3W5SqWiCUefA32
FC1q7ogXJP8A+L3JiKNcPNzmaUUgukfY4nekkh6tpo8CDVO8HToCjedeMi0RAeHq
krJY4C4R/qti69I9E5ULPWBcwArVAfHaQ0EHLPQ+XE5Bo8oNw2o7gsgB+9OHb1qG
ZYKDi5jSWDy6C1SVF177ihwrM0fl7padQloMiz1lPSYvyZIFSCNytiysIDyI3iPF
UOsv6n7LJaDGeAmnK6hWf0/N8+VURXi6vLpqcxNYdXyXg1ldegzgxhqOB/8q+Cdh
KLmES2Dp5fslCQGLRNCOBCoqzGM9Z2hJ+tW8l95fKhG5R5SSep2gZYM6CUZ0JAWE
1TfBz5qvnggUeKtoJpoOPHwVx5RyC5gKVcDOvXKQkHah+Dqkg1N7P2656uic1K3U
aA4v9meVBqzaCXCMWpWLVSjF9BUcB+6Vq74LaG7kcOKuSxP5qTrQR6HlvrjR/OT4
fu5xaUOGEwaTr4vjyyOXjLvfg4ASe5CcywB5sTQL1DyJjuIbtmRgp83LHA+a15hv
PT8qq05TWLG1jG+BoEZTzqCc960gNPICBhr2BFsg9rKl9W1qLixIyqOYVV8P54AX
X82rPad2GWLYuJQaZFnbEdx+DZZISQVvRt9LKMNYc3+Jq0giCcVMAn4Exkj9xKOl
Vt+RaYplIF5QB8S8xvsFRZr7XvuEbaef3Md4H4SZDuVBFdJq7lNejZFxO5XH/C5I
oGiSbNK3x2wSRbwTzntCaJWBi7j7sXaSg5HpF/l7n/42QzA8Xulk6B0UsVbiPoG/
JlGgAQoSp495DVYLGpZXEohqGQ79ZgFWSW8ZxjzumK9h2egF0br5YVkmzj+6DNlY
pu/YXIJZkIATz9Ll5kixOtAI8LA/Kd2ynoHrZCBsk3cheNI896e3FdKV3ITqkNro
NYwBd480Av+Tjvyw8rLcl2/cBgMVF01/yLUVt8hx+tCc7xo9fSfmJUZ7f2c5gScV
n4ZCIDMuywy5ls8RlfHsi4T73sY343KD+lnU8RL/i8ZxAac1bDiQew43JOBfki5e
+/Cy0oug20oSDGAod3ZXWFFLJuCYCKB2uI0weKckEApm2al/ogv3c3BWZy5FjH1K
Tk6BF3ot0HpPWeCfeMS8FUb5+U1CmMRtHje1hyYB1mPvyNps1Xrf+ZEN9VK/l5JT
NtNCON1jDUaUgWPeuwywq6/n1JhnJjlNXioQH9jtzS+KEDa/fXFccFvswXWe4clJ
5aDNpxjsIDxFMG1GxuDCmeG7y+Md1LGpfrL0Hz3LCB4CO2uxr1p8fyP54TQESPxr
G48KwaQhWJjXh/kHr7Ur7U2SeeS6IS9QOnLZGYlVjFLMTgTi0xQjgbKDlM2ujREi
n48RCS2AQTE5SU8tv0AFZpWjs7dukrMiQS9l2GZvBS/5qT3B7QHQPLPjamSmZ8fW
i5FhGyHsm+wwmohU3dvtgk9QwAKXX7qri7Ax/3veVzwNemQildUCylwOKpI7/mER
Lsv1J7b06VT+yySUBO828pf4PwCSNH53nHu+gubsCyo1fi8p+a6vPsFcNjrm08Tc
w0zshYbkOlw0HrIm1X8HybmjfbiPPLtojSjLMmQS6Ck3VelmM/fieyF3ewP9iPKP
50GrMwiRpU8WV1hn2ZuC4yAvec5/e6EkD0xN5eP4RiDNbTahwRyai+gmylxhHLnq
8+17n+KBawvw/99V6BWXvwpzdT3p888FI7HBCy9+zIJjwrrUn1BLymQ4gmRQQ7ce
5PbPVk2AcS1sO7v+dMVEFKvj4cPh2k3h/SMpAVWxW80DWT3vfIim1G/uOoHcDCBe
PLVAjCYGasX51SM1++bey779wo0nMKDX2Fd7xr9hDdKzb1VBbca+y0bu2B9O9SZj
HtydzgfSIvlRkbheXdtGJ1xaMfz7glNXVtbyaO6bVHaf2IPDevqZxvOJe4KpP9rc
/rwZWwczty//dvaA8s0ERgInBLLlHV1kEbpIFJ08XBibcAY99axo3lOeSIZEhauE
CMIMZz2o/BqJqKSR1sBa8zKjnAn2RjKeyunkLnpYJFaj6wilBqv4bsg6TvxhSM3U
wdWE0DlMSXxvzYksI+bxEHOahzSx0c4NorbuX19vHovyPvGnt535jrAqPe0TJNvj
jJFh2776jBkvf/lP7QBsG7HZtbj/bW4OeMy/QZKCPqMtN6xWmx58jtHLy/o2i3s/
pw07fV1BD7IbYb32frZbSbjkVZcQlKF+ocGRMXzgf0W/qGcD8yQM1frIVFxPf6jL
waWd3Dl8Hz2yHRI5tvVUT5+uiUBBiBay66Upm3HF0leVyDjC8VDacvYhfAyaa8t5
lv1fIXj8CxXSMZBFW2kb7m+L3UAWW+qiS2qNMKgPUc2n+ZAkKzA9s2x8iMD0GWdb
izGLD2Fj9ZyVyusAK/MSdfGQVQq456XTLBcYSIT7AnpjumfwOxJQ2YTY2dVNLnHE
SNrZ3Sqy5mBoMiPA+6HDj2wA4xBstUWKI/p++6u1GdSsueJtH4qOZiaUXROQdRSJ
WH5w4WQoCfkStr5VmTfet0kbZBzlyQYDlaLb2JEY1GgCh2hL6BWp1LWIL8oC/KSo
Nk5MjZW3GGmKxKG4kLqAq8LDH85zxcK0Kbp6oRwcsDrfHkj+yaVAZycgxy2GZB4G
XHADY5oK7evGfK4pIGbg7qrZy13kx4fl/GVtYrtBQ1ZkW3OXDPahnvAE8UgryNVH
IXtnlsYeOLxB4lWDAGSKjFNyi+RrnFdMaVghaM0uIn/XPZqfWJ2Q0Q63LJoF8Rvv
QixglgEKmivy+kbZMFM7s1Y6DOEYm87dSpB+g/iCc7SgrXw2H/mR5qKzsZZFhekp
z9m5kqqkubufpXF0KzWZQtLiTYqiId5Nk+QWkl2M3uGnYAOL5h6DVYc4r0M2C8qi
BaQiN9Ltn6IEq9P65Yf64zwsSsAdPO4TKSWEL7OcaFXP7xibF0TqwrX/+rbhCPVv
ydXDMazb4GlsiHIxjAay5nitZ9u+2L9WXMcH2mz4vLGkDCu0/Rwhsq6bh+B13vV3
JZMt1uKOTX07lOw+w15IFEqES4wDEZI4CUb/4HDGzmvjG2KJM8bGeQEDQXFQF2Qq
/m63VwBUA8RwoO7PaeJ0KAqx+pRKRErc22A7Bj8q0pAvZKSwuZHJQHB3Bd74Fpzm
hN80G0mpqNrvaihhT0U9g2nZt4OZBl+5/3N0h2xW5Xhs9F7Go4gOaIeFcvBfjUjY
AX6nEuwZj+2HB4aJGkmzwPIi1RzIHPhtvQQ+jKmvj2QN6evC9mYPlaNY6w4r9Mk5
VoEuknwb9po7BEINy5IRNj5WveUqZRXu36AZirTmrrnfpjhDoTCdyBPEUfLev+Zl
289QgBeCq+8aoGXOlrrVqvgnyhL/nvwPASKXhE76Ae/3ET2KP4pkUn/y9R9NcNQ9
9SizwBPiMNvR2+Gknyf5iRzsf9XzSK/ameLUUPyDPqr309h6K5Es9nnYMxuX6m+k
165pnlIhlyhQrxHVDfY3XBlsWZ4fyyjhsx3J62KqfaFm4J6Zc/ISYhZbmfkEzXxK
11RM7FDD4PsurCl5hmJiyJZOI/F76/Z4ZNsiNBRVi2LreIgKFhrwUhvAV0vE93DH
MMw58oJZcb5rutnBue3LH1wgMcaOUcRhu68vN1Rn8sCaJq2+eIuTRUvhUWBN7KYQ
CmhBmVeONrs6Mo1YP3zV6eABD/82vUOkejfQWuS89hocQhuVuuxAdEm4Tgrg58E+
TOAqMjZrA5HrhDJ+6pSwLBtAjGo9nWyXd496tqTidSf7KW8rtQytHF2SEq0YMtrA
idEDCKLmvKnIxwxnbvNpTrJYrN1zInQHM/omIrlEyJguzJPmvXTIU7thqw8zrOIj
aIK4+Tp7WMAkViu+TGwwCCKFPVykopVrXiYkoiL2Qrx71976eLuVS6XxquK31Ltb
zJios/6xyYp8FiB2P4ehHo4SnvlF3RuXpXvpHU8+EzXX4My5Nkt/Fupbr8FXrqNi
vPaEfuiMmkuCiJmo/ZHQrPzVYB68w9bf0wtBrVhBRigcFLSJZlk8t3NvZzwv/vMf
h0KZeeZ46s9ywHCj0XvBOQaH1Uwlu6XEJy66TdJYwZaexWgPV52anEyinH8x9V8D
axf+S1jiPY20t9wtO5rAUuiSoZUrsToAzw8AextsYLy75UXjsfUM93HliwNCfKUG
0tBK1Jr36oi5NJPD7lJJSzy3aVNekI6/7n32kqIJeyglKW0EwS0X/iJFskZl1j4T
ty5fd6ll4WMTW6dsUSnLVCrwshJuPZjphoplstM7tepTpN+HUDQslMALcF3RAayJ
xDLfq5epaeTWQKqAZexCO0/ARU6e8KpON5eTHWd5oWr07mpiPHsh9XQ23ie9ZBc/
+Q2/48glrXF4iM2IWcUtwG1dhIqRvxhDg4oocmwaBTl3NTYFwwa2jwV2uoc6Uqd6
l9FFc8IiNr3R7a8EF7w9kxsJEgO1ujabX/NYsTH6ytIGZY4KPVxbgkMJPEtlZZPX
Xr+yk9AU2z6eGB3xiYUDkERtqtbVA5ELprHCmPZ6KRgLSSBwtZlg6Lg3IZowLqs3
OkJVcidZqWTT6zYExqsnOs2zFrHPPsuQuqHJywKzb/iYLHXt476pz7cVXJE/PRTk
kdNJEnL+gqVSx7IK5xzSOpKUrqPFu4qDwMvhmbL4W5gutjFs0eZwa5/UWjntCjcL
kAPqOmQrAbT4sUJVYgS89onhaW3Y4nOucnBNHx4h8CLgj5MQCoKjtgIcel+9y32i
fMAcG1wVyB0jhiFU4S7ege43dhpYPHrXz1d2nf0ATEQb92rTewHWp0utDmux8Gag
P8VG/6nPgcfoLQ3RgApEumE6O4gw8ZNg+VnA012uzNzXTpB6sSCgGvKCQtgyAqQk
1kAKQIfr+orVPubfmqi5BbbC+Zd0fjcLuW2ZCtQh9myXHyuMKSkMaFSFjJeRZOR3
dP+QEGeYJdXwGfdhTnrRBNnYwDtqXi1/Z5IMV4FWjseh1/BVothZvFl3RkBOr6zZ
afQ/Ch5Pzmi/P2eSlwf2aTVdMpZqHh9Q9csndl5o2zS/CX/fmTXH3hb2v0ZFpRqM
2IeUpE5y6xx68D/l7ISoJWiB6T+nkUjTRlq9jVEwGkFgS74QC+OD4hBto1Z18h6n
29htI6PiP7hTPvgTlY5S6O3tcu78AnDpTz24HcxaDNkBsdn9/lgttoMdaXsyAd8S
yAPslXLe+RfPQsUfCMghwcyIXhPk3XGZV9RMzUOF594KKYy2gQWXSe7lgf1WJpWh
8SQ5gfTaU8yCnmI1lEFw5GrwxVLjw/TIMrFZA0/4IUBim/k5AFK8TV5RvfPQjJtq
H6kZJNehzknYdtM6mdLUnj8A0ldBGptzqkzCXbzYnD91k8I2SbMNdJa/yZ0JTONt
FEV5/A1R/1aKBJhXohY4P/0uQvYJqBnW3CfD+mzp8BhKCBikfDe5U2CqZ22zVmW8
tzZ8EcUWK7bFB3Ehh1jZympEGzfPDoFXY0BiEspQrwYPXZGyQ/WFPr0zmsnc9/0g
b5bvIr2LYDmkaNDmHD1yRbKYpNRPmWBZQfXHAcJqYxvfy0Y1Ffzy/1sIuVK8eXUo
wMVsfqaV7g8e65W0GF7KHkLlkItEj2gIN7o/cY8NAkeO/KoZpzVSIU6KpopG41X+
I/orln23HQXg7Iplhw/zf2sXEJ59ODIDnsDNbyQYVov/J+qSDdoDaQXbSTQca3dA
rrOx5v6WVfmrUJwSWO1rSpXRg37W3XtqVHVUtSqhamKtCXunlyDdQhI0G6nzLvCs
Tk43nzbQLenwibygaH6L6N9jsnCZzWG0KJ5ExrJPgQQ1LCajO5CZQY0oh1u+vXjM
W0ZBumDAVDfqN7RocKl5V+gLR7nrL7dAm8NL/ym/qCuptNyzl2xfiB0Jk1L1H2BA
zaZ27/inAFRhYjm/XZekSaWwPlWf31cWOx9zabwm52wl2BOGY7n///YvrzWzzZRC
XIOPQ7U3wTvsy9j1/x/VShizBPWxVP9W888teh5c4LH2DnBjQyrWf0VdsFBZeJZk
uk8jRN7VF/VrzAgQaFdLcfxMSxb6o7gaPLtyJLPUPKe7rfZqdK5ZWIzHz6rZZZKl
NiMnLbLBLUC3Zfhm/b6C5GFiACI2idoimZMyK86RLdEnI33yOjenF1XFrgBEU1zF
bgD9lXkohw9T7I3kf6J6ov8kwG8ECeoxeVvtN8zCyOR89abYSpmf2bZA8cc6C9wZ
uZGElGlmRS8byiKxAf1WMhwCxr/+qi57wTILv7yxbokAasZD8u8ZnzCt2slr7NyU
OLynbPe0m1N/zYke48Otxk024Dnw0AFjw3wzKNhA8zXfvUy/sv42LevoKQAaLVZr
p0/yz9yr/d9k3Ok6+z6toSqeBuqWj4s7p8LNmlLrR0s7CLVLTid0lViakJLfmahh
ML5YFcga+cz2mF0WM9rf+QYXdxn2+sMkOsD1f2s/dlR62mz3hJFOT3IJwa/V86x8
3/YPkhgi+gdrPTeE1jbs0ZOjR0D5m3qx8mXp1iMRcbdgqoxTkU76aBTz7yTXAXa1
/74M1K3NPMiy/ffZ44khEwAogQN/i/XyAN38+w5XBAMfvazcwScw5SoDeLazNFR3
Jd9/0YqtSGUKx/2CXHxObEokPB9siDO3oxx/SM5080yP2w4d/l57Ejmo4ijIcIB6
dpoSPPu8GkTXHPtXs8IVqy6jPs2lEazPBF47W47w4oUUK4Uz4Tvatx5UnRFdlkS5
oA6HI1CezHg7Ze/PgQgoECSL7XZjs1A8LCQbjz10UBQKDnD/PMbb3uWVI232bPtw
UZwFlzWB+ZS3YGInzDdtg+SQYIW1qv2K+N6RF0AvV7JFPOIEP0ihkSjNddLw6Gek
sHWKOo9BimMjETprG6lZHs8sqWudNVn6nG4DRq6WutpzoKYRhUQTos8FLcGt2vew
OHjwqFIqM+gGpwNlTKk32bkQ463kwoNXlQ3MiHxAn32LX+GBnUPnePK0XiXN38ek
KDmJZd3grSEnLm/b7yFhFrvxA/bw9713TPDD5aPeFiBNoH6JNuQ5mghUGkjbJDXI
bF4JaNThiX4bt19uZzYyceWHQrm7sutFHFjqmjEeCUU2Jdfr767yg55AAqEjeolW
qs69WADuavwMwse8eZdwccatd2zRLCbOdS+GJfXGUOXK0vb3UUV5RrZ200LOPO6K
r+irRg5bEkOb2nGbPhEGwS4qhkvVEqw8UcWXTd7oZjcUM1BHP+pfGps8u5uEwUq2
QjOXQX9SJNB2QDm/K9vsA51Vx23UyZV0t64OFDaKk8vI21pgwWTkI2UYHqGuxAF5
qbI8B7cA1jIRJ943cJBIdQJ+586auh8zZCGT/G8b1VMjJYwmqZiC8cGSLdtSxFMH
YCWgXxlxrTndyixxcWCXToeRP44V+FO4BrHNGBPvbLHDrzBjFpNM4w2b0QMVcybT
fF92mATPaAujGshl/b+UiUp09sS1eO29GnLDpGXMcZoE0SiEIU2YR7MoapZSU2Xu
QMqCFiLKe+2NVYV3OQUbyayYhbEMnFjN5NOa3j7lgjuMxI0PpxdTyj9cQcyStc2t
G87+stl/OXmTcgQ5orWEtxcSetFRgwoOK5FZd06a7T990WVmvm3f5qYNNahT21TO
RX2IhV5Impv456aHB89dIGbWOb7dOJGcsPfjT9mVARvRets6cVLPPM+RShovBHDo
ZjI3NK5/e29+MxtJ0HE36r+lVZTbx0D3fouahDJW2fhvzmdjYtXBmz2biSkeTN9v
w/b+PiWtuZ1dZRAs5R/Gx3YFGbdO+4L5S7rp5dZKFg/VlzLQ/U2Pr9Ou3VJHXOgK
5XqYXA+vP+slc6Mm99YfnSTrr6JZBnUqcl1QXGHQBmSgyepea1t2yTMJJlsHvp6q
jss3IxCzkAOKZRcLGjwg9SnNRZjh6MY4CnNgfEELlUUdbHIEiLVLdeN3hmOF/3LZ
A7y3NgT9Of6g3+P2mpjfjOQBCDRVUTKXToRkx7N6pBSJia6Htfb3GbIhumL0r3Gy
GnlNPBQ1kWGoTFhOtRlBIlbiSJL6xQeIjhxZfTPW/1lcXXaTS1osxI3WpC2J3PjW
fD4mZWfENSEWGIy/VDRt0sNobLI2NnkxbZvTE3wS9JtOrWc/yalmhFxTQTkVVDSM
DHb2Ky/jmfVi8mL43NnxhDoR7yca9dKHrgTBQqSpEjfeHwtuvAa/UccVa3o+x1bs
OdeSi36P4+4GOFNX5YXTWB54cMf1u2pCbYEYiYZ+prm/YSUkmibMerI6qQbq1LNf
GCGPrPMRI6AxNrQI8bq43mTp9s7ueNeaV2PdZJ3ZF9Olfcd1VVgeuKJVjX90RKhe
MdabINTIlJyZFud7Cg6Hf61DXP+olU+9hVCs+HgLepRJErOdAcJAWlZ+mY1mlNfQ
heSpiHPkbLCRieJkC3kNVaA/lMI+f57X5EuzCj8cS9Fq4kGLfcGbgQpE2G02C9T7
wBLAp8ta2VBwtltbAwd1Qja6J4TQcI2Ov3cDrNH+8JWFAl0I7Ur6B+uSqSiafjBO
CDuQ3yfY3shfY36ocfjPi/Tx0C7t14Ni1MqvvaS+zjOWidT5u5jlKWMXJn/+axUZ
n/bRw8D6Xv5WFYS3ChyL3/HULtfu3IyNoZgEXhERPZLzUmHMd9BwKuXl4/hfqAhD
ZcfOhGH02Cz9za4cMV9zfjiTKAs58rPqUfhk2SunGmPFqL+2vYf4mnolc1nZuG+k
wqmR5taaErrEFfzq3FyiAYjEzbCOeGnMsaSXo2UriydhcR5YDZbKZNSg5ONoHNPk
BDs290yjtvSw01ZlKZsV80XiDd21//pmFVeCIzGuWHqs7R18+fetJEziZoA0Fvdn
TZiADMoYtsX2wclY0PAf5t+vuJKpSOoJsIkFC7NrZiWcCZWPpYVfFL4YuMn1HLVf
TPw0hBDKUAdiloiQBq+8vVqgiyWbiNvfGXQPKKF+ZdMIwEs4UytVUrvAqHmAH91H
UNvjz0A2sd7K5sETRs9zJz9V+BIyvaaAzmjQ+2r4/wBjhrxsM3J4a9OmHITsyElN
W0Aj3W8ARSyqZ0Ft9sBkjWVe8GMqto9PenCCZjHDSeU6Ci7tafa5GgAmaYeU3LXu
ZqHpYLiZ1v4xRLIrW1QzVReNlzzRaxa62MqfhpuRocTQpMx7B+AL1l6PyO3OOx1T
RyaWVmdk5tFuFLYszzu+OHCm/08MIKqEjuwOPZo0kEIdjjY+vtRIemhPxZ0yeLa1
aHJYUqwAuZEEGuMjIJ4UoSLNQunCfAwI8R6qvXCH49cr8LvXSjMkR8m443M1sVTy
YgDrjkg9cVpWshTUkMXsrqlq6Q/9BgQ+rIp428bphoytSfaC3PlCs66jwybzXf3v
ZSAdC0sDgmRJCCioz67FS72UnMy3nlUCZaVIfB86wgx6Oo+KuVJ/QWSENwWym9Ke
ToxodnC6YQ32kSIMFH16Oci9t7a924yDueEDRpiiKMo0HpBB3ZO+tiTLOz7zMJ6r
hwzfsrKOhItr95iSG6axk7+xhbywNNQH45R36pRIwLGlByFFis8s468/XpwxbDNU
60B33kpl84fDnaRnKw5FRLIy9vucZJuzv+Ci13c6d1pALcc/AxSYT5Q0g+7tMBSh
NBWzcDLY0veIyojM0KkkVwE2+0p3heQatCuWQov+aRAyp42pdLSv5C38IuFVKN6i
7yuBXYOXgn+M1y3T5mOMQFbXm5xTI9UmOnrS5tSf4L051dWTI2dG5Tu9m0HvvAVc
31pDQ+3Qlq5WJnF9xpEJpoYUUFIgt1GpuLsNrw8WADRXsdYMktXrba02EQ16bYSP
cXgWUIzh4jq6hjniK+qmJckXR2ABrwWdEWwHmt3T1d8TitzD1dY8fkZRbC6MCiZL
pMkcC4VZBPUzQV3a0Obt5UxFii7/02NEU19bLX3r+MRloloXLKZHmOW1MzCWzE1e
1BNrOakH0089vyLJQTeyO+iLvZNyz41Lz/JoKD/A5+BMmlOs6C2zfXljtvNsy3Hu
SisivxW22j7nJxQYdN48degQX83CfNtgrFraLlw5gVdjcYQESZxyR2NRAhBiOzZE
eT0wEnX53abeuiks6P1XHsHxD6EgKD6JtOr0SewiOcWlPs5YoeNdxOB+rrp+eWTt
jpVLb3w0NfC6rlSxxCGicpbHB59wD5b7reI6zLg91Cmym1O9FI7uprd1C09X92/X
8YCVHiyanbIcpNdtbHvwRivT5q23jGGJchLUuXDZp5NVmOVarOKJoExyyd7a2dTu
RkmoNOyD/UY0DndgfUuS2bAU9gAAnN4R+C6j6VhZmtfXjq5Z84CeP5rem9jK7wzq
zgkOR+2w8TvWZqnM2srfnPaqpjMfEybQ9IL7VzhS56hFueB5vpZ3tTv3uI5Rp33H
CIDu1w46L1qS59HHXJIrSaOgajCYON8JhlpmPbsUiiQ1inWA5MWsl/jVc3nj4nNd
ppVk8LkG/6/ka1IcgngoT84s2pA+q9GOh31jBUBNERr0juLQEor6x9ri0jBfRVjs
Q9ufQe+HT4DMka/8QMiTK6Nlnzt5vm5akE1xij07xf6SW8NySCJiMKcXope9Pawy
rEZ3gdohBUarxOYLi8jDhlk7oLejiJQlrPBRhY9DMrQ9SQddATlbhW9p9QJsjX1d
dJ+p8v19sj2VEtNH3U/tiVQU0OK2UBlmPe6Y9VsH3e9k8qszreWExzkf06GMam/S
eb6VJIVK4gVw1EaWdROkf22vVHOZO1dhfA/xnsN37Vamkb5nkqg7/sOsYewXfVXA
m3+TgzP8Rih+9f1VMeqUxOXX/aU0eZZbm1hrhDoOSvng18KWb5OWJ85kVg0wC0UP
+Bvafv8FGLQ9z1CjfrArksdg2soyGQUdC+zaCWFWv8YUg9zaEalECN2HTKhBsNMV
97jWsZLdBwzINqnmdqyRWN57PdCXeUm2E50ZfaNYGaprEs9ISe3OdWo2IOr8yf0m
xVo5xMVJVV9m73RwmXOE0agEyLjR3ZIUd6T6yvw1qNXgkMBN/iOdGWEvhNnCl651
Sv20asTs0E2N1aYeektCN8up36l0K9vIcv/fVDX6/sR8uaIZrEzswJBcusjKMK5k
NKmVLp7NJaMSHVkJDdWcew4gflMW1o7rZTvc/F1AVp6AcNFRcwuBIjxWjTf+6LXU
4YGZhiIPFNpUyWb+n4btkEwWLX8TX9SfdhlwSdKv5BRY7rEL1u7yktzuPDBInoTU
9sy0AZHojYgoPa1SKde8GcVRwQ6TiYN0302pV2oLUz4H+T62n7g6VBW+uCIIk8pJ
j+AWtWexm44fKCcj5A9cIbPlnMo8AgGnxggO9UfcYYzH3pUlFMjbj4wK9AASq2CM
oWFTWHsfhrB4Ub5L5Y9CX808nNKZRQHt6mGwTIM7dZ9hJ3NWeazFxy2t4kncqJHS
2mjOdYKhwYLDRq1M81RvRYtfpHxaeEmrAkpkjlrz2vuObXYbP0lmRuaTHyk/Vri9
oai5a4yRZmRWUVGcfKRtJXPwMHwbG9rU+DR6DvkbXTPb+VEogMMC4BQZLg0rLBkU
LfyQuZF6QrcIjsud6Q3yZAOT2SG0XsoEJZCKHSOTE2omHCbY/OLMXe6GQ+x1EFXn
b0lrYvoXkbeDAcoN6zQjtSkpNcauUj02+sp+3meVf88TIMXzS51y3gWnqU2Fv03B
VFmPXIvTtd5a7CbAx+2+ZIoAUitWZsd9Z+nok8nz7w8wO2dRROKDjuhvSeH61s1V
I3XV6YgN/KS4lhmu63qX3lwoXyFu5jXsNqgg/LpyXhQ+ks7+tJDymtVMIAyEXfyB
x4zOCqVlQvDr177T+dMNkmHkYJMIYu5ohdB0vQ6Etf3/nFLC13xbjr68h5fBz3be
omXshqCzyZGLKr1Ba0WMZAq2ExX7UBfIvl1t4TE5D5eFHQuOLqFvfnYA+IfImOy6
UaBnWkx1CaqVBk1eiUJ/ngOlACya+iJDiqIg0namzvS7/nPqHmvx2A3kUVVKbX1f
fjrtwNJuSXp+ahMhH8Kg5q25wp2Myxn55NIro/SP3gOXwF8Ec3MIrGII7fbYjbeI
dfQQCaqlQOEzqQrINy2W1tYsQZiko6Vuiawbgon89bsxuWgRNp2T+LhWRIq3hmhz
DvKKh4gWiRgJuW+PiuvAMxi76rG0pl05+1MVlsYm01kxXiIr4wvk07BEyiaDM7B8
nAEvwCtwPOagyYWvmkOdfEW5mu/c3YF26ladRuDzKbwB/wjbTm0DLBkiJD1+FQbP
UB/vKg6gkCpifMXQCARBDJSqhMGAiZUW3tsOQAaRRttJKqRNptGx0UipT0QrjNHW
as09xqQL7AHkf53m9SJCsieu/3zA2eqEx8F9H4UPIjmrHnjRsQhu9B8KKtvENWN3
NuM3p8wDOU+5TQs140OE7Kj71BbCkXD7Zyi1JBTIsnX/Kf/fFvjSwtC7/qbHbhMi
cSsHIlvZwOp/XzkEpWMlv/eU2AMgXr5/BADI2WUhD6e6NiDyurrS4Zf0Bs9qqMqY
w2x35iBvp2CE4lvZcylNLSK24pBfWk09LOS9IGlZ3dPABs6SMdhOG1IeH73pUqJG
uEu+EO7CHLBUKiWbIK/iVN4Ffkn0GF/NRsnmRrzZkPZLD0IXHm6PGVrNnjTR9/ma
2IulfJ9KHc89NBLyWy+qha1KpgjuQc7kx6JASuOl15PnYVj6vaNjWjoyDqMT4YOj
FDtpT+yLMRkjfB5SK2Su3M35E6/0mMFlnjH9lKwh7jsg0U9fhBnFhnDWX0qB943d
NTZ+CTGnqo3mMJSEhXFoO5Fm5vfM+OdPt7rzP5uCbXFg0uhtdCLIbCljoRhGODm5
ogM3zD0xsyPJqSJZf8aDgktEFNv4jFirnoG6ij3dRQdWAZKsRmrsuCcjlLGxt23E
oaBgFWFVJTj3CDhrg3tl97JcLj+W1ldfjS/beBj2JuaXyicA7Cgz2otHIAT90TDZ
W8xqnMfvA3aaC9iZTjasLLE1JtwwQP5mMEiycpnDPsFIHZT8IOn4vlwf+qj8IQLh
tmNuSRYGJ7X98ZlK+kdwA5shtTq8+qfu3g4niDxL0ylCDfQqpa25zu3yRuWkKV8P
bG/I0E9pTpyyU9Wl7MBIcFn0Gv+M5Vff33iI5lK7JDDYBfk5nQJFnT9wumS8tuk+
hjGoOTWFKKh/fASrIoSNzEUqRntjYe1YHtqIg1JJSgxIm5OmEkv7IsZoOKQjDPYG
Z2UFelZTXGwQy6qp37/tkUDYmrUO2k+414xW1cnJQZyj3QKu4z9Q6LrVxtjwWg6m
ck7+l5AqzYiNM7k6cKZRdqW3xdiAs9fkod2T+BAa2mWZ/7gtiP5ClrfrPenBC1Da
ZZCjQQUzX8wX9p8xwbztmlhb1ZFgZ2aH3n+kNfsAhsucRW+Dr57NPg5kVGEYTuii
ChFTv7IJI9nRRX5O06lJBuxRvq9V9G4556yoBPXGCeVUEefqcZrXwEau9cus0NjL
Hiaj/JxY/NH8TbbAUn+wvZB3p+hgTtsdVE4JEpbNI/ougnKJo5aexjw3/B1Vz8/v
HrYjBm0Vfh8uZ4QU1Txdhh6m1hSn7oh/b+hy/FaMDGBZ+6TtSrqunsmWPYaPho8n
dN1xrZxtSJGqKt7/I+wHhI/y5gzN9kRT7jgGUA0H7yvFb2GzvncB+x2RG+cL3Njn
r2I1WLrOZe/Ku/1Yup9Y2L2JF1Dz7JwA8zyJtM+stz1oGbUAmmyzyxK73kn7wgZa
qbljS/27XAE+CfX5jyX9luF6v6nd7utP/GxcvRjnfFTL+jyQLKv0MZcUJSbblHwJ
zvGpWRyVo0SHnKwANs6cpQKjSywXOQnR0MxKt9pgZurGnOICdL+YA4yzScbqMQ92
8f86L90sap1EmL/lbKatPhi+eSnfYpEuiMQDGIzb71M4WZhRVUl+4g1OlEC6cepE
occ8ibaEUuH1WjSK1TOoDwRDU2RxtNrZyQHddTtsRA0XcJGji7VoirbTFJxmDzu2
rgHUulddPfOYOPVu8m+gtBTaCW7IDm8dyGflKY1ODDuGzgrDrRDrL7VZJa9UVXIa
4GwOB8tJY7QxhBASey8vpIAjZQfVXMkv4iQ9EI6trAwra5CJqx+8gbQHMyIKbGCf
nl0xQEMYhkEWP5XMLP2TYMfTkvzb5BIcoHI9lps7yUrylsO+wCIwu7zZNJUhvFYr
1MVwCqtEwX+LIYe9NWB/qz/mp8YwTk1tRiofPl0RHFHGzHOwwcqoo/TZt7HtPT/Q
MtUz22/fC4Dxaghy82V3Ty0aYM3TvztuL5P6z5r13zGzc0cgClZtCYTPGiJeH8qB
LqsQ3/mDgIhQmRL5mWlhoOcIsJS1mv8MH/YIwGeFFSM6H9w5+MwFWZx5+z+Ju/Fn
pNiXUea45jm1df2OwHa6ujJdVN9or1k4BnL5H9r0ffwvK8MrRZEH9M7sfyoq3yCo
NeIY260xKGPmHX54YBLKCn3UjGGGcQRAI04uqWA/PTSEwHTW6DOp1MWLR/Z90Zuw
Ou3LM0y0/NVy36LirUzy5SMnr79ABlc6h4cMmGLsOebeG+mZP/5SNpC9cDVYAk4m
1qYPFKwvcobP7kMnmFoJoZeKZjpkXCR+NZGkZt1QGeyrUE7ACvTYbwU/JWxLgFsn
yDe1MGoQ+sG7t9OOkeZr+kYrH2ZPShs2tnQS2dzik8f0K33E2sF8Ek4wyAgVg7QJ
jUdBcn5BCtVdwe7hKGPcSNg/yfFsxey044oxlmyDIg7oCftcBlqNQ/BZht48kuw/
CPSFVt02ev8cOeAzzfFuh85f9xM49Mb5m/NTGdm9h6ZZuE9ehjEL7uQOEMfKhlog
sBG+5ccW/IfWrQ0B1p+JnYJVBCFQoh9184psPwagoCJdB/HSBSoNP18BmaE/T5Bc
T27cGRjhSjRJVf6fTGjNMARbZSBzzwwIa23hRR8VnFGpLbIz6xUNciljcsWUQmVt
1Kh8IPXzBZ1ODV/eKgsjuzJMMes6sKxkFsyoQolWxD4rKf4UeA4srFBsGM5QA7uX
ysMBvtXMCn49fClqdjSvXgDK7EfyhDNVyPrFTeN6bk1qBU+uFRxvAAuoMA8nESTA
U12JnY/hAaEBg4bAIzOoXIRDyr8B5kTLmt4QC/lxcCZigZaAaCfJSmdFJKnByT4u
qcQ8DYV1zchumEbIBqYmEXIQMYJaIle1QIWWrM39tLOVIZXsBs1YFkiKznVA1M5E
b8bbVMyNTsoKd9JwkxJy61xe4NFWG7Hc1pBZR8jmWsvuopcd5zdH6RZ/vl4oteu8
8fHvr5NWT+kA9g5BW+ZHBXL59B5T+USSvcN+VL60UJFV8B4x89zBlcRuCHCN/n42
RVYH1vteuo44dDnP/OV7saiTHOyx2Fk1dHvGyd9VsOf0MH1l/mTmRCCmtnLWT5jk
d4xM5A30zaD8xCdKDgmNKraLyx7eexjy0ET7y2AJrs04+dyV2PuXCv/GvMqCqRy3
/Mgd2+iugVWQatwXIO3dkB/TUzna6Hx/fIbYL9JWsowjEwDFNN2Qn1KkcoybW/S4
tC/R65M5qwgz410duzyaHqFaSRhOgguyU1K0nUTlFn5r6gk2weseM5s/hWJbOYUx
CqcCHlWWdsD70xJHkglE/J/r+4vnA36pyy8QMn8VO6hpaGUU09hiBHtNXTKtAiRA
s2eQ2xbCB3gv/NSio3hF0WrqyappqVOD1UfAVfRKYvMAvyHk0quwNG9Nx8yK1toi
TRdJae5MsosRBNw9i5bL8zCZ7xCXLvAoNJQKsWFgTiKc6lRruCMzR7/Q3x0Wut70
vFGrHmmFopQdfYoj4kYKPyv23RKNNuKDqlgJjy/oh88nkWsBAVKhm70ir86N4daA
YYDk9PPmvq7Up4fuo/2KGc/oBahMyIWZ5vdl8UcyUzHBLubMvKyjTWIjCtWUs1xa
rEqrAABP44u+nyN9Nfs4jhSamXb6lTGS2G/PBw6bZCSxhDKMEKw/n45hHjYTO3gT
c4jKGIjThbYygtTmw+ZNP2DSPEuHHgZ0pWhS2E5nI1rU5NStccZbNyRqLkjgeIdx
Op8ZqhrFHsOibgB5krp8d8WErF2p9rNDIEmX1wqV+Eeh4bXop6hKVK6RPFiAVKKW
paDADzhf2CxruTGNHKsvNmWGYp3Xew/E4yr6RtRL2OrKyNwMgaIRecbPMXFAPL1L
57141+wimgkKCyNMeJHTUpHGyLavBOxqYG0pvHAt8ZPuiPMQAPq6GAU2DJRUXf0Q
ARFgfkzIXQcu55CA+uW8AQyyjFj9Fu5zhg5HM0ZFUbzSlUug8yjllXXBR4wT/Z0M
OHqxP9CTBKAEh9nnj4Se/YqaW6cnyrG8iEMUkFmkLBKnTdtGw1UxtN6B4sb0LpWy
JaKMUz/lRn/lHZKrL8ajRazJe7Fwsd3Q81hcv+V9c/RP81vnQR9BHx3LmEODuXlb
qywr+wJa4wqanC+ln84m6zOLG7/1SVBgmYuF5sFyEJgD0KtU5uIFcyI2QDBMzp0u
CSvX5bKwmDr8J8wopMfm/4xqKv5oTIs3HquXHllo8EFLktgDO7e6bantKP2w5Y8G
zmgI99IVIy1OdZJ5cYG3qkDvxm5RiMT3lyMoUWNM/+R4qqAK8kx2kTusnDqloXzg
/DoQ2AitDDUdVrWQCfiJlyhUwuMU2cln4HkuRPKQ2pFYsyTAnoZXQTJqfHkqAi6t
WM/YVm25hVilIhwTzFyeeYsQr14/L8NhNxD9CR6ACwkCTsV7FbuO6Hy8HoXV2w9v
j8AP880FtVcpUhMpIn9iAZ3Y8lsS3q9Nrs6McZbu/VDQ1jA1+a4Za+Q1qsFwn+tO
taBQVzuTuXZdOHogfqXVmGs+7LTldhrCpiiks8F4jV3WsbvsMU19SqtG/HwqOinY
LTtRjAluI7Ama29eqDwC8WqyGWZ9IYGiQOgefI4GRlLHaVoiv9K1JbY1Ugl8/Gcu
FSHY0gEK4aooUyKCLag4lDdRiOWmTg+/CygaYEg/+6RQpCJJ6mJ70wOtiGuzhlPX
9jeQ2T03hMFPRAncIlyJ6cyPmRPBIYw7owVIRu8cHtIH+SElIssYnmmg2Us1fRPa
E/WXe1c02zKfLVIQrFRPPs96i/SAb08h/ZChGqOAIYAMKk33/Soy6TRb2DLMH498
Ia6h7GIeF/hlSrT4CtkntMljzxdTLvlT0ggXMx5laD4z6Ob08aps0V6oVSx/ZyS4
Vf6r6VHsTtTAKPu7jQsTBSSGMEUb8sJ5YaCIrDgM/8OZzTM5VTXkQEuT2LRHYm0C
31Fsj+7+WWykrHwfLoN/CO3BdF70OIeXykhYEJ6pZv2Vr7SWNjk1FcahFYomprvL
hujrhcn4emGVy+pXsRYPlkSVzlIZ1e894k8c3dNqbOYPsg4LoVsV5tKWfjpzw+/T
cJT8cIPBsfZ4ZGtCVw1/wfJaueqE2U5gyfFzpLUyMamvJ427GGwwZZkFQwUvfZBt
/MGHrsJz0b4N13DPioInXsZNS0JltKxpQiZSKlAleUx4VVM/OealrOnsN+fIyPqX
L5Y5W1vifzqwOtZB1SahOpSnX+8jxUzSH2gZC8A3qnkMXSHTmYTL5ghvCNAqsr1H
VSQGIbEGfvV6XbfQ5XVTXe+wayrmkcXcAqyow2PUfWR2oXcVIP+NTsWvKBMYW+g9
qXYPYiIhfO0ANCHGQE8ygj5uMDfciz2OeEHNW/qwHf2UwyKFbBPqEjT2w9ysEv6y
aGdMt6yThfatP6BY17TNZms2PpyIMZlaH1qvFX4DJ+y2nJudPeAKcr0BP6eyCGpx
FZO0CxYfhKhTXUKXoDGNo2dWa5NTYSzdJLClIhSaD76caOYsXcISssBhxXsmguP9
WdXiY65jYdWoqGgGR/0tUffITEKyjXaFggihnvQnP4OfELtbYTFlOyX4LJ7uh0/U
ehM/M9pFs0cJGwcody0B8V4DOJE5g8wJmzhHQWUUrZm+EAYwxmb7jvRPr6LoxhmT
mtfca3phnsyu/F6NjY9cmvy9vb3q6lH53e04UDWluQ31JoyGyu0nMzwre3I69DO9
GcJt2JhPCS13E8q13U9+Ux1Fv6GMvJ6jzJSVgxbPpo+Iz/cDpLVhjarBxkpAzxTh
cDoJ318vTDN1zss+d9bai9kBOe+F30y1VD+G9wMSPlIol9hym7VYvddFNsU71fx/
vPAtzRFJIT449GJPsKH4Ola3qbqWSqpSeRcrQ8lQOUuL/kEnJ/eFgV0xUI6qkP7Y
lZR4jeAsB6MKGHC61gYLY+P78ciUMRhZR0/vr8kUJ8JOBFtIn0O/pMQLk7kNQQHi
ago9SIW/DQBBfr3nauQ+bSfro4q3kz9Z4bVaFd7/9G1LVX0GwUEGIDraMVqjCfPG
RPrJ7gjdHqEqUjz0fcefOw55H48kMKxx5d4ngCgzPHTqpIpWBNI+XC5IeylkqOX3
8MvakyS47IATQY8Il5kK8Ihj4uw6muwCfoqQWedjUQ/ip81gokxT4jh6a3maX4rn
CIsfLtirX+84vIMUxopzo4WSC8LF909O8BNHrPz/u4bCoRDQd5i/0CKNiPJZO1VA
foz56L9TQ/1i7MV6Xr0ZwLtGdJtAyt/RbSHhDBmBmfV+rEt+6qAW5tT1sERQokFP
AdiIA+jp2Bdk5MI+TTHfyxp3WUPDz9mYWO5ESWYbVl2G7iHJy3+oR/J4PEM5Thn2
+a7PhC3TfjWz17X+mAeQoE5qkh4BRPIJoeDeqYM+yZlwRZZTyMvqX4vqDc1+L2BF
6eVHr6n4VH7uDRnS+HJ4hON/PqntSlSPWPOCB68XKrCb+0sd2jIs2hj3YiqywrF4
FOtHHBvmLsGxpawL+JnowlTSXKFQVSQcc4N4/eOY3RqBQO9fYCTAkfWQlGHjYbxr
jod6vxiQ+/QIgaNZshZwiz/w5f5xIL745q0tqO8TegnQ4R96Zb6i6rwPP6L9wFtW
0n+wJOTbsyqaqjfnAIRSyhOblpTfMHBOIQfQ6hm3t4Y5cIQWnFNyQDPJnAj6qfWH
7J49TjLMRiA+adihxsWP6Ex1d0KY+mMLnHU22OnlrdscTUm5JZBIfSgKSes04euU
qe1qyUruzMBvtmdwc+alJUMmkHXJA060qhhZ5Q8oUbkYO/HXGocQY1j4k7sPXZGt
kyNpIcNDMxXDx5xxgWxRnzlCJ+exu0zHK1PzI+hZAnQZ93yv7LT/jC1BXF6GT9uJ
t3oCidl40mlhTueQqes46h3A6zTcjoi4PjL+TPwe4tcGSMr4T19GDMrAe9G+Xj7r
xUjdjVbx6Xd7+U058G68e0UzgrCraGVAPmn9c3mpzJUx1qtTfzx8+mZnxWo7sM8B
StJEa40BvQgL4kHwo86BslQM8PcAcw/pyDYKyilOf3crFEVrLk8Y0pGcvKm9Gj8F
T+Ozo/a/qrX7DylBbF2JZ4tFrLtrtI2HzDbpYmv5FzdqNWHXti19d7JJKE2FZBga
fOhNKrwTel0yVOXzhYVngHVxPvHPdhkQpdEumMExs1LLLQ3n/Y83++JV31Iv9YGa
+7rL8Mvt/jmDf+yvaj2DLsMdpQh6OpeBoaYtwtSdZZXx6xINp0mWO2kPv5OQfmNm
fEIDfYXn0ZzWrI19xKiyIjfXLAzT507me0yoW4962C4D6J8kNCn3a5/oJSA7Hc/V
xvJbDdEgfA3XQNSdtB5/pN9v7C3dVLBxmvZzU4wWEftiOMLR86KkMfTzeRBs8UtL
tIKeMJximmuzvZI4PuJkykm0yoU6ewsNechDR3pBRsEgDdIp4JdHJ6lWyk/4KACI
U8mKXoj5fs2w5vRivh1sD7ClqavfyoysbYgKtoGu8wv758CUGTPahj3mvrXz0YT/
wWjQs9ykl3YlrkpMdY7ZdFyjTg9BdLuGY4ZSRHd9+5rW2MHQWNCtMQzXKZozLdWv
hlsJRz70vwHs7Ur9w8h7REyBgVgETnLHvk7iy1Od/20JnJwGrEQBGFcvFO1hDudI
qc27Ks1aDjUdrbDiSyoc87scFTCoXCA0KHD0mmKeYPpjsnNHQcVSYD9w5TEFx9lE
01H/wunBjbZIS6Axh7MhVO/n9Z8NDGWjP9fG4V0S7YfECHIZ3oHB19tCS09iLm1r
MCYxkllnocyOTNB1LV2sBUf86QlkBdzOPn4NJIrRTSZJn8Vpo2q6tBjsj3mJh5hY
lZkWU3jQYD7mOIzv5f54YcZxN/EhfW7MjgwaCPMLstkA+tlXuiNALT0yg5lkl4j/
3aF8MV2jPa91MABH9FDABJzSefTr332qzQJrktJZMCwfrOIVS81+j83D6Wi67lMB
GnX2+ov+dFj160skDfcE1pkwrLvN18VS4pCWq4fdMXGqNz8rxOcDS8Db6Sp7myud
mDWI4rCCy3xZDH6wQt5vun6npMMI1vHHVHE8guMD+aUjeKKiyc7rds5idqggu3u3
rVXvAmkC9TSY6to10ZhRMmTsTXZgu3x0tWjdnVZNqXUCyO2DoDReAOoBvz+G2A49
oYgNSSSn6fs/QokIr9vzn865eLs7wmEeXilSAhSa6UtkqtQHKAKaAXqhVu0MY6sO
UgCpRud1Lpjk+NGIQFqXeKKVW3VHTtVEiDlfHRzMgft9ZoUPxFKfVVbbxgUf+F/X
0bmp8B36k2Vq/+P9+cxUtmR40cv9+oi7ysjzCM3UFcrsHqPYDEjiNJEv5uKtoMVq
KTfxJwZCOMypDo5JY+LrmKfeGJyNqG6+RqerQiH4TeM5IcrY0iMKPZXz3zHZKRVX
ri9FQFIYWj8PWLdBj+bRo12lZ3kqsnOOT0hmNw4H1xQgFQ29R6TCxFtBwKRMM9dA
x2q2JmCjj3JgT3pxdN4OO3RD7So8NA5JZp3UrbtnTdLivAPyYi6ADY39w9CAxXYd
79cRj14jC3Qs+0GqDBLeVpJvSDzMZ5b8isQGq5mb8RSzRouNi+SSTDgueN3QVgwU
mqQKXBgW9VsNsNnP+1rELaMJBWptB7E1zQLI80lZMW0JUV2Pxu8M7AqQ5wSslPKl
HAXQkzi6JT+nE77onjcSdehjA5Cessm0y8aMBtBmRikReR4FGa8PEW7jaApfPZiI
SRHcW5TnDnE9bG+/MbKbcxHaipIKqWXNM0Pc5OMog+X7z/qnZ2c5EqEGeQCh1hwz
0VVJnQb5mznjyKdc0FuwRnxXBQlanYhNuDxEfN6cx2f73qrE9h63FYZSuVj/I/iM
siJPzS7ToXF+9wKphbNCiT2lYsQx/6JKDpdQyPWMrfCsVnz/fJmpVZ2e9kO1ixx/
lB43aYsmnzC/4F3zAYWfweTD8H4gRYXACUgozVx3jtB9HFwPFHN3C71y1avJie0N
HiFHU2IC9/A7AfZUNKBEOZDlrwUlrh/JKCqdg492WXU6PLThiXBlUwH6VF1OQsrE
qa4RXxHOUuoCmtKP2sNVJGVO2YbQNe7CHDyR442UpIJUVrILwm+Cu6TcKRTsCZks
+apo3sgqwiokQ4veX9Qiwk6IxrdXrt7svTqHhhqOO92wBDu7G+VRH/+wTxTNPT7i
iojXxOkK5imaXDYbIOavmPfEDU/0flYayK6WOcZcVV6ANIIUde9hkX1YWO7p8uhQ
IvZeB7IuyO7YyxFjijQEoV+79jjYGpMvQ9UwmicL4nPFvGmYzVJxAfpcO1XZ+OA2
H0ZUT1o4bmW/67hcoAAU05iRVlQm+DvyVHUR6ks1FomSAoloUFx8uozrsdJIpYJS
ZzAgu9VZi45TLhpvT6knj/WHRkxnoaaxYfrHJUfFJeuNLnmOn48E9UNjY29UQZjr
QOX3edWb9S0t5FbkzwDRaIWe3x7aVcRZ99RbdVsG9FWwpjcCtm4SYcFH2PoXLlpR
Yw3Y0JhtPfPlPP/sjNPALDT3/y+owN5DvPTj43/N/9zJ4TMJ+nmjTjR4CfA+YY6k
Mzw54mxSfGZjSvkhYKwL3IOOVDI1wic+yhOvsBNK6qdZTPtuGQPYCn1V+9/95wEH
GCwjdNqA44ZDxF7a+bLf5Ms3fmiYbdkhr8ukqEAaGOvcD+FkVmrcLtUze9GfD3qE
A81CQvWVJGleLZmgS/8+qAaIaKq6ZOv3aAqbSdSw5m522PRmKIYXy/ggBppz5cgi
raEbX2wttMsKnne0LWexvXGdZTk+0GyenAO951Izn8dTDynCOj9AZzKZ1bgQJHK7
A+nUToKwTKOqkBkOeXhOx7P84w+A0ivCQ+YqE2RjWDsezkmJ4iExycsKbToNRp2w
oh8EiCIagI0O1Af2JmykD1EV7j6+Fxfs9OFeE0juU2qc+fl6JM0wz+dg6fqEIJ/C
bWDoBx+JOH01lX1u3Q7QJcVuJk7E7aSVmBdQZ5GbIKGo4ry43H84YLFGExoZa9ju
uot10OHa3eqBeOCK+BtrqunDn6db6aJuWv7A0cBlJxdiFBcOfuutb8EwAZ0Fn8Nw
R/GkDEPiT4OQvD8NM5C0MsWiefD4gnBYusghUFQdYzZnyl6TWYpAoOAR0rgNHThX
Ppk8WPY3UqP4ZQyEh/ordtdnW7fYbv6pNorr7AJSkkWmZ8BJf7WrphYl3HswWefk
WXHvc/lmzUuNOKmTxAZUQBx7sg+tt6EVWBUzKj46UGG2SbdloBYjKiQccpmlXzPb
UAvgGrOAvG4Bm5xDp/gxXIkDCBh3YQZ8aMtWsL1dXqFO7IlC9/f9oX8hXvbRQgEg
c5OvHuStkEb/lu3Fy/foviKR1vol+WQSZrFlolIaevBZ0pMeqMYSX9BWSFAmhTAX
36jlNmoryPrb1Tu32TfN/vz1aVycSnlokgv4b2pYAvn1tlMaNiO3LN6uFKDDUIeC
jIJxwkm0cvxjCdoOxwHr8CPJX+mcFpXZsI5sDIimn2zrTALPq/jykcHYcXju1OJb
lhUJrm787cP9ZuodlUxnNmSNui++Sb8ZUmg2t6qJn7M9PgybiXXLcYVlLft+C+sr
OBdaR5ooCL3ccX/iJjirB6zSV8tWEXH+IzO6tIhrMOx4YxCxu5fAN+xRHMkVWS9R
1BDEWtOsMXP/ZUUBh3G9B7KKA2JDpRLE6mvooqWcBtaF1eLEcSIMznzNRODGRrbq
9csABFanCqTPa92yokrEyY/191JETk8ouy0QN1PwUxADeA8Zy++AEqgbaD2H8M+f
uIUqH+w+puwZ03lj0z0qlm+Bwzn2LJXRI7tkZeYRUSQsVjtFJaXCsMQYPTIPzz7m
W2AMCYT9FrTWaUgCBGZdOHoSN9AjYaZ/Jfp3HY0GCl8ysFqvm3pREn50aL9S/TyH
p0CW9r2GZ4EtSYEKaDkkqrhUwPHmeztv4MU/0gjgrO/rjGcmfD4XKHDkznlrS5eZ
a61SFXr7qvMVFmmwtH7+K1kWAOhiifCjI2Z5mYzrXbRxfVcC494UbZnRjwp7mqCD
JgDi5cg36n5gbgXcZh0cnjL50tvrycJM+nbqPwlJwkVqVc0aclYzwuI0Z6l1G6Ak
fMiRWQdnvGjxq7iq5RjtzXZH/g1PEHZ2mNVxgJbSUZt0+ONaguZEtNo7gFobYwKV
qu1wOW0zzIurpZYsxvUgJHrtJJ+XM83tgHv6iYjLy0VTjhcY+P6atSi7osz7azpk
YesltoCHNk2hjaLQzsizNR2FiqpnJ0tX9m0WtWlPeSAxl5H5WpBZQdMgVNEXWeAu
A69C0VTx+A0ei2QnbfOvPKjju1gU5nHgSrBBFtoV9CQeR207Ucw+UhCDjehncXrC
y/An93hBLn0n/2++ywjFkiAnurC9dx6GPuYn0g3EV0i3PYvBt85SkVTySYpRTYxG
IYcVfBr8SN9K+7VlTEqCzmaTFKgjRb4U4Rjw7TFcNikCWRzNawhwtEC6LJVMICxr
LalC3LIn/ir7LWxcqI1uTwJI1Exgn3V0p08Q1XG+vNP418mAl5RRm42wTr9vc3W3
vVhnVwyK5vWODzqxsWeXGSTxuD9JXWrB+raK3IcsvA9KHwi6aQzAG3v+UnN+HWC0
0eQaTlROAlrf2DS36AmaSJQ/FzAztlA4MYDQayeRfs4yICXf3YPo5uW2h2YHRszX
XQQCZT8FJB9p2n29othG2zuX9gsOv573ONlL5mtP4MFgCU23atsw5oUw9zvc8SXi
znDo2Xaj3nT8m+E/JAj6i/nbB9+r1+2kan+yWVLkBxJts5lmAySqLsoPcqOK96BN
+X1D67tRq8/x1kPEXR8AZA9CBYnYs5jqDW8gYAot/h0rlvcmeWQjKVwzkiXjjLzm
UpWeaVu834U5/X1FJHL051OdPZkeg/TsncjKN9EvgkSBquPXuWWnPsEh3LZ+P11w
vpGQq0xhMh4ozNkcFMkL8A7qRsu201MBINtJkE2iqZ08mo701a/KRpXqb0118SYO
kT1bW9TJMspu1Kl33fr4dfIWKuVeEL0Dly/e6G8DkF9hd+gjVyxn+tJGjB+ysN/H
zdAXdJ02awLcy5i/IfXPntVzeP2XmM7IpjaC3NU/ffHOc1HY8yjGSLz6CB9EIkL/
ZDx5VCeCBMTZosC2PDQO3TGFkqAkFqYQhPY0wM7nITR18i5zvbecekRPnO04fY98
+64tb6QiN5KpdXpgPl3RWabZbKybGSQPpv+GT7rZT5xBa4wByJ4Q4vwC9Nx47dc6
VU4wkxcVLbsL0GofKwN5jw58zGxmFYpBrQNMvi9goDsxwafD2EqV71XW7Ea47NVh
VfoUEAYx/17pK3Q4Rn9FX1oIKz1tPNeG7HlOVE/XCr3pxbWmxS53I35SOlL+V8OK
4nVBG2LXkhpFz2bf8hqHGKeyDzsY7TacK7OFiRJy2xBAP6u71cap9/QATLrd5RIV
A1OtTuajxHqbf+q4WSJW0iYDVv2zk/1erinMvXLWQTqTodyggJtPSP1WJV6w8RoY
pkWf6lkC+Z4WtsZk/+u/Bf8QgfAhyXYRYoVFNPQC2dV/YD/fWSNEN4iLpPrdOUGL
JE9iwch1Atz0rdxNa5P0VYin5ZYhghnrEkC4TMgPUy6k7E69Dpvdusvt8+xqPLoa
iKWfiCZ4dn9RehdVMH8NAKsblcyuIIDdymXcaPoFZrV3FFybPnRofTL//rUz4gqQ
3dfSB/Wep+olyi2b7R0qvLpKf9jP5HpC1k7FITYBfC5UtOzVwhms6bkzNe21gtov
o5pm+XBbbbsBZJBDJGForuHCkfEu2QusrwJlNBL0g7Zr6d5rgrylEfR1eqDzZmr5
mjU7I66B+D4cKIfgQE41YcHNNGbxEmLncCU68VELpF3BsKHuEwFByNlB+HaA0BUF
6fP3ljpS1SED27STNhZaEl8cGjf0tKyHO+9/ilH+wGAJEWi2Q5ZiSDt0OxGIjU9v
kWwjFzK/HMIoO2yGr+dSCPqULaFFhkObxy9oGIyR2YGt0Xow4VC9vWHNFQ+bvyxi
/uku+jBVOtCYebp6bwhzirsmR/aIpEwD+gThKGe7xAyb6KrjmKVegdVX1B2vJJzx
+1kvyKkoM+IOA/A9FwLbX34jz5PYwslpH/u69ukK2KwKC1u73rfN47hctURVcP9F
9sIy1zdU8p708GzHgSzE1RmhtTfOIM9U8/YmeV58am5YWP68zDeJSJlKtuQ+I5Pd
cg6wa2iMgoLKAY+FJj4fJNSYvbJCZ0pdIj64HgPkP2d42jhhVlpkcEUiXc1CN+f6
MorX7j6hbYClWdH4MimnQjxXAHXYG7gDtXBk88GGVht9OHpVDaGI8Z1QQzMsP7pb
phDZsnQdb8fONYA1Dy+Lt8n7lV4gE5LXSPIDy4GLFj7mGBjUd7eMQF0Ln4G3bFlW
jKaymMFQyuRq04KiN0EgUjHH7Ki8aApnb9XE5d4jds8plInc8p1Sd1/RocPUu1uz
t5HCdLqLiiEC2V4cCqlcSwOZhrBBNMC4I8KWn0it7u7pe9hb7cKlFrUIzaU5E17j
km67CQRsx3nI7ky73c0aM4MhqcWyj5q48PxQuDkaEWdPTM8RjnPe2ueG8aVGUAQo
dUQjs3v10hfjf7sIhgHDzfhCD2sLQ/UgntOuXVtoiq4wU80//v1gE1wtJdli5O4N
tV/PkQzejonGJprwWbccO0DZCoarveP5zY1rdCzqK/Ea6kgnP2CugPSy/kyArRBL
CKMywcxOTonRTZSJcCIL4dewP7ms1HLdWdnwxH9qBC4rSYAe9dXy0g7GhYO2dqii
bQZnM/c+SxaP6Jyxbf07MXWu4Jk5ohYWCn+2cCJvUrUmhp4v+eYFTS7pM675mv0p
+0004g1WI2RABQ4Izga1kolCg+xqahUupzxo/s6rJXq5oTdgcAXniGnx/BbRy344
rN+L4h0OYcpUmhgBYEV45npFJCUwR1B6WbXPp6IE7AIzJhMGLSSJVTBsdgEblWeP
xv10PAYH+g+/nVRfi5zMqvfs2gW4iOV18Mb3jbeD7zy2cSFnnPQYRGC3WGSPwN6X
ushYSyd39nyq6qvCDyV4iRVZxm+M2b2yA3meHPDS8kczbtEzYsCV2M1m3GyuH5Ta
zpcqAkSev+fT2+KGbaJpMyp/m+aUjyODJs8tt8qcxK+LY20H5boIIucTjlAMI+2k
+8H5EpAQAltCTj8Rj3/rrNYhyhGgzyWVOhtJCJHuN8OGgI4viLKglRGhHpnso5Rt
fqy7A31NaSI+FLjSLFnOR5KOQo3Wm7jMwS/a1wBdIV97AvDGCGwUHfTFmvW7ms++
SoFVSgZw2t9ycnSiQt3pkEZZOA+gQoQTOcBhtBrNsEEC92c2/el+Sw+DgL3DPXEY
COLid2N7zDaLTCOzdSlO7ZfcX/8TlDRisF8+IUJ9Lb5Bf6U+tPiOpYSabqaf6weZ
+1CdUe6jzE8+uzs/F8Qn936nhFh8sTvfNY8ss/inyzL/S+RWydvM+Tnq22oz7YhJ
N1mcoVUpVqBxYm0FxjfcP3UqOKSfXBpcPF1V2eQgCF2ZPBai4Dj6xpQSu0OhAoGt
YCWhvXX8wQpuwXNXrJ2h5aZDbR4IsYzXa78zGe4mwY0jEQnqFuBfMpeCyGiTGLeE
L9YOpSxdeNPO4c/ujL5MnMo8hyiGLzOh7N5E1MWNH3DuQ/tQ+YGFDrjibrlAE82m
bNOzRaxYwiWOFdkdIkk38m/HY2YW7o8Wd/ZQ1BGGTSivcxYRvSL55a+2ParSF7af
27F1CJ4p/Rwd0nHDEtF96fX4qfvlD3fBCOVryV5MaM/KtpQULGtu5xgGINy6ccxC
VWtxD95yD8uPO7gva8scQ7uOU0bsKLDzZU+KUYQfGgmBULLkqYJiTZgmpXM67rI5
OjHWi2xnsQtFlMbMhVr/W57il8hck6AWq0vtsClfgSubzGhSLg/KkzJ6w5UJZejy
+naSXARe4Hvoo6BNzJIABQ8cERsFhp/zGZueH8NaX2/YaVYV8vRFXY0xYGIXiKU/
IGcLZNRBX8FNQ82u/hZCHPrmE7htW6vF4QtTecA7L3ot5KMSz2Y2r7i0CHYq+hHp
x5uyVEwHlwPyjvMWSuEBlluHv2gO/54YjJQjyQz5kRrZ/NcZaAogMXyVQbmPEBzv
Lnjb/Da+1qgRZfIm4A+zyoEDiM9XMJtiEQptJr/OnMM4vCVxhh098XkOsnvQzzWJ
UvkOxukUtOmnuc9E/k75yxD7veVOaMsws9CMzbQaSU6ougBNdqmIfxLx+7/Etw0r
/NlJjTz1qyRhUe3DA9bl0EWkcFRaEY6CGv+poWqWYebvVUo16NCgwObp8FJ3y0+J
waNrZkC6HNwsnvZU2fs+mmaW3FerH/7N4sMSKWeouFaXDjNjT6pLVeN8t9dhi2cq
px+YVaxBE9+6w7QfLijOkVpqICeQBzJd3VC7hzEWX6Gj9WX3BQoOVKZEE6P/OXTP
ptWzujo0xibds44OB2iOTU4kaovknSgV33tQnYszGJ+jPyxXDQWL8NRWg5T/NvIv
4/psafxcbolk1yg5veL/H03MhOP+C0VByrYRHCl9PBY5TY0MU3lC9h9G/NAABWlb
VAarG9y2FMahLR1Y+6iRi7wQnBRleo10ufSA3tokrGbehKgh2D5A6fxBeJ6rrhpI
yr4D956YAk0+33lSc0HEdHXAQlKP8Kpovozi0ih5kd/e81+c6qotuov2+AXg21nQ
ZjWXJnBpRDNwdy1PfC1x/iBkNBuIZU7HDWFHN8l1Eu+4n3zVyZhiEimCCU/no22g
IWJCrLpeGxuZCjd1DG12P6zSJYfxsVXJkD2LoPpE7ymYsvkfLTPOu7jXrBANTDyj
TWr3lNs/zO3pyAfvWL59MXNr/n3oTtexpwofXDSlq70iJOKhZUC9xCWZNgQ1M2/K
UrE65GUVZP9E812k81iR8UjMWXdUHddAw3rKDRMREK+oXYWaNVobc/tZCrFvpq0B
mSJZAVQvTfvFBj78XKdyeVFGHO1yS7GWEVh52aqa/Y0ghx1J6M00wB/IXZ3/8LqY
QPKBuR5LldyAVt6lQDaaHRK9DkNMRRPHm5bNfDSBHSJeogEcfSsHt0fS16xpdRz6
ZTBjWo0cdxH6lgF7YhiJv4xQXXpqQeSBjY8upMS8rJRa1am6+N6O1242GKAaoCwb
Ar7tKNcnwFni/6VCKv5dNX464hFudoeXjNWVYDWHeT1ldXkvOCS6ym7VZWlqNX5o
NZT4J6aCZg8EgGdPi2UEt8tgWJkdbBQPac+FJSfL+ZfU6UwOLmVvuuqoVW1bTMv+
iz490/TnCSAOV3sYd+m2sn04LCCIah5lJDXWprGB2cJMIjDh1ow6DAe8AazfeJJN
cJGFQnj1GXJNQYNnlLxhscYr7I892dcM70J3NWp2/utLJhxoeH+TRca+Yo3HQHoC
g3aQ7yjNmlR5H05L5EyWUlYwq8QoD9lLBs9yvLSWyt5jIHOut0Jb3pZ8Dk0vhpQC
CkwNFAe+4CT/ZYKkQo9/+9b+eHGPiI3JhVvGeEzRRw9WgGi5hOacUz2qCYxE6wGY
aqPn4VDCWx+hYK1sT83rZvkXF0O+EziZ6grUBjX5a8mZlf4bQVwE7puYwENsStiY
/EHtXk0BG2pjB+4z6DVCKslCPTNoYBcI/7TSIhVq6dHcyQVmcwoCLWn1y921sYK8
EupUaTObmg9DpQZX5q5WdOEp0uDd4uJX5zUrx38/VBDR44sbRob4HUXf0M1PT4FT
/pukyXAPMih7/nBIMbAxxY5ixrvjrr0Wpf+DFqR9Wb48H8IuyAUcZSrUo3QY/Oy8
I5/3rlEsI/acDLh5CNsqeVLKq0b/ppQDkg81lbBDiOkWziuVDsl5moAa1tS6M0tR
oFu2vbHX6phE3nBtGdVJYR6hMz5RzBV8utGdQW9D4HR7nGizTmNndRXUicRv5ueX
7UPIlu+ab4ltfukDM1Pc5XbtZLHzpZdBFT0g2e5wr7rnK7/v7EzA5S9Re0vCSV3Y
9hZQoJFd3GwCXgjUzqipkAct2z+lgjOcZjnRoREeLhWsD/gPXFGTJq533ZhPEDPo
QHlxjFv6iTS8vLjTwKRGGCdxXajupMxLUUzD3MmmCAXww0O7pPF2CmahCSQ6jkI9
UBRp40YGfEQn2nBbRjQsXmUQNj5YK2Fy+spfDzAf8N2IG9tcmsiYFfRe5Hp5mu8j
wglcZx3LEK4l/iV2GrLNQla8GO0IG+GzwUFPiz2K2IZUy7Vpn5felsMHEqo+BiCz
2u06gi3dlNdh3JAhQKJDqsXM/IT/84pc6sAWzkOXt2Fz19HoUEEnMhEjGg4rp17z
+D6GbptpEdbUDTGGXPmgp6OXteFolB7JCwNh5jc973m37Mrbpt3zwYBTEJWVAGWa
KJwANYWgNEAYIqjkRqElDCTvXm0xbvrvAaE90S2t+szkN0htrd/RdFmkC6YIjZ7R
9naHnu8faYHIMAy2SD6xCkf1j/Z/8XHy54y6zUfcj2DrUho9AEU6ZBYkN47N9C5E
/pykL6F8ufx/9nN4AnreEJjbcv+rKThfJIDDSmi8xr+IMj81YDc9eLNcAovWfs3k
u6eXU3jPiuTxNtW+uWvh1xNnYfDWeQnRFqtjKvM087nGtrFyLUsz4YrSocL4BPvT
bRNk4PJ1PCJ2h2e87AXFBhSTs71B30oYNhHB7RD/wdVBuDcV0FNET4GF0873MX2m
uVvIhcvYOLZ4rKzJc2T+lT9CQpmOb5HsOSvcwbj2/fLGY7GbEUHitmHvpj+ffLZ2
ubeaf9Ni43wFd/jCcF3/CMkhYfsbkBnetvC34wwZx8i2cfdRJSLWrVZ0xPLbIO8w
iLl5EqjYSSfz55XtErig4+aDH7DtdoiZLmn9iCWITxX1atfSlxGCZ2X+zBO1EElY
CaneCB8nhfvY1d+ci0KRrU/L5+m3sE8z9vkB6VoSRf16nwC2FVTNdwwHo4bODWEF
ngvX3s6rzwFx0ii/MoUl63JowVOcDEuVobwwnDp+BbhNkOUagBwo3H8DKU3MVA4n
E4JASxN8uXW0kSI7wAR4qlwYBkaVaq41EavzGsFHxOSxIZKg6bYeCipHMgM9YCoJ
3qp/n6wZNagrwcUn7FSLvDaE4fP8A82v5nnQ+UvW4OQ+R/oTnmPVyf5/SvG+Q4XA
ZsyJxnyT5U09nRhNEd9xIEk4u8QVN7Rd0faVi5XcVads7fOTasPNpXihN5nBRqWz
kRcWhjsBZO/UCFPtSP2eW1vESJdqKdTmaP6bEodH1a9IsoedsWL5Wq/w7+Mb8q64
7vDF2VAPogEknG4rLGZQFnFM9XHBq1F1UScatAhG/K02PgEwh6ij7q0uUfa6sFS1
dYHGi8zeiWNcsKaMnUK2L/GrxYvxGo6wM6vdpeOrlZjOIV5p3ccbqlz3y8vpo42t
yCEglufWtB3aXStQek2ODnD8MHMO8u8btIWIXMh9Jc+ycrZYtoRQHP27aRUBAgxe
nCdEUVz1mwOAMDFpgEWLaVVrvHdc3ApKd/GUZ1pt2AZa8jLGwrkM9reYSK4rw8d7
c2y8r7o2/oEtki9taiJRn3zZaQV4X76Mv/jjVcFsDr+Y22HwAR3ubX1fXPorj0Em
8Goc+NvMVy+JRUiMkuFLLfaUuEU4o8IH45Z4kmkR+yoyBNOLQ5tyMBGj42dSKDgX
qfulhzse4R1GD5vmDjwTVPZGUWUGezb2am3V9v016JF0BFuXQdEDCQb2i50rgSXL
ofaJxmsNB3vlofYCgS9g4msceEHEQxD2YuUwAoBvKMNK74mLISbWSSKfOyosl/Gl
VTVuhkf87rgIbQ8ugJVr/PUk44J4UlJA2QG+R6lWDtdS1TuhIqE3KCbfP47Fk3HM
nbTJpg4JgcBBtRm+q9U0UObEcMIeyIkOmnjborhddfBiLmnoaozzqt0xDUQork92
h6u/a/KZWey/PDvRlsurpffwgGHKoMmNRq5Xyvruzu9qwlNyh3A/1chHOUwMaCoR
lxOttaAyT8/tDSNfwAG95d7UYyxHhxCmrEP8HoNCxw8gCosx8I0PBh+9kmhaZIPg
lANbcixRE5XJxKMwz5OveeDSix9yI3/9rLv9PYyQb1BMjFWhD2pCZoO2iu0Tm+ug
/YzVm0C6Ok020PCAuJvUmFLSwbG/70LAtMWvrl/OpKG0V3TVggzXh69aoFGRZ0ri
9O9tmVK7ATVre7/tm23ZYoJD+2UEyqFoYSRiFF4sks6yYPEjeRDJGznqti89NH7I
AFMLqZnpBy9lep7nkIH5EciS1iZJDTWzEP14k1Rd6155DhqUDrBX/3rqMADRToDv
TzkCN7imrdcp/KdNUmFXUEG6sde1OjCsZN7WHcjVsCxeD/ZA8Qz4NNcaJbiTkl3x
iw2NVg9KDXiPEr2zDAjH8REjRrSvFATd5PAku0nU+rJjjmRMDMKuazUPk8h0Vn3F
cJbo+Sg1dtAhQVxkdttLPSE2vHhY9nj+4N+9aHy+DyTTlX2x804d+9XkDZJzSCbQ
OMWBhMcYY3GPskllPBZ3grz45eC6u4PC38c/SWnouGQwN3d2A0nY3CA5LWJ9RpGt
dxVn967O3fm+AMz4O5iXcfOmBbcCqXCiZMdKprskj5FfY9mf9iV2aXAgHHJwG/ly
dqZC9OnsrdlsUX0Iw4mnhiUywwPUfsKAYIDvjJRxusB7UujRyT5rrjPmAN5JhMyC
fVW5+KCBzSivBA+h2BtlwD8PTLj9iYHWZ6EYAWCqzqJAASTs4HtYtNB59t5NW+oT
N9MJ1AYjW9eYB+VpX3Gu8xiOU5+iJpOkhjxx7OA/Nq0in9J81LmUtyMxDOBt7Jw4
HLpBQ+fiAAlBDZD6q2EhfYPvrtM6pWzJWZwtgwX+eLpXj8evu18Rf0b/1IMeqma4
KCZVAF7W3XnP3SHrU170tmTtCtmXyH0bZ40741a8Vxarl75x/O0qH7cuSIs0SL7p
JZ8vdrSehcsiTeG/ptXqeu9h3fbj+4RE65LMurgq0nbypjp6L3dvKs7glIYspv6P
H7YK5IDKjbNJAmM8EY6+nRfFfuCGfpGNVKH1XYeOPDiZH3PoqUti+F/37gJMqYFi
92Ygbmq/0SReI3ggamPJnVqTkPhqIhNTp37Kk3cgppBdWlrsl+mPaGeuzS3lRw5w
wMgHLEZQvwhmwgqdKz8kUPwdPjdUdirRR0/MZbnkq66ZsqnrvErYTnVvJHOQi/rC
9ex4nHZ64lAyMTLWe37gxS2CmsM2/k1RZQKVK2fBVUuVsWG+EI2hDUb9bQo3F8f5
xKMOgU2RxYs71WVzsJJAsISLut6VC9AV0hUWEMag18ePtpYrFdYdpK16ZjJKu8BO
Vkq6AriPLRPMTzv7RffbnMU4/ZiN166Lw0QjRdpU9ClvqxLRq20Pr68V6JZ32zVK
JCIUhGqHcySOlSLrSLbmB9rRjMf46CNMYgl71pTQCHHs//9brfRDEqGVdv0Y+BaM
oZH25K8fR4wxXilk0odSVt1oXgyB0ECHNChYGepgD7i4j058z+Fg0Ha5Odo/k7pf
GXizWKfwqpLi5Vt9etn0z43kpyuROhn3dcBH/LRxS0LZZtjJKuaF8zEEZYiH/ygG
85VdXuWWFThSYIl7AT9TXUubCIN420LD7H9XQ8k67dDjmu8/YL175ymgGJ8U9VDO
QUP06uH1neTVztYBqW0N2WJyXra1YbghYttXZe0BZaoJaGBi8HgVXgrMfvy3sOEP
UKfzcjNL5XW58efpUM32uBnZG5qnJsswHs44lkstxsXXaOoCsnH1+QTnv3qVQeKW
e53le1kgnuc0JI+WNoXxz3tDKAPRBHHJvBqpBH99iQNkk1XeUYU+kQNAY2N99J4P
SHEUQxYi92RXf684aPy3PAVABiGc2JXXpJ0vqcncz8KU0iA3MsxFiCwACiwgtlUS
UZm3xx6/0oJjGGI8V6jm90s+L5+pktyoizdLuHQ8lNI1FV4irkRXWxYrOIlRTvnp
8HtQGh1KKhyLcqO3MGUDClT9vmpxY5Z+JmMktpng9DZXdym28ZtDzjDheWUH3tZI
8Pq0ZbqLV5xzf4jQ+VgnOxqOK3RoyaS68zfbk34UVaPuk+b0XJflInZ1Bbu0RPH4
kiUB/vNCmdsffgO5N+0WZHEkgmEnByhXFoXeMwIxiBkmMcGPBWKWYtbw7a8Ayg9E
HGbA2RJJaNYTEUvFAzb7o58vboM7IA2i+Fw9KoZ2cQ9GQNSL86X1AlVJ02K+zeRb
3J982IGZNDonF6MnUg52VqUzdtwRxVbpPsVY7XRJ8xMab/HWQxN6BI6m/0iZRDUt
zK4egkKzR3L4aIQrpB9Ydid+UUZcjhGojOn/8kDkFIq2NYFRUIXSCi2xZApxAmJ7
2AAEnOcx1L509hUS1N2l1M3eMFzKAOFRTxzQMMr3y/ajLRo9Kd/KP3GX3Fz0RFxX
cBmcKsRUQxb6czu/yOFLw3L9XSvMTsob+2AOrkUohJ/m6ZtnMN4XNVU42Jw+k8L5
gzcJkycHu2uTzplSdvznv6lx42tfB5ondinFWidCYtAGxS3WVL99QMxmBVL3sSIP
uq8ogkUq2pL6xFdlMnvk8GcBzMrHL1hNcY61UnmJXA4lR+6XMUsP4D8SaZdfhERS
SCOe6DKinz6wRHIgiyXH52AidOtFpPNQVsZa+fBaKTMsbTpbYevPi13/6FX8De+e
ITIbWOkM44dhsFk4wuZwB7NtCMfOdiZ5OGUTaVnVRGJJ4pyTQp6fButG/X4WapR5
M6/qxUFdmuFP08coXD5F1WIOnd2PY3jcTOC2nSgs3aoO7lat7VYMQqEmXVOf+wE6
m6JqKecD3TA238BYueMEny+D5h+SWZxLPAHFdjwTAZrEcnZztnBiJgK7/cy9QExn
V3A695QYy65HCKDHr0QyuBeDVKl2IroRvELMw1sUE6IqopiTQmyZ1XsL1B9TWVn3
nd+jOX93+h3PcTAjMo30kAmX8kbj+x3e32u7G/1CVV2yUDlKHr7NjUPSKHJUIOnb
KE4FRR3JOIabpRqWzE8NZH7B6ZpGqq7VWfQvc+/tFpGkNNthcn4nHLMUyd/m6ozC
Z+TP/JTBIqYEdnI9K4AqYtj6U5Zaw/iC60JX2YY3ci9Lpp2l2i6LbJ9eEDmTHZNo
F2mPChWLq/RqvolfcBlibCxdnkdHcpTcu00BGTR3Pld/bOaPMW9T/7hWM2oZo+WX
tiLFaEee2MuOdt83nCd93muvG6gp35N8XBNizORA0KgEx4RcBDBokqFb9nMJASZC
RvRPefSQgQ8mUf9e2fn1TgK/6AUTVEHE4nbWaQWMn1irWXUgxFExb7cnKs2ljvOD
X3E8p1EKkxo0wn/YFAbMBmGsPeJ+CO9bIj6zYxZIM6HOGP4LFBxroRcz7vYMAI/o
d5d085AnqnFv+bCsbXvklLT3EI46IvrE98OhsWXyu4Qcg9sjbj+oQ2dhHds6SnLr
sDUAF2+TVtjtwetGRMP1SHoYw/2xOODKNLZgANk2M7sqkRoEBlCBYogZ5ZzXEb74
lJoEI+WkQq4WAl5RwgoeVsusCP8lwVLiv/peOl5Yv2P+w0GL9wRdzVEzINhoNJSF
Cpw7bNxR3MXCUZ3EpixgcuKss/eEj2tgNKrQe6B9yQDlWyWP6v2gs7qvLtPY8CnX
33ymtNXlxjylS0d7XGnkZWgQnIVYTlSKR6Ac6lHr0iOMnsizY4AjVcnW+NTLeP1O
VO71Z38mE97fyzcNWaS3ZRPW4XvPDBlU8QZcioYphaPCFCHD2SUmPbDCTrl1g2hP
VcdNQlCZEukzT2/dkN4B1C8vtZ3A96Ma7WyYx7bu0VbJt/X6qR0hdQ8ncx7jByMI
+V89pIPX25qc/Qg0TY0+5YOZfaptCcpS/hES9dhhXp+A5M2XkII1IKN18u0a5zqF
xXqhsQt7zBifg9wQ4HsVnRauu1sCVkLJwweQ4BI0quFu1t6961Mq0UOi9GD314k9
b6HF9VM2VwwNk98vdpFEEPOghSjcvX333BEToQbDmJJ7/7qXrpwtKQpe8MqNYA+8
j5lIYsQaq0b2T1IsUkwb5dPVOMcVnz7yWcC9QpO6tpPhJZBmaawydM6xfFQznDXk
L4pEiXh2fDDPd5TgRGRvZy8Ag91JZvPMxGYgKbJNd95sEgTyMD0BSJ6H2GUkV48p
/DdfZu1u5ZxtTDFd3gYnZ7hXVDLRaii9iXZe+IHYxAUMvWglowXC0RoX/ucD3m0j
pCT4x2MRVqvVbmapv609HJsbwvBzEQf3MPMXgtvTpl8x42WN8M+xL/3be6shavHF
gTVJOoCm//iSq9mJgI6kl9V0c8o3s1ogsWv3IvZObavF42ouZSdv8ZKL1FfYmJZ4
as09kkqoMYcrlrVSojA9UO6mBJ5+MnOIky9bkRF/bZ/7viKwF8rAMJRBgslgOr70
n6GSj9EI97von1FXIgwB/X0a/Y2euGW7JN8PQTJuUEH+aPCTV0y1tiW7A2Y8T+Mv
QQ1IGEaJkr9vdu9bCSayc5SaOayZs1tiKnbcNQGTt/uc5UXCLGyxjf4B2hGoA2fD
Rv1RKUng1cOL5bjN29sWc/9tXS5tUXGM8+Bezfu49BidDKfyRCoGwMEfKuxUdRcz
6sklYAgViUwxL+npYbegnQ0IjXzhES9mEWoLs497Ax2miogpMdF+XTRLrH/Ty7KC
kn5niDOaN2+3Y0XpYd9/LmfzM2Ze8+4vx+xVrQtMD3OUGYcB3c6DTWphOF5RFYUJ
3PJOuYkD796Dv08q94K8lT/59IbzkTnqgkmMxd2dYPIuwhiU8ru/8zqSGaQ3AY9h
mTr5imPLECr5bF17deANhTHm2SR5a/JAnO4bTtbaCvRR267WgZIY0fLUYmUf76zd
tZyHl81Svf7iPbETOpxDGzlctQ6B1Qkao1nkzu0efQWvXL/HGHaIYDpwfYIgm6KB
0HPGCTyxFkuJu/9tYJlvt86rSvwwlkcGLSedWlOM8qeXURGElCaSRtOEvQ2a6efB
pH4pnwweO9p0xWJMkdy+URhhpN14oX9dZyzJrLqzxKRdrmZS6AZNpsSTjfRxIq/i
3r3S0XeruzeIQ+m/91xcJGjolY5PqJU90r8GNamwTS2RizFzQe1DkrJJ+7nhKbDE
7O7fUTrqWQZ7tWg/CIkcsxNDkX4snjvE72gOxGzKTY3t+AouIrHvKA7dhZR31P11
v2EPFk5E8THbFs2O9xqDIGW9QqtX9ZxHMbquEOBj1A6i7Nh2WcS9vPzSgCcI8aY1
p1jnfG7nEwIqwoqm38PQ4JVN1sVRW9ndCgRhSo7rontM4KwOpiCVFSAOhn686IjC
k+RMzl43uGl+1H/VQ/qfReR01NTPmnMl4Jz4SQxwEUoPGnwE5Hm9xzLUHXL3je/y
sKMbSKzS4wOXLeXwtxjhTuSMjy4VSwSNCdgr6F5b3rQJCPHDtHY0SJVGGyNshmN8
Ushfm6+dsGWuwjaOFfFIq+PmHJA9XJoWItGzhkcbjl5LFYBswrI7UP41xuHWLLxK
OGjT9sIgMVqISC6D31EEA1D6Vq06m24rqhlD0W3XPSNoY5MQ100Mu4n+rH75e5Gi
btZPMFhlQXwrr5rwGFxq+ng6By+4h6IW5GA5RLLbxQ2PD2HQpsiIhFKHvBD2BvuW
8Xd0Ifl2fEeAInGJ4irJo94k+ygnKeUMoN8b2rnzx1aLQFt/g4J/muu9n+BNe9Qp
8sqSCZbf9aba/641PviLgu0eR+x2Tu9kFdBjmYJv1F8qjz9HFX8Qvzk+6Pq4mMkQ
RMj1Vzq9F767Eq8y6zBadGt1Fi/glG9BAC9fE2HsElQ8R+Fc35AnPtUUF9IQoe6F
Z9RDi1u4AQy8v7YIszuxifj2Faf7IUUw01EP6OwTUyLVyRvbxXbyM40ePmO8Xyap
obo+ORRWaM3lWDQccwSNz9Wm06oo0jVuKKC92XG+jYG5oI3hemx88Kbq9U0GOU66
R4Kj7U3lJ0lRx1w8lRa6qbNP1scYPG5bMV+H+WiNN1Rgqq8l6aBDZTng0Pya7MpQ
hmA2dqteX0KKwCT0SzrjVP0eIPCL1XGK2S4p5wrorzvD/RkukeSWxIonwN/AeTZ5
5dSipwXGhDkodzpnuH1/ClA8j7ov7nXVYUq0ZyzxK7ftrS8WAUl2kwmf4HxI6Yit
rdXYCLOyBZ3Gvd8G5Ub7a0qDDOv6+Xcl4gDpd9HsYSH9qcId5KPG7i+XE+2GTEv+
4ODDrsnD0jGo+W/yYv4ZTAErR4SiYoEcCtDL3uKLK1R2hVsnc8W6uN1E49ggYjEE
XiEnPrNdDeYyXbj03wZwi0WayvoIScACFF+Ag7ofn+IwS5aJ7j0qc/SxQruu1hIN
jYbUuMzbhS9maerNJs1802G9ejefTdJCvqF9Glt1HMX4GrSwPLCdEgcUxDkIiymQ
20hCZumf3ICK+7trRJz6Ad8zEc/5fA4J41KO5hIPQ5LfKfW0iqDJzCAbzeKCiCT7
iaT+QHnBFVO2S7XKkLeoqdagXiNIqf3/K1KPofoTJXk1UL47p3kOuJ7Bt7xpHIQx
gFVHAcCV4cEOQoRTHO8acnuuvhYnzQGrHi0y1aAuUfn/QiJ1fU0zk2lh1BPZ8FPs
2cxqEnTA0qj/vFAxYbP2o4eOE2L03gKvZm3oObaeay6aUaxeKzhjkBeC94bEU9Ej
bT2G7aLrCz8LJDuSt7ulkQNX9sYAHNRRzqV9MbMvn8mh7kp//rvWyoc33Bhb1luY
GJAPgrzUzGsvSkZxTA9kcuSAn9NuLn0jNjHFcqby71sfmwrXu6I/qjZHFN76cPKk
B5gxBkVWhN1xi5ZDo7SFYV3bp+i4NHC0ZlYlGZcw+RsIMm3mVyI0stH4nBp6XU8W
lptPZuMteWlJALz6Taxm60Nlgu0eos2xS49yUQeCZw6T1bUPSdyRF1QL8pOvDaFl
8ZTm/jwPzk5BgldnVX60FBnvfGJKAX3Y8XurOgFuUHvAdHLxdXFiJ7W/6lZXXHbG
2d1CHW8V5naSns31Zf1RUn3K93dc4L0Rxrh+HGtnr6vtX5v0Qd/ngKqSUlbRYyzE
p0QtJSeiVVa4DBDUGNytdTzHwdtSyohAaSxVLUUFJr38P5ASHZt+DFuJy4mMGFDE
9v+q94G4LPTak0Omb79C+Tt60aGiVRVoFJExkf9RBGMCxNrwnm92pN+g04f5V8HZ
Fve01KrbWkc+EwA6P7zM8/1fv5tsNHY6+i6rucp4Z/RwsfX7sxlwGe5l21eCMJyW
14ZxvEgHKtOwEtQ40SdhDGrz6HT/3q6I1tdxOu+IoansQ/ga+sciJBfIU6OpPiVp
KSfwsVENs5Wrde/VutfPUXEdgsJC7oSuSkmqthxlz9PmOwRl0BS+RitN0PH86JKQ
5YLs88Qdb66d8cpnRNSGoQKLZKgGgKXCfWECHSQYSCoihdV/Jmk95/x0IO8qqbDC
Bzb3r0iTYW97DD+c4BeStImZ8dG6C/TsQImccQJ4z3umrcVH3cmSWTvQlNj3syPv
K++1UVNwh/LCAi5zENfSnFamLAI+Qf7OWByG/sVfwPnPg9Fsahd4+dLgLLlR/ZrM
n1lzbSUW5NvJQDgQJ9K/YZufwvFtRDpx19g6fJZD1XoYXMKFR4XAADeXICNwrsWZ
7atdZ2l318aajLO8T3jHuVPxk5yISLnGB1xG9uhYML3heE5hWnp3pUETj9hVmhHf
x1rwJtGZsJqOdxu7I2ya/KqiNOywSNc+/cIOW5PsHL03m/PpL+9FULSk5t18l5wf
fkldmsakDebVK3MzraRWLLsfSUn8pHQ4I1uxM1wVQzwmOq4vdtfDMJj1OTuaq+uf
V1i9ZGvR3pMsvUBiyp4ErPpFpDXUA+I7LEK35h6BaLwLd48pexPB1Unwc8dzemPR
wOJ+RSLDajuPaovyvld94Mz35Sw1pwdE2Ru3fdAs8JzAxfMnAZEtHaDsHis8ojEb
Y7uU4TFfAG3M1gqYst/GJXZ4wusJtpy7QFBX1dkcH37ut+csaOOM55yYvpTnWHi+
TkDoQ2qyqjz29dHpSAWPQNX4UdljlgsO+4xQiBbmBv4WOzjIEm52WH67QJ/Tn+EV
8ZiMEzWbNyK+GGtSrguJslVBhvNPb+ZyvhvYT5ElMxU+uNWwsFEJgP4BEuVGHQea
gRPekisL98rPE8Fkvv2xfPUbezumZLLfCJXgSWvZj4zMpaOxOAC9uctz8YfENKNI
dWzZecff4CvmJOxdBExmZtxtrNmuzhoGr5v7BQVQIGsP3Fn/pj+rD+zMB/QLtXrG
yDb323lbV75pdd+FHBl1kewJBabKKv1rEH9qM3VCNlQsMPIzBM3qyp5FkviRTj6S
FfZdxlr2tLx1WsWARrvtcX7ZaUB2qnnMKxo2nB2nw5yNjEhnJAzZMIUjYSSbQsfC
XN2kaymdE2p4y5s0N+7Q61n1Dcu4UeRmtIQbYQ9Kv7Kglqny6U03lDboE9KPkAzq
W9rX6fYIiVFNAzDbB2ZM7mJyZvwDTfmiRHAlBrk6Vlca+7ljdLR2+4gzbTSwcVFp
+csAtgRDv9ILSElCWUP+zH+c1a2L8ZKqEizqeIAg6QU0YxVOOkYrZUvZbKYq7uQh
kY9Q5N/uwLE72vU0HsRq00qMz9GLp7dMi2i4NltOT5/k2U68VYjrzy3CUZS87de/
vTqG/Ieutbbgv0vfxm0t4oF4XNrktrl71K6JG5oKYsDYI6gtJaq+5nAhEjASPXNG
eTbGRAllNX/AbRP092GH7mwxMW9H3m24c5sOPHByptJDFTJJDf3/fuW+PdgDOekE
U5VCSeZyyqrXvz4iIyaVQYnq5ChlANZMsNayVpPymnE2qNr7fAYazDF5Tj+oyDxQ
Q264xMW2Mm/+XiLMyds1Hda2rOoS3WVRqH3KKRzi9rMdMujH6e7TJSXrULOQ53+T
OEnln1+FL2D+fk2OxGdxM7XS7d7ptxYMj6olmGyc1AktOnJ+F5s0s03Kzrp6ithW
snXkHJYUdjf4mg8sqN5my3tWl6ZoJE7MPYwHQDdxHabE2OMzRs0OP+SvhR75wlSE
koENHOBRPHX7HEiZb2j2cLMA4OANkSGU/cPGr/KtbZOggCP0/I0peAyjo+dvq2Sv
WH6sdumbW0NyRmpHmYji7yQyajYbYVXucBd+FB2kqmdTA+eFontli162bqCPjRgw
8B9OP2ck5o7zWEuSB5Th7/Asz1EGCVQIl+/UhBaTdcrs658q5wiBR1El6+H/Kdo0
RFe4+0wAj96oveSIaikGVVHuqsTNyqu/ns2+ltkHydKXzaf7yGSh187pNA/ypTiU
x7vBG7uhIuyvV9OIw2QKYD82UFugbul3VFp7Q32ITO/mrfRjbSmX4/7aj3Yb3NJ5
cQlU26iJzOJjNOKVex0OPMli7sltcVVKEMNtbgdhE9D8QDAcqnK2I8v/ybjzAQ86
T2/CK541uySm3ZtjwsXCZmgfTzOLowXnQkTISOEWQnneIz0k75FJ1jzy/rrqwQ94
43S44OP3QPb90dYfATsxrWKVELpn+9iUovJfn9uqbJlyp7+mAGMvkHHzSHNXGr1K
9cZ4mhyV27BVysjX60O+8CU6mXPJe2+AjSgkRCfDNyB4jSE6RsUtl4DLnuEC9P2z
tLQjk2vSBdlF+GGAaRsbh0zBR1EC21Q2oDJFCeB/Sj2Q2Iab+xIJOFuJwtkGbAZN
VV/bOchMoPT3l/aO7cMztMOAYBdRznxItrnpe7FLzCbYn8eUDLHSO/+m0QWPIAzD
MCCxj6OTdBhGVAJ9dmdBBqDq5x6NJZbdIGvQ5ccYuUKJblT/y9GBLSw81Tfn4W5H
40SBZXpqucD1Ppv1v2N0Ro4W+g6bFfzwdiB5V2HrC5qYlqLfAIsoGyMkL77VpVpe
vxHoCEtno2JWi9pKFCo1HGeawZuZoaY9knq6msQIToIYkFx+qnt1+Quq37+gDGOI
z8hFZK+TOTc52qAtzLujLSJ4/7jQgs07TOuaFIjQ1SkWFrrvfGnKxv5vjxqSI/Qq
hqvBD9qyzToFLUg6Y5ck3b2Lc+RwcH05aTPgMMIRgTclY3kkbMUbrCt/PfadFeCK
8vHzJ1WL/8Uoj/hw/YZYoj5B+joqcrYl+S4U9As9lqjT+i6x0vkVNFt2P3Ube+DT
yPQ+0sep1U4nH9nsJYMKaGf9W83sP9wPNEr3oYAXOlqWtVZDNxeXxtnUn46GCxOM
BU8zof+P471iIzxBG/hofYFJrCD+Weqp78tLlHL5jXuQYNxb52jI5Pp5xnH7jtV/
FeGfR+eG3rF2avUF61rKiszbGiaRik4YBleTXP6S+f+wwCtxZ2cb3u7mB1x/K71L
/LHk/QG3sF1lAy7sM9jjyDfZhLjmYW+z83HZGyNtVbzLcXd/utdDngcGcPUCMNLT
WmQG74UpqrFNcOTVIuS73Bfxa+NoySaNm9ge1ad3iOUJLwRPY2wW7W0OnMKisBT+
yM91DSUODfSCovpQS4Vnzx+K2py5gBXVeAz6BDjeZHUZl3k0aZpxbr4efhmay90h
m1kg8TtcJk8jWjL+gl8uQCiUm5qYVn0X6V/7NPCjNnXT8ItlR6cvHKVvswcZ5t/z
KfmmAU2p8IFeYG4/W/w7YhfI737eqGTSWiQcaPnuay0aluoijJogc2/C9gZnh7YA
s0+nglbmrU5xaWD+IQ6fSNYDLzii91o3OAg2kr5XcvfhIaiKFKG8lV7sD6ST0EBN
+SvJce3m+R+Yi6ffWSjXQN/Kar/f7fZNBEvQ+aigoOE0VYDK2fLZgY9HA6e+psH0
g7aWaGXkWCToFrlJQV1VUuOggAFEr3/HaatzFn8m66MR3z6hv+GCfJj0/XRTo96U
fOjRz7oR/SctT+tBVnNeaZa8gLzyrOiOSWgX7untJ3I4IokJtuEBsyTBB/Ag0oEj
ozVPlkaoF7QFBTYtm1bkpCJuQ9wETf9uI0F1J//Lm8TDZZjmyeSi8V2aShi5qZlE
sleAiQ3GwCU6NR+WsyIH96KdnuauzKQM5Mct0OucU3odTEP8mhnytR71nEeCTCaG
KsBQoL49Qj+f00nEDKzkYP+NjgtcwQ4MPLGJLCY/2IFow9bX3r1dYOpcnJ35RPhy
aSTGXK+xGi/F3eRlRRvWEF9cnP/D7iWq9ZNDN/5I0cK5N9K+hUcLOljpSyxngEnM
TAJEGnvwheFNwmpJX4WJKuq2MQjjCQPS/V49keVhX81qYRslv41ao6HRniCvVcEy
LV6QgCiWes0mmGY+53oBt2jrQ1CPxxXwtiMroGLZV5yl8MS+khT6aDK3dxJFlmTB
vw5zJS92fwUDA8cFtD2rnnWILOySOIJ5pseAWp07go6Pbt3MkVHSHCgH7QREsGSF
B0XavUbe0cAT7QNS8TFlkcb7uARmHVNdNIxw18ozL//wT1sbex14CHhxhNYXxce7
8ZHYcEzt7nwqWXYqYeYfR1qcv+VqzAZYQvosSURKhyInSPlo34SBMBTcv4oVsN/A
4soaQVmepQ5+C2/bEKvYLTqzc01W/2h+0jjNcuuX943MMoxft7XHNAgU13Z8REDX
t7V3Lnnao7Tn3opquOOvBngEhNgGKkdxM0yOHJ8SHLrpEdxQuZRHHOianqsmzxli
AGSD9A2D4GQfyANmauiJ0GxRfkmnfxuOOA/D3muhTHROOdsPsTek72MtW3x0YNFD
A4iI9QQlg7TbB+id+AyG74ozUnzes4ibFmeQDbrPA3MYv5LPGpvfxJTxW0ROtamG
inKNeV+CWLqu5Mdev0iGmfYZ8RS4Bu2TlXXoObh9Ej3DlqjShlq9KLZtKsJqdqEp
bErmNI5tF2GOZ6hT0iXNAbAYKmfIRZ9s+Xp9lQ3nD6/j1WGQJYl96b8bNUF7ClVU
GSpWiII89idsWEEvu45vFKj/jNyqkmXuD7x5s6ncyxpnVyKnr67q1lS4/Kg244Z0
W9YEs2VWAwHEIuQ0e+l1tjRgYGTqGLpNzquNLyCFJnpF//ThImp0UvkmkVybSSEL
vQvRc8VGzPasg97r/W1ic6sokMCjGd47w3vux1b7xc1W8SafenmVey9T3FiCNUUS
DNTAAWr+UlNEzPGGEy6zCwlYgka+mQVduFXzfHCLQ9Es48m2P0a/fiS4UPLceCRp
Ee7PLArHWw2CKsohemsvkbVROZuyhOOKSRi9CqDE1zkHU/D1T4XTzbGFO4elq20t
E1tQj6mtnCVxlWktVw+aBY1n6xC3jn7YZAoBHBjWHkeeP7mHSXV4tbNN8h94X8AL
1SNCD3tXaA5J85wYileS/vkxbq2ryFwdcmY7K22AhU9smviqtJLD+ExHwCPN7Z57
HkQY9ATTnXwL/xC/TBIF3Cfh4BcXjQjofR09fhsh1qEn1Id1YUkQaRK0XAdxAR4s
scqPWq0t8sWnbEa/quhL5yHO/VFLVFQdMZpQtUWJHjvb1QgrgItonMVq6m39DQaD
XdTnwXMSKL1Z91cqK+9upyK38hg5sqpYqfM/0BunrJWrHCsaPdniXFicoYQ/36gk
/DYD2O8p+sxSjCeUxb4VIiTNXkC3154i+Hr0VTxrSSALPNV7reYUIF0RSeAWEv6E
WPp+Yqu0RrlzDV66OTRwVHQwgpuoF4XumDRNywAdZXV3kX9kRHs3m0OGhkfDlSyU
pUgU+F8dXwFOs4hLSLD2xvb49FwAjYBM0Htf+ZzLE62VDF/LbqUmOLuA9RP+kN4f
h4Gji/KTAKrIMitSnRq6HPcfPxf7m1WA1ojAqxfluJZ8f8nzLF0GGdIXr0f5wPnb
t2rvroEoEBhUv3PcgfkXr9Kf0Ud4lOhUfb9CF2TMqEIH5imJx7rC+w7MhnXOy9cb
7YRDGWb1cCQx+A+EdISNNSvZi6M2YjwG985SSuzU9bwginp+5edJaPLFpldehaVN
v8JRScUi5xd8uL4R4BVD/LpIDIeNmN97GsWYxrH485HNt8cw/MCp9DkIytMrFtED
OE7d0UuIGxoa4XjYgbyrf+WvISH4KR/jwzqIdGWqRv1e7L0qWJBgV+hVuL/TXEh4
T2D9MSjpObIZC+iZMINJSqaKKcsH3cLlOY7SE8U+gJ6803IXlYMi6prlkC8wg8BC
T88UtYGnD0aXSeFleUn+YvYznTwNxORTDt4uJdiFMSftzJLs3o98p7JVhfdVfKPo
eDfZa6PQALAOEFohKvo81fg+RPuJUuWy2tdYGGaNHgoqNHwAIG+bsPZ20rZ6yD3g
q9B2Jgqz6ZVYg1IC6JLrjg2+uoXTfA/FrrujzMr+iluEnUqx707WixxKf0UZPXFl
eU9f1XINbf+2c09bD5Nsa0YGRQO+iwN9ICU9OUJ/fNgCKBsV82AfZlRgoN+9oF0j
qEIp+l5RTqdnMnM2IwG3S65yDb/OEUWJsJyLwVUHstXuoHLPCC2X6ulzcKaey4Mk
h6fLioWeNeYiKjCGTuokk3v1iHTHToj1VxhtI8yQlJTbuBvkz12kPiDdR62EL7Wc
TZQwgSb4K1+a6VfI9ITBfhUX8q7ZQf32CDSl0lSdQjJkXJ/hZfeRQAG3Bpt90fBw
Y/mNTkobXnJaFCSJA8OzE1BzzMQLPfZ3PEQeb6yUYdP6UBAp9Z05pYwHFsfdnxr8
8pQs2vpPe0v6qwKRur+k1v+tRlzFxQUI+BOCZuEev8hi3I5x1ega87KvPKVrKH//
DJioSThIO6gqe/jjXZUti12KyA57XJbE+U+dpDo2hFpmhnronx0ldA58/2nqsVZn
wbGgs99W4HiINBuz1GyV8lC1NIjKmR/COg5f1AuBKxXKv7In41qWFU9U0/EbtAhe
jWkBbfN9+tB/G6Etb/lus1aCFQPnkwNsfudS7QTNhjXMNqEABo4H+FcaKKvnnyqs
am+vwQvd6ICXb7329o+5uagDO6CvR8B5IJaKQkoxBlhrh/EM1pgD3Q+M7JvrJcj8
PZYizjqawB7pYxcoxDfFAY6BG0pII0ObOiR4DI+ghPtYGuElLB5mqpBnWe9INHO4
S9G9IuTBCHH5X2GkTZoseRaE61TtMaWYmnkC1PFiHGLNVPW8LaBYuy4xMcD+wSEh
Rn+BNzRv8PETSrW/RbpyljGpPisjCm90oJ49C62luo84q+MH5vaMai127ywm+4Vh
QRIZKgHur8PeU2RtEQ+4Q5upNrHKXKspCKsO1hdzaG7Q/a+HX1jVIk+imbUDrqmW
HVOVDagpH1Q3cWCQ3ypvaS6olv3JvbKJ9CaG5/V0NhWrL7cB1Z5Y+W3KN5aCNa3Y
1T5+VBWJhnHhLme3SmwE7zh3rkFZZBQqAxOnYa+pw0djoSYcUxw7uZ0BimNk1OLq
YDDE3uy9XDCwVYx9ti8rhRa5XN/wSpMR9XRXJVdYI+ZoNvbw+O7vITYF0IpKaqTB
XHxnLC1nwOLDQDWTAAiB7wnebRkYVUEyvRzllo+RJganXDb7kbeN5ysNy2zw2Mw4
kyrpnaBS02F+qxJVJ23kkrh4flQxp3BWvqE1qUe/31zLCchLTiLWjgED2XNGQyx5
lnrehcef1UMnoYIFWgwGppqDtg4kWrMlAAJxYHCyicUKK5zlsc5YwgEfG9Xi/yot
U0DaBL7Fqw+9mAX6tg6FmlCGvGgX0eTOYkdoxrT4TvSpHkk9IbbMpBp6/dxYen8L
UnE+6L874KSbmJRjiOVxbdqDxmTqiAmxwqBd5jFrOQ1i1iq8yUJ6PLGnjnTfvgQD
CX3g/Y9uiVROo0MTxu7BM4gFUeHw1yDGRMjhZzhOfY5ZkhTdEnsetPUZhs8aEX5T
o0HYc5jOutqDOhmHwb6WQaZcxS5dusIYf1AwBrJ2A+bY2KKGo+G4yRYiWci7AZxG
uuZuQoQk+RNlACi3HbIJvqgr6RqK0klpQRNpET6xanvvEdIl7OYSt69JY5SQYeOx
0M1Tvm/0gLRilvEM1y2sX2B1VxUSDOlQNi4nm3v+FtBIQ7YSUf1INFy4kF9KrGR6
5yWYqjUrs7nfs6hP6mkcYXSFyx29ucmV5ahjulUrx3bxfvapFnAvswBIl7vNpsvv
b0Tp2iOQ/yId2Pg3AfeDs6k4VIKn8iLqfCKgSDhHAm0MQWZXOWVVpUHvTpMRbVPU
fyTTHgZEMWmR/Xf9hG7zpx8DpU2g48QgQCIPYtGokB1pAnbEEpiHCE9yM43BGNkf
CozpqH0seIQfyqwR5w7zyc8ec+f8hzGS9MQk0PeezCbXjpIBMIc9bs1cpSVR6+th
K2Pu380NJD3vqSw4R8NXIit2im3JzXUDz7gL1mEjVoDZs8Pz05fCdesp77Llhx3V
71j8BYxOV3pxMdibcnFjv7oJqT4CJPilETIzH1DDTpJfNZkeRS6VAS80s6yLKfQv
ONT5uQO5uoYV2z0KAaqEKkPg6V2RbdPoCr1wi4PE2TFbVnqMelJLryrvJ8UoJZpY
FZoZtSa+agtynGi3w6UZNhjI13Rudvahyvsy2PbjQs26Il7jpO4SQcLRR3TWSe/o
Iu+CoKWa0JfpnfpJH5SNURPMInX/n629tpgVfk8BH3qltLHmIeiNgd9cVYa5aYz4
+X3pQe1SQelUrqbqWZUfjqEzbcwM4Gi48NGe3JKI8zhNjbGBdHacmgH1aYGEU7Sk
e3Q7tcMwsIfEwx5Y9RzKer+qZGCA7jQdTQhrh2W2hzAV7pf7sr9QDgGr0Q/TB1OB
gTzAQwNTRsLr/fbvXKCJD+79HSf09ij5rOjbW1bIaPdyFPDy82sLRlHcc9++xAAQ
umjPJyE4reHDIalMBfnwBgHAd22wvTDvTxs1pdzAAPC6XDyB94mdIWGlXAxE7snh
m6msgSsIT3dHYt2psYLpplMFEXu+0qWG4eIr+TSEFEpcEHvSQPstzLLqxPzc1YmS
jwEbwNBYRDz4T/aDasUZsOHMD1gmaj88+uz9zdLkFAs4zISaASkncidI1kHvVWUU
Mb+680t6bUUAyCFKCGX/hHUqzjlfAGpqxf9U7Zqw31uwkyRBdVnpSGnIpUCWoCO2
JiSjpRQP3ATJAbcm1RZAfRTaBSDPoKrc5Ef3i/sSeh0plQlODCT55A6fyQW8jG51
+/xnoD00lR1LL3yK3ChX3ywTfeMEKQ27XkP1M4UvoTry3xzcJyrBt4YyFvBa1Mng
D7lGJN6KSzdch9yMEzAOygFcDYUjknCYjssa5TEAq84lvAHUbyX8jYs+3mXzMPCy
Ot+79i9Kvq5axtodNqhsj061xABxJtTzi2DdU5oFy4WRenq5RM+Edcp7lAQX0afF
pBN1JkHcU0sYqPMcXE/zi7BAp/OwXctPJNf26jcSuMGCP0HrEmiQvng6CktEAWiY
0g/oGJXd9XyHfiHPul52NldfBBhFEITASnZJ2ycsc6FNfof8wGYRZyFLcBU8N6Cl
9E8uITDEwvslzm6/24PUQc8bT7biTPyRfGd0ausMFjgt4qUzT+JAzOkDfX0xL5wf
B65noHSitD0r9jn44hBG/vyTjIvwjJX8sAXsBUD9h8rvTySPXSXo7kbrHzcbqy5G
1WatUeAUhl5UfqugkADahovxug3ndLTydxGHVNgKbi/+gjGnCPxNGdhPr90KuQz2
ikZKSHWxAjmf8eAUIQLCULRuy0e5AUfUuCV0MQtCMgejlXZy1gHXBX/V/t2Pyxc4
hfAbDvXzMAwf8RIc4jtiR573SiUoKAK70avrPLyrHNA0p1eoMZ6bqX3uHYQWD1JG
I0VijuV5VwyUJMtqIig0aC6vYPmXxbQ4WLqGpOQaWRba+Ifqu6fhTVFjGlRj6d7w
W5sVy8CAxikcZGUmGHbQm6ugK0GW0QKKKFEu/SlXGtVHXjGRu3uO9Ws33+JXD9qb
nSAg8aU5cAyEv91NTeK7iwa+8x80lvDuJiZ3UUIeyN0ygkapzuVIna9DQYzdh81d
1tzphEVGgpdoYqsHKtZ36FwBG9jYykgPLNpWbrQimR1Lz60mXoKDrrPVwK6uctvF
b4OqroN1EWQBFNCTlJxXaJR+BKtvnL3ldP0pK5cbruAflh4ApsnHQZFVhc785l46
86OsrfGzI1GwzvSaT+C45AZtHO8KI00AAbJWfLWnvCwcE3vVLurFurYhsI6oJgIT
GUrdA3JixxQqF5FvlFbyIIznMgoZzpIbVk74HtrsbKhtlrS2f0h30PTLSH6zfDsQ
2Aq9z8dKsWppg722Q9QpPxs1a2ZgLjNB2HmvAhV7KTYSPfUwMgTpbZBd7VJmhHlT
V6l8p8uUBNN0KZQg15fbD3O6AkaAX1cUYvfsBm0ZRpBV7c4FA1LDLpO8SHb7rj0W
wUQS/Hf49j/WtriAd1cP9RemZV1Fl5A56GWkgohTFUd2SWbUTiJstccPd2rGatIY
z70J6E/cxwPut9VQ1y/gyR8O6BBdmQ8rrB3xsQfhAN78yKpd7tmmcZ/mhsmcCzJr
8xd4vtyQhX2dgaS1PShcXkxiOnAtSpdiYq6UskrrqwjRu0U4EWBr+EhK1TURz6TK
Ne15xUpgCwGSNBWrANeVhU0TB5jWqGUtNIksl8q7RxDjKv/Y64XVV9Y2fEXSFION
LqiqgVzYDgaN8yq6ISYCqGcUZDPUSpf/pchOkX3D4nfzSp/KxU/0xETm/FMPxcmV
X8BQlN3nEwQ8TGGKlhuKYpqXe7Gb1AGHi2jP5W1TnSLlrwKiYJixmWQmmLcq1frb
nJzgdekdrnOAhAPpd5iXjYLeqjILxzgZxaargoCVd6E6osd5izmWWg7F5O0178vz
ssNJrIb69begmop4T16x1vgFYXF/83q/GVjUHXpx6VxUc+8gXvcXKF8n+YsoCQwF
2yi2qvTUp95DwZZryTX4faV72iMsh6OBlUev5EqVojHcSwKAePJ83fckeD7naOTM
Is+IWeRAJH1yt3vBGRabrT/IoJZUySOPkq2FzmXIKTnAjELc+zcyCMUjvkL5bNuQ
2X2/Nt6hbH7hNjCmVZS4Br4V9HrlmhzCGqcVb0vNvSBCeeuOgx26ebdtQkTgKI03
u9FdriNG7P0gweuGHfgrLVcJXWJrWdfHhDlA+Gx20y6SSEk7dWKqnz0AuJhdoI+N
qCo4goJX6ki3BbY26/14palN9PUv4varnLqCww/woh5UAFhlD9TFs2JK/tYMeoXf
PcnMGCR8RYTn5CN+1tIvB6o0NDpuV/Ke1G0UBASX+AEoDrlsDerX7Fok6Zg/8XTI
01wpD6pmUmZxo5a4r0EY7DTditsPRM5wv16RfiyKlUC9Le6Cx7LsnBDrsSkLn/Cw
Yg1Wm/bkScHocTIuYH2H6JywH0OEf7WqwHfWMm2mYyIem9xr+Bm5d/oznWlU6OoX
yM3JULC0pSIY3O3mNh3M0S651ikEpoInNGFTMZi1WzxNolOZfOwezZ6LEXVzZkyI
Ye/2tLE2O+H/J0NehG17a5kP8awgca9Ly4kw6EmshXk4Y9u7huoqDDKu6dYfiaFc
kBo8jM42ikqnvD3i8fBhJidzsDU+fF9SDirZki5T5x0ROudfdhJCO/fh1vVyc4+z
GGdGXm90sMIQUBJH0j59KWLmmhqzbHhs/SbZU7if4NsB4N5soANCRcdZQ5SvJf+v
ZrPKVEp8W319hGc7B2AouSyodSUKYc1aZIDqgY2UU6C37H+UpK1Kuu/tWOfQMykN
RZElPjyq+WE3a5f9wCPTQNuqHZ0wOFn8V+5Gcg4TdEHgmi6EsLuNxY+byDf0GzQE
SmuciRuUqoTbMnbmOJboW6LjpWoNDPB11Yvs6a19sWW/VxevQrZm6o2Mhqfos6t7
Hxb8MQbgnGg7N4kXzHtk3h36YigalmH9XfoxJNUT2BoQ1RKMPwupl9aa1is8VOqT
6tp3w9yjEkDxtweCMR1q3deUtwMOwE9iAFoHDl91wLjCi0ivRW0P7CExBTd791Cb
fGOQixaIEJzhOkyYlexvtD+k82mmEFMQtHvjaaDVRfzdBJcKGHbcYaly2L27r+e8
eB0abbLgL529DdAk8Vwl5KpWUDFTNkRyB6WTHzUb0bqQTQrrUkcNy9lcMjWTLPvS
wwOaLjCObM6/9q/3MAeMVDxdCegcBsGOrlxeWuovb9rjRCm1fuZQ0n+onzaulS/K
CTGR9ACRZb6856OydsgLpPeO58zcnr7wOng69NCOlux/cc7zjPdrMXrZZqVlTIR0
WMiqXTM0D4/UzEM+rlyCT03qogXqepRUCZdNwHdgGky5hPyTsYX8zY3GF7LpG+fA
hF7Pcp7Kn0G0wWjOdxsp/B8HPOgHsGkHw418HCYpN0eTVlVGH0kvA5Y3eoo3mRAa
jPFQkuDS2EpP70XoEFYx8Uh7ve4U6ql3yVJKulWluEl+oBvk4lThIbcTspeadNg6
1JSSnlPm26Cust7AIYR5LQLwgT6QGUTpIpVbgKPwOYMsE23MxrT4d/YccR46H4ly
YCCstWdlZw+i7grbUTpd6fOfJ2HyXCzEzZ0ElDltRxRvWnNwdVXbj/L0Upo423t9
E4X7erXpf07q89n85u1LLzix86rg9/FFt5qxdh7kdCH+jerKzh6Fxza3yn4/miVP
5zrURzb2241VDWiVqKhpadNn9wByd0EXMC+QgkIrQy+feuuJI2E2mDW0OK2Kd1Dg
hZ1ECUbw8VKwX2Qlep6470SopH8Plmov8MmJ/SUUsPfjT9j4tOyPVVn+5VuJMS6g
3f8WXjBvvfbcG47JQTB8pClOT2wCj3mOeNc86cGKT+MAEqPODfgwOrPtVqndJQ1H
4uuHd0w9vQMQiArUgp2M+ejN2NWF66TDOyQ+VoX9q+c7Os2LwwdabKUM1pbwU78o
g2KUbfUGMe57udJhnGOuGyFUKHhP9kdf/V52z1T3jYEpsQa6kLylkkhXU54p8eR0
3zygQFsmuXArgC3OSnnUI7A9BekqFDKjYpVvsdfD0igDA9OFIXWPnYg8VoquWDiP
1K9aiMHLIynSgrXnscIU4PttyYVXsC+NfAGGePcpYTs3W+WCp8vTgmF1Zru393mR
741KFHRMJUyAZUnmfDSpMUoDpjZu89feQnuyO5Q8l3q2FFUA6TFWVTAtHd0bq9n0
7wUU+WFheKI7wsti3IzYGMjnyo9sxxfdsmWPx1jp4z7E272Z6CP+4eji9u5nvoJA
tate95tC8R5GpJiOWbRf4T2vq72l+0KrHIllUat70gJqZywa0vhQqSHs6skL3D6V
7wR52FtW35ZIDQuI2dg8Wb/CRXH1IV2ywWMY5SvtTaCmg95QUwbxtT0s8eaG2p7q
wzXC9b7wOHYWJI8niy6xLqw5jHE2PdaH8iScBGhD98GTvjFKMynYwPSzYVMhzOUg
MrcrpUFD7qovuPe/veaCKfSLrFgmyMXkP7AFgGFDng1jblmKGLXDa3l/QUoKnaKV
HQ+e4p5WX5ENQTHvUffz26DyNZ7tB4UcXQGW8fLr3QaW4/wI+8mPp/LvEoQhviy0
XepE8hHfI90jjpfhpVeLLlIBAcuaCZHWnvPUC9GQapi53kIghjMiztni9ynsHm1B
odpL0y7Ji8MREhJjCPx7VF+uabMIom7dQ9DEXf9rz/p9xbAXa8tBLjNtrRnIYg4n
DsFkX3kf3xQR4g7UcYr9F+DhsxeTZIfo9ix6NEfpPWoNAffE67NQEt6toI0hY1u+
jOhhTdTKLNM31bRnX1kOIYQvsdLEEp467yl+jHo3NEbnVxPHUyHjvUGJLnI10RbD
3+MARu8zEea8qpZuqCRUuGB2EabZ+djrv5AMonZBl7Gfene/AGqyrFjzaQCFvhvK
AWqw+Dq3AM2dS65PWOy7sINYX2DzWyaGFYmwN1SXV7etUNfGqqDNuegrMhj0XA0t
OTg7XsaRvfUnDxtU4lPaBBrQWY4cCvLZHHt8GB9/5fdnGcGSXZkOteXifBEV2xOp
/QL8pg9UeoCtRCI9WuHDNzWo62X5ZeQUFJsOUCw7MKcqhvPRw3e3wnIBnQN288Jl
wfh07AZaCah/JdKaB/7r/HvsktAbBP8EqRhbpglqI+5Smc8qMTrdwCvwHDJTDj1q
Oi2EcDJZ3gLbsmqNp/ikhhaZnWgLP+vrbI4PbtlghDE70u7QIpDz/ucLoynAqcjb
Kup4+3WNuQk5s1ntprFFSK5UGtSPTC9SRyoLd5mFyi9jZG3trsFqNdGNBdAchF9g
mngu2AVdl4YXS/ObTFsjzCz8voL2kKDtC8TxF4E/BTN5bM3oEBcfZXonVqyf99Ty
O2+EJF2PX3UcUltJ52G3YD3K5A43ZOnRSDLitNIH8ys361EFOhxSr/ThQv3DyJkt
+LBPS54cHSbVX1Qryjp84m86lYE9iKPaLHIyUZ/ccA4fFKvtcJA59X/aQY2SnHpW
KQcn1tHPjbR0qFRYPO/IDHkz/wdGMlmyp/cM9HYY+c80FlKPQzEJg1rMqwLa4pKw
QUv1zuZEJewicRgCDTEomM0fkVipDimzHlBaVU7ULBq9uuOY25VaY3stod2D/aad
va5r1z5rUvYO8Ns8Z1PN0W6FFme8mbX+DoJe0bBL18vlHzLakRPZAboODW8S2fiR
edK1LougxriYGPBdGScetx13spQUxjomUctKqNKSzCXpExRPDWoSO1bjiJqv5Nxw
NMorIBeGFcRsrVcB3ey0+hJaubcbQfHHfTsaCmjmg/Gelg3fIZnvpAD322RgEmzD
l+fNDTVIPyD3iv4nStYK3AQAx3/hnYCzcmXjRCU4O0hlKe/qli1KjQRK1OvSOJFe
qtJ3WqnzrM39dofWB48Ytks62r/evGeDXk9jQuNfuIP5W+GKjKLCdNJXAgl5GQER
Xge4Dlz7U3nuO2srxyL05ki9aY+dW4PFhiWkTg6TGvfEj8ajkqEecnbmq5ZtIFRB
FJk2r0PNu3hYPRfonVn+XwyvOapa2FGRcn7kCSMM3yfCAj7wajPqwMH12hOy6kN2
cdT846ZTPax91SHbVKDDB34MJPos3I2Nn90/eoGWYG0JUnnPcDoEHshgoVbVUSNg
vPQ2OBIVbW+BBE30wEJCitBaYedJCVNRQUzXXq5x9TSe/+R3QH0EWdZi98oIkt4k
0z3xhkvqFw3ounqKWACvBUO9KIfjlcfMtDREYLlW5FpQZYSDiAQcM9jGdYQCYMD4
APVR6qKH1uDzGCwzG/nU1lLqmZ5944bngH1mMFhHFZ6HBh4QxEc52PyMS+mqp+zX
7P/JhYNeii2aeUABDWDy2kVeyte1YtjSl/WEAvBhNsameqiL4pSny3hggUJHLo4a
O0zvYvYEFpLIbamI6+QDgkpvasoNRH3+JY+RFb5VCvPRx2TjK7eyW+iRa3cmNBk/
8wnB2CPGAcQzosYd2K2vy6n884YTvLquEW6CZ/d5uLKkf+5pATTnpnpuq/L5PkGK
Nl5y8nHSvVKqR6VpgEpLlt4yOtCzvMx424xkjosACOoqC9PTh0fJdxgSj4QOIiwF
5nRRCvx5YLaobzL4gscuwmhKg6AHNSYhJkh52I7r9wvUmJN6KmwI7lbHelqLutOI
NhDcpWGDV+EPaQvWD52UkX2par/2Ikjmeb9prGabQtNjEZDk0vZIjDvSawMzI5Ft
VRcPfihm2aMwUqMdVm8vqNhyIvAZKhJRB1ag1YxLYobFWC/1hKq0Qn3UaFmqicoC
uS9v6VK4Ika/ErLGk+7A7cX+fKtqvLYv4igQre4q/8ofpwa0sWy9Noh65QBNVX5S
16DT2E8NsptIxlzh8TBBTC8Y/wKxswtcDNj7n3h1T71vAzuN/um3we0IjuvSuQqT
B8N6rbHj8nzKWIVmiFuPvH2lqqrv+6Q97i0xD6YUwAS9DFIBJ76oTE4+k9Bnwv+v
LIfAvML1Gi6CX0jC2PXHOO7hgWk/bZAobqKoh16sCI3RJM4NxLtqZETFfYXmaC3f
cPkOK0v1Av4gduNMVPkaMz9uqYpH+Zp81OKdjjFxvIBk2Y07O1Er9fIc3Y0AzbJm
bdUYtYuvTdatkKLX9t8WHwa+dU24jP6BGEf3srvKkGPF2RwqT+zBRhFWC8pU7obp
UnhfdCtH5OPSZTOIuMYt5qfKHbFzeP5gduHxECPYsZGsTBQEDHPwew6V3TkCQYP2
JJccEMJNcpDCWsfVG+wntpEIwcsxjbaULiN3rfsjwjbFgZ1KfKjHyghkOGIHOpxa
aNRGp6hEscPtNJp2zpNpulnLxkQEouX1yrVmZ4G31IEn2pSFbBB3wbbZ5hh+H76Q
/XM2qx/NDL/2vJeU+RRnrkHBDze8R7Bre1HnUNcsh+mQxdnys+TLK6hu3pCE5ZEy
CnQcttpm8hALpfvJARXXPbCvSRtLA00UTB4ubAnzgjz3QDJm1GffYinUXt09VXoO
kSwsZ4d9FlUnCTa3s6qQR9yBxQLopOPeZP6HJ0agztflvnz6chN/naIOvkVvHbWn
FHLhcopkhCqfRwAvKnIZH30G5kIrEEYtF+Fkcumyl2hbCid/6AmdEDuQOEGBDUk4
CwmGhRT38meQRd2pRl8/YW5X5Q/p++M5QTczkHowdWLmhk6Ju7+eRZzKhPfhKkeC
z9MZY1oLVepEfgcA8+dEe2Ob5uqlxcVizqQjYH3llVb+y6hPn0Xb90WVudeyqfeY
2MtxuvenHFaTxHK97e/OaWWIbh+6cv5OKKRmMPzceUK8PBJAEGE69kcJ/CbtLj/H
n/pcB/+iRD2IkDrUzhC0pthMXzFzcmtbRx5D3kPm5NCxtnzEJM38GZGNse/Z7QO8
qTePOGS0HV0STArR9YfAcBzGV7A9FDmpI/3wgLZJr0XIijCuRswXrkiAqw8sRPvg
86CoOg/mlCHyFzfWho6oJ9TQrM8llo3HdRAcbIZ9N/FPS98FxAi/MvHL/Wrk+WEa
UJiVP3C35un+Z6/XrRhEQ+ozkjzqg+Vm+2e3B0JDswIMbBeHU8mzNBtkEb/gF3k/
HQ18rmOHPlyVwCsnGEmufQfFbmga7xYsgd6J1BaTK6TYaQaZtIuBdTpteUP8yv+O
YwfeDrGzVCv3APZkO6a4vwk8f9eUNLlYuqsY4rg1Hqk48JzoPXrzlSo9Bo28Qm1a
nzeEnTfM6G03BJ7aoRCABjX96dVPGm2a8uL46KD98YDK/yJfH2RweNT9JX9DDcyC
ngJWgB5wiyDIkXrFZ0fWysmhrm5xxvt2VBsfw7kCB19WkPnRr6UOvbyBD80CNZzq
aSaBg0jCGIrM4Xir8bkCtdNNCDeZ2HqSllrZgZA1Ui8l6ScEgNt1EBhps8KtRIqo
x6KfxrIGC0t2ml7ODkDc04Kpsi+NrBi93yAQoApatNQdeLP5g5bYnXBQ9WLW46fm
GSB92Z+T0IEIHI/bekOB/z0Nmm93oEpHkTeB35z9XCJcPEI26wp1kv+JWnAHpFbl
zMkLxQruWd1Jys9YHiIXt8P4pNllueIoKLUn+JD4NolIK85KfUyzCZ0tKg0qSe7v
LxoEdz2OALWh4jam4KCo8Sk1mjXqH9ay7Hgy2ugM/enkZea2NDlBir1S5oOB30Os
sXzvoeXZ4Foh4UpcegdlUfDcp4LypaCJcFi5QdjdfDRG1RHc36JnaeksjRn55Y1M
X6cQghq5zbNzaU8ocEj28TAXc7zx8eSY5D+Hb0YdyifSWIHkgcU09THr4459OYoU
5GObH1jds14LRJcNiWaNsaYC4rB3uzk2o37SPlRaWiXJyAcMYo9a/v0B9wLszvY+
IU1BDCoi960PpREzNgruoBYCSaJeNlGyziSxdD26JOZfain1uHCVbP7IEaqFDrX5
m88G375ripKwYfNGwLFQqxUfVl3g51xqEg8gzWPQhvfp9IBSqRxst8tjh2NvhErE
PwjLTg66roBz2cXvD1CtQGXXo0b1gJSeZYyET/gZHJysc3u0cWqHlZ0E7JxkgBfY
u9U9wypY85hb1j2gAzFOfOtVRLTY6dIYGQ8gFP3++mlQebT2HzC/umCmYcnf8+/n
4IKunHPdSSHKhW+jAwVOhgxNPryR0T3EOeRqaKMRNKL/CaDWfeN36O5mW/9q/qP6
gnTwtqPXq+BXzSLdKX0Mv6HmXHRefqvn9+Dx2zGsdFObK9Pxq9xj2pH0VryhmKA4
1iUs3u4Zfj1CISSL7h8097VVXG/Hkag31sj812bt4nNlpjmg7hz4d6u8D2ephIFT
MxfH7U6uoTg6ux1GP9aMyzfTJ84FntGXp2iuBPbBPsA3b4v+LfvFBBHGovNfvNq1
AqyTK7ItNVV7g6G9ZpEa/tM6I1AozUp19pgfXEVw+jM6Jhmi2KAmMyJUtNwowYxz
Z64k3k2RQ+S3TUU5/PCAQjzZyeq/3kIuVZZL0flNNlchOYBoDGctQIlvQ91m+fnu
8zYB8xK5SYxbeGmWKipMEGcWr88r5uIoyIoDL7Ao8gUgyIXw2TvttOH/vXFd8ZIp
4c81cSkT6Nq5rWCmTJu6XgqDtQQhKIvO4gUpsY6uR8s4Em9h0qJ4yuIKk8azxIN/
EA/YghEr1NSGp4znOKAD8E1hmm2BDh70YCX7yrRwEGI/DlB0rZUShptW4t7hIL8V
ug8CdvdH8vhw4RPy/CnPBeCWVENRJjUMGNdzrfR/AcNiZVwEIWR2cubJQJ1WAQoA
ER/bniS56UJqAcbDGX4+Eq4+UWS8hfFSANwybB3inSGmsERHC/zTCQj5xI/JfYwv
4JFESDUxTZv65xw2yRicXSO59PP/SMezZWXhF/2dlryNs4lUrx5yP76ggRf4nyD5
lsXb7oQy3gjmcBYxlVFN71GDJJGigQTn4l5W5zI5AXx+pgAuoUKlhrs/SOC8UO/l
0d2gKMKjwyypDUOJlMlJylMr33T8Vkpi6nvA1fN8cvVbHNOHJGnBLzRr61ToEihp
1n1fWgzORtbVx5Byesarsu8Yeb3YtbkSd51Z0RTug8Wfij0ODY5unDCsQFx1W5lX
8StFImZX6DqMn87HCyOl4V7afwPsXda+nx5SRVZqMvr/JN4FNPgF9fBZY+Z1bZMI
opX3m/l23l/6JhlwijiEDtwh7xVx3rTkMhzYC9o4FdXcsxx/+WIaarAddxlypKoJ
KMVmjFhOQQfNXMnBjh5DERBp4ijAeurGaNOztAB+AIwAdII+LEiFP/hUM9Wd9S09
orrXVHngEnQFlf1fW1qaUQlkG0wmlh4QAzaLjdGVoE8EQP/Yg+Qfpi0TyWS6UAqB
MEpHHsITbsUXYuE11WVBpCltaK9B93g9ITRlA7b4uD9xTPlqYT52+/ufDHIgRLfv
cf2L5v08cuD6hotV9wTFbqTrstZTlf/BFYXL10EeMJFRFA8KGqbwl7WBcYpnMLFc
E2YFfs6viEKQhF0SE+t/4Ywe/JKTcQCY7nALFzBTF1O4axoOPXBwtXjmzI1rZUfs
cXI0FjMGS/vcUfW3p/aDovi040tUfbqj+DUK3zH1M/mu03hIPJWkMSkjziVDIZmd
yiBPEKr+Dvfygh5BU5KrmJ6XFQ4Hfyyvs/KXUEGDYpvUjzynejZQIfhh7hyqa4CK
9du5Jhriy2ehdR3W/2bMJuU2wX0vnr/UryYdQ9+FMSqZbKzulAeFjXgrQy2SwLhz
+wryGzXkcadbMPTZqYAfb6PQQTaSGwCdw+Rf+8I1W3watjvxfP2lMLZCidYXVpg4
r782rmWowDlqp0SdomCnzJNvz2q3F6Jfhu8btkY1iUtsCJy/zfLfBl8pHNH53Wj7
ETfvb8H8oEFXavHz6wI+BN7/RCBtePpFWfZRB0AKX/a7uiNvYKU0pOCP+sjHOEgx
D5keLdSJjvtT0p+LdqhIEOAgBp6LxafYKPDZSTDCjfJ2Xp0809iLx6uC/PzgvgPY
7zjb9P6WC2dVy5yRlRQ8sxD01yxaLzwPXMXxQui5Wef8JdoLF9ijjvHDLApT2NoD
JBusCEVEfL44zZh+sBojy6XGbqtcol814F6gdLvMJP/c+FW5/gu7TolHbp+MT+SE
t+1jeW3yOK+Dwvf2I//ANmEJQiBTYpiT0t4matDj5tWXs8rf7Q8QQsOYxYbU8l9Z
J3Q3b9r0a6FBf+6DpeiAGv0EEbvftjjOa0aGrDUWzUjLb/9j5iYLkFjZWRF7DTmn
wSH8XwYcNNFzaD2DxHvog/La1hjFI1yw9ZjJQe1wjd/EHCCON9MbqMT1qHW9Vgwl
ZLO1XaSQgfL852xx4xMEfQ6Seb3Rcdu0Zo0udYdfHX+GdL46GWSO68U1Iv/zMbFO
r0CgINY9k8dT83GHWL6S3DllU9UTr62CZVFHsbTP27RqBj8GIPlGNJSHgBiHPb0D
hVv4FGgipBrHs31lhqQkJro3bQkd7plpSgqEA4HurUZO0LKNfyxxw6lVacIN9KhK
ziRzjD3yOIDBFHSRS8SFF75Jt2Hp+rFZh5BR4w4sGvHOxrJww3UNmLFmnhj4oSdA
nyi28cAns+xl5PKZ2j5MYQT3Et0/370EvmD6PRo0s0S0Hvfs3n7VJxsItpDvLxRL
PMrtJY5bx4SXjQ1XTyh0y7GWicgcFnbAWYGA/oqrFOAmPJt7T5P9BIvXCmAbnaMp
ABvYEnUM82f2fdGlXdKgfNcOZSjhbpX9zbIhBCA0lvdtEENGlORmF+0Xg1dUg7Sv
FWSfa9oznZM1NWhsecPWJRzMQtqmXFIlDU/3CUHwDyYvPCLiY/kNuLpH5pRPQVHL
r0oMznbaYpcj9tUF6dzT9q1TRe8xy/S7g7xMzw3tdP15lGHep8XluT08ad7EeeMO
GDldQiCxAdzMuTk+GGBufKTa6SNnt6LSHvy+8yVnAT2JzoVqTVDwdxmB5VcnjUEU
lYTZVV6CHzwVPDpQcA57or7EZDvp/HhFJOy1uf23NNa1xHipItT8+gcGgTXL6ZoT
xrvOQjBDPUUD41OLpIitjy69t0D6+ZPaWPR/ZwP5ii1kublmuQSt3M8p71d6RwGs
u4l9FNuo7kv9bfOGILfJfirxr31FJLEl3vYVoyQePowGeq8DRc//jzMXxRI/LiJe
NU+a8QxCS6i5zld1/W828u7xJXNktjegjTJF5rluhQl0r8suxBXqj74mAFaQSLeP
5pLXfqVUd7dzKCTBP3wfEOHL/21BQnP/QSo076QeYNTbg8oDYrt72U9QFZOIMsfn
kH2VNpDuF4boxCw0BU/vnkKp/wYXc66J2ulSdXqa/+yipiTB42jXnJROVyUm0Q+r
LQUGQgjMLdJQdtfVMPPll3zdCC3/o0MD2tH8GN/E5YAzpWfhRJfpCq6yjxh/i9hI
UAUdv+yCIqdeRDPDzwRXqpnqG0awpz6/QyR3JywjZ1oSCtoSQqNfzI5axViQygWi
NGlvZcPAgKHXdtcuFzNbgIlaBZygKlTC5Awi3/YUvHv4wTIDnmsNIZhjcviVqsU3
DerfqHcjIIEDuHuvMsgpbGn1ULub+ZRKZO8p4pTvlv7YVWiQKG7FjMwg3qMtuUuH
17dHRuvYxBi+9gtYsIO5dvS00/b5XM12kEdT9jXW3TeSOhwKl1R7UAyORoGLGMDb
KZIvXVlYuAaYb78N9l6WwUR0es4LtTomF1wZ6w9KrgXrVl2N9QEDlz8q9v4F4/O5
dHsHyMYcK9rF5oCb07o/xNRDtmD6xJKL/E4dfpRbTY/7cLV/3jbuo8CJknTFSUsH
TOXNTuG1KWgGuC57BQhdoszPy/BLBRnPRrwHe+FVrRf9R+crzDtuc/qfCzdpY0i+
UO42epSKTOWUuTuLC0f3AwFzl8PlD+hLz2w1+H4sQCd2L/ZHi1pWeO5E3A4IfMko
ca7PhaQZI/VM/RublYjbtJoWW9XQeZ2bPevC89i7LXvksCoi7BQQZT/7oIq4grqP
coBZOLSheZwppp5Yktob8VmpDqbEGWMWaY2dKzW6vLOtuaY2T+KtPB6OFxgYWnye
x5swuX05wFW4JZp3WORYQpHoRkm89WnMtRXLdcZPdotRd7+ke/zv/2xiZYzNS0ym
bACaLaWTSOAAQszXAhcppGkAJg82VtXCelfvEUDDScAN/o1H1lGbyx64VhCv+UZL
lGBtQUV6M6JuRqof1BRkxnMq2DJuDNUpPgV07McCw3elXmFzd7Ef9SVg/KwVJHnM
WaAw6/UTMErur8V7kXE89EB3yve0ah78P4qM8tTr/vbRHn+b153pxLSvjN5+Oeqn
smU+otVobG2LrsGtJros6zdP2EYecPIJqVQozRreM8w9ikJqXdSIJcHa5rQwq/sc
f5zL6Q3cObnZzCaeCb2pcwENVpZ2TJrHXXPtRi35Znw1SQkM+mc8vDw7fGsVNaSX
U8fNNX3ZFAJXmdx95tzNRwEvxkS4OFlHvrWIRK2hXMrEtP9xBLU49i95USUbR8Q7
uRhFo081oCx5i46dYLHN8FgPArIuJk+HIkY8nbX55q/AXUQZqgw2VVcao7fMnoFv
zbi9E0BiZ38hgtDsdbAz4h+N6uGVYjJhlTp4zgilep31cn40OTVHHhrnyvpPMDpi
z/yJizThj2LdoOD3bkBIirqCD10lJwlp3YiR8xJr5bb6rdr83BvPErQvD+gjpENZ
bHCuTbg35C6IHwDauNa9Etf1nZIuMgLWn7hkN5kw9psM0CbpG2LRpKC7A0gHyErR
79Mif14V4jIXuO/86WyBf199E5LpiP6rLstFKxMd5DeEjKdhzN4301gQfdpIneZx
O/0lyJLnz9ITyZsJQuJ5M613McIsKc4Hn0CnqXCEuID0ygOR7pa28Lukr7zaE211
ISchgrpJxrEYqMkmZglKpgDNZhUzLK9NeDUsasWJ14+8NEil4YUZ13IKRflUBKP0
USaexJ+2wTxa11Los5EE4N5OZj1o2i+srrcvd0VtW4qABhSMCYCayLNP+SYO01f7
or1dQEJZ2O8IcY8RactA0i/65lEq4cWr8nznEXagiSCpBpXftWXtVAO4ZGxl0Ipp
QKD46VZd0YvCZpO3G4jJtCuvCNQDmCihnIEaWBghUfKq5kTB4jZ45t1jkVYneBLn
Nfmy9ED+BIN4Fb8NIlzXS4pP/RX1cDByvBtVhqE+apGxUVMkQ1bm5VFMkthTOVbF
7jyCOChjqevX7fLB7Ow2w/MBCJcBzWNY3lrrZD4Xrsg966gOFqTRs8xgH9AKa8hj
dnUhrjYRBPK3l/C3agASOYyrZmsh25uZTkpzA+72hBOnFe0ghx1XCNgsYjYVEZKT
bhgUSQFRkd/jPvaI8BRKPv3BqIzrFyM0LYoqVR/1UToERsUc/3e6zZNIehDs2vz5
vZqYNsPOOTD6JTTaX42I/3lxJFNj/LeU5ijS20EJbNlYc9mQ8NH/f2eVXmzpAm1K
jrkRUVWknWvpuZgKzZU+yFARcjr7DHMGM6KFzqcDYLGb2NGhhUj8o0rsW8VHKwQ6
DNjJbPD/1lVm60JPMgRNXOAi+tl2ErLPMW5he87FsRfqhPxOpq4abYs4Aq6a24fc
8a7lQx9flmo2A01XIPVJFGIBtGQJKtm47hqvj3JS7c3XtgFk7k82q1ePpIxHStdg
qMUAFkCLznZ8uv/ZCTaea1xLbtaNT1h/zyUe+8QHRsoLd25aFRgv3QMpW0zMMuGE
rNWftE12GUuoo0WctfQ4Z9sxozUu1cs3z7Ck4efvHFQB6lX9KGYhwJ9ttpADYWsK
ERMN/42WPaaSNRmfszsl8Y2XePDCadjZA3hpkfpuFiRpkTzY8t0JlDYg1gGmde3G
6NLn0cSE9/5AT3y0AQYgowjdKJPlGelBkmM9Ng5IJkW6xlK3bTdyrQU177sV+196
4XY8EfRwfdX67yokYaigV4CMRIGroGq95cq2/UanAE9lCPcVJdjOTg2sviMG4gQw
CtWGJDTFGqG1/lnGy5WlwnLOfrhpI0d2cRZqjdnP/SKA/QlJnepmWdb7pHd9YZfw
d7jg1OvHNhRdWVE4EHLzISIdNFpZhLoZEWdLJm4xYVFVR7MiDK1KLAsqlut5AbaU
HMo7DbmaugvVgQIj8g/vmQQfukYcDdmW1S/dZwt/n6R33ZHAiGPQMPX3UjOPkvBV
fm9hxsr66wypc+OAsrMcMeIxe15eYlYwWrzKyOtVbWY9ht+sO3TRjJXikugtMMAG
32CyvPSaVTFAASWsAa47/66YGzozR3CNJ9VH6Yd9VhlExq1vDrXuYufe9HnYpMOe
UEgqZVxEbxh6irF6414vRCHgALeZ1xzDzB0uZ+oFZdUh/bBeFAxXXhePFV2bJ8sd
10R2riHdDXJUz2z83Mem8rLUjQ855rBm6dyPgg3Qe3gcUDWSwXy3s+8b5m+dw4p8
HGrHGxFEXr7dEO4iQRrI7R4dHnF8sIu7ox8bGCQMPHBtiAgTvtzJEZ6yEs7fCUdk
65p2yC1FVsGrgOrviPPTUq9dC+CQfKRjDScRQpechIJb2dwYJgncm+x1+YoDYXu5
oX0e/Xu5qiMNlVCQ1uRNm398mBCCiXN2ByejJonzBTbAeLMNZpgtDNwEu0Fdwbmz
Co9MtiSAivAynuXZkaQ8fjaLKnSoUoEW38Fcll52j54VoyMllrXWa/apy2YGdG9I
nnEBBtUSEegeMcq+VKH27O8Ie3PGvodmVuZ5P9C6Cx56KxeFnQP3qzyD0oU25mzv
ryjtmDpy9MlsS2JWV6hiwWB0TGIy3Jmeqwvot0ILtr0O3BPZjiZsrnZjCVUiQ8Fx
U1/WcrJwZIobwGD5TLlMOymvwfFbMZduAHG4tgAJ8Gdqx0z0gzGFE+3zi5jIZcoj
TDaMwA6ormJNEI5Nph7SP/I53wlOb+vKLWOwv73CNVj7FInqpx7zfqbAsLuJXngv
f8/D2J7VFAxWBWSEIPDpQUnqgeS1eHEdm7MkyPR81z1/igLx/8w9AA9gzWP8c4QB
DmMAQskPAXGvvrcrV5CenQuGWB/gfcZl40FDOYpL2YW3fPud3WOYicgACx29lAgD
9uXy5DRWDhvXEF0/w5xed/M0+RlO+Mr7N0rNvbf0ugqhJxlf/kXP/TB9AQ7L+dJY
KNtMQblO0uF+JyiDk63OrEfb85xjIE8L5b5/1MD8SSWbcIX9+E194m88odKfdGfW
aom8iHYoWm99/ONpJTOCOlBvUCX6vYKTrXEEQU8DIFbbRU2WWJIsKHwlA428KQ+4
PtQvCk+vREJ1YP+fiu7aNW3xUCOrvbiHPPCVVHwTH7P50lYKb1ZCaf+G36M+f1D7
iZpQDieZcNgIpaM7kW0c/sWCxtppYoT/NTWRs4giBh6Q2Qf9RYSHS18H2LpOjV0X
6F+dth0qEosdHwUjWVQRMYMCeOu/sl5hqPBOJza3bF2U3aUnYu0wi9qUbbku3+vE
eQ6QLE8UEWk1rhNe0iPhSztEUgbat3VOgsWEyfWEPRKGveGlH4LpDFQmypfm94z+
KjqGsVKQOcEpzKvMd3mzPAQE72SLxTyC0L/Ny2YaeI/au+fCb+XJeFdbBtP+nqyH
GO1W+03s1yhSrXrAMFkEG0d9Dc04/Z2hwBwxjYjPEe4XDs1tMdXmtauNtxFOgxh8
aCxGyMGA62SYoNUhERlPNMVmY0wDH8pwk+cCx29AFNXFGx+kHvAClW1DubX/OOFJ
Sr2ovlRN/QSrhfTsDKsJPTWPPP/HvC5fL5s2wXEIv7cHN4DZX4mh0emsJX7D4R84
q+/Y+vbZ07MgikJfcIM8kaGgN2Q7j2T9GXTPnzFTcmTUrmvhUgeluSQtash+sLk+
TsG+xgmmAuY92RF3lCEGxmXBRiL1K05GSlUPwYlapRPzt+3J/iTa4+J4xpAwMnO1
1mE4OsD/9X5gioQzYNzwXlRg+mEtxPf9/M/5M7yQDrLRIsCTyzEy2RzNSMeWk/Hj
5Jh9fhxO5huYGWEb22WDFXsE7Gcdso3rCqges1+BmrsTj6J2/F5bUS5WjKxre6xT
+BTC74WMW+k/06u1IQl+zuQzEc3vo8ufyY3TVYy5n6/0EztpOIHvaunavxiixzJz
uPzov3TuO+uZGdWwqA0s71gnckE2knizB64h5aAUc+r6Ma8CGKc/szHXGOV7Sl94
OcOpr26tXAZZp9h8vusVegx7J/UP5oEdAR7mm55CvAm0qVYyZQp5xkLGZZ3ebyEn
V/C0SUM/J6juHjKrmDIyBxWc+SKvW57Vl18safzaEBAFTJkab+Lv5sGeX4SJ6nIp
DuTH3vxO+u3skByQiTiRehuW8ecToOz6JsXq0qcHEo1V2bBKbqUVa+hMoLRQPwik
/nUFgMR7YUHp4adA8KZNZfVsVu0ArxiMPwO4Hs3MRvd3lbhz4zlC50wI3G0PhW6S
skIuRxPRjrgW6fMjo02afyh7bl4bjKo81UIYhRbtZGRe6a+PWURH6kcxC7PJ/4So
eygzlEREKzWeP04GdVhaULXWBvmcylwQ7kTjszGg2oU/vMzRFnSgBUotKaIRZsL9
/vn1jchS3NnuV0IrkJgo/kUX7RGUoaV658G66v/NGmd0x9n+LNf5R/pDxH8yVKgs
kImWmt92kho0f8x6MPvm9G8a6+12IwR3q59nN7+BGbKNoPnXzDankVx4rYxPhK4T
9iZYb6P3MPTd7GsObf4XH/t8VaFYkzekx/wJ6WbSNWvTc9uX9Hi3Wt2WPvR7eizO
GxolIC5X7o7yeGQVAL3EnhpR3UWp5cgCP7guCg/qpASO4XSSkk7mPceIwiQPPaAX
JrKnPoGwm9D9aHpEvCkVlX8Sybhnt1mN2ZOhRLjb2ij+Jy8aVZ56nXAcm29NcOnl
kQ3dcEJ45PeUREZG0bWGRmG+nCQtPySmY7NSwU67M7IVOTIOm3sCu7ne4Ch+9oRB
d1v+Fl+6+nb0DC0gRneYm6orG6NdiKGrmBcB4gDGVuwcl1w9zOj+AtsXjia1f5gN
1qGou+eHSj2PwyoqYwjdyJ2BdgzQIAb1EgRj+2iDkRT2G/0xIHa42iyKt25r9jov
D94g5Mvs+Pi252MqmDei6tA69+ufuuuR0OY8sdZu51MuajB6D3aZuqiYCYylMegc
PwZkrg9p/BzoQBMNssSjcrWb6pdUgeeAkTDvh2l4uqX42lipuLwgALxcg1Ir0edG
FAazvFxkyL+kaFmOt6KWP4jo7Yo8N6VQcI/9DBm6/06WQlKpakBeSB0VWDqLNqN1
CejNDt6aavKjwIfz9fPATbiFy6cnP+7Or2fg/143Fkzv3EyAPFkUvVnls7GbisVK
7+OhIcIL085+yZlKSi+yEzPBzVqQVjdP/cgNsUVPkuxxosEKuoSLIJsWR3lkUKLN
ZskOSEI28dyPfxHVTCEshaH37vI/CrcPxFpfhKLNxo8PPDKG/bdLHLsBqfxpaHVs
5dzUamgD8/ykNOTxquKiIzfhlNgGgVOjRd/d1LoifGujuo/BAkB6qNTORGSH/qgI
h9fPwV4OubGQNqZx2rGWCl2jLT+i8sAUZGbdKkzJDkY2FUMWkx608LL2+EvQqNUJ
CgjG5CVqwWMDGrlj26SggXLNOxZ0+fPmarDFaH2PC9tGjKjYBZFu/lML9RXXbcy0
r0OSCxsQbn9FbTZJ+QtFG9F5MJJTeBMJBIAcy+4PuuR9qtOxbrZxADVOECsjsDSk
8qEv781aITlb4yoIsM+vASG/TiafPNqUnDhpN5Ufh+DA3lLFVqwEdkLlnKtSSicN
rcsN1/voQprjm+1DgZDco3sYoYyGWoKeMA2ZZIY7f+K7Jxx1h2mz3Ct3Nn08zgOD
CHD7ZwBHY7i6HzIzjyjCZQqMYTFeGOzBHOTnMCFAn9G8CL9En6duIAAvDGDs8xwv
v31T0Pmt/zn8O9zy6XM70x+DGTN0VWJO8PSx4DzWODX09FfrAhygCDeFHW2jjQdx
RRoFsvoLq/DXmj/wEi2Ur+ErDXpM8BLn0YHOBC/FcGRRBzgK1oRhNiQrr7t5jzGf
VLlQGRIzjUdmGxTZwJveWGp2lRDKKV8hZKf6+ZLoS8/09dX0BmyJexM62wJE5Eq7
2HSeT47wus3Kiu3uexW+Kq4miCWwn1UlfbhSzLqJyQ177rXu0/JROzYvzFOVPkby
P1z/pqXzuSx9ZPh6VqYiZ67mebJox/r5V28t5VzReGl5OL8UHxph13wNY3xy5Xor
aAUkM7UnQeS8u2zBCFFF1qqQZEsha+nOARSsGe8p+zrOnChPxsrw4yzAkSfII/lQ
vYU8/TNQwzMRDrxHRwll8IObt5QKxPZdrXHyEux9HZqrf7bRYeONLUN4ke3kwL6E
lRqiayukUQYhNPCk0kAbey7ibb9wOjUFswc9nRSMdJILD9PUQEpGvxRT+Psfxi+U
ipIa8Kg4GhaGGZfM/MElWYZD7U0nfp2dKi0sIiDvxrpkrDxYDQEGNLHBxF0I+/NY
6TFXGIF5asToDwWDs2Cl9D6E8Kncm+ESxU7RRLCOgjjwz7s4BmysB4QlzK9Wu2/t
e7Q3QaiYY0qY1FA6po36s7I7bnGZiTfhj5hIKmP2HdqxwcsBQbIpQOSptJFVv1Fb
+C0cnbPwDRsWY3GHdDp/EIpDCt0ZyRp91AEWv1/GB4EFdIM1YgP+mTVgSJHKaxx2
8mLhqLo80kmwUR1r5M/5MMTSjEnzhGpCpRpxaR9xcv13GfnhSlfmQmFTO45v8eZ5
CLCFrMY+JO2ndUJMtmA1bQyAacLaBCA21Hv6LkH3vJe81I0bM1WlWtGi2u0g8yRe
P6G4uOfCOj5ad4NG/WQLDqUZps5w7fu2Y9AncYz1DBEgkfeqLEV5PtNS1sHJwSg6
dTX9uhegvRopK8YWK1eNxOubc/9rWmP+22Olu7maVmUOXsx9QEFo3NcFEfr48wN2
OgnSUZh9vDUdHvGgaiOz/NIjCAegfkIjFFcm60nbho14M8BoBAp6WkT8aI33xO7M
RTTEeh6JGVO1HmZgzYFJfPhbpqTjYUYHPzdCcdFck2+TTIKHNGqIzHFjJ60YKFs+
SSWG53Wg5mIwkNvZ6s3ISLSeYUPU5TTzcFecGxyPG/QmzzyfnttBEyzuvxUoLZ47
2/+3NC8vBXddU1W9GOrXfJBu6hg3dOjBHpuGjLZ3w59Dajs/pV6XNizYJYSvvFFP
J5lf1P8wQtE5swHj21oRM3Bcb9/fRpjmvN5MaOKkpuDkI+igupVjvRfAkoS2MeQ9
Qsukpx/Ah/jhDjXWggnu8ALOlmiBF/iEeoTYbVXvBN5zUQWO/OJPJTPbufvtZVXi
TArYbeJdugz9yviJxFtzd42gqfK7R5mO8JfWK0eO+xxMN+1LAumwY5wMSt4P8xgn
ldAMoDyLZWEr4niE4regGWlTjmgSGBiJBRGNguyrwoQkV9zazc8sbht8xKZQ2RCg
3vACwoWo8If3SXLia7Y6sMOcQYiTp2t4zYOg0aT9h87ulWLu5I9JF0XtUYAv28XK
OyWZoThLv3SAYRy6J5Ck+ztPrMCoG3XbjoSx3edUlm3PgNij8FGU5Uq5/um4xfBJ
NLYmZ6P6yumYPL+qICVicLGSQ5KqwdsLiIsf/Ow2rrvwdcmVFi4+dwVd8gmkshrg
0Cuy7nitF3+xynoqsi/cpgE80nA6d5JevKpTgIGRzvlWmP0jioCrWU3HjyixAYVD
BdX7VTYmhc8NFMUyXU7dIfj+hro19unaPqEvzagRPTkPaWjlVNOemmfPvPqApUND
mWr3uLGkGc13CvgQybJdPI0r/PiKM0ewFqIQ/EGmJGWtlOJDkcPAUUwJIgk8rZOK
W5oaMKwNmkLdKARju9sbaktK+NuzGQTKWCPdRTRz+ExzIGOxHdUIzMQM33cuNy0/
iXDrVwzjrGjnTQcWePrAXbK0XplQZV5cRNvTJzB8gpItuhfpJNro0Wk3ZgpnnJ0i
MTyugtoRfKEzcTGbgBuKUda4pb6aVCA4RFJJopt+KyeI9RMY0/eSoL/nLcgiiuaQ
DnnEIR9hov/LKJiAiqnTYdz4FW4QqU/JZEmgkhRzBgIH3RnB1DNqCHxV2NPesZCQ
kk2BAAuS8vPpzsE0K956goeYadOQCgy7s0GjXwiTEtFbC2Zs62zWtaykEEyEibQ5
fMFH+lYnGqY4J3BRLa4yAjugxcLqx32TMe+sUA1zcekEhcUdaPedJaZUsbhok1ar
feK/XcK2/xpuAlVrA9ZPskNYdZzB3ww623sZNTj9xv8+e8YErvA9DzwTSOjkTXbM
kOBzRfxJXIwQuPXdocSSDi9RcRqkgx7EJww6yHEBoamE9J/Q327kRbGokK3VDXON
Gjb5WUc6k7+pTroSqb0JGzjRosx0xOaOL67oUzHhwukQ/sO9KnNzVIwMrWGvsu4U
0Gx1o23rUhXq7dn/VriJnDPiqoU5kEYIswhy9yU24aqL7rt1wO0TaOM0TPLNPL0V
fEkFX4Gdt/ZhHNLggNZgGUeNClmWQPuJWC6DYeXGc6ef10XLn/UnsYJksKA4KfoM
kKkyYMxW1cET9PSwHodSEm82TkkKKG4Xdkx97wqqMmQN1c0OsR/L6Cf8m+iycg1H
NDEn/BB03AkxoOqLu6/xeZ3GVQWbLm5+bf8cgeO8THUWibjMC6pwHE3jqBtxGDfw
KCWIdt/eCkg8ZBWf2Id6scAnb7u2CXEMbRtYNjVd/VIemZSJfE5mqL7ojM0usFvV
niWGie8nGEZkxBy+cOzbF3uC61OV0juj/VBhtFvZNhOK/XRQtFuycXhTJPSqtRJX
wzx5K5Z96VNfJj83DLMMRmnR45wCyPkoUdSLuvDfHiKp+Olvk8FoZdhpY1QSoAPx
tj+Mt+vxher8iDDsBHk5j25rieTnNh2t26Wl+psoS0C3di5b186uot0DCUvXTSYc
4ZzAwb1ICXWf22AwsjsGIK4bisUjUN14WOCqlrVc9atcdIRhAvpeuU+4BCeUbzwE
ogkoBYAOcjAsJfb/n9aSjp9fnc1POyoHFXmeo1IFW0d95QKt0+O/C1KlkSmc90Wj
QI5jlK3o7+FycG+tTwiok2M0lrz41xRzx8D5O9xMbrICT/opLQm83I9qy5dVDZCU
bssHwYDCROllN0xnpOLBZ5EQS1aj50iMXxtrVrw+svQdZ+S4kMINrqZUbp+ngKHl
lK3qEKkaaYhs941SnYv4B0p1kT0IPyb0esJkRdd0WYKXTFhrvS6gTl6qNLcBxSwU
AMrJDManfRRziUiCtRXyVB3vgf9E2Jr5bkYHkgi2vkJXZPq0yyWD43g88A8daoLL
8fsLJr7xAznpasVhsr/X3vLyOhCxKMycSsrv2qHlVrGB0HZwalaMQh2KDb1uP3kL
n+jvZa+7EG+TQTbYcvyzsnbiwDoHN8AvPMMm6HhmGJSfkdFrbwHj+XzivAvh9nXJ
3YPfKxosxEIsyWAha/vV2Bcs2UEAC1BxwbVC3xh1ijXkbwzfQ/5iIm632DNdgvBg
KVfz2aDyDetEcv2qUfhVHxQXulf4YMXD+ejG4P7ZkduSe2cevwaaZnqJJ54XExoq
aPw7RCrj/RI3uBBdM9vejpMKB5NMhDL2MHlTj9gKMVz6uspphRVLU13XPtEKfL2g
2YyL+bLrJmsOdNV7TlM1WHph64XxZwg9ERkvoCYPV6jknW2RKvwBYEE0WrK1imFI
CRbBriYpQ+5Y5Z/lCwGz76PGXlXw+oY/EDnGnNyMIlh2h/OdqcK9d5bJ7k0sWvsG
ZVUvMor6rpje19v8S1SAlNPhfa5VKszEDaYmAi5a1V4qKECZwc1X5rOQQUJzpUzX
lPFdNl0RCbGyTQOZGqGwyHZg2RsRbBxjuiDFnJykwcXnZ5x4U1Rr9DeE6a/x5YUh
WkWlAocqfpNmRsPAeSsywx8Pp0BCdO1FlxmqTavMhtUkXAQkN7/TvzB8RfkH/R2+
IiuwDGGr4cA5hiyJGsND7bQFAGkFFM1UBYxkF5YZFJVssrrwVSvJ+aV2ggIBnsai
0GL/WSAFkAz4pTiK7PWRREvlUnNGpDAzdzriaBZwMYqhVrkhMUPUo0gydiVvXtPf
fwMJSi0/56EyE/ewVFXB/oLtOe+24zvVTjGD50Xdyuw/GftLzjU2IYByEDX9kZVa
aR/t5gXd4qxbIS/Wz342jgoRYkwIViL3a9JgxHbKftNC16rVKBwkFGwuzTDsOGBv
876LvJOpK3CekCdlXzzZkBQAg7dYqdYGE7HtItK/jdRRljgs3q/kRco5hPIlTn6L
egp1DSlX4S1NH/iqlGskvupr1xcC1AVfV5I02rJM1NWoMiAGo7PWNxBwVyBb2Jrt
czh7JrhIh7ZvfjrMDFU0X5q1DXhFI7ZUqGIlshGWHTnLl0mHWEQPgzw523KINSD6
W3sQJ89+PTSZjwLirZomur7Iw1gRwdoSIsUblTPQlxdy6wtY8v7fFk6uY4GPXw37
wywcyL11cBT8mFtN8t60vzQ4NDKFJYJpPjmXbuNh148AKp7Zmrn1/t6j6+68qF92
kEjpHM1DUQEYyW2qSUB5/qWJ2hZRbzN7MMtUp+KbHgsPAV3PIaaotjuazDvZzx/A
pkW7N3tc9mUrbeS7J8lvBOVQcpUZfNTphF5/4akMn60cmgtTunW9UWJTqhDyEiAu
rjROF0vQzTwPZ6sGJO1rRjokCdYn3Gy24k2Mkn6twHV9NVWf0AZwWWQFv8ZDZ0tA
y4NbpCUPH2x8vu4hF5/vUzyvSrW3GV/cd8sYNBONkUCNGWQ7rWZeHyDfHZTvxky/
TokxNiJAtawBBZdKw4yslCCbmwxsIvsDVr5ANS53cPN0mrZK10E66AV4MhiFIJ4H
WPAhr8B2k4ECKZ4/i98c6v9gW7agBSLXFfOtsQ/y//BHildRGO1nKc8tcYBSxUZV
Z4B1+LfaZr1rTOgFAteYzxxp/tFWZ+36YHIylg9cv8yDTeZs3exoaLEZzOu1Msfh
A6hZSACa7l8/GanqHgq/Q28BtBP9GwDjlciEBtZuEALW7T+g1FCsLbKbWt2i4mMw
nd/JCEqFddc5rMEf0Lwtyd8LaC8jeoZZw/bwE3BgqbTyEZoimSd44KU+TG9cVneY
H6iY7kktjJ8YkKW10usdxznMl1rbDWSGczRr/Z7s7AvEpFjypirEYEOob7pqM7Is
GsbJvxyB3sLaT81ayVpbqIo0zXZdAJPEfNS9NAlnm4iAh3rj7Pn6aDdF6FxZ01ry
Tqc9FUtk074VRHUP3MGKTreMwzeald1z2qfdfeHnd6PibMctUhmZ4oOB0PpGhG9o
J5w61n2E4UAOmW5eimStbsnUXval7xetQOnGaxvcjZCJMkDEsqHTs7YTuDet163Y
GrMKMbovuMX6KpMybk3GQwkVuXZY9EBZxod7bYiRzY8yoE6Vjo4E16n+gzcb4BYj
SeDVoEkcjTGJbtpW3re7RiUHE7flSO5hW/WryjLekEPwts/FFluL36naboydYMe9
ZwbMlmoXKB0iFCtj+ywVw1Gsq6V6NilJtTV9TlLdt+g+8s/rc3Typlzl9i4s+pCj
lDDE1Hb8Np6hydZrmTX7hbW7JS/b+jj8XSeen8kT9Jlwvfqom7d2FzfeIFHPKcFt
7yZ8bT4weD9iAOypNPVGagDb6QYz4KeW4Vnjsg8R+dUkbM5ZADHMZcScecj+c3OL
97oZ+pqJDD8uJ374H2HLDZGTrT4kTjTsD+rPH+5Nhq+Rdn3b4nUjXQSZkbYG1Ytc
zHQLQ4Vkc/OB3W5m0arR2Ag92iqTbOapGWfWUu7AxgsMOwCLlujp7+C+UsjLSObX
xG4DJ3acrDjme9wRUhy26JQzdF7rHi9Z0udV/vJAXO/rVsVWbzLNVs+RXbZv0gxR
nIF6v08ThMBuNiwhNxByXa0V+D50mBotvssLKSe/aiyz2xGH4b+MfYz3Rd8VPLmr
e91YV4zGLy3RnFAsZyDGldRuWZi2dKN/PMfxj42s+piDkwDdm9LsaxWQ3bH0znmG
It/nrK24PQMCiqBYcpLcQ7D+Zry4WsjL8a/UI+Ns5eLDMz/AVU3FFZiCj2rDZGve
VRVyqCvynDTxpasC+FSQt8EJAdcybB/xcT+Vijy3zqXMrPh+dK0XmYbakxXYDPUj
ACGGwgp04dE/qQ9pzFOdaJIjTvKbZNNjSt+g52ZkpF3K0e4MRnBg4T7Kz0JU1gAr
o5lwfH3/HReXejugEf0CBO8QXsb0eRzWxeLtc3nNbrBOgwyQp7NEt3LlPe2XLon8
0rD9EwOi3yo5XVppXSwbNGbnkpED67Vw3K8Bh4EUXvbk3l5k56ou6LySKRO/O9oF
GL7JQEVqFXFp8DkDsvL/DX+JqHYqxu2ZiPkgtsgnXOrVvELXDHbWQlpoY3G6dX6y
yIKhuoE79gJX/8+Fyrf6CRdhS8ZpSyX4R4vUfCnTf/HPVqcqYvfu8M/5Y0C2zbTJ
1f0Ex0zGzBhlHmJum1CokdcvPbHMw6rZHdCqVulesOpne0H4dnm4W04aXW5w9rFD
6E2R1Jw3jEFbwaxAp272bD+3FWFD66PZwxIehncK+AjRQiYWFR5nQtm7jq95jU7H
MffVQ1kJPh32AJB0YTsdZcONDhSyyeY8qDunY6AmG66NhPrUEXZkq5TMnifOP8MW
jf6umw4H5ONuI0UMHZQ/7LoTC7PgAttwFyU/wUZ6QnTY8qb8ZOodb+NnSB4aDOti
2XpScX7yzyRmvStuMRZ+sbNCxnhlbTIjVzrwKOHXvxLmTAGLvxdTtYLKNwhDSw4P
4T/SwE3D5kwueBTmpHy7jxWBpQaPLU2iHi7hiwO7mbRnC6TzPeoAewa1GlTxCbt9
EoDhNFH5gxfOfqvQzdYph3p4BKdvcZX2mqfGeca1QtwDWFj+UL+ZlLvz36CRYeeB
l1+PvSqwknCLZONKhaxbNZMIUi8V8q0Dq6m7rKc1T6zS0a2Z/CTqiSXfap+7lxk8
14eO6iWEuihlYDrud+b+q3ThgcI464qW+WyQWddhJCBQb+8+6Au8JQWtAHWPF3y7
ipV4rwJkIYwgH9Q/LVpCepUkG7LvljseoYg9HRk10xKjZKxVocZd+28pOz93stXF
PbtjLMCaBldNXB6o5rp/cxhDfNJsTQzGWAncO37NQ/xTPQZi/GbdRiI3UkPbowFj
8H3ynN5lkcIAoJO/TeVxLpthL2BTBVPYeu5rv6yhE4vw33GAPlnvEYHZ843xywz7
nUMcb8kgXFresOmVtNTM9SwCq4b7wJN9QdiIGif0OD5vcgZn3eAFbP1uTHdXHM4O
i7enbIBNxOsH54fzhA+ewAsswwShM0o9jJLkQ6f+JMtozeDjXjldH0BYQMNIcc+Z
OUIXfM5B1k2rwecn4f0NMJHXdy6jRWfsbs+PDjkIf0UiJ4wrl26Psg+wIoOEy3Qm
ev2cWGWk0i7pHPnCf9wW6T0f7cTcx8klCEo35vL9xzsIZM54wUdkQwMHKpgd6FIQ
EAbiQxkLyChZry6eKciyvCVtSAmeUcMX/kodk3iv1sbZz8DKyExxm8xfQLsFQyMs
BYZY53OJXDsmPFJTAqiXiOb1K3WUGqy1pFHWm+fZIcLLbCVnVIquItc1CJupUsOO
iHCjCBzKRO2BQY79/2DYbosXeudxVnK+VZ3X+9Mkm0zowyGNf7B04D+l0qx2IRZH
dZSSVY65wYbYvcP/IWstNGiFcbOsufdtfRa/pu+ruJhp1TskF94qoxd++455Jz+A
SgyP3GutxFAEswp0lY9m/3IJDf7vwFLgnknN/PbtEDur3Zc1prEGXHwQAyFEFRdx
UDPgAk9DlWfjmgLShrhWoC4kvoz7fBsBB2SKjJUtFLbMjVI0i9f3QUWoODhURDzQ
9UE3niy9jjHpR/d2SULMPq7TLHMvGRQOjKoDQ8iHLVDGh0Zr/nDTRZAOk6QeJF5G
2MkYWquLVS6MaaTR9fb3Ya3BEVq15rZOdwRMSEq6b0Xo/AodcjOXMFWNCwRgOSBJ
j+ARpEn4OxfuFGaFeQqtV0zpI9EbqiHmEPRkScOjixBZlsUeSsLAWHIN+BIQDVE5
QCjqvMMFCuQgFZGg9YjGpYJ2o+huZvqJA5/IB22LGGkSesLdnwJ1wf7Z77wFDkrK
PUcW4OnOKGxpfR7xQPAsjcL5NoMA2LEWa+Dss+gkFto8NCu3Ourse472es2/VovP
PDk5/V6ail340PTzOjXrVhu+6E3gjEsSAOPf0pi8seV6nERRYFpJndnQWm60FYRn
1p9o7hjLSkoHyn51R4tjKyhAtmDj1uo9FbXN1sxjkbFJEskN3piv+dputp3IemcE
AsysetcpbSjhz8hxt3ki4HaxNaAomD/9H/pk4axVMj2iem7bZhw8S9fN+lXuy1VU
HLdEJEPprwTEXz2HDBMI8Ee9KoV8QDOM5XMpNmfShJppB+fY5DolQeth+GS8DyqL
Bl7DxoDylmjinhlBt5XVNuWdDvxNUdG10oowOpf6XODCLaMd4zloeyGAYVhOMRHD
B2u2g1W59SfJACZvvtbj4bN0I0fO9s1uOmwJoF9a9eIZJQu+U7xmR1q7nBXgM9O8
DsOMR5dMEEndN+1kdXxQQULaClo+7Sd/4AjcKDIKXoT7rSl7rB1/Ts3Gh8cEYLor
kWQ7CTnQ/HkV3vW+nijRDWTNN/kRcziJRREciHnT3eL8m+MJgS3XXtUXZXPEqFBy
VqRTHUwmdlHyTE953zU6PA4qTXqER7VwVqnUDehEjlgZiqBrCox/38+8kyUnv4dv
lKg5QITYIbxUb7yIsGiuZ7FMASaBNK1xhJLzZwgVYyn6cgTHeHkima+bfCTwqwA4
fHFi/hhZZ+r1GBD5YLJg1juu16p13+Lc364j1CbKB5aGQlatOOXfNZsc11OhWEHX
LwqnD6GuedOqGsdwpeW1Sua2UQbyuy43HiZCbBKicMmhhk/nOoXm8BhuKIYgtcFC
JbReMqtGtWF+5geJbB5rYMzhbqS57u1T71LaaVmj0aCA/tkxPqbYz3l576qnQgo2
qKWg+pAXoIwIVTUHnEzDRd4NFJEcYoIRAdwWlfVsECN+14ZNbtAusVYcK+pYDrQS
oiUExZmkfrXV2CAauNhcEblfn5s+Oq/pWjiHZnLZ0OC2tD9drP7ZfS9lcKvPTP0V
v+BOV7VNo+CMUEZZthi73eh+dlIWztCu0ad7uWGgE7EAZwkkJdlEQxW39jid1Ina
Q+pMpYHOr+ytniJcIbAq/mv9C8qAD7aE5TlEQVGSJNpfIojo4JRbtu1BKrRsX0lu
bAhUe6BQb2wHi7G/r2vkQZsgoN4ggY2ya5Djz9TRrAjSq5bP0Cvz+IRP+ousAKwD
mqAO6MU4yQR5SUuxe9JvGFANBScuri+t5vbEBMebQHAYIhIdDMV0Sk6jS63OK5as
Fq5oZG2elkV50y6DjDuRpxLWg35mbQmON0FY6ICRdXw7uGNE2zA60iognsJKZXpY
S2puoDQ2BRQ69WOWEny64l8/l1urSqZqwU2ThjkZko0rAg5feqRCfihIUMggkW+q
YyouIzwHEIwSyloPUDHRiqVqSV87Wz+P9GvfoFhqptSo57oFeUeA/LM+YR8Nwe8h
hrEqdbE7onDOooqXfR2d9sESqg466nSNfULs+5ukqC6lfxNi3PR9L4h3LJwH3N8e
/PjIKV4BEfP6p2fsW09gmVWFzICMg80qgGp+O31695t3xoys8S+LILVjwrE/o/f3
qUqVXtzIDM9p16unEUxQF65tqyACbyzgPaiVTo9TQI5BRRiSTewirbEdXawmAlYU
XLLqVmFd5lmr8NpQnJfroRTsI0HKuAaAGYotqxuBcNuX7nLU1yr2ZKA+wC1mYjDz
kbjY6/INzEuRlic9Ta1nshI8f7YdtUG4sEn2XrXKI5jBDXEgkMkIWR+rktt7l+NI
DYCvCQNMR2eITYW8MtoQe8IJGjt40tpTD0+BIJB3Zo8mAzSeIHwBiVg40v12fHRw
ak9Uf7ilvFFeKVdcKZvS2LFNZD3rbCZUAMdcBsdurk460QQDiUyBJR1U3vv6S9mw
az2NAa1cpYZtLf+y3SKqEy5M1YQp3hI7WfB6MLLm5jG+v6wydzjepINOsjhzInv5
EYPzC1IoCmb8ZOdqgEYEWKfRVYCSB7AvJqJYKzxTr9gDgtgVqGQ6Dt3x6QAmZZU6
WmtjLs2bt43WoJZaLwLrM2cMRz2wVMpyD4IrgzfizB9xaREnredZVdGOcrkKApap
zf1eX6E/dNJKEQQTHnAjbbFo1Y2dkC6ke5Klel/HGrJuU9RIYeAbnSH/ciO4VA7G
unEv/qt9rU+5HHlerXpI9q08ESRCpsWIsvOEw8aqzwpMTJrr68obGLhf4ML5vGpe
kT1qwWU4Ju7cca/O+pesRelHkdZl5eYoAYeBAoGC/Z39DRwnTUaJD7VL32908BAR
QZpQGOJUTU1OC25+srwvqubbR9eijNXyenHLmUJUyI6tckjFk+WBluf8bi3puBGV
fwiWdLdzFOlrlpH2skflCxh9lWY6edqsvuB0bNSJFi3iI42zkeTT5BUzjW4vy0G5
HgNA79NPv/4dsGPC+yxSotCkTvRV9b76f5r9mEz4f8rpkHxzQP0r6iY++sv+9LKP
4AKfaU9HlWwwvaMsMCzjWkBWg4itdW1lkPKu6LOVnevviMwphOLZjDqvPXAhXM9a
IRMnHFjQcuFbtEKl+iS5xjdF3ZKpHXwFIMo22ROMHejEHaTLpedaxFRDnlgRc1nB
gBtfb7IInrgFHMa+vfAcuFClqTAfgelhsBvlTh1p2ZP/TFRtXr8h23yXtlAnscLN
nRlkV3w3Tl0Mb07JnetUMpDKyxSLb5ZP6/eWHI1zD8F90NYwfMPB/aBASVQBm11i
an78Q96Itz9U6G4ozqZLX15TSgu8wEB+pRH0JePxMejpMitQF/IR1eUsTcGoeI2y
o0W5/VueW2Q3HzSrEwZlkCl430m8WuUJq85bg4HjBT46ihs8j2zKi9pPZd9SBNbB
HD/2uCxP/WzaZX0LBexPZzppczj8Wm7/Zk/K1U/M40bxJA8F3JqFsR/yS7JAoO5G
PICMA9Pame8hiz77wn4HlDK6CmlpDL5O9w7CMexsrdnKxTxRQeoNRKGVWEjBxR7r
RFMV1pJxJ82VxXEbWUc6+0FZSGeAoW2CbCwKxlXi0FaVH8MEGzHAfn12W1Uo1Vwa
S14WQYZv74b3K7FAZ2uPuPoW71u6veyaZEkR+FfRmxofxGlyu+HDt2H2O5cZ3/2v
pRpW5HMAegHkxiaNXNoxlewh044UKWjXb+99rVLEZkONCz/pYkPFnXsr+SB/sEd+
FUP8nd7A4mrQWZDZrM3QqY6YRqDVCoDwL9LX31/atHwNLYoDRGEjb0i3dCOehDiR
VGq4fDi0dVEJuHdWS0uMFKdrBjvNrg1E6L+2DM1LtNr8kb1z2RAVrxFJ9SmEBFCn
ZBItcqhMn1QOoFr8BfzuYNeUlGZg0cWmhMKEkAL1btmV4KAXF37INnSHz0R4Xs9l
3CEfMVuJxdR5FuMOdlNOboz3zOVxJEOqHznAi/BpYTXRu7YB2iMgao3i1zngRj2L
pLg6Ft3QR433ooR2xyWFLHzxaXZPSQVMwGFjdG05PpP7pJlrYx4bsufVkegcajt3
Sin37vrG7vZE/5LhNjJlVaczuyavz4eC+JUxw3cLBHUcxE439tYZTOnIyavmPfg8
elqYZeKE4tRhU+B9N4cwyHpPn+IX7qixpjD29UwH8/xvLD0/XUjefOL4oHJnTUWd
B0xWKZ5GEzT2cV9G6iflRthZJ/04bLsaWmJ44d+h/cLrYmHqp4BxWlq4bfWx6lFf
uaqIIw7dGLeEm6kgCbIuUuWwc+sGi6HEarXp6srk6uvdJiPP48YqMR/0MYcXXeDc
JV5srgfOvPi3xdgUyYoIPbC6yb5u3AMcXEurP9vxvapxNfLQd81OPdtz2kfGl7i+
o2a3EmL5UhF1FpeQOeqpEQXe/J889xwn3C+01VqqyupjpUmTmr+FhT50saNNy9Kr
4tzYf7nZ4GnK9JTI5ZUemFb+m9rb3bDzVJ8ym0dF9qxgPbBiPgyyN1MPXJq89WxT
0NiWF4ewuSjtO1rrdCg1PJGpYyk73SgdwBDJlMHfnkbGu5XXWXyAMegam4sbycw1
6DUMzpIznvdxaatHh+EdUAichndxCR2pNYxWA7ud6l1jedVyQvLtaQ/2LV2TFTOk
S/DxTQQ/TE/ggKqgdKf939HGXB1C7wGzQzCLnjrTec52h2+J177do2Nlfc5iWhGe
7JMovPAOacTOM297cfkMI8IYRG/q6J6jOAwg21Ua+VeCZo4tsSGjUKRh1/6JOiqR
iwwwr4jtFrfc0vVsAUIHBVfXbaaUIleqFXQcb/57wxMqWD8asED9bk8a9kuKlBz9
+096AnQOL+rG6sAivWRkYyFR8GgdW8NwsDVK8gWo93mY3XhGRE3w9/t7R7wKXOzF
itVq7gQA0jIIme2rz1nb0LmzUPhSCLWeZrXSUVVrocGAmmCYRCwUlYfAfP62zAGa
uXB/pRxj3b0D/oRdDfDQA8vz+3Tjsyst961KpoY6BpX7WPF83Bl2wrsGY9/We/ql
LapzhxKkDyvnkg9DqsaWJBaPSaWZOUCRluLWjvC9s5XZpfVVe89zxCmXXmyTzRUi
7hCX9WkH7F4BY9ilt9qALnZUp1+FDPSWBOBP+nVHIcmqH+Q+OMvz1l2dekodr80q
HuVgHybhpi3jXSeHVMBvqwhnPXE/shfoUwyUNPk9jPRuusj7QYyBzRIPomxQ0b4o
iPPzYhwt+PVMdjIIjxIQNiOzYwfKmxHkUmunZLQqXwH3Y9UOIY6Umj44NSZE7LD0
ymyo+ScfIpU/gU/oyh2b16CCqlYXYIIEbPtHGU0GEpji7N5x+fxpGhEN4uEmXAuI
v0+c+64a3a+JgIfaYM5b+cHHLA5C6fzgFV5k9wbU8Am5B1+U4YZoFnNuVmyBHBq3
NDayiio8XmIXgMD2FS94QNN9fFn02KGzjh1qLeo2czcFuEVGtK0TVHN5XS3E/DcR
zkXrOuLTyE8Ganrm+PvCNerhcJPmzsr3+AImMP6n9yVSi+7KHB/oHkcQFZk5cv/e
TQo9Juh9+JOD9IVzrc+hFuZ06JHWwDBlN1SI4NzHzFwdarZ0PpOMuV77k0CpGLo8
CpVKLMDonnCDflaPuDPuOU87v2KorMPXG/CmEGW8erN/eMnQlpQpYRO53c7mWiLK
SFV4HQXMp9jm3jbK5QyowPHlERd7grPdB63cZuX6RdD0fWGLgUqNAGpip3VW335X
11CO7ICHIOKsURkpFXRrHoPVkcpD885Mhf5vrgpSmhZqVHw9igbr55tkPDJN/hgw
o7hRvV7c33540pL5VKMeIsEAah8cPGRrIHXIYhp0PPO0z/IdLE4XTA2kfElCCXuJ
XOJrq4XNhvOIzBCDSuXs95J1h75USdaFlXFMoQkFjh0DIHPlKkvLWsTzPILrEzcg
DfSSkNpMSt6Q7bIV+BzlHJfYZNBkcDBmrZyURQ2ExIcgA4OKwMvSIqZH0XcG4iRA
FAK5BoG5Kw4lZoxEvfouB5hPcpb8l745kihT8sGFfBMtIO/kODUAI4D/ZS5W6RVj
/njonqpgsLET6xQx6xqmuxD2FwZZoe+dQ9OEs2K1Zrhq6u3ULNV8KnNqzSS6mCL5
nNPClMYahe8NNm/Ce+/RSOD7DwfL1BmWv8Fi85BradlAmWrQnlwveVcaPyV/4qxG
WPoBHflV3vme5LsUh3OqOAcnwfllojlh467gPxt9EK7ErvGtCkufkTlETODLLDC7
YVtorAnLWZMAOHM1rnuEewQs7fv9lZi73RSC0JH/qrz/z0Di6wSaB54Jndv3HeVx
qJN5qws3QEV1LYIRjlwe6bZm9G1VtoOnBqbwrjLu0dZaY5cIj2F0SqzM3llg75wX
wPRbHr917UGTRSODL5ipUU9az4CWW5jDNT1aPb7IfLIGF9ilkLILWzD5HLsNVZhC
n3R0pmkxEoQR2lYSEJmJ9BMgBn5tYUGkQZjH//0PwVpHIjgKypDS4gulmCurEnc9
VTNabBWpJK25Bi1+XawrmDQHeANBlYUCC1wzuM2QAJ+j0j96aIfIOpW7/lcpglWJ
aLgTxYk17ZWZy40hV+HZx2L8phv/ed0fGt22TMWYVuAKGOG+NCGgNWjVGWNb+Zeg
ocDFwh2bjiyOwCcggIaqq54iytjrpvB7fEEaAblKILiTMxTvvWWRAHxgdQNlhEgJ
C9yRkX7VVC7rw2GLV6kpnron7YxB0z9OXiFblPGOGyFjKCcb5xWwX7CZxK/C8/66
oYnyA6RvwN48P87lFut7fX85OsxC6Z3qUzw9B3PRM/BQbB+hs+pC2GNbtaoEA+Xe
zO12X4acxr2mX5Ug+uJkEUgIB9vy+edI3urtbg+AnBL+qSUNng77ZFrjTRANPjE6
dObYfb6l9PSdyq7AdMHXyE6nSO1PTEhWbDCvy5UzLhFDN42X+XZgSp7EdY/rq7l5
65bN2aBNYdO9akf3Asyi18m/HHyR4DnzvhWimJKJcfk210q/xlTQlV3jO1jxbxtV
cpD4FinLcHKw6iPTi6x5TlSsvudDElf/GkXK5QQyFehspmrU6xx+9M97tqTqHSE6
nWKIDIRy2pxQ1l1RR7O63awLVw4g2l+8QYeB7CfJ0uwL7oYFYeTiN/XYq/ByniDr
eC3E6WsDP7aYQqq78HoXFjf8aMyFO8l6sQory0tJtu/M77DoS8u06Q3gqwzAWUi6
Nj/j547vPaIV+ErXOk/xwEH0/f1IfSJxGyRfTn92FS+QuBCyCjXBlkHB7EhZGFo0
eivPLGAZBVnPxO6XvIHzCQiKdeVkkCUOjJlneHr93d2cROKcfed/WteGQqAs5YsP
hTOi8BlUZmJDzaKVthSz5BjihU01ZrrKcgwj3Wez04NPIQafc9+SoNbX7GCyAI93
gGkqSuknVABEB8HKHTczrdDVuu5Ee64KMSpKliobc/eUeTzNsxTATBMSkOKxvmeU
27yCd4ZbARKEZufyEF8bv3u2C16e7yrdjq5aFVdWW1Ia34xh6R4FmPngax+ZTOoH
O8n3VH3tVxIv3TsM8REaC0+yvU33WRFKUBmwj+gkIdP889s1AOzG7EcaH2oB+BpV
nK3JzA8t6OXNLzmwH/9L/WQqQGWnCCdLOoCRjRqBn8fkiZ4RGg2EPw5S5nvW/Cfv
N0v7jyMwXdwy4GkhwBXyWfKsKr5b0Yuv2lZCyER6JNVmz1NbTwJlFx4E1iA+yHDb
lQwJSHsGfkvuahVXOguIEzNaJ829b/eMCG+fzLDTqC/8RupqN7vlKSqWGd23gclO
vhAUzq38XLGP75D1r6qc/R4Oh1bUXfYLGf2698y+uQtriLREZslB7FvEYToScYAT
WmBNYsnxGUzVJ9rpN7O3/S5VYG9bnN3RLgLkBAPEnROFl/laObi2Wwory3+1Qwwr
W1vqY6F9qiqyLqpKH+sjXM9qOeH3ORaU4tQPzv7gt9r9CP1cqAMN6/DovOdQ9osT
xN6Vm1R07dv79Yy6AFDxv/uF6nABuPouF5yg4I7isDmytWCtD8eIk+c0v9jWEecy
9F0t+XEQNBSLLaVJAxBb8AZMGqeuDYsCLlmSoSy5vEHl2wpXI1vvplt6VfOr3ZwL
huzUy5ngzLX+bzGfXkeOjtXHuOZWHQ1tLqG+x+5gjXVQhujuxczYSpvHHBC3rShl
rbEp+E2rzVgBuzkY8+hJkDFnT7T1WYDqeJQpIkU0+VFl273AHbSbdebeXlQZV2xz
McSldd+bQ5+rwjJFv2vJuTxUUsTKtCMRvW06gI1Lc/3ZRit5I/Qckb+D46NPt11L
WxKqzRZfmporzu36MGz6CHl/uA/GHg6gnF3656SCo+ltvhDj2/gRfvj3aeDtfMSi
3RZEQFJC7C+gqMgyUbiob+fKn8XIs8zUvRbnuaTFs8Jp7d3vXIPqpq4gR2OaM7sT
HGG3a0MjsTzxMxkkA+U8RenPTju6yYFEGcAAvYWFc6KQGXuk9PG4/ABGzTzT5K6r
sBErIBdgQBiatKG0lppqSsjY2Ic49kbvvztF2NtyP3r6ZACPpGhkHRpN/ZlCHwip
7Ru/SFWaner/bBCCdoMq3QrxvOiu4GRaj8JiU6orz/iira0EOUnY8h+SbMlOrxfl
/XuP0tQQiYtLz0thuGS4KMD9AqZqa/ZwRvZ6fgafRjQFD6/+RWDY4jNkZqI1X35b
i8SxGBvlHHuIhv6p4UUB+skbCRike7al6LG1sPRBOSwE/pSMR5mStLhyWhxppDe3
Y/ML7342S/+ut/GcGtjGh9NciJTiHErHSlDEAS4j+BAmWnb+ncp684KZeIarXPrT
iXJL4J7DHj0jUnomdo/mrw7NUZSm3uecoRCInLeJvQS36g6B5ouKuXZNc9BO+oKL
lSMD35sly39Hx/mOQZE55fdsPPI3Fd4yU/D2OnWPSX0cFH9pd1yC7mMNLzUH+66z
zsNqeVttxkBSVGFx9QXrWx7TCb947mCKXA/c13Sjh9UvtsQzL6y8Uno7RTU3hCV4
ZCUuM6vHfyDuB9zYaiy+5qcpc6s0UrEHhXgWDiTRqwL5Dmov4zh8NDzO6ut4+jAY
RJx7fOLirJXqP95ZoNt01Cbpdqr256WuRbCpTs3zMYfj6gIV++ThHqxi2pjJEqEJ
eFnvws7DYdrWi+QEG8WQ/Cqj1W5Mpvfu0NsOlL/VXFRjl2KtFBXnG6Pxewl5NDDJ
JX677kWeC1DRtg4zor2nHvW2Hpj0d86pe468Mvr+oJg3NK5LemgzUAHU0azPd0nn
TuXyQQHxY7W0xd4LFM7nUtGIvTgE623bAoGgT9+Gc1CWPteAEKD1uJ4fx72gVemF
H/AfZmnPwindNz9Mzp7fIkNdXycj2IPIEN2im5Q6K+IvKalCrhCiPf+EQobxg5X5
GQOy2ZCnuFkFepkNM6y2omvP0Uox7mb63J3hwJsiiR9SsJWJFIagy+uode2ifofW
izd0dQnBqHh8h2kiXKjg5WQb+9s2Ym7NFORF0bsTS3uosNEKgL0SHerm9ffXvtQX
YNV71wlXjf5U5eFbYNi8Q7i2+LZVDRB7oBnrpYL2+RbW9hduOnCIyVoAc9rvnQiz
GlxXQMxHR/eGmFH9VGqxEv7DCn0+LPUpfN3QNH3dSRSJr/J3ys/RFcI6q607d3uY
zSfaF3+9bY2aY+HqAxcvbqqJVk1/qkOCQSFE5ZamAe95j+PdBitrAc6GhZK5IGxC
NKEDxowM3QznmYSao+99nt4AryAcGpugpiLCuAScfebJzdlgX5WNaVTQY8PbziiN
2MH/v8IW0n5lCCS6OYzL97X2ddkAfFKjlJuAYcgLG6fq+5JOtLJG/+MZ1V8tbZSn
A2JrMgKBhjkb8YAYham0T/gLT9UyeAH7wf0QW7JgX4cxyURxIn+6mErWFoMFQbDc
hay2MOvX3gKYeWOzqYLPpwf5v6wSJZ6UlUN+H7nD6oXzzes6M0N7afuGvZOfIdjP
Kxta5f5sRFVoo1qYh3I+g+5EI8p2Ib39igT5VdsrUAEcfA/JzFFsic9DGIQFCvZx
kL02PsE6z+Da4wkj1gpLenNgzBPoajqDvw35upClJ9b6/NwdI5SG+SjlK3epiW7Q
wcg4KNC96mvtj3v3mf1fAk4XRtYq0UUREP+vFrXGrRFZfbiu3ky5/xocQ9lqkOO/
XmRzppnJgfWh/F/L+QsyeeuIG+/fDWzFQROhQxC5FmcDT4GocsRolhZ3nJhEhw21
NVGw3gFmGdI9YFzATsmgp+M4onot/TDdPMddhYW45aDdnrTx/xNaRd0HIP+Nar94
7BGON73mXqw0hpVBvPLuz/3fy33FSiH0fPRYOR2yF4m0UAEDrTq8k2BRedwaWE5i
tcEGvD+gpoIYrNk1W8G7fpNveluulqRT9zBDdymRy0k5Nc/mMVdXjSn9A8Sdzrtc
ZQPGgH1z6Ype75vKOlJ7Dc/cZvdUjXy/eTsIAzKRWyvFiRyhz5+nXewrMstDh0hZ
umk4FvsdkCeSHcgwJs7PWDua6VPJ3xMVDPK0MJpAJ3PdbYbkCykoVR26XTzEkDUD
tLfvSJtkdBTREbHX+SxwAxZqQFEd5gw62kEgk+nPhIxiIDWRbY1qhIj35QABowiS
nTpnZtyKqyjdvfIJ+R/nYqbyRkvAvAXNe7h2hUXRvufe8XVHEuL9oR3iGUNcV4Sl
ls0ifiUjfU/2UL+ubs/FaMrktUm9SZjKoKO9SW4r8xTrjVvrNMM0hKHWpweEGZlX
GX16H0Z8zXXv5IF9yzusRhaop8f700m5aA39TfyEI8VJ71B133PVTCA4Y/w0F83k
rvTzSwqKbny6Wcfmj8rBOvwA3uuPy1nQ7ZTpwFsTjjCh+MhCC3QmZn8Ze/S/bMpD
nmpAIAQzz0sT5yV+lNhLKYsVVBtx32M0DTj2HPb6Ag7Cj/IPkJE8bcVIGcszcaq8
iuXSE8iuXlB7YtjY1LPuyiu2yKHKxHPHk3Ln05hEFIfTNlzrO+vN71TSMyW2JKbP
GmlD6uAwwwsaIZPR0CNgneGhZ1gMY8qI6dU7Psv3QdIT4sTAa4Ino+0VPy5Wpw3W
VofU8vw89MwBbM02D9Ig/aMQlDGLMtqdauMxshQjMUvlobZ752TVtgAHf6K9LqsD
PyW7vlL21Cz80Nt4N4tOn6XIEkxK+jb6rU68mOOu7JZCfG7GPocruisB9OPj5wCe
M3mO3lCxyw2tA9mJba2oM0CslDTeTfRKmZ2texCYK4QgVqd9/yI4uuc5PHZ/Ei+5
GYedH2lZR1rADuHfnt149xodXPc4UL7EAySykWp7bZbcSwZLFaxnSPbY3QD76vje
nXNqusezJto3Fa4VHBvCPWuI10M7vsBmt1RZqHb3LNQSe5rBMKiGxuzd5qGIxBFd
4AgXTs5pTeMlxXCQnZYGi2JljsTeoNMNrZCQQGkA83eoMdDhLZB8ph8J2soHolHM
0nyfngqsJZgfyumchGz/jhgx/+ejDN6lXLxl2GbGTxfeJwYE3MPkj7FWd7f6zRq6
UMmCfzAmnIxJdsF8yIo8NkjwGwvOO+kARNxfwIQf0dLlkELdLmCpqqwcbnDb0r6V
8iMzAaeK857W5hwaXscayxKpWLwoxgk5VOkwBafze/NUPwt+EDY9MoA5UMvPxKIF
GTMuONmAKRHdieyF2j7xTBNuw7DPHimh64eZaumkoF4VU0T/BFCGD/MgJbidwk/5
bwv9QAcOe/C2e8x6D4IkRc+ZNAu6mQvarRLeNDetIwcxjxJRTPesamjuRG6xg8we
eChha5AdUXsq3WIGbnARjjgzbdf2/KTL56tL5xkT4gbMA8HaOLpBpOkdGdUfGK5Z
Za5JGg35qqhCZhw4Tfcink5Xe89mmrBOKX+8vw7FMaSQQDmuCax3gW6hl8dExjrC
vslqzcgge5j4nMhoHh+Jjlj6vjvjzliHzvoD/XXBVo0NXFTZJNIGRK6QGa8mTyIZ
Prp+xONBPDAee35fTzxHv8OVmX2pgh61RTbOb9gS/I8i25BBNteAyGwxF37drLeI
Tvnk2JCsp+ZNBgG/PSRxpXumdt1yaYMe+kBDxtp0JgUCM+V5VZKC4haeHC1UmQ5G
S/RMSA5mxX864eEmOZ0iHfN8BSjPJTDTVMj+3uzf1NAGaR6ElJFhYzhG/t92Wcdl
uh2OSZXe4b7L6Y+YU37lGHj7DoxUObVS7orzI4nw/l2qV4BGNm4/CSmeMxdtZdQw
jAU9LCIbStdXMRnpJknG0it/RqgER+tACJjehn/ykEyzIZ4dScvAGgBDX5bHMeUz
MppKFq7Wu3B4VC7ShqF3nHwhh5Hyouu7fOejHkq7aGOZ1ZtgVIQL7HoW42H5wZ9U
t04KNKY+vm3t3LAdFn+pnF2/ErOSaXyJsMOCrKsY3kK43WpdAB8W0tEjTAIYxg3y
yrk2CNqzjcE2kCiA2+rA3FjmrKWh9TO2s69GK3nMb1BQ8egvQYGm9OqpYZAEKK70
9VVRpjsDjmuAMCy/i3nsmjh+BiQTXUvsldNINBVPz+FHjEXo4vdVeX1VhE6LESCb
VYu0jfDjBgymF6R7d0jSyCjcTn5SpCCcubxxbtdkGJCbFG0HdpJ8ikp+ZDeIMASO
BqqVvxAEdECjfpXKpd1YV66BLOTFjolr2nvqh8dCKliNbPj0SU/fD5rWsmgUKqLy
dynlPf5XOK2j9JKcW7YQmuULmKiG2w3ackkj8iGjKlKbl58DN3KW02svcYo5kBMw
XBj8vN7UmTW1CDv5LD02oXMjaXt1WuJbL7pS77RzhD5D96FXa/EsznVzciRLmY+y
NsfsF2IMC6yKgBoue2v0HRdLL82qFLkQbbmRkCrHOF7mxCXgtHQNJ/qmdORzujsm
k+j3tLxCJhk7uQiU7bRo0VN5zmYs/DMg7RV+m0a1z/w42opP+qIAQc4mt3DBXg47
fpTR8rNwgPBYWfTPdj/qB2jp+jNny+l4jSIrY7qum9c8SJOki+0Mz5dyyItfdv7O
DOJ6gvMs7QGMMO9OgSJEYH3FMOx6k2u4dcACjLoZOan6M42r7+TASWc0mSuWyspe
AzMh2K0A1DfNl0OjS92dwOYv7/zcecMX12YqGBBdHeoO3EXKaMOM1ESt0AYbdv8y
LPd0YsO8jgaoM6fW33h34VoF+gda0v+rbEUVWVxuCKE3fpC0dkwZnzbFI2nULC7M
NI44P8wKipaDvhdS/VBw1VG5Pkuolv/h2WCmSbgKW+dxyFfl6UK9FiuQ51MlaM6B
j2+CfzR5XjT39YqqiScDtRrjrdXxP/HrOoZRHtilxI/LQzfK8/s1M91/e1x96a48
0Twx0XuKkt+PKCg7AIwrL4k1TUkJWtMBsdsOLc++r44ras9VeM4yMfWAOntUBw9h
vwpewdO5iJVFmXkANee9T0XJ5yiizs+MR3RyWiAutE2OhtKxDQBJHkwSGlbrjkSa
3cnI0WYThAdPtd+F5+sPmoai60wVI3/wzyFXtz6mLDHNA+uRAuj5or97l1Bh6F4k
KOCDypx2f8VkHkK55o1hRq7wvhd8H8epMPWqx69uohkLGH3LgrKsICkdoDgsZt7O
NipzsiuREgOMUWMdC56OY5fuzedM5fJjU9mx5O6uVMHXw9tYzQ8HJYpOIFBbzTJq
lzo1ljGXD47/q6JIo1P8V1qB4UV3KoPiaFVWVL2rIonhPi+yUZke77N7djN5WyG1
XHz2Od5o6aEz+ilo1iUafqswgsvQ+8/aK/ecP9puAiMi7TeH8ETo0nBGaQHNsts3
jskVYOKsTpUZb5Tn+8CBGdDf2+793M09Xc4PRO34heRNC02PwuwwYyyf19hLjvsP
dvirKby4Ak65f8Mf1NWnBxmVUNv73dPgET6kHBqvfb/sdgQy+4uGDC3WJnroABF+
tiPxTCT2kH+R2tdv7RijGOmmQPts9lyTHQMKXYBBytMHZvf/sfqAjoI8phMEh+8G
t3kXP7OCZ9NZeUxOxt0RLra/myxmOJEQXz+Bfwrhdfr9DLLtgdtGMiFGwBEIxi9R
+44HwDvultQ1iLvF1ArpVeJ9Jy1+6Kkuv1cIJFGUYjsdO5QNKKG6zEr/N3LzOHxc
OT1/SJmtjeub4wxCy0GPnRA2rFmnnpGrLkHhVJF0bmbr/tbBMqOmImZ/qa8rvn0O
z6zRhMnBNigrRSb1LcjlxsWNjMKWEpoI9rEo1Sb0YG5dVGRee6Q1oyV4lCWzbzFs
95oftU4yPclKA7uC1R3gGbml7nQ5gpbWNEbXzwP6tpVN0Nioy/m1wDmg2GrHekJN
jZ2gCU/zaDcpyVDpRKHG01HM0puN5oa7ohYegfb3m5Zw3A3JnVe8EvIatChy/ue7
wAV8wtVAVwDRLaxiVs5Nfp/6OJcVZLOhzYGcpmncbieVFRKJ9hEvFibbvBKjBZN9
RrOPWA1R30KEcNqPDgpB7XF/2nv5K/eE2+s6j8ZlvALsOveSFuGF/yne8cipMIc6
J12bvh7Zwh17CJyguqxW+d6GQkRKTaM8m/VFenW1TGHZxiXlUq2fULqu9urTcjXF
J3IlrNqZp/wKTibCrdR20C5kHStkWbxHUqWuC2botyOiWt3tOh80vKUZTwlxwKO5
2CyhfpuZ/vdEk6SkFtwZx173Pbsur0GolYxSKTG7KyDLsgbeFxtu1iodWAMnopTV
qedjSmZTxPm2CgQYd1o0wsdbdsI9rMMMtxTQhedrcANOiU6eDNIY/WJ/tDcqhP9N
mmfILBdihuwYqrOOPHgDcvJ/TEGBgMT8/pSRaYF5UVhbQKhzw3NxFHeoM2sjUuKS
3YsM+4AzWhIoHuYQ5PRJXJsoK1ts7HTXNr4/9iIf2TQZciIF7LbX5aOPE0O+gtTN
Eju8ia9C2D2IJCiOjJcjxzY//1NdOesSeCZgjgm0twP0pu26p8gcvsUsox8gSNrn
rjacwVMVVgtEZ8i4zypMpsbksnvJlFqrotYGIDtSVFgbJvdEdN5ITOlagvjhGdZS
voANE31LjB4g8x1DpV8LH8BCTy6uJ6JHsQO5Q3V+Gsu+KiR+xWyzCw2CapjmnW10
c3F6Kx1QycoBj8QzUWAmJIgsh8iAZQ+dgaIOHVM2o/6u+bsV+uXCaTphXFLc3eC4
DzZL37jYe2QGbliBPkhBAGqgJPpWOBQ5PFtVDPfF/0IqyfKX4ZgQAA8hoCMgYvNm
OuuShTFKBxiIFJ5/sPtKgrqPrulB6i9jn61W+ABLLkSY9xraqSPIxZz06xXsXfDa
9ayRa4oN/1cow8CW5M+GoGTuXhPPZPm/clZL85yeyFopjAvwaiz1aU3P9J+nhZlB
AzDUGN36Dh4GhLeNTZ8tegmBVKOnQzlji5CkndZHuWAohlDr7/Ng/4lmD9ZI31CF
pMjYJPpsgnuvfW8kZLIHvj+GolnqjHb0Qzpzvfcv1TI+LKlpa3M8M2BEwDrg2DwT
bGsyhyeU6evzOz3vPUboNEjsIV3iEALk6Z83ZHcdcYG2ABN2TWIWDtM2Z+9fTq7D
Phc3/Kwwl7cLTQLedu6PrfzAlCd3i+Ib5JM9s7PIpB4a6N5sFQIig1kV7zxyXeWd
Xc0KGJTgM5VNYkgc/E+K7JPd6Q5DgIYj0vwLx3SfzbBG17yHFWeG7mPr2n/4e+hC
HykpVQw9DiTIwXr7NI1PoQwr1nrIRLUwXnJPsb6nVKUQcxgFLadQFnVs8WNPqMpy
gxN2Nqca9OWswCZ9/sjbiHfbneQTL5EVQJGXccLNCA7rD2ny206UxC0mUDIEwMDM
bQPitN232UUIGWNTGduSLue6WsEnr283cEiPSsb9nQVcDYu1H7QPv8MUy5WnrYnd
tJS82VarTmZ+DHTSTCFL2C/DkRAx2SiquMvXcqazf6MKn2viIapzNlkyIUvjMHp0
mH153aN15CPn/DX9SYmZsCYeWhBP2TvfMr56oH4HFl64bIfqurNKoSX7MShlmJqW
rDFpsZ25kEp0hGZekTBG8u6wDls37TsPApw2ikxmhSUl5il4wTij3IPJgQcYpWWe
dVz1z8eJKoZSFso31tvBzedyhzY4t+iAflIGrXcacVpgyFjtfNAjKbpHIwKPWscL
h1JDySUK46k7rjIwseTdOMcqZivIeLMsvC5VDyoVhSOPkvRPTSlFo7FHFEXO2oe/
D4alrZ+q3mN8qmosI9KWDDgCHYWMyVrecmURmdJhhk83etuuhVEjKSoFmE6kWHoY
LZ4VpIp24zmKxX/S7Lw6VUchJnu5sXJhVpwlyc6EWYgbXZ61JpTUESdP3Vrd+2SR
BkVxcvYdsIYGIqJGtCw8uoOS6mlbBYg49yBHX1xMvx9OHunOlKfo5k8gud/c2hSu
h+/I44v4iURgcq0fgWrvkllgvkWtJ1X7cG5hNlIbMFTVPlvLYNZ/9PgZ+w9YgPd/
nHTaLRwMlJwHwrXw96Pgl29w1w2nvkZHednes3pcwjPm8G2Klci6jIQL3YQpZtPQ
coCyW2dWuO2daHxlj5ZMIsFglvKIzzn5j2Hyo9BNYuSdeddTvy7HAoaYJMGsivCx
cKl57d4Be0Q06TU7hDNh6+gMM2zum3XDwPWWc40B7nxrIULUJUcEPhM7PBGqfWd8
Q6rNC7CxIHImEQrqOod9jtbond+AKHc9p2ZNBpYiSt87JeYoHfB2rSUba0hjcaD+
kIgyknVkU6HKk8dGQaiassre3S+8YolCbdaSDwvLgnr0WElQAdLbQCt5ZIZmRN6K
yK3uBTaUbfrsN8pia1ta0T5NHZGJeSdidzVwrA8Ijl/OXy3q+mYocFgnVaxBYCM6
JA+k9x7WIh6GKdpRQrDju2pjutYUtZUBvbO5+2OhWS/BmyZtVVxPwm/IC6XTz6AF
BdsbMY/7hrcc8Vt9JG+Qq4FNNx+JgpLZrJwcRF06z0T1HMZmUAMq47gTkeikur4y
vrnn/1D4Ripn9FM2S0v7PDqMdisH3ZYa/lQZlGb1ImJtswM1R7zq8Puwfkcc7htf
3nv94v5jykjI0srITCWVjGJLh2yelce0OjasmuPKh9NDUhpo4UyyrcXP8TolHGPc
FWJeSOxCje/c6hZ6dXF43Ug0HasOrrrzb7J6PmwRtziRaURTQ28YlscBQ/ahTcMb
SO40Wip2HrcET6zR3a35GFsc/yT1vuFTw7Xp7fF+06R2gmhaCU23aYAVq0piu8th
KiuAsmobdMmE8S6PAcZXyj45xyU2NOXYuE8k/FrL+vf8Bhq7Y02rXaB9fHD4+qoo
pFy0sl+KB898cUb8IHBWldnKi7JX+ibzwZwpO3YWu2BDGZvV3LmbNjA+SX1pJkJg
ILPSG+RAUrQXh968ayxAmIryhwGohXlu4Q2uwPzSnqAOgKiPtKIwN7037RHPqWOb
mtZxcDG7Hj0wmzXUFuxuu9MFsUQZfWCGlL7LmOfwBAynv73cs7+E+PdoUk1JUqBX
HmNG+wB2OijycLVy/vb/fr3nmvkMMHrgnHLW6gz67qBcXQdKkDfUAe+eOofJ7ABI
DF5YAZgmhBw6+oH+26enwU0VNRDVcjVV7WaT/9MNrdQKkiRHvE3pxvTzpDwVoxtz
qqRVPDpuU29Jy4dqzjNmMMNdybZb94c51shFJ4dTCsa5mJCc5174jkYpc2FOmt4V
xP3bDRwDa38fpgQS2o8CmATzNPKdxBRNoYNmWqBQXE3kEM/fwKgeyMF2hZnEkEL9
ElUasgFKAV0yBQMjO+ti6VzfiIoxLRGEt1qK27MWJe3c+hqh3eokS66GRjaHyPkB
oISLjT24rTB01W2tSLhN1PKIhD7FyIxoOxLkegxtgf/zNWzRBgLD6JjoTDWDuRBd
m6ii69Qc4b6cVsrMQAshmmi6gAA0n+A7E9CC863zaMqFT47qjMBsqUCAiSNuzvU9
9yNcqrJsw88aHO5Hr+N+pMfSFhLfyCITzArOQs0CXGX/2+xIRSaLLigHaGQzwAOF
vn3e9RnU1XY84FgFwiQ9O0xTmQ1EAtpyn8e52h9NuPwMSg1EoLxzG1D8vK+9Q52I
5t3/0fRx5GEVAV2DNddh54Gj/0F8m1rfioH8TTVMu1RmH5KksX/pLH8ZjTPqKFt4
euBzlWc1/wdXgpaPgwK+4h75ovvfcD0SNWJOQX42HXlqRKaDndtiFl2xbhq5uYtc
1jwyW6mHVgcuuX7btDrdc3zfV67pRlszqd3bInNq5H8VIXdariV85EznomeSG5Qr
AQCC0M1s1TZhd/uNyX16UpOZrJROL3MeNPVoRlCScevtHG4LRhspR0ejFStWqV2B
awPvf28oAg6GrltPKdB+IK2G7RmDqo8X0V9uhxa4LEKohG19SMI/PmmefKTKjaJP
dLo3R+QcM1SFfoA2/k+jvQ20aoo8w6QA4Y4K7yUqEq9ZXqkaTuquJ14xPBQT2WX5
IMHZtDxcg8wTXoRmEzcqcivc4Ixh71xAyiZwziEaTFfj1PzOmyEYr7fJeTucJrtG
8dlROpMpIR8yHVw8Svy/0xi/brMiB4hNqhwYIRXmgk1N1bGVUQOwiMN1vLwdNkdd
sqkpgEoPBydxJ1i1/fp6BIRkJvQCQ2j5OpDTEjJ5o7x3l5K1r3uJC7MB/u2CxlXJ
hZ2Eup/PpTB2ls30mCMUOs9YALGuF5W0zvtUC34r6F9pdcPOo6KVrieestKASWVq
2lHFJvPWyZYwi29xIInGWbopqfGYklwcCGRDo0galpj63qrikqBN8E0gW60dS69D
JPo2OPu1FO7TxYAocCh+hDLXJ2VYw+6ViTBljzkhwomIB4Ng78c/t+DtFxiAEpi5
9WqaUIhX4xv5o62B3yCEvyN2gaGRi91Z7k+QOnYNAvkyllOoJdidQyFEYbM/eOj1
/HJWopPD4A8pLuqNll8f2Z3Ve7jnXEts31NU6zkMe4iWhYWI1gIHklF7cqJJtG8i
e6wH0Yvz/6AHr4kmsv0gDpIcVvcYE4z7bijem19b9IlxCtjrm3bHMFxNfeJmV/7D
uAWKLjP30OClvOOK83QJzNv6VwYlnQ5ZdXsMGROrlFeRf56ZBNR2jStLaFYJvsOc
zmk5H5pElD97jElAybZbiBoL3ojHmn/x/lltmnLRll7NEr6XDIsBWE81H8s2J8GP
EL69Wxw9N5R0ohZVaww1Q6qb6BuqBIaJ5C3LtFB87m0MnsQkIz9TYf+Lj7DFy/D4
p2iCrSM8GAPj4ybinUG5PjMB0K7A4dFDcWNn0pxQqlt8g31vZ7O325dtNis2dDAU
RmSGVVNfFYRH/36+6y7HC98nYKEbzyKSGKcsWjVk2p2v+pXfW3yBdbr5yKkagvv3
rZEXJaAqfYpvVuPkV3exC/rb9dWJVYj9W9PFUMOtyvZk8boM/0jaPk1gvMug7xRT
yG9NRik5je39M3uL1Al3jwFpkKDbqub+/TbQ5qCN/VNdlbdBwzLm8bApOegT1QHs
3S8Dof2n0S4SkAUfA1uyjuq7iq/jOYcnCcUMIsGhN9OKs3KTZvv625o55Nq6SCZd
tvHZigXyt0F1fiZvmG2W3fzybRoVBg9IN0M30JXXPatYxoR9xTMXfRLgOwvOSI1a
mnQkQZPooc2jM4d/+3ZHO4yzysTZ/nwgrnjvC6zStk3g2VF3boHxgWpG4RBhDTG7
2Mh56/18t3XM/Ps5XINk3qF94SMdsDJK75sAz8v88cuVew8KsxMID9DgGnEEipKS
72HTKvI9gyhZbuPLPfaUDWKuzPrsKFVmT+swdkD4eowetieFzJtWCjsSWZ6V31SG
2WWnR0DAZrmPrDATfSHaZMP5vurniX6lAP5mUjkeSlQYuhlppnHM0nnsX6gmu+KF
1FRJCLNZRlB/XuMpFPg+GUuTvZFIXDquLrVZGSOK5hn6Rv4KD4AOMCkbMMCHkxE3
mNFCT6fkB0clwNZzuU2O9zdPFJpHeTAUSTNT7swJpF+gccQhAsRUhSMMQhsJ1XxL
VFDeSzta9aWq6HrfGAiTtjxbw3wFUvNmXsZ49BvvL6N6COQRQEZJqtgQBxdxbBC5
bu8Yc26lv2wtUlXXY7xj1e4lRXmMu0ZDSbXJ0GnYRJZCrQa6OXY73H3NE11Yn/Ck
jcl5EyERyFNprmVBs3t4m6WE+tqFeOGWV9l17hGJQQdB5s7LClUiTGoEbILm+TWT
mSmAxi1FvL+zrTHkZlxnXNFoGoRNngQugnp+ZnR3c2PI6pF7IRoS+csetNN+9Xbq
94AePafdPOcaOusiSAPEfy0L3zfjro0HYVUA8e4sGxRKT7rOPxpg9VGUyzKtBdVy
24M81tTUCgCT8jcgDGKDsZBBNWpaML+nrZTomfF+JHTey3mb+5iby8S8LGv4/jxp
QxpsM6Cc9608Bo0CB4JRR5YClQafvRClQuAztx4MfdnjT1TMmd/z6FWieAndgJTC
MgjQVFdYScHjhPnkA1dunrMfWx9RbpTiLOqxD/37mYAhI5RsMgqGVGr8tA52wfXz
cpw+5tWJUzwMdgRNsD3gF97XFtCrMU1m0T74KduRMyIguDGg8p2m1kL8TyAXJQYW
a0Jrf4A1SWL8n386CVK9aa85sygpojt+ZKu+b2ZzdqyrS37a1d36jiyJgu3fpoaC
cHebO6bWsnppgzWzDRv3uj5W6RWI4y5Np0A54CVIGmGw2MVifBNYw/0HdmoasvGW
dQBAqzd8feB4o9FhiHZTOsQMHeHRL8WVSNKiZPH6AI+pgb65yDFKVYz6GWlW9/zZ
Y06fjYw6JxL4kwcEN0JKzGSZftvAS64kbtvpxI4zpNwdne6VLS38NMvzBjf0Xugq
+o46RWBp+vqzEd/ku6WZCxyzvEi2EAx/kD6SuENfWk3F0cMPv1xZyZsD60NVXAbh
SvWkZBZq+iZq8LGNkf5ZTuivNGMRUVP9ulJJB8Vq0Jod9RZEToGabMf/sQ+JwT63
3N8FQ3XBFcan2PsGpB/ZiX1jnCvGVbJqXXn1Q1mnmoV+Z0MyOx8evNhhL0QFVpLX
JME7DyTgiUula9tgt5FShPF86JQRk5zjBzQkODmzwZ+UlZeL53Ya3bs0/lQUdDP6
GzsRYNyk+y1lFvlFKbX9oLHq4OJuia1cjcrGSPsUA35fp/u4f8gWQkBNIApNu9K5
GMsJ2xLyX98NA/zzOtAztZG6ru7bYmKy8zKWyMt7anDBkrhmQy+3xYJuVDTrq/Kc
ZFGFUmBaf8XfpfPU1eK0F2BT+9/NYxvz7EU1LWWXtJhmgwYXO5YoQtulVY3Z1X/h
mQyJ+mWQXzqLTIeOBqR1v0/3hNaFXiBV0vFm+JZO8O+S49aF8P0quoK6sZT5AWGA
6fQl2GI2tHmWGDfa2RhVFag6q8Uu1INSnT7kwywqPmavYAQV5UhhNiTUkSQU5JTb
QkKbFTlJYdfbB0Z0G5YDLNo/rAQZ9pHt8gqcG4AcyHh1QKdH93pwgdXYONzW8Iiw
RTSJ5cPw/6ZpmGLl0WRWthxsyUUf8JFy+5xeceKEPBk6grDlNHrjWGNi0hDw+cjh
OvGSvo/jwh8wwj8LoaaOiucMWz+aixsq+BHfwZZQyoLSGEn0Oi2gkkonCQfhKdrN
khc9FK8EouclwyC1oQXwbehBt7J63PfWYypONnpPlQXGtOjQW/MCYnHzy/MiyrpD
HP56HvSa8rmZmGx+GHqUDriRANmIXRdVeViXl6mE8nusQWcmRRSHA55LKflpcj4d
ZtJOEnz/wFG+zsIDfqZj+jPluMOplXcDj30gI/0/KRny6IWmOkdfM3AqlLl97p0m
vgjpB8FjZI/0AbojSLmYMJklka69962WAKlm85y+JXCIdLBvHznml8JDUwTeRET7
OFy8o4Ur4Un/lEsItqI/XGGILmro5A9mxiKwEDoIY/pSNeJNKttKywctOe4J7xds
72OMmK6NRZKbXDwVm2UbS2wz2ixGreoXA3ufv6yxjwLedZ+k8eK7ZYybsk6Zgf+p
dkDNtkbX8kXswf6cjlgiIOD7RD0sDsuvHfLmbtMlgBNlQBrRfbQ/qHtyNouRb/9Q
U0hRnOVcRAiP+WfNBFyIpPHwoNxQRmkfHrQrrrcinhTzHiFhQ8JSAkejZLa/fV8a
xMaBLRJOf1GIlYHRQgoHPQjTmpZ4XiHZ6J4f1dkEFWxWPiQIRF8ZKa8I+fBzHEtu
A9qyGMCGlVz937uMaV1De5qT4kMCdyLlCreT34U/nQrWfQX0wiIDo1JWzGFovdd/
hrTYJIJk5vF4Jm1VhlB0KYu9ojBMyuOY53dr5LarS5D7jliZca0x9vZmb/VKfCG6
Azt+dZdxlyw/mfxmOtFE6712gwNXnEIlHoQZO0DzmYdvdEjmHnxJmmFAYN8VVkLu
V6lm+g4bb45Coh+TatF617BQVNJTpLS8fWIrvaAxDg6e9Kk1ECZBkWXMDmuNIasl
TCkNv0VInK+o0Yvg8Kvlv0G8sL+oU3xbUuqoPvsEdw6f60y3ObTBiSFnjGwpWvOr
Mj9L46YwYuXXjr51RRx2IxNMHyZzpM2lTmNUIgXKi3E5+OziTOfKMQ68pYEJwknx
bX7jJujh36r1DAdvkQJQXV3lyE3ebjZSDHpwVKKqoqB2d1zzrDcTvgFWOpHucfyR
I2f9ZazPURGTr7r5Z4c7W7FaawYlLiyG0q9ZZM2xImzNygaBrNzFpndjNXYts2cV
nFDtTEq7rsrE+7LODFVbNgEMZmtffm/9IgF9lKdhPMJpnY1R2wNdwicD41VdCRff
/24aQdHgkqAIXa3b0DmBXtoAbykHiyCFUMiBKYiXQ9lopc5myJFMi6xsRJnjIvXj
93p+WG87HutlwLy73XS3K/oFHZBnAbcfocn8tQiQ24X0/JlxlO6H9u3GRpqXPoIh
WUW1l/wtOSyKTyKIbbBMmOnffqFZVK0SWux4aAsHQFRFAwf54SGR9b5SoEf1BkZy
OiAAY78H0Pxizng5qU+4ZlcHuCJpVxOaTr8MIZ5YJnay3Y5Z8meG/EqxPEFiKCIO
BQuUEdqsooPexHHoKXO2kx63QNo6RhxHSkFeiLSid3JEkvBH1pKtS72i5oQ2I3b3
z3GF6Q6ckXx6rqAI/LqIuBHb9rByVdzGilBtWI7fgnreNP5nUfKnwH8Lb9ywVKyf
4p/0WSAsWy4vuNyQbL/mTsVEfE4IRjUbwrRrkaWDyYs2tMRGSvPR4hp/gVJLQiaM
OoQKDqXZsOGtib6c4H4HWMFDTXAPsNlfSKorSCNmcYZZgC/V3TbYKF6YCRSsJvP3
22MpsTh/xyRkH9r5AUD/lTNUS5sAqIPqm4Lue/2fdufANZ/rrtOuJ5SQR/UfYzG3
OgEQfj/DmV46CtqerzDZUy22sswTLbwoABA7+utTJu8Xqe7UrNyZ6eIl8zP1ASwE
oE7awlYX2/bV4HO33zyzx9K6nLYgFyYbPx92rTWx1go3qxfi26P5inJrB78Rh64l
ZoWRn/VJLn25PepU9Yt+ZWhy015BJj1ysRKA/xnsrseDUvIc+M3ESVdWY2PX2L6y
GD/g3lDCkSN5MgQW4M82ZDQxtGUaOmOJf7SPWXVzwPP+qLuR4qKCwhIaFX+cmP30
ctiCWuxywYkZzmsEUVk7P7sDuGYvgx2VvxbxIKFvlWBakMz3sbzNIAIe12Xyor6j
clz+eDGrvTJ/FKUfC24wMjWTo8ddKfmQ7zoaGV+KLe4l7mdb2eRWoR5Trj1VD+gy
CT1H75X3Dd0df+IoGdLYcs1a7Af1t1suz0KnaoHuup4jt5FG24u0vNgIXleZpAGl
ElEoQXdjUt273YWrvz4lwupcLNI9eBrNTXRQkVgRIeB35yQ8WCkQR30zlID3x7P3
7P9XMEDzjw6utOmfyG23ahlKKV9VVuClAC7R4lzmy03Gj+7Nlr2tMKjTjeyKXJOF
cb1jwxqQ0zlSuq06s11d+kQ6d/1hv9KZcKUeHxLh9H/SMsNPoGRkCUGCdq/VAK6g
LTatFp4MI+gTNw9u1+6G4XjemkmCNmliO5UeBhMRN+ryq2fnZ0ksEgl6/QO6L5Re
OEBLjJ4pUFk896bam4ypcwp22SY3OZHg1uipW1dn0sfYu5182qOT8efBNU7vdr7T
ZDDHDl3T1hn6j9toyKghX9GhOYcxmnaq3mr7a8dUUFiKUedWRw6zJdhNE4Q+G2BM
aUJryK/bLfpO3+3XTUEoraOrnpOjlSplgo+X2MtPI0SPDe7OPPPwpzcQvJ7JVk0P
omAIFzUR2rUqwvJukfSMzkcAUUKijaPUQ7P2f5i+7vIC3uUw/VkeynFrFvmm+2ou
dtxvnEDc1t2VHpJpO7e8ntL/CNLZSUt9fa6kFyMSjxZvcrND1Bex87RAqon9BLme
coUlxTFmGhMkuiFPmfHowQNGG2ONZ6zBG3UEyBqNijxgdw1YAU+nuhA2jGRc5AAA
SFDntMh1nzRkoNzA+GZuLQPRKqFpQLjVEvgJ2HT45+huJovjvWD0EzF60NirGIpE
8jZVHdQxhwbc3dIll8mdk0ZUiUqTH7jK8XruEpZPCS7afOMaZXHA63YQzx2Fn+fn
Rd5oUk85vVxywtpUCzOIOymB1A2N+fTPrSElWIsdhXLSDZU1fM25y6H05UofTft/
FahIetOhoI8HRC7gKEJkt9Dd2uohhxY6hCFk6TdTERc2XZ6mlwgkvlwYDmH9tVoA
xcnOLXO7YmCA0EXRMmz7SyHWPOeFZBALTYPwxYuD+CaI1AvURsYPjdzXC72r5OA3
FedKUeQGtv+st97AJ7Xax8/D+Fx1Y7as5K1dvVkZHd1ZvJMZQGVULcBBsHKyQgWg
w6xQF3z0olUHWvZC1O77EUwjoLfnQOh2L87Rd9hUYPYVyEENaVJ+uvplYvuLWjLr
n2A5MKv03lM8m8zi8Fhz/LvEWumpy0ltluO1EDxRT1XrhKStKjrKscj2MMwqPjH3
aaaep+x2qsM4vPxuuu2Za2axgtAC+H3W7jOohFjCB0Idv5dEN9WbE2QMjApqdT+R
C4nhUQ0BNM81jYgRSMzsH/kJx2rMG6e+fD8/BHjXE6POPbV2DQtbnFI8yTqiw53u
lMLR8TaabOW/VX2mQf1WCCkAyJYaQIMJi7LS0mOeQYp1CA/BG8gf8iDDfc/aBjXN
jeo+AEydCR/hVuNcNXRZ95TKN86YdMJvSqH8scw5AaVoXwXNoS4sYQ1weCAG2iVs
vkYjZCo8xIjtG4a08Hi3EkNWp5HgLXpgYHqi29B+pz6tDekeMXerGi1fmsQkK5WE
IYzcR5ClSQYgGLaoYiJvGMcgyebNDjfhKuyuW50Z5YVmjhbpbx9qf51vv4UnONza
Nxn2iwqVXIjhdFzseK4wSwUqIb1+uic6/OKkHeAkbIsN1F5sbSdA18aAZ4BfAMnL
EsxX+AolhEBBXxB9o+ck4wsnMy69//3PHZrEZMgxRTIskbdIqxY3IUVPu7+QSwzl
rmHmirjSRwudMuNKn4Ps3PAK8bUSqDV4pPllMVTJoans0NljEkPNug0dPljCZTR6
jEKqzkhbBT3qM0D2z9OHxONH9v2fxJY4Xm/t1SqTiN8zw9SyvuOVW9CwgwiDkX1A
PrrwdPlpxJeaqGgQnbbOMlBpB2z/+w1HQbu//ZyJHRd0Eyuza8PYPXrVGaGjbvjg
XtwxucOSdNB7yHbiaooQR3AtYKkR4wQLom0tOHCrACh2K2yQwfylIvIUCa5JWAE1
ERdut782CifIXiMyWdCF98CjJonrtpm8Pf4X/cfXFpFqhnZqOi8PyHXEGGDx7Mcr
IydcjosE4LfKTaR68vySm1x/BQnNKtogB0r+vfuQOC1PF4PA5ZR7wPrcnXgWFDaq
OB6SeXeHpfDlD8zUULcVOzFd3e7lYHn/8CWwGWupgOOb2gDgZR/cx1BxhPWzYEco
tuRxN2Ob0mjilrFZE8AoxwnQ0nB3L+SHWwujoD43xBcFEiPFYxTNE2cVzKIRdb2U
5ccBw3vujbeqHXjXshB5zinyCnPd7nIJWgQMHIZ42qBmxNfBYiAYw7BmZeFCTYeI
F4vFMcFGWnUlhkLyS7dC49wIP8ikISTYYc8wo8XbJmsBI4/+oXmC3Vefx1gPhBRV
dyS8XejzwsvMBT8rG1oy1QmtVrdrERm/GjGH22gAXxARtMP57FeH9tm++8ENrLhe
skqrfpYG6N+0CQcZHxIyNMWdvQtUKt1AJv9LSLz8hLGAIXtAnGU+et5MODY2uzXf
9ikmIhnDkC37i1Fw5ZFCkogkrxYUuCk5rr58jV4PVOBma1yccHlJMA+b5gi0f3OT
Cf4j1OTNkuFaisn9mvY89UirwxSepW/dr6G28ykuOtmC+N+HPkZGSEpwLDoFCaPu
XftMD8PmF+xFIanEbvk5doFOW0eheUiMpP7IujRo9VUklNPd2kjckcWmsCNoNyIu
x2i90Lcw3axFJMKBkO11SZF1FacEU7yqBxQHYBJaij7ZLFM0On2b2EGu19MIW4Xb
ADF5oSiGrXXWiAs2uCjoyNi0WE6EfoK9AgUI9RoWAdl7AZhiVayzq0EQTR1YczMk
hLYlipU78og3pjcH7Jc8vdk1Ma7wi1eCy1ZP/p2T4TWcApQ5O9YDqKIAcBRCLwkd
3hGwDvSTukDSxp6K0RVyEhdpvo+WeDujGlE42jfX2zKGBFuGgV+5W5XnzsmOxyMS
LrAiSW96yFu10Z0h5r1PXqC+XCSaWiGBWzDMhJLEnmsr/K8pAsGhNCH2O1MwZbh0
U9qVHH3fgnk5vDJsClNGRMpqOa3In//N22E2f1ZzWgpMR0N0v9rCuCjseSsemC7i
26+GNimQJoLMVsUoCiG5V/KsXXU4FlJejIcIPY+RMGZHO05wkttg8eLXfP5+x/3r
8ZOeYbqiIAz2yQoIaPIvpoA3rW7pN3D+uJlSf50gVKILwL0xzU3feYIjvuOwvS9K
EyzQUWbTXJXZb0jG2A8AnIyTVDNZaaZBpJ2sGtLK53JVkMvJezYzEMNVsPbXqljP
Yp5huVaAxmg149zUt8F3VuhFLdhJqFSY1pdwJm1cZDK5+/tvFzQVoA1KjIovXv7+
O4Wn/XKFHjLMWOMDhvMJbCfJzmWzG5CCfK/oQtXr3kfZS1/hEaa/9zZ5mUvcdOUG
wkvCa6/tLkMPiTcS3B6Ckge64LKXPAUywwBFfqdH3t3DzeYKgsd16NTWImGeIBQ8
3qS9Az/uLEC8mz+dhHeJJ5/puAOOna0EOL79slasbk8cobgLY+p9cYkob/nsCsIJ
gggw+qUWYShUDjE4dp3NuXKELaZ8b3UzDol7bxathsfkUmBt4spmzob+Me3pwLjQ
qm0QHvTahFhK0OKjjeu92fdxE5RxpMF/+SnqWxjRfjN6cf/h5tInZdRvAlXQnY/q
mA8e4d6DmEF25uPMOcfiYUZ+QT+YWEeEhO0JE3CprBwGbgxyDIiBp9Qh3eRv6TCa
C210vp3LTqago3f4/j32MqB1s2ZAQ9nCGDc6aZE5ycokee6uNix6KESzM1do0ELI
Ob9fvNhXr5xW6bgAUyK7VEPwsvPYg+Lu/cO0wE7kgNKei08THOeTwaQPq7bN6Peg
fZPgYZjgcg0+Xvg1dapaik0LyRrxDiMdocx31M0fXtTEqaqb2ctW1EfKieNS8EfQ
BW1YFLCO9MwZ4cIrGvPa6G6mCD7sVfFfQ78anh9BRBLtmGRyX48+lnPqliw/dA+W
VHQ4svn6tUoinLyJ5aPKaQmgGqPN5i/Ru6g2QypB64yVkwtg9UZ3+LzdjgntiV2B
dH4S7X0EPVRhmScZLPzgmJiB2THm0OKRM3pqCHvWO9wgJz0eC7+07hPpy7yv0688
OJWm6FUwXZjdIeBl9i9njrFk4Ffpm7DDv7gJINIy/ds6V8AdYsO95Kdk0Y27Y1MG
lq/P6G2Q4CjemWUl0SptZUj2hzcOge7ZOvYJzi7gTAKJrcIcXI5M1L1pLnGMhh8W
0idaPdTlHBbiY3DbA2SDrVcjGh4rMkV6K3Dy3zh4HU4PF2vtISvJpWdiWkzpoUKG
YbggjvfTtDRp0lF1nnotn3RQI8GiQdEvUb3O+/oaNj3h6K/jcFs3P5bSPI8AjLjf
La+64AiN4unmQzUQ/BXOmYjvc5ic8lkqZXF00CCS6UByPrDVnJmli0AfRYtn/9u1
JG2od/msNZ5FswtcHbEKN1a5YghHxHTeiYW8ZhnF0T1AviwutQqJoJRgI0kBiqS+
r0LRhUcHkg3IqBQiHN/3nVvmJPzMT+uaAsv9tWl3Eh2cHbVqFU3vszT7NX7ue3ic
feFyRmzp8xklPttA9tWbIs6iASKKzgEQTouuKabhHe77ckpzPCWYKCn5lov0yzJC
TevqHayiX/Vg3qBCKaD4DrOt+phw0HsYrtqy8K3wFdPSbk/6vHkLAgOzrE42TiqX
Ileay3NmE/GT5OosKk0Q7Xt2TtX1xq0SNmphs3zUpGEipqgiSpLGku6XgY/3PDzn
Y0tdziYqSAlKE5OUCQ+FyxbzYMVLMXg24LbdxnK7nLcrdwSsoAhzmWt3oEaKydEt
j9AvQ+SNjpkZhVa9sLvKv2YFv+n3n+Ldq+V0Eq+f+r80o3/af77fCxgZrBnUmrL7
1Oz6O20mxFQM4EX7UGYCkEJmqNs1gmQ3JTNwJmCj4nD5ifNkhWnQibzOmfj9nt8q
iem2snfW1me53AtW3kFfJwt6z9AzgSFxfRrMc+pJYBZOxFIaPQ97pR41P9Es0Z9p
EPfo4sbvD1ZZ8eakdwksjCkPG+j+gnTHvE0DUNwqBcoT4q8osYkyM5JlXXWYDRfz
pHkfg6brQ3qEeDVSos9sFB4+5SESK6bZQ1dNLg3Ps3E7AT6G29IeS+XyEyWgtvEU
C5JJ6qy4vEdtAftnDgpfJELbrlG4S3RbvhzIZ8OXhmQbrlOi2VX2sPUljCQgOdZZ
rn/snuX2elL+aNbbSlIb6eN6gMjOkSBSDZqRZ+N3UF64DPSU79Rb4FUPqm2uLbrq
6z3mSMxOjCFMorn/1RfxYYiSuT/e24D1AX/vXXNEigFW6tTgvHV8S7SqcBWD1u/H
0GTQ0ac1Pzf1CpIGH8lctfm6x3sSrs9GZEhLXAUhK9/1sCt5zJZ0nubOix3tYf3e
lt+ZYKW7gH9UKDF+1XbppvF9bdtfL83F37EMSfpXgiA9pZDqUI6Mvn4e578LkEeo
sCaaSYzyyOvkj1hAMbLwlnvhFL6V8AnCnQE0sldOsapLJB71CnfV39YkeEBEBrqH
/xgLYfL1ahIp64iYy69SN0xt9jBhpnhcJth1qZo9FwhR2Ri2C4YQkQuXWPABXuAS
rKBJHIz0NIkMwT0rbsIbhX+d5vGHKLo1HhwwhURN8fcbvV9tkwIg+piAY0buNtYg
Muvm2o8HX+hVMkrGywfumHTcv4nUQ+2aj9iaYylcfunYiXFUioLbKYvTNx45rFD2
/aGktXqO4XF3ahEhEIcHR7mYAiMEiXgUOpRJzchvqLTAGN3+j6lCiGXodezCdL8I
NrF5xqFD989oOyk+draoEz816+81A/4E8roGs5Vi/DZr9oeUPTI5Rar8Q9pFhaaC
vZdJ0X6I9RTE0P2lZc8pZWIXgRagmBk4rzO27T4eJ3yEc1/Nazaf+RmY0O6+q01e
69549XxR52K0UdFbKiew1zRea+Z37nY0YmkHVuRjMh4z1l0BLGU0XqgeGBreoSMA
vGS3zHuQo5AILqvwHMJsiUJ6fI5QeKCrlv82d4OtV7hyXXXEDI0ZANtNNSGC8/JW
lFKpSL+Mc6g6CWimEGViho6+F0qBmkGlfssJFzr8cQB9WT+uKdC3GbwCYnI0cEnQ
xMVNVQ8an0HfyjwIB/+dG8jnuVm4fuDrYmQD+lXZZq96BSEznbKgHMzUaIIWRwip
GiX1TPCROYqHG5kDVeYpw8Ci0zTKPkwprFdRa8Ao7qj9ykg+2XA48XvP5/SPFkNO
zpdgpFsWJZF/JZ/Pcjvg2maUASunC3EtvnwaNF6bussa0Do3P/yZp9wAe9dUglJI
+zoZ3KLiXYxVzB+D7P42bHUGl5KQlKBjugzgef7ls2Cnp+5GmBwaRsYVTP7V5bII
rhDKpXTT7/piFyhaYGFIsVPEsns+w6C/8ZenS948DIw22V2gclpLr5iZYuEDKszz
44dX2gZ0JPxY8gzxrfIMgmTdT7T4uCL6LkuKoSdGIeXWsZKhZA+kCOcTVkUzmPWX
ueCR/zdPwR5BS4TlWUaeNMGfp0NVoNOo9nNZ1PxuLgPNZMBRH6qSQVGk/9ZhmDLr
DJdWUNvTslAfojzBIL7UyrO+TA6ClvPAj+Laxb9S+mpJkzySS8/ROpX2zbmxWR7N
0Xo94F1Oibxrs+CQQ9qvxN06eg5ku7SppbJziw4GfHRXoc+bVcJMN+2lSpn3f4sA
I6806a5tGg6D/KlwQccFg+wjDYXSo1n/HTOSB1hkA3eeHPjJ3FWvYIda/LQaNtvO
lrxysIViJltAqRtVHDwBIy5pASdN/Gnyw9QUzGgMFarxd+XeLoqt5s7TpkrpgOzf
38TOh7oiGdLx+bh0Lu6vdaqjM/I2MvczugU29S36NzrTYA4DDKsUjSsyUmKkdLru
jKxg8KP6bh4UBIUpO7rs03UVvp55zdb8OlIDojGjN5SetgnaWE1mxufGi0yRowg7
9I4L95c9vFKd8cuypa45t/kXtk7l1ejpEyAubg8hQPNuvVQgnqGZ490YlIBIg1Wp
dTQ2VEe6ewqzlsPummtqweMM3YUEm9g3GRSUdaCml5fUQv2eob3qhAlzo2mjMCm3
IWoHpxiT0xJKwe5QEPtrK6drDO2yXgrSSL4BLoK1YWSsVfIRUoIV3rtfq+V/oEtS
hROCYPA1eEUdR+PF54cKcwm3vpGKNP+gcSC70eE97siGARVzNfDywwjkdiHQmlMx
Ht3GD4VzRnI0FmUzPbHZVlm/0f8+8lXitBF41PBdpRL84tactxH8h3AAKOQr6oCz
1wRFC28UzV88M3P+DlYByLP3yfm/34W1M+051cbwY9m60WC4BhsKpkLcMMwCtbe/
G3p7tUloUD5+zyb3P6gzSpbiCCvU+s+DWOEtydxl47LUXc2u1RjzC9dH0rNbm7K8
J6+icCmODGUP3QsXiFHkgLw0mR+wFVP6oFW3f2jA9RD+16pkpfBxTxMzdnLLcQkj
WlP+d2TbYqMqNG2jJJhRNkTlSwHCsKRp0Nr8bLmu4ep1KLLuybukgdUGeKc2gp5K
EZylz8ObPOBx1TVgTUd1oQ500Jyl+v1b6fJDpD3Pclm7D/stVoCPQ8iDYSQFqQ6T
NZYPWaroDe1wX8hoHOH/LDh7pljwvlkx4WNVwmTK9sj/B2iWv1eKMnwWSgFdzzQG
n7N5NkoYW7TKBPXjC1yi0g38xkNCUfOGz6+39VRwsLfEiynSF6NnTptBKtAFj0qx
7ES4sW19pJgHyM22i9w/y7oJC1D3Ss7yeqPsXoauoql5lRxnWJfT8aB2h0cX6f16
ZNBCQn3gOkDZfc5BqBEE8VCe3oYilQQb4b54qw4ttAPzHLrjjzEjjLxd59Q4FVsD
uE9hk1MtKVe3CwknBOV9IaKNak6mkJB/Uo41LdRnsSJK3kxOWJrfUsDWlA25xc/I
kX0yLWR5y7RUu0peo+sJBiCToXvj+y6Hw737ns7+QLct1D2Cb2P68a3bFpo3IioA
5mUZhv7XWcjrq18coTKIB1bVHh/RTc36tfa9IoaQUMqnQV9U73Cb7X4D/B6ljZt0
O2rBSEubt9YppF3LjoDpAJfs20qCK9NssWEwUxN7rew/n5uA1XxoHZ8PZHXXbjiC
sTtCsczE8wQkJb93YOBd+neT6fMu8X+ZNTAc71DHyYXRcbF4uaX5hYpLqCEMQqJs
7EaqRxU3KE/NGd8h6ck/pt+ARbekmiKG2673JugVng5PMKAQmkygTFzMaUxIpYZT
r80TXFxtJ9p9O9Jh42bf3D1T0dyIH38TpJ42PN+TVggxIdFfZy8u5pId43MQNvI9
kEDoxiOKs2iFB0C9fkNxaISH3wCmzRu1YEoasq9fEC5v9taD3v6mGEbTCocOXW0G
zMP7krdqsPzP/B8WbUwxFh9L+ol84EvGTMUlLC+zneKSwqNCj/qEX3cfuLcbkiG+
v6HhmScxvJnJvaxgQq3cZvxuWARODzi9lfRtExYgFaBXLqZ43PhCRa+51KYxWo5f
CIe7KdtOiQUD3QgHWpEM4V4SmnPrC6rbHYhKE+VPCG0M7c11P9s+ujUjvTjb3cor
GfDMkZpbwxCCWtRPxkvzFoBpcQ2N4mRZxyFY5k5IbvhJDTAQh4m5lB1H8e5BnXXX
VIwN49pv4vQ/P0UBgmvDupWkgt4GHiLIXggHRVWuO/NAXm/+zgGkAb+3BOz/qcRU
R0jgHBYSS1ix7sVzch5Q3afOIYtZ3hxt17rtrMfKScVRrs9ae7CfAHu99NLTCM7B
IAgaV8hkrHHbhZnxA6wUB4Z0UJrYs3jDYvYSiTewmxu//pjuVzCqbZPGgkulQulT
WcSXPJvJg2EFxvyLX90Ail/Izk70BgyFYlRVgcwh5TVwTchTMb2NTcA/hY8xk6bL
YJDupbG6ePPVjLCvCgWdpbhhOBrDO2gsQz/+UIdTP76K5hD8G+w+uXp1VRqTa8hJ
It2HXOMUWIhMPsH2ksXkjZh/Meo8NKOC6TghIf7riWIQhyPz4bBwnQdSSbdymre8
YWZSBGnLfnHlrtINGdcScNC5PciPMR8au60QB5Fh0pbUfDn3rJn+cy4KYBHBReYn
1uCX0xvM8VJLR33DGVsekT5wFxi4PeIOYDvyWFaFwnZfRb6eoVWKC0MRy5kenMLK
X1R9sk1xcoIswQWCBAZrmh8n8KAndrDhxsQc4WtW8gIHOOBnxo5KtZTT9lbFu2pE
4RHbZjtkQj4L8CKPD2ofCY/txepn+mLLNECGIms0ptHQm4Oigs/7t8ypFbrUBv52
57zzYcCTTa5l/a5+ksRBUmm6Waj4jvdm4LzzNL44Xz57w2PF2sdGXE9It+2ezcz3
ghEKjHgMY8a7sjSO1JEUOXA7QE4ERoU9cLkcaLgmFVFzZywpaxcVmQgsNnSIksP5
oVpewHF05GJJPgKGycCOgbOixModzJ4mSTwlhSmoKZ2J5fxtHos7xONl5FMvycB5
7fzUJwgTphSZ64+MsqPndaJZWOQTwKwRRu6icdVFMAnp3hvMS3q9pV/1NUBRn1Lj
ZWF6u1OoY6fDoi18XA+hRHO1D2H2vvt80ZL6AXiK1ih8ajR0U38mwcr2cf8yBeiY
0MirpaewUa/Q6HwZMQoTWftvyzx3Y0PnNQCJY9KHp8lEKbCju324xXqTgv5JKCnx
i+VqDeTTNZgihK7X2Et5qtjWFxpJQlN4ATOoGS+RRKjF2uAlW2rb05hYJdDMWTWo
nLihZlKUgFATLa8UC7/g0CuHfWYehWxKHw4nhKZXdT5iIM9NgUAhCR6k13a/53Kv
hc81bvGyqT4UM8XD+xdjLIvqmIvnaSfue3mQfeAotl+askPpzWcyoBHt9gp414h6
RXQBo8CDofJU+WciUqlcWgMBCduYtaGlmEnrnDKecQQjxO0+nlyd7sYeLklG+z0i
4usiFns1t0R9VLXOHRv4yZZYxxWZIUshMqvTg1t4Y3HM8ciPe275e8N2T+++niJQ
CoKOUL31ylg2YpFcQ1jWLm7r19oPsD+0CORK+FMWwTy+DhHiI7cdVItiV3GjcyhH
nCWVJxIWjeYwHi13Jay43eTt6Xx8oVyVJTJl4vVFBpmOEBpt2ol5IM6DpFleWEPk
o4vhivSYaBY/yAvoJ2IOvIwnQfCHRRXkVikEZ9dn9GTY8jLoV7l2SLElYjQiI/mA
O7mhV7ZjEqn6o8bLdzeOA/eNF5R2HMpR4e4w8PxUmHX6g/N6qcbmgaXoAVKco4y+
s3fttHAS+ONkfe0jbh1mlMzlSLibDaBodaDZ4pwA1n+llp1oVC9nIaKWf2M/1kKQ
Nvs0Gkarb+4ZrfWoGFwWG8XP2zBqcUJKqBB1ku7YHpcm4gund7wceZu3jWIuEomN
0zjtDKojPkZYiMBAg9MOOM5L92LjDSHVVR+z/IRZjBM7d4CqN0i/FyXvSy4j/tLP
0NANMlhn5j1c9fIkQ0zyFVjTVACYWXTN0fg00idGCr9AazLmbb9Y5Q2kvlhzueEO
xDuOSMYwWNqCQ1asg6lLqIYD6wIM2f02zPSnlHGQQaxT1imxlUkwHueZVa5Yogbe
qf1REhLX68wwJAFAeD1T7TGXZb918Kn8iRpMAwsXStG8yrEDapsTzC6Hthpkag5N
N7PGAsYip47H0Zo7s5ADzNZP+aZd8ZYnV4ZJ8SLex4HuwT/luGWbIPCe+ewgM99P
xDQl7R+jTuha8I7agXslCG2L5k7miOgPtVf5QkavN4uJEyCSipeuujjOAEw32t/5
Uq/FjgRJfJhuJJs5iLvvEdLJmjSaeU2p+4+8XiiWUqaM3kufSo0vtaiUIMbWYWaV
mdOqywdG3/eCiyHLgUEx5frUxr05MsndEumAwtzC7UX9/dh+eem1Dm2XB1xS1Mwo
CCEyAxo05oMra4ERyotyF4JAnADv/SiH/R8puzt9mfQv/wlhy99EYfCIZZz3L+4z
Q1mN+m7czu3gd1t/XuR1WtHJPv9lAjOcz34xo8v7xte2FLBCruZQj+QKONyKb5hp
Ny1SoDo5lewNmAU8KoRCVkVJ8EIKZT0jAKjxMHo4CD8hvB3NMzfnFAbv/ZsHcAR2
oWn4vns4/us2ZtnLbRR3e9PilPYJm6/vC7VuNGQEkFfFSOQxJ9AJvvzhjp3nd1fJ
fOZ6sGYf0pNzdVFA5sHOmArkaoorB4CVg1RYKqiOUnv6K3RN4bU4w0qBSlRnmFsW
6m1wKK+veQRUwmzBsvMsq66dy9GPjGcaFXNUQRE0yeaBHOFX99bPjrkeNZU1UNIp
4p1DQnRZt4hZ3wCLravrJQyShUrhyLVjp8m5TqJhBJbqbchcYoLTPbjDDLPc7EbS
iuQhJWuKbKMLOL1AqCfSBJym04l3832k59kUuxojVUhqVukCqNht+ElkIqOYjJk7
R6YNGteYtyzq4PD24AJhwPzJHbTexl+V6gsyctHF7JOG9h/M6ZzsIueVv/g0Adf0
A0EjT0CuTfPayP38XZM0VFezyuU6s02WVuIhLfOdDT4Rrw49l8u3qv7VQfI49/Wk
ssJF+p/Y7Gx5HAuw1lLeyBOyHWUxWRnDYB7UCk8UnCTN1QAmyHPdDQKMOCQ09kov
vP2R4rfwTuQfKDOs6PbHEFHuBrV7SepHiI6PFX4BWnrm31hIQ1/qHW6sm8P1Wbal
HWKqLwm9Lxv8O3IKglULlh0uOZzWLT4qgBmr5aZAWCOJwf/5t93N9ir42TZugySV
a75ZV4ZotbwJPTJAUoWu8RgOi8zGaZqiMnE6sGqKCYbtGIhk2Ooe43ETN9kirsfS
upxX+Jk59WkliTTRzBgD1b5/h56oBPprTHK3MuBCpqcJEQob25IC/lkKAsfdCDOK
hfUo+Ydfxb1QH9DRIpbtI8rzg2u/it3lWXZVr0czND+ULl1Gh4w3pO3r5v6O9qbC
Z2835gVjS0+aYIjidIYPBsVpTCzpwUfqwZ7+R9HxgyLIevykXUG8tYXgY5KS/owM
Tqs0a2jwEVseQKgoqS8uEpi5xbinKZII9rkF4s5RZO1L3MYhJT3qI++10Ni7ZDbT
5KMVX6FCL7AF2f0NjKI0wGKg2zxwI8DHUwV89RBQqkBwRBr+mZzbxMqslG85dy8z
e0YqonWUUYu4qELJ4+eR7Pvof/N2vD5JNzE1jLuk5WAIMdi/fJatATf0Bs4oBFlv
88NNVb4gxCJ7AOJ+cdm3Fl+W7xRnOT4dimht1b1WF5oAwVy6eIqtqjuw6Z9UpyEl
l4CAQ+dRNwu6nSsUquh6hFwE6xBgAfFeiiiUhBLMqjxWBAhKSDbWW13lZaijSgpA
LjEape4/rFrVKCxN/ZSnfpgln7I5VCR2XeQl/+CNk0qY+X5m0U98dK4XIMY47dI1
STgaZX7oGhrLVMWaH8/lBDGIbTth+WyFzjrX3CcUidhYimKECFAXfpwfmwEjja6u
SD8U21KYZ2zuBGOoyplELECHaCbSXvZaE76WpWDz59DQBYAgKQfwCsoFbr8hzDje
w8iZ5505L+bieuo5DnvDp5kr6dbRdmPLN1dEOM2DbvA3+R2Zj2MbxZYpWL/eDIGw
UoO9S7JO3eG1WdA0siOZG07Wg+Mfs8dWH3JjkUSo7S07m1JUEkQ0Gt+RehvU+OrZ
rAflifBBFIwk5xR39tMzeAwVe8SGmvPT6XD5mMkK3N/kRqFzthM1Ey0fa1y1PFgg
zPfB+dRPg0p8vaKfe2TPpN+1yriSRDzCcMx7az5VwaP30ppMj3CFoLoPdJsM2oI0
/U5KImbgzvn5XQfbuOQ0c1bztFz+UH6g6ngOntDzGSmz5YB6CfRr1vwwb3b9ofao
eUBgKo8f3t/kxfvOrsiM9UMWsefbRESMi1Id4QFAVBIM7jasS5fYWQoHAg5t5K4L
g/guB9hIHG7oayTtEJlQVzJcOilVSZHhrxzdQOWSLf3ZnKS2IRyQsMclpJ+HFuo8
US1rPYMmBLRDa+kpk2rpIHIorqVlCR1SldzPP5Qw1zM8fb4eZH67toD9npKrFWN/
Eby2QSTiU9L+Mtr+hKdjFcbk+tc0pWb3cGKV372RI5vlplc8GAhH+8P/a3pSDGpv
roYR3FHSQ1KKjQ6ctAz0Ch3ATvlmq9/zOlEINctZkcR080HmOoJTYOth60p09Oiy
Q0WR/0/3RULFn2FxRtceDC6W5cfVnfV+G25grn446R6or2XumPsTk3voOdXMWop0
Jq9zAkgicJRFL1lSqrsbMojyyoEH/lc8v5gQUDS5HOgg3hyVa5Rm77WLIAAUV3My
FTU/1CY4ORNX+qDbe5ATA8TWP5oSdHerf2iPzStbkwemTq7pQH8/XM6DtCBOXWyx
RgAA84ek0uI/5usv/ww61MJd98J6+CUuIuh/59j+dihDAMSNZDNuPgn6zGVLyqc0
OzQ/kLcJe4diSitMeuwWd8ka9JGJ033DMud4+d2qkRVP1EAnOXNXo/CVpu2xFGbt
J+hQEP/lJmoQplJ7+PaZ9/XozHeZ4oD6wFgNYAUmDTudmDjjm/5Ck/Z5E6JWFjhr
ojwG5iNm2aLn4b5wJYDv7Buq1m57K+qdaHS2m6F3jVW/HCDtw/smPu7unZao3XWD
K94JLRC6jZpNGa9n184/elXpA7zeGqYcps/j9r1y55WKdO+iSPZUs9yfj9p+JtFo
luhLRQHNiWVZ63rpyES6Xxxal8k2NEImCzHEgRZm5D7dVU/Q4SFqdN6AQgYTDh4l
0ZJ3Dn16GKiG2M0JbPpPSCudIJlbvxuMQiqSXMMbiZLOc0b49FCqbJyIc9vJuLqi
l0mpQIu9SRAq+3X7UMxjdhW2NnPXpkrPMqMXkhK6nl9lDmJxJ3lc+yUg3c3r+whx
E8xf1k3qoNYJIehDhbSiO39lie8DJlUzvsPxXWq5avdNRk5bhh84jfKiTH87md7F
MDFTxiJRzlslQuOJ/N34eOesKfdta+kU29dxHa4dUo05sWPAFn8swDBl3hXI5YIh
IuxGHJ8/WlCPfvgTB3+hTTVuTTmTbT13pEpo2vsAHjqT8AuI4uGwkPFSX2g3t1qb
/Ze3i6DJ8kkNleNf+r48mmiWUe9iBnoPPOXF637E9YFfK8Z5vXklLjv8CZFrZJqJ
/FJ0SIc0H209vFsVVX6rXHSHNYhMd97JJqtqLO6Yk1Kn1nLd/M3z/93/LRSR0vk3
hR14Wbr5bztY6AU7CDOoI4rc+UwXt0iJk5oF0U3QnnqSQHIv7eH0Z4nc6HzpG6Pf
DD3u6XY6ahwcWj+372ZsWu5/7kjm435RJudcJAKdf2c4uaJAK8nl2xYZZ97QmI3R
6KvmMW2+Ikt/XBqcxkBKGTsj3O4X98rpzyYNoe4u2LLIgTstX/V3fQuO5OK9/qt9
AsniSQr/Xm/yXM0JiiLA2xqXAUXvOOX3JsE4oaW9enk9tOC52T7iqaaPwwvPtzJS
ymnNPdrfzRV92AmqFqKIbwYpP0xtT61yJNjxsKp7UsVUXtkkEOFkhiCdRzmIecIn
YU2hw57A8n4ezZogzl8C+fIhUogBPij7p4rK2fJD1Q5mE/N/CzVhA874AMBBBAen
Kiiq2eV+r/PmiJjTZIcFAVx/D4DVZwbuDSsqokojpb+SYzhIrgVbPvM7rp9knGll
5aLT67HfvuhSffcpcT922Wg9JxVSTsXtS4xwD/t2q+rCwCcNAtX7vgokmZVWalqN
+YK1p0hWvZGPb04szeWKyendZuyeJIgmCo+rfUiwLWXlsMCsOPMT5Cj1creRS5G9
Cy0zlHpcpXqFf57tKFLJD9ZPjdVRpeqlXK9O0lCtkTbMYN9UNifQHKMkO+jFBAts
USzNDbymab24gERHcZVM5raDYonfqWIuKM2ZQBvo4g2li2pO4g2vOb7+hZWI+Qlg
BV8xJ1IaOAhUubNsbwSSwfv15kyJu+OAxBkJ7jOgf+zSh7nwB9EYev8b9+m+3iv7
1vdYsQNhd9WkMKkXeogQYgjDHlbgDrIG8b1dH2BHOhWMbWHURdI3kB+mtQk9vdhJ
IEN7Mc7/9wM3owrvuIEbse+N/QgQ5Jdp3S5aqjtytrc/35kCBtXqhg9qzg50eZIT
f/EpN5eNxkNGZWrTEVF4eVhmWQb1J83nhQynMZrmkenfgvyk0sLPAKWuPWbsYw2h
qwpULPCa6bud6ucG/TI1TDIiilggHHIfg4ZRewKOt+2DHaquegBHz9Eky+ehcnFE
SNeSnQKE4az1FF7w2rLJNMnXuOTxmeGaDi8P/dkS7r9h6sz2tlxSUJ/Qv3gS3i++
yby79hVceCm1PWlZMOHHXS/Azbtbsq+jC1JSHgL2tVuGLIGA+TR9CQV+gnOQmeTv
ipilPew/BUOU63k6K5frhs9UJkDxD7w0l5tMAle3DP5s7l/ie8go3mA00juEjmOk
18hCl1e9IwgjVe9t2luiCZ5s/82E2ZJNzVLlFDe+1QWSqU6DbSI7ahlvJ5t6ZPoK
KjW0yYDjaAohkoq/eoecuYzMdLpK/QMv8zqtrVmS37EK9bCokPWmcyAXYPVxL+Me
WXYi+Mm73VZqCEBuVJbVnocQgdHC/uiBvwPHGDtpTyXfJ6740k3DbdEBzOY81WC8
c8Qn1PrQrN+1oHspaRfz7O3vkQIaBlDnIxPrTQFwSVFch62eOA9OCj2cGyqRWE7l
NxLhNS83iPShk8+Ap/E3ZQhwugVsDIusWtijGdtX/5B3vs0NPKeqJ/uqNqub3K1R
7EauLrN0zY29KlBJeO5j0MXJI2TOBRlGQ+17ubxiaRAtZQYjjLvWP8+qvQk4Okt8
tCqOxqOkj0ZYo4qCuuYZVihOB212nUeEpaICSRqWEn+Jh6nc/dC/5L+MU2oJ7cc3
z1lviBXNNin3MMCruIhMlKksMRbg08YpgaSyr5bBnATNKOZSmSeZT9vPCxiKzs/5
ovXjT8V+QBNn9NCf9rMScjRYHUR3U1+LQQTXxKjJEmIpakm4GUZ1ICrDxmtMNpbZ
+ybu3C1IIrcl68G2ON9eTmsZBsLzO8t2nlo1QMa02+R2ydih7ttW1/1w5ErxMIGf
sHAZBDGO/h+kbuIaEOLXCXfMXer1X01I8+9MTnHX6Qz2+LvnCjCFxWkwCy8CPVu9
8o0eWgLdqdX3milCDEz9ZQvDMLtCbgCdxOeDY3S14mG+ZEmmeanJfSDFZTALPit5
eYNIIcux/DOS8UB/ETicD0Psyx+0xbNXZROzNw9cED3kKQCvnAs9ASqObn0RZlCl
g3gn0NhwM5tbK3SJ1RUOI6Cm30tqbEqs6C48OI/mQXqHCttLyHmYPlpldWmJeb+W
pSKxHvm4/lsgv4RDxuSc5sD8WxiynEe4lmQP0EyZ0OVs6DAMLr1oSEDnbiONqslS
ESkw/6Sc7zpbNbsq9baLlbWE2cvPu3Ou0GDfmcBODNAJoh/M6g71RfS+E/auC9HI
ht2XbmfqeYVybOh0fjICMDncHSI25m6XLGuCqg+y5Ruckuzdt9WK8/uhFvi55jPg
8407rBkz8ZAN0kfpLtLaKALp28SP1E0cgoB/mXEHjCkAefhGp8ujHqQOXV6muRwk
ZdIJdfLUWFdCWJEO56RQFGLFYsG9sauOqV8WmRCVmp4XU1qDx73jp3eAM6NwqLrK
dcH8ddmdz7INixue4aCaPGyIBdvtc9FNKd6hCZm/U8e3r5/wVvAGw4PzNJqwSihm
KEWY715pnc9ZxzFZmsZHpUM3Kjg0rpr1gmjJ9Tc1J1s6ES3vwnwVOWz+Y3l1/60d
wf2oUEZO2tJ8LN3sQDWwxlqPTtcaKBc2m2QfrwSo/edUXmP3AwKwUmXE4sX+OOv0
Si6MYWvt8Ck1MQC0zstwze6IPGWy+stovpMl2zmWY5axHNOFp4gfMciuRN/Mtxnv
UcqTa9CLWoieGRLfoM5F4nqis3d2GuaFAOYg4VH0uRoeOWJv5uvmts4JZkuQjUfZ
e2Wj99n9gB2xcUZFG7zrpJJKN7K8kw9jNm6a0Yf9yL2vSb8SPFhy8I7v3XeH8wqR
MJ09Bo7/y1T3j2HcnBZetaEAiKNcVYOGnKwH3mZamil/yV8Xl6Z+cRacxwchLlAh
yRI/gbubRb/EIh8svnrL2KcuGseC38r+86v6IKUSvBk/Y/JMvm9JCkpBEv19Ove6
8C/1Q8C9gVwxdZcO8niSoAKanLzrK47VuyMpQEGsahimNxpi3KvJyvQZUGULQzM+
sGIzdg61DVoeJ+rO3woUp6wN9jN7RAaNMjoAyN9UhULS4uB62KaqtZPo2e4XRC5Q
ePxmn+H4TN9kthFpGHEZnoonCRdut2D9rgwLEITl2M53RE2TQZao9HTJlL5fg2BG
Kv5hKaCc7zbWg4fevx+pn4WXHRfasc7iM2TFDIHVpe7K+PK4CRzVX3yadN2jJO61
VmoyfnhnPZgRiCZb9nbFG2yz3vKj/Rcyh+SrW+GKGlhfV9Dz+abxFuQbXATmOeEC
3/2ir9n0NNxy+tjT/JEFs9AvQ2IcVto3hFHIbn2ZnBciFJN/ed23WXn2M7HkrSUD
DiwxoYSURfBVFQVf1sF/ivBFYSOw+bec93cdMMORoqtBURCQAOhiCEYK0ugYe6Xp
HGNSmwGHvA/nMohNwGrq7PJBqTK/i/ez2zRJlOEW3zBFUyx+5xCZxaw+svgptWiz
kji/VzPIiLxfKrDMaDnqzZDKDRcQ6gTcG4E3TZqb/eqdimMwzZRhtj2BkxNwfT3H
2iP14q/Kv+As+toXVLzTo9es44dYLU4N9FXX4h7T67hRQ3NZYVR3j0OyL71ommTY
VPEYDWKwm1uWe0iZlDmXqPwVzIcyGyix3SF1e4SVR9Lq0qG70H4lZvUAb/qyrISP
kvOSU5OeibgVxxp8RfnRFMWEmG84oTQLNNKu9lj5qmw8F3k6WnmCTdDZEcfanTXb
sjpy4ejKTV8iAP9TAVgOXWfYtFiJMGLn40EPWIzJ0R944R5FXoY7y7vqKBkF1X4O
TszzHx40z1SjhiF+vwY+951u10++bBJWH08c9YYuPoEyyW3crRomSzA+ilv3gJ9B
cr2OU7NFTvjcjFpD1LVfDTEJzaz9fO31hKKcdZfHhAblOi/rupYG5FTI+E5X+rzv
1HokDfZqJ0jtghmBA2fa/CTPeVU5CcDFWAn8bO990s7O3u6zKYyEFrlL+1m3EuoS
Qx7ZymIhWgPEXBdWIeVss3bZ0FlqFt4yDx0OiWeh+RRzxoFP4OHaxs/Pj+IToN/K
Dlaxb55f4b8q2/28tBqDu5JlHwAG7rc8JmteYVmd6fW4ureLDVmSPmiPfkndOkLk
fAcXUZ5J1aFp7i/CnPADQiZoJvqmhdAx6rmn//Uo1lSFKLaWuPwjvZsP9SxKintm
x5AgdQdrGDJntdvA/SyeU0NKjxlWfkVb6YyoDgn3JytSj6TeoII35XxcMRwPyd24
4ji62W+8IwO+sagYpPCh1WamC4ZmYC7oWpY9Hy5uodyY9SNM+mMw04cjyMt07hyt
vR893dCD3Y/fwPKJPgw5+/2GeyrlVuDEvgNjNMxsRElIy/1eKcIh8jJezh4BdzXW
2JmO4rxOCyW+Svn96Dk+iIfEFKgWDE1LFgmgsmsrrg0aLwJjD8Pk2h8kAdCGf0tc
Ig9R9Kikpb/uqTHojlO66pZ83WLlYjHkQ90aE7iSSLnGpSpxjHmV2+2DrDWdFh1C
fXeugD6HZS59F2I0n890df3qAbKFedoyBxeatCiSSTq5KOMHwUmQNCTcPofhanCh
ZkPIOgkS8WgblfRkcA2TbcMSKXZFJ5KG4L9d2b9zsmofj8jcqTCW+LLKgC6gR+Pa
nvDvwhgA0ni2MYKBp7hZ1VcTYWH2F7YM7qytn1uMo24084e+YPXhW2YwSEz4bsmS
ATQV44GA7/wEMM15EMuD2vPJnlLzq42z+JSt4pDa2iQREx9Bt9Vylor0lvlyuQYO
Yn2aiTBIFwzw7JZzmmAMXh4QqpOi+l/9KnZUU4YSOa8852EzhqALKh5HN497pdNF
z3ebZ+6RZV33kY/2QWYu7zoXZnYXBhc5PvDjYs62fQWg49W+1Vb1v7MYJ/fuFYh7
6iCtNnnpGi67RJeMKq1nWDK7PhZgWiMKqH/M7ievuMkgws2zb9doprFqlwFfjJRE
/ONh/86BSw6FrUhOYWZ/f8az2+ORioN7cWlrSU4LlzrpagEckeN1+45eHvi/g7xc
dIyDxlXynQo9ubU0Z9JniJ3p9kfhkpqTFb6nJYiZjb0XxvNQvUE9i6BTRMO3DXnT
jXK3rXNfoVoIHHSnE0gisuXN4OlgW+L+M/H0f2QvBtVdWLbz6Q0Mf0BSsHpY0crU
yTeHcdoCdJKr2CYfSNSDi8NgOMNh7r5sSvzXkxdJEuBdRR/ugyAQVFGpvLel9KUH
SP9dDnCcfwvAU13fgERh0HpS4GDu4YALc8O6saEZWl6uA/qGHB4doHFR8dLJXfQ2
q9PQ7FsBK9YBHYyJ8+TrnRK4fTw9/iA0DZEBMVGn/Q+IH1dA9+7L9o5jzawH8Nbp
0QsXbqQzT4UsbY6poXzJwlN2/muKR99JB9iInhdW3bgHo8c72hUywvFpenrdD1PF
QEV3Xa//WmmK3YodVb49UYZQnfOvzfn0bqkq5J5fxulw+1Vo49o6A3Os66olbNoH
nc1G1NO3LmDi4ADCIIMUxrEyA6dIjxGuwHLnPwqj8veLHXNH3zy6CUFvZJnABZ8w
hSU9bXtzCnkWmOkNg0M54bbyqbxU1YdFbUMHWz+owIl4u+QHOEmivp1AAGk+7FBp
nk8sfJ2UK7q1SMBRmL4Dqz7woq1w6VZs6IrVDKaZXOH/uVL0ccpupF2Eh5n7dqsw
3m4HXwbHbl1A1aRir/5E7TEx8itb7MeWCaG7URTgXpT/niAshO1hfL9qjVlfBuaI
fXmjis8VEgJY8bZKNmQiRSu077b5YnWBuyagPa6KfpowBYGMr0e+LhpNGLXzIrOp
cOdmlhEDoY4wVfDe1JfxpDW4rgOwJCfEm4b6ldDkq1KksYSfL05MV9uQ4Zc+1l0Z
wkLklP3OMrCkPC+ZfX/ro9+9r5xjyoFYynviYPzAi6Djn0t7T5D1eBNZCNPh3Q4C
PziN+0yaDzZsfo7vMygekuLoOVmzoKUMKY79YE9eZeXDOga7Z88tLsGk2yQFiy+A
62s44M968xgkPlTi2qD8hXy2TEne9RwO+3LHx87OpXTyaGAtRNshAJGzyXVnndWi
B+xK2KJYeAfTuAbTmodvZTLxJ1v6jygKStXPE3yMMg3jfiUL0QWVSAi002pROKb1
TzXgJ14Vw2Cs8HUxxsb1+1C2M3tXstcObuAMJoFCHQQkZxsEKJgGO/5vKGzNvRdR
5RXd7wjCtAt4piQtXTB4kLWOZcK0jI71Duis1sLAAi6y0XB5g1aObveHMRpi36Mc
dJb+PGAnlOuL8qDgbkc+4Oj8m8f2AdvKca6LAgMT/ZHUljDTWWzlRYSvUGaxI1Z+
6zlTmhTaqkJhQ1gDvyM0ThaiM4aSZun0aS24xIDAlmq3n3KD/GM+U6SOaMH9OEtx
jJPGlkqohLO4YTdByvQK9K+jL1C3iJMxJifOfabd1VAWYXyJTU6gB42qYOQkMKJt
6pJg7zzFzQa9cngN6wyPieJ1uranfVNosBcqMyI/KFBgmwQ9yd7cEBiEgt1el25R
JDt5q1Pt0HepHaXX2AO4c4xHgvmkNZAX/XV3eL3h2CIad0HprAxgqu0AKzFRyf+F
Z0mURBhs7kF4E+O4XccfKj2882DOEL44d2VkGC5lXcWxWdSFBQMUcrIj+6LIZiWC
EhHsPnPL/In40SqtgAqxLPfy/VyQy0DyX+0yw1/ZuKBp+HQ8Lc+inlaRwkr8CKyx
x+N+O2stnl618s/qx/JRI+Gw7U0kxSAXP+syelQpEO5/7ssuC04RwNZXm0DvYDlB
fbk/i8euLGOz4KeOfCpMmPqQLL0+yTpjr5HHwbAkneo0fM//NAcwN/wRiYQFeyFf
sJRq+7vBk6QbRYhJYhi/6dc5x6wxuebTbOJum0DuYkTqxA+Mo9yrROdBqWAg+4bM
V93adx1E8Sf3KMTMRlXyWtutCjHH9SQQr8YSIhHs1ojvVgFoYaPspbdg6+EJoS1T
UqG+AqklyDD0cYoXZHy56gr52rotgYCC9y+ptRzKNi3fBc7AQbF8+JH4WSJxGm1D
yJFCc95LD4tXQsB9uRtuOuLjHSd3xIidOkoESvKBnlIOqZ4V4ZfSTJwUb4GK+KQn
CgackIIxTTW80jH8QEwlwXg9mZNxYj4Kzaoj+D1UswDppZ2pdL2nite07+7JlG6Z
ctUi7ZlLhnZnYyoz4Qq5uvThekbD8DnonuAbNCk9MqCTVSr4LxtWwEIoI7pkfedh
/GtV5kxI5C2nCHdm01VjkjhMIE25HUdRFv+rKphDy2JQzS10ZAsXXtUmi8auk7ZQ
jlqDrIYqC+opBWj4fpRfn3fvvyBduuh/7ui6NFSb9CPUtXrX5krb8yruzybwv9n3
s11xBvN0chHXwjuL63CUXovuRGeM8gitXYSngZcl4jPTedBtQ8R4E+n9nruC9CIE
V4s/vHD1bkrJFxwF4u5xvn8djFKtDMukTcytxaAPcdvTY2r94nNRZIadv0FCYZoT
cStgrSS1Jl0CrnBCqWERiQ8IHaeTblutKFNe8vNpDCc9d5cBSjlC+eKJVnM4XaTq
acc8WQOg7jo6erIoyr+T33PfwI4GjNE/HJPTcrJuM8vYu6dj3j/LEfQbfKOlx72H
joI8f3QBu20x5141zNOuEmVoSzxbKlDi6axxemQWr/gVoydBw+v48hXrP0r7EbJ2
oWXD2VkOkfTbICBPr2A9LQhFhseTaW+9VPZKMhVlQquJCbIYKTGhIV/sGTwnUvB+
4UjLxd7/1/gJmUJYLklmt4Z9Q1WMQ/RdHM9oYK/YSlreazQyqoOr8HafDE6Yw8AQ
9s09JN9sBrSJX4iegMxjJt1BpzVaNtipbrT2lodNwOIbQeHr2yfABCQ/FWkDgJbb
JL/eA2/4pSwuJHuQjhJuVIlNTzPTtoOieh8euhsPn10FUQ0p9GKOPHEKqxSasrqP
1xwTNqBObG+00K+eQ/RWTxfdg7qvM20NsjCei61F35U4SjcgCihLMGrfQlOwZMIz
1NTi8NZOPHqtpYkOIvbuHGqEy7LfRcAVwwQg5IzB7hPsg+oR5+jk70thy/zEPDgr
ptAMSOp3hmkmEUmm8cUVVVUSjqqVuiadQxs/+q2yvUJrBVgSPXajUbQ/vv0X7unJ
XtGgC8gKudy762mhdsdbFeyelS2+vvTHSrle4ZQzEpCUM/oTIBysDbqUt9pNXbDR
2DtGwa5FGmtLH34hW18wxLM/0Ril5Kd74Yk14XeNO5DPkhPQJDdyBjLKfwpDC/9H
jufL2VSi+o9hRKumRM70W2AiBm3avnueUJRcVgVn2LPRVe3pMpSXiOvf95DKuJyi
bBDXgvZkGoN6SEo01IdPMGyilSScyS+tQ55WMLxgiRwbfFoJTLXNUKpl1bJSDOBX
kezOxBQNinn8biQ+NUbUG2qsuJYzD8d+ZaswfpeuP4LXAuw4iLXE1WLly0LZnTeM
TSbrb8EDmg6+nKiTL0iMgaav4VO1EYxWi5//ZaPY9WRt8LrcqyB251bUnyqeu+Jl
4m8tSDqqMNv25C8h8j+Oc1FmaSm9ovTcsWszmrtrDV2fXfX2JCqPItvB4tt3xA1R
Wl0UWjgHY8eurWwJJTNJ6WQmC96xOtSDrkgqEUqC8rK/aqtmdkym4KsNHB3dfH2Y
eOohMWntHJ4jrX9FR2DDScDyagIycixRVb/7tSIkjO3ybdweGgt3qAURl/rYcPmq
zzxDfFEIBfCEvXNaT7dIPElagttKrkoD1ys5RHx/oqdAQt9nJyyRnGpQ6epJS55r
EqgZZLt5+G7WJAg5I1F3TjML6l8n7MD9LAS2cBydmm16bTa5OcnffjmfTAZSc18X
uzoSSRz/Fsv827IEzFp9ZAqLOg1SkXrekLoG+/cQsbmCjFEbwzde+yHc/uHbFkpb
52fnnuXsIRNbTuJMPzok46Mm3LNgEUqKaxcWWTG5OfI9n8jIkp4spGPBQkAotw6f
mcDqeBu6sPvOBQH50dX30/89Qo7NJHI7y9ep3iSnWnMEVrolD5G6JJDOFF0YKZaZ
Y8WS+e2oHYo5qy+FAqe7m6zPjQe4DG/UKHFsG7pKH24eqtLM/QnN34bIY9i4wass
BBOilpGfa7xtstFJnhwdzLOui7tGIpOTiqWeWyuKOpueFC6CLQrg0DmLL8+3+/wE
BDCTerbKoIk+RCGfEpKOHJmGF4rKQCo3ooeoZ2k9mLsu6/3kSJxFoScNTvp14i7k
5Xj5vY5PjIQkL2kcpg6O98Q6/5JgYrJNbH95vUS9lKTU7FSJNUyWd9dGtebVbJQV
Jl5t20DH3AWG+AlcQD0Wlz4Oix9AaXVC3w0LRYOsSNIhCe+tXWe01BpsEnWhQXK5
6fPSR77brA8stkux6kYHl0s+EylPT4mlevZURJqbq8bYpQVswjV7jFgSiZPu1ZeT
xtJMjuuNPTiKS1Py9QY2MKP0OtpBtPFn+GF8O4DthZyok8mq1S1QOXOT5xTc3YI/
HAm16Z6tQN8hyKuahDKn3AEDeGYcNDz32GI8Q2nxwRi8qvBBjUbVDu24nF06vFtU
xbRZB6gIyXI1xrdfLwNB02kqyDGZolkntbfzHcD8DSqwArJT7YjRspiVJZt+bkmt
LV0OcWMCioQpXR5FATeKqF0qEeObG5NHybDKC4ur47R+yaXafmEJvcN1rY+ef4qM
WB2D3osJ5ZE2LLvCyYtJvEWIsRO7Jjl5GN0Fs46foDywdjnQBCpvKkORPwi/0KC8
IZjybk777h1Ip8ZrY3xN8JzvFw1DurWqILp+a6okXEIp3wTytR5PmAtJ52siISqI
1oISfI25iG9obrtFrZ3zwYatiyHWX43VWG2pf0PLCxB2N+K/utD0V2dj/c4NFZNy
EdTI6tPcug3JP35Hp39vz3B4vITGMSi++YdeOYLU4VV2sY37cn8O20eoceRIr/j6
6K6Xp3TmWMy8FqDJLAiDt0XBr1h3bfMr8DGkrQGglD7iOKzj5Xg2hhqSgnNVGqGe
PlmgSgFmI31OQIwIZmT/3ojg2qORaLBlaY/Rqnb3SyMCuvPXfQkwJqoPqQsJZZje
neWyMXMhHoOoDcf3MuRLIIf+g8tegl5SBLwx6U1jZ3/k59gIG1EAH5x8TrkAyuI1
CAj1eXBx7PAn3VHLtTHDCiPgY6xTXim6M62JD5Hm9CZ5QCuewcc2ySmHQcLiQMm4
M2YyqnxdefIYWhiTKEJxhhcZeAxgKhIbbuSY2vPQpfAdqzCn4fsIwyjoVJITnRX6
H2cg/fpmnEXhQw/3yGXQWiIR2+rRMyLQKmcsfYi6pCsdKxy55qqC9YCOfWHZBIXT
MUVUwWlI5T00kB3FaUDCIdgNDNR4Ey51VCOXPWFGbkSH6Xdyj/nSh530PranFPY8
MIYuKvk7ULtutqVpctExI82y2IAcOay3r7XXWKytjBY9vkUZevmikH8c/BKmwlVg
JmfXwtZ3jc3aBZi1wEDLYYpurPxuyu39AuJOcexDfIJJABQ0F6NO9GW0igUkJX3u
twhe+Z/TzjL+p8pzpb6H4keXtLtwZD4sBi09C4kXi8CPDO8qWHNjOsyTfbu5bB4a
DbKo7UPbwqa/1uKg0Cp/hzOTqzpF2GsIDljpNEJ856D3GImKoHMprZybdaDcGuyK
vxRndki62HBwKNLHjBN+yZsAX8paJJA9L7+1hIOouSjODc5nq2C6CzD2Jj/0hoiF
mdwZF/tVy4QN6XHjLjoTlSCivnZlIUKxX+bV75gFQuveljZIQFHO9bOxZXLazTjM
P/IUlxcHagVbV+wI290m4PkNlz5qEhbxKlSoQ6fxZRoHbtoKswDopuzr13VlRvhQ
jT6kHO+pECxfr7Vq+KoAwBGXcU7kEd4SLkd6xwH+Gafri+SKbnJW2q6+exWQcvyw
kSAZLpV5Ub9ERFw9LaXs1QYDoUIv/5RwGIJtDCHI1J8RKVWfLShSQhfiBVF1qxaa
DGfuYtrMAga4n3zF5FVXxLX95kblUFxF2n9tm2o/VOTI5ayBFxHwKVSCjBOOAoVo
x9kv14EDZXYiLNZtAX4AapMJj6QpNd0ApTKBEuWj01kbSvxShaHv58CSAA3zwSBs
CMHGc7dtHhCli5hKsHM713qeEzSXfl2rzMfDryRtFLCxCwnsUxHlw808CXxMOWpI
iZKqy97f6p3GtHJX8KXfY7hPqXy3mbT56zsXNVMo4iK36pKPGrV9b4BJOBQGeqXG
rZchw3vcwJcYIJPI1oeffh1qx1/XFHbtgI2u0rj+D67TEWquRstbf121ksU/pVQL
s5bRAWaQ8VCcb/GsyFNcow/hKtNwjq023yNtNpRMZ56vVbiRqBMAy6cvkE2lYdW/
Ioy2xV/NtJlzNNixaExxhj6vtqnp3TxulkoeM7BaTjlL2UD8mZ+jeiix0BQmmATP
438TjMu8gNmLLK69MNZcsinZKd5Awb8cEA9ygh4xSxtrxfmzR0KuZ+OL4UVL82Nv
qXTMjInm9ASoJ5GXHZZBkdAJj7L3I9NE8jxDjyRBvGpDzfwxDwUF/uS6cSqVC7XU
EKvGodI5OHReLJUb4peREcfqX+DynY2jZFUrakVeYg5oUc8EaGMDUjnN2UMiz1RF
qlUQlrg10lNI847MgLUO1/VDVmVxQh9tqvciQ0FZruWDKBI6CboRp1qT4/IClYFw
2q+/WwpR0UAo1aZp/WqutDRWxTyB2AYlqRvrleOvqk5djOK/hsvR9DlHFzQCtF07
9R+SERo7yj92GuSF3AZ6t4ip2/1LWMZokog/89pLOVsPUcE1g1NmRcntAiTDJbzo
ZG1Az8TcA5gImDuV7sQvmqWaCX8xzxsM6bMIzg6VVw7+cEakeCy+iwqrfQ9KhS8j
iDEvFLePKmXjBaU79qOl7VnahF5z+ybrsoXpgooXJlqncvCKgeKf91XDk/iXqTXq
xQCqU9xBdivRNiUychcqs3Kz1PpH3w8VEqAYpZF5bdZvm3V1W7sqTnpd5mQgsCoT
nKJ+hkJWpSjlB0S3iwDOI2P6CsBCo/Com5O8e4m9QqhdYXT7vePPFfHAZwUznKZO
YKN4rebs7HpPhH6xMPrMlmeXdbhOOJ5LLUKU5P/zTt0d7/uHb9Fe93l6Ng/qvY7I
MmtqFtslReur6g3s5KTOI3VKMuwJaNmwukMTsmFcmP5gjEqiJQTU4aoEeCc6Lglc
litHJlZv+TmyQ9mAJqTEr30LXCsd9yF7567n7h83bHGlVeUncklKrMSVuN/saGxT
RQ+siNI1aLHA2AqwtxzQK9s96wrZpFLkZGqd0z8ELr7u46u8cmtVCY6qUcoFCGzd
DHXlS0X6fkzQ9si6CmkVvfliLDjNjEc4A/4v0b0chNehbNqCic450eKHD/INjEdO
E0KdEAPuAxV8+hITyQyb94ct/VAdFk6rXiMCp0D7HJwj5bV3szz4ahXr/mP3ICZH
f46yokp+TlHyMu36pr8q37oUjGANA1qjZ1qQ7hyn06fKEFnDhbel7pbQTyhmCfcE
VObnmlVUPa4YaJmw9Leht9uDlnhKpy/masZIn6+iL/LvmTIOI3L+6/mS2ZaklJ7B
x7/goRnjxSvBr0OKbWXYY5GqVVDZO12uyg7B1e2kpK0hGSVAyyc41dgoLzmqrSTx
3QdYf8AXYDELRUS+OocQGgcnANMM6nLPeMb2AsWOMWFaNxDmU7gDS/R/7eOYFwQe
prn4qFPBe8Hc23F5a8IXCn0ikO5AZ2PqJIsbf51n3N6CoMzWzk2kfOTk7Zo4hGH4
s/THriBOwmtaGnnxIUgKGZux1BNmV+iUFsC/Ygze7xo17kIHzsURVzR4bi1tnqb2
ym6OevHDGtkWKbWyGogiPTPANRgcmSxbAaLny7rYqCcyMLspQnjNqmCbYjwZZ1Ph
Xun6f4XrWPOz5xaSegqUhiJCueaCFLShFHiRIRF4+rGgFK5lsATVZnxeoknfT63P
eskwQngbzbpuBm/wSf1+wPIGXpvOtKVKjFadXUO9DVeLjrvJy0y6QYVu3sgDMRrm
YdS2uPGj0qXZSKpbNV0GJqHJeqr/Z72FW6Cy72GbV0IheakNtRBTnsKyyEDJ9IKv
vrYvDsX1hmWpOvQ9e1Z5iPzZJMDM7eNwe9Q9bPW7zVD81XY/oudd+DgiaeTIu9Zj
TyqYmLdqV347yAOzO+r4umeAg2FduD5adpv4EYDwomCjmI030cFQsI4sKLFKrNSU
ZtvSukLLRNxDsmknwHZOLY2uUjEzhg4DPHrTLNmmtlL+M3MHjOGMktmyYMC3Di1A
7QztnGGLNMcDmiMJO9qbAFkHdtER1AF0WltDvL4VfUAfkSbg5dPZtoSfl+HtT5wV
QzVmI2B3UqwCX4XSWYMKL8NYbDeGLx+J99vj4hcSiBCKIUnj4gX+mC9EXLImE6rn
MplX7qGx9LOWGI7IAc0TWEzhN7JhozNiAAf+Cu+x29KrIfzw7wEAfPueIqDbM24p
eas63eAVD9ZcfdtzW1nfZf/qh40b6nD1M7ql16w+sqfy1fKn7/EVZv31nBsc9OXz
r33PK54GCkVhCNfb6hBiiZUhRBtlhSWcpSHFEFzEnrzUk92x9EPBWpyM6JUzwfKN
EWXXSbocGZWflgqxJlv5BeF7CnbXuI0a+9X4cUiZIWacTnWYoBh91GgBA2Kc7G+z
BdFhWCuqBq97XZxpZgHKg2t51WjDw4YpbaIkGnkFyIPZ+DfYmQNdYkqdOIhfKwo+
9uOt1U4HR4RcnM7V9Zn5i2geEeSK8npRdY4B+OzduqaBPXvKc3PdQcT0QR/pFZGz
rTM81Nifm8WqIp5L3jqCjNqrL9yibaX+3FvA/LynpWj04WlObZddsSx9GyMt0NuE
pRUyfX8RlJlraLH+ckZAUdYPNcPjAIy0EXLvPWO9iaiNjo2+kdhrOBl75Wl8hdbu
AF1e+XeNS7PrNzJCsn/ganoUJEMpd+NteHadu/ievNx4+Q5vY4IV6D0JBRLOwJgy
UXgLiw1Mm+htNxLpp5RPSbxqZvEVy8WALrMoqW2f5f0hSRp7x6n8dtpWEyyIMa8Y
lDJgOdZNzQmqdQYQ7Ml2X9oOLuOpiJfGCqmbAtDQhJC9FpTQmJM8VBtSlvbjNauy
91/SbbnotC93o/NlDmHznR2a4A/dPpbQVDqy87eT6zkuhQeOfFG2s3Au7ZNfENB3
jft3bsTuHbGhJXLuf6EWnpFydFj5IHdttU9l47SwBln6+pT1mEMazZDVovh0Fpbe
otFY3S8J/1IA3o/sOnTqxCJX9j0Gxq51NcwsGAAdmXPG7oMZ4Aqbd7zyB2SbmNfy
D3J2qjkjzuqeVdu5PYMWKvfvv0SJkx2GHaGekCrU1bhaUpY6zkfeigdJXUS3NQrc
9PDGDCB87rZvlRlt92K52X/sdn4VNgaLWZamuJBz5znisOn23X6s+nDwwb2GOFk5
CtswWD8K7FYTXDDw/T762nKbXqrvtses1jLuDIddpiRd4LbH3Y3+soEf9c4/Gu7f
sTCfG4zPyTyToyHkfPxQ+jowBs0Iug/TA2EsbKJw6FxPpcnlT7fYkwvT8zntpiGp
hhDy7dEu1s+YODhKbxdYKYG2pcsjKHOR9z/iv2e4Dkc04fxK71MmMMyScEyv7Xjd
rOBGl1wKt0LHp8sAjEjtn0i0UBPOmQhVlvHv7hPJYO2rQnHFwpKv8PSfGr5GrxF/
Eaza5NEA38ZLldAXf1s5eC2bJd1RsuQm+9vqSxNnRUW7ZJvzdOf2R02VgJF/EdnO
tyKmpPdu9VLWpredX3OYsa9uvaDNUKV5pOkrPD6pgOmCCHgz4x/yeGOfroS0rwig
kJPw187tDz5xzB6dVpI3b4nxbA3mz3Ag7sx3wCuxXQ5WT+H3mv7DuOAujXNIJ06i
8BSQv3zj2Zu4PyxaNemDPIeSFz4sJIj5AixVTfS3GnOfecjUetMNqJ+6fSLAj0gn
rrRk3s1QSxsq4wDkY6JT2TTdJ6xXwL4NfJe2mnxIuzv36lPMLPl7lHWJlIljo/dQ
gqy/Ye6f21UIPGZsLuVB+7D08Je3RP8KD/tJvti20lSBMSdbxYerld6W7lEGJ7Ox
RI7zgn8QfjWTfaEYPCDqzbQtWM8FPCD93b9KOXRu3klY7bS+gzipYNl7z1MEbmiJ
RNjlr2zc2JRfgoTtgsJAmlm46xzCChFNFAPTL+7DoOEjr94p6D78sUn7VQv0uvHh
e04CPthlicD9ffivmuXJlaDl4cfm0cxIJ7MdZR5Kx27OHs2WENajQSG6UQzYtFQi
ktJpoHg+GkvX2RPjqfgdirX0EoWFAA1432KUl4MR6VO6GlqDrtnPokLVPHLZ+fUW
kiovbc/seNVdq8oGCJehHcu2TmFSpmiyB389aganPaVr8yQlcmHMPv2Yh0hvLdpI
lMNjdeFdGLfQrGSSdlRnMGwc+koPwVACaDCj2V8o+oq17NBKj0veURtqVeW6/ePm
onPm9K8kqKFSmmKCXGOjF/xdi+XlqjjVwX2xSGJ6y/V5gpirAeJMOjavepmqMvaT
SzLYFYycsb61lxk5D/0yTGOQRAn3LW7y6bYmMm4OTDlzsyp1oxf2upygCwI5hUXq
gRpClcSrXEoxF844rNv7dY3MCbh/Ee3QCy8borX3Z0iEvJPDP25Nm/hVzH2c1zEb
RAHYWwzE3wv8/GIS5nO/6QJAOyEh6u4VJeB/yAM7ODpJSnn3GGwhXf2DlHCDh8g7
xx9WJfeqFWox8AbZ1Rj1r5ClJVZ43F2hxtbNIP1S4dsXXcnlABEeQnGaZ9hXFoBe
eIrR9wmzjNjWtZFZd/SraHIzV/XwapmysaHcksa6xcbKwyJy2uLjq7B782rGvEwQ
EnRWgo80VeY3kWB6O7sW1jgRWdRQYpX8YB6k4ZBCEHQhkOTyZdPmDjv5N/3O9JsE
cZkpYpy3FQpIg8mUZPy1rf3bvQpz8Q8hNBLXcokJUCxMBJwwwHCgN7Augu72xnc1
HaNzjbgGa1TBeZvsnLQoG3MePEyT+mW2n6DCjBUuh8DFWFfDzvPyR7ptDff8vcq3
8/SmBdAfYWWOB8pdCHU/ZdIU1yTQMMDjHmwLUXTOqF99rhkCVA60tzHQ/AJpvJl7
VnjJJodqpM71QiLFXQHDYMyhBY+7TT1Bv2aBp+BhPE7LLiM40FJ++AShqpmdHcFZ
Rxf851GwDFCs/onOoECXtEXHsEFwP98xif3a4dnJsAJ+iLdCzZKiS6pxfG007dgc
FdGWm3tWFuvyXLkR1KCb9/2FH/EgTa0vjKwcBX2jIbKZQbTobWuJrTZhxSutDQUJ
U3mLMg8wbokMTXRJaEghiu3VkIrZE8jf86SD+wJ4JAZE8O5biBtATO3d7qWN4oSt
+vxNF+P8bS9qvCw3VHBHoSOZpNhZi7sAl6Y+oa1ycR1KfNqZ/0y5PjgK4hGgq92M
hHaZJd0o1pAZF287YckCMeVhs2BGn/YZqz08i0vwTGLL4k5+nzhDyn7LCpjYsa0/
aq01vDrvnxhiQ2YQOv4tX9vY2KnZbiLL51mKtE/h0zyjXxO0L04JZH6VhEwSKYSE
X0kIAG/K1fDUZNfUn1FVhezzXIEiWg1PL8sM8HSKMvnH8tOnN+/RbQm7LWs7YL8h
Alqy4QRCDDY64w8+M8lmPKkOMvsvKfNZrOF2lJuG1BJs7bbOz7WoVSZMstn3E+4I
o3URJmYyQ+k4RGpCnjIucUYA174yLf1nbtEHhbQUr+uHr7sqznUVwUDJ5W+HYtA9
Vt+y32snepxwFl9OCdokOGdoMeKk7tFyw68oCFX8NOI17vbH1EVSkmqg3+l3K2Ey
dvKHWN7G5ZemPKLo4IQT2NFmn092DRI3bw3aj/CdzzUMWPTuVMm1oYbv5GxQzj6K
1gUoac8JMelxlXd4Gio2VzNW8TsW14IETzCuXkxohoXs+GW9JMcs9wjUXPmYMO4v
tk0P4jEcSKPVwlSSsYkEKkbr7fUW7aX8Tmb5wWibuPKZDPqPsophPMR9B8PF3cfY
WnMYHXD+dSPnOUGiZkbeaknm98fkZ4eWp9oqte7vP5+6RYQmnuY2JuQD1fVK9EjV
Qm5tHmUQR9pN4z7G+wTwAiej8LvB69sekVmBe4lRBQX+M7SP2qjIZFvnUBVeJWev
oXJJVD7OM6CLu2D8ptGFN+nwhv4ehTQK+sH8wJzCGzPkyWQFi677DtSPKqGhQiFC
3bSuIy/EmrR22ZZcCfHQYkRV38/xF3lljfR/ElQxQlEJY6p+ci9g7jFnzU2YJXjz
3cEnRpZZIalImWvftbeGA4njm311FyVZMkUmX4ODf73uP/E4nU/wxXxYYFXdE1hn
NDUNiFf6CljEpwXoKFD80dgSat17PuDICj956tvqH4y4viSXIay3V6+/DxKRXZqX
2rLIQVbMUhtoGEayOvSukB2AD2LBQSJX+33XrFS+0TbLmHnf7J8yWTcw9larP8Vd
FADkXGpzNT8sT0GKEW03thvP6jyeeAOw9S00meLrmclnmgw816l+qAak7uxl2kR7
k/0QhJXWeV/+kTva1xBsuwwf2OlPGuwE4dnPayAdfqkmOVhwFYLghrKEFmRgVDK+
ruP8rxA13fvUgYZk3qHlW5seEonIo0QVv2U+Gz5YJjT+Tr697tOXATifEQGun3ku
wIgo8WmInwd5RjiCm95v6elaWXSRr/S137MnNpBPhGdU2cW94MGKVFYpsCUeQ25v
XOPm6ixAgXJ0vjkxqW5KpgrglWzFbJs7JkhBM0D34mORte2vGiITC/ipg9OhYeGn
zaiJsLAQwbLJmozueH/PoPw5mb8NSYw1qvY48i5EXiQ9aMOO8pAypwJyEdeX5YFI
euzdut8mtKD3Ypa/N7o65OeO70D6UxZ8kV8VtfpDFRPWr097mJVLgW2XdWwHW1vp
a1GZDVERsKUZ5suB5MmmpYsHMhHAXv1uh8AOQU0AsetH6URmpEh9QD2CEqPhkRcZ
mn+Ml4RxXumFtRdKsMD1Z7/K/JlXsAi52KZFEIlbFsJWp8bEKErmw08wxzANmf0Q
3zxOaSHb+bZFjRFCZey0Wt623ciAsPuyQlNJteCepQgqEwadiBvMZCLJaddEh9+P
4GS2ULyXwJdzuHuGBM2nmAgg4yWRpce9Q7w1HoiOTAtE+KfSU1FeeXus3RSMDO0f
qKa579y3bWIr2sMvMAm51+4wf6WsLSJg9qPz5qwoipn9T2nYZrKX5ieMhJzhgMq9
1E/WchzpAAxi+8Zb8g+F547NJtv+ZW+YRWaHoMa0h4LPgqKBaqfgvW5UFwsGrp5A
8jV9CXe1vGBPBmPhuBtcnMyGnc0Si1dsf5tXuKm7wGP4AGeWh6I5qEZaNpWWJyTi
2ZvQOZrj7mM1QdY/AcrJOGGrup+DrttvYD5gGRMdiYO45Ujj6bnzuhMqI+wrXXQf
hkz7ZR245qYfk84s7ye5gCgIquZ4kGhHbESZbQ+YjINGuuONwkx8XXfSjyCYeH/B
lDh+89nepCHdUhTOoPVbQ96DyVWk4/6/Qt1nMxFIYAiI69I4ixioYfRNAVWywpw3
vjy3unrK1mOYM315PhRULL/vtp2o7gfbZDCCh1B/nTgCfbwhkMGbIbGZTqueLDRf
2a1bO9GmPNk0zHrCoN6neajbhZjlwmnZatJYtLR2+J8qS5UsDnUvQgxf3bNXfzuv
U1LOhwGQmCZX/pP6/4GEvHHoqE9hosx0gZqNtrrwvKusWBl6W2hJLIH0XJfA6/ad
elk/4SyOyPDaf2esD6L1rsPNjgef84LfVIi1dBNYlY4jesaOtMza/zs7GT6CT7P2
7smn475x/UJzImvuXmLeavGh5oIwk40k6At18RxtJw/G3l1KH2oVHv/00Pfwx4Hv
3CedeLoXBkpEagNHGGq+43XWpF2DWGqnGJD0CjLNhujkKatayw5aNFTpRYumiJc/
bc2RW39Su889pxwq4Z8T0Ep+dhv0YlgU4tS1TsFw9J9P2tMjrb8ItfELNB+KbWCd
JNCNq/tZmwkbEZtxA1Zx2Du4lCilZWXujm6AwV80TN07FlUdN5+zv8ix5c2ojQhI
WL5xO3k1huiUDfuPbflYOsMEjZOM/ZPGSaEkrcb6FEjkHoIO5vx7GTGylOot4ERK
TJFEg25Bhwfd+yYPYZdNRF6hNYZpPiwkxrOEDUZ3Vb62qnaTLw5oWEckzLefRDN8
Gp56CR+tVJkSXvBAj8PtKqlbwBysKT92qqgPJVND3xfnPcc54Z+OT+v4kN9gxbXH
u3T9Jlqz9/v1KTSO2yxwXsDXqb5CYIA+VuZc3ZxhCuuO0ssvJD6OrNeWL0dN5iRq
GAK06U/Z64IFF1Ah/XzRSkGJxfek4uduoLCvB/y+/C2+ypcC8DROn17QoMb0+8aS
z/Y4V+R9tMkO34qbWEDsZYwvcEYrdcbW7BFVdhm0KjpzwGkbOceN49Ce9URYLD15
XYPT4rnBEwC0a/gLCSucDOyg37cFl8ZF+3thYgRprvVYXTSWJ+NG4SPZriwQQPon
uvlpSLoarV0anpxwdMLyqiHiLugaxo0kW0hiltaJrxWgXqJ8hQxYCdXCDkhb19OA
YwxtZQRen7bjIa15Th6ABAtvd8Onjr0ntLWgJ40tMaW26IaB53vYMD+hnUfdR5O6
jar9F+0OA8/kDZ9mvaQ0sB4efleEk8i/EnDB6G28N15SD0heqBFrIyVAaoqGYG6Y
sdr0DbaL43TB9baDgvlzfWXz7ptuw7j9gvEf3jgWigh/Ef89tDWkUNQxs/knJvWO
NiyWfHFVgzpxVspcyOnaUAaNBhmPyVL4CzvWXv2TkjJN6cI6WEvhNB4dEAwOmHz1
ywccvypQYulRgwkdT9KT8lvOHDyzWJHhihI+eeMvMOu3DFdSlKUt81uGZYaiJUcr
SsUQe6tog5iScY5jI+1hRXSX5B6xgytngzkPJC5NvjpFO/BMny88nGIoH9guJTJx
tmY0lYpYnX3w2nsl6lk4GKLsjNeWkoD9GBB4TNhWLa3cXxl1ua/bPDauAbWqchjb
nnjbVjIOE67bbCP2ncHzX6Hoo0xi3LdxEPKc70Ik4YyeokNI65yYYi15RYb2lZ0T
79DiS0bnOQUIyr7d1cqQu7gYh5lnAmAi1FQ2KSol92HitHS+ovTH6WkLBJVCVyrJ
LUzAdcNcX8vPxjo9UCZo6S/3Q+OJgGJ3cqVlQ6uZ1of9OwYe40nMSPeDxNvti5C7
aqBUu6LhD7QDLg+1zKSVanIpXf5ldDmhi4MDMHGzCSJQw9oTsxpWdQcgCuqfS60w
h7+RsB2kzd0TlL8G12SavYEMRPIqMXw79oAeb47u2kLJKocEmPDxjdwPLzjRyn9x
aydd/nOVEhjdncbJP261EodjeyQt/LuD9ffhTnX1hbAaDfhb+GpX1simYcYk1QZe
l1RIu8jdizFJRARPpMOpVMwJNMHSarpvbsm56PFLiUd8mrZ3QhUtq+QEk0EPDJqS
WVH3bKPpS+xlPC1rfOuuKKx8OEKFd9WC7Vd92BWUTMoq5bwIDqcZPLDdBG1ul6mr
yGYbj+YMRZSud1yLnnm0nVuSn5bIf1Jnzy3tiCsxv9SLVFmy4jMTJxsrF7s+HrRR
5ljdqPZZAhlEBhUnNBxTDa5poDgXzrEJjTNp5YI6aOIPu8Pb96DQm3OCEzfaGma4
UFjNZNKPtXY46kFOEKuHT0/yEHbrs+z+88u2iWyxOY4ODVqdG5PKa+VH+1G1s0P3
FYz7w7HVWLjjKcEIpL4MsGZ6P5ccDhxCjxN2Toid28Qb3tURnyR4vvGR5kVoel8d
hfcWCKNi5yx3CAP+IixPGVZiST+v6ntlMfmo2g/ByoKNgvJdC7HYIpxKYoPOsi9l
LQir06gfEIjUC95kpyT3gnIiSl0yaTWoKoGvktr0daX7o0we4BxP06XPTpyGpuFD
yrOXsKF5bByww0vMiwsCeV8gXvjVoYsm+5LdWoLR4lPRuZ3HXml9uGNtFTbhzqey
rxb97hAENFn6JFToRa3oMpt3QY+kBbZKgh0dGr/GjmtprgArSox6bmP5SGV0E9ya
nYs2Lz5H6uwFzJfIhNa1RDqhZ/or6IfDrtkyFPvtqq3+Td6ulxsnKtAFC3tE3Mxh
PD5IROukIy1a6thHmo9NVR5yJgoJZSb4Avvjccu4h4aHVf89ejifkL6QXAX1dBPX
lLGpnQ6FYJwOh5kWwYjpcPHbbIBmA2fYjAAf2VuOTsofB6p7eRTJvwYLJAEU0LcW
vC5MyBYlkrlEpPXtnOYwhJAzcmgeqtcoBV/AppNlgLnnQkEYquvo8LaFIM/O9fuk
5V1lAWjlvJYD9kDpeFio7NvrXGhCxdW9U319msBih+MKAtdqH2/q32FhNtkIljlM
bZNh8QkohDQ0hsxctZfeAAmOvpOZgIw57jpIHMHXxIdAcvWPsiYYGICkFAZHV5c1
FuYtYLYCRXa7GKV9R/jNV608iiBSoLhBhKXWphf4e3dM48LwHvgXBsKIHUDmFOim
M6ytFddWNTTvMv0bPV1iXnjjV8s2Zupikx9CAC+v88PFqWdjx/RUD5nJOV/Ro83e
eh0JKihnW1WK5bF5goM3DdIGX20IxXWYAtkyMLuBMubIgr+VPdI23VB4Ph+mwgUl
3jP5xj2O5nUuVIikr7TSybMowJqQYIbxSMqgVSX94hFNgLHFPICA5NWBtsdFLmOx
prtPHEEW9GfhpmqaTlDw3JuVIrq1LX7kQZBAvXxwkRLet5j3S3tjaN6HwpS351NJ
xvUoRrmDgkYoKHPvWpDecTWstf9O291ar6sWr8Ew1vH0GhlJ/W3h4zv06I/7ohNg
gKrA9msZ+6fNqbUVhn1r5LOwjkxjcrlpMfMDonXC4KKTMD9YSYmQllruPCwFFGcz
EhMUK7eQhHYXXpjKijkVqbH26iibYvIc5PsUcmN0Ug+xoIzWHdJNnDUf55RJK4b8
U7bFtOglkBVQzDonESX5S/sMs6peIKgIWMbb1qtvNY3/RcAgQotvpRFevs32eWC+
7/OoZ1luw9asAYVtl9RnpeW874vaxKGhDVHuM/uxrMz9cAUebyogrvs07BSXHkFo
GqPBkZyXJww9uvxoFqJQ9EtxPt45i42vUCHYPKg6cf5/3Wx0nzNMFeXsGW42Jfe3
74wdPIZsa+LI0kAOW6qHbpJl9UhBWGUfmN+VEemQhBm8gs6Xyoo7exKSnByGyuKH
iM6/CTJnecfg5qjpa/V6HmecNuCy0/o0wqekFJbZaOvod+UIZ269O8iqh9RZw/+t
vPrV/Mj+4y5d0FOZrnVFI0XvLR6bhwwlXUE9P49YhJgFK3fk4nKvOPKBBp6iLZ3T
g8yA/BL1Jy2ztERuZKPZ4W+ZqMm46Bz4cYGYPOCDLqGeJCMOsOHhzEGgF9stlYPa
py8pDNAs5NB6iBhUPYKyHDyt2w8KHW6xNHY/GVAcylYMvE4K1USf+GX5AUR3ePlU
WFhMml94YGZi/punicbGx7e6R341YlIytEvL8R4NcFN29p2ak7Ih/DnA32lxXHoj
UpEmuOdhrcJakTCzak0g3b5h7VMBISWYuKHP9I1+AnWgTomJpT/YR+Ci2mGLOk7x
EWLhJK3esPczLBp3CCMO4KotCbZpPjHgROxTWznrl9DbrbSpRkfHhnTOjQ7xaIWR
ulGf7H5JFyI9ueZSQngdvlLFmKizEv5w0zeglPsyl2hzvceuNBQMrtrlD+rFsU35
FYGYAe91eDYLsVwJuK6Gx0cnFXLzx09qiSJKkApzj4Ahc4juAlTCM5O+5kxKFDBh
M3wQBHeoHmCfZWzrnLBtF/tmEA8uOBjE3qVqjL54h3yQwyVXW5WHH3J32lJZN3We
L+TnZTmJZR3Q8LSwH5f+p95HDp1DuMDzAJraUDaMsk9Ol1fboJ7gNdjD2c9gobhb
j6tCZwlsen3hu32rdyID4IFZKZZvj7FN4G59bQzCqYlYydSa36QMbtg/ChMw2QnE
HRkUy3FaBqIapdqlWBI+MkuuUQu04+2vVXxiSKGuwBcbFYg3Kn6p+tfSnJxitg3q
SwsdAod5G0zaw+kFhRf3BOrueHz3es6jEnEjCHWw6J95Aj4akCJIxfmBli099hUq
UDAIP0dqfg6E42xettN52iEvsiV4w5S9vlzohdXmv1gKVT2+gDn63STDYmgWiBcx
/St2tyJ6dpPHhWoj++qDBc+qWSVSHl1Zc/7B94IqYJFaEGZO/65C46ENdztwLCWk
eeYtFiu+FS6IOKmgfhH8j8ZeDoByksaqmbRr/5VJREEnIVtew+8c1S5ix3SZ59WT
vbnW6Isn4tf8KhD+j98Dywwcxl+Kqr+EUR2CuvPBEhyJrZrmCAg2QhgAky923Nbs
WfzRHBTd0QAQQ3TaZ8cCX9NBrisgrF9LzIx2jrRcBbe9qvCfNTXfeqohk1CG5bm0
og+Qyqud7irHiJAMIPj45aMIVONxUBe27Coq7JDheVktpSMDpB1GXShib6Jj/52n
qSFQLrE012BofGWv7+x0qDP5EP/XqmzDkh9QyLYY9MYX80tSfpZuRYTRub1k8yM/
Sn0UrNi2EwGH0JewwGtWVxVEmJK25MdgtSp4c+RnknS73KEUlvE3iWQqic2ZzbEc
Yo/Ui2j7QJDJsyFoopt93DFkz1qaULvvx5DZZvBsGYTCK6bJZiTmpe7qzr+e0hZf
QpCSzVlRQ+wCoTW4BFoNnsx8t4SFSir/2CHhd272Mmdirhb3ClNFDnpJ9dkvntu1
uec0pXTbWD1UNiB5UN/2s4EwaS716Bn6l2a9k4oL9tiuBXMhhmXQHNuDqx7sA4nV
U5MA8w0187XdamiB1PhLF8fB5znEcNiPmcFoJJA15NpQ/ZJvN2XF64J5PkfaW/+9
2L9BV8Ni23ZgDMrA1svxaYDI7q3R18cSp/EUhWNc4ufADNE01wZxIebPtNS+cIh6
LJMZvcKWvPhNImJyCNVKvn6/MLHmxq5mrZExuwlFbHFoCiQ4XPVhk24v7KfEAGB6
+i3D75DER5MMeQv87QzMRKUnnZfx2z8TvUOOAJbjKg5S+sVwCO9xhwNtXnBlCcQ+
BQXCzhpsdPGZbLC0hiTcHnrYiynJ4qKIz7kHQh295VYmjjyg9gDcGOJ943gP4dAr
1ZF58UK1vtuYZ1AVzPJnCFA5bp0z7Ujd0BmXMGGFA6eNjWmwo277AWSeefAWqKBF
+MqfxJWva2EwFyvpCbqkoBrH16RALZOq7Hnuek2EhKLkBrobsxiUWSQyQZTimqZr
4DewS6rVmz/p2VmZHOJV3759av5yN3N/T3FsqcW7N9ZNiPnUQIcVbkDxWDrRRhua
WVbIIrV5CauJEfr2rBcziSeFFC1zvBYoN1i+OhlQONs4Z9Ei977uWx4rvNYFj6Wi
KSkh0tI6DD303t3zdjVelmwFuSdTrDihjBOltXG+wEyPSzm3JIfXhhgX0rcMnUN1
g1Vq/tUIcx9dKh3yz/9eI4YTQBB1HbnwhPueripIaP30SLUhWeVgt2Io0oeyvUGJ
aPbqHihXJjSEszurGloqDAyg7Us4WWVX5znqmx3cyfrKSGC0CpKGHYWfh09pNaub
bG7NOOWMiwCsPEn/A2SyKNT6PV2ss09cyBNhj7r+rYhNZcTzBezHHfUos93wbWUf
ZWwbxtInlfrYA+mshOIJOcKqewEcT7aoAA7pGjvu82pC1qp0Vr55X0Teixixe2DI
Lwt5L5L+beaze5v8erhRAz12WAIt66JIQyE5SjgxUqpe7mz0j/plUrxsXaCJynAa
fFQMEFEU6/KrEWbSfaK/RM5lUmx6POyjcC6MgM5ujkSJSiNO7eqd/qJYPntQTRnY
mVibzmS89Javd8xW5qIou2lbZ9hNcA5f66wKvHNli3jz0NZJJaQUl3QOgazP3Pfv
cQomPAoRh08gGuu2/Bt8vzrmDVvci0e/SagdHtxp9h91PIzM3POHNIa7bEn5duXD
5DuspjBQrbIW1kEpv7BxcoKfr5A8+AbIExwIiKmW0wEPRru1aSC38MjzQUpvbuFm
/8k+0ZYeLp00U1T4Y3KsLZP2yqLScnS1uCpeFNYLuCSbcqpD6vuQGNExYZpmSiOy
4BduLAlCfWFMqcZkB8yeC/jlDLvogdlJRgAJoct7B2cCDf1tMb5JQQmlbn3jVwsU
4op6PpdIq9u5qt0aUhOwzuAvfeGXRCwMBMZo83OrZy927WgO0qsfee11JUC/KJQR
aY3mpxhqVrXTmZLqw8QCYxkjy9aAwp9Kbq0Tj16k0d3bD7g1ySwr5KAjX9roCTRg
NT28irARvtEr0IH+rBUEdT9MaDdXFTUwWspgJx935g7+XEQ5kGBJi4XTmM5oodiS
bzdWvSfUjGsTEpST1KARfL7YZGJ5jn7XzROBLpEdaBSLJSLkb9Gez+DAMINhkBEP
vnR7PRKcvkeoFBP2vYp45XFdC1X+rCBw0BYZGT1BAE0nfcoxW9lITFkPHrrLvuDz
/Rdofjy4aVYFZ5lN1G9hPcru6CcPbBxWzsCxCH+/khdmBNdf5mzR4wfr+pqlDwjm
9NR5bnFxmxFFOpMUoudS9Mb0JTIgPZtRa89v1a+NGAvdv7A5sivfh8G5xaKL8LCP
dT0tvh3q5B+wJ43QglXgW3Eormr4PLWvhvzCHTmHjrGDOlgBySmPVxbYVXSA2UBx
HLBXETG1UBGdilF+aXF68Y5kOTkMC7OqDkkZ+hEiV4R6ufPv9bkXHty++2a2BEp8
S7TQQ7vjk16LP2U6JPZovweAgGZkumRIYq3fNUtPvDujHkjzK4NpfJ042rrR1FVa
Lkj4HmhV2gyGY/YxJCCaL/REPC6dhbLBwsFrgDl9UIJazKad08p10XILd6zJNDgX
cHaKGh/UCmZ3GgqXHW99CFVfDYqia7zQTikQFdLEMbkdZcT/+zaeglOCyHGvPVXL
tECn5tq5BuCmTF5r/2ipoHBtBD5tANe96eqL0iTCtsKX5rojYComs0OeGjxuceS5
pEKBDdGmidC733C+rpOf+/jgMWnNVhmPpPdrdeOFaS0qR+wxzkDorPYbz4HhHviw
rsC2SPAU/nlgnmRH8w3SJDYqPOjfSwgiiFCfWEPJSCgcKbfHlu64TYMRKI9RDM+o
E3NdBCrTq7DzoapHVypU9807kuJmNbUaH/wh6XREESLqXBzD0ZVx7u3GhQEEdnez
wywHgVbH7LQgu4ErgjH0Y9IwMpuAuqU+vIV7jKZ6npipGcRRZcNJr3pmSSK7SI3+
UFccXOnmWzpFPNjuo6gCZXZ9h2sSy/IOQEx/pOFsa9JLW1wK0vAI44c9K51FhlgA
5qeBVSZENz032X16SbOGBvnL9Eb8dfHdM5rD87qZI6Vna/11Z3Gstr4G1caoyuOz
gDljzmT5fbvx0AAQVgZKLiFoy53a2pWpaESpFecZ3/lGDRLwpwBxFKVqa4V6Kivg
2YAK6NR4CiPORvNSt59HGx49pzk5NlBxNSnyaG4NyaClNmfuwnT6LCOh1WnvGUtI
u7z+R++IGgYLgG5FUQ8O0Mu4fAU+oLC/fyOPDQrBPCkeIMZZvIHvQm3oYIeQnLz3
OARAivCWqlWs2WdjqRXiRYER4OQv4YlHm+tXLj+jabjyk1euF3jmhEnyFH8IiX4u
dmfX0Cy3JVIdclyXmggF6VD2AOGACISPkuOELjRfqZFnvmuVdecBdwHpbFNW/hlU
MFoVfi3eN5Z6IqkyWhp+mAfNly+HaWMLlisl/FvXr+/ZhJN/3RFus+MkbuOQlp8X
LSl51kcPMtztUp2WD6aTK7CQBduNeMUtRnISfU/2I80B2DUpK1cIimN+hjwRNmxp
LVQkJJYq7/k1EY9Kb66wgn7Qxiunq+ROwHpFWLqhvMKReFHKxxbJMOMzkR9PZiCj
M7hPQflidrKTilBu7FJacqnoyKOiNx1sOCz6+J9SQA2N3M5P7yF+OENCx2pb8E3d
bK+B/t8rJneff6mRI9Y4cZ7hkthY3mnVGE5Ho44wgwh+tj1qGmjmIxmhgHoK5x/E
z9juNSjGUwQRXbqAqhr24Odg+vBNY1R+RQv0boXajAe3CBdRxOGDycpDzRpjsB7n
YcBSpdsV6v6oiVKOnkIeqi31VyxrosmL5JIhvuiOlFN/bVSnuj8DuGWNJiwCJse+
DLrXVUJu6+1xOl0XJPW0b9Fb2fKB9YdPrbIcDAuTAw/2T4xxqVgALDZOUD6uL5jR
yvNh4/tKT3/J4w3ESSLgEzIT6oXewOhi/S0bFEbDtfT8Dir/8oSyEEWAZa9T76ja
Ll6Lm9kCNWVEO5955IHBWIFJxW9VejaPPHMVpCBNEijfxYD2apVdkTt8HYXOIVc3
KDiJtJtjeq7B1SGxWjwhEutMzFjXcM1Vakx0kO8KLeZah9l0Fjqz/UHoaPQHuQlG
PryCYhM7nRwribzETVbWzR0W6/fwkW4gq9+jmT9ySWYhIVDMl6ka321OvHwQqk9O
5m0pM/Z3SYS+hABXTdIDbJTm4gGSY1x/vQ/Cp4tmhvAUcQTWpNQ9HzOtXlGGzbaX
daF10oe9GWG93RupCt4SdhWbO/k2ojbix3vmURvAP0ghQyXEdYl4xp8XzhjMwsQE
1FyMQU5cejOVJNQdZCllU0XA+xtSrcijZqMAyPo5GqyfUz7Ayzi763euBDlWU9fV
UW7xOf5OvIDWYsEJfPH0LqiRS7K9f4uNgrdZiuFb8VahUloyhsitf98VzOAEPgK2
YPAyUs8hl8BRcQSs+P80Ca/Vzb08sL47HKH5P3hMNJskJSpGUJ4w/t5YyXNbcD+u
2r+yH6Sn96Ll4g1u6S/7ABVTbq8WxEDD9IK1g9lodb+fvFJ70M8JZxKxjoh12n92
MmaApIextcFCR9mGcPBybBsTSUOi/J2SgxP0fUkzFgcXs67qm40tFwON1rTt+9Ip
b0UBsZcaYZyXHAR0E7sbUtiYf1yDhx2qroStZntvhGhRRiP3yt88FFjLrz4wCISy
SW8JS+57yPbrcO4QLZFo+Ua0GPFGe+YuSSu5AscryuACE12EaKyoxX/EhcofGcvi
JKRf1a5OkyP6E21RcMmJup6zVqH4ZsPsbKdtWLZjtvAZoXEAc0qaX3dcOsuW1G6g
s8HGEWPLpOlmX9nPI2Wh2fpI5JHOGivf3dLWjoderR/IUydgKrrUz0yhYxY8S3s/
CxLIka1hMS7giD8zQRYMiu03rIUOAugctMktK9akoRcNWog9B1NDi9KxyJqtsu6X
/YIvcWai2gU0GzCk5tGLlut2WLi8RGsCZuvOcujMFUl8unFuu+7Hwup3Gj19JyLV
0D6zHSHcucj4UHMjzVPwRvhinTuOcjvpJ9WYR8vWNd+pHemp7n1n24/CPe3seFhJ
aHEAymUCv9qgeshVFyxH8wqncWMS285KaJXdNTUrJmFHKbPfmW3pvDJ20eu6SdsK
zRKWCMbgbuDM3/rv7Uk8q/8C+m4aBi9Ey/ysxxzMSVKzHeGRSaAemkho9S73TNgV
bEpQtOCG6z8Hu7cr0foHUUtlhUONyjczE7RU0snjaQC1p1I3pySH9JQsveoeA4gm
aIe3KAnLKkU58msEua86QNOD3bVZkc2I/3zhLP+Csw9DL1b/E2G7Rol3H/uM0Q/t
ktgp2pKNuSNWQJU10Q9TV/uMuypK5DpCcwerd57dI+q0WAk7ZptEWzluXGT3YHYX
AleBsdmhjsdZx0Ckx5F1qpKvBwkOlLA7vUjy97Nur2JLZgLHNIajaOmt/+FBdtde
p2K+eiIEB9RNMhEKiU6OQ6YECOWPyxcbEZTBcpXXJHXw12CNW18yfbHK8U8gW0cR
jiNKqUfZQwF5aK70Y/hC76rOmjCf0lXW0Gy+SLDwNEKZt5BdTg6tlgplR9zQv7Be
zN9jl3dL8Ou3Ajq2gKfrI4fwlqO572fw6tJ1mnnK0GnoYXSGPQYbmYr07ddTu22b
s8s8ESCybTgDIZECgJrHPauB98TJ3YjTFfR6zmkg3mGRPoVh9FbLoqVUfK5Uf9zx
q0dndSCM3eC+Pt80eyWg3Q/uZbqDAEtVXNkBN8EE2uHvpdPq5Bc72y76qr4eoLHx
+vCGRcTGYOtZ0Ouh7gg2zsbVd5sUz3sjwiVILCQh8zfYHGGNc/1VaO8QdvymRIDB
V2cSjJA2L80JO/cLER9ARdVx2Y0nuxz2XWj94VbqQAtixddJggxDGIrABptJIjye
/GYC1TctI0ZkvO2GScp123iGgweoMbq4rPZ+ZRbjuPoNJ80BgULjOUTJa/pjPSIG
pViANx8O0BIDz1XZYCgN4CogLBjb083HJ2MEp1gkKdQzJx2H51otIft60Icb9OI9
I9fB/wnlOo2XIrj/HSrpcrW/5Aicn03OcRLBq0zf4O+5tSwx6BpWGz2X9e4Y0rn8
t86QtMpJ96Wqz9QI3RrkAWBX8ywUiejdYU5DeCNNV1DByRxKTmxw3Zh2tjkpmTjS
7uDXB8qsrUr5xIBs4j4na3rkkE1Mv4l+zip6jwNNDezUNvXo/ukAGFBZFE+EdYkw
FFB8JLhg6/qmrkJ2bQVvYVSoKzxYdz6ILr2lTmRGlQUpAzvV60drtJPHcotu40m+
1FUT9Nv4knGHagQ4XEahu4cxaW2sU5BjYGIpYw0F2MlO/VcYiAXOG0ry6rfxhKrD
4xxyVxKAsIGbUTv1lzUpwF9pZqqL1c/BJSDJ3eVLDrj7Vhw6bRAzc5cLvYzmJDQS
AAzvKvwGBFLk4cYq5jdsp8WmVpmDgC3r3HGy+67D/yN+dGsIxOXbhpM3RjrVkEnr
WCOpm3FVvhSKx5DwqQomt4T19MfsNemvgFmsXr+yFQTw0dPXvhkWobQDBUDuvx9N
eCbcMDv/JfwkfXIz1rG688wXNgfUpotybK8J1tRC0fi58lqDFQZvyr2SUPkWyMzp
bKV0+S1gcYLvv7oEV5RNHHZOjv/1iiIICzQ3vFVcLC0O10lfvrhA5aBi/PksirFJ
X+RIIyqG4bjbBrDviCiC7EIpJiOTpdqhHuQ69EQSWDGbIpXODXtb6tAcrazwjGkx
fTwp7abK468FHKQ62VqiFdQNCQM/HAHypiM8T2Na9EHX4PesbQGPjzUO3Zg6DhB2
dn1W52qNHY2JN3wXJnGIfLHxDfoYPvIbRHee68ivLWeIe2sVX/DCe6GkRSRHgBcq
4jjD9DPKlb1B6EkBgba3RFq6eSVuRf6FyI2iQ8bQwlgPMv066/HxH5/DTl0KdJ6D
VnvYiqk5vCFNhkKw2+B+JdyG3QYBYxhlaaC2fLpFHaY7rvmf8s1ZpEv7EjNS+msa
QnXlkdeYLfCI78P8LaD/7+dhzwmpEkmcJO884hLUcIKAWiaAnpMB+C/+es0DL/mf
ggnRxdSiZ/04KU5cN8qL9Jqs7FYBpCvGljv51rqCwGi/2bWXwt0VvdvjzShEWX8J
3Q7kqPhJl7LZuKR8lR3ltSjPq+wO+fLvhhEwhXxHEESClB1Vbx0s/AMg2AvrzBOG
ffITs+gcVtFImjNcmhV98w9+sB/o3/McoFvCtQ8Zsj6WDa+1+5ZHRf/+6NYPGoEm
THayQbkZpim32Ugbg0Y5zyx3PHATU+OepDA79C7yzUmIyntxXZc8Yhr1gCviYL77
JkvjQOXRY4uI7n5JKsoeDF3rLodhi4cIGw4GEu0Y4jvqCc2Y0hNbWUKTRVmAGzW9
zYo5ma1+h47CpdxfZ7Kp1HA8YkWRF7vIxyxo0GxvfHrx21MqIfwc9oPwf0fVMZvu
wZNYUth69JJ6v4nqVJyozCLt9eptV42+Q4LJhfzn5BLr0BtYrCFx/qdtvKg8IabI
W/n1R0s6j6SShluCFk7+7T1OO/Ze9lRd6U76RWrMDRSQcyU+CfI37RK7LgrbTQuf
9WQoeEdA4ApgJxsrtEEsNOzkBrnhsT//QNr78aZBxW4UcPFUR/HVlKNGzNdmyqwi
ohjYZCtVYqioVmm6q1XnoxPGKhVmIJrqXUVRwy3LgXujqAjjlNS8kvK3qnaDMlXW
V1MBMM7PeN4mEfya3XRVX0D1ZfZQM5YT3No1nXkX/wGHHBnf/qs5goxjQuD+25wZ
7tnJQkMtd8DycpxGTrro/l5A74h2r/FjNEgW/bW9af4XfEH/jVhPCxFtAa+Kaecz
kGztGvkkh5BPYXZgUUqh96dxQlsEBW5xWGWpVWIoUjk7e/TWCCRunLNd+mUM9soG
oj6mJzj4Bhm7L7A2ZqrG1fEo2kNZLeDjzlUp6fLMI2t7QcyCoKLf3qS+EitfzYsW
p2am2BeeDWE5/JV5cORHbmI2vuqKmUQRU/lDLMQaepHhNJjz5GggtkyxyzKSMkyk
oybAekj8r6ZiKQzvRnGRtZchUmSPcSxAr5DO0L7vvDtmWrfwj/SMFzC5lh2pk07d
nVSs2ghsB9b8O1ZU8xKOEJ8HW9tGGCaKJApjUuzCIghWvvhPcU05+1TFhyke0qOP
o8Zkiw0plpzLLNAKd8zevBQJpizeqX7ltYLjvtJZxC+3EW8ivIslBBW9yluiEkC8
NQg7hfcvlzmQpG/X0oLfDY5TVfgcnSMH6aY7fTS8MPibToJlUBf/BESwJoQNOYjc
vUYuLex4ygYnqJ7nCF4p1haR+SBqAp2odWd/T/Mt8CILhmMsVAdouz9vYlBS92dd
Uf7sLQKjPXgUn8+LJpL+yo3homgA/CClNL0ifTeZcdd1nReUYehkeuyMD/psj02k
fPMTKtynxI++obN+qpieSTmBoIOH/htNbVqIKpdOK+OSx9Pyem2jsBDeaBAZJ8hP
HVLxwM4NzYhBrQcBSSXlL4zrEzVjKv5tta1HVyyMaPsOwKTPBcYk9vgQkGZ9rYqk
jITeU1aU61+39Ihp3wvAjF7Um6Ao3qUsDcgKe6ricGQxR4NK0ya1pQ18BuArkgpq
sqqxHJLHw7ZuJmWZyYpuKN7vbM6S1jC4iC5Qng05mXImuuibjBIBx1ysS5ARevpo
9AAMCUrWqjacSBPgizDnc89reIOdW6sYchf73H8EcuyuMqLU5aj6+EfNMr/689in
cN+C60H0l8fu4B0CdmWbwWkjr+A2n1cfVkxmKbQQx6fVKCG2mNQqxiiVk+oi8BLd
WauVOyVtTsSI3S8MRg57sdN+YZhoilCD9oStmdpVAluW2VqnQkBfdh9weguky/4g
ELQj9tswKSPjFSgCWdQBVYk5571tDIiox2rJNw3upHYtqJInIcbJOJG/DxLH4etT
VIw27SvDp3pOFDwsIHhaBFcmZ/izAJsccvD8bbT6wyKzKn0GMz4Cxq7WAzeUjTs0
j3CnzmwbskGvLMtn1EW3V9g0Mt3ohOa42fDhX7CMYsmkWVntlUWMgqwr9Z3Zwcem
watfQI+kWWq6sDzNGhxPYWOqreKvhQvgULOnQmYQCvPdwCXop3hExn9HJI3I4N6U
GFOcCTZYnf8xsTfj/sm90DIMbZkv60iKF1/t2pYeqSh/eFC+aMqj4OK57OlAnOl+
Qur41jodaJMKr1FEVYPO+vsb5Zw8E1z8q+cdOHKrMugOmaNxyxNmnFjUh5FsT2hU
rvksM8Bkc/yh40/J4KUe9Anko+pPeqB02aWbWRdEGA3e+qUF4dY2Gpc7UHWkIA9V
hNEhW3SyxgQl+vrAtogj+9sk2k6uaKsuySIBXjuJTM9HSstL1JS57BnhR2BoiYdq
bjQu9Ht4LMXrVsNiayI1e5r0AIeoO6bsZhTvyfT9iRoVx2Qyc8RwemBOP2Fa8D9T
nmkL9Q+n/zEk5i4lx/kiEylAlfgOtLIYz+lY+0DikH4QW8CX2+E0zSmkhu+9HJnj
KuKjXVVfvpqrXvZV8rQIYe6Cv3kSrCB/QcKtYgMnKie8mb5CfCHjgrQyqAJqexCf
5XIXB7THv+8j6QVY5tSzgQoZqez/zRUksYgScZmbWUSMQqCGauYt0ye8TOCXOrz4
/R2aXID6tq+sMXBByePx5ePf4tC+hFh0WC66tSDh5tjUymU0dvSxQyUOdrRiqCsW
PMmxb+sOk+K71rBT6i7zoajmMS/FcxMrON7rHEecoYU4fEgo6J9AUy+ZiC0A+cYa
vz6M+dAREu4DGD55shpTdKrtVI9qa4GVspue7WNyOBhVX87+vq2+/mG54021Y73H
PjRq4SgkRKd88qDjHuqNWW8A4LyeLpP1vZ2U3VjKKG+tyOd8CHBRXXi967m1xaBW
2PrM5Sg48CvbFlc8Fb61QoR65/F4hsJmJObaV1fGJQ437BJ0NbRRPNwcjmb/qxg2
vqFXb1LEyq73muT8Nul29HAsXFJ+h1wJQYTc7OdmV7BJHXokvh7L1n1eSsSLmakX
kPhKwa3fp+IgAA3UAcvcRV16TZlxFHCxMZy/G46j5tPlGz4H9bpGNpyCpkL+gj3b
g3EM52+f+mETyI3fX0CyzZ09vYVkHSRJsQyA6dUBVe6uDFgZKLD6Ya7dF/mhkBEv
3hEohV1Zhy9T4X7LNhaW83ZH3SkvAE+W4E54jniltEJLyxOJuoFdREWiZyaykXbB
oEEa6IFFnDFXnWBIA4o/WOxFQ13bpTeIjomkkM3flZCE8LonvVnbbqEVv9ThVtWT
pD1LUPT6pmPDtc9D3XBarailU99tvsHCaoGy+m0nFV8Bv3QgRc297MqLXi3yWj7p
Mepk+exv2R1GGWiPJ9Ys6LxJj9cL/BYTQgHriSGruv28GbKUwJSD4AFeJbj19ElM
DnlMPcie5JxFiEDhR/KiWU8xGOLE0cR8yI825HDjkimjFejQ0FgNiD/a0ewDExK7
F2AGE/l+/hj1ORNxlJolZDcEgYDNg6NatXHK+jWtlMrrQ670JUs6zHD2BpHkd/fq
0Bu5iwYc9fd8hA4ao2ETRXLZXuvcmvUM/eqzHpXP+MDI9mLypaCWeX4GoKr8OR2P
no2GPCdQfLsFyGTVvUrJ0k7DMFDwSiugwuWFb8LLQADduffGzEelG57yPXNddg/o
8Nz3CmHN8R9noo0E0VkXM/V+7fYj+pIPkI6dHFdX3lddDo+RUPxlCyGmZp58x78t
pSBsttV7rCglkhFKB0vFWDjJBMS0gssPoKbCt8qUQeQYNQa0RB3LxtYcy8mB7zGU
BsAhjTuGpbpZAKNeH05oiMNX+KSvyGBvGvKuXyEj4VXLwsC+rXHck5eZYD2mN9lD
6TYhLo83B4rSjIlCpH2fm85UMGqpDWqqCEZxVYevQ4L9GLoRh4wfbEiyeinVilJj
1C552oO5YpNOETHsizbcbUyW9IspjBF60y2de+VoVjvtQ7pyU2BnRSWPYIXgn+o5
cswXDl/G42czmdP4lCvHrKQyDxanC8kIRdJvP4NUkAPEV1HXtaYsDhXEZ3bzg/SD
UgH5vHN7zxgVaEmGrL10HOVA3r1H/ri2pmn472HXYInuKKKG7+hiqiqe0hjeRtri
vaqhhejiljkn8w4dZ4JHIiK3scvgjI85iNCF6L8ZhzGWbIdN1pGni2z6TNU7wNR7
NzySfCzD3bT7THRm9suy49Yt2UUA6UEP3E5S4KLXW75m39yVDrksYUcOh9nxd1yq
+yibUOI8UQoCfnpypDL7ZLR3w1hz8WOnuspJ3fbV6UA8AVhSXj00zzvUo9QWuA4V
JqcOiJp4gcvoDodmBp63k5FCH/BkKGqYQNO+4GSoQzFgSkauBHDOovorLm9n1KCa
7MGIYE77pw4iOLyoj3tJ/NwLRX94clm09a/Q5uFNw6CWDxtdfDLaNzp+Xwcx6dTK
xkcaHCpGJk6lsEDnRboKrQBEyXgnI/fkii5XIyL7oKztL6DVqlAJUqEqgaDT/FBL
Zx44mZhXDg777G+Kqlfe98l4jP4EzAkegIY4mjSWTC8pOxXibW0DFTrwzgioj8Ad
H8B/O/N11TW9BQr/RHyCdD/e6Qr+9PPTfZgHbeqO38ppeclyaPqbydxIVcqCsLAC
DI5aObGtsbeDyEw1rPO8G86KZJ+uCFJzhIzwUWLFPpifq4vI6UKAOpLppU8RooH7
FoDaK1Kr2weO4gm7RnBCOqcWNt7E62FC6/N6MoEVeqTTMLtqqaoz60cc1Fc19LYU
L6ktYHDcAFg6f1d60uVljFRdcn4GM/NxBBTe8Nra98V6BrYDbFiBScS+9XonHua5
rYCgGV/LoEfS9oE7+3aUrEajOcQGah0TfNuT4mldPOShBJeiISd9Wfb1dx9GPdth
mvP5yapzdkeCjnA6Z56Yy2habQzDeVFygDfkzPg7A7RLCQRBCVKBmjsWsJ+XykLe
F281CQ5CUbsoMXjj/iJ+APnpIEYcDW15UrBohZaOJGPGZHZqWGg8LvqI921q2UiK
h0liv8b7wwKmXnemJS6D9dXZY6VkmnSKJ93IkRSdWLZfoXDdqJOBiXNegpB58twK
6diWQ4+bAjJYkYygThP8CCoPeN8/MjpDqtbIJB8J5Xu3D/JUdqSoUCBy+GFcIf23
agBkz7wH6enYKsL/hCyJgm0q3JgXTPTNEBDw9rKq3BHwhix+ZUwlKWM/lZEOqqEw
NS947t8xjXUlbofNFOBKWjnJVb+8Rs3uESj9LTseC/bq46ufSYJ6z5RkxRUybIia
NTlBra59Rvb00Tb1TI5UJEuJV2LAsGGtIQjqQyykxxCiE4b+cJBETL1MGaDpMNRe
JtjHVVvpGfsy0K6jpe+p1o6LJSmu9a8KhoplVYWtF1J43X3ueu2WVSUwo0t4YUba
Sjep/HhqwUVisWNrS/2d71cEI35D1R2qc+kJ+CO63Nf8e76iepAJQbFXBCl1r04y
Q/Fnq7h3c3D6tvWgw/IRiKN6t4o/h8ul5JV0mHsidmGrdbvN8m8ECc6Db85+Td2U
rd/Cbg+TufCZZ9GfG81LOX9odAK8SKaCjGZ/6NA2amgr3PKSahL6GlrEZDH91DPA
3GQ+LhxbeG18+iMSb3MRQb/AWQZOZmrq6qWmSAAMRANmBYUCY/QG7p6Fw8j5UBb2
eST0Q3WQC3voS+Cfh8dhbr540cMW/AZ2FOUiWV7m2tlCswRHSSRezkoCJ91b7KKu
F+5od4MNzsCEXLe711T1B0SLHJTNhOB/m8IxW+6zly84pAiZ7Tbt8CkzG3peWBzq
GPM+CuzFG/tPoMCorIw4vGBXCUXQtH9sUlBWZm64rWRFBNKsQESQYtRj9OF9yIkD
zPSDnnrLAFwe+YLR7/sJ8m/1vdOORu8LRNEztCPh2Ydm7AwyjX3OFunhOo9NI5U/
ewfUcHSLYd6+17rqiEG0isNh78l3cmJrVXA7hBJNTJe4cXsrgPApEJlydE8bBD4i
z/rA1X7P4QgFDFQiGpE66OVAvrNbKRxKYoTx2RxVV1p0LM2NPt6y/pgKgIqf8MBD
adOsFMG3RyUhXiSBYikoe/BIby2HUoBk7l3gOJdh+sUKxHXH94nA89Hf1pvlfyAx
DkLDihpVUEqrkpf9QNY/uG/TAkJb4SwdnsC0zddljnD3iIPfIhgKvjq7B0bJl3HF
lgNfrhM4g96YlF2Hbk+RB0psY5d6dEQjqDwbvsmlD0jpYO4T8RirR5xY/SXpYU/W
nP4kJC9ZvpGgVhRwEKPEUFurNEGhQ2XoXqrnHyZrCRY+qeahF96H/a4QKekfi95i
jKZDOcVBoAtAcKy1+yjntIeQbt1KOqcEV3gfC3EIvGXn//8hB9wDzW2xGr0/Vl2v
26JIO12bHz26UPLquGKmOfigypzyWvOWSf9yPBBSh7lWePd95dawIdQXxAZG7u4Y
NdAMkfYKancwR3OFmx+T66mmnbJQekc37wYAbr/piQniqpNIwtZbWDFDR82r4AqU
KBOrht+48SvmrmlCmMdg0QCd6vx2NozHr0BQTCcSiRwh7J0p5aJpimHf5bsgw6OZ
7AcWYM5zLx+DcsTLEKppMqI/SQHwufbnVcD0u8BUcJyF0lrdXiFaXnJWID8i2hto
f+8pnCSag7KZ4NTiSN8+6+/O5g3ZfW1jIefDKiINbWHNAV5DWITFUteWwIO7uSu/
I71uS5DFTbeUtmCq6QvX4qWPw6qyVt/AyVAHiIaBx9hTYadMgQ6VVoM+o3ec5RCt
3OB/y03gFVz4xinzpSfVMgL8zrOgq5SJ/9fLOSdg3yM5BN1KABKTz9J0FJvNo4GV
0SzukJl/f43tXgmKUEUmemwHRDWk80XtlhYGSWTbZ9/irkwvMgxmdrcs0G/VHqgz
Ax0IMfdVEvXZrSsP3RItHijLVWsY6kctfCdG01buDm2FJ1Ws5Bz8by8H4HALARYH
6TDQ/re0aKytmN+2xqpk10fpTf9HAhv6THbEZUGksOmGUbM7SzhA7b5dYsqdqpOr
dYDVpoizzjawmxqlFgTWAydtHCD0jtfrWIU3I5bcX0tq29vGs4CLfHWHiaRAsD4l
Am5zA+7XbY1c+6Z2yCndbWQl/jJGLatxM9PwPU1Mqeo2hJXohneJENIBoZF4Heh0
7Lgtu5292NNhZlnFPbrQjpJUCFUK1y9md9Ebrj6lOlzq5dv97+Ypx1BOfmGjVu6E
Vo7hk4WCoiA6VteH/oj7nYPDo0QiNGm8e+xyaT3bHBSF+EKrY+u/+oXZucONsWoJ
ILmVu0K1k2sfTKCDo7jnhPBTEhRZeluSuy06Cl/jRXooof8W6tQIsCnUSC6OwkGS
dFTKOmisJkRqcGCN5Y9oLZNhq/7fm6PpbEMhK8FThcSYtxf/eypYHoTa3WlyRO4p
cBk9DOV4TRWAHSXAk0ASBNwR45dfVL2ahHY7tqLW0dqh8eg0QLjqWVB4NReV0FX7
AF7/ir/z3eQ85iRdt5pCf8fje20Ao5qPKOlcAizXNA+oxKltA1A4SqNUUDFOsbtP
j0ds8cjU/sH1EFgTZtIN5H2YnNCD/r3jwwpi4I1nLxCzzU3ecQTx2HKVEljIEpz1
4kAtffjQ6s1Y0JahKJWDG3YaDPjb/eIG08RmyWPkqcH1I4xnKuOnvIjjFpdLiJRD
R0jLW3+gJQszqrhVP/B3TEz2fO1gKblCV8Vwsqd3F4+f3XENdijmRgBqf64Y0C/V
BSrqRI9QDKlkKExOX1g1wT9t+7gEp0FyM0/SJru4axreo2pVfOTcdfqQjVs+byxO
8i/dNVoKAp/zv+toVS7lh3Bx7G85077IZqIW8aeHuTzOCvDvcqOyZYrbXEmLuXlg
DD5LhfrWfVoB5yRcw6lo3B2iac6mWdQScQhWHNqk7JDCOg5Iil8ugBhyi9Dk6lyJ
4r7dYujo3XXzi/NX9pmyW9+JVfoo2Bt3Jzkp3a9pM04Pq8xnNvZzLN75RugmBFEQ
ZQBOOsSF1/FONG8XLt7VXb2pqFDuvGtQPWuyVCTB7GrO2eFkm+iT5tdOEd1PdDS7
N955H+SYSdpa/UxccOmjbJ+uKOABzH1CiYAT9crNPrikH0R30I0f2OgitK/hecpS
Qzl+DHR3mb3HsKQckktRB0D8yJfw/JkyMbcySIkTa8ydixX67hzZF/pHqIDHwnjU
toQJuqJmz2NvhaxAnGYgfZR1D8YlRRCDurob8DxTTrrNFEXq4wglWxjGhdToVPFR
pmolRGYKvyOYaVCMlBdS+gDsgB2sob/kA/OC3JzHMtEii5Y/0ej3jsYFh0yGAP3j
86hezEq9NVvEZ0MpZabom0F1OvU9fAnrFuY9sM/9ADmhC+gHm19Gw3adYI261RNa
XC9zle74YsfN6jdG9gS7yE/UlLO8QheNK8+sWL4EvVbq3mGFAKxuPA/MDKJv+EPc
uVc8rVvI2Q6pNq/vv9uuHD+aHY0JhCXSH9bxx4ng3MgrzeZMrqiOA9lZWRBq1TOj
SD8mDQbwrHBJz0hYI2l7FJMmnqejtskFe7bhR2L8/tO1CRvv/AOcgBGCRIgxUXCA
7NGhq/25U+2ZveBTWDRLooGYYcmoUdN+mCH98Q7soUiyiLRftXhu1ixwhQTZ6OUa
2X6YdUC9m5BbUWoE1bRbFiXNGMIEOPRxkdXUDARYfptbVMszEdfcKfJoRju4TFx/
fN5xUIlKp+QmJ4PWFPE84RWDWFkW82f5iScsfH5ATAHDzl8UrxUvj45kS3xKryTP
gTKYvssmdG6aXgi2C9TeM3AaI2tTAYK2c9Y4/bBgWaW6YLECGpj+w9FRBoAoT9mM
gCKAaubWI1YoTlD+DoinBSMbaHaOjw7TO2FqR6LXWi91DpfBFqQGc5k+GreMEQ4i
iNILbDbjKGE0S78sBE7JwpVl2I/QiUU6bmgcObxRxuVTJnRIlgA+jpfdM4MbebCA
Emmint44uk8yBEijzFhCKzX3APt6f0twLZl0oCfAGtNS4hpKmP1N/TteHUeRcCf0
vBYcb+aYY+zItSeyqd8FeNes/l2LWV419I4s8tdpKvaqI30j+F25o3R9AmPxafXn
bdmhA+auaKO9QdBCvg+hWtohmlZ5hbhCLKvn3lSOyz5LHUGR0itOD7L2RXf4VY5a
YkPGGt/qRINHysFriwwyUdFHZjLosewu3JWiutZAdT6w2cVT97h5z++xYR4eLe6j
r5NSX0x2KtV00dY3yt7liSDDDq0uTvUaRc14mXq+vEf1YKE3c9oQkVcWEoM6XeCB
cprZzhW3cznDpE5NEYMWOqy+DAyWzCuPsRHwghcc9uyNEVbPT2MC3qRVoL5s/fyg
+gksIcBcDCcWJagVb1MVyZEHhlgBgr1dtALjKS4ZSoxT3QgFqYK6Qi5ThLAxKrRA
DEIKyh23RWd6xJgC6X8yXCWO6G1mYdlFSHG25VUiGt4tQV7HZH33gN3tgenllE8O
81OTYYbA6qONXlvjhMGsBRS9nPGzJh6STg59vSXrRsy7Xu4GykzOAXenz4GHmIL7
DKv/QFaJ2GhFMJoFSd6CvLrm2y5li1scM5AgNxYk3N25L+sqdjrZW/Xak8uoACA1
QHVATg3WSXhP6QNr71a90maaDamfEesxDZ/fx219eIBecvoUqDrJJ29iAjoGB7pg
1VzB9IDmKrMA1vH1p1Odu7iIadazXRn/1IbCXF+lJ4Ujw4ipR6V96hv6D7SuarSq
xjKrasdnwFNsnKcsmEkVxtsBKcVw3AEKoeA0IeV3oh0lXPWPyDWsLsD1y+gRgE8U
bWWoz96cYVScsstX3rAmzchVVNkxNhtrw0GzBDR+abD4JTw3D3dTacu4Qk/7VxLi
/EDDGIBlMA2L0br+Ch1+1WNfRwji73xm+DofO8rwo3DpGsaNSYHzymVIKLlq5LcD
CFzsjmTmFE3RlQPzXyQUzI+k/7OpVjOXrpsIpbYlnp5GKmsHWWwLMcPyrYHLPQc2
J/d8ggcaWYjVrxwUZIyRhrjyA3PXJ7qj3wUuNj09p/UnQcm9T1JJiJqv88h2hmmi
Uwrf1as+W0VzFLv/RALAphuEQgE0u7q/UJ44YM5sa09NlmJqZhOwLW8kQ1OBw5uw
GjfbYNn2u/ZnwMd6ynkJHDkwVAGDI18MkRbCdUvQhdljm5zO7z5/j9QsKRUhYSla
mEnpRyk9FR3T5gNKqmqMZosiRMJ+t/F9FVRmyuj5hiXCyCn3/c4ph5VBjo907Aun
eyImxC99GbtlOYyu6S1ijpGYeIWSh1qG7o1cqmHojyF5OiZp2u2PlM2W8YwCzom8
QQp2UnVRhKrSu5jZOq3t2WSeM55wADRyPEIZ/WRF4tA8871kJDbu3TRrpmE9ppkE
e7oI67uZtv1PiV/v+ZLpAaIjH2b7sN9JsAvUsT1OD4gSy8G+/kgIKEt1vAXtdQVC
clWVpuYs/6E5qvXikArq46i1LJ+36t07+QJtWoPS180ayk1UWCRjSO18oi8lvKUY
Iix6wlI3YGopVa4kbZvx2faPzY95rnmw8ZhNVY6YIW9wAJO871x5x20pvGbdqdV0
3p8QqS2r8Z4vc4ZojwonuFYnnzWvce6Lj2CUg2X7R+4VeN8jj+eGvUVhXUhRDzWz
40uGJt0O3IwwcmkJFfOlTwyEVh/Noo5u4lFm1BHLMa9RVvwPWc0sJ5Ey49iRdf1o
uNwKEqBWFNU84b1Tk2gBluB+hZ8MfIGwc6TwJW+IKm0TqiiIBkM24w+rq7uHX7oY
J21E0FDLX1mE+iLqYnar6xA4TZC5SWqvGjuODo37AVEIr+gEP2MT43mLQJKRzbQI
jDC6MWZGnmsNsKTd+lIRWUtzew5F7YOYlSsGYkJM8pJyElw+jwkCebR29xI+Rxzt
KsNLaUtm29SxxOVF+ad1gqtvRcFozSOOFitYlRZj+6ZRvWCnzoamrPmRJphqObtw
CNW3MvyQHnsWtEqJHyN6GyWihagIwFQa7IWihgD4NdeCGbIQ+dNLD7DeeR1Re2TV
2C2B6L2mr1zOcQUTIsu6zrI6z/GD+5zWJSNEEoCFKQ3Yz290b66V0jNC024Y1hdQ
7N6Bvgf3KiBWaCHiL2hcsIJGoqebP5ZujsEakYuNA7mCwwm3DQeM/GrWVhoM+zH8
0AgzrUL1DJdXJhx/R3SIgy3H6+ajGHWDIJazuRKtS5SfM4fvZV0eOk8zfTjZ8aee
REN1axIKZlRlsOcLp7jjLsy58ZYl+MwoW/wyJ/vpsXonpWCzdOjJdKxW5b8lex9Y
5I8Rj65PnXB/zlEGkIU741y/KAjmCojkv//6TNScnibVoJhpRe4Pv0N5Lmt7H2Sj
vtOu06zgkIs7LtokhC2X8TsIEFND/LvqdOztE9MqQotaDquzIQjpEDWnQaqrSNoP
q4EBzNkyEhejBpCxSAscisXnfiGz3s7y/hrah9cIaSxlxQfVV/lrWFtmsLC45TkY
4haCW7IhFYPx1Vbn5EvrPV8LzTRVjl11C+oWyJS+BAa4cjDl/F3Z1igb278u7gtq
FLzL1yHnXjm8vfxrE4STtYKIxmtfaYE4+ZiBVbct60W2D/iB0MQ1Zg86trToq+ME
77N7XUgfE5lvujn9mSC+5it70D0Q0HFL5ugFsDm0dzvlIFCr3hi0B1q5pNXV8uSK
WNcOyCmmdBPkipOGxZYeEha2qp5V59zGLC58hPtf9V/BU20yRzdN6grY9cbY1wzc
bCHZY0WTHWTAZmrZiN5qajueq1HiXQaZTMGVC3WQ0t3W7CDbf30noKMcBokXo4Wm
KGYNA4/qj3uIMbGBSG5Av1W/bQ5rRMOqtTyglB5Z7r+IFglTYiVb7lsmb4v0mUMR
zxf+UmrnClfinYSNESqhexR7f+LQU0bXcDtaC30c6F38FaVKvOMFmkAQnfu79+Bi
2vQcmkeBkVS2Yjuvh7LO1e+4/xaczjZpSFVjaR9DJxz/AQgmt8KraOyWCykJv2m1
D3herMJjHdKAL0U5LzkU9OPLLweMfWRQGl9ksVlRyHQnsmmltgRu5sHECps/NGTL
tJEeF52sGjb/pyJtMHd+lF0VRVVo+8pqee9s8A83qD0WcHZy0xVZC5n8dZosvrBN
vQy9maIqRzy7Wzwu3tk0aTEa5nTb8DA7wrcwpN0eCR74AYyzBZwzcep4qEbYIgp5
ukC5X2DR1mjYgsgWuY+DXh94GaREwMVPH+kGUU5PDyzxaH7krq71N+keX3yGfXeF
s05yyy/Xp88hg0HRxoXE7qfWBYNGFLztCMsMEKrVcDDC/WuZtgNCea0ax5XVyzJ+
PxK3EokegtgCczNbCxqnLwJSXkQ/z9xWJ1qD9Y9rOQoNHT9RtFrnvNQ21nKSOEVm
iqsKKAdAJw0zP4BzZVkOTOgKl+DjXkIr/DCofnRDjRXQWsSZWAXhfreFPveOapE+
zsMD5cICxT/c8cS3sJdUomdBAaMARlDRgRy3d2IGjZB6Uufhnwh3J7vuUlvas+ju
xwxeyABOV81rvYIQoh2hRrxPWPEqXWou++9W9ACdRatV/Hq2NJ5dDF5TIUS3wCva
B3efPnul7w7FUqP+Ebgxa/+wx2N4eZu7iivFTHJlGf2HcMEf/jmltMu+iF49srNz
r3vcKcWgv+NGvk7wj/DwSuyiBRV+WWlWLwHtD7ml3mWs4fa6TgPr5i4dteBxIRpA
IqzWimvXwaO+iE39CMkr1HiM671BwKBAH0PqUQ7G7hLJlH3YKEVOZqBmuLafhG6u
lbCZ08tLWOeiP7o6fexYtAAlgUitSMCDtXPdJyKri4EoYuGY3zIMqWioEolq4ASz
yG9OCAcZCHFeEqze18ZY2NpoFInkGcJAf0bzLXxfKRsvK+IXOhDG9BSSWsyfklm/
mAF9WdHmaU9sXnMe2HTlv5+bW9Vvoptqaavhgl9Rgta4qUwbwN+aOa8UHYuOZXo+
f4nwSP19AABgRlM4J0FX5Bg4HU7Jng3fx8ZbUpz124skDnJpxsauK/f1F2egE0qZ
06hJOqPJb9G5Ftvw/KuI4F7TPTCqqmnUyphRnD4uqbeJsYuJCCrxEtYu9oMmw1yO
gJ30erbekvpiViqlZx+m3j0Tx2NGvbWg/ykpfZp0CvJMudpLxbr4ngE7hyX7LNMW
G7y6nS8jXhR7ixV50Ff7LunWNyg9zyBX1FmV9Xxh6Jj97jC0t2Aj0nUCmsocFRf0
tAzNRb6/xusoMuRDsPBQSTeknn3tp51Zl122XqK3t/N6kD/UXeERhMOILgXgMvUU
amacKMsHvuy+MoqNRyUV+PQf5iYq3HGI0OBPi7ysa9NJfUlDgsmwqVZujAxNwLKh
tzGwQs30o3cj1M8PdnOVt5mL75BoK6F4fXl9oVc5xw4HGBCxCWEGla7CUWpEAkhm
Mi+s5xN1OYQR4T8jHd3Zpik9wweBdEZ7jrpmiSZz9QW7G77Y8/Wpy7S8DEu4GzxP
DPLmceXGYEeXh4OXYxGcs+UxssVjbhiOWZUXiJxAiwDoqC8ZeM3pAMGapjRQIyU1
njn+aKRRqL/rKkAd7vVe0SXGLJbexNmOir3KRxenImMpmG+EwQE9C+WsUfJiDhTt
fcshsR1AB9g3qnaGLmkCZGelETNjh0v5FqdRXLAJyKRCFVGPDsFoabDkWWt3SzON
b8jJAAiP7+cBiWlir7mV9XKUKFoox4dqYJ1FhK/TXnF9Md7lbioPhdEDywVWVHA+
ByXLo/DlTUQ9oNxdoayRoE9+0CIJ6qvn9K4LOEaoXniZo7OmGFY1Wdahdd0X7Gbm
it7EL1/XrX8CZQpUxHD4UYaLZMlMkvDAQly0b8h6CHwtrsT0ZVz20SALydn5o6k2
YnSlXDNX9Mk0Mo8AKwiWW0k8XcBmW8NyEEE2tNKRt5U5o7uqL0AzNvq3qkn/empb
sVU/FfbqJwDH5ndHOaFM5JoJYUm9FBoMHtAA82QVZKkMcViFVS/e2T2InBG4Wvjv
A1r09J2h0M+gBdcfpDQzDCnoM1uqmwBd/USJhaVOixS0bGI/A17uI/A84skpXxC9
Zgk9c/x/mfaLcqNJYmsV5Jkjhbs8fOQA/92KCtAaW/1PCEnAkmV7+QeK52u0N2iN
OvTfst5ivehLvVvA5MPmA+tOcOYKVK6via5LG/r+LDPC4PNzEFBlfwf/KJDmMWYD
5mL2/SpkvjySvDI85OziCMa3msno7dtDIlqFu57otPJEL9F3myACcgQ0Ghv9ivfz
CK9XocoQ6PfptHCPhnrf/8dT1NKtYiRbZiLIl93DjAdsPtkhxzfHWDH5JpoRfqu8
QMivnaMbglZuNC6NxJ8KEKkSLhNNKbW1JTVthfnY5lKkWht6etP0xt9iBEzAZjQz
L1hp+xgc9yFw9zIYkfdnNnJ3AAZa+Yax/zJpNy6AsztUBMDpCtz/MWnfyCETlqG5
U5HX7ZiunY2dlmNPxiQO/B1hZwLKofB1CRBFBhBvcPks8QvnNlWMaS2bTS2aWF8u
HNk+/qnzY9dwxL64uItsWlA5iIjCoMan6sp45T/i4C2sajocelFm8+QDVi0IX9Sl
Xu7UyPBrjHOy+u4KQANfKsVgJ4yJwKt+BBEAN/GPO4UsS876lC0+QizmpoQAo/r5
qK2EE6x4VWPlb8zcdLom0Madc+bzt0V40T7HqhK7uljQEQjuIs05hxwrozSm2zT4
RmDvZYD7F65j/W4SumhJdbhpUg1kFx727uQy6lxAJnsacRgwsHHlPPcB7sw0gl+7
wL0TrOGTvnhupki08yZLYf4WmWAHSJgCMWqiL18xsFOi4a3/tupMbGYeXAIeo/CZ
iKQEj9+6MJyr1GqmfR1cBkiDGG3+3lpbMNpJKu5AsoILhcVaDfruDJ1RxqlD1cRS
mIe8OV25pjWGciH3ww95RPAHwDskPEPEZebY75skF91CeBdu46eh/ZbgVYjr+Uil
YSorm4LvuvyRVx6B3r0yA9GnyCnTF3YhFKSheWxWtmkI3Y2/CVsWVGpsWYp3Snpt
hiQn6rOGwbWe48orr7p46S5GRWU62d0KG3UOXTjDkHL/UrxLSDV1tjnE7KUb1Bv1
rrbqB5dJm6VIiL9IZsebSHgUe8pfQlnu4Dk6G5muEXLJeksHbCtvg0tukLzVQCS0
AyvZueoZ+xtaXAjVIcaYB0GwK5EsFwgXHdcazA0QjqFSY7A+ska5U2SJIovxTcSs
yDL2HssBGncF2Cpv1Ua2MN0tCao3WvDvhzOJkQUtFGYC5v1yXCKZ95ETdRKCg8+9
dv9OZP26w2438um8l8WHo+nirGN7cuWPF4iZxt7Yycw1Kzi3uzEtH1dUy6IPNAuw
vlo+R1h6tewUGtOuISuPUpOUxcZ5LRCb8IqO5C/nH+5/UrQ7d7Daam0uKtmDMsrg
1X8+KExti26y2VGv2Z37z7lQc74WRdWpmITkaG2E0ev4bzHoPtIAkQ7KDTwlbk4j
vLhBaMNtITO3hBAjbJTUuM5wMexcEiIf2s2JWDgKQvVlRQSNOvwHHVJM8UTsBlZO
roIp5S0dvT5jNkDrhQifNORbn7h6PIMFjFfw+Z8EptqRFKNA8l9urdBYCOty7FRe
cOqmY+l5DbmUXhjC03NGMcaMxywzi19aFBwGtc71KzEid1jROUEcypceL9ChpZ1r
QN5eE38OGaQaXpwPIjlcyGRUndqSbGv96fDITQNYELNMZLsj8tHkBemjNTZfDrO5
5KbpUgcshts1LFFWOPNkC3kJN7SLYacTMM0TBu6YyC34EXIqGkM3/vYf+BuNUYo5
/dRwDztYsao/TJfAcugw/0RSP5Wcc9TrktLCtaiVuYle+wmVpHvapWcOm7hkasHG
CCS4eI+rS3N4d14bRcsU4Rr7hFKTV/PYlxNtkXvTxQ+xWoQV/whx5bSL03jeiYXO
fQcO+g2p9MfErz4IEmwwSRsKLr2BipW88eroExOCdSRTn2uuXiby+WKtTmCnzo+o
j74QwCz9eL0ZcgaUx7sSI6z2qNGHK6WJsBs/KBIpzsqHJHXFegdy4FbRhJVMRYDl
+YzVUjSTnzhTiRZUtnGuuBdZT+sXldVDC+05BPGh3SKhR7wCQAt1gOpER9/f3fiw
g5HhlT8dNbMc23uOrTpexvSJ0BDGZAAUIXTWq00yVxYOAWmO26esxaJJNw36lvpf
Dlpz2DhZNXwUwO3ce2SlPjWSly4kPPXCnr2WF8+B+dy5hyJNVqwINO3ZFyebKdUT
6kNm64u5cOWau0GKHaJwD7zPunHqlzUVbN+LIxAKw31XdrjOEvYx0tGGncTwU8FH
34820ZFIKl232/KXWB5X7Ng0Qcq4bvi4nPF4c27eA+0JTR59yrNtJ90O1ww41c9o
qlzIeWfbTgSZ7vaccn+s84/mAVFZw3yqD/ph4NqQTjRRJcYDN8jD1yROhnEe/40d
HCROCj+Wi9m0jA2WM010QSXMPPVhSGyqoIw/oiSSpPvYvRU3Aro/f2nrwPdgcmYX
tEcIibhxaFr5MMtbUr/psHF+MwKH73PSKYdAebatKAvTZTqjS9+SF49rOSL+x0B8
z/AawDm7c41Qrj+3BpP3F/LxZ/O9wcVDXCIZ2G2DWR1uV+J4MqOc1qG74KPsvs2y
B/HasHqm0nR+4TNoR+27bOR3dbIi4dIdUvEsToRYyJ0eik79pbExdwux+4iz+vNG
Lul0yfKQm+qr1ND9lzuODrsk27qmAtjobci/7ktMwqGsn/VI2a85KiNsdJdzgZVO
hJat9k3JNKiRxTBHW+eSHiLxuscb58ULVBPWRHpzDQ9nMcMvHwhGNm2jTq6XI5dk
FOSiR2ECKs6b1vh8ZE4U89nm0oktEBlwd7h7VHf5PkMHKVtAr3I3r8kLhBmqD8ot
0PBvdBx/zgluw0ImNh8l5GJOUvW5Z2LDWa4WOGKGd7D4j7qZmJmPkSzFf76IV3Q2
oYBc7pBLiv3LY+7j6S32vBm2UK2f7yZpbzGDLJ+HaVhyBWbZ7S5z9xQDcCEwtsTO
Q5gwmK73pEFWSQIl4DCD54JWo0LcW0g702x6sJF9zVcbQLJ9dvHuonRwwbG4c4Si
N1RRWRF6DpXu74WeZKoZ5P0XKLH3jav48lbIG8bHw4Zak0t1UCcwm7xOjGghw4/2
71kDf5TshGfMpZab5QwFVyEPtyZg+T0wdoYRJp/g8wul0ZMWYuTEvgC47aZYlBbM
qUjkNkNMymUxNt2Fanp34+3i9id3mvFiTaN2gYbC5m6llCL3sgBRkYTrDlug67MT
AfQIOCqgnBIZxx6L5wg8z55as1dtVgffKfS53VDUC3vVSZ6O81cjRAWEuls884Ov
clnKKLxdBhmioXBWVezSLcU2k9Yodk6cZXOmrOt8D32BFO8In3P/IjW0yDOh/OtU
o6Gc2zm+tB2WiUZVUVscbeEu2B+31spAzLlYFQ2+24MlrDvsoxJYU1650Z10Ebhj
YfzSgvcjKXCOkqaghfcHHonRJ8YupUM6f9JCHsTMWYYb4RTIiyhvuLWwQZW+8gng
9w4g0BlswVj4rdNDbQ+kGUhXOkslWLBxDCtBAoTBPV9utNhcE3yljv4dnMwEGiRo
tWTthZsSBw8/JB8wwxUhEfWg8qV7KHKBPLjk/umRdoN/osx6ne6RnP0l7fbPQi7C
b+v0twduEUiqM03LtzsgpJz52Jjw4N3BqH2okbuMo64hIGYci9JyXhDWmv+7x8vV
B3MV89kvGDArs8GIv6SDqFX06kUeenxR0mgZBYY213XWqbJXcL/E0EwwpTsUbQIP
3At+DbGmv0F+wDQk+q32Z84OByPGaY5XaQc9IBzCU9KmRgZ2fQyzD5vESQkOApOD
wTgnB39Wb7I9BQEuTYf/NM25/agA9GoqER9MB4UupcwwhP6+WglNxlByTqqdJmdc
0Ld1N5XW+mL153pMUdOlysQX9bwj58GgyE9HuR5vDanMbMOHO/pHLm/qaQkzKzhL
C5JelzlHnekQ2kbhlnBhMnjr2cyjJU9Eze7rIdYo8jNHKQnNYdbhYGWyB4DNR+WM
66FL0sFS1PNO3aqw6aMJ1LEx2nRmnpoNYbqR8ksxUNafJicd5ZNjrulx+fhiUnfi
rhQbcLA7T3P7XY9joskycxTIznslbUqS8pzojO04cGTJ/AEz+mzMvbODQBcSB/R9
24uvw96PT18mFQqH87bzvCPpeBQQOOx+WzOgakFZbdGyFiRo/n//Pk2N/BZDZC+H
OgVNvVWJRf1Rcn+QzT19UXBmCc2mgx44HSu2X05HwcHUKAVf5AFT00iIdEqmqdat
+DBdupa+IAlEi9WqC12E3Z750oHxT7DDFfK2rYBBZNDO7t7R0y0hmJL9onTuwUW5
WaPJx17Z+07/NcL37Wgze+b/dX+/+04aol/aEAilQs1isbqp+0ZLfKCeuomQDw/+
ZzeWzfPkE1D1Ut5xlAgElfvFQY96xWg+wTNMxXHBvZ9xuRXtnwGfshZdx3i+10uU
WMZKMXkd0kymu4Qxu1kDinTauD9rGDCpKxdDaVlmxJczGXj8/axsm8uCQPPtW5FL
eLoMEdQFZc5MgEJDiAzim/ZHQ9FTcUZoeDoyXa/fYNza0TbQfeslXEauaYQ0XkmI
p9ugI5iKtog9LePV3RjC/kSQdl3gYEq+j2n+irgYVY9T2GpjVinHGhTLaPnR2qRf
GGlstMDLWi0um1noqfRWiA/g2vDjTA8ZhEhwqLRo1EhfRXPCmIt809i59gArDo8R
skSGIqb/RlI1pgvFrZgc2XkjHLq6I7fM3SSB+jrhZL7vq6rCSNKTavlUCQfwV3MN
gHBNYlyqUov75XgjfhKRJf7ScMNj3aB0T5aTNZ5GoA5Vc6ns+4zfIGOyDYvC4AKV
dgnMTqVpI3KtHC3Z2UfIP4330mEJHy5ptz7sM8NLWDQPYMDSCAW4SrnxQa9HbAiO
Il8RoiUwauedgxbXH6z+fTwHVyZU7g2EAEQL0twQaXe4Rq4j8skYxjun6NQNXI2U
XVP1HTAqEozCufGUOnolwjvhSZIYoLXalf+t8sFSukvp9NqW8t2ghoVGul8AwDN1
acGjYaFYMXIHfTQNAJ7gzf7nDOFxfHq88StYeUS5gEGm+gmbvNWw01lFze526wmd
iIk2CcEWiDL19RfFOBGU8zNBC7tEHfyaRl4YOBqtaE/ZqvI9seAFuxhUY6UrkVXG
LKeEPyXKzYJwPatp/Vr7XfYypDHS24+L4Rm4fFG5TTQR4Lz9Ptp/+CtF+kSMGhwE
7Kez4rTQUlpLov8leINMyyoVCeMUhR6HaVAWaXVS0mEfWsy/51r532AWVo2T3HTO
/JbmPFiOfhXNton5C0EXA3bV5d5FuqgYVp1lTa2QnQoBCrSVvWZV3ZgiDjlJt/Gz
mUbHB76Xxeh5lvoYAT5lAgDGqwC7dlJlKjs0hWhrA4vxDd7b+Mobn0RX+nF24KCa
v4Hqx3ZzVBvuC48kFbW03Jo7+mYdA9nte4rS4KO/3pVJLYYSP9xGyf+nUp8y0u/A
G4D0PFfmo1MBv4UngMAUbBtcpcdOPij6BBkVDY4FvcT4FBQmCE/7V8uGa2pNx0qJ
+xty3LmuJZbBA101I1p5PXFCLhB1gGRtQiRz1WmbKqdVshiDHBjRsHpJEEN7GUc8
XEJzpCWgBMqDf/I6BFlGVi1WeWFQAm4PnenoBpq8rXgJ5TxY+aOjtTeiJ5AePgMZ
QSgDykveC3RIWmTB3uDciUZLZi0uAGO/bs+KFJJhbFDHQPaMSizz89uZ7eH6DhVe
PdtNoAebNJHAXlqLZsByReVIUqFPo55HzS1sI/O6l7gFOboWCCje2qYefqZijYcV
Gwy+SQ7e7gLDhYcL68OhSFPZQ7UHFLxA1KSoewAmjPvgixqKD/I/O3/ML0O4FN6+
xKsgU1ZOkZBn4yD1jssJ4XTtX241fvcRrAx4tuJuBRvmxCibbbf88QnNRVgzcqgG
523qDoLC5pCKB9EcoFb6xgwi5JbtklGp0vlrKrzggC8LOmW9B+j9ucbSnajFYAAF
beg8hffD8ofeXdcRygWToxMWyjjLle8OUaZ7WZkSZ58YtzslxWQiJZPS+fmHRWss
8mziYNvIGw5dltZyDuvmAER8wo2aVeyjhOYw2/uHxm0IL9kjnjVxqwjlccaO8Kzz
p1jDWPT/jwbszpa1lQZ5OJyDZNGrWgsBfgtdQe2Sn5E7z0WWz+BCbVifE0Ynj1ec
JU+VONdxEpfE5Ozx9uX9CLHh0Sxr1FVUwr3Iw4JaAy3liEvBP6iE+kRJQoJQnUmA
ItrLD7Fat0dqhh2QgUH5ZagvItwkG69xejYO17nImx/MrF4vjld1acDqGnYUyzlJ
MxuroFlrNuRb8rscjZtRW8AXft0ArWlbct/Z2M9ZmvSgOPFEMpV/AV8bjEyUeulh
4ouHXfDHide6xWRrxdn0DIgo4dZogZ8cU3rneWXHzmXlvZ2De3QiHuefu2dRntsj
DU4ESTDnyqJjYfLUjuXjj+ydtDE2s57DrdWfQViAohVP1NYejlYZjeqQ2S4DkfM5
ywO249I8pjOdhny/UEJGEwLwjce5SPCSGqzL/gCL1rsTxkmpMLSoy4sOEVDAa8cm
mRTZGYsSwznshH/v/ejO6mR5emOzkT46iMuZbZj/thgGHy895kKGLnu1O7BaOhgN
OzaZOjfDWS2Q1uy0BXUHA6B9u6seczyH/DOKxLwrdY3D1RKhyPY0yAHCLm5dtxqw
DwheAky9DDQ6HRP8l5e/8WNH5djBWMg0rjKGIZ4Pln9+/s7xVgh2F7etO1H5csu9
lkFyCIl5F7luH4fGsM/PxI2oO5Xbhn93BGmM7hmWyVyfgsASYLZq7LgAjxgtZ4LI
L+C0e7YbaMjWGD7csgoft71fQhmTXiwIJgBH3cUhCAnrwU7l1W/n0r1RrK/fN6sj
JGb/oKV0uxt7lsNJyhBLVH457t3V4Oir0Fc5ElWbX0TLWpw0SAhgdd7qghWD1Far
KuT7PtKzOXf5G5e5sLfbFZSQMSLR1r2nruVZf0cNJUWPE59ixdAQ9oaHhRp+QHvq
5slcDMq+QxBgcZio8zfxXvGl1LaHTvZ5WB7XRyVmyIfm9Mgqng2cxuDobJYeVOao
hhUnZhrvZvklT7TNstC0PQxA5Kvu3EmKkLYFmRwev4Lhk1RrAC1BUBkJ8yON5mQ9
Iz/5RW1NWU0RLWxLOhBR1tvb3YUmz+w93dxVSco+GcKWvC5t9x0UYkApH0SEX5At
fzkC+gn9KBIyr4rpQ2jnh9KfDueJYQ2GAwlCzs5Vr9GCQOCrunPc7plP+XZSD5l2
71fbTSNaZVd305USiqJaflsMuof3IHdwALCjY2IYhYU7u1LQ44+pHVu7UhhGZ+uM
yu5G6hPsM0umeQXcBepsmPU576/MyRUd62e0YJVk3X5vpnepIv1Qfp9oxbgRY+1n
86yZQmp7gLSeczdN0H8o3yqBnaAMu1X9lWbic3le48mjmOQK76Qo6f25D2wkn+Di
5m3pmcCt3rsQN7rMxIVpJ4MxJJqpBKlPMFllVuTF0kmSRMUub8ZPGX1Ja+sQSV58
wm1J6PrVq6aLiYrqid7D+a7xigf83XN8kBE+Ul7b/7g8lA4bmLVBWcUk+cqCpFpn
m8DFat6WNuIaZ+G3vwa771sMQfkNIcjkCPLjMe31dY2y47zpTUUsxqFqlQ26TQf9
4wGsM/063iRbSky5ZaDgIb8icx6VAWP8p/NrC4oEypG6gMoOyIIuhmg46Lvfbn8d
IMddhHEEdoLYm9dV0eqWR+HB3UhZpyjj4PawbH8zsUY6lME+ltfH47eThrPMcKtM
knWRW3s7vN+7c9+JSEMNiZZG8kFmviDr//QUUigIO7fUjRA6zbPz0BCcC1oLkaHB
Pquu13nUpYA8ULeEfKAVofF9UZSi09ulRS6iE37bYRPO0tY3LCQPBaHFzyKlV+eJ
pAvTXYuiB4QFIWkA/pVkv+vHwHBD7NCjM+NHPSpfUVG6gJpGYiHSLOVRhcN3GX/u
CpMK1zu6aBm4Lgw2WEh8Zk1yuA0yv7dWyoqEMcMTMHGT1zMBVd9af+V8GSvLLyH2
3tCFR4el+tKf2HadYAwVzpRZyAianizCcTXTCNw9/PF/G+5joCU4MukSYKuwuPb5
yKb1+oe+uzQrhdukxBzs4wLsx2juQiAHu9+UuTOXWP+ykuUPIQN3Gsfjdcz3Ekq/
yePe2oKKHdfuBd/TJ4ZP7peNZdnD4BozAN+KiN6UhluHgR4W/dhSCznpJgwtkP5D
jDu7B5F50vQ2GKoR1tQU+9pup9Djwnm3Vwc6UCztnhwkEB5rDqgy7B7ujujVxOYz
By5I0hIGHOpEG2gJozGKcHxoa6qcuLB/xUk/H85CwahMJVvylwnmVIRj1BTBCn3s
YC5w6nTeXvvZWhsK3yKXKPXQwWVScPuq29EtXj/NZx0lJBB3M+iJVCWt7Qlykm7G
mDmg741PCEdku4IfCfOAvdkpSh24ppdU99ZytWH58yhOs2xDj9WNxxYPQOCxqLLN
8N4A3IN++dLpvWmEq6dOvhLy3opRrnYZQXRaeJjJ7C4qW5+JlBEA2HQKEiTlZUVG
EJ7r05lmSQVxZIouXTE/IIR7+wfPlMCRYZ91fcPxvX3iwsrsnYPeYvOHBf5sLBo3
DdUVwu4Jl5NLKwoLkWzxrb3MKsZEJIhi+6zoHsINTJ7dYmPoahsuvsqcRmetev34
6jDHGxRbbSY+M/efhO1g4C8NVOarbgRlZQTk0zHFVJSZ4Xhm3q/qPWEqnABllpok
I45hMUxb7Wg/CKSoyUkLIVKjA7nvCAYSr5tmdUd/mLBUM31Cp/J4U+ThtxGL6tRp
DpFYCR0h60THEDJYhnKCCKOWx3OpMzmwLb8RmlwixfTXvGDwgdcYzkYDtuidM5cI
yU5mD9kI+W4WZKCnOuIjfeOu2XrIHyzG4nPKPhiIVLm/+YHel/ej9fXTZCsj0Z+p
jjoIY5f9gLJLxjvbdalJYFUP1UZG2SIrsT/rLY4UQjJ1N4ODvp2phlIXUkoi3F9D
HZB+aFfQSA3E+g3XrZEkhiMv/Bu69+LXRgQkfGXdwSb05VuniaDU7RGeHmrhhUOx
h/pKEYFGT/YBAFKeoXVxUW32Nj86uTWi0qjn0ej8y6nf1xZ7uTDLBf2ISsQlddwv
bL+NxQ3FNPB7Cs4dwHmPmhdTzXBKhw6MBZB46IBLty4sBGfCFkMRANj0rrUg0Dzt
ZUwEJsvv/V1zQKAuBTOspjcVTXwEaznqYLIolvBpcMXHnSH3mTDEuCyPKpyRYO0O
yydX9XLGfA/beTMDLL14d5AlkNr2YD3C1B8pWote4L7X/O8RBqx5aUNqr8o1nlwu
PvJp2hkkY33vlnyC6LPDQlsuaeJ9LaZpR0LrI8bILEikThtqboyuRuyyqmeo6sBn
JVytmqpGDoNIzicjwY2YL311YQFigsq5qW05V8URYNMfIMiIspirTLy8sOCDg8jv
vAPdhLG1BqHq8LfcXalfgDSio9cbkCRHAsemRBmE8Wr2fE+a1jgf9/o+s4BPjeoZ
vcM7agUSOJCcg6Zr3W2rrAqG3hveTGdHCSglCUghtPNjtAoJhdKrfT9z7NHyvfta
EfSCxX3aalTA1VqMmZVReMUGGnHVBEbleHd5Rb4NQf55ElyRi3igOKHtzhlOfnqF
OjKc0/m4PvqGhDe23fP3s5t18bKUKcnzShlfgTfGSW+rr8a5asRH6SkHuVRPKjTB
XsXEph9/Ch7rtVdXz+3CtKmxzMCxi9EstAlfeU9YtAbLjftjqbV5mqCW7F9xFtS3
evNUMZPKMrV9DDSoDyVTO7FZUOO4XFtfvWAT22eDp/5wpeVRzAlkebBZtGQ79rfh
igPum5bhhvyc6PEWml4ICR/euk3nePjweDu+p/TItSVytPVvtnQu1rJcVFnIzQ5F
hkQKOUDHc9KMI7Ew26SH0dVT/Qvtr9flaGDJbdSt0KW2IwZzE8Homstt/+ceAZmm
dU1NNkYmzx25gWyBwuayFLcIM32GXYKKRkdnAn1io22jldk0jcMGx6kbEohlhADT
9+eU15+WQ8J9KtOXjMf1DjUzKB+uItesn3TAlYZ93rvBdR8OQdabY8lXWzquxxa2
hBUkSYE1cUKC12gYuHB22wNNbwDpYADYsyPjfGtHAIBuEcQKjpCh8aDB3xznxquP
8ayVwnXSY0MlZdEIVKeoKfmOMUnUruxrLFKc0k3X9gz5A1cNis7qMnHK7b8Wd9P8
mOYncSTMjSSXbgjudppvJjs6p5+xWJHF9E37zGsWodSUXpUpXAfBiZWdR05IWvmb
67drtfXygcGgi3oefju+CH/gfo7eufgOBw4lZdqi8iyCQYx7tjUlJDjT+2LY+3aR
YGsZK7ntwhATvCeGlMIY/XepPz+d4qB5kLdssYIfruD3W65zVnFTbssx0PMp8AG7
5fOBflNVLedaztfAgRfoTYBq006Clu0QpZpkNfLDTehfqS29Vd2KSapVsdVuzCzX
/+VrN5skxngdnBEsJIK9CJZGl5oe5I/8xDLlnZaykL+uDclnw7GMWQMwVhWUrxxD
e/tYY/86NnjgUhsa5ZH7wfDtuqyg64Dl0VuA6KNrNBKgV72iIcrsVGRR19pXzBLo
45YhByP949DO4Mk7Jh/C0BtIaA7re6EPaubwvLtEMHiHH64/qOKnhjngoZL1xpE+
YR+N71lRbxfm3XgSL9iBmmht5PIg8LGjqhZ/0nbYxUHpDkBxoQk1SA/HtYGuZyHF
0HPpt66GGdkvhlmTsUmXP7FrQKzGLAMDdmjpYWJxJr/EzTRIWhmT/QjYpcwBX0mY
429HjaEof09xmYaCE/kZctvtWTpTDT/h2IpMWa+6zhgU+d8kLKQ2MBySOnyxuah4
VbLnlDzIIjTJq9Dg5JCkIbnrAn5QkQr8x+YJK9hdcx9UoxFAIMvibQ+5Y6+uwxQk
Hh8Op0X6izQYyLqaODlNpNF5khTd3jI3/sLQC9FBIgneqvxmy4MjrkUp00uMbHoF
6w1hbcDbS9uRhvdlaPNGkAru6CGtVIsVDnYyDCN6mxBN3CN/W5GGi+7IFMYsBmZp
m4K1oNZcRvyvopv1KLmRng5KfyhWs3SWYgXzyUErKdh0spNrxFQCTHp9Zmxnq1Mj
hzmk0oEQssqICd1xmz+ZHiCqK4yUU8gKCQvCeleUdvRQr2S+vxvO/5JLDLzg24U2
2GVS26yZu9lXkZM4jzPpqo5CKM+yCYC31GGIfB2bphsuH4G1NUA0R364VCzg/VZO
NZh25hOB5+S5X2lUJGuc11RgqcUS2+GJSh0Gk75tT8iVwmZmeIKTa7Vm/v0cK4IB
WsofdUG7mNjAMmkcp/IMpCcqvmXlFvFW2l8BgXTLGIwz8CIt7FIG7Bjze6jejbc0
QsU+3jh1OAC2X3zl6Cmw55d6KBH3gVyCZU12EjJ/b7P4OuLQJzAvJL3kBsWmmTtq
vG0OFW/XUZPeBqJJ1/kEOZxcnfUCGjRwzYpR93gktYarJyEFgXYwGic7yhfMGeDa
/asQnUvG7chPnc/5br10eVA6CK0HKSkIc7uuHopeGsdz7b8tpdrIkIaqFNWehhOd
JsIpgXvtyp/cQ/nYqndtJ8p/Tk9d5blVU9fOZSIbB1Va6exePQP9XN+/8EJD/HMy
Q6Jz1EkA2ka3zCbGa/1jKicm4WkLgGvUThHphqpMp/SOgtOD3PdaT/32tUi98YEf
Oxd+1I7rnoGonJOcnAWxwJCDBpwLri2ut2PTFwnMhXRL1BiwebZlyKIG8jXyU+Ba
j8Zykk439vkqqfDLG6/O1cj2BktIEPv4k6+u/tbFk/Sxn3N7bCbPcYKdIXGx/Cdl
971zFhQWAiDw7ZrA8i+/7pMlx33VncDsidSfllM5sHFPGPTiZ9rSUeBGpDBOdK2x
ed1bQpaTU8Kqi+26QSMGAVyFjK0CD/C65hvMADESMP8pK3xq/n5Cz0Jkvs5Z1v4I
BlHsmENEFML+1Qc/h62a/ZBHji4dZEJ3tKNbngfuMIoA4KZfhghXnT1oHjlyqPm0
MecPhXGsLUIbAlhoyu4vDXcYHh80/5oTEJwrhvb1FToskTadMQNAqRhbXdQyO/Gf
et/W3wnz1GD6ZtQdyZh/wqNbOmVU6jidYpJCXa7znP/46trbIa5A95k764E7XRN4
YwfDAMhxzfZeA1TjIJzpQMbSo5RGSjM0ZiOCOA+NShKUEOte1LPYOXnSqQt1dvdB
LZMAuwD2oLqBnsPSbYi/QSTZ2Kr5iEZkjfU91Y3mkFTpkZKRAscMHlgYovvfS4wI
PbGIqKATjBm/3iq40Eth3FW5gCgiF8JD95MiveQNCxDNWQ1krsuRYdvz2SStipDe
0/Ijb22gT/IcUjNZLJMZi3pEWQE4AmPZ9rAJKoXPnwep9kR2yZcEr3lQCczDx2yy
n43hUmh9DQ7QibRJa/vGS2+7JSTN+NrZKSoIKb0/MiypEFy0tRQDyLee5bfDXbzZ
UNaimoF1jhJeatnmkZ9njwXXEOo3SHUct/uDjxQ7faoz809mhQw0M8qaUrdTbm20
/sRPcx+R4mMnhzs3SU6xan+fuA8cpn7kta9o012Y2oc/bZZej/C8EBy6i3MhNL6L
ofJFsd2s7b8oAeBLvfM3LrMrw8Hve3o9WSNYULD+ewhrsTxEXKVsc2dgtg+ClnG9
Wxvj4wadB7VhvzaZLIUxYfC96MLTQ8EWfWcDwIW6uM+Ju2wgREIPmdjS4ndrnL+a
Dwod/qxgbV2TmvYJlkJTylcECj5KPeJQFiHM/SRQL9hsVJ4LyIxx0uY0EaOX+hfw
37UMT3HeB5TPj5TeHioP1okResCfCbEzvdAOSo/a4QbCedteyYviAaygqJK6qqnb
vHOi6CkYme9haIJzNg39OOVoJLY/RD2mogZVwD/qpQzQew5s3JkgI3wNc621fTuf
RAfjaUjYDOD2vCO1497xeVVxIKB3+O2jC8TcNkHYJoE3cFysfzIcEt/fNOEXlskD
tqv1WqQEvI7J9fAzlnwq0bwB7ZAkeFOk9U1CGDMHo+aUna/RRO4eRhQMpsOomm9w
F7r1P60oOuBQVRBk5fWEXEdmSBOyR3cVreFAdycjVrWqMwv+TA1lE+483+CaQWMX
cyv7xOV73DL9Ps3+XHHt+IvnquIEO7WA9rBtIzFiWPm30SU6ob6Nlgt+dWYj15oq
TA8daH/aFHNxhOjYcKrnsLbP13F9bYAPdZfGOzap6Hkh74NcRFtWmd3oGLrt4t16
2sWaIaFWGQDQvrwN2cOPuwPHZ8yQt8PPajnzPLWZW1wyb/1+rwCoFr64WUas5HoM
3Xs4oRCFWMFGvMM3I0Kpyj/uTlfBoQ5zztLZxzlSz0kg8gL+59JzCTrkzUxTJZYg
NSrTDuNkJSfTG/qeLBPDESzj7o5PNrCwfzeJ8xHZ2NTRO7G0E6tEfNYQIO3besSc
O+KAw0TbcME7/HavzIKOwF+SHIVwje9Ll+ejBU7fDnfLzhbhATzMZGA/JgcYerBa
xejWuE/Bo8kAqiv57rB3KhxWM4arbeBgPLWtjE9yzSo0tSexNUKX2wZK7Lc3sLBM
55cZmx+5SgQxjlm00euW+KPAm3tYelBH5WkabPftQcCRot6XefdLvdEp6s5EXhrG
jBoWdAKgHTCBFvmqB9EZmfOzqYhrOjjwUgLKaoANMsuZ+qNK7uadKECkSrM+ctQ5
fPAIjruUr1gwmS51oBKtE+7/tI7kyP3252e0Z2s+9AXDdZJ/yZkS/E/TNEyb+pp7
GE8A9DE4uob06aIL7kWWtrzkgtYqTApOIOKKy+Pnx891+OZXAdMtdebJ1rN6wkyg
k7GePbUrfF0ZSYLIw4WP9JUdyqPUrKTsEvIde65RlV4Iac2/uR1PUMY8v0VVQU2O
MxEebFYYGPSURmrq5NunEysCRFawAXsLIw9KU4NSCeYEiJ7hMKaaROutOVdi9jzs
MV/AK0JMo2Buq1zU1yX9Vgd7pNzuofMTEr7Ihc99HEla+61UPsBpVAP3Qy0iulhy
bqEercmpYBLZzggjvjEwRqPn+RZ1uCh6ouSKUgG3m+yIc+gLrUn+FvC35mvOmd9e
6tpXKs8dE904u7bAF5R3Jy92GUDDLlJL0eIwxTqz6eH1bYxnZNh98A7LG9v5oonR
g+JST514yZT+mCXaXPSGZJ/dduG5Gg4AGw6+xiK4gvRtoTo+d+dzBdqn1gb6Bh5k
Rjs3tWudH9V+Vx9nof6Mvuy8HJ4Nq3KHfiEIMiUUM3GW3Ixv83gQ1dIJdLs6fzDy
L9bYGsNMa8Qk3d80boyldRd/EG63nuoVgCIXuo7/Wo4c13m4/xDy20muMcZVqN1L
7C4kurgp5iNJYN0QbKHZTvCNk6UKO+kNCeXE/LSvFSXYCXALgGsYRYLZ5RoYf9QF
G/QD2//nsEUOEjaWnRRkL5DykPHFd2PVfq8Ba1zWaP9RbuDiTVqJXkMuoBBfomYt
is61LXiKwNLY0FGP6p8/aQuUga6UWUqMUYJ3PlMkQ+585j07l/4axvdy51ZMC5zD
0mBq2STzvVsxMZEVurHPsgtzCxzGEN65xgKaCf4e4Kblg7rQY6k2b70J7ms3kB6/
YXqWNnSGoZbrRSdMlmDglEzZaa9PlmqP1Awn0erqVsiHvqwwylauAufySUGoh1H7
VVi694p9azm4x+9Jf13ENGyDWBzxfMSMO+KaEb/LhVheM8wf4ibGhVkH+KM+YLJF
/BqXZTkq3GwAMY4EpOQqEdo1kd9pDr+GRLt2iiHTznqG41Xt92WAX2ovLjLtgn3F
44p1nIznp2YLge+iuqBPd8EGN8kKgvHl1rlvxkrzGqJ4aMbrhF5JtFr9uaoUe8tB
bmoP+fYXegKnvTjzh+joKrY9fLPRiBguTEeMX4e6btIXJQDxTbEYObxbA6X9r0OZ
hJeh+Gwex6awFn2c5UzfFpvzbNQ1s0XQ8y6Zi6X39iAFzmZMFsoCHAD62l5vREIz
I0uZ2t3kBjaM/eqy/hlK/lrh2IgfSW9k0SqNK8ssl1SdSCendbxbdiyywPiIMgF+
XClmmfLJO3USu1twmcnoBIqh9BdWZXt/QBrs/RL/fgt47ZBQZKQTyddzqVBinraA
bPmyQtwRwcaj/PE1zVrQypQvQi0Ymyk86Tt5tIvBJ/Ia4F+DXkBo+jsW7xoi5I26
rDStG4IsjbtrJ/LO9pNvmtJTg/A0dK1YwRoc41Ipor9bHkVSogc7knjLDtcLYmIX
d8mLZyqbDVr87bSEYQwMy+JUHxvRaIt/dclhpxvJRN8fRCIYr9VLIyIw2XY75YQJ
o2WkuCRlUyUtz/bPh/4y1AaYeTTFKGjLu/DU1yEsSLJERyXCT30I/U2VDtZVGFaG
nJRDbquwkdmcgJuAuQL5PQcjuBScQcXNENRVq/hrkkPTd5rMjVyG+UcTjnlEXhHq
jHpoI3Gzu4G0oxqgojUed06MnaKy3BMlSVECI3+CqvrYJdkEnvkSxnWD+IbKevSm
8JrY5QaIE4c/gdysHfLBaWuLvPNWquRLqwERl+ZfvMI5FE83uJYmB0VQDEuURyvc
q49vaTGgjQ/BDL7e9jniyw8bVSe1B+vwVLiOHN1Hill9jGsT30PHuOxx2iykaTIQ
lnafUDsA179l+lvAGxaCG/19NSBtwSlemJlS2QJ9/FyyJ+abD7g4KsaQsAl5o3bp
TxmQVGKK5Ah5HE5nLLsIwCeR9Nj3GsHJXSwhgc0kBycVw78RXJ93VmBCb8ozpOE7
kRE6dqCuUfdxy156BJlCor3DF5tKj3cUT7yzKtxY6sr5aackWBEUmA79TXjK6QuT
TwgBvSblzg8lNmbHIcHxzt70FTwXUd0RIw/BQw3QUdOjttwEh2jmgbucVdAIHf3f
NyrLA27MzvqZkLx6zEmW7SGkOm2LukfPaIPa4TDrF2Ui1SneNC7onKVAYpmZfLSv
jB7wT3v/JUWOLEWz3D5dd73O9uVAp7MlRh5w4X//f5l040F/jhAeygLH8BsWaJh4
KjvAVyIitkCjdjhQ7/bclWFERNFpNzRPC8g8AdkfnMtIX/qnCY7BAoPV45cM4wyr
eaToPR3d/4HVrMk1OuuNUEEw5GnzAQS/kOPzbKJpnJzpnN2ADUyoqLpE92xpAik3
zThQ4F4C4sPkMQJCdbX4iMR6+NqT9Qg2XzBGKHSHfeeBuSCjzwzsogQnbWL6n2Rb
0oyYiiuEnciQu89C0tIvZtPZsps5oQq1KZq2JSNzLD8SonsqLw0XmrRR6CVQuEmP
dBGZOet9LyQbo56G+sGQbJQw9J7rs6U+LLypRgm2Dhb48d6iexQfSmSJoo3R2SzD
YYK1owvPF0EhDdA6h8oP1nVXhs0eDendTLu2mzciH8ykrDVyldV8sKSNGy7lkZlH
hEe8yzQpXEKnhgFf7ng+k/OaBvd4ntD0yGspzeo+V35d1fYii2f1LnqKdwvknsnp
biqxoTZQ1U4ckstcXDnLyALYP3iEKHeYksNvdSEiEmazpl2NFqJxFUteViyVwakY
hWdkzmFbkRJ9drSSsO2IRoQPykPrp5J6nSyRoU8kEOf9r7g6PT/zxlLsVXNCjAzl
8NlXQC/SVWoeL+f54ko36299Hg5VwmK6rf/Mol+p0rS3XDiVnHwOvTiE+dYelDyH
Im6CDUNNz+/JY633W+j2sbdwwCWUbhanuI6R72xCO2P1918baWHcX31FOkG3+E0f
UigW7zRsE2gIAd0h4USRNpVlQ2wjbCdrEGSQSRMTjTm3mebx1nDt0gdJ975OmTG/
ywHy9ovN2u9AS4v4/7a0s2ecnL/WasCAVrroeUlYpaK97+3oxRZ/MUT/NVt+jP4n
w7P71dXhG78vkjeieYq+yjS2WY5AusPlxjVCCmadzJtfiu9d+0DgZ30k3kuJAytE
5xd88Z7JdymE3kBIn4SRqEi+vSyt+nRKMs8q+lUH+tnNOgxTe4AvvhZMBeJ5kStG
90heWovwXiaUYWD95KJz8GHQnTkrIeojUFp4KdiKZH/j/0eBQUxQLdUiAzzQFO2U
KIjegY7jn9P/DA3d1+2wIdUBXX/N5oL1riB0n9OWnWUTxPkeF9ZDCagN5Icx9OIt
n6eBpHhsgvr4d/4AaNX5mhjJj9IhaiU2IDDUd4DP2oXesjTYLCqlR3cJKsivWDPc
AXS5A4uDunO8o8iFdqwD5aq8jwKcH0pNquQP2YAS+EEZUKDu1XVlxB/6Srzeldyt
M3cIJKpJ/0gsaVs1SfKYWvcwkP8d7xbLgpgnLrqPaPS/Lf4q2m6y1vld3Chww1Ac
kS6Fq7TJIgWMQ0piD72GdxXX1oFXtfUPISLYKPHhdE+Z0C+HrFiy0EsLo1DGhV8F
i1ktYuXj70L/0iIZxhJ/mTWfpMJvS8cSMS8uHBkW1D39eLe62at2dMd9hxGtc8Md
tc7bcoKT7VtXghTeim/l+a+As4EfEn137wLZ9ZhKfBbvfqx+YzvbTuBJKDRdodY9
+z/HJ9BchDfFcxMyLMNuFd1bWcZ+G18MXF4RbFVbOkIKO9NaRFNdmjEYb/kpUfu7
CJZ6MwprLxLTYl8Q6nJ9uTp/s5aiLLbtj1E8g61SL4HKvlLyRRezVuk08/nXKogB
hH9R8NvewefblEq17FsT8/jW5MRhsHh8zo1yeQagE2hk2NyV9T4L2yMPc88OhOe5
lnTLXCpfb0iFRydOO4vUGTKyvfrqhwvEwr0cA0j/sfvx8nppc2u21+GLA56MDvju
EpQzgRJ+kpWPfzfLk+MMm7ga02mSfxig5M+huvm51M4NPgo4PxEsgfNFni/oZcRc
g8nnf9SNfU8DTbUPZI7TqNyckzmIrp1VLEr8yex72+TVkyeU4y6/QMPrLfjD2BvI
+8HyUQkXW+3h+XnATXLmJAEd1j/z8Nr52rhZNpSHJbgk2gBWgG1i4FfdjaD+DgKK
GNkMGaO+JJyYuC+7PRqzqVr4GoLGg3D6gwvaL1e7gOyWY8kDEJJNkbnT5SOFpbop
L98+MpZG/AxgPtcMEH4oNnNQ5el5tFZtqzdvLI8RVW2XokKHQbvelibOSfB0rskg
Lq+rEWcrcH/kWGetIrQ3/AbrgdrROor1rYMEUt8poUeIWXoqyfTe1KQD60jwGCzl
CcvtccD56PMGCyb0rPmH5nlNkG94AiESboTY/kdak8MmypwP1CSKyqWaV1AnLzR4
OuH/r5U2Sc2VCoufPyAGLR9J8jrxsJQIsX2TkcbwzVLcYNTEN/GdYS8LLqFF+k5d
cWB+IkYQayAwOBzipkhtGIktykToJBdXx6hOQ0pzdx23V363Kt7RfEo4i3AyFv8d
vm36IvHEqYAoYQOPQLVYtVMm65Fd0tKM+MiOCOEn9I1F7Za5wfIjVM2zmzfF6JfM
NgyzUwgK3tDe/qEfrAnysiVP2C6rMwgX1gYwAqBfHKCd6il5Bm62gj1xpjZfTCsl
XSB5rnmr+tsIXmy9U6giUQGNIxASU0ux9jCDsySCOUqsWfWvEH+BaPQWB9t/2esq
prz/SXVM5MGPX9Q2Enhd822IMzI5Sct24K9HzfdYCmn541zDOZ/7xDb5lWhSoFE8
ITWhB9rsYx/c75gN8XMU1dfw2SZGPeppnxjtAqxUdANF5v+CdVzYK3BQ/jOkuZVM
vh6Ozgkvv2YSD0cYnS0dN5dmew4fYrZzP2PB+SRWWHUjfhrJRdj/ERIHPZG5z3i6
G8HxXZZPk1HHwEYIrp3i2xb2lv2VjlxbN9pAjFRU9wKRGmyI3D0fzkegW2DKr1L2
HPo0MH4Qsv6unUl3CY53oCvJxWAHdCrgPkQUEak4k92ElGPW91lOoPY8riStcSFz
ul6uozhaS+QrGKEV3cFQuXqvgnOt9/HZv9R0EdTT/TWmKi25Qarqb6BdMgoWI77q
F0pFe8h/nBBo0z8z82d4KNzxEPzLCKmK874EI+w0nYGQuGVOp5Rywu8jyKLR2zor
IkMZhR1s50OSXCSkfyRJl5pc4tcJ1dGgTjMCQUptfv4tMvdumnCMxm25jPKTsbJA
0vepBxV2/kKEqGASivtblfN5jRbKt+8LzeEDG6M4vKYUvWzkYzqx81BPvYoqgktz
cAWckwWx9M7IL3NgPjyJeye3+4nmY34P9cp2rs1oTHeX5j1JSXAjqnfH2jmg8ILX
hQbU2fQ95p6TuX5XOFOSRcsWPcRrQ7KnmDh8b1YdYWd/i86+J3vNOqxLjeqMezi/
j5pig+lL/HJysjsY0aB/8s99zQWcfSzp3+wPS8fj966cY0i2zlAG5xD2GlBQFdaQ
/SiYI8vm46TagWUzNiXbBGO9fqRgaRcxMY3TJnbgVb9UADuwqRkNSD5hFk0GQ691
W0b5hgkXXv4Gz58S8wwD4tpKU4y2km2zvy0zl4Tm7YptdHcsjQeYCNEMaRALh/iJ
C46AyurbG+TmwQ8IxXfKc0Xp25zNSUQW6GkoL9RoRziL0uqsj3dUIMaSlNB3enlw
IcNSQ/kxCtDrixa1rNQQlIGuxhVLU1b0TqJGQmefoXkZYK18ST/Ma890x3bKeBIW
ybF6CrYNa85dNNg00GJY5bAwWNG7VOYuPoYyKeUefpFPQBz+8dD3qOTVwXn0QBli
Yah56tJ5zfq8l5qX+q6D26VZZX3mybZ8USjl2hHsCPp4A9EV/NzJa9Wgmr3beHHi
NkQzCGWgpJ0zmO+793WZCc8OQEKTYr62Y6uTfnRttDc2f4cP6viEitkIFV7myDMX
NeECXtlbrJyRJDbGJzBoTzVXXSngltcCX3Ofoh2VWWyQKBmSflhXwNi2jV17MJRJ
EpLlGiJ6NAfydxdDwGQBtId/1rCU2w61vZR6jx6+z67/9e0EWKMdmyHT6cDzs9Qf
1Sz7SbKfjdYx1ODsgKmKW253L9Pk9SSV5mT0afYo89xQdXFijBniGB8swx0Vye4I
ITlJCwo1jU/qH9C095RWUBucgG5Z1G/aBeLxXvCku1Ro+oK3gdwQn6GoqHoIFIhx
LZeZNcGuOB9UXLWoEaQTkJyJJj1f9B/PsEx9lzDCMS3uc33v5nx7zdpdsYHhgyev
/X+1hg11eKF2zMNx7oJknCkZ8fxlEWuVM1IaEijDXrlCbjL7TID+h0pU9SKxNB/Y
nDOol0AgQceONumxU9DDYBuu54JUW06wjwZYC202xGbai8/+nhJXgFCninBEN8hM
EN/0LgbJDzjL+YvFtrSapjR3S7DQzxKXk/KYA4IFA+EB9Q/YRxVp7jny4r0IEugR
s6Acd0behQw7/bcWIWtFUYiepw2bnscfREJtumGLrmII6zdXZBDfouUvazMGUPc5
VydMXW8qo3SfrV20KWWPb8WRV5FrEpbUQHBvubF6ePEe1DWXpLdlXAozheoGQQUX
9UOT6qFMYNKtFAYbVThkSEJtPmIeRKzo51K4K+pQzeBc0SsQA78dq5xfjxcf+dyM
aThchmVfqK8ljezgLVetxWITpYTtAfyWTe69nSYQDWsBNSC2GKQV7jd+kmCfBTwd
NmGIloESI4HyPnAmhoRlJP9J216XutGOloCKjYoNe4OhP5AB+84vNd7bS+JysOcm
zlb7AvzUTf1hOKya6sOfTiWWLRaSZ2l4A1zR+6M1E7O4h7ufF+kztn9+uOe4KEGO
CHFP0c1lmy2IJoC5k1U+uu8dm1GiqELvA0AnOxlQUOSyfnCoT3j7yr8qtB8IXpDc
jCiDxd1yZkvvyt1UQ7tpg2gNLWJjHZWO2+wRQowIoX/MZJ92FurpnWpLzxGUo9LB
782M+dVM5Dj2XSdKp0r9XM9YJUKlZIQSSzSJYgP9xZG2A6NQzQWWJ53Fm3ZHXT9H
5uiU19HfaI/JeqN++7/NPxbkRC/2Fqgf6+93TyWSFDKGsU0wDnzt+7TT/gtnsCYe
MFMFBQ8Sq+1lDa2opM7cpRwHQWCn3HAKmKDpcwOO/hZxO6wYz7EbzRCdd0BwWtOt
yxyKPmkM7OxNAYprfElkxddXabrlPddOBfQRVur06m4nSkDOkqVyiVXJFXcHs29V
YaKD65xc0im9ozBdVFUkcdUK+U5er4AppdpzATNzXKvssZfOhBKEWTy8OyqWqRpp
aw4DwtOJ/fPucYcnOkMm2Wwd18Ca40V2Jst4cmSUQ2ZyZyAQCvgDgHti0dQGMUg6
xoPVmttre1Mx5B+zuAcWIAJEud74pRpy6QKNP/gaepsW2jJ3s42o3VuC+k7RyqWL
4Sj9LKVbP6k8J1H5nSKDyZdT0foE8uuylODdXIqqP/Oz88SSwgmUnnQA3JVKQtOX
4eGF/BlUmGYpimS/cnCor4abdVGihUEqhivUDKEASopL/YgrS0BsvCpXUDk0YWeY
2oJ1wjAg9W7nmsPMU6xjbhmbaEbR1NcrR71y1rUKhbyWji7z+soyCwrb3ekNGfqt
rSJXrxyBHF3iGPpbsCNh0exEFFui1mG31P5WRcD7K35YqvtMpVYVBqnJ81lgtfn5
1JXK8DkdGbN5sbuDCG0XUvA2+HTckVjyaRwhqu0+tkxdPCoaOc6YGKZIcQsgTRG8
DuFNzd3EBYV2DwIbW34E1Rm9N1xENW+W9bjpR6a6eVz0GRHmOCBl80vhO6xqnAam
mSmlHRlBBSQIPEPu6iz2sUffStpdBdRexhLMWGaKVXE8hvKL5KFxDZPBxWR+Lvpy
aJ9oNJfD9KTeqlBpZxJFFTihet4luG63DqQz/B6jcQMuztvcsIyUq5/LPmJl+AcN
Kfge4q8xohEqbO7Xti0lP2uhO+rmhZh2nBQ29Hac/Df4gJpA8t7BbCJpbWpASkCj
ZSqqbH+VNOMQcKKh/5x1fCseTh7Yag+EyXtd7rKDOyl2Y8xiLTLvz2g7FPOb5zkO
xrJYfpCboxPKMVob+AMtU/86f0b/MJgvpq154ED3mb/ARMMpKpVw9LMFyGuITnvR
CSUEA9WvmnVHrec71xnTPxBO2yASqnUuPe8kmWLLVwxEslEysR3r9d24bxVcMvRa
rzKxnrysgD9tbdf/ChfPySz0Ap9KFZXPEgM2dVmQkSwRfs+m8usr50v/7IKJxKtN
yZYlUcRqGZGHmY0lFnZQBOJUuqAgYOu7KmB62FWH7CESHNWk7lvY3h/K0+wWdsDX
VQOkscdDahnLw2MJIeEjDrDH/zr8REkCikF6x2UMhaGAmyU6GFnXhWScu10tSMOo
OX83We3ZgDkx5rrnVYgmELXtlMEFCIteeWsdlyJm3jVpiCVQN+Sfv/IQlpYFr2fT
Hr7tLLhbhg5IfIswuo97Oifi+tFk0nZ5ppUtYnPR/6G5rflBNXC8jD2mXtxMUOmr
hhebH33Jvqy7rpJ+t+imxXPESepaeZiRjIV94L2EoDBKPEfPBrU8IdbM7yQaaMQD
JhMfOtmRSgtyNUrgDTsQul9gzm89xS4cMUnOSOfk4xDLzI/Dsd22EELEoQXktxPj
zWo5M6OxW91n9/FKNEeaFapX8g5sA0Gd1Hxn8qWCDK+7Kyk5eNZgAU2OyCdgL/hX
2RhBr4TZz29FjT0RGW5JwEg/WQhXRegkqNTOl+k2If0qMwEGt9dGdxZYjUTMgaph
Z2bIHEMrm55uDJL6WU9HxXU5yZza9N1jWzGwnnXHy+O2zQNcwsHpVNGU1YP1KkwS
QFxipfgYwSh6vn3KHOaYESVu7z4jX8EMUSf6XSpo1Tt/rZlSmBS9hrtaLOrradey
7x+5bCVD3SDSRdSU2E3MruQxROQcUl3L1ZCNX5pFQGBpRHZBsrRupXATNdcSxiPV
Uk1k3Ab0OSaxeyL9GurIEvoKV5bzZYnWuLAv3Vtjp5lBggny/sNRsB4OdnSe1c29
SaODFHQxSM5IxBQu3FD8abzIy8JQm4bhfXHuFhVGOUK3Htt9CADCj6UJJsjSt6Of
HplgLm6RJ/NDsf1sYzwiAKWOlJ6kJo++XsIHRRKwTlU5ZWxjT9qmVesW5xfGpsXN
XkKjgXbrLlLL5Ze978lz3XEWltiYc1Ua0iUwh1uA0wp0Y3Xj6QIJd6gdXiMeiRSi
mR3ZLDjXrfx8yrFv0olkrWLRK11BJ0RT+4wzEvZmHhoWom9mGPWYzH16kprr8AJc
DKg1qP20CDrfLp67hliRc6nyfpYM7iej7KGZVPXxceECDkCbQefjJaCHZJ3QXgMq
EdAPMt/mwXwl7K/7jlK8gnvs+uK9JFvN7a707CMNNkjzmxB8eYjrjpQXPATvCPLN
Hg0byCRAjAuEJHTOho1BJSNFqh52YrWTkCxXR/lz0UohTc/ecftXOu5uQ27aX76+
rfPibz/iUrDPevUpGv4+Vbzyc1B5bfgOG93Ddr0ynzNuiuZfJCQBiMkJgk7mLrP2
T8UGFuzwv4etkeQAmM04Ol2qDa9l97fylG2trMn3Lqq760QWlw1VnLnAGRub7I/f
AZvYaD88wlKgxkFYT/AngswjS4Xj+Kn3FEV9ndZytg5h4OAOgoIV6DSwiNpsrnNh
g6NMDUZ7AClvLNIzx+KLJzyiZYJ5oDqEU7rvUCSRe3wcNvZy4cLyieMimBy5EUqM
6gCQ+CrPXghMChrOKBnPANJW3H8t80oF5cLG73sIrf1N/Hb0vK2JXVMzHzkFrWx/
9217NPA0tV1b/mb0mHRCnBU9FVxo47KTQ261TzoB5nRwmGYomJEl9bSKAR+kpjm3
Z7YpcrwLyJ6BAzG8EvMBJm4TotZ8FDDb6CvLAvLSJ2GUlCG85woMZCKAIZYun5qy
Y2XQDjppzDfgQyrHRgcLLcroaCRgjn8svt963c5WH5g7dSHtxwxUJy4gP08gf8S7
O5hPN91VngjxkmBfEQ/0H1RCkpI1IhmMHoRiOLvEbPdFvkjsd4CR5MR3s5ZJk/g1
RphAVLNGsmKdGUi02Nj3Dj36V4KPtr4sO2vSE5ojZDY3aoZ06mPPHhsZI48lkRlZ
5etgCCXj3K78iI4gkNzeMUbkredYq7Sr0Usb1szc3gF3gQ9LRtOmN6laGEfVHI/E
Fe0wMi1uZaprxrOnZlnQnYg2nwRXFaRASuUpWlQUyKKiym2YBa/QE6zADXh2G0fe
R3HVXhqNAvlm2LoW24GMvAq7H21g7E0nreBY/AAMZVG9eG4AuoRpSNGmJo/cygwa
aAACT87J0goszVJyW/+u/d9kXo6EgDSXbhrtQe64bI3kqUshCXq8gDDncLjkQ7l9
wimIftDaVH8iVuBugdN4trWfRPGrMdB9FiLuwfSHSpYK7k2bWnTwq252GxsJ/lWh
03rUvhYCoPcZuebtukWGUvfXQ+Z5Av/1CG7ofo+styzxIKeXoEMV58ox9X1ZmiZU
l8S/3q8Stun4ZRE8jsv407PFYdJNGPqtsf2n1D7o1V8uBrq4bOF644guheg9JvEs
dQCUATqMG4Nxi3SzljnxyfkkYAsRQmx5ozleIHBdifh1nQZ3EaL6o1px5rl4mdIf
dCx5zqNuXfNIpESogvJuaB72hp/ucR36L4N5NDcMhG4cVX2SQHerYauP9rmMzYFR
0EEzS3km351VBK9EBuvD8L3P9+aemT9EP3WWMMR0KbKX++v00B+esaXbhgTCJu5m
MvUwoepB3EI8ZQP3NYcKqva0+J2Ug7FUHz2MhwZYcqHoIyRZfj20aZXzmxS54iw7
a07Mhf+kHRPaJ/KT1R9jvJiOWPJoLfeN2eq/FaXzVl2nDT6r9noDIbp1ognKy3G7
uoO24g0e1nta/v5/+JiCZVlJ2bAibpFEGRR1CywlILc5GZmyN/i8b/g4OQ4CEa+C
cSEUWsD/uS1EetpPvynSoxSUldl7TYGbu4Ual1O1JmZS9z/ccA9gicmYb4VJkK2E
VZszafha9z+/z64HzEO0j2lEglvhwbBJOqHMNFz3kbzFA3OyyyTqKZ37RoJua20/
+QkJo9TF2jr1UhmSu2sj5P7ISnGhN55PvaDLuQmVBuIq+gGzmBa1E2Q9Pnq8vTbA
Dst9JeGxZ5WBZ5KbLG+zgZyuPtpOAZg3RHVGKC7vlEfd7XRn4Nnq1iE29kGNaslt
UzXg7lMMWDrl7yLeO19zr7o5bBMCxwKEkII+dIVRi1SVGvy/1EALyWzTkgblqOgc
aaTjeLXs/bo+QuvZ7EqPwBBRSvY8W9EFPEx64MadH3dB9DapiEd4m+EHE+trAAdd
6zPEkZ4tJlbNVbbhYexKuIx5andsWb53ca6GIbRY8gSbD1Qidril410F4FtBo4xK
ZsveMraiTvQYNB2KgrJ1EwBq31i3wxyRDKMyqgBnx/s7k14BfG+UfPvd30Zoxhjx
TIELgDOquur61EnQg8sFxpXFwwByqWLr+5q0p8BvYApo+07KY/d3nu4BW4at0lO5
LC3++Lav9iB1ubD0GgM5/2iMJLAyTxanT9//KgZKYk8dTX/3+ZTC1DRCxtJW3Hgr
ssXtc0nqOhnG/kobL7P1DtveBzhpT5OHVPgn7Pz7V+niF56ndcDkFjbHWqOEFVkM
0xBhL97jF0YaUB0NwMDiRqCPBsBZBtA8nIesXYqyvpUgwnv5E+v7HK2KGsQ+wt0f
MoHi9m4aIkmpShDKQ0jClAR0nY2Cqmf8D+LE7go/3Z2MBSfUZ8QZ9/7xGNjsDAIY
NgasJQQBr0EAp4ulte7RHstTN3c4t2UpltBqTqs0/y3w8Z0ko89qfcLWD+3KpgJw
TdCHnBM2qI9+tqw26vH/3R7ykROIndOzd0XycF5qob9gKxbSy53wJUXe3ZLDKdZj
J5ZrhAy1ufvngl6bCh37wNQmWRVpdnUqyGJev8ttzRfFV11h/bW8lHjjQWSOS96o
74MmMLsZCpqmUuOGjba8kpJpHtuFqINp3+UVttOoGcd7x67tRJB5a0OfsEaY52qZ
BUMUO2HRmu94Y37l+/aL55X40tggorTopWso++2hZB2GVV4w4UnZRyO33fA4Fh6E
SQHSUzqQj339Nij+lLzEm6sara/hyP37n0nF4kqtbzjOuI+FSipSXaOnW/Qid/33
JCQo5Vry83CjY8LxLgm1c6rkOZ4w4vDd91VVOdOlO+3BqF9CYOwQeuieeUIAn6mR
tR5d2YHXC0A34JuDrfn1ZDfGTvZCqhdW1nFBL9DMMcIgd3dfUT9uCXRb34RcYGRq
mrUigVk93fvyy5G491x3I7/5L1wpBMOU3jLBUdx9+HAHRos44pWN1ISTrdAzVYLG
qRhcV/Raa/T5OYgNYKcKb6n9ILcVBfOJ5R7HV3GROiAtrK+jDIagMK4vgJ0toEBA
1Sw/sL+NFPxsCSZ+NRHU1+z770xVhwqLOocJSZM19y5XilF1T52dOnvafKU8FlVx
fzgoHExEOjw6gN5sUgwjcjF7lGaFPP8qP0V2CbBR5KbsndDBjXPGDvQzpDrjQeP/
w3RtYw5wIm8jeBKDAG+IdqxzLCZl0yhq1egf5sE4x5Tm4MXFeB3XuDvixaX+NCq3
t4UArTf0WOe0HS3UJzHkpTjyyrEJFYGmfF33hRZSe+6bTLxY22SS0dQHndB/6fQz
5fBzWZb0PnK/F0LPKOJUlb5+ylrEBoKlX+K30T7p3RiviD009ij0rMLO645Czvn1
OCWzycNmvKmVSdUnZVf8dZVPOVIf63K7vhPlWCx1j70U0h7QNhmqjxtZj6bY3mOU
PXdyctovzvN6Hwv1gRw6z2fiakUZitNIyN5R/P8LfOuWgTBu2NckcuDN7238ZqzI
FFash0vBQhzvlhOVB1M1iwWiusyBFudTcRsexziHyhHugnzMH1TxLmclXAFgQXsJ
jjTyMc1jm3WnSPT0b3nFmoJ3ZtQPxFBAREOlA7uXHM+jIw47jPzPKmwwVYWUq7SD
3SQdi6fwSnYcr67JBHCeVBF311q89m1OEoR/+cxdLSJ2NStGw0Z/Qwk8AjK6C1Ct
a+Eec8pt/zJuTVLKn9mVlfMVTdsAW0tyHGVJursquuhgLviRj0dK6fEIjCioiHGU
1hkMVI/9El6CgSGJ/14Hh6CjuByU41xGeI8d7gHnQzRmDOVx+8RFp8wp7AoMmFh5
56Nxc41jyXWrI3bmAVBCkyDGVTX8detaSUIjPqZar5CcODu0wICGdLSA8bEcS5XR
xQ7g7SGeNnZZl+6ddJj/B4Nd1PoY1bbM1c+MiQ3qOGBrwpAb0okv2313K0OAzuRY
egPHnlBMV11vYGn+W/1LFAg7+wJyTb/rITOmNNOjpRwCE4a8octblEodHljHX2XW
sSyceDD5wCEUSkOU8uPNNlx5nUGByKMKVeen5WYYjcmhqykpsxFNfKHuLwKb7u8S
HRQhgYBw9FuCFr2QQ4Wu31N8WUfrzPDA2NJqgul3CND2x2v0AD3vz33olAY4/pPs
zSs0R8yAD45e2SM8dyqxOe5FiR7Z/oR7UE8Duk28ZGYIPmwIBHSEo2RL9Xyf6G06
K2kAcjeTsyMrECOegvCtwnmqNa7v25vrgmFzEP5S2UlOz2SQ+Wv/1A7TUbI1p3r3
CVAPxeoBZaN5o+AEcuOs8xYoIy88jO3EV6zGVbWUiHN2MMgHhcsdWJkCE9u5jUtm
zr84nU3PkNZE1CiirQoaPc9SoOR9KcMj2IbWU+8Ar4Seswo9fmHRC42+QhvwMNiL
upsopXI9Geu2w39u3XEd0iZv1OwZtbotOSxlZgwMQEdSnfEGmCU4OGtGBdmRnlfb
RbLAf/MXMtAJhD0wxatEvfAiKmvNAPuUOSTJy0yX6oMOp9NcXOeEKvZT2/YE74NB
seCzuRnKFfkWGieANdakObBkuPYwQBz0E1jWJDLz2Nha6EEf1CU84JVp7bd8Dekn
kYgrGtO2CcopTTaPDRRNUFIT9dl/BNws2AK3+H22xzAxPHq2f0LsC4woXASLbiKP
zf7UxLGI4RQ9QYQ3Ad7udNPiPHf8z4Qli1vKdDIfvpiKLigFoxTjl1KSpOh+yQE9
B1TgFf2+DEtjAwD7oW4LagSLSkLD2QuK7lDEYZ3dhMKM+pVkhaoZIoJwwXnfv+sS
k5uJ3BHXilH4tl1iDPlHx9febw1fuSdchEUxSUGkbwitW8NYG4fXj8u96QOA3Vlj
NDjR4+5Y3EVjxkVKW8WP1V4PsdwTLFjii3My4U9n/3tbwvovJZQnuhz+aFdZtmzK
y7ltldNv2g9TaeKTFtBHfGQ+hMtAjp6rTErKFVX0nTKmledVg5mwIbUguD0cUAIz
+uA/hxH7/mAiIfoD0RvcxyY5+kWtColxq/7M5oLxe1C30HICwv8s5cnNCdciR046
uhzWnVNhThh2Czy90+h+lDXU5Xdvi6jL8AageOmtF6HLmgfFCmWBVSm1JlhHuXsj
eA/W9IzlTMJTuHBQXJjcLI2U3xb55pE0GU4Nz3W3pn4ON8jzLB5kulQLzBf9pKkN
krKVAzLmZrGDKJYFQCrAuy8w21jSdwEO5rGnUQCHcs7JJpZglxW8TjWYqnN2KAYK
+NU41YUWmun5dnsx6BZg5WhibdNDhQ+C8kf+PvmIJCt5KYV/0A6FYrUKVMihEFIx
Cz6rf0tXenaROVKNkGucEGXSWKHvYFjvVmciV0A+bJSFso2pG/bNAG4L/DsAhmi+
slp9iRNAeWAyt7kkWQqNEBrXfNU46O0tn6PWFKsrJYagNy14Yg+Y7i0plCp7z2dk
/pccaU3x3kCdvpcIM42IZXSO7QwYWi7GCDFfuj69/++uwvXUkrqP22y1xCghXuTk
8mnLeCyu5G9arNceoL/5lNpdgB/2nTo3hzduSnu5agEicu/N7L6RPoQtxVImcjgk
uBH3UjjGj1fZDc0hhmDcg8wEN3JxwCPEUXHWgexT4u0PSOkEODxC6RHBy8UGT1dT
6aVzng8XhsXP83U51ZxIrMM1EMLYWF6ZPcjTOLfOxHLvG5HGavomKZUZFQNAxW/g
ij1yIvRLSB8FBvllcw4OWopVF8Er/zx/gWvG6LbFPueG7e7hPwvv3tpBHtEkW49B
D1KcmoHnLAXLhnayYFDRzYm+UL6obmvqbbzHOAwylJWyyPGcUcknHgN5mI/dIfa1
mElgG6Iiwo/785JqW1BIdlTF7RTeH9WgDQUMHwVsdn12+nMh8rEWnNRj82ieYofH
epyKV25rDXJuqvv/5NT1OoGazwpJOYuU/Ha0fnSFXjOKlyb0ZAaxtQ4+p23rW9qO
u+1PekJ1tCB3lg6whPeIpkQBDfv8vVjObSweM7n9/Gcm5r47U3AfapMvt1A2JSDO
RMtfS8/DPNAuSC6j3MPHX/I5CR9xXyq2mgbH95+sdC9XhYC8cyVz7gmpx3ut9Jvw
/cQfTEyQT7/jsN50qH0nHT7hb90v/SmGPrR60CEuNbVh0nU6/bJZFaChGhMIAnaz
l+OV0MKJBz2cxHO5yfxKgKd0bS1inHgdt88uf+Hta/QIzCdu0Ac5g2niK/3i6IQF
2DacgTs91qEV7Mj8CFzkTSvICqML14aMKEa1od+Iq2aeq+cL8GmLrKThsTQ4N1gc
3tmUn+3HH1BQPW8qxdm3kskmcZnMT+RE0b088e3AsOOtW7/ERZpllUR7as7neqdD
me5UHIfOFK+z6sUbdkBrHgZ/GdTdGLv85KaAurk2oRSWOzdFOG2kfrBEpE/fKMs8
0AWIAKaa9Gj6Pj+n568N4frbk5bRufQQiRDxFeqgxk1y1IG1pIH8E9NM7sLUuwTC
3IRjeHJN6TB7Lm5AH6db7Nbt8lDRtcyC0ryu3CyOB3tw1X3B9ha2PfUHnhzZkYih
307tqFOb2BE4klFrhUBE20UK8iYvYBDmjLnVecnULmvmnfnEUDN5SAWO6tRQkcmP
Fqss3rRtFWKqS/wYU+HM1zvRx6i2NtK+OaaFl0CgjUtlAO9WjmLScuVPTmjyFw6i
kvoeecbloY2zwlo7mBvrGt42Sb8f/FI64PYLW67zN24EQnpDecIG356FPgJrL9UD
bWNPG4JUcRSPGcxBIhLUOqQiW3y1tBNBzf2wlDczfz/Jo3ZCSWomLkFEjncyu0zE
0pNIGZY8qf62cXn81icYfTzuhWcr/I1qQJIG7iavDqGV+J9bBlK4In6FiiAxD1Lm
jD+Tppa2PuGdsIWVeomFcCQO1LhusQ4VqvwzbMNztSGd+Go69N4gXK5CrghexuHI
4IC8UGjwpkmZkj/BLs+2IM6lqkpJ+P1v4aEcVEKPfdLWtyLTTkvl+TKIP2PJR6uS
csc+l+Pp1Vmng6l12QuDVcRgXFDWIxMRIRzyH1fYIJr/OguOSJ8ibHUTWDuDOxZd
vqVrl7ZA+97TRvVPkS8nSd1cAS8bNVRdcPVjL2SdX06EKrOY4uFuXgPCKrM9hxb1
rpy0sq8XNQlvSzhWi7tTVdZlsiTz3dcdXBba/FwyPNzLPi+0M/74nW7/Mtg7Cjgy
RZVekVlvD9plDEFAx4IHTewO1bUbTUtXqz8zsq3Szg6/W+RgJCx/ZsBOy4ZgLEiR
TTVvi/08G0ZM2YuCar0LzOcGe64+VXA66kTE9XLSKLGX+Iw78LOtqZD8QFjrmosx
uTgdbtTb3/lDG9oX5bIoKwAilydORXfhPa0g7oYI0u7pGRdakiwElpkYoDdo5Kt6
jUm00f+bI+7ELT6jor2NAZ6Da4GDT1b/J3Q3Dxv06BftB3046Z6n2vAbXhYGxd8+
pLOvsZx9ltDAUKB0wisIQESop9K/+GrOLq8DB8xaUqXjJg2LkymwnYPT8SUkJOxH
IY3HQs6lwlT4rdFxedxdwgiJPsDj8U0xQi7EPzQ0B3vSgYwlCc/SA6gfgdcyX+U2
anQOUmfh5zSZ569jzoDcLmV+vc/g1nJwg2ExmvgZlxP+Z0/v3WthYikZ14LBm15X
FM02pvdk0Ro9APBYimoMlYGLBjkKH31H6xZrkwvU0jxSxQrRJk9A/4rh+r6yaEzN
vHVc+I3ciO1sgNht3SgpV04Oy7gkJwAmjmsUOaXbjwIYBOtZRv5utsoES09kreWZ
98nOkZnxAZXBT1fLwmhg17uX43+YVM7UrHLumOcvntfUVIkxWRrvXMQk6tFpIqwg
CpNYWKkKxI0gQr+DfsAG73ppMWR9ONveLrkdboJGRWh0+DKsOkBipu3O15N8fXLf
UYz1GJrGYqPYF4mnBnlrakvJImOJ1glgPl2OggTf+4gfdi8BYIaCNZmTgvTF6LgC
BQsbitZIvg5L1lolitGc7dZjD0FyNAWoWMtOdvATYn9bEXVJ4i8T794WUMmhboyX
9+Ir+lrWiCdYGmGQNe72bhcxv7iwuGYrSHR4fcUSCNMuym3FbRnMblmA383Ona3k
QB2nGlaUx/ZKCnz0u9nxqIe9Rso17649ISUcnBCtFUU/5hZMOQq33b3JBWu7CQIk
sGH2HGqf8J4ROgoZ69VHx58TRLhdopXdmDT1I1XKsmJ/qPlHxEsv/NH6Xo79uQMA
KL1fQp8VZmUBljpbJ+PFls5rfuQjs5SJjB9X7BtGTOnDG8u7ieSdQDqTEtyOvW2l
9RtjZD+Bf5AHdQkpX/YK3/gRh/HueXw6sztwAOWHHoV0E2DjXsgArWjiBB7jQIRe
iD1IiUjQpsqatY0X1Y+u7ktrevC2rKXcHWLdf0vc2TPdF/C+E6UH4DP1TR0nIUal
CHcjP3dx8ltAwN59RC5C3/sfBUC3Dl+XWV6wTF0hH5uoX+L08hUQjej8DOQFshHg
yVzcRqLdfI4snoPYpHlzZhfTVapRezXPBmwJorkEFnLXtoqOIGmcSk0jp8TxWq8W
sxJ5YyCqwAA6XHKdqNQ++BChcDzYaU40EyqU8U2y316Fv2697bZGqW34uHQNmVBf
XGA78M5Sst/zynD9jEaRb8r2oKZtLITSS4RiGPyZdMNZoOgoKolIAcajtJMeuGf4
gGlRR4rEoAErxqI1c6E4F+PoI/ud5BxDc94VhsAIOoIAxEBco86Ltzxv6p5IzmOY
fHvSLWmnzn2xmQMDBi9bmzvH4BNSzT5p6Uyvcwh/Gn6zN5c9WL6yRy2HQH4di5ag
pcREM2DZaPoEn+Z6xulUUsoLhujEBxXlLZvqxJz2ueUx+rWVXDfftKAHNkz5TNUv
CkUKSfHm6dBv6Oxj/DiZ7W8T1dnLY6FBRg1zbaXPBxXqmjdYOnGxQMIYqBdDJZTh
s1qOmIoci94xaZNF229aAZrwm1jJasY7hjlRSUTNT833AQeVUbE50zoGrR6xKa8c
MJUGLmIVICbBc5M5YS0crooG0KvyOlzqAnQzCpFuuEDbiCW2Hl/IihkXrz9V1ecI
FKXib6wAw53lWXQ1/TuVok6RWMWLP9toDCwqXA2UHBKbdEeKqsMxxqOhzMJSOuiS
KqsGIt9/NASP8f8VMAfwDWAhVzNdIMPQxwcxdv5+m9K9Uwg1UoJgwYrDsOEMabpE
kB72YmWgSVGxR59hlQUdK0ZrxrOgBQHonJiz+TB2fw0Fgf0zxpsZedzmp47jSTor
VRbC+M+CKj1IvVBrzp8mygRWELUxVdl65Iz4Ji1Sc+lS2Bt495MyzEkybp24fps+
I1NKtgW+6sm4C91b8zXYkV5NxY2gGjkNBMATt/XA3P54sIsC5kl51EwgXB1If9vt
j9CkKZo0vZbRo1YJDn3+D+6O2BQjAW/cV2PzrwU317bhacszYzlVU+bopWsJqh4A
NurKJJ0d0r/W1q8t61loZF5N9YWwfyzsW/44q2BYgt3B51HDTMgV/f8e9VqgObQy
CybKQYOkpMSATamfxYZ8Jc69ptzIz5Z9a0jhALZwH9TVLJ6Uby1iZaMFf8ZSY8N/
dBChdL76RcYIAHRuSYtt6yojBfEo7le6GKWuFMA4Ab+kWJt1EHXVmej0b7+/TIfL
ytsFCv6s8g+ed9XX7L0FzYnpD4YkR8ZZz0Af27L41i4atsa+337M+O2VhyCV2Pcv
3XxEivMxKiwk20mxRKBTtcViETRVU20KIm1GAhrm1m1iiTlLjUwuBFH9iwKaJosY
JPAFaFpsDg5oJQB6GF/kXFepv+2SUTyxBk6WFamQu4qGG60enPnSdNITh0HHZf9f
0d6t9u5RHB9FksMWfhfe5yCJlQdS4IXHBlsEJNJpddeEh+RyBXgY3gL3/lOkhluf
+I3glU81u9Rf1gJIwK6a7pzeoXHSLoatkmnYHYA2LaFX3hUyGmZaWFJTA7PUHwS8
8Wc9kyK1QBQWi4uv+QS/Xkw/Oezr59GDGs+VNZnmvgg6C835Qm1kBTbMCWWA67QV
tsYNkEcSbEkOciSR6BmR4rVPrHlYZ7BH/H1B3plXgde89CDvnPg3F27E7T35gu02
Om3OeP5Uv2WsZHx83M52/x+Dd0ziOJ/Th3mKWtOJfC8UhyYqLFXGqYNr6Vkjfhh1
HmcSCce+dZrthq2uEP5H3YcuQvlTKVbAoJOFBQYZKEIci40GZCmvlVs5ueaDn2bB
4eckYtY+TvciwH1//9Zzqv59d7/GtxjgptVaQw3tslbLb9scLU0UebrNZI+X6Zsw
qC/WtxFmNYxSd99L4fUQ5W4yZHHKqgwjiQS0jInBYr+7kQVFoZZwQEpSmg8qh7A8
EvL72f5w73++6muQJgCh0GAsJ+29bD08ddEXy2bvfAinIiUES5aLq8Efm2slNSPH
0twMA/audaiAbMAzR6Nc+A21Utswrb8fh2gAPSIrKyFB0xqzIdDNI+fF+ZkV/y3+
wjHfrt6dG5nbv2ZoIe8yS5X9cf1m6xDgn9Sg0SG5+NMLdFBOYHJFm/kwpFJpAAG6
4kAKDeMTOH5KpBRithVzYQwsoUvwQbvwBRr0BOnQzezbOD1WXvXEXrWA7/H7e/Q9
QozCidybOVzctNrdVVG5ad/HThIMxfHQJBUjDFOa3A3cO4Wmvhxaxb7FIGSk1oXX
UnGm4jpwKEdBP6mO0Hm/jFD1cTneqgkevp7tR8/DK6fxGBhqomj3R3JmotdjjvOn
NU87CvVNmtt41h1NpFOYaJcK4mrlre0R4ISkCnhlJyBvyiqt6TxxaHfGK146Zrer
XjfL9ATfNEIo5jeVnguUS+BACpSWD7e+dWXFbSyvRbWFnBCXRy1VoCdMIu+PPE8c
eEYnN3aRH3Y9D2FyoNyWqFbYHlSJwiUcvqWvAIrm7ksfGZcP/gKbxseXYCb2n2eV
iZm+dgLm/+4Uxmz1coK0V81+8b2sAK1i5TUi/u1C9mEGnhhLnj0nNoLXgb+Sbf91
wGmZTxg7YtiT01SsZEX3k3wj9n6SO51BB6zzRzxJX6Kz26SLGiIN1HQWzhkZB4oF
taOsLd+JpY35FFFrYh2NS5kk5guA6F84hrDyyk6QkoqpUnzD5icPkiAqJnnXLGrV
wPBW4U2zw4GSVpG5D6j/EqlG326fChclT3cDSweqZiGZT4w0lvAJcu+zljNYXNMR
Anv6lmq9oOPwkQbJheF1y0EiqxXHhdpCBFi1/kDOFOzFoNcMG17rQM0QO1wzDXLj
Ykh3v6lhpM+utxU3qHJmxbjKsp5dtbqPwRl23KoiZtJxwqQ/FDQiw5y5EXslw5/D
hjBzPRWDuVDmYLBjxuLcXO4E6e5Z/uYaqzaXDXY4GI47C1hrLflj3wJYIhJJenIm
uCo8NHfEvPIa4nvE0vZiyrxv/67bdKXAfs5yzazdxO9OzAUl092GR0Ef6Ceft5EO
wYKSvet5Cf3gtQaQx+fILnZfGBXtiOZ0kQ0Qi8OE+nTBtruUyZWPLRMbzTr7v0c4
bIAYMGt+gv0qsLwIpqo9VYQNPWjAA4rTE1WiUaTjbtQuN97OO0e6RDWEV3db39bv
nsoIuQWV6WnXkoCUiH0XpuCG6glaAx2DjlrftuzWLMEf3NpwwFTzFJOiefMiINwl
43wj1zfWaRB1BYw1Kaj8Cin6rawBeGU477dtu6Hzp/fpKS2199ZspfalKQxBuE2y
IjnpKBEAdNrvg6jrVKFrIXqqAw4FQPx+0KufQ678rMgoPQC4ssVaJYXNLtMw0cH4
7XV1BZbEnmeY7jqDpneI0Q/LGmOE2Y7Wu8meSf/+INGT0vHj9QAwloPZDE39p1Q3
ZMQHPkbBQ/Iioa25WAwTvH4yRrBZBKI9RgWttMHetf3K9/r6AmUKBG8cW6YcTApk
GdwVGBnTRZUpzqkUegfpjzTDnwQ20YBblKGlnfQnxPhSlxhL7FYObjXmdIRs31CN
ggsKaEn1vqXTle9kwrnpPVlCKx2FHOGSjJh9rC/Axm07uN0SxDK5GXWnGlvGJfm2
euPu8iS+XFYFte1ThlGP87iPVWVwWXN4YbpVbgRB34BzETLS49H2vgdb88t/WJgn
A+HMAI1omOoW0cfimuXBJfrHK7HSEPMh3Vy7NMIgEcVdWqnNf4B/r+MM9wLV2Sg2
5CRB3Yed4Yuwjwd3EsK+SVvB3fltgewD80u6l/vSQ1a1sMQ9Ol8bQuJYXbN+JVRo
r1HuzHKDy7eP9AEZI5lK4ZdvurnG6GWR7jCMy5Y3HCpuZRjHLnEeVzuhdW2RAR9g
/VDFDDRDFAJ8y/uy59EqVBAtWtn7cXop8IDn0k7lt6jnQk6C31Xub5OkZMvLTRgo
qSBAviPA7iqB7NsXbbWuXks+b21wM9qWJfgAub82lfl/bBxCy83OW+zHjtThHkpO
jTNbVRLjGwq4UiVM666wA7jZOUZXczrlMpsdRzSPkMdRvwLA0k4U2eBeBsvpiASA
FX7sEDafqaBCLjyoWXqoqxJCIvvyd/bCFR2QOtl/QhXAHCJKSF2W45IU5KHfBKql
k/G7bMZSgYHmsWAyD5HKLh2PM2Y7Msi7e3htoz7R1CZDactomuT3WunR8X2AYVOG
XSBZaUFD0kYvQPRSd5k+JS190StDwImAoNkgmogoWnSvXUnNpl3pbFN6axi5I9Tn
HGJZlBklq04lFLGkuw/KZTgBEzwzNDvvg6qyil1QbFvJz3P0JDgHCRBuBRYOIlB3
KqsYnKuegiSVTK7JkNkyJm4byME16o0Nbk3XO75FuCRFESniHrOc2mMZ0hDeRWm4
EYR+GtTxd1kNsVzVKPpSBbjQuCUYjPIjKE9iILxYEw7IsD0Y038i7aNT9hN5sKHZ
vcoXxTqajbIv8XpTHQXKI/KJkfhs1WwcO4ov/aVAf58gIfVn8l7fNjo67VDDBLDt
gp7T8XLk+dcShsmiV+X2LM0875pkgdFvx3uOz6sRY+tzD6Jp/FU0FEEItCJav9gr
tEjhLLO52SCs9RPlRv+ILFKubQgoGOa9A2EuJX6RPBIPVHtOqLQS5+VAdOIMSAoI
lZXVQBYXBgtkYM2UlcG7tPr5yuM+ptqVHc+At38Re9K0sMkx75gdrn+SLMi24o+2
ENyBi+xUtwCDMa8VCb901UF8o/JkXVvCy8P6YEoHJPI0blmt6TObwAkzKOVvQ5zl
YVumHZ6VemEZUk7axhdwj0cw8ahoXZeryY+WYE0+wNsrDIFKAHvWk7emwBsEAmCt
TCYAqi50dVxTmS5RNZ60PVDkA/A9NoLAVyKG746HqgN1kCC7fzGMutUL+B6ES8fz
mBRD0TAw2CN3oVXCG6aetyoVld3aboSyAzrP0KgwsKT0kNvNa/fQ3akCo+SgHYaz
A62BEtin3P7o9prMOun6dozrjVbCfDw82MdLRuaFD3p+3ilTul/u5vhe3nwsAS/R
J25eLEXN91btlaHx+vgc3QFqB7gHqkINuuwSaqhaMQ+ZHepiLV1wIoQ9XtJkb0/M
l2uPAwfV3nXhcHrKJvguRa+mdMpwiOAzNmsUXy8VtqbtMaZuupSgidyYKBuK5Td5
73szTpYpMN6+0OIZOoGHmQyFBJbUsZkxI/5EiaqGjfZMnV1GN1bAwQwC1K6eERKJ
+FQ3MxOnEsZx8YuTWDQ9Le6NjE54Z2KtsAUuAXAkfMBEHRFhXTPPcfrYfIw1TFOF
IL/0CaAxwl+sEPAJwlgWtRkS+v3t6ISPw1S30S1sRWpxNHf2ffUU6UqcKVdBIjqO
187b01+yH7lSxCDbr4bLeI2LfRpMQEMelFJa9QGBODuk4H+lWcXpTuif4+RkMpdK
WuJzMDWuTgJCoX7igPbZ0OTKr4PaJqD7T1dXVuIWBTLf0yNUwHhRnTVpW7n+wFeE
O4319OZnwlkri73xCICL+4bSzHNzxfShBj+o8L02KNQkaIQAdnRuqEC7lcX7UKE/
I3rFmiqBAUywIo7i7DHP5KRZhHQha37OVZo/U0ImjzcNmX+28C9wGG21GzQq3ZKE
pI1XBsCUBTnh/oaUzMH+61UOMC5gTU6XeHb6u8Vn+qeeW9zyeuqTVydsFJqTDSqw
WVOLMTBhaGC74UQWbiBfpSWszIR56lHDgNshQw8XUmlFed/29YnHeYCKZvH7QlB3
sTA5G8loX3aDNUMVMwkN/3Pl8QR0KbQuySc0avuphxcp2iv2pTgsgM/fiiKiCBSV
d5ReJQbrYrSl9c1Y60PgY23v9Pehrhid+ecQtMExc2RMD2ppAPan7PfQTC3C20YG
lQJaiC/wdB12K+DMZ183D5LAQT95ugG4TrveD/oRgiJUIzJH5Xrz8M9rmoYxi6X0
Rx6gQDNw265hHLcVMoBKGuUIffmXD+DD8zUJHibUs1Rax69UHCp921L7wYgMIQ/D
7uocw1JBBKwloA3xCYqr0gRT7NfDctVhbY9e2Htgz/oBnoRPBXvM2ZwPHwa22r+v
VZgDcL60a70upgI/2/VfSOpyjy8OXNWfC8bW+sn5eFvdxrIZSJdJqcRsuvSv6DLp
2ZZiULrittXrhDvVcgVSr30zkMm3LXFvZHnLe1j73Mc5KX7kZa/EVc1g+CHdwWNb
4LrZIK0qSQy2hQQpQJkcQ0kq57+W0h951t2IQRuARODDqLrYuFCjFCoXDyM3yqJj
ivx75DZR7QgGbZFZkKiFPqF5100DOTbjn5g1MOQqTk0eUajBpzccDPy+WjKDpnCw
66HJqyMqwlmbXVwzHTovHv+m9Y3j1Qg8Ovscnt8RMFin2/Esjewu93UmSYwi0zbG
gSsC7o7OTb+ydWaxFNNkk4eqVXJztPP9jbln/jTmJvg0Ct983L8A1kQeAwOwCmk2
+Zy9k9sfkdQa9s67Og1KH4xEp5idCfJUqB1aHm4iIJs7JN3O2gUDITqEv/tG1L5P
6Wp/DwYIitYek4Mol2bBCMS2whrgI9nSdDykG0RuC2ln5VUVgIHDpUPEW2fXB4Fo
2ECURqV42R1VkrA2Ecjm+TSsLqa/D9lopRXuhqfvqnl4VkVAtz7tRAl+yMRIi4L+
pfYnJf4J+ENcGobIbVd2M4KqTbMQTplvc4ZWWx7SrLpDQXW+j8V0651MtanN5DXi
lfY7Z1+oK1lemQXN2rYEEuwAH3THMOELHa+rECrGiRdqYk1LJzvopHQKidEJa0PM
TMefSex99qi9hMIigBO7EQ5GtqFvZO9KwJdpFEgrEWzmEEXKgXwzQ44eI9GEtFSb
51gonjkvKZmDsM1rqOwDk905L7kab4h4AcGzFcpTiiyU+qakFaXwIbpZq/8f8r1c
UmhAahC90kK5myWtiASOErPRrgvE/INBisJ4DTZFmqfGoE6xAgJfNyV0AViQ97kW
6p63qFNm2gcb6hH3H+33rT5ex1DkrnwTHr8e3QqUe+tVfHTrV4RcQdrU5RMfzSHv
LaP+LAe9vukYiU+vyX5s6Sb+Hv2jd6yH6mrhrCaMh7lLYZjzdpXNUjRrJ0/TvvP9
opk6xeEHL5h+3eWhhs3K7b4R3+Wz5sVgshFpSFeuUSJRmJqzl4RCmIXsZIBGVSmU
6g2o5VIAJdaogvIfG86SzZ3ZXu5O7edgnxZnIboCEB5Rrm1w04jx99JOe+GRfi+R
thY8OHrNwVxR4ENR94L7brG23r49Jiwjemt09uQsVvlwJfysqze8ESkGy9XQNJ8p
HjV54rzi7e9rFcV91OAf9DVqecdYkHamDEdt99aJ7OSNML17/4b7IJ37ZUGhW+lP
vGyW5i7BhwCajFRFYqO84bHme0D9Zv14Nh7ptpNDsbv9zoZLY/njATYcbg30boip
6GF7g1zVC8mhn0u8gz2AEl/b/UC8l72uVC4tcfAjdFMOME/21Yvr0rGgNjw6NpPf
EwDkQb++WEZsqYfMNsv9ZGBLt1OBnntlrXCfktDlyFf40fE5iP/qYu8Sp1t+imxB
JaE1jO8ojuhGgkMgDAAPwQZsNPloAFVSNGiP+A4HISkYnM3NKdghXDDVcb4W04z0
TBtPLsYTEncPjhS4Um4LJXljQ0cN9YqhnI7t87u2VOVPLP9tKJub06lPGW5sXiFr
o1S/Zxq80Dp+xOfd5UC/3m/ZvodaPc84rdJAr/XqmcnfhDwy0MKpcdoigeh4RZte
ZFKh8X7vpbqkdGcv7p0FFHGEsbqtL3gY9YxsSfZQxDilU8KuA7zR38LLho88CXwr
skK3HjRzbzoXUAGpsdb7Lxoqnui4OyVEAfMJgHViv3j5YxOGB8UBd6xY7dMtdRhs
ZN7LV+Ahr1E7B9i5lo5iNBm3yLA5BA7kTHLlD6IXtsTKLKhIOXN5yub8VHAaT9ic
cudgT8pX1KP6XIiYEzZHPdHSRluCprhyoNyPKdQOU4LVxro/Oug6Hse554xEQ4Oq
ootlbH4QiCDE1TpyGx2YaU6OWV1o7rQjekspgRdtNXWXKL3DHfA+3CXNK5nOq/tc
elFR7oMVRXPQDRgvD23wp3LUAHTGfD9gMhCdgtKTjhDMvMRFLRgpaL8O8p3EmjMy
TV44iRJ28A3kneUyU2KqSIuYVb37TcnehbHz+Wy/qAr1Pa5iQRvpvrki649Ij5NT
KZeylNVrwX7dEDKpmu3Qcn9zmI4ej1ur5LHBXJB2yCxnsw6zMgLUobx2XQUjcNKh
6Iup3mdmqL1zV+vgDpQaFsJXq1IDPKfHAs3IVOxts7jvgdlk3xvWmeDARYTavB2C
Fq3kBGXRe2fOnja1WgbqMxnDm+Y1Zu40nqZgNeQuXbMGFdm2fQd21QkTIsAJCsv4
1Dm3GCnVefU1D6+A6mopCZztJjrmrOalXb20g6hU4pRPUCD+vj+89rodWrQsscuq
uUzR+NfBt93BK3kq4i5c/m4XP1ItjNNRd6EfphnG45OsitzjZKaCWVsRm44yTjIf
CxckIIWUVvOtrNJMa2BOPvD1FFG72OtiMDYlp2T4VPbBT4AAEjQuGwRwXU5XphxM
te97GqiKrF9FsslkhVZShxTQKNkOxvMb6QD2HDsqLeOfvevYI0X+JVK+NR+VHUEk
sVEMQfu3LwYw30RG+D+ysCYU26VRYzNhzbn6Fb7qelZizWe1owG1kp0UAa2Ih92U
lM86I2hU3ZIdCTbs4DDdYX2KUt+zefewFBYeU+KLwe7R+gfzQxifVngwx+Hgtw0V
6N4QKMjH8ButN33+ovUTYXCVJMDFC6fkLCnlb0dRAhFVEdDvvmfxYuR6rMdHsCJB
QJBoLvAdAp2yh9byKYJDm+uKI44CPcYWgPXQ1QdMNqrtmbHBODYbLadnIMNZ0cCO
XePVgu26lC2/siuF5VHodUXINDUY1AhgATk7x+xRfZS0lyabCVp6F8XQKNnSSpiw
Z4rzp0500CVoGbsVnZteyHRsh5EORqtPiUyidl7YNveoofEO20jBMXlIjaJZY8Om
FjWcq54Ezzvw4WQe/0jgh8UMYSVd/wr4Mv2KYE1tkc1UGUVBidjlU/aFdHouvf6j
wlOCqSA1TFGTTM8UXjMlYSk3lZS4I1t2BWEl4hsYUUNRZX3LPr8bmx7XOOvMvd7/
83uN8OjCSs3kzRBG/zj0lU7rsUcghW4T/LKvjb/g/uzKL9YlBWMwXPPFyKY2MEG9
02MxAG1/q0WNU4p6vWD4v6HeS2Hvfk0QzpU+JzfXwYvK++fdCG06YvRSoMvAsfmJ
Wn8hgXL2imySHS4vsMOsEd4wcU6Os6v8aKIL0rMBIzeUjEpC2KRYBz9nWt83cUIR
sIbdLvs8taJFygy3W4YhbaVeRrFfyu22FRBTWUL3d3/o8WQp+IKWIQzTzG4Zyo9K
o4V2cg2KwxWLqJiRjxVjlnLzqUzf6twmv+I7g9GslKiihp3RoWRz6+nzrJ5nAm0e
5IGvwTHtCctjBKLauqpaUPJEU1KIcO6eK7IN2ZliqJN0aViLLd5KL6dRwQNkHx1j
p0tasvHI18JJ88PjNfcPkjQzv3KAGX97g3nPc8zSIINR4U9WLHfLESQVe/TEG7Rc
CpY89eB7/+6YMcpE4ZwyoHPYnCNdGIMBpYu8Qi3WysqwcsNwpbPHGDCKHG0nmqMI
zRppUYUXiqKCSclCs880/RJdA1qiFsR1iQh3UX1H6Mjsb69pSVKoA8JWiXFDlr0E
pFvN9l24ZLu0kg72k9o6m2wNRpPBlWqt+3AH2QNF/6X1vTXukAdZzV/nx70h6cqA
W1N6WskGtjGNdWIspFbMgX3AZ2qWcd1LEsXaVU3JMEyMWxEzpVozcoxC3OY0O0ix
gm30cbIVH0wnqVQ2llWz/2H0NhCdh7aSUoghPOomXRHxZ4mY/fxgLGNAmBvcdzGw
TlyANa5FYHLbx81BV420mhTUG41Q25nG+gUrESksoEWEFXBQi1MTJraYiYX4XPv1
0uaGcYq6Nbzj3m3MfTmGpB2/6VmP4yVZo6YtrLdKg/tymGnxd51/8oqzJxZpkKjB
bNhRmRHtKVKyO2B1AoZRnIXBmFo9NbS3Ddg4u+ZJztS3iHRfoqt8zFx+uUvLPsyw
P4YUKqLu6+uIqkgLerQLZ5fzjY7P5nLG1KGfH7TbUlWYRtlJJ43i30KWn/q16NPG
saQiiFRlNGiMEdoywjHIfIFWAmCUYkfzZfUWC8G1vxXLzMpP6hjrflBo67nAQGUf
Zfe+IXGagjm/vbJ8+JwbCiPEd5RCV7R49W2P0Y73+q9P30gMNda86mBnpbVAwh1m
5Ub26me3AApnF/h0TymztkoAiQuDLLYNyNHgQIGnA1qpURgfcDhoXT+vw998GA0F
AVmqfkyOrepayvr1cQzAAHFW7PkQX+EG3X27yUJPZnCF0BfltvHNYrhNDVkc3ju8
GHI1lJKV21X64/SMNHT1b4zhXvyk9cDWML1xdilcMoDIisuUFW2TVVGBJzweolaN
6mSIUdG2q7KJsXPl6jmBvxCDa4hi4L/UBz4Vzf3BQ1ILtK/4ER5RfqAvjM/hZL8O
e0Uzs5m1XHepnaS+gqSX2CTk/iQuHN4UyC7N5JkEhOOv/zHZmAY5PTmewiT4KMCt
1IMM3DoF2Q2Bue2t4Tkq3pniX8JLc6mRlRM8gJWRkWCH2LLpB7/DAssu+a82uzy+
PZ5NpjMFVS2MC5hJF+/U5Q1fBMfAOIXdXe/Vmf17zTOZH3hQa4703A2KGEJ9cVgM
j3w/QeyJf5tH9etYC3anEgVJe3hFZUfzO9ECsixOSL5CSILZ6FeKETOFOobN4RuI
Mixgrp7EiRfIyIb3pRdLwoyCVQLVda9EYJlJ5bKPkXzSjfUtdUjG2WUAdP5EO0Tl
hYpr12NZbBB/OFaZpDR/fgZab552Zx3MmXgXJit5XbzQSbP+EgA5G57mBWbgKeLq
l2H+tZpGjeRDq4nOm5iAZUhvfO1fc/+Sak7aKDkQ67OwpcJhaBRyMN0jc4kVZKmK
zUEDb+Amtku3CagGDglQ8b9Pj8M5KbquD6B9cm6JpufslOHIzdr8znktrx+d7Cao
Yma/eujNWWxqpISRPmAK5le/6dlDDZyj2fFejOxfGu0SM+R/RG7a0X1yK5WADQQY
Vi7eCOAt9OFN9b8cpF4QUmSGaJgxkNKAy7rn23rrVZDadXD9Etmo5S8lT11Wa8GF
1B1Zim4iuLj5LeaxDIqDT220OI3kg67K/ymVlxEQzNz79H7gu17mlWiaeb70qxu5
7Zxe2kpo289ystEKULh5PxApbJedgsWSGbOXvLvFM8Cjg2dVjQFeuOO1kxcWGrVe
D1bPcnXwK52Md/AmVbOTEwNwjwt24qbDovYfX1rPI5+UR089iVvlhnpwiwfgairw
0m3gtrbtt+gnj6ud/N9xMt/ZQCnQTjhcBuJ6w3gvZpu7/gNe6hwSYWiFmpEZtfcw
0dUFdmI1VyrG3KIy4kCWfdOkUnKsyDv/hSt7P1ui9PqJHqmMTUcBmtzXTElPo6hP
3cPxg5stnAFvG1/jFVbVneIz8O3icP2AHg0hFkgGxzPjiMMXDxnwCCXMA45PueGw
7ws6Zin9oufA5dVIeT7APQQdsUuv4TkOULdJmRnurQZD01FfME1FNRemkw1Yay2W
6yPPjmgyyBKzNiRr8uxGXmDdqNCxjVyd0JzUoes2H/SUqQfBYZW7Qy9YFA6zPMHl
QmJzec/UshK/YvUS3czzvPVDS7xk+bv00coSZF0gFgRBcirQvN+txhdfEyiuVOBI
/w3NHS/3aqOXdbB9TWAs/1dvDtJ8YnRopJNXi5uSvQuZsAmw4qQJNDoXAN5u7+98
7bmXow57/PIMyXOG0U5f7AlF9X9eqpZeofy2mqPG0XOanYXeXPcpOD+l7wNIeg2C
sPij5gLnxIObJtf79FRU0vqmlsMYTAYLarMYWN+ce3QX5zL+aSbc7aRaWeI9+aES
6zd1mS1dpQFbz0/arSgDuDXXeD+38OUDTthe+GZamCcyoGl+MrTC/9Q+IGROAIdf
PGb4ixiz993gjalZx6hKXEea3cagIRNzkV1QvG91XcOH3QN9kWvL/CuxmKo74vSQ
MhodhHqdvaDc0Fn+UJbgMIZF1VekfSJeNzSHVFbWmI1dlstOW5OCi7sG+KiPM8A6
3V+X3eOjzzcUlwAzVypE4GwykSd0P9ArB3e22v8SzNMF8TDral6AVi6FxLx/1QVu
SpMqxqJSbDYPiuuKlG3NHL+VlaR3MnV6t1EUTCqnV+viWodWaF8O4p3Vw9QHM2jn
JA+zws5O8Sqw0IiwoL/IGNP/XpDdWozZtS562bxLdnK7oRtZ6XE2vvHf6n6Niyx6
tmKaoIurDXJjqhhmtDfExazct39Vl7gVi3GZ4mD93/M/VXRg1c4/qaIHgCfoYVkz
u2Hl0kBH7klX4NxxuCF4JV+fOLfhIv1NrdV51Q0ML90mdQO2N4zbPNmKiH2RUDhJ
zdP+IJGEruhvxiZFIbIOSk/48gED5h+HLE8+beu3fpLGQtQNbsmKOKKsIiS9CQg0
ML19Ybg1VAYcLTdQrBYW+8Q3L3o1hIxShUax8Kg53xi/PkIKcFW6/NS35h3pana/
Dh/MgJKHlzwCAm/P7TfsieMw+T80UExkAzhzv+SJJaXEzF5ZhXx2eEea2oHgrgvt
QExo+oDoV/08EoRhF1EfZga+tYLKKrzCa5jpWd/03VxUZdjZJ0+WBk1jiYeBsQxT
W3HW2MwhZkKbR/0TOYslBBu1CNHcgZLO5yUYjWxcaKgBud5xntGfmOpOvSJDFUvh
Rv3+uoaYP8XK/IIf7HUFSJWP4NbQcPGLmq9yyxXJPgME5fLUS9zWTABnaLqjoDBO
Nyb0XTb9X3vZkmUUNl5l9gF/ZtLPqQL6Hu6fjiIMG1+Dtl694/yRjB+SWcijVIwx
zyeZWTjANSjgf4M1+lRkoc/IqhIMTBRPRR3rtXFKbQYgIYWDTGW0+3kEtCYJI7hg
teWe7YY9sEm+/pdx0kF/Eb91pA3fZNoYGhmy7S55oIgQfuswvlt3tVP164EzxzOd
KVHQTa/8ExtRYSvzZOfxd37kYY6SK4D+XG9kwvWrdlCk3kf1xaTpZ015eTu3x/HP
QduI6zwOZnzmg37mqWYh5KCItp53Q21U0ZsIUeuJQhFPjsBsZB/HyxBahbICzPbB
7VgTNsom44r8Q2YNj1tDtY0nc3fVZwtVVoUVc1/fZTdIz+AX0bm/XRCTfjkw/2bb
JwBS+nq6+adQOME4zLW/ABIgQjtkNhVKxw20xtXE6CbU/l5qTCD7vLY1xDHMsPeH
Iyssk7nEMoCQhysJhGx7QYdPlz8OD+jDvJb4PdPBHKZyqARiM6yXZ0D1RN4YjHXg
7U91Kw1hRcWZeXSgnjTTZVDwpFhkKcfIwpqEKOBloGrgVTnRoXiAF+pnhR7m8Wkm
Vc2e2QRoDX73JOJUApTmCyeuTW6nQSZU8dSISzOweGOoSn70FiFjM4v9ZzBXn7DU
2/CTMf7JCKtScOwxncg2e0S687kra+Ey0fLNLmm9LTFTnInX5RuJAAnekq30febo
ZaOAa6oviGmKGf2fjCpbxDPDNAuRJ1ITPF6QnbNzHV0ia3pqQ+OYKtBGqmuK0WRa
jUheE57H1t2EQwPXulnKEKad8cmfDlRyP7NG9TYWUsFt9OsMIGAM4b00qdYM5RpK
PyEcLCI6vgxdzzixGAt1soalYV8HdZyxrWjaCOwgrETQSR8pOX/NhTnqZyfOM4Hy
m8oHW3GLCMvmI5Pl44Unf7EU3WhxDaGf+cdK8rcr8dIJQV7rD3mvcLfoocDx4JbR
Z4As++Wmrwb9X7CEU1CVyz9bFXUwkltsl01+7c1XZD8AcQa027RSxoSOOEsRcKf7
b6YNBRwimrCPUz8jTdz+Lny8Yb9clWWgqw/uHcj0EP22KrHoRZcScY6c5PNvAHUb
mH9fyjQeI/PY6xvZ4N41oHjbTgtfakjJTqaK8Ki9vgqLuzmZKOMcGHwsTikcLRiv
WxBqwr1IR2EcCOu+hsAFWN2Tj0qIl+JbxsvZ0omwGyecb3/RX4LiQ0lQP2SUhTXK
Ifi2Bo78snuqceSddGiMYjwgV7U9Y7t1EkXgSR84vhW+k/M45KYFWhLfsjOB03X2
o2puFB8WzWgjLwSP/53y74vim74/ORwki3pJDJABW4D7rS/w5rgk9EDG1/kzDYEd
c1WkmJWR4SETpVrFMknBT6xolkuvxSdw2JE3Zi3vZ/BZ8xAaXOs6hs/aRN9q9aXz
uZYWRLeR3LjQ7hedweELeVeC3F+Ut3sVNw4D8P5GVSUlmykMacjcAYUZgslQcWSB
FBb+z5HmdaP4FmErRXbaKx9EdSC5AKYVVwW2UKoZ4lxEW3KEgETkQ7N3DWBhaq9l
RAeydObvgjGDM4H0gh6GqIBkjDM/RonRdJxXeiCBcnDsYvi/0JuQ+aI6bWWQOahR
Atccbz6TbngB+wrXkHYtICPkMyNxrAIJ0VUfEd2SdS6mFInAyKLHuWJdVFGT9PK+
vi34JFNUwCUzMRFVq0SKc9Do2fLctsBHDzGJdcXHXr7rexhdIORt3Yl3482lQ8t/
VJ9INFKD6Xd4KzLPS4O4Eu3KfsT/v5wYoVvBzJ1TvgAMqzn7BzUacC72mHeo5DUM
yc5SSuf2asAzdnHhgZNbvohzkFSLmdc8yLKpdXnT6fXPTkJC4Cbu+ryV1QVmQWMN
KFsrizbcwtLF9EjEXliy29D3Q49wmAL6CiPV0ulf7K2f8CYynFemXfzzb3MIT+O3
klpxuVmIEfK7sz/kbJmgKTv+4SyuxG+9VIat+b1RKG+N/xJaoSJStTSHu9RNDQp9
Qcji4U6Ozj5QnaXEHi/k5JQqM6v/EvwrlTFjBx+D8RK0o9iAuqMUsMe5qYRWY3O1
e7L0JmLimjKEtpkm9WfsYk0V/AnUOP7Tn8z+Z8viwhBSXoKiejtSfIflxxmkA7pe
uMAg5R2KluvbEegQQJkmYmWIFq2EIDm8fdxkc9jInz2xhF04ZHOFM1EkHxEIKzAr
32iPMPuB8NNc/lxymmz4HRdJYVBD92IeCuqAhfDcHOIfxtPOFJeijuojJx2fezjJ
HhjsdKnquXQwKLIayJbABUL6eVeYcswhNTMVBZarjLRnGU/Y5lyXkABcjaE1r8AV
L4uFk4DPX5HjyVBKwFiyO955n4ZL8KdN3WQTlYKH+oD6aaAptGaaAkKAusnZQEC4
QyEmjDvH9RHfvtefnuLNIw0X/v3UDfCjDTALIdUslmPdkuzfPjadcEm4vBpk1Rxw
pPfyyG88hacc/vh88AZs0uxmkEsNct9xUcYn12kX11k4lRx6WIv8R7vjx3V1ouxJ
VXo72jApYMz3xnA4LueKi4v0GWvBDCMJHJ7RbaYqXPUAFRHCA4iJpXLIRwY2GU3+
PIFLeQQIlCVbNbFfqdTXEn0epXAqMX4XRUyKex8KlWW9nI0qy02UOmvjMsDqsI1z
62UJoaK6BJP52C3q8qkj1fzuqBSzkdOrtSRbAEVpEpV1S7LdOaUPe/W72uTTSRa/
PydJdKz7dXgxYSIHkhLEVybEQwjel3vLc0+oTFnNS4INDGdkt/n0JK08QQiRDLmR
EDfkbRYGqgVRP4CpbKqykxPc2OcZ6rREUbfA/rPLTkOIBmTuWjlAdIw4oh3Qe+ew
6lRbLzGh3bvXUS2yxvkxrKnLyc2YxFVKHsPFNXyExH5ezSJyHcE6DmnpwHBzZoDp
1yAvEDtzNJ7MEn8xS7bLpRERJz2enVLrqytKFCfetVWuQ8Qhhn0+5fc52bBgdqEa
E6fi6aAsBTMTZuTqqAarz+nurjHiNt1uz4ztE0PBJbhb9YabzUMORkN4rh56G/Bc
dkfx4/wUphdQEdksuVN/MKMC3/JIsikAXYfqH0UxHUs4dlL+KvLtUT0iupD4f65o
7sDRlmteHfHkIOlFpd+Hj1BE6d0ErydWl2FutnwTiO/GwQpwtOLa0dEdetCRytXU
7ZJ1vK6gNPHbH/XCogrgNvEeqYz0eZdSoLAJmG8/vgbOMeznQoPecW82TYt8FmuY
0fw0iuAYjxItRF43ZjqVYUsSrmqFC8sX55H4tZhwQe20N1xqkwIH2iTzP0gGegG8
Z56PKv2WR1tAoaXpCIzoHWFCjtzAiGZGw3tQA2HIrELrErWY1dNaOaYG8jpYYuJS
w8NHybqajz/SOLyrTvl4XUYcbPX0tC08s2Kt/RQDz14I4lBnEHmGapbfhoIKWgct
pvQDilC/5cBt++QpYdfOsf+5xQw3W5jiLVBuNMrQouN18vRfX5elpOo/NdM7U/8/
5f47pr5zfZmkKM6nEIs0HplikElEvjCLpgJli3incMjRbRQoPuCiKYoG+GBhRn7+
U1n0RNPk1FdbfsxWD37glv0Y1qUlp+5JWc3bmBq75eSvjzlLjmU4YH7IsH2coNEy
1Bkjc5hxoSbSnJPgnx0FviR/ZgqXT74EbAAXw6Ry+ZONaTV5JtYG7WaUqyy6iM38
6Y5RNAvEzOUrBbaT4pAw4JACbJ1/4BC0WIG+vcf71kiONaOfCit5zAEJst5yMJ68
g5D9Tv4Rzed6w4bQ+UxdEZCF2NmEz1YcgiKH5+TlSsnKIwVixaiB0bvyZGuwlwWL
9/0e33m5TmT2p2VgRtwR6SwwyBaIr8YGcI7iT/KibdkGXFYZXACz2ZCfmj+BjVKT
fFCchS33OGZRHxOFSbGQBiYj8UBqlqxWwRRKhBJE4uB8CD7rirlGl4/weob9JBBL
ZUsMc4CeF0u2Wjdvf76Kdh3HTPeHveNieFPoU0/RO5NTLw1bO4L75bvzKJCYK00S
WhqyjVdoN/+wgtV+2LJAevCMeB0vH+XplxAqwSCQZD7cs2Ihf8KV0gJX5mSZSoSw
PIlO5tm+mb0lJfI21A5l4zPrEqzn4s3vyE16UkJgwCLNracTIfNs4r9k8nclNv7+
gp2sua+KT7jz5Z5jRWp2NR//DcU36EHwacrUxtTvdN+/WkR54m/3xulk6/P6eU+p
O35Rw/n92aZqDs+Rq1um8w0d7C8opAI9Y9t+w2hoWZxh7ZG+Jp+6iZnP2nURrPQu
QTHKtg6YqDsw6c6Lh3PEPhB9GeoaHZjcQP2k+D2YqG9wD9U5Wy9cvADC+me9Vqbn
H6XRAdBj9QZGsPHHEHL2sVYLwTCLa4IucUwwHKXwCdUan6WteYe3CQdMyV48MRMU
8CLLOdy51t/7I6FLKK2wu5lbse66plIFw9HnuDPXgU8gLy5LF7NLEtgu8Mf4ynTH
IqMEzKEZzwoyZ3/mZvYW/1X14s7fsfI0bEVa9HefYKDaWK6tnpjf8v8+p7mWHz1+
RCx/h4ADA1w87MGX67MsWEYMGtEBxrC38qXKOdOYjoSM6tHLKJZ36+ZG+oXRFuSD
8OEXW7vlu8A5MzDjjyvnPlf27TC9JSyR7oDhlok/4igqE+P3O4cj6Y/nwO5iyheI
/seDptcpNXPLQZ9FxzXLWB0QRHfbbKJxwTr8uzitp7LYwX9My/iwzW8aTSiM9ekY
OyidFAWiZFvh9kqCwi0KUu+G5T9p07RkvuEzWNnc2oftq8Oq2UtdGHfsRv7auIQ3
cHOlBlzpViafhhjBGAG9m+iqXSzCfmCjsRo64OtQ4T2VRw37L0z2qliuAgjPz00G
JHreh2CN1V6W6DdokmFo25il7oR26A5k2/q6BO8VVcASnMMfiYCXHhhCnxj7LCEg
1ytfM/3RX6MoMmyJ+iNDt6yafmdIBdmx9/pstmYRs6RdrjkdEg/ICRY1p1HJeuRW
zY+JEG+0uE6GcV+WekX3vVOflRJTvssoa0XFegMYuXgdS6SDgr2PFiR2zbZbYDRo
u5Zv+Mv4giRG9b+JEWvtJtQe478vfpye60zRVeh4wHHa2kNX+HP9Gx4PyEFocsMK
hjhV55w1YSdll1mrhvPTCjnlQ9JqVIHZWtNRNMGQ7frZznjHNh3u9ECoGeCovX6z
OFHeW3s29Ej7KQ0maAAjXtv6WS4wvchsi0gnsJkEMihXTs7ABkYSLlLpF2kVnBbO
q+xXq7I1TtDJA87L33QuULlDnXqE5H+7Q8Nr8ePiIsIVubtGEE2wxd+Zpa9Om1O6
HKGjfs9djLFIiI9Pad7YOg+/KvB0ZqNXaBKTT6ZQMCd2APjT+l97ehNV4tS65Pzs
gqlvqV2Q+pd59vxPjw9vUxeSYioRrJ+4ZNzqbPa37VxFOttLVyOVFpQEP245EIi/
UYMyR4vMY9UmPHC42EyRhOFMfcBMxlYOuNbesmudgxBekSGc4KUid3PkwnjdB4H0
aRBuyTBW7laeH3X6XXU4QJQidmvF/Nm4vPTIAJpZmJuLAehSfwLJ1OsurKwkRNMD
07m1Z7DYJl/IrWc/NthyNz6286bHdzSx8QnuBQ786a1vsnEZq9WeyomyXUMcbDvp
2xH58P9wsG8PihX54jK5kxNX+CI5CfYzLoRUjPVsT5FP11VRVra0AYocfJbzZQ31
A3uNUTO7Mr2cjZ6dWa2rgMhVbMsq8RDFLb74/0DR3dAz7sgsWCVuFVkhFT/sDSZi
kVAmi71vtxJUgNJnGRvTN++eAKNDS9D2ga26jfyzyr6AGx8LkNCikNizokEGw2Pw
2z4+b2Uy/9pF9YXxiXo17qxRuWNGSbrnqIRCAYL/NwyXfEbWke4HjjBCmLAWFZVj
CgmMqPDdLKPsPv6cCZ9XG3b2Pvyt8tLH0b1eBhkbgyCpru8pUmoP6l1sGLohU0ho
hnW6Wj5+PFwqEd/GwqqSZIecZpQte0/4MU3IVuC0ZJGEsR1f8sC2IMTxzERpfN2T
JT5KpNZ2/IUl6WP2mHrqivsxZMKQR2pz+uqtGPCg8lPBssU6JX/adHkPg9nc4Q0I
QSlzQK80Ed2qcnSRRJ+qKwafNeVdlRdqZxsBAI1SxJfy+Vuybk11NY+cVuCfgdR6
OalRRmBZyR07p9cd0YgO5p4v2wZ1Lqtr+VnQ2eMfj+v0Mo1A3ARdFcn7AAypnoOy
KckjTN5rawL35pn6m056ZbkHMoNl0tKUhcDTXHApUQrf9XB/AHp4ZmRSggQaER9m
UcNqRkBpWYAXOCR5xFxXp76SF06aunUZ8CZ3Gd+HXFs03ViZt6rvY0U1oZhnMLrb
Ofu4zdb+SDg14XvkpoPBI1g9NT74xAnDJJuYXv4Rnkyjmg862WHVuGbjNSVx8JEt
OM9V7xYcFyfU1h9Zsk4ZV8kjX2zyLcZ0Q4GQWfwrcrNJm1upSHveJyMpag9mgi+i
7SZW4mlBcSRt2tfyORiKxmG93+n6PYUJI/1GnJtj46DeX6eZHc1FC2gJCzebYXV2
n1Pbbr3c3JaMEFndTHTq/zEpkeEfmj1FW2e5XeRKVCWg1igblNfZA/7iG5fkdn1B
oMYOsqYn2hkL8Gb9I7tIylmez5qx7vL07wqMW1/zfzEmD2tz79ezNu7pKuLxMIw5
xHAxi4Z1L6uX4RTTTXkIKu/7/MiOAuzPpw/GiG4FvQQE9pthMBJtBFjiGM5oPwqK
TcpjRb6degpheMhpFM6AzAkRBr1qEJuCWnJgYkd6kSWrYz2ngA4wTPdM2JUx+jnJ
HRzc7UaJXLJpJNx4BeQ6PwFw0bx642KwWg1JC+rjrUzic8eSQJUR2soV75mFf0SS
i5ocuWKsC3OQEsOF89uGW6Hv+gt89b+ZQVZAtVFcXVRRHOdB8LfXzKE+ad1UMw86
sfbl2QS9a0uzoRYAH3wFxI5l+Oj2x0pefRmFCJ/Xpt+ycB9Pr369IqN9rA4oCETX
THuLBiCCNHUl7Kira+m/PcIvKOnsSuYQh+UjekJ9tDOtsFcEOHurJJZ1A9LqJdgn
36SjpJOmaA/EHSzZqFnyoqhc6SweOJ0Dlwu/jSlW5xe1AiY16vOykKTbBh3PYJxt
fG0FlXSBhpFjTnQgeKGVAvJD4kVYf1OPc6TFJWf1BxfjMyTclUKyJjNZxrczcsDm
GoRdEv9mbYblt856XtfAFC2YCKlImVgoaJPReW6g29VWC7e0YjI6xNMn0gMW4HpR
CqAwDBKaHQna+y3JDnv0khs/22Qr6psR1y2jpfUHTS3o/8jZ9mQjUKl0z59uOjmF
o3RrclxTbFCan/1nV3K1OV77eSatvCbSrFCOEYHmRnoPp20kzreu8aWW9dhiIW3I
XxauUvjIqrvambqF+AtYufh+igriVJ7Vltbfvr4jLnyrpgzSfOjlqhwxE+8u9DIA
u8L/HVk0hvFH5RA0Ys3G//CeJjhkk34EpOFRwPevADkrZJFmtQ89+5W+P2HYqXyu
9jxSpzF9l92j3jpUquhPVyHo9talzHyRS0og8cWhR84lQvaaz1k6AhSUGWDc9nM5
VHtqyT2LfS43B3CDJLNdHU7mmmn1oy9Eoo3LD/mvdlu+w8ALy7Qfo6fdThD1g/5u
XBMLcfTXeRXke7jvMMuvJcZ6PJyp8CSgt/ut8ojTx8xKopLA6ZUi4UyGj8Af4yP+
TvR+IEl/R4X3ggdTxYB7wtuRTkm/dCanCm3ofQHQPoaTlKmkO2R0QsX5KzvcqZF3
NDiyA85lRjty/nQEQMWLmPmMXJYj9K/ZI+h0eCKcqpL7vX69cWHjpfQsSokn1Zoc
omUS7NLUGzpa8kVD71uGQQwi+vo8lPjoNCHftX++RXgYmbUBw1s1OurfmaznQ7QE
BubtVCGXPDd+tBNKPpYSy0HxURmnOd+Fa5pqOBsU0S4CQv7IZjQRdxuk99EJAvy4
BcIHR7w94jxFOvUJiPECa1cIo+LYMQWaHNseMzx59XS+OxpAV1alG8HjMK8lv9QT
0tmmN1f0VskBiPX8OUQgJ1sF9TyEuVd96B8o69K0uV8Ddxo2G03fNtCrWbUe2+wm
Rqm+UawIZ870Wuj6byt2RnFeNVmm0yC6RWAfZ51PJMQrTVUjTYL5/y6/2Lyjuyew
mv9zKyUtilJHFYjnQc4+/6RedeKnUgsLdMpPcR1VlJ/Fp5AUIiRjoyzu2mrvmZes
5NNzXMUtVIaTW6H7WIgezKqIfwZiHiazTcId09K7LlLBxBBTcDXF/COXzsJXnG3e
ULxeUjinSeN81YPjULhEqvCoX/dL94kjRBusSHuomHVFIVcNRgtXIfiGtRH6sllG
jVmnQs7leY+S5iXJB1Ggw1+kI3V4WHZsSiSL7NK72jqKMSI+kSj0Uo4weHzfRGp4
ypg0OV4inIm+k21XCi07QwVfbBuA3GYP9rh0cAOiPXz3IzVzgMZf84lmtJCmikyU
+VMaBAxUNwOT5AH/7rPavBgT3UQbWEIdV+RV3zo6XRAP/fGK/RKgPEJNiN1g1wLQ
42L0DKfhqGbAyb2FAs0Lt6IpI3e/5xpyrwSDykmm/Gg5zP++ETdGP2M8rRZZwZyl
K/E0hmeE/w6NKO9fAoI6DU2UJx6misnG96U8OE84gUbazNb/eEo/qU8Lkxm936Ix
SqAZfaQ/L7Ls+zQMFxtCy2jR7FODTx/DUBRKWi7oaYLZ0TajB/1BBAE760jakhPU
micBsvJYikqi1Lr36hFVtTXjCrsdmdyfcy+VKT+xoEIUxgkS+w2SUgx317GV29Lk
ArcO/4o1NaitIMQ1Iwk1qSZxAAg/PymoaPnJU9mMKYsU79MFZE3YUSWRv401oES6
ddytFNkhaCzxq0WKtszPFGVLqBtC/Su5siYzvJwKNweaYEPJDwK+GkcDd3XUwPqv
iZZgSSSIto/CKCWYWN+kUWW4bjwKVcDRmn0gDYYP0H3p6S+x8ARpPnF6dZznhNPH
0lEVvzUHMG7jQUyt+MpkuQClkvZ70regy2QAiWiSAIOcVajbirifgaxk01JBEQnd
wFoG6gek5pAcDzkG1iC7u/a41vx8YAhq0nSB3SK36JX3DpgTnfHrFGxtwyK2bVuL
dGHxiA5iRldUHp94GUzVBnlv6Sz9ALfv49k3+Pvhe/wA0hfZKOT/uchtGBEsK1wA
5FYTTJdwwfLE+13kln2kUBn5Z+BDHx4bw1oeyXIBE2HF62qyd1qjf6XTJYEFCJKk
D0oUzclegLmdQGlZ8CZThfg10LMAhNyDcKlHCNmdWoF2AlwR7rfko+ItEf8P7+Nl
WGKcoJVGSptuc7NaMX4dz95xl/gZe6SNssTo7zRYme9o8oT5LiQG3wnY/HdCl3OJ
FIyoaOdzs6fUFbonYSx8TmNNlVrIQXSdzQraANraF7jh1q2MwfqWEwxDiGqWTVfx
r4yMdSAaeS6efYGyhp9TU31H2BWw5FRb3tSwn2vqwNQ1n0GdkObnUB3Dhwd0ySXX
byL/4MlXFzUFcYgtLAxpIj3/2vYtwZp3I0bSexI1oau4T/YmvhdJuJj/w9CcGW64
+lU7DK72iR19LQYp2KqOYNM9cKygIuRAlNwOFRFD55GqplToPysfmZvVGoptwyHv
JLH3hXoz+1lxHIuCDTvt9p62F0qvv3jtpB3iuELA6OCiNX1CJksTPK68kJK1OwqH
viXo18jjWxhizTSLksghyYhCsqeexFtWgv+FP2NJziSBHFhgx8IR8y10Xl1YJGX4
c+cmwYUIbp134xGj0rOfA6FKzFefFV06wletKN9/xy/H6IyuFFO0oqbR7E7dp1Ke
3gHz1Ps9A7AEOYXurtQBMh3NLhdR/5jP9hdPEl3Rt3OVU5q4EEXEcA021Tg+5Vnd
qWWkinOisfTHhOftrlGyDgprp2imGpVly1tmuri+8vGw/PbOAhJkP1uxUvGWMP47
dgZXZo3PKkTNdqCny98Zs7MAyDD/ItZBaasMcwBjXjbVmHOitPIZHXTL54sfwzqA
icCfnWuq89aAVGNGB/XUsyBbieo7fHziBvbdBG3LO5YkIdJVcmqzjHMczYQAQVqU
+jv27itNk8q7sGCTlzBm3j56UjB/bZZ7aK++y2jYPVXN4qkibM9hgqcxXwje8X8U
eHzgp89DhS4Y3SOARH8SR0w8dhyOMwU4RJNPhBguq3ho96f96gxX7Oa4gszVGKpZ
XO+SI8f+kqoxsqeVfTuxQq4d2kjW5ghJFaLwB1X7Rs6NY5akcDME+Hi8RWzmxaL5
KUB4a9nTj/ZwVFMu4is60DWulLF8+QtTECmmcPV5eeysRWyq4AGn9CKpVt3donWW
e3EU7GelOop4eiMHvdXf+mr1gCNfKr+l/ohBdv4L4XghuGjI1YM7RFXFPoXITYDD
aXWMgwGvM0grYDCY0mfXR9axBaqYtnRbT5a2brRrmhZAYTqapj9vP3WYPC9oF0Tc
1CVrsDNjlSye3F2tzjRBIPoDpZ50YwzlLs6jFJ/aa/FenXINkitz/wZguJooy5TU
WS+Vy/CNXUovcvgcYwxqQZ9n1H1P2AetXm5s9JSlr9ne0YENy2HTbvPZ9gvPUchM
55AhhB6m423ewC9Hz3DS+taZpBa8s05+lKqDiDAz8AfpVVBd/uxRXAsmfRle0BU4
fgkyjaCEAoAvlckwkGHbyi9Jy7ktUjZyMwEXgN0ytIjyg7q4R5fh7g0xESSqHT/U
NZI5FKKxnb6hMBfj/0BTlII0Khgl5ZlSDgbdz6P3j5iaowqrr6tqyP+2ZICKMdBl
ybt7KkMLRezwln5+MeK16btymyAmfFXRUPRbbk/trRRAdEf5rSsiutVGcOsFsFc+
o5/0sBMObqeawp5AhtkI/eQedo9VDLhwwYaYvc8TxIcthMmAWBu9X8W+ntjopI3i
RCttBACYfOSqyb0B0ZwpJjayyK1i8MUjkUZ0xU5VYw0OdU0rDiyat8hTNeZAtdki
0gFE5LDNp6aIG1POpuTzMPofsZ9InxQjNsVQf7ORw/neL16eNZISVP97Ys/QVcyw
PEtJ+78Qc3TirswoNw64MKFB26QNeQ8KGBizjWZoIEHtjLIoaBoeRJXGQsjSvLZX
+0hG7EvDgUsu7fcOxgqhjxTLZsLBF7ZKRoIXUdbiZ5EflWMOc2D9gXtWrnLE9uDK
JMWL+1WmsoirGp2f0tmeaqALY/lUOSSrClF0/rBoPem8SUg9s1NE1Xn+95ZnhqaW
to5nRbulXzK7G8n3VN06r/SXylS+FExfU9F2dranu3ZtnIaravvR6DQb4YmkJyEA
P2TdaZ9DwI3d0ZGOyOgh7zg6Z1PV2WszmuuO7v8mNhNJC8hD1kArgChFQFU4HEgF
OtSIre5fU56I87uFDDNyES62uy493qRRnjTy5jI13Om7BCNlsHc1GmpL2HGFAclE
5ER/zCiB1mtXyeIWdbiONWQnMRLKKJbfdumtwsBkRpBhWsovU9fRqY6DGqUUqIpl
zQVya7jfACTNzJo0atBrUY9+btR8YTfSyoCO6J2pipmO/2Tv8ACrY5LPw9e7Ipk7
ePS5NRvnSG71o3EEFIwVQ6pAuQlmsTlkA4Hxy9w408hvOh+dItr1dQExrP+rRG52
+bIdQiqMz2zdAlcScqAmL1VkXjbDSfDMwp3wZ3J2co/hqQ96Kry8Uaa/NBqyAcN3
91Mn1dNnhaErku/9z06D4DiYHb49zG6Hu7UksnaP2MQ4IGwQM4jLqi/Pfxg8jVMC
Pc7vgIFW208ZvZrOhudWjT/h6IWMLInALpdjqAGyMW6Dcle+Xq9Fm1LEeZGvSjR0
a5SVTifcJFeXZWYGwPu/27qhJDTjO5J1eH2AwatQ+o4mFOgdMQo5egIMSFj+Bms/
z879sf9a1TA8bMDfTcn7Mp8ThvY/uv6U5e9MdYbsE7fzBwrtGDXYuwB1hxPF20Fr
vs+ljL49F4gxxneI8krOaUvNMM5SH+bwMpDV+/RhlhCmQ8x5Ij9xmvmj7Zp4Fj2Z
uDIrT0MGZ95u4/ZCsRFGoOvZjecL5BIvqCLP/kH5oICSfmmqEiE7kPDcm35CS7i0
xcXGn/WavVexC/Mv6kIPdCTX7iUX2pqonLNAjP5FifuwTCKJXX2JofkEJotPKgNb
v1oSia6VOLTPITp+AVPXfZyD0P2zrEr8dL2pb0gbzylGmBKM7Z38HdamttkNzUBt
Tl/s40604BlnRsmFusQBzwZ1wCIanbXALpQuk9g5xrQZ73tUkIUAFC2IpnrrsemR
6I9S4VEVbXPX7/KKy1AZFKtj1GrskVPxlNNQZtZaKnGqtYU5Usy67UEFXKRvcG8m
n+wJ3heKpPkauwSQV6P1Vbl/aevz21iSaWC00jhm1Sj4P1g6UmdE5IOb7z7cFbGr
UxxqKUKmwc0Ou5exzfVgsksfJaQHFbZP9fg4MKDK+X6ELifZ9Uz6kA0efIs+Yr+L
2OLAc8bPLfhN/Rmtx+i3+I/DNxlDtfuMtddGK8PEheoF42bAsEd6n6gpKH/BCIzc
X/QWQ8oqn1sgN+hmuR4Ofj8pfH6bxkheA9+9nHXLpS8bu6tzMJ1GKMpc17d5lxJb
/qVeB+2nv1COvuSRQoyldDljcsWJVMVVtoorbw+U191gF2e1Odv8qPtTx9xcHxPT
jGt/hzz/MZNAjtpX6itTTmNkETBRivWciU/esQEPzNlPwWXXJRXXS6Yd8jRnB6tk
AFCnxXS993j7gUJ5Byd0Gp9nxkLhYpRuIivwQDC++vUDm87V4QSsoK4JGltuVEG4
8tC2AobCgfRmu2d9FJIiQbRvcibPhl0rdQ985dkOfQKZR1Y07MTb7RHyS4ahWeKU
eSuj3o2GX0h6Z0CTNSnLJnODYMM/xH+d7KvV5VcnvCaGNvvYfUYstC9HckuZ7MhN
bYVIKiyv/x29hzeOD5HpqOyQ1I8mAB991u28B1uh3MEZX+g4ig15xsCfEp9GCF6X
T52kNCwH8rj2Z779BpGKJn4600LGcZwWuit5N6qh/fHpR1cAcvslqHKhPkjS94mc
+vapcKi6nxhOstmw9R1HlGCNNzAGNycYuO/RvRSwVbXgN8vWKbwBHFrGD3+NnqC+
N0bMEsnkz0dBYMTlcB3kqAFWrWmTkCHfmlPIjT9a0QmYcBgOT3mme5PUytXdNe8X
qTrsIkNNIMMKPvDubA+6pyuE4LSsZtQyFsy6C87yvEWO4qQQlv+TtWGwhcwSMtn8
yq543bRybreqoKxJNqpIp2J6CHWv37zjMcWBTpkfIGMJ1Zovpn3/+cHsPDIu+2sf
BSU8eGQbS8BSUr5d9XuuY8k54C50cWySBqfMOHCFiwmx62iXINcPZpnhv/YpuSL/
nnrrZGkCJRmtPh5H3TABI6GJBuZbWLQIPsSnQ9+Aj8YSAOUAft9e910yMQCqPPra
9Ej4N5GNdDrgHkZyGurZ2x/RUzpt+pYlVN2YuamRcE7I4xuU4dSh/RCy4MffL7IG
MqV8W0mEV4Hd6TzIlk2hfY8LCFJ9q0rjoVInEw/OSYL0WMBTPEXLTYea6IKttYAL
Z0wp0X7N9meIlaOLa6UC1c5+T+4YAcbffC/YTM3deY8fThegas06PvD2ibihtsnv
jnQxHwUoGlqtCk1TRvytwvo6xDwSPPlVjSHaQF+t+r28BA7UgvhB/g7NwzwHQM2h
DJ5Il6TEt14aTOs69AFB0HgfnNoPhCN3lRVt12leUg8xl9/0ZfIii7jIESlf5wIh
UuYfSj5sySSDKeSscmQmBxi/AaeFm3VVG7OyaLFnRQbebfe3t1tvFF6YrjgP5Mcc
Tbx4SNv/6DxZEifa0Gi80L5hyWKzmj08uLa7Jwvv3zuEnd4E3aWwCQv7hjUwFJKh
Go2BPPfVGC1NW/ilLnS+QADWQUZxkF2yopiO6qq/o8cCU0DipCfyUQEo08QZlv8r
/GTyjgYjeT9hvjLx/5aN/9uk9PllElK13eg912AfJNaXZEYKA0NylnQV3jpgFvsB
jbUG8uiqI96W967NurJ5RZVSHsXKV9f2LwlGCYX2XqeZt7ofFrcJMNZwHNtya6yw
Asw5JCBEOCJzDbYcSXXDKcP26warw9H3/YjFmDeQBFjtt9T6DDjxAJbQs9Z24i3Y
enqQCrxbxzf0RIzme8xJMZmfebT4aobNru62LrqYh1kxRkmZcR6bM4I3NiEOsmzU
kAUoElZMBeFMUNSaGxw8tI4mYA7ADhLoQdToSl0qYJ928EpD+eDWy+IPe9rIulYh
ygwW3eF8EUQAm+pyFnDDzfAokis0V6IsyY1QViQrWfvz6iyygirkfY7kvfI35CwA
IIUqFDq0K2qMS5/k2KyTdHzjdQp386mXbwgMkFHH588lGmn304+pvBg0IE69GvY1
ElTNjV/e9xNLabptQZ9usoFNWl7lbChjD9rMYl5PvlwS+d/C2upz23G1epvcH8pi
99/r9pEmmuSUHwaY4R/HNK9FWEm9qINXQk53jWio0PA4JCxXRccNjERCq8PGEL6A
4t759D5rFIG1WtCkwrBf8mYS+TXdGBymYaOPD3Rcot0q0KjzESq7CUpW+43epf2t
ej0du02bA7jM8OQoD7YmrSYPWl1Yk7yWHvfN+BBEEAzp01ytq/cXKnX2hXmr4cBt
6i7AvtQbFG60E324TrJeOF1lYpM4qVZNFU1cpa4QehziRwWcwvWwPJPToEuVfy1K
6wCaSNNP5X9NzIAkEW+1xxIOdYCPt0oUU07l8g03Xy0hUVhDHDHyCtTw0Fz7rBWD
1K/+k4aUlDU6cQym78v7zps5ZQjx98tpPZlYaXxAVf5fQy3wFPgZMzZi+27ImLaY
x5dnHZMrwp4evZzRoEFrhSUxlda4p88yBBdBZ4PcQgIelsO9P/UBp6SNAFEXqCWx
oZ4z5sdwxFwwi9CRwvgbSCbySU+mqJUDMZf1+TtGGlNXJUYDXO6gt9znge6nmkhG
L9mHJwDMPZguaHaNQEMN5SfFUDW7XMvu9I+UYCFiYb6n3yRLRfYoiCjx+k6dS6ZH
ii6XYtQ7kj0Ry0fzG9izEdgOKIjYVMxoZXw/U7QQe9bbdR3BnRrKwRaoclKz0ji9
w326PZdx4eaQtxRPyUQ2DkrQzz6+/e1ecLGA8lH0fKHBuhq9bZvGS0z3D5t6h/R5
r1STSQPkxi7PWEGkFGIDx5bQfQLna8dB+2mfnZBojgxj5xG2qidN183goPHkqGN6
bcbONaBm8suRovxUDa76MyqtLYVkGuwCcWXr4vvyVWyzqAaDMcVYUcp2bDILuHff
jFErPpgGOjDeoK8p+M6Xvw9zdRgLOpydHEGamSu+5J6MS1kV14Xjl+EMCWSaYnoe
nL4HVT/Kk1Ng0annjwlEI5UKqMaMFlqy9VSPZxPPWBpsvB3P8sgKS3enJ3MwhHQD
gG7BNps9CWsYWFEaOYws1am/r6SKX8Bqgdw2rO7tiCmflApfsyYJ18Gv2bM7GmvX
cUwMdtDjmFePVcvO8pyCLqnS3ZwLnEdxTYtbfdfgcxPpC8mKpdvC/633w3pktcN+
o7S0zu2QoHhdacVrw5OLiFn2unT11kODQCodC/Fpttsdfvx/rlp04i4GLgfiJGAQ
X32vQO89p2j7kEQ3pilwh1BtsbtFAau9eGNiPLhKv9tbZN8/Ot0xpSvZL42gdywm
+oAyf9fiC1ZEHVMmH/0bKD4TsHeb4e5nY+V8fZV+3ZNAOnxsC3uNTXDPbVFS7ucZ
rz6Edf+UUzoqRU6rpazjEg0CwrB0dRpPet4Nq4h/mmGOlefNpEcDVggRaTs5lYru
mosc2vCy01+Cp8UMJ+NJKGunz1WgEMiTykaZGLKgy5R5OnQgKrwyD0nhhUWhydci
V314iZsK8pbcQM2Mg7cU1Jh5l1NcfDJykNvQBvdXj952ojftZj0hm0GHBUXIbTBC
JJYrVnzb72jlT0qZ0gp1TggTwq2dF6trVJcwzSniRQIO/2+ckrRwC0koUP+PYhiw
MbrNnUwufANcdZoP8K/aQQyozaAGoHB4bJHBI1WP/BVqZe696/dlhKJ//EVfiLdz
+6OwKZ888CEv/f6KFFDxqqdnOfKtwPE0xzrgc/u3HF9ZB7XFyWl0yXCTAXOuzOf+
CV2FNnonDczkkIgWedMVU4zG9oPEwTJYba6/oe5REmVmmmBRAbTQUzTauiKhm3Sq
EJxgA1Po6o4Ccl2l4xSRaBQo3KHmCB/sCEAzo2kewPdacqxWyE4ZoWcM4qTMuOha
nE/W8cCoYPHrQpP0IW8pwBOy19+KI9KJDa2P6zemxaAwBZICNeXR8+XHJ2IYIqaB
WXlG7uA9klDcQ3FcyDrVaFFBzQNN/1ZBWWWnXl+p0wxautaEs8gZSpL4+aDrOv8g
KiSuGxqwwN4Uj+lDKKnHQLBoAB7j2Oyb4Q7B36aqtbVkMg1vzioUKlvdenBCvuOM
DmKtJBhtEoR+YtyHRxC8W8l1utdfxcXj16FQGFPRJf/UnDWcRcj/52Y09Q1DivoV
TQQd69aQXurgoaLZDvtJdTDcKbzYitMfZfrZPg3ufPYzaG8JMy/zX1neQOPzinpC
lF1sOpWbnw8B3f3wSGuvOw72R7zdVy3qyWTIJeRJ3bY8XjPG8Yge0Y/O4G5QxyCJ
HS/YCP2rkcF8o5bcxfQj6zi3can/0vdgMtcYeZ5ms/Q2TRKfALjyyslrSVBUJzPq
Vase58+oZOpRhDVM6HgQ2vMjgPL9Zbqb3Ys2lJ3aGFOHTrLc725ljQTVY8XeLNLT
ZfhNj52w0/i0qMz4idlVFRtvdQdRaH1mEhD0j8JYjmhOTJ46GIfwBh+lqxBr1z9H
MY7CJkin7EcepiDwMX7NLV5qk4Mnq7RViyNXD59Awjm3lk2wnLPHxtocqz8587qU
ztMgF1ipt3kbrq/gkCZdMgbZZGGmLmfbGi1iXzQmi+i6Mo+f5NQiFfT+puRIojjN
RuUNCLteN62KOvcfL2Ex2esgnlpznh99ctyIScJmH6TB6Eznfw3r9H7/C4ohj2Qt
JTr9UGXkG9haKqF8qK4dMEO/e10+0d98L7cXFLWBGDIc2frB8xin7TluW6g4eTVw
m5eH3RLGLbq8katKjQ+0zZHS+UFIqhas/k0EKVUyt6FJLIZX1kLwJYnXgrhCSXt0
lgDh7Wv9qVd+Nuu23C0RhUYMxUV51AW3JvpPalZHjqGsP0zA+ByLiZ0kkeDbGcjt
1LT+qbeVcwP2DyjMKMIfyCvbNNUGh+eHV0KKk2lyOczlqerzg/jaQesG6k5g4ROP
1RyG2qs0UZCiR/wbrZd7DTAqa8/+nB1S5yqROWQlxmHiWtztKn8KWLDTaON0bgKG
/75Q+A0A17gWZrAUBduHFEiYgs9g2NxG6+pMIZoGYXutdJ4f6zkzqYnjY2HfIYns
M8oHSK+hezLdu5Q7ItqIqiIrAgQuk0Dv5Iyw9T2IrZLKP7bDY+R2fIGP+E7AHvp4
GkxYvWioKXPyPsJF8FLNJOnzz3x41Kq5WzPwV003vX8JVKAGjkweBngWF56mmvqj
+mbxZNeGulKdVY1UMaYaNIlcI68iA9ez4kwE3issIWvx/03VKBOEFfTprtTnG7MG
hV2qBizJwTvfTeG7p7/vilcSJcMtUenZ6PoxaAjLfS1RiQ+GEEwHka9qI8HxzHYR
Kk2p+hFq5snCS/l6vHwIzeuJgzupmXCRaWBZmiY8VFpgEVoCDSU+B6jcaMhTS9xH
c40z1Vn490NKH1hmJV04VcBId/K6B1EqEKjJlNo75tqwSFAa5TZrsOBgHPHzf0PE
q4U0I1J8XtKNWjXCsJfo5bz5ZiqpV7L+qEotZrxhV0LRvjOAe4R1JPeITVnmSkvl
7Utke7SlsctMKmCDQl1vGtwTJQAEUj83zwspLa1WmEh0wQOyz0DJchqb7+0rOnSa
3jG8l3RfGSmT/2/xPZjcuF/RNG7ftI/JI2+2eifVezf6eWXmRaWDPASFX6hZ2sot
bMP/bvSOER+X0b/VqYmlBiPzhz4ZRN7nOpLXe5b84x/JvXkd6T3DxQH8DTBXU5EK
iQ8gv76PUgjDI83GdTcIySpYJXRKuZ47Oxj/tGHwVfZuKVOq8nhrR6/PhzUspDEd
+U3J1P6etKLRV2HjinQC+srRXHJ69miKwsq/v2GzZABipIquorhd+qTTm50/U9/q
Z5BLEW7FMenFUkbfiptGCj4k63+7e1I+steRYa9VGe6y2m/Q+Dve9fjSV/7A9sUZ
W/PBoStm5Wqzk9xcysZ3bqK31ZmRYzPLQ6X+bVsFt4VUwDDa4+fRkUJbzLW/8WuX
1TxsbRkRQrnHRoLZqke4ovv1SNM8ZA6mSXvwhD1Ndp0+RyfLrZNid2oMeG/OxYz8
MmX4PxX/Uw3nlHMKnOnAd4ubNzOdupOvbjayHVYbB4BkTefFgMhMuSOvI59Glsg1
SxL0+gCT9P5g6+VQYLl+8xnIAJHsVig6Oj8pdp9dHgK9DiSb5D3Mor8mti8XIcLD
Ki/+vCJRVwyHr71z8IDYzJOKBUfmLcZMoC1HehekSzrg+Ma5bAratW/luM6i/+jp
PpZ72gp2D1Lkmk8aUnjQiqVRF9jaZQANoemAcJS6UYnC8qsg52WfS3qrIxS626Pz
HOab0cKt1prXeDM9BCMwc/YptEAVEEbJnDHt4TVHWk6/7IKuzf4N8Jx6i6eOXVm/
VqNBJHhMAHFmlM9SwhjevRnIcPIZPgcdj1d+ZmHJuD16QBj0vpV8yAqncU/SC+ge
9RXscYm0Ch8gJKPJ37dnpYfc76SZBL2Fr4aReehrz9pfyv8GzMMsDuq1sbrDzU8P
gnIYfC0OUglosnAOtnUPIdNQxrhEYQpPyC+LLHxHYbgSWQJ3eN1zQkan6w4KJfdH
uB2jYw+z95OGC/l4t91rgh3vTV3upcNNx9h1wfakt/n4qTis51EVezGzjGy4PAfd
4hFBQmMKrzt+/LXqbxbXaPKlmzn/YJJtTyXGxVXjao65oetgoTP2b14PmeDvTsfo
vBODUjG+ng9sJIJf8oKh+baSD8cqRIbi7iSCaaZjt8LqyXlJ9CYgYN5uzUqdmyPf
dxK67ngrtH6kTqs64yBvptPlV7t1BdZ1DwRp6EsZjDsXvLVvAhjho3c/byHuGlx5
4cFCZkRvfsrNRwSQRkCCCoLI60+ah8PjQYAin2wnOmdj+7y7IR8bSccOiFCuEOFs
gHed7OGpDBP/rtbDKhBK0X5olx/jzcAs7EQxHw31VQz2oDUBk6tq71safpltAftP
o2A1dTgxWXYDDYKGGdOjeDCFYDvKK5fyePVskaxWRMH4zYo/8or7kk+NgMTen7u6
m6yGAEd0IARdTiiPKJcCbzWk7NvJ1uTVh8xopxd3IkWZBIeDmfbbcSE34bPo8THu
2zB4rWS5QW8MF8XHtx3krVtk7NqjhsPpu7KZghRjcTJ40hxtBNDVjfrVlqDmK1rC
JIG7LeFj1kSi/ZWx5uet4eUrC3KlGqBNwsnpbZ4S6JJNhBQWRYdVSXwPNKzaubhj
koxNujPfaMZWkKUOAvdWrRWoluQ/Fshb3cxUKxVfLlufV8gAe9zOQ7vkZ/ybRThv
Tq/S0PiwHW3kd7G/up+5XTaA7zOFDu7ZdbDQRaQauuXvg+EZEn4i+I+7GT1aw54H
C+6NjB0huEeCQ3vgXWsm6gHUkDBaC2xOJVtAsHu0A165KPeJ+VzZiVJ5AhNsubZH
/Ve1SWm0QIoXGcvqQEoTWnP8Yzt03MlZOQug+keJSmJ4lczq9lsTdn0mIdP+csXe
UbqF6R5UpnDDWiTOiCfJkfkKuMrnbCVy9Rdp6C2hqUN7JSzs1n2Mvvx4zEZqkymF
QtBOcvYRYHe8oy0IM4QjbR4lMjkt4v7d49mgjvbzQyVFbm+9byxl+3m7Wp5Ffegb
rHBLdxiQq8yS9P2MZq1+QkaBHGrkh8gNIoEDbksKQQJlXEYJC1SbiNZfj1TOwH/K
wiMZE6D4hWRLxA9+C1XFAgBvRBVPauq8tVbJivcSzb3IA4E9JnWnK6I6R9jW3b5q
ytogy9xExK4p/JymkRVguwootHFGs3/TFiiNJSJ2lZo9WLiHi+sFKVna+9RVbcWp
7vBRjPBjFX8PNXpnoERapBIrDN6D9CSMW4FIF+zUkAOcTDCN+uKOA8r1DNfTGIWY
LmnuB2+IGvce0ll32pg6CmfdnvOxQJMClcaM2K6VXrOpzEWzw3AT+KAj7NoVPnj8
PLxuU4BRS5iuXEQoy2QpMXgTxrSi1u7ZO+ij4RvqLokHQO1rJ1S4wHdkhtYBPHnG
1Q3Ad8B+KY8X8402vvAdn41o8Z1tJ2raRK2enunuUORcVkgPZ8dtO8nkpTWs1cHV
GdSN+hpuvtYPUhFOPQoNBnNZnytGv5xnFVgYcDxCfq5eXjM/oNPJBCwdwtqGBlt+
ZGImZchBi+9gp2qQIFIaxeVAcMJjXbOX5jdfZyDRgXgOBQaRFNagM3KL1xHZiTly
Cch52MD2lZEai9/6wyD2DBwxbKhCJql8yMdE4wiaqX1upgjgProVu7Iz5VBbt+to
1SEtvb2CqwFwtdEo3B3riikYvjmnEJxTWvg0XJ8pNbLviD2xzPJiJ6Fl+femDG/e
i2KMJ3kvYUzMFu6xK1DaselaOrhtg2PvrK62yP0/YI+3HJXli7+yDYGNsVURBCP3
QvO9oVpTc4dyt+YCzfJd7OWv4i+imWVNVk7KJg905QlTJcjfqBs6HY/XIdmkV1Js
QnqFsaiTAvy/TijsjRaRaa21+t5w46DAarFWNZI2WKF8XAx3uBwRCgOdR9MS9Kph
YCTLh3uQ+Ff5zLw6RTy8PMxJCZvhB2K6ggUTkQO4WN3iKLblwOP+pl9n8yAUTz/f
ZHJrCvOUQ2dU32V3Licu8UKkihearNNAYkmsIwt9/69a7OvnWraBZIA1Fx/XlUDR
+eA12ha8QDLWb8d1Ty0J/uCIsUDQ3j6N+UUOZbRKfaVsm71V3jQLq/zl8gaRciDb
PUk9QsIZCCejt99FIlfJDGJ2HBErFl+kdjbdiMbxBlrOz9ilv8EGi3QG0i3sdI87
TXwp1RZDN5LUuoXEP/IaQp2zzQIMbPUN9lu9hwcAD4i6mK+TX6f2CTvPpzBINZZO
jN0rkeZyj4DFLYC/0i5fyeIynUXbyAgAHQ8aGC05cOj2IS9LW3VNeODL4xj6wdN3
/pQxDQxUacughovy2waCd1o+8iIyoBLFV/PIlXVPeXDmWQCwgYHKdOWhj844VH5/
XeeJA77wOekJ/kIYCVlltxbjdZK6/EgQqjaJ8tqyoI/dczPtCAP5+67lD6JbUpsa
/ziLotu14NCaMiNQomDzPO8mkSHAWtCCg+osDjpV3j69joUpDduTKkjGpYxFG+V8
g0tss4amn4xoytNgBnQFtyhRQKYtrOq1SJmGcarFnvAQvBiL3UOf9DEwiDIO0gFw
37qpPiqReBx+XYhpfFYO8KFlPLb7ltPFtUr/TEUJ8Ia1n3zjXgUtDCfYQ8IbUYSf
2C9++8ZBuBVQJcl87UhRvfcrpL7MdiYVvYjTDsKraLuDtVOuZ3SG7R0nD7siUAuq
SeAKEo3IvAoJLBy2PNTdGVI0d2JU6LoddzSDscPvt+BzkV/lKj0oitVO/R8L3zlD
7DokZO+cKy+vqSR7txOh0J9rgkjGheO6Eh8AHibB0nYTtR2Kd3R4CmjvqXgVDk4m
7tZaFJX5EN8MKSlPJplrKTA2hMKbMCQ26YB4AE3CexKU0prEYfMuFSOTYjl6mGyy
aXh7u+SWCNZB56NTKUqclQSn6F9hUZYmul/xemgSM6+K1m3R0mjbpVBUiX8Um+hi
yuoi5FNiEro902zzD8Vv+Mk3IXsQLzQ1dBR3UocfvKRr3qb25houcRBXwiTFk3Vl
KhPYPZ3Znpy5y1bVWGxhH3hK/fSdyAfHeWWqFrTi6qdn9VlHMNUEylaSFl/ODGh0
yg8a0bJmJt5nDNrDjMUm/u7JKoRvq9A3nyak3Bet07FNjAuOhwnWz/0dQNpObFV/
ub6zMxeTPTLCD7ObOeVpFHKCQYc7EJ4xdabMoBiWJ5G2cxli/EhHJeEUz0XglIEx
QQRkhb2a07yYh0xXJZIEoqcEogy/TW15GdE2GMarMPYpmcZ0xRnZtexyUlzr92lP
KG1nXPYV6lTEH7YQk4fyX+M8hysGtYF/iGZZlVQ6Z86cqTVig2Y3t0Sp4xTr+dZQ
ONVSxze9YLxOG9rasqDF6yn0PTyWqWrbre0sp3ci/U0ejL7DVpWfvSivX8ei2kDW
p4k22pwUn/TWkB55tIBKZRIZI2d8qSxTUDcLYmdFIC8FFvHvukBKwe/JA1cuJqfO
gVfO7RYyQb8+7ac9dduPK/jJ2tP2kt6/Bo2bMsJNUVZkwmgTFghT8APXNf0yRUdr
6gSdiupoqGsoyBZA5lEHQtFQ09RQeMhDVmJCNtAGgLsBgK07hsluaCDFR8RgVK4u
jmqVQjUn1AOXhPnE7Txs6BVb5tH6V9lyoiIZPl+bs6JwWD4oX+Z5d/h36D0Otn3A
32TCHH2bJt/K5vpJjc7GqJqWzVJQUh4CdOUA0bN54ZP3e5vtTFgWhX1AbDperBZl
VIQr35zDpTsQCFpu17hYJPy8BMC9vlSWoweWInqFnfcTMnPYrL/ktLM++TGQZApV
C02x/g/NnxpA+U7VyEZosahrbWaG8QfvyBnQSlCOvv9k6U483r7REw76KOpff5Fs
FMpMCEABGqjC2PAsrlYWDzaEaWLnyLVM+voJQe70PmI+ydpQSRZHM+yBG034RlTs
0gamUb95omV/Zuto24jejKNs+4YcBQ4JoK6c2wWGjpl6MhKYZDyn6Vvbl39Bg+bZ
9ya7oGzJS1ATrG7I1VwWgYjEIWfh0UEJkD0YNYNpn7J+Lsc8VHKSgB9+vCgN3Nt7
Z+pk2O7RWPnQf/RQZtS+IxR3DYrTzzZ8Qd6Bdw+nZ94HS8ofgIPJVFaX8UOfx14S
sx+F58KDVEBxBh4hdcM/G4JM453nuNLrCs/rmfEanbl/N1wBtOtEVu1Q6m0FqV7L
Z1dIuaZPAwKxVUFFy/8e8v+E+SjWbf43BzsEenYvhNZ1wJZRuYsakh/kEKd90Qig
OV+bDlfBWKXmCZdkg+0BS3kf8dw1e0fgaTmCygnykc8gqOlEr87s5lL5puavchNC
lychjQmFbEx4NfsIJT9uX7c8e3xdl4kDwLgNPVewCDM3DFAuHy2mReIh33DhE62M
UkyE6se48paJ4UlwknAPYhHJo4TC9efIVws1UfCvphA4X0JoHHdE9r2peTqJPOFE
kP9cdwIh68Q9CrLbi3W09a+OJQr3AIUPry/S6QaX4JQ7NzUDfEm/oCEC28rkVnaL
ezfUUAMZXF7ubZVnzMTgHJ7U21dFIfq8g8pB+9oVe2m8cqVF2s/jZbl2mR/IzWCK
7YCmTbHVU50THeHh+vFB3E9K7+TFLYAGDqdrSbaMGud9H3/SjQgjk8MkUJU9eYM6
SmxmFERiuln0WAVURcC12vbicH8uNHGccbBrnwdzdGVF1TY5FlFLgzLcbs/xCx4F
bvCUsypkn3e8gt66GwQon3IRrBTCCnOXPwYTtMibaTX8aL2iemc3QU3z1ymgILw5
XPaW+PAzlcCk/x/zFgLk7OYRCMCzsR4g+ODcd1whsRSk2kIwpCmUtmM/JNUqJOn6
K3kobL/L80+VqZE92/5UDYq399w2DO26PB4XuETXVyrpjplSvcGeXPsyc9J0+e0D
ALo4tNZ4PoeHIb8gPfzqkz0Zt9ucvgR6w68Onp4iTBhXbEnOPUJPTq+9Kloq4ccd
eNhC4R3XKjaf9dp4MkSKhqYgaMfDXPQTgyRwQzKT5YF+phouH6QTva7UxqOy5rtO
5dc3MALr6cISZZ9AFpAzplBM5cVRBM04O49TSM6VJehmUxokfgeUMM42Tyv5L7tW
LRx2tScvseXAG9Drg23uimLoeoRSdj0ttSLSJUZlVC57Ri0T9eb6nCisS4XA58gC
8gp94JjB9d9H0/xzHQash2pdcDlSqaDMPJjxJSgsbnFuq65xuj34OCOuMQJl3qrH
Q1xm5foqXJrdyGJ2vqEiTSj3d5R9wVfMI1m4aaoEL/ykEIyvTIRuksc1cuf/FCZV
HuK69YzbSDi+7iOtsVP4ooBzO74Pa/bmN7Ju0FuwBoZpz2oDbmh4Y0xvL1ZVBoTD
0lQDmjL/XauZ3k7vTvaUABRAHThVsvn6XT2TRtLnuI+cgifkUEHOAHYrTvmPiLBK
wB1xxWIwmDFkH+flWKiRK2nCwzkv9xo81KItwVtjMHHaKyo5sRiMn5LQXSXoql6L
DagxLNiLStCwfVmTMRhZelWAO+mGZ88oqZGPTa3owhG767uPkazHtwKU/50GaxS1
nMjRkoce0jHzJRqHHlT6bDAq19/veuKPYLbgr61vYQUCsbao93U0tI4OeF4VTOdB
p0Y8+dD1kZ6SFEl60A3tLcVtcIyA9uNd4o+zSFtbROhbRgR0drWx5vGkmRaWegSt
ybGyBw/bc0M/jCJLL8xpYSgdSChNLsYz04MDfVYLHrVUybCzxyFVnGhe1Qq9d65g
bf1hoQ2qqxmGrToaNcejiNk7zKAcfGwI6WdjV+UaqnQQKgxo41u0WNZR+0PC6pgN
FkJch1NAFYWeGphsXm0RzyZht2Ah/Y4U6S6oIEIEFJ9HGHH43T/DblorTfOopgw1
WVUm0J2bDtkjbQ29TLrFV1owbQWN05V8dI6/OrTbuxn7L2NjwB8+uyYMTuKzX4X5
MrPBwoSLeTM/vWyyQbUXxHU/1DwbpBRaF27pEBRu4/b2DYm2xdRseeeNen/X7HAI
L2C8PfnBj/cLjRwuqbBpNI+1cwK35EaZg9qh6nN+h5y6f+YDLZHDgdyhksLpqgag
r/WHjBVh+1n7yD+VDSne2duw5WmPzrrpxRR9hSVuyYYUS7dlGtqOeFEgUJEmfKay
jWFkO+4MIQ7tSmnMphYmD6W/uNxuYGUJjs+y75aODBl8dfNxhYLuNPGYpu7rVvOd
CUcr899FS0FNS4UeIZdFZbPno5LXBeZsOeNuB26zBcdhIm4gY9lOSUclNX6xBEO+
4mXtTWIlm+m7xH2oMVhXaUy8c60gNDbsmwGKn6uVJZ9i1xGZpyy8dbus+89uiohq
8/Qo8hYO0KLR8OhTHL+qEMbPwsumqvUw4vA7orU4Dx9uUnjJ1EoiBNFYhK2ir49i
bZJzY7LP1Za1ZoSBFvKiL/F0bz330x+K28NDxy0h4pdvdyigoVMJNs58V03qOYv8
XSb5cEKU9+ZschvvwnafXoTgeTqUiddZCBRK0reaC1aX39jv1LoMd8eeoK99vDps
YUewg+geElC0iaf8Ypo0OI4MX2s7GcEW/jChPBpFQKu5MBvI6ReEzotaOLKHV+G7
X9XOzDcllr778w3vEg1HjOgi1zfJQCBCBqhoyr62CC/jz5DCK+ufrqB3e85DEA6c
mjj4a9WcRvU+5jmJlEIfFuoyS+m7euyXnG2hHMtMSgHvmCxAY4hRhvaH/AhhUcMn
jkghtBr8AqnjUReERSfLJiNfmp4dboKyR0L+STTN4GbFqTMekIXnFQXuDxqpJOTh
QtfHqF2yE27y7KhFCMqDtWSW6eTHIjwZeLqtd7l5q5jQoeWXgDUOm1FyLkKPRgVB
uTtEi2WIOS/b4E1SXuF9hAvplaNeF5G7Aj+g1TOe7LJOaMSqLkbXdp4ySEwH454+
VnOhRRYVgkrD6aXL9Yjkd4GQm+KVAZUfYirmbIIMmugBKpf6wWbuyrDQwqZNqv7a
JxWhGRtDPYVwfCweKOpaJBrxEq72bJ7aSzyteSLtjAytXD3GzfPSdOy59RrrVoMT
+9n19mfC6WWtAQxHn1/HMYDWwmKldGqufhMzhIgL3LoRsGDuc7oox9BilzGgC0W3
UTtNg6hFl1oxhmyhrgLjCfliq5b8fs3h1ShWNaHjKYnOxPMoaDJ5tbtugPqQoaVJ
hwXwMIKMSbKwNrLqBW6X6vg0pzaijkiiFXJAM9eynz2Rju8CEhlAUvIl9nXdj7QP
kg5q+Ix7BSBadoFSONlIiFQc8EZP2AIYZUB9o26ltwK9l50xwN5zzzQlPnuiUnEv
oeDktgPsNsfzHEEu1CLHhMvxhPUt/iUps4R0LXt9ErRVfs7TdX76KV41Ck3S71B1
IdVGkSaKX5ksSR+Nlhvq1fnXmk/4xw/GFlK0gkYe/wJIoFgJcd7UWVHN/Qayso+2
cuzESzfvZnD5OALlX+855mLUdwem+qncztIjj/veyfFS+f+ZpVrqyGRFh91ed57d
qNPnhd3PsuOE84tLOa4fnyVkxiUxUTl0hqWHaWvFAwSYtiqIPIwT/gpXuZrjBV/H
Kb3X47mvEplBj7KkEMVEi3LWI9WhVXir7J8n9KeuYZbGPqd6lasvCWKVYfPqu3Ac
MThbTSfaHpM12b8nvrwMbMUyDERU8Z/UVnSG7zZu0eow1WjSHHbVs0J8uDgy6bfh
Kl4UcaoFgGqdv5NUiuRJgvUdShioKQuAAcb2s3MvLh7ANo1962my6Clm1dzwOL2n
n/Xq4wXyL7R8qvPgS2wMciLt6sYnphAwQyAK8sO6MiVM3DzDZTmkb40wKSxjWAFc
vsRbnNORwAEz4QaMCu08mW5nbBAh6PJL0t2H+UI/jldvb9POtO8o0jm3Z8b2q+7p
2PLzU7Z+DSXcCbd1QOsaJfR4RrFxiaAneMVOz0JiL5LFSIwoDEZFnNiE4uB9N7Z/
gwKNtgTNGiPzUx8HVG6KTFkIdYRSoZfftgt1+wBDMez1cXvOC3NS4G2YipaJ/LEN
ZO/KBzB9tT+WXi6EW1eEc7z8v+JsVLlLj768U6rZmK6zA6ErbD5a0ZeyNLoNKVf/
6TDY6MGuwvbuqkh+Bf2GAajhpwQQrk+kjHA0qvouv6y/b8BCXUsg8X1NH1aYFv1V
+yOa12ZXlW8VuyngjAITfZPwaYHAPxZBmEa4OonajA2fDv3nGxlhdOjiJAP65lq8
3NAGkKa3/MWpVtjXh0FwCZgsNikM4l+mhnb75ukwShlmstB3U8VT+6NM9xzrL+Pw
8/Vybo68uq+lHHsKbbH3V1DyIiUKS8mdWO6yWAnIlZhIXbPcVHhfHVZF9V6wb3hq
iFrJb0bKRRQ1UsyUWD026YBVfLtvfEX2oFrWpL6x1ALk/1oGGvdcedYydAGemlj0
xiQgTcYBeKqbtnMZ1vSkvabYmBU8ZIOVraPygN+clnz/wDRtRM6e78DOlJ1ObNAx
7MXnlXVzFY0zYzAjTjERlUDuYSxmWk8LS1MhLr1pwSLD+nqsJtSKxrN85KL/R04U
/h1kOSOlGmfhhyglLnGnkhOmlUTz7dX+qknFtpI1bLMYl/DXTgnPgJdZH+OlsDl5
Dl9B8fyFvd42qyHpFWnlNNB6PaIqO2DtshZhsplJDR9gfM8Mds1SFlUGLZqvsZ3D
nsLaoSCkp4yIY8REj8swjWJstzqCGx6y3n866LmUwruFwK5sB6eCvRXBlZmCOXgi
yxlSEv8xgjgDarxkU/grFONWSQ5l0xfZNBXaVMHi2xNci8IZD8qOStdDOgYUXYxv
DkwFYTgeMObOUBl25U/vFg3u5oJ0INL9P+A4htPjMz3+2krHrDsH3QK8gglfnfHS
hKBrzHnoTge6lIFEYlI0MShfUHIo8aL89Vm0jCUcT7uVvLZFkOLEnzGF/eaSPrQk
7qbJosfJUVAXZFOLB+GopnnPMZPUcx65IxogAb6bD1Q824mo7p55TqtzO85wTU1D
OIdu/DEjB4MS/PIm0bhX3bJ9I993ROVFCSdLcUbpGrk38MdFAAAVsPwBduEhFI7V
0OeMNxI0PSIbpjSan8ksYQQF0w6RlbkAcjxm6HBrQs/sTHCqDtumdGkBWMtM2gpi
cR2eTGN744clKGsOma8TTGc8dM0zOGjl1b/IMmXtljLkCz4bCes2Mb+CW+tqYgfw
0XromATYOgGj/jLSR8DU28rRmFH2CKPyApQk/oSY2XA/xv6w5EFpkA7JWk091QXO
xizx4Q5xP5Md81XQT36XHX4QnqpNsKsynxA85cxoQQsKhv7t94DdkNHdNI4dWwS+
RffEiw0r1GXlORFDa3nkdJ5/dM+TnxBOsmAUuqVPbPiVFS6w5WUFs5HXS9xTHgUj
eskPRUmQYq3a20PlqhBhJWhwR3SoiPMKeKKbjuFK0qIg03GHjIwW+CrfllLs4/ai
MhCIBiuOdZLNHdBb8Ns6Mqdd8u8hET9Mz41v6a71bou4X/vSsQu+sFoNjzLWO6mJ
oigcr9zO+gQOPT7c7/Rz+NLrnSfviwVHQQaK0F2c9KBTaH4V0dgZv5Igh52KcyUX
WnSguRml0A7PU7hswZxLTxN5/r4Y+Wi/Fv2QBA16UotVD7FFOgLwhXhMNQUXkLdq
PkzUtBmKeIgFAjx4opn8S9//oAL74VUfXPgp/AX0+gVIUFgzGWnblvXRhKxI//FV
uUWjqbcInw3PP0e/gzrKpgzq7xYvEfF8gvaKBfBJjtxRdbFqRYiLuHosi8FIfNtC
q2VLONuklQpYBpt2FKh2Ire3oxSqycy1votmxaA4RL3K+ssq6zowL/UAblDkWhpt
C/W5sudWE4WylTktPpBP8enc6tIF+F9drAEluWKAK6oXG5x2nMLfCZVdtorpjkgl
yoynYVBu7SXJhkQev/FCppENOFRNltYC9056cYtLUKtb+Zcr7ZQL2RH5D3pS+AEe
zKQX3mD9k1MUgz244oD21yUIRo4wGPCEsFclMztk6rvaVaKw4eX4TeAm2T3cYfJT
0eaw7QURVPLGIltGryoxGuUH+9+lCSQFtYSYUw+id5lZYxmOQFtUnY9xLp+OZim1
JAYj7NpHI9qIVQWrjVdWxXL24JOcwl6DZw1qXA4z01HIlmfJ+Yr76Ss7shN/lygP
zup7J3L4/VgDfaq8u9lipxr1rgD5Rmoxdne8iW3C7Oiq4GGPAX6VZX2zF7+7QLA5
zk9iCkDviegJXqNuBLmNHXevrbXQftJN1zrgBRusjCajv97RGX6QyhtajkJMZ/tX
YnZe20/R7AZpVv5x823dhAbwhkZIFBn4tVYoC4ZKbar5VsNEv0GFyw45agBZdV5p
TB1FSkZZtk9Pfz8FihzPm+vAB4nRb6nVIxURV2ox2+cQbZp1NzhZZOL13rxgbKNX
MFGaELjg31imEHJK0McUKKsPZd0u2x6K+vj+wzqzIp9LA/MoYii7d2AoHP0UZqvF
yncj3Xa93gPRzLvmOd6Xl1FjMRx1GJxi9yAhVpJUe2nE4wDrqHdbWW1mFhPB2zos
ZwHTZ/Xr/oFFFjqX9BrHoUXpeF4eyr5qkG/6JL9hj3bckuQ4DvhNXPjqUyiOOYO2
lc/rXDoc1tjF+o7xImgLM3H9R0FShNk6SJTYbTmK6zB8DH0e14zcWgouiDy4qrI8
r8SEydaIZV0TsvY75zs//CgPeMxg9DLlhO+GL+mda6f854F4fRa7NQcw5W8SiKia
af1KF1TmJmCl+PGlzQYpsLJFDLc0riqkD9OMMmPS5sVZ0B268t1N1xYnoTtuob8R
I5fz5mL176hVY7Q+rkuZJgPmJYDkXfELGJNrKocYS9pVQs447cZw5M101iUEzRGA
D+zhjyrNhuLh9bM1Gp7uerYPwhqD4d6qK+v9Apl52CgIAO58fUR0LCtGudRELyPS
8XYEf82iUdkZ/VICW8HWBaJDY3YxlRBNWxCb1RDq+31WaBaWumkS/PYB1EGqtytf
PCo2MHNoaRt26qVzy+fQJ/0xjNLIqj/CQWbVqIDH6XA8plnF9NT85a4HCaWhdOzt
Yf/oHoA5TMviuRD43QiKEEBsxUumVwpSUQSSf/56KKXsOTCYErlSnmqW2QCP2g00
ThiIJ22I7x6koS8ldVSa9m4wDVGLOCM1xfUH5LGX59PD7BdbyW+Hs31Yga1hqN8H
i9asY8HV9dfDc3XemXI13N3rbo659p6iYuP5txTLIopkEgV5DKZvrj/DTZuwwGbG
Ofb03eiKP8LvG1gk7K+MyB2S0swO4vsCmeXri5Kwp2oyn8jZ5YOx1kYcYTNMBWcY
0MUiYSeMSm8BoiO+yZulClUAxPVSMmDBlgw/6yrIZOodZ1GFpuKGmqV0pDaK6+G6
g+hrqp8sJvmtOYOmYWy0+cgMZ8cr/TWXw1wJKWwF/XzVwKm9B4xIIijJqVywHbx3
nQFxJrrb6LemgxSw+2K3wt3hSzF0t2IN8Ky8FADaNZKIHkMKMP5n2VH8L26oMA8F
DcJZlQECJEKQOB8NJIN5TuZqzirybmhdcREQhr1OobDCg8pw+maZMyiGY2e+xDOQ
hR3dRMPE4Y5goCzjPxteaPSxHg0Oitd0q/4w3Z/oLGz9UlPpQJ+N7LPHtlH2k3/U
iRXAHFCjg5Zqy65S46O3WJpZc9oc6+7Rg/7NC63hW3+S858G69mex5/NwCjoPx4X
jXuj1pX/A6su8wBwTyP5Nv1BdY/8nK/38mqifWD+KKQm+Exaz1fw8QrduXeqxH1Z
Y9iJijBGghtdwx53a/fRgDf6OKhUGQIkzjoG/IH0Xympm7L/6akL6XxkVaPIn2lB
zJFqLVsU+NJvLkLPWNGhsmWv79xK8Xnk8UFrba1WFsVVQVcU6Mr4sx74xiTxrKRP
13XolQYL0npVCPLx3aA0MndXXhHBE30FLL7D2UVXByv4YWhWXRwcAUhuXjKog7T9
la7mHIhPRCiug/Vc1ujFLtoNpd76z6XqtKKrOslRNDf+0QTyx239pJ6OsImrze+9
K4SIvTfaYtmEPPw2Fq35tAfHwSe3wzXoFhORtWe3/wLQcvacpg+lzciYZriVMANr
g/o0QnzECI5WfvrgB3ZzEZnZ62LTHepqBrf6z7GPwb1pFy+EpVvkGSMo+H0gWMDp
Ho3nny1tTFL6+L2+ARBdVKVHQMpEuRsFjT7ya2FzJAMOLIIYrP9/B4mGFtdlFNOz
jDGj8SUaTbBsbVh+ZwA9bW7cMxbvDhn16YNFL8loYYwtu8ni5BOIO07jV1Y4GWcq
a7PecUq1V0vDoRaOTawu7SfST9ogQCzwO1mMcRdmcuwjBV4bRMp3A9+l2s5Lzz1D
hQd7beESUBXJ8peWPCpgqxPxZ1PUwy1lvGnniPwG6utyHU5F5JPcXtovy8c6nE2e
kB9yXbeWaZoMKZ3AyHOZf28QfwMfFauaJCfYCCxSdwWzpeVahI+8KzfqXCTyqEDC
SLEkLq0fzLlrQe/4AgMfdVJKnEoOM/c82KS4O/5i9c/K2OcphGEE5TUDQmKQlh0Y
hw5s1+2SdZVQzCmGIWdSzwKEbXCZE92K/oI83SDwI6EbgqcVFj6FtCCk8WLwyvMG
VhGJR9/4usvD3GPJzDixnxPig7pNjzeBDVieipBfW2D90FhNQ+PKT7dNQeFq6s/D
yP6gn2m0CykV9XhTZqOWGrlollI7sjDuM0ajw1z1eGe9KHOt7NBQxWV9Wi0GR/4o
C4Dyxh5emPS5ptOperEm6TTNkyB/HHh656KBJcdzn6whV9LIPVEkvzzYM3cPyMFx
tBmXmpZrcmhetsSpEgBFeQHUAOS75+F1GmFmvMp3Pnxbk3EBDVIagbEx72Y4ppI2
z3rK3IAWvRC9aPk1+2qhE/BGfvPIVeG73adPv3dGrIy8StSMyBJFF4bLsOd7nR+O
WA5skhNSVWjYuzSjsFBjTze91SCI8aTPGiD6F1DwDPCI2GFAWekxhDgeLUxo1tC7
cA92jakQm9oKFvsEa4vFE1T4qorUqEkl6qwtoObs3ObDltb6pgZ2v3umV4C5b26X
MjzKEt7HS2XJ/ROgIriMYIFz1mW9ucPj+QzwKqrMOdCDqVigPj3Qqq/YOGeb4C/w
SLmgWKtwKQ3KyNTVUYwxzSUlIEXaeeH2n0BzmCwuwsNjkf10JGds5Kv96BPIj15M
iCrIiP0CyVbEnhQem/sUpV9DjSmIyFkZqLHpHX6A6eWojW7zpujWr17iG05c3suS
jVC/ZGDOouF43rh2OF909bLh5G3Cr/AZ+IydYcd0acQuc/xGYLiO45NE5Ccfk8dq
bfW+I6Own2mxHB8uw1M/XUORDf9YORTjtQ5Rx80CEwmgCH4/8up5nsU+X0zifbS5
cCUAN0XyAb9yErGiUMRF1xC8wFUvDxbGl2JgO7G31Bw7GDoPDOaqhCE5sT/ULlVa
/e9scLNtoC4iAORBqIKpLcfqkD2gEijcgjErdMegL2v1bVnDzPIvv6AYQ5EEpJrm
KTLHcw7kkO3FUyPSxrQmsE7Mp0xOhOYukFTxdKStF76dpg7SlenbP3RPiU0CYh66
DcJLP0nMC1pTjKiP9GzJSgzKXRfrcbfBifC3jRk2d6WsjyEXScjdKwB8rnZE1Zu4
rrAbL7izHEFsvmwvi2RwgS2HqDF5HDGJPlTjitnl/kIATV0nGAOnH6jozefDmALN
vL737tmnQhd5mwkZTQLH8C6fpxmUci59Ur0lmZpPz1Aj5gUaeEiBgy62IG3/1t7x
jQP+aVq9ti3tVGVOU9kPWNFJUTVL27nWisuy0WW7k+cKhAd/AnyhPJhRou2/ii1u
PnDIKSR05LHugfg8hLfp1bqyq6plvliBoyyFt98A7R28AFehvtwf3ti7TfSwTRWe
N2ykhO7+ibda+ga4Ny2GyfGeS0sgv+2A1QVK81iMc2l4JGVPuMA/MaLXdtpIuX5z
nHieRWQ6lVMmD2VNG/Zb8Oel6UbqbWoI8ZiELdpocX0v+aCuQ+0H3IfLqFeiPLOy
pR1pDPnmlVSyOY8ZVVFOpk9moCcX3ObwXZ5djSpoEfA5uXGB3xrBOQYFxWTx/QDd
aIZsqiVqDDT7LxwLW7z87CdqUwhmBhIufF1jXRj7HWatWaNYr0g2m4PpHcaT6n6K
foTsEbpx+R326K9SNUfLoljmoLqScEOIhMySxf/5mp7B6FerL1E9JvSKp6JyU7Bm
H18N32qYMfJsBeQTNKJIxnyKBZUIh0AImWxF7jcwGSMjKJV0d2MlIiTAE6IqnPlE
vZYcIMN8dllfZBydwv6emzbocjHUGovU0aXrQH57UtjXEtCU9NalhuRElfSulVOK
e9VLjGev8gF5nxRw8pDp2Dqs1ziomc+RICCOJPA665v09gVKEkPf8nfwgNqZWxrU
T+VC6irDLNDUgBlp1P4zuv0DkWpezXHMhUAlDz5Ct1vpmgiiQWHctGIUVuIBfw+u
36AK3bR11IGHni0KSsTlNFYXgZWjLpqjqu9uYBa0m81R69Ew6KgecnxFqtC1R3kx
6P6lKbQ0O4SfpYQJR4TQ1a0NXmMPcc05vewtC4XNPbMemYyChf//8AT6TbZTE6ar
mcGOmJNp7spto7P7GoKBaZ4M6LllTyAZWL8bIVHfqCuS4V48TDpiuQStd7legM3n
ICmZ14DcUfgbkscH0BE8fBAwvu0sDZaaPggXLeTDa/0cN4ZOLGSJh3/tiF5jMeps
FO9jOgyffOj3/gKGNKPvxaiDM7esSsaRhsnaAPyT5zUJeFCIVa4ALiB6/Iwsxdan
nZxukV6r6CyUlFtXOtdzl58520J19yfSfiDvgKgIK24Cxwb6qA95Hl+NFivwOYSJ
ioPVnp3F15vKctoz4j7Z4QlLEg75r10yPpBujdYkMWYGooPZG2tNexPBhhRVxFNJ
H+TCV5tTvkCSzecFLQrA3quWTu6bCKS41FadybPZ4D2xa7+Wge2FFcNx2bcDU6Jf
sXzB6fc4wnNfyrD/H9A3oV0qPMOsyrTrQ6kp8R/5aEk2BJxB1PjnN5nWoYHJ3rMK
7hz8IPrJXsomp/sidtQoTjD29urC/78ANXJjkMROz/OZMIY2wrTfW55upKuftCpn
fLFRSl5AGlGqJnwuMrQQEJpEP2aq0Vna8TRYt3r1Pi/KyZNYWq8+jpT4rRS2E8xY
n5dCd8RsSCLnrhOyrqPOgiWpIr/w5vzxpf/vZfzw0BhIPUuS6o74CnYips4/A26n
Mnr1iIbHc2RWRs+KV4qzn5/zWDmb3onEkh1ruAXg/CzNLhz6tZM87c/BzoxiOCem
hkb44m1qdOl1I8+wyleHw0zlxN4NslMtawZ+COECkaa3D98XI0fpr5gwCMzpzLU5
k6N6RmxM139h2FewA5yRvAHmaRVOd1j9m5cti8IPT4ZOLi+aqEdfIM8xpige7x8W
jnI9Xwmmaf1kxJOVnxu7+7V43iMjqGIWr9o868EH+5W4f+Mil3Ztw/in/Odk8Sqb
RrLzoGmn31+3/E4lM21XXvcvIaXzpkJcQfXY38aJMhPSkB0IKqKm/pP3mn+HwUXn
n+Gua+FSRNplt397ExZI8vQIv0RdxB38fFvBA4brTN8UmX/90S0Iws6LTgkXOX7X
12Iarpzf31j2n2VVXSjxaxR4KmiS62HzhY8F97yYrNu/25SKIimq5Lh1bDlT5GhB
WgJWqcs6juppoATPLODqvjTORP6ivM1hlKhCUlwLYcFzIcE1nvOeAH9T/w2M3UOE
okeU4/4ZhUZ19/MfIwS9uuOkRgpI4ZEdiuFBkwjwYs2VsY85M1hJWG6DgyfdEd5x
gRNAwu7USVYKIsXz8UhWDfNbGWjYSe3Y7+SmC4zFp6y+w4/sx0BskuP22gjc4sYd
thQ/Uq/EPaq75f7Q6xF+XfpKxLp7jEJOGMPZ1enC2U3OW5hH+VDL1v+AYlgJXRum
JEgq7njTw1xAR5oTZ4WmTVNa9+nUfi3umCDEsvegR7uoEfr3oUkntpo+IiSilDJe
6GPsnd+YKd1JYv/srWz2cGgugJlervQ1jrNJ3LEuf5Yt3vymcWpNLr0WssaqIGes
0GiOMHPgYqwp3uS2GWjXpxQ5cg3t95j2IBJNiLLZIu+tozeBcnYRA0jDXMHz0my9
KO94llmYJJNrlpGVJTgZC5jl2o0nKTIYZoudVRyrBLSQM3rJPvW6xTuAdUvLVLmK
3gAUB0lW74Aaluktkdv0q/b+LzAhnlE21Xs1XJ8XoK6hv551J2gf9CdtTNSpvV/v
7/cueO2mt+InY1WoAKl2H5V1UK9KfjSKLBXCcW69DelrNQ3cu+j9UaP6QNeAZfRD
W3m6angyvAuqGRzdIJTPFGL6CdYAbwDM75m2ti4whukwWA8ii+dOUVwLrYftYSy3
Ox6MarzYFE1mFJRVKhnjhc0rFrriY9Oc4492HsIRxIdFtDGY45+3NltWvYzR6gMb
KY/rLC/94sH12zaI46eTE3JnfJjwunTe4a0vC+zQgN2EjoO98Akyxq9yB/WBw9/o
kgWwEOz4fG+lWVC8Qav4WhUMF55kowJmEiiBFXOjOC42EkYvGpRZEj32kz7fjayu
887+qPrUKE0URdFKXX586h9ExJjT8Zt67kbfQI4Xkg0OexCnEuj2JqehL1WqCq21
iSxKNtNKerqEFTB659F1g0NVXvxxOa7Ss0ZrTlwIl3zTdUwzp65YS2nbCPR9PfpC
1D6yj7XX/Tl/zC519mkbwelvmdXj3GiHYnwBAZyNSofB4XLnPRF6uDIBrM7Dr57B
BcKNsdGnxWssEWOfXF3kbIW+BqhvWiATKPK+O07m4tv1jwDdG9q0b2C65pa/XPOy
Y6ONv/Ng1PWDiguDKkqie8jjg+s4s9ui+/kM6TzjDMtx7sKfA1J0G67uP7JY8x38
tahrHsCqE92h5GD3xiuIJjarwHnZkOeIcr4+vo+rULJpBlaNmSCyk/FPFLUz8RHQ
wPZiUQhfJxMJ7BiQciibnPzIlU1z+mMhxia7LpoKf4XtGPzk3oaj3vuz/twjXq+a
AcQidawXsEIxtR1hmx0wTsFgpK/sEFSnYo97a8BEyJ2+9yrDCkncNs95xo4YuUHB
krDhKFVqX891SZk/HPw78RAOYs8v/DB7zfr3bR/cDtDJnptaE+b++C7QCtcytBqL
3eonf6JfFwxiChSf/ph9FeTFEr8lsjbhNFTjPL9qapEzFF9ME/am6OxrPIbJ8XUf
xvwzAvVmZInuzulOkJwK02WOrRGcD4hcH/tc1Eo9far3xbHwY2ygRBkjmvDNiWaD
t1ZT7To2IUqHN2FzwoN/0YeIEN2UJ2GAWywpf/GIWsAkDcdfNpbM3nGBcEgWItdT
NVieo3d4Ey68XdYrvFLCj930cLDc5y99AiHPQ6QiZSHoPZrgkuRNuZZ1Ze8UmSyv
uzL0+HsPHsKZYRD92M3BZw06Nx03u+QVwKUp9sb2rzu8pj3gUQmbXhWgrjX/LdRX
gAP7dJOpXtTGvB3/vPPPvY2j+2buURI1zncTa/y/x5l3nV2WK+dXNxL4U6CxKHt1
cXq2r6ppu9scD5w1zztP6XVtMcr9uFARnQy1Yg9MEEfQDQzpiPpmlGc27zHihlWp
O6Zctc61KBY1sFD8rENhpy9AmB4M4c9rSr5ZZbtGG/RtliydWkSILAFsOUc8MEDw
jBE2bnklVqfd/BTlHGZPpjc9fwS6m6bMb548MtIHhbxZO0pV2YfPSC9buT1a3Rsm
dMRBHRFnYcevt3g24qd7opyIqR9XlBTzXriACPtaEmWHedMAILdPyAaw9NyEwCAm
Crc09ZYXy34DUs+ZCRuuWOpIgZjumjtK7MPpeBa9yehkx6O7rUmYWCZSEnX+IOzO
8JtjlEDRNZk1LL/3WoiQTauRsoAlQRyYmB0r/dI6qaO5BxOAwUGlIrsRd/2Ch0EV
9byhy2D1Y87kDFvbLgw8JSBv2FIJIdLQL3jIkaUg9E4zkN+nfPweGpOr1s4ZOPw1
HPP70rq7AzUYSOga8bAvBS0MEzIeNN8D1zaQS9b4YtXkF6tzBj5fHiefZbbGke1f
5MoLXkS9XnfAnjwY4Z77/xwN2qWL8547CACPaYjDY4WT79v+hJ9m6nGCBoZTKXGh
yJrbt3OREvbRi51fOhskSJ2HpCT4b9Sjzyljar6twdu3e66ugFrE+nhyD32PVVfn
q37KDCSFupbHMzieJZ5nSCEbSSVY0zGn4G3qFfTTJUWhyrxl+LB3Na5/TSHlG7q0
YFIt/PTWvLvbEPlX4WWTa009Sf2D0u2e4jSJrXo+YvoMFDn8ge/btyh1spr2m4MK
cji8RcDbmfHYPiy42GVxOBStG1BldEJLxDemsNU11FTffG2aEby/oaj/HWU5yzxD
ke6vyZHXIuoYZyIjtAVPpPT5BKxfPBSCErpE8H+SCgERYw5I65AgKWuxIc6iNr2Z
RtKjxraSc6N92k90WSwT0DKNnd3uJN2dXqPHRSze+VWIidYfb4klREIL2dbK04b/
JKLML1/ApCTirqPPaMBSmX5AFmOAwD1TMEh2fUEJdVWcvOhCgFkwaepmpfa2vPiu
Cq3ZYDqewsdhcYQvRhlaK6X5yNKHrGz3PCn4w1UXOB3k6tHiijhgGU4i1aYCDGlo
m+H6aZwtXjcU2FN7j8jCCIaSqz03jZ068i+FsMfuaQqFQ0y2tYgr7DvcgV4NELGV
YM/JX0gE9Zp47nPKsnukmkA0iHvE62tAMNj4VswZSilAukeSuYddNZM0Y02+zeNE
JWvW2nzBMVCN4/tNUBVNaJ6rS3+mE3aXcb4m6B7y0UipcSI+fHJ7b23PXHh1C1Xx
qM3NLc0gmyFfEedkgvoJRBTQ59GUrKjHwNXux9TSckryykuV7AWj1TtCMTm/wgJi
kiRzV1lnqj6NGP3S1CLeXjT3iwG8q3jArIfZWuoijVqfuOG1K26HYlVWUyNpbbi4
18lH1QMqmLElI7vjoRXoIqF2nhIX47x+gK2xtHt+xpRgPT8QoYSRxVkeQuZoVO4a
OtuJX1hjeoq1fYo7h3yx8U2S6QNFFBHpirWFJ3Bb7Q/iXFhdu1g+yflfMR0GKXOU
fJOKMLQYdUcMyhAHwGoxfvw2KByX2z7MXa9BcCs32t8eMwS7NvMFRwUKY5AxnQDz
brDU8vvS8AnwZ5V7nQsxUV/6cqOtzpllGojNQZVEafdfSmNKuvnjDF+pf1pvegQA
FloP50PGsC+g4HSrvKj9c4OC30IlBZnZlX1O5GBHTHAM7Yt86str6IVWMJL7HDrf
VgaP2jD4I8JMeaHlJmBAJ9UMuHLtoZ080ZjGgQYLvSicVn/HhCgdU3l4j3PNUF9O
S/lX3JoXW5Q2W22VSrs1ll0anEk8GTXcnxP3nu3EsYiemsvh05/k5QuR+wGSYs13
4jFit2LS+S4jNNBeuU/U73pTrGC9iFbu9UJhvfqhuUlcjk/Xsugy6X5GtbE+HKK2
WHMFAnUu/n4eiDUqwgn7f+JD3Wb/9YsLs9rpWqV4I1XjZNT02zBvSYL4QkHrD5yo
M1yK+5Wi85JEBi3FP4YzAw3FJpaLJFmrD8FF2JjryXw6cYjOZhiySkhZuH9AqLza
omO1Z6KgTGG+V/15hWoBr5HlJ618hIg2hGcVOvWQLti791RbXmDiEhdHBFXniTqF
uz3RyCzvSfSNpI5U8/zoV8JboVcYBU9WQzAdbxkgqqwRgbVPmd3WF/t9PNxvEpn+
ctIPndTqxQvVQIiIwVVuHILh3qIEh2DmtCfZXlCIHpIrKogTyOogQRTJy3sasY0s
QH2FuaiAYntdLk4p1sCJHwll5tReKyPsE/G77g/l2D3Nj+Mk7Q4fxJB6NBykITfT
75+DgcG9d8l27Siy3RCusrcu3ZUdhidT85iknzHjpBJR/jKtoUwbWJHXaVlOWDoE
6yqPGDtMJWmUKjrjjAiJH2ARrGmSDG6aT2rCwN6VN2sA9P77FabuzTSH4wO2Ve9/
EqUByP03OXHoSmfAzieKby6St/sIH0Xpnxzjd5ylt/upYg6D5uHD+M9Q23d5ez9c
AZyeT40RYS5kVnB3jfGwoAbg8wDcDu7J1zBMT2xegKW5Z2wd24Jxoch8G6dRQ21w
g10lMoNaqicWT/3Rpm0LC6qANI4lZsXyWn8HoT2n5uI3cWXEM3GApp2iI0K9w8Fk
zylrKWo24pDTXLC1PLJ/QPSDUzCU2+lu9x/3vL+I//htj2r+MTutSaU1mWNUX9kv
1BpJfqpeUAsAC2V/AMcWLTUJ/Rcjop/DwVLI9H8byksvYCraSKrv8yrA5SobY7oY
VFSIcXZUapk/I4IftdFSFge519F831RFBHOKYg9L22vmiAZfurY+ecj0ds43+6u/
PDyO33HQHkkgyMuavMnu1V2ccQJv803HQLlZ9S3pI37XTdPb1gRwNfoqpos1cdW+
hHHMopiEbMRtYsAzzBVoErdkj++d6duRaq1la6XaB8a+UxwuewCGRSxAd9OPacXx
HjI7i6V5BSiJknxQ2rVijXkUTsWBvfvwIzmyPlnySnwoqWivS1nqcfgoS+OHAX+i
2c84AN3BmEtDPbOCZWhG0WTJrjcHBSjbVWc+sCIxSenJG0ELCcPQWU9iCAzLELqb
X+YZoUTtRe7G8F9POJa0ZVdy2GTqbU5mBBmhNjbXEdEdNB0PYdhO3Vf4EwubcrrZ
LjJFJ/8x9NtPoQkxvXuzD4XikSynqc4RV/Dp/3Wh/+dpaL3Fg6gdYJDeSzNQr6eS
NyKjxYB56S3NiC727Yx1U6IRZ78MffsadDZXJkC5xzbgeLWyuBUre0WZAc0l+U+x
11BU0c+jY7f+tsTUr0XVgA9QunGKiojY3WYMyN7IkQxB8KUO7QhEzPCTJzpU127U
5+Aq6VO2j65rCFm2uH3hk3nljej49N2bO30ti4aw4aht7HJpmtmr7Uu0u8/C5DZ+
4FAwJbbo/PiN1iLutVSoozx06JIVnxlfbolhb5Shl+HcHgSUuDeLiUcNojJPhmo8
xtL+tBWZzIc/wt2uWdDLpREreqiJso/2afS0RyvIqkPPY2eJI0fdGsu2DQbT5CSj
fD2qEgJQIO0CrW8dMoxB3AJXIDXsgi1UPbTn2DqTj1y2PHTr9//nGIFE7cdUiTIm
u+F8nuGuhjgrOJXaUeDC/wXxQKQVDsK6mPPjkx+FcgzbRJeVWeljJEL8gAogP7Fw
l7nuynCrKHW8ehFI3eOvvd3OBro3Jvgj4oPNEXfZ6OWCt+OKe6dpiAwsAjAb0ViY
k3j9JR+xbMDZNvK7mPE/+pQe7zA45n7gckE2rLaoSwRiE30ZsLpbyfejvBpKb2+P
igOxJ4rUGAawksRKe+UO1cMAWBVIGPRNGMmWKulQzMqHQnXk4RFeAePP1A6v9t6u
UF1Qphu33rRgoS4SqY8ifCjlc2BJUZyybw5dPOEf4lS323cPy/TGt0hsirP3CwOc
KW5kP1CdM6P+VvruNgEydSk5XIu7nE5KkE0QKJLNg+sTypM2T/oHKobLWuuIb/dw
jQkHwQM+DXAv5fn3Y/l64KIrUIhhSYfIEbO/RQdfNFVh/1vUl5PCbbPQQajiZGTv
OP0UIm1KAuvEah12GG9EpmV6h3G0xF+/koyLxHFK1UN+Ri8pxxjMwa8DaCqc3gfp
m4AQVBpEpqK6OHAlA4h52DlMzjTPcMcoPOSNwHdwoQ7hAmKjC2Y6vXyeBsuDcuif
efU2ItiOAiRdf77l2a+NGmSFzbaV2IvuC0WARZSL/ol2kZaTAZ20nLew2Ao6OKnc
U9ci3shpPUoHWW0Ow4J1gm3jbUL5vuYRnfdDOr3rSA3GlgSLrcfEcZvKqcYfeiw2
xlaZ/SyCBAVY9TyYxz8Ca0p5RgFVOzo3J7znvhGMlkvM4VF/7tafy8pN9B019yMM
ALavlYeLf3tIYeZT6JpkTzwOQ+Hrelo9ZqFL8ee9JKQldjbMTzZzU8LoITIbCHoA
WCxug5cwhvddhfueL9sg6ZKU38X6oOJIQX/YbX7Dn2KrWW93trqDx4pcQYUZzGhu
bCNjAQecOpBH+3R23uFhvFoP1QUVmtbtiVyZszM8TrurHyTlvZKWHldqiFaF0wTo
GHmCT11rMXJz0VGURnn82KxYpla5zI6Y5TQBYFA6QJBnYEQ1DrHcKfIGh2PtOLK5
UvNrmWmkQQQ3KAQJYn05Ggz9D1ngx6pWBhovHNNp644HQOh2ZvjalLZVLpG0eAng
s1USaTNDvN2AQcFhAYP/LQR2oceDRP0XB3c9WYHDPQMpff/gdcdxbH11IPngPOYT
zL/crjwhB6VBJD8BZpWmYc3713aD6+6wNB72iefRhFHqusw166hF6Ai12Y3MRtoY
iRCzXC8hjGr3jN6RuzIZoKpe4zDplOTKAyQ6L9xKVq9UFUekWXXj2mPh9KRPpSo9
kzE1E1DMDC+bDQIG/z3ow3z6C/RgW0F/+vY8wTH4pyDlO4EmfbUH03aUsLQVCDTG
sZGNpO2tpYb33w7aRoJFfgxuSX4xa/vjO8hIWrVlzsrzUU0n4iKCgnwLwpOafADL
6jUuXVu07aDNQHl49ezyX7veGhLXGslW8TCxiAVNqYjR9NOIzg2Cqc1mCMEWUZP0
bCKJvza9dE7lZZOjQV5j28qJbmzybAg63PN9kPZUg418sgCiVlTg6a7C/Czse4sb
tReCCVvdG+eD5BKZMzgPUmq+5koQzfBIvQ0msrLme4SZCPWncsmGwB9WMtHG8vS6
zbsmPCa9BFqHJTGA8Cpr7o1fIFO4SOzUjmLaVdcRNsD3xk1/fE5n4gB8VLZzjhvD
mZEBruSM0nffGKG4ZosdDvnosHtJSqfkFXewBmum3FRu+6Aj/VJfCg8ktwtMN7cA
WX9tVBth4SxUi6NuR1Tm0H0FC3DJWulIucJhA5SAlKZsJjlMwHZKaqxNHkreOLeC
9Cvx/AnvVP0psUHQdVLsovNGCOChzHEGtSkiXO7BsYX/XPuQiLiWavCQ7ckIpl1n
x6Z7GwXJ1Y2Dl/ib7Do2HaaJ/IMagonPGzHor1ytrD5N99PD6LFf6b9nA5RANikm
KVq/S6grnFS78pu5eloazKpJOCIPANfjukb3GtVsHVr6hHf3sZPoE4B/bw9nCYG6
p1MIh8pfzkLMlsVWvXwDikEKIWKrzaQOQw37VKLEeVVbYAhlm16pWvq1+HAXeDU7
Yd0oYSZxmwsnF8rLpzoCMXipzE/dyGEhPbDmUicUqjYFZooWQULTOtimcTgslRvL
E+WNN9fFQZx70phUnWfoQPBJMt3txD6+zXQ+EnObxPcvx/kCta/JtTmFPqeEQvRp
fkF2N5RTGXrGMKw+IUopR0/Qh0W/RBKReq451YdVodqzl/NM9i5GsbZ0sL7yq02e
ZG3iLyvj7o4iNFKvHAzsFiRzP9ExhEl1eTbEr4opIjrItAQUb5UdVdirdFNbJBV+
gVJMPXCVZNkbIvh53rIRImC0IzcJ2exsVkzUY7mXSew/xDjFqr6w6x3qBRLgQQOR
K4st6Jmtekqdl14tA37Zuk8qO1hPqVHpIIu9S138oYnkx1RmJHgMmoA5flxEmJMh
pOUByapBEHKUNhF1szLJ4+6PfCbGXKyYlyzRGS+qTxZXqv7/71nLO3Ij8941kX1B
kEJEvqw3VO0Kg+WZDxknbqQMDZY5dcip+A3XiiOQyTzacDgPhWSQjoELRTnxbKX+
t+XdTtrAP5G63TIOwDqdJ8yrtrz9tviK1sXb81Vr78sCwI9pGZ5KDkKWsbqf8SzA
fjgXz7MXgGZb0W5/NeIyxDzPKEqESvtcNWoVItWtRNQ2MJMAD+t7nN3WyTjGs8I5
yZ7azVZuB6UOMU1sIrooSLEjcGADjafNzVNogqQaEZNVJAr9qYEJTENs/yuuYx/N
24byPtj26Rl2p6Ki8K7jo3N6isOkfws0G8ercmkG3qZstfRm474wEXHT0IT+5lT0
An/wDKmM9wi7zElxYao8hEoc18JLXVDmziXb6jJ9PMdhxtAVPXzwMOsuDOiCsiY9
siTKiF89MBz/gcOXXk7BoAhARzjm+1SfimgolRwNJvVXaUk0EPcQ34q7kbzTS0Z6
s2kMgfCDPzs1JP1uifJwkJjrVejLntuou0UqBsqwTrRc/oOgqSI/c9b5SLlvrj42
3/QMw/t2X2FvPHiOPtcI49W1Ep+uU6CAUY04gw9C2DgKhGgLCX2KYJgP11iV+Bwb
pVF3Z/0xVA8axzf0ulKqBpXB7Av3xQdCc2VvaFDuYKxi2xvyGF2zRvzJUs7GhgBo
/K0FH11T0uDoPeVCd5gdHDBtLq0xfb8jpoBDjpjdFIfL6Uwbt1wdHyWqSknxVe9i
RdXrBGRPWKXBtuRXug+8hH3G6b+gq8Upc99sey2vVmFweiwWmclpXnV57lztpJbL
PdVlECQugD+jqHz4rxCtK4mu9P1Zg83vQLQ7wnLPvX8uA3VA20BWzqHLeR6tOLyd
BxzDeiI0IqdMZOObmDnKnd+4teCBli13Fo1OSwgx9jzy3g2DfKuKk5attES+vE/a
FSH7BSPw321c7hl1RVfYrGqA2kkMpaZkfa56LvDV6SRKkyI4HuQQP41QGiuRm0Tx
0d5TPhA0WL+TJAS6FPNCyWzXitWGhanZve3bEyriL6eXe4lyrJuyh6H7PATgqOyf
K72tKYvACmmZ8kxtM5W06myTMlFJ30qaA9nkAl6hSqPEM8Pjiz1A21XXvGb6Y6XW
2UPxygwhNLgClKjrYpZfMrgvdJwzxfL2jZsMgGxHOvpAOb7qxQAOhkiU2kgW1OIY
OQtRPV63i9tZBhB138KM74srDCMwAxv1XC0WPkBVwxiaLYPawND4/E4eJBI6RX4i
UX4JQxPOcYIl2S5gJK09Ald1k2mQ8/zvdnlVTYlr8P3kXeRNPyKB+QOMN51/1DZz
8NfHc4Dx2uZx5ECh3dFPdaPaX4AblLi8FnHe1fGNne+x59L1cWlQj5xQbz7Wpb3p
5B8aq7SfbFpeH+2jHpsb/cFkvypaRCvhhD/Sb2bZpPC+zWiPmHqptcrexJ6Gj/M+
gRt6e0ZhMyrP/3RVbr8GEX7ifP3A8ewf6JiF1uL8uiBLwIrKoMsV+VjxHXRE9tEN
JIiB5SRMiCq4Cd5NiW/fAgL571vtYo6KdDs6bNRCHhwXDg3jZB4fLq5d5oB52UST
joVHXeboB34ZxSL1u4rioSPzTYp7Q+c9+O44N7xG4aXrEWO7lYK5MVqaKJesUAsB
38EY2KO4TckhglUxxRBhZvqSSr3DWnkuN79iaNsU8yDOApn7B//C7zqL9N0OA70i
eI6M/wF4P0ME5KAF3SX3t52CQh1lX6SymmkluXa8MPSWwNCyEQPXtGMF/abtcjCP
1YoTEk1NJIT8JLoTw6XmYxvAXKl4FM0wqsEEoxgM/tpIi2Itln1l3jEZU1TTVilf
1pJLk2BCl4BO0LriUZsXzMAwgh4/Rgiu86qNtsDj52ojqqgjUFX9FtuJ60vK4h75
rBEknoQ6qxF8p+drbEb9lIYuOmdOsc6k+yxYlPt0qtFqnga7G5bW2jOFRELB2i9O
V0MCUpaVkv+fMyJEL61tkA/E+ZITDfJujWAnNwxUbY96zzx/aM+A443txq+eIfaU
jelaP2wcXoAnQbfh0TRPVVIhJ8JZktLdto3eMZhG7wnmofch1vCnObcalzuSnsgP
QxqCaz2ACsQ0iOzj3MYEw7FMObsfOBbd28Haxa0gLQw3hEufOOtQHQC2wurDxlJK
rUrChCVnEz4VnOaT7GgDzDKz7wmoxuSZ674nH6GYCe2VaUEevmO94wsaOz2vxRCC
lOtXKKWqHxB2N3Iy2m7BbJvF0J5RRC6n66AmQ2Pr0u5v+Fj0wOEkDSdVLZ1GTwmH
cLoypAgxiLTziWrNKJ/8Fi8OngjLbaWo9Rb1b3q2jnQx3k9T1ROINk6ogQtFRoz9
NyRp9iP9sGYNIlcfgKYrV2fd/ZjDF/m2M6D1R47ZelNJ2QXNWypQC0xUHEq4OKC6
1CIst0+SObh1CF0LBLcZR91nZ6aBoI1xES6Aw0CYSC4RPpOCkAcFWeJjyJzkWvYw
28d08vr605DL6rsWiXLLLUAypxJjDc2+yUGu53pFQ1WKfmMxcNwugrg9ESVwelG2
+bLDba0wPqSO0qaQIhcPU8jl3i/XprmG4h2MtZWQNGNqW1pjfXoPZrVowDha9DGu
w7vwk6cEXajdhAu6Amse1omYltWWOG8mo4kLTGJtdr8vvdR5WKAz67gwy5U/wOHl
v8TtWsBQUx1FC6N97g9q5hQW3qWLiKmMstzV43t5rF1arFxcb3nDiyxtH1A1QBf2
XlGE265v1YZcadtgjbWFxiZB4a92Y1qg1n7UNAcLwt47nTCCI6gaM7eLgSQcTAkW
W8tTAEzSQaWiwxn20vyKYuEn40/nzCZaoOKV/e7/gqz5akBqbOrxVZ6wckLKTUlK
aWbu8lJ/DF01DTc+R6IRTEUOtxF5CG9pnKLF/Ts2c2cj6e3IbBGCBE8eCWnOxstY
FNc4cjSZiL50axUUFsDu5Q/1ksuJfS9XiPcjfz4D/6ZzK3iAzHKiRdZpKlDbNspW
xHbRn0Biu1o9TsHurZqWSjn/fnEyiaDuYbR631qaT2uQisszhlNtf2OYoqbNnFgq
QHdIQWAUVCmMvFjLB2v78vFS29BbzJZFwzH7m8KpuIUDulg6pphV+lGj+pzqN66w
x9p+7ZifeAhM/LNRSMeXu+0IzxsF0LkQSIOLmtC52iFNyR6fD8idN2krUiYCLy4/
iSf1NTN2UVewbHWYihvyC5Y9JLZHJ+ch+NUyTYlrfzJ44CgZrT21ZQdL7kFghTc4
YqHjcXRsfilQ0lY+ISOGMxRpOihtpLpepFcKomjQ8e7ElmzJFspvytIL3RDfrM3G
8d6XgQSNNAVOozQ3xIfpuuICU70DhBq86zDFik4sx1AouPUYjBG849FjufRdu42B
lhdpEGRVTeeqbw7NtCZxzomqYEdv5Rzg4Rj6rsUKky9Gkc0W4jsp5DSsoZwY74Mf
EY2KG6mn5eqFlQ19oZrY9q9T/NQj+sEFy+FFBr9iBVg/v0XU4Vniv8M0Z5OyxbzV
HLlTqWKQ5HlhgEenVh8ZyCDFRuCtyrP1GhToUdqkLIRBotr0rYlbDaiZgehi2nJK
wc/NMDZtD8bY1gJdTlgVNKC7nYWQPVb9PBCs/5XlxVx+4YoFq9CxrTtgPGV7BaqM
CaU0F2wOukZb/ucCfo12D3FcxDpKRsZHK5q1GDlIa9BQbq0fTKrnAwcfCljkUEGd
88qVziF/pA8PoVfBUD0Oum/X4poF5DQqzOSxJbF+HAjoFImmerOJDaDbEF0DwJVu
QYZ9EClfdi9hrsfDHgYyXXLSv2bKcK3yoJk6wa6XJ/iJru9Lpg0QHRjbdGXf5sJ0
VB1bGGVvAf2+rvWwdDGcAEb+BHGe/1C/lbgr1pfCK/Qz5vVnCv6C4rK+zk78Pfkf
xh+a23YBYpoVvL7hjOPwNPVp8N1PrYAe7PxN3A54zyB6Vn/uy0yaWb820ryHIesj
OGrpolS/sslTJe+eR3lFOhgwD31K7onboa/pFfTVmtJQAAqk3k+/lta6IGqsA37S
aOpUlaGU/WqKApxuBVwjJoBg6WtDZBHy286BqJwegNe+SjSUiRcnTCE/Fv4W4yml
aOLqrdIxCQnm+0edDiOZDJaoddZ8XMiY+hCWJBLdl+BQQvIqIyr+Gh5P5/DPLOjO
sa1K+fnmBnzwxxSPr0OHesx57wnFyekEmeTYn2nLWyGFTTaDxLO0K3ZGEJ9TkoUu
nHiFNIreJ24k8TzMT0M6agr1YV8CV2O7XqBVBA/ktAf+h9rq/OPU6IoPrT7uKC4z
xUwk8qeJyD6wSjIA/iWOM3NIabXXOMgUt6NyY/7gN6JquhCo0Ltd9tK9m7TSOYiX
KRct2FuCMog230ceqWByLI6wN5qEnJEoBqEAM2V+6y8tTxAGFwMk0O4KhXFkLGJq
S3myBznvfTlHodXQls8RbprcYZ2DRudMGe2PPbRL6R1t593bLQ3XtPRkParDjD7e
PUk++KUOZ/U50EOMbpJYVXOvern7svbGMb0aypfFh0ePpoqpykqWNNgzZDPUJD1c
Onxh17t2TEUnhKFkABT4pldyzfkkg7l11WavEHTow9ijV7xHIrwWlSi+d4SuRl0M
S8KnSdt2gPe0MAxu00Y0ORt8XeWq1I3kOW+gSpCQRR9mldEjEq/VNXCjSqVhbyeS
5s1Tf+D0GootmrZCjY0W2k5mCyo2VAjpblFnlv7Vd4KHfx2Onz6M6PN1C6c2m95w
IdRBZf37NJJM4swQWXCvXCTadkvf9NRk21sDmEUXQjZq6IhLQ8fTtMecPWbKlT8x
XVuzl7fPDkPIIrVrcWF+IFcbQiLoM/EzrksRREe1y1mnC3twa07bfwkEvz4jrv4Q
N2p8mF8JyWKRIlwuiSOIltmfBeH1RJ3ROeX4iGtR7vdxjIDWhIoJEHygXt60LLid
7INdnq/SOz0xxqtxdrCpOyIBuHTs54y194d5GZ0AK7ORIlFzkZ92iydaiDOQo9w/
z+jif7fZHrDL4+thWz696uJoUecFSBuHMR87VmBCbswc4N+lDRdpIwIWfCs47ENq
mLTspDXp596NV9GJiNrm8eN6IIRAk8oHBNmO4Z4ZDwAD/TtxRl5XEnKmRqgifSL2
4rq/t+y9A5NjD0z3rGI8as3mCLuheiYrhJKG3fvnqjjaeSM+D3UvZjkO4Pz0pTSE
a3wOD9J8urBmAazoRSKZOKBnZXlfKQegL9yh+wV88jMUJ/8hLBW0DNivqPABuPAe
ZaqDf4Qwjp+VzVOTxIH8djf2SJYq+DICoBZ1SU7fCWRpaZAcKjFM2kVu8I/FqieH
4Pqcnla1LGAuSYRmf35BYHWO1Z6Cv2N9Kg0I2TL9oPew1Fww6fClThUOV7fSHUM/
7xxaKSIoJnb0eC3Yh0eCBHjgyql8Rf4Ni61diLLuRdIFFAtFkTiakCU9o8MLOvXx
Y+7rzUDYcZf9/0TqTa2R3sxFg9OLDBZASCwMQIyARMj55doQoUiw+SenZS3pSKWH
2LRWYWr7zP3/H6ODouXh5WYkyNdzHQfF1q9iJv1Ot2COIgFjXiqjEbzNh6wl0SzL
w+wRL2140U2pWxVgTssP7aWgnbF8zXtVm1XZnWKdS0EkaVgayAz1YehbJZ+bYtkI
lmO5EhcT4nGclB8pPW5qhqukhwCRKHgLmrRvDo6VxGCUOaGcJgw/wD8jVLCEFHY1
62UizmZlf2jyafCCUDobUyhkaV65f2H1NzxJREjGcoT91Yw3Y0IQXNiIMJgdv89f
70J7tf1+A5hrHPLPJ+FwIsfmBYxLIy3h55xrSj4cxbNu0XmTh+UUIVKVUBoPLByl
q/3bNonyMzHYAFwsqKNjk9RfWLtYDVtJm0wnvf2DOl4NNxvMoysQYmExTlJWwOm1
V7u8qZEhXovCxRQEPJJ96Z39Tj7o1Qig4lkKtj19jdFMhwBaNq9MlwFSq8SD3khi
JJokNXhIqOw1s+WhsU34Kqk2Svai+Kj3dy4cY1TY0+VMWnbCrMlweJkjkGaiQpdK
7evLD3tozdYPhlnMxzN93ui5ZGkLXLSvIL+u2jscZtRUoocw38JEWt26zQu5jdqo
W+wjC/WSReyQ9sApF0mF9vH+fX6TClYUXXy+0ctxxBbrDqM3K8LXcLrXdCBDUdKh
XTaD6Vy7Mb3DNR6uPzhMW9sO+oKT2vUjoYJz8ZVRa0PzrlupUig6fGcltXx4ejI4
mRhvpTzr2ukEIih07z0QVmURyGH646Z25tpAkA6j5EYaCc3mzJgh8wlWS6fxzffO
wNPDb0YP9PtEYKgnNgR2z2+koolkYJNQRcyseOBWiDLMyfF8B2KCs980IPx4DjDB
h/rghXHn83fg80FPo23yjkWschjMHxhPfNv8dU4I0BWbbNZhvkFrH/pCSPOa8ulX
nj7yp4mqiYICz4/lJEF76RvyMEuGreY4QX4x6qeotnZr3INjH4pEAKfR7F2X8PZL
AJ+0nnbs0eMITRu1WfoOTTQAncZ7kFMTl1cd8rtsbFcEUZ/p+ZW2zYymBoVkh2DN
v6amOhYYLSwAjQe3vu4Bt5QITHZq+c22XJ1h7qWuAN6LiWF0DskD6KXFNm8zTW1M
79I7gPBBgyXnJgYf1SkE3gOlGk3+4HAfrGdKvBp+WmYFENXuVyGTiyA3KNuUgwHN
8A14MJJazUvFu5OG8eohJ7WrgT4bjubWIpoKn5WSleOci/p/c2lKXtqe8HKN6X8D
MpQ2d5Qq+8fEJqm5ORkmSPr17DgnhfXV1zUc10SMNZs1RkOFEpQ+pbDhxw1ZWFaJ
qf8+bEgruwVMvNfEO879h/X8eJ7DBM6/uiHMNZE5dhTux5eyndk8ntOMMDF+Aj5/
Kg3g13SFXT7fw7bc/2n/0aLh/wIKkXNcjXOS1p2tPbepHpKBylVo0Yx+J/sLTqcR
gbjBsBigC2d7cD+X4/tdWDeufaozNes2EYfBAk4+I4GWPdiBlVuh5r4C8JREPPE5
YBYfV4zbIkeEwH5Cd0LvImIBVQZ5oDsYHHkg0eZABp1sLfXzAAguCv0Drg9bXtRY
HNnpwlFaaXfPlkqiQnrHM+awC2c8IEIJEpeQF9TkKWvemlgfhRgAXBEkWOGUQdCc
jFKiE0MV5aMy/5d4TYVw6ZR7hv6x7iUGWBdB80CgnE1CZhMhlBFkzKDt0UwVVrCb
/MnVwx+I2PNA4VuvvjQi5Q85KJtFf5foRrJML64SfZhXdf5sIKfL150O2Y/kPYL8
+30sI4Opqy5iTwmk4T6QI1IPXR/kF/y4/m7+qDm6qQDys6Mo+v3B9Z0cdMqaCY+l
grt/fmyqSEkSW2zyQErRiwwxu6Sb/Uah3FJwqBON3WTbD7ZiF1Gs6Do0mLlyAhYK
hIQi8FHfT7KJaqXsdfLyGYidPLB8FZ+5/eX9kE/nZc7Shf7mLrUmfyJslBZKptK2
HMRL/vmi1UkTm+O0UpO2TVbqy7ZzgxiUktE0jeekFrZnTTg6b8NVq2YR/9kzxVXL
6HbAKXrbltiSuysdSK6G34Fwe+lKpBLKL4xxy8VjkE+zx0cf0DARyqjCJa46JkpN
MkdfM/MJhILk+nSdwse0sR50TZEMrQyF/4BskcNtVrxC+YpMIC853+9ipqWoiTAT
LKmLXo1x/kKcVLDtlkqc0QoRvZdmnqslbzYmHgC+ZsEAwpn5UM1jFqgN3Qx1/UTN
2BH3IMd75RRWpkdOczv/sV4IpYob4trdJyCdeNhrGD5d5xgp8E2MlUJDm/Zt+3Cb
HrPRjb1IWRpOpwLUL367fC0h0Qm6xUa0M+voYh1EItmjSdTVSRIooTzIVmAhquFf
nuznj3/t32ReZwtOfflthRi4LmNkyE3ICtJrz2XkyRkewdNZYgMWrP9EIS3O8dMa
hwsVJjlQIHcTw7JmAO0oeOpfTlbYuXl5OqjHSVaNxbImIKxsn5Qg12ZWwW679NTH
v5t8mFJwI3AvtCq4giprIPgQFRQfwZ//QXZVUzeUBHGUAN/4T8O4z+qRiTSYxLkU
VQV7g6FDpJ2qsdWQsmXeDKtV3dbLmr9VA5d8Vtl/mgqqEOXZaRuPBbpyobs8b+0t
Qmbqz+goH1GGR2xjf/70iLDluS2F4+DvDlGQhD5VBXiK0g5TyRuS06HrxU4BsFGP
9+RqTopHbOxMIaYudI7AI+wuHyOincWvLxSJ0axgQ846HFK9eehZJ+ZMvBPIG/P9
S77B9jCpw752ftRUTaItjjyrQfvZY4ipzgJhR/dvdNZhInvodpFd/n6cV4VK+qyT
WApFyBB/EPCVHavbNyyvllGOl7GrUlC0ii18a81QUm3zhjNKUw25re2120Cp7anL
0sMkkapQ9T5nSff3jFRmnDIVDa8PWjYuDh1H+faHJpTiEdyD7KtlzrhyV5y3GmpU
YCxBDkoxlSHsIlde12AXyCI2zX3WBXjhFlmCh+bBl2pl6afdANsm5n82ls5VOM1D
zf8w4AI7+rOizMIydxcajSBVbU9mYGrS6hb5XMLVw7C+zTs/E5QIxl2IWYGg2gme
D0SEV45MHb2WwoZJmDHLNu35UIwe28cLxt5CydDDnqSHeEHF6sMtCvbPUX9xnq1P
FImPE/NNSiUD2Wbr81mKsxiv8hOlPKPjYa8KLdghrFoSv3GqSLb+Zvp7pLvvjjbn
uO9OVa8u1wMJOBZIdayqfWWIuYvbnmRwgvqe3MLbjm/lFnq+nxKNnwmAlF/eCNza
/d2jCUDyVSRA6wqoA3bmMYLSqDgsYfayUsqB+nznT7S6CIrYZH+kVXSD1SZojsTq
j3swTiuQw87Yk1s+frTMm/GIWFhQQfHhXn8GoGhX5Pie5VWbmcf+ZIljGRe7b6S/
JPvbZ9mDhr118Fqb7SR05loMabqftPJkqxZP/6YrK6cswT7szxVC2nc3lw8slcq0
ctfOOhVS4iVN+Zs3jldw9LHpJ7lrtE6vOCgA3BbA7MdmYbx7Ax0OLhNrDIgVNHg2
KBGAAW9aCwIOWGcs3Jp0V+YcaRGii3YEU8em51uNFFHQ0byj4kDRo1iD/mJwXdLH
sw4D42HiOg9ZNfVGSR5N7vhYm11f9ApC5lDcp/ZKra5Z6+eNFThNcYEc0h/ZRV04
j3d5Ma4hDLenaczY2HJ1KIXITdJgOsh8VnDIfESZLDchwjHfq8MHwBqyli4QcFk/
LrvRv7zt41YHOFgseAqvrRpQgI0pawGGOVVp4UzIHNG23FNOKDWGTxtRXiB+Bcpl
1OZt7Ik643sJa6aUMHoukQ/vjMHBw2EBsoDbukyDuOwFV/1m+XgQ5C4ZyzeTlzij
tMIA8HQl21R2MiViPBNRbPHEp5biWgRv+jx8CBlERd1CYEFcZk/c7qnm9mHDpdE9
rxEmNDNhXr5izhjtLsMBmA9eREjOG7XL4oOvkI6imTxqGXYEutOEdF0jfjFM1YzX
GtmvOWl1ycRCrqXrfLSjWJZIUnHmhYUiZRuXeH2mtp6ABMjZag7FFJgl13bCTtWa
dSgEmaX1/A4lXxaK6NZhYGRnyEeNSUe9HYg0ghvM1yc2owIT20eWtPN0y0AobPVP
SeJoD+woIMXWpRAlsEH4w5r3eeepzrQaPg+OLNcrT0zvQEyFcFwel8/7kC/ZENZL
FDF1lIY3ih24QzZtbz1T1/bQZcxUrcn45mWqqZ97VGjMAoJDCY2kxqjAEr42LOdZ
XZAFW14YeC9CNeirCmbfZshmt4PVVqM34SdeOtLCFuL3Grq/rtvIIZTBv9YsqAHx
7LUG1cTYzbXdndU6p+i19zmofSeG7xSy1VWcLO/eHverObstfR7icwUzjxANx2s1
NH1+J8poT2J73jd3HMOaE958IYVZWPFEyujRCqJHp07OFRjMa/jjYba0Wz4xbNVM
Ir/NdPBdkulOTKAhQja4AKEtVSV5mkXqGvd5952Zk1I4gTPXgO7QkuQeImnUewC8
DgreqmJzvl5VChpRh/bRJToNhbMmBwvX83MiCn6WLEkffMgFi87VBTOep3oK7Agh
JxzXM23BsSfzHDMkjSK90tpgy5RhJ4xxOxTbJZjztZaKhVbk2xdSFQgwJT+lxuQz
u9r6Ie4bPxeOUvSm6T0PVik60JRLJBKY270GxgSzUtTLLCppv+Deriu6goIFg5ss
FmIewbOf1VUkDNMb7n0Mop785utBKI/3v90HyZmeih5olNkJuUZ4DI+Pe9NaglAN
yWwJ+UaWwVmuPzn4YyuQP1qKoN+Z4qkwIoN62D8sin8vYdI38f4Lu9+k0/LSuoO6
wujOq+zdjxjRHijscsazKL4T0SIy8BKV8og4pHLJMPu8xCw1ilGd3Sfl2ZcXRXQg
AhzoxUJdzJj0d0tFe1HSQuxSz7Q5tlZLtZ1lp+UmaY01WkceR84P0kzxRY3bOZjZ
RQFr/Sy1qscXwNhYuodPJ/REVbSjAQVmHXzFFnE4N5RJ9JcVNPGIVQMg0ym7fcJ1
+HWanO9B875RoNCjhdk+AzYZcFfbvxk9LCEnTVxI/hxea0obNEzZH9SIOq/bsh8e
o2JNrt+iTDJeFgjLv0a9L5OwHmnUK8IaSgniQzfJ4RYBUeR2UXPhkOLCx/2SiRaA
G6/NBPyg1pGy9wH6ttvzukXN8USXt63yz9ddRy6SSz19hltgHuokoN0SxBxEAocr
qy222+5HcVe+2GSXXJsgW5BWT3FfC52g3+zDmYN5Ux8JPjMbfQ3I7gtKowNfq+9k
DCbjdRrPKiTCCSFKTizw2OlL/1IE3U6kKYP0I/ovk25E0RKLWQggub+mUMXpXUuF
o1GEpAPwpo7eXbLoCuDaXdGA+HJZ/BUx1zBPcDV9ET5wE80iBw8nFjOS7ftjm+6N
7hkN0AR1M8x09OYNrXNbSZaigClUQ3f1FNicHtd4uYibIUz3TWsMyLUWCCPVHBvF
XnD/YkGDNj3IYgzWVIztX3RU0CS8UQrch5dZDFPeYH1qn4BsxHyhXtB+JLWxE1CV
IvNrSWum5CXlFVXj5hjCk26LiiX+UjhYNT/uvDGZdy0iZzGu6+6TB5ajRBS0+qQz
fMvFR+xLrf5i61P/IIP7MyWS0meJrFawfvWpdQsBkPxUvdZA0GTRizvOiVGJWyYk
5xCsX5EmJV7rKEku2mBjPN4MTZP2KsK0fbpey5DX7aTaT8WfgdUNmCz4e2yM/iAb
Vlcv9Jbz9MWAU2MimYQfaHv4LbR/mNmqe+B1wnWf6e9bjNKJm50yrKoJbM86jxpa
Dp827qePw3MadcgbKefjbzlyihzNnY/QMqYJkDdBhMB16RtP4arDuAUm8lEGi7fq
8tFcyScaABFqdPd7BsiJBpZMWvqyXqykI9gJE9BM8A9W2MJLoweCmTzyCcxog/qY
4TW3HitkAFyiETj/P6TGjv8pU0TG1p5SI8ifPBuG3y4a3s1YNb02j+TxJNlsImmk
DmOQr88XIU1hBzBIP/37vDEbh9dc9p3SLHplaqMr0QmRKCE+rxw0H36S4POvqifQ
M6SIh1YfmhkHSAnMJqOFwIdwkTONInJ6FRpxc9W6ispuwLmJ94OQQJVD+3HGZMpT
ZaTx6/UeqSDazzY45k5jYaeJQyT1Z3SFvv3G1GkfWgy8RqNCLzaTTKTPaa2FxPFA
P3Wt12E4VVzrYLbdMdJCQMpvBNsDilImUrvqWhmZuwizhLLFbjJizPtJCmuuuVi8
Ldkt6JJoRLYPR5G6WXdpikDsHqZMMWpbjyXT+yRsZeBVeQUBeyiI87suC+P9TUPy
2XJ3kO2GLltEfGUYKHS0+efM1GYyOh1AG1a81zMyS4jcT0buFBQb31enUrWMJCB0
e4sQgMyVbDZI0+meO1AQNWkUTvbRImbY+RNwBZBtwZ8LcoRW8mQ3sE9bjOQz5d0Z
GCT8QbRKG8CtKQInrVipJ26CGpBusXv3yQ0tcjidhbjLj9Rj45HAm6/0dfbb6Wci
NOhRdvp4rDycSdOVa5cSSTUz2p9/MK5PNAIg9EEOuPR4gOO1cFSv3KTE9KYB+pqL
pQcSAlmKcBfruAtdx5gd/soLVudxRESYj7byFnO9pW93DyhaacxWnoOoCDwb9dcD
jsQrmy8FqrEVWVgVU6cdnZHXMdWDelTIlT5dmZnZqVUX5gckdbzkv7zX+bUj7gtw
1gLEAgAhMuS7JsmRRy08AYSnIqIxzNfZ0XnfupGhMvxRBZYDQqFKp+/2+cu7Tuxo
7MNjCeGZ5g5Y2fdn4rZldfE0SbiQYHYcJHo+6L7YmikwcVb+2JqjD+N3X/NH2UiY
Zu5VTgfeuVUWqgHt3FJz1DU4hsx++TA6CVxmnD9+7J1GkT66EaAzPk7Zid+ImX/o
F88Z4ThP8j6g+dcnECwCAvoBRyhABXpw81pP09WDBl5Y+3dsEFAFhJZFhSZdp6If
u+INPtbITiZAA13vHTc3QLrXkq1YLt5P9fFDvkmIC1vO/CCnUqrRvEzkzn/QbNTu
FCn8Jl+0+rKvQIgJt+argOh7jhl02R6BZ5GshAqNzRXNZ8o+O7U5iVmvS6D5EUY7
ou/2og/Dei4GgU3J2P8iFOFqUJas9EyricPpaWXnyRRsZXRNcjj/98GwYEh9yPbq
hDy3d9F1LNo6qJCT9HiF0RmWAiLJ+vFEJo/sZSeROVXB0W4BFMhSdXfAtVOmarOj
luD/T4I2PV2PAKUj+mIL+osr7S6NPIprCwALaxfaVWZpE/C1Qy0/3dfTeLJxXpw9
+VuxFsZwmO/TYDTjCqnORk1zMlgkTh1am50RcBDrHGKv0TCG0+O+RsH/h9i3oZ/k
kUoiTJW2LDmNr74LmJymcXTaBa3S+uE9uxPG+FpD7o0V3RYkGp1s3pMMzsujslTU
ZARRITo5hMuofuQmIOPAuhW1MN5DPN7DQ8Ume02M3GQ4RpJzNNLnTQLIUI1b2KEZ
JWeSyYLrg9a8aTqvg41eXXM89zfFmt2aDxk2TBwD8Egvy+vkjYcFn+X1dL7jMBAd
jfpNeMrEIaS0lLfG4wF3un/XPF/rWZDf0sz+gPE99IlxtShV7XO8YrkOtWzZ7D1O
imXwOvO3lq3DrvukyzAqXA2HF5HOPxNIs3D2YR+syJhQLzMVSLwcvceuWSD13etk
P0AFwaYFMjiZWosr/RfXiLXRgWd65GUwlr7vjBvgA+mLtDycXhskm54fxhF9LPxL
LytfRe+SmnSIIN6acCLCLQR3cssKSCdHI/+tyILFuJzTrbuZ0h82GlBeMqAa9RxM
NRZouohGiJOTbsz2ZkLLMAqTEYOomGTXA0K5VikPNiy6EXFM6lq3674spJjgkTT5
Y/WIaWgCFOLes8GYgCLtElm54ZeyVxN0lsCPrJ1XDlefvSL94rmyrFf7+yuOQ0sk
wN+EeAkeOHtYP9zmRBU83OwK977004Dt8Et+gV28wmCBYEMSt+GBSoOmYXs2EdEO
AqXJW/YwqO5Xgf6wzumpQyfVSdaxcN2GrOWeNRfBUfCbrgxa8LBTZzi5r+UdquFs
PyOghFZoOpX/N7B4DhFlsmDhadP9gbKijLwL3y/qMvBfwYXcM4k8u9WxPPj8wo88
RbjE1Tkp1fwm89JYp1YTtca/10DSPcmVPzrrldbOwei6udady4+Cx/wXpe3LH9hz
agcMWd56cxegY86CtWjxCWi7rpj1IDlv2XkHNIgp/6IO16MCmdtF21jFGW1xWq/N
9uikir/WoOKErkbqoc2djsLgGgBRZvrc866I/bgqKzUk/uiPKySoPCh04VbT+SHE
0dY4fzpEjFNIfgZE7b4DRVZHpL4VYHCqdqptp1if1i0um68h6lhb2yCeZZGW4p3W
m05/+A5ckE35NKQEFgZ7Y8jznFYQ8CYN+todXViC4NmR0j8bJoZaYc7Ctlk50gVS
3VCpyDxjac5TXGOEkJ2Sm4OXy3UJTbpdrJY7w1rDdRRgxhxrwWfQKD2vfoHmn3Pb
xN8a7h/hDcxu7F93/b76K2oLFn6FUHVaBecAwgIR9TRMxtjU9wn2MKDUh5EBUD6s
+0MFQ05aQvr3gmbQ7NIlwbA0vHMtNZqD19bECiYpeK3inji1gQBlneoLzr1j4RSn
N+3fPrgWjUf7dOvNr6Pk5CiyEGblxtRMVqdEkMoELsAtMfjxUaMUGpb4c60xTeyV
HpGHPzNNROXl/BLK91npI2g6KZfk0mqsizGchfLZAqieGCMEOjRCNPX1NI3wE1MD
R1Mpz6LD0D75r/5rnGvWw0bgXZfswbcIqOk2rEbRcol7M0HrWKZabSdmwjbfYmix
v9pVoc8T4sr+sO7+yTBb0u1c8qDOGydLVjawGqmlbwTP1LWZnV43g38UVFs1qxmu
11U+TCfx/SEN1/1IBfv0bFHUNDu2YKzL8hwOF/4bKYrCqmQbVBfoFtOgwx+rnKXA
TruZmaYz7+ClFnxh477FNWdHfeHANXEKTVR+sR8LvrrIjmikwS4Y1Q0G38FwWQ5w
N4SxABDgjHjn/cwyxnQ4a7bb+DUG8zH5dQovtPInIRUzJU481ouJy5NRQ4YVDeO/
MY2s2Lf8clYUNRt18byyxeGU42AWfDhBdGBQV1bAmb6dd+hCALwdgktKEHmQVUJa
rrQAuEEyJtBhJE3XvYUfcPFdiSOAJmJrp19xxCJMDLR8ZT1FPztHt6MVWwMsPcOV
Qa/JJqEc4hTVoiUNvMXU5gWqldUdmbNEgPxgXrTg+2XVumKmUMLH/048mbXWbK5G
/NiNXqE5XrgklMSJw+OPujaC8oaCRtKoDZn2S+2QQDTrHoBT6RgT9a3Wpoad+KTA
FQqz6tc7JGdcGL9I4MJIllHXDApjVRu+miOQmnaVkgz1HJFs6KA44anUXHwEMHKl
FZ99NvCANv1D713SzpGPBMWhVrhu0JW3OY277cdA0wNXQZek86jOZIC9tUL0npC5
JG1twMfMBdsSQWbUxnR5kqIIMDbNT3gVgP6XEO6luI0trCD+Bh2MOwWebJGcnjrr
s3MGbpUZxTgBBFESaSYwRUvq/Wy5CZkinI71ROav+M0weEEDNVxsf0bniwrFs48x
SmUBzQa//J3EGSwdxGlpgEtEskrNiNseqel8KXDQ4TvV8pF2cbhJRjfPf7pkA2o6
3bauhz4xGIy/Ns9bjfTl17WGl9bkFzh13j5gd9SVD6wDzwEuIMbn+608Kw4Vd7Os
PPLvSOvzIKx/Ih5oKZ2e5GvCqnE4meqyMHZChq1nPpohPyYkIa4m9vhwT1b8hwf/
sLHgJPXT8v1eCwT7bdVzDliDcto2jrug8NNYn9xfjFOm0YXfs8j52H0fiLGt9CNH
S/C9dO26YcZoDM4m7pRh6jSljD6XcxnEQtSyJM8YtNH4xj9DTAvhx9CH6GDhd+76
Mr4wFGTZoZCKTqo5qM+wiWHqr/fINm1y0/0AojQoQbhiYS+v6FTmjTD3yhASCjWJ
K9QbZjXIHwMUF/gowbaG9ltxWfnw0oh+r4zrM6z5N3RZfZZIx9FU91iTx1bW4Tt4
pOhMpMTUo8YoBuWEykoJeamKWUKq1e8/gIvpuwvIZV+r8gkAoCopZZaoQJYrR96b
BUY+AiUM9H5dMZTysUE3CbhZS6wWjFUKrJbWV3ol2aodMSbUvEsZv3jSRDLjTz/o
FR6LjEmTN5nG4I/GDP+aIe5JLdv93Ch9F/0xKJvYBIW7SiUwXtWbLm6uy9xyU1w9
4D6s0yhsC700ucOdI+p0CwnhM6eGcGQpZlm0BI8O1pxQGH6OQ6CU4nmysVUlXxky
4lncRhZWgbWI08oM+m9bN6U+0Om/9f+NpIbKGnHD1iVqZHG+94/eTkhOEG1N2tvo
XC3pDPTrxFNbsO12OeXAv9elk18PIlOucFeo96NY7DaayAlexP7XvktZsncq1tqW
PZNhCzbV+WjssLgBDW4mW0THMNB7gUY+KfeUaj3FMelqU2M3Y0c+pi6x+yRKSpZk
9pgoJWoMSGDpEeXNk5OrXM1AGAjPZDpWHqG8/2ASv8Nc0tlyLdJS0sFGCUIaCkx/
+EK0g/8zDWcIEw2UrEBVgopnSHs1qtoL2OCghhUHNpSpEtKZZTda/P17hpdY6aT7
0jRG7rP/q81V+B4w2h264I4Fhu5B2+kYAx8g0a/96cKpRd6gD5wooH4ySdx1yNaN
62dy9zW4YuXjyMVuhtosO6UJJosZsuIbd6lkuMRRqpko6+jmTqP9J7+iAMFWRGzl
7OlxcpiVpyKxfjQXzWBPiaXjvN3ksc/d7Wsi4re5ZFYaf5RBRJed/Vw1tKEGs3eb
V3x/gXfRIeMwpmyOWMazMLWviHZ5iasG0DXSGk4Sa1gcinNYsCeMLRNUNnUgA6En
q1QgOVO9HVik/L302zhyhPUQ01eU/58i4nMCS6ISC9xTYoDiwXdRMakryyfyyZoG
VpRZJJzHOdU60d69PBxoy2qRD0mYiTOY4MNN9eZN9MJyYMcOTO4Dsp7dv3yTJPfA
opNCaXMxJCwDVAYyWSsIhs+7ewYeAXoOoyZ4p/GDqo8YR+jYZyemOikol3GV80yC
CtqCfAVFnDVancqZ0/KdEEgGNg3ZjPv2ee1AjpmLNWLRFjs1gwTr69TYhtWVNtaL
nFZXe+v1TP/bhqZ4CUg3cG5Rlc3DQrA8YF23UtabiGIvc1AeshBVZgD0/JhSHxsW
HdYbgj43nlXDzBne3TfJbLyA/00hHp00bdLDZa7+pl3ndE9WvIxjhx8vY9Pcx3x+
9LhrdqH1vH6CD/mQidwi79GuHIjw4lBreNB9OfLzPhND2qGugSzrNh3OD4SzzPOo
YQTRciRIwGMHbJAjmnSM7xFp/tNhp8wrh2Q24cl4n83wAsIN0hZA0jRzmEBd4RiZ
rkUKXSDJhKMAkksMDpLYgZwr2Gb8QF5u9usft10Vf73zip3MeYjP7gaf/Lt0PhlH
/RlAAXeXcH9K9dlmSLDREo40gtwCv5dOBjpEyPYfvUvn/NGrIzInrPMBj5fYF+CN
TcYaGXnYpRfSSGkf5yOoJFM70TvmI65BdwJuuGpNCs9VyQbgYS21ok8G65a5+8Ne
VJior3DOK5XDUUIvEtYtQrEhcm9by7azTdM322R6qN54NEtki2Md1uI3KsW23h3A
HQsXUnnV8OiIcZIan2HnNArl6vHDvgp+g+RczZUuJ/tGRoxOoLxAQCbNa8G/bIyB
hQhxTE/+JSPFFAewg5Lx/l4AhxIugxy2+PesH0c6+ciUyXrX4mYO3xDvryph8vx2
Y5c7pQUySNhZoh+47usV5vi6i1FQhn5Ja18CTOacsJmsfUXGcSmEFpjVvtmSI9OT
u+WAXg2eCgzVsJieGjfw8lZhObVAoaduzBbLwxym5XCf2sB5HvFqgpEVoBVkxTRs
UB4qMFSdKxs8TYalqFw5S9jPnyu6siDZJPGwZXqTZ1Ja45Q9eUct3spRX84ISgj+
Ddkx4GfkJEBW/5hLn6KKfKP4ha5msWKoDJsTLS2eItTzmKP0I738ygNhKQpWhpqA
YKT2Ixceavlr7VgV9Kit8mECoM/4IaHaPn4LmECRkSTTlcG4CxrF9U6C4SuQlJIi
347oFOv2PJ96Qkd0YybhIGlhjnDe5GOIUDI9tjjsC2jz/d37mLEfcLzjYEQaw+jF
JwfYDcDguh6Ncr2y7cKLf2WPDBE5cr5BEZ+ytEl9H2L//y9Z9qwo+2NNRN2aq2EO
bd9nZ1/iAq7dVtmdrEa7rfRKMpkdFaDjFDdssd2QAYj1BFpO4i00PMT8E1ExBnDA
I9+DgpCNk+jlXHsRSdLkjNG5Rvb5r0Aqi9TzgSogq1qV7C6MOoIwXr32+FyxfNqe
PIrrLlaCnlvvtEHX+T+DPep2oJHN/2Aj9CgOtGtfPJ3WXuWFMY8LNUYC270wHQpy
Uf0CuOMglQS843wQZEYl26q6ZJAdXMe227tIP0fDHoRQG51R7MZDdnPDvjLpKP44
6C0m19gEEngQMYelYjQou9Ch2D+CEpVr77JFyfo4o2A2KGPp+drb0ZJrN/alCuEu
ORvlpX1M0zjOyuIjQvD2Kt/8HDTxaSWl8uEi+slnbWvqDuL7Ig/cLtzYJSKheiNw
S34CNeKxtJvtmJIwUN8DOZlrIRlAhHM/c+QXcieYtG0PuimH9VQPioBceNpU2gZU
i3sCIkREsFyw3jeSTmyaDIcA26PnXYlFw8yvssy+M1sGYblmCN3Y2jIwQcyFb7ml
omRi7uXhHA+L+NWNRvIGa80rcy4F/T70cyUem2viYdJo+vqOVdlFx57irYpODLHT
03m2fTb+KAORoXzkXz8iPbdFO3u4+cKmbceD4TMWa1hQ2Rxk+ePX6ni26kr7hi8u
AlyvXMQVyahoiP0FD7L+H0lSoryLmsCxStQFKFXmjubrpFTB1lT9/BO1eHpYWjXT
otbdV5K1wN8u1RWa7ckzvs5fmktkwV9Xd+Y9f45MqJPRxz/LJGcl6Jcq18hLtFQc
qybjbkqKmPf7oWD+VCTk0jH1ful+NQN70B4K6nbfTa5Z+V/yiQ4ZFFk/iwAfJfUc
ScQIDbFU9NbiKO5tqdqbGXoVrEaN6y+0Iya0+Uo08AEtfHf9pQwVl2/z+V4eZPdb
L2fgMNmr0z/cUL+U+0SGJreG6Fatzq89ABC4Jxplr+cC2iZMihiZepWh5U4vZBXC
0GVmBrPvogs2JnVlrIRdUagG1zNTvnoVQo3DBm4M8QMI7faLNCeKs52M2KVG9GIs
ab7trAvPWNZnXNCuwUTC+NjTCGpQFf/Nfg6aD+Pk7Qy9+tPtHm4b04OYr7WHLFT8
0bu93iboR6g8cOFnyrzda82XuxYu4OKtp2bSTe3ZWfhmqqHquuYeFCw8lgK0AFEa
Mfg2W+UCgsTQbv/2ssAAipFie03fz1p9VaI5iDOcIcz0eDIAMmTZdMwwkkch6noC
yPpDYmFOEKLe0e/xV2EJTRtPDho9v4rK6e7Hh9BkImyZtZ419INESuqAQIB2MQXZ
W31IpwxXymY+4Q3TbyvUZireIXgYIAraybNvqlhW3B4SZtVhBSbNwSA53TMyrB3X
iE05KdWKdvcKIo27bRgDMQqfxnB6ASirignklN/5uv7hpJ6jmeQ+X2c6lFCQl/fb
1QqqAC2cX/mipdCIWo2kYKiZETsJUtgSBGIIJbFvmO/hj0tk7knnQjJBDEKmn1Jn
Xg6SYjz/GZH/ad7Gz9rrm6i69YaxxFkICiJQYg/yIyI96wy/HL7pXK7mLibu8bwx
bTj4lgjvS093qUn58hBQSD2tJkS/fdh+uxvtG9C35P7l7Fmk9ZZrR1u8rrbHU4Sm
0vioI2nUff36f7VRn8Hju/pEXKrfWfdE8+25Zb8VSJoaB9bDrWbVpPQ66otG+7wC
eNJAx8i6x/KMeiKzLMvcjOt2MHsHE+Z3S/F0HloXZZuGnN4+/HmGasIGs3/Ngr/s
4h7wShoalrpzGl9jpSnEznXw04DCP7gYotTnF2ZO8h1pXV+8epd3Zwt7wLDCZtYa
JL+7gogQbS+J+ff6fmK5KJ2wKTAs6ierStLvXepWIPfjgOYWY/hkQfNh9QvYDASP
UaTOi7cKqOePg016SP/o1YRCDBv2ollpLn/OZ2oraZF8zhAzTSOdUQxhVbBlcY8N
VtuPISMLUjkxD+Q7auozPMgx8W1U5CVVcb7Xg4Lv38bx7nUThMKxjRaIXf9xXbIu
cA65rClfKubrDUCOz99CFshNGjgRPTTUZJjMWNWlNL8TelKVZqYX5MBVLYhuZZoL
1QVoWCJYGGNOJ1pnB/gxML1sWgUVdqH7oILe/ikrS+V0kRkNwg9pdot9Dq7wEv94
OwcKW4EADHjLmNaOR/JTKx/W+33hWoNkCZlaAbid16QPpJORDDZL46vaLQXJAXFe
Dd0M6/7uDrJi2p7WJ0vnGhEGb9K1+Kb9bSumo1S883pU/6Vy5pYT5y9K+k6k1xyA
kX2m4P8zJ+ddnP1obtKoM3ICTDSkgnyi9FvEyTzQb2CLgRnDkQmwuO5iVzD/hOYG
Lt7HsWIVudOtW5fEFcnJyvJVbrr7oIcF+T/7xClLStcXBgFMzKlwqop9KlnETibv
dEtw5x5OjgZc8w84k63WRtNmCsQs1Di7tD6k2csdC+rfd1vBDsbu1Dqsmrf0dl53
E+A8bAvquyGpDkqvGPfze9R8CKDN9KgbyEdO7HiyuSZMLITZIpvfqViy8zzVddnC
eSEZySpWzU5QSar2XZHfyjwpaKBzCGjpBusnG1Hn4Js/BcPHLDMTBuHGhnbDzlOk
WO26puXTRbchPnIAz2ky860mzd7l2turI2e4/B9ttZhD2jHh7toaxsHgPpgT/mP0
+r00unccRIv4zPyCQfBk/cu5VubM9HZqKIuvnzu11zFQrfetuPHw9ugGTyfNDpui
XoFhQiFHwEh363AbrbcRINxHTQASgrTC6emAZIIJxIcc+tv91RIGlFHOKEOMFZ2G
4+uZJlFSJ4rI90o40YxJY0/kAP+f5kLaENjnLjfYWhDMCrMIF7XZfAG2Dd9kKfZS
k3gIBHNaXx7UkaEgToFEx3I13OcZPtP8vOWUMPBLPKg+TnhUxMa4g3hM3LQ59MxG
Uqmn0ZUnqJZOnLdKMVRWkc/RybMAuRIfL4ejFLMRtHS1Ly78daqrUHDKRCDjubCw
wTgFiq/gPS/fSquo4Sj0+Jz2CgkZzNYxBFpoYZAMPyjDVhNSZa+YOdrwYsgbfA8O
w7kOuAwA5CRUSbmwKus2QiFoqMWNAbB1cpQqUynrx3qYQvNA/q/63BzLtvGSTvvw
yg6Mv87Bt+2HY9rJVdDvRpyUn6AEr5G0aGmCbEJdvQNW/2z2BnWTDXZh9SfDU5bF
fyfsXtj/NX1PhGHndDSknPC8wn2GtUZ+8ooUi1VK789yg8LUDplwVR9DXazEbOfH
8GqP89rD3P6pNDO0ITMh72pHmIUXOi9UqlXxyeqqABUzz8WMLtftaiNjqB6dcl5B
C9Vqr2KgbiXkzRRyC0qc9IIeRtsPs1Y0RNCid1Ec2k3jFC3E5DXgiiMxkWHDQfiP
+PcxLu+/BJdePb3DyDRrtqT7arReGZImeJwlTWhNMSN0/ocl/4AmF9tFZ729NKOU
rhQKRqKDGfN2Qw6ibv7N6IK+AWt7aqjozo8acLc1MQKV38yO5bvyjumCuc3ANNvS
sMCwzdUXjlIGme/MNVCPDFjw374rPxa8W0wxFRO071sIa1GoO/5bz44sEW93NARU
9jEdc8dPGICNwde8nilBy5+sfDx1ME3jpZW7lqhVdmveJVF0Xvpsr6LkYexDkzH4
Jznc/CFi+oR6cxYrImYhkoaJjLdxsDMwiMYkduFHSlLVXd3iTgRJZq0HLkg99l4k
GMhNnXOz001hIQYff0i0Qd/Ogsac5j91+TZt32DYwniQI8r2Zm3YB/BQnr2VYuuL
3DxUBicCd2hoVxdFw3T5qmJPS+BTD6o8B2qErdv4RCKyOVO8TEnPb1e8HdNwi+Cb
+gEtwKcyaMLevicPDvSTyGW8gqQCk+04J6vbUgXIKnUuYQXzJFlF9j9AqKqXDYX2
tC1yOjVzYh0no1bVBI9OC14DAO4EAt6VFJyXhuK7XEi0JyowNtGvcgD8aHucURxk
Djop8rlnWmV4FPOHeUm6yBZeJ4gg+ZC5P2OpgxiKMVbj7fmFdj3xyekl4/94l1fF
AuPsIEpi/xmgEVUoCqA5ys+qTaq5cOMqIek/hjHmtc5ah/DLPasgmOI+Fy32yIIj
+lJO05ik3xmYjmXx3fQ2oVbzMXLhFOZd43F+xOs6Kqrt8Eq48aqGCllyn25O/7bo
n9dIk3DRV8JpELEjzIrziIUVbFQATVaxRKBsLW4gOkv9LAl7s608dD/g9yPhIOEc
USjgyxdrt2sW1Md6vCWAkCNFBBLW0wi3+dOB0zeTc1Dh8TbnrRHfqQTzvZdTiOK9
uR3GoEUHxPeIhmk3ZVqKIedk0HgQhFXy3EYjlWIqkf5dri2uOD+vWm0an/vicQkL
gnssJYpL125kjE0SXxUFIqSoM9E3Pg+LAPijE3Tb/XZjif6rz6+x2ZQD5IWOiBeu
QgP+ygRTUq+f6k4rUZgFQAiza+xNAV1ldZ4LFBmzpUl6WsctOqn1NKQqQAVY84hO
4xqi/4EmbVa3cGpWPt2esjWU6dBfujy6CDkNJ8cQoREmaIYqz/fpbWY7HAJ+SLs+
vc0ORWcnEsi7pflDvdg3kmZUnJPZedXna/V/bDesNa98a3Cj8qTNdAPz/ToPeZim
AY3eWTzUZyzR5MTS4OrcYwCLBB2bf9HnPvofsJiyWeSNwlPuC+4FHTNMFT/4AU6W
E0UThm86OjIpS1IFNIwAbXGE9ehQZlAxvFXa3JHyzd5te/Gb2M8CfsVdn+Hkhr7U
PrQT67Gk7LklJbY+Ra1FqhSuCIRqjVndNT/PdmJk7W1CAgUK/MwrOelx8AGo/uKd
d5FGPJOPThtumPkEKF880jYHYDXOOJSC5Hcbs2Sepanr1ysim9cMLVS2/5o/vKLv
VsEb1HhjxkXsntrSrsM7+FPeW9VTf8NaBV4EAUHhRDgoYBgtHGA9IuiJo1wtKnvn
shCRXG/l/kuHFUn65P/ccNzaMfypuPzPNXzQBAsAr77ncZtorBihg/XXGK84g50r
hcVurgLcivOxAwfPmWAn+g0NCxtXJmDa8BcBN0R67nYzTJ4NVP1AvgISEwY364rs
BmM6xNoBSFJTkh3sllOKMqVKIznU1Qp9HNu+o5yBRiy/JJv1M19dy5QcChIJDF57
PZq/9k09hXw/q71GtLYkBoJMEkDR4IJDN6BjuQzHWhMm+oAdCW7Vd+ieTB5XOjV+
B3rg3yHP/msA0EBRM8rkqquHgUPkT1REdXnT42jTbTE+DDzzedY/x4cgOvZZAJ8u
vl0psBjhlQinizY6/oe/HXnoCIx2sWlkWFE1RCerirM31F++W0sl0kx6ZpWc07gI
w6IcWuTAdzy27F7kU+H5AVKTVDrapucJdouhNoJ6Nqje+xe5xzde5rIEvybz2sdr
qflCGFaBZbe6OVNbjn4rMJnBYbzW+NzU4H2SuOME7a/cICqAITaPB4vdMm4ZG0EY
OHzwZ1QtjsRUBUPqAt2o8Pxg6kqqZotqX5x/4zY+KQBuzm77NYjJxEik3P7BCRIY
qK80bChle1I2EstgOvqM/MPOzj5wSxj6Sehkt2FPLMuyDecVlG1tVyqzA0wOjn6N
o4txa3a3u1F9+9L87B2eLSHJgTpq8W+NACuAQ0PbUL4zGzTht1uyl839IcihT80k
vNIF6kZheKLnR6GDoyzAHfDreCtv2VFk/dfVG0CoUNK6BqbHWlpPIGy5sHoLCyht
/B96sRupIIy4qoq+DWKtdo7wHMQ0YTrf+ciysyb0C2j7Xv3ku1nZWtYpiSuEZSP3
nL4DLl+BsOfU/Q4HCyGqHQThsB4ouX7DpPzQ0F7CU82GVWEjoLOvwvGQV5o5SmCV
1zfdMD5Vkai3cB4nNuaSaCLN870EuElGiXjkLmffn3jfAMIpDVoxN5erYUjSoGfh
oq8pkWJ8dkya5BIerH+VZh5geRFPngZSCbhJerI29Qpdj0YWf8EsqWC7YzegRwXt
Fy++YnBQyHZg3lEk1bX41XyZ67VBnzyxan/MNo+727SiCkDNz2hZGl6igz8wEXnd
iscq8lPgA872qxppe618Ki2y18PEHVNXRBq8PQcUS7UywrjS+IKe82YUS5PIJzDT
BtLDgfgOpgu7Uw6X8oR9M+vWnh6LJdOILB2WWoYc5qoxYfuKW7KhQZuy9CLyR2Xp
WTZFBUCKDSbHuxG62OmKRjWTXwvGE41takEfvdEG7l8qOXDmqFSO1z1Y1qR3LBON
MyyQASIUjGjQOavHcwgNTtthcHeEPKkaEe0rckPHGcYKC5mGLxWcWRsyjcLU/Zd0
acFM1C2pCRo3nBjyEN4JJelg5coOQ2YFbIHf3DdgWN1cB25hMewwF0slUs33L/4P
z3JK65eXz6QUYYqTJHOHt4KFkTj4weXwck/iUowYamEdwVEja3kC6xwWjSlx7ACJ
yTBkyWtr2FsG4DpnGaGOpTtAEbwElP4cljqGvUXbuggiQvsfY9GGoll24fzyGHPI
AInQsr6sNQL07NPnwh2ldabQz/VImkVE9b3m5/1WxNd7tiyRoxAZn/hQeKXqjcgp
AcKzsih+QlfJbE2JTqxrJi5inrg1NB8CD4KFWrd7l4agN2f9ABv++zorX0UrxR+n
b8xni2l/BlblRs+oDsWxCamaBRsqCzFInkDUd6K1rITqmsAhF1hXSJy0ibfcBiPu
5V7rI7jqAC+AQ25uFufNT3j48WKL90IrrMaU9fSgPwI1y7VvTxmVQplMr0igrFJI
OqsFzJZ6mvVkx2jZgFcknM3l2S5dBdu17OLGG41C5LrtiZbwKBmFCIg5b6Vmvr5/
AxPsiqm3MjwIuw7B+Bx0xpDS8uN09zOuvIkZ8+N99lAWPVvscHwnAmDPJTQGbJuO
WbKYhgYiKx9uRYcBzg+iwAVnNDrEiS56322OtUBkH54jORcv16+Wk9w6Bpjao0x3
Ix3T9xawxw/orEstGYq6tyfXW3X43Lra2fCg/fnZyUcDFPrAXePlkpsln1ZdjwNy
vLUrzXAg8ppQFjgMibyeJbkqHSHImOpevCURPj3OeLywsY7N1I/oHyV/rn7QDxfw
Jo5rvw+WtQLjcKQ92U+ZUYRw8Vup8jpxaRMTeER60JP23rOcznvlJdAhEsGzfOKO
V9cKcjpH9phESYu7W3KZuPwuO5K3tTZGRCKWHCfxBvC5E+r8gA7Od7aSs2kTW1Cd
UwLTS7rU7qi4Ai4MfaeYIm65122dicvQyAEp0Wbvyomzla4w/jB0xoF/HVXdMcvZ
1Q6iY6yRPcYX0bUUGnCtqTwEhen9n0idaRh4AVoemwG/9xS2kbRuRUaYMsuvbOnm
myr/ZLfzvoWp4Atk1BAUWijU0voAxJk8JmdCKTpnqonPoFFrIO/XarQrQjsScwKy
6X1YcboAmG+z5UIAbYl+7Yf2zpFv1pKpZ8I3xdZDpRhSl9Ujc82Ps3xINWT+27nW
ukYLmdHNya3TgOma+32aMmJ/nRGgE6TypyzrMBEP2I11Mu5hRPYR6TYovHCY+qHu
fyrdFV1FVjVJJLovRK5bjEpW1TXE9TpM23Ygrb45lnIxqyEC7gUi7zO2TLXkTeOs
mJHXl2aCTFndsEH33n8lS7u8pQwQOIB+3W1dhfbzqzviVGy408U3rs9fZs4HHoe1
kZQmReZ0FZz6WFIf/C0BWLKghEL8ndMe0xV3+kOxzEQiEzHQ02i/SUJ787D780vj
az2HtjjEPPoVU4cp5ZEVxPdHcjSZx9nFgJKiUiUUnItmUti81wEhNAOFK/EbV+x9
BG2II88LU2eaLT+tl0nYP2ThGkAAZ+ErtHPHcBBeTqyiCT1cbBCnCsIybUa7OhET
wTkFjWMIGTK4ZRrwC4dBzl50s1k9tFUgTKSK16RdxqF5oqwi0dM79VGJsSXWYGiK
muSUVFESpLnlRetA3vKhvcYWIorTeX8DYJWpKPgU311a6sgmFT4rFbZbp2KWh5tC
0CoejJ6JhvwHmlEIhWi3hEk9MgDs3IHCgYGP7Gk3NKbuBFw22T+LMuOJyT4JKJS3
WL9J7B5bp1XVCwIiSS9rKeRTLxgSew5ewSVX+np3T4DL2jOZswwvFqZYAnAw9scN
rVBX3m93E0Gb9fpEKJAz+rEWqBaBH0cC+O1GycunSON7AyHR7sLiu8kfmLi00V0h
Ui+xoFN52NFIgziCbIMv7siLdH92Q1hHhEQ37g1NYvqfkVe99vO+VB4wBWc+KUr2
RzNtxhWvs04jRWlfEg9gqgBkwLC+ht0Wtw789SHLSzgu0wXXjawok/KZ9Z6lnH1q
DVYoW/BDSD/HtT5tDDk8ru+VBAg0N/moliKVNXt8wlhDw8Rdlk4io236tIdsEJKF
00XoG5rZD9ZzGLLyvsHAWlmlzb5r0yw3IM/GYTtpplRFrSBppk9g2Z3qxo3b3viJ
8miKwjVjo8PxjVJ7/rzCH/XCDIHo+WJzh7X0xFUQr3KzLSY9SfsWTRM1IQNuYrBw
tDZwwQhhoVioLx2mAPHMXmM+W7+Fj1T79coQsST2wbvT9QgmwQxJIaKx4Ah+TcPh
hjNG3iBHYh+jsk48UUscFTKYAo7HdfaxEtCkW2POIjLcp9BB0w3B8wsLmAGeCxfT
Mmq/pSFmetFZ1080hNGqYGvpAXGNuBD73ULWpPVGbIlvq4pDWgo2etAFRdpKEKK6
EjGm9RxeRMapzPnLMCcuGwBB676VRJD9rwVVQBkNFAzjMTONloqwLmVu61vALvwe
2drKPRIWmpqCKWrhnC3mmiuHAkCzU1WRUW0POuMaUpbmC9Qf42ocrnWHkkYrF6+p
6t1XpbQaQNwGiOS1DsrSW6VgsjkopvxuPpXP8hFT4Fkbv0x6EqeGW78SFhKToU2J
yEYuLdEQzqmNbH1vgdzW4emTBL3lfNYx8apQD0X8TOWqHFzJUXPniwHt4Jw6um33
7t1qL3CdmI5fIPGZVNHlu8IATHeVjFszNfX2AvU9Y+u3JJlJaWj7AuZojgDoezgS
Xgb9GGuKebEsxn0eQkAQ8HZaIu6ikS/vPbZNxKmpdUyQEGFQZKsgDTZHce8IVrcA
LhOJju0BI5C3BuHnYFJtKSRrsOOIU/4ntLbvc29rYTBgZsmldyqkn+q270ltUDrF
5FkJOQ3QkrsKURrsW0RIROriRj6bfYqJR453Z+s5+QMHpAEFr+ZOO5hXrLkEm+9L
Jlw1dm+jseTDAxvFL+sAuPkE5CEU11aA1rZFeFrs3HwRJMHUH7HSmqWotqo3AAMA
TtT9briSha6dBj4FgEff6uMPmoucqGAXtr0H0sP3ektr9dnAnu9vwCVenVCUXt0t
kiUeQAHyoo8Vry7Lf9oLbr4AYh9g66Cad3rl4jHHnLpQFALdnbrg7CJZIK07fjkv
XvbVyHvzZ2a/eQOaQHbYCDA35XAQxdk59foL3E0R3Q5En6aJL3l6c78LyTTpung6
mEBHIUARzfFSe5Spk/r9/ul3GZ0oQ2h69O1P3Yopr9pccpdFQSjk0JYrmEFofzLL
0yJrKrTVa3tlfk7h0n7ngrcxTSnhL5zWkZgQE8lleG/xfzmxqOnty0WYuHQbrEmp
LJ+zju+KMbL0x5FSXp7LudlKjFmt65rvWxPPl5i94Vdzxg2OBmSoPB8KxhVvQRDZ
zugYlZKMDQJADkvUMR0mLZcFJzz9b4voYrNH6EcByrVAYkzHRXzIN0vMW6WX7a60
xFI42CQ9S5uWS+JhQxPUn5wHxVKwqulNRITk8kDnhetJpDr1pZt/FCCPbxhjJ0O/
pXLwBPjJdn9NtYVJVCuk/phVPhozHGIH5FSPweEDNnrNQJpWB0WmpkG8zXoX8PUx
QiVMvqVZR4ZFBeunkUzP3xAm6ttThYkXiqz3ggTaAzL+8duXMQBnkSQH9w5Nk/ik
OBEdTYqukLCRI4ZEQMnURfnviGTBGjuqw2ikbxH+AdiK8K6gkKjp2DWBrDw/Q7JL
Y4D/1gY3m1tH8LE0WZCjscafizTaPmVy/bO6p2pw43xOcdKjqfMKG8uKep+m/i60
zDp/bqyDK3wD/T2iV+vxjTPkITruAvbYpwPOR9ROGzjVG5bsD/E9et0KbrQzPiLW
MjYKnm9zMCWqq8+j4G4VYc5LEgdCYDPdhkAb4ESC/qadqSNMIB3eCPaGWL51WvYm
qV4GQvo5FNs24YOfb5KfH8rvJgtMBtJwd+ksTGydyj0+Anvgw7q8Bqt0c1LqV8zT
PS4YOasWQx6dupiGLxyNpBNWeyYe4/UAMn8dkf3r9wTZ4pi77D1BHQqphZ3RsU4V
aGU6MZ0pDqPe7HqywMyioJyTzWld8n9wd071FncaYJ1ZGjjsa26MxKdPCkMhQND8
QBa83CeoLZ4s9H+xM0+l9y+vgFNrRCPRzKf0xgcVasBe/R1meSqhEOPxIH0oKjuO
9XZgjmjKkvTbyTYgkijCDIDOfOfw0cD4q4tLjEJqB7cFUHSqeyg2P1OxAGVHHsnq
tq8sIJELS5Q73K1bx8jb4z9yUngYXBAo8Fjd5oKfSF/BvGkdTeuI+/RKBBfPcwRv
CxVZqoXJtEVYidXuUAn2C1/yx3zH8HFXjcKg1UQOOUHglLFDnAzCGPnA3aeNk/Kq
uXCXiZ4itmb2d1V5oc1SrYlOHk0X3SHILhWeGMKmjIsAWgQDF5mDFZnpMhHMgzT4
oTmVjM5Pg/Ao/3mN2+KmlqP/mRfAt4+rlqcHyknIeDA/ORsTHw13hmdRpHTaPEBw
2M9y+FcHbgO/r1tLj3eUUH5MMc4/bPz98zesbiMS2toEAj9glO1esIqxzxDWMSW5
J/swj/6fYSS7FLh+o/Ppd+7SRqVRDp/zr+p3OLUbv9ivBZK29vCQOOKixVCb4oF8
8WRWcCptCPQ4I0xQ3Bl4Yw8qmc1I10OnpjDIwdLq88AAXCEpzIRxAWIKnIdEhdsV
4dq2CsbZ1tR2KXQBoJNoh1dDkOWH5CEy6nceuPHpiPkgreNpouht3q4fUULJ61Oh
Ob/Uewgyoq2Bm5olMiHbg/k8pKITtc0ZusLkSw5V+WlDOhnOhv82WUXPYOWnQHK1
GjbH5ncU/poKv9AniqFv5qr4AqWoUnTN7hy6yMuKOLLnaV9NvvOoYF6Scx7cZYmd
0XvE7TkC0R8P1ny4gHJW+fpWV2bYXQOmFvmnQ94lJauEEnZZgjBs8cRI0A7nDGso
m1fGESqvelyeCLkt9DG/F3U8wsOSnNUIHXrj9qbQbi6EfzbARgSJSy+6ArEDlQPc
UNfO2X2a7sd7eV3kmum0FR/zYcbnB/PSFg8tl5Ajlic6tAQmqllCvUs1QGVwYEVD
r5+McHnyMYshqkU4qNSCGQo/JIs7k93aGgUtiaapF35Q60bjimFdPzVjHrAJ9Ce0
HYSeOHTKwHUPaxWTw/UnpT9aKzt8Z0rdWbpCSKOgPzt4N1tiF70RD7epUpIi3VQt
sGzW6viPzgYluMEcPC8vERZhAjz9qBSFgVFb/sTwJSaMJ4koSMP7ud5azNQwU+V2
dkHstpq214tvMcbuFozPBwTFpV7ljy7XdYaFh+OMD5bSCpnCx82j4H6XtE+uft6s
ZWP6kRwn4dhMfHmGNmj9PhEaR5JWE5tX+w4GY6nQZsGNosai0dZPaZr8RL/FHRL6
vYH0necRkDlYq5ClUHUJn+f6u6tj8M9Q8h9gLUvRam3btNate4T3/Otr0+9cyjHA
sMJ2lTPfflsx5k/2YWMgv78J5TJB7bSHOo/7ieg4ZNOx/tl0OQDlURHH/Nrb4NhF
HXbQSCmw0NjAF/mael40KN20Y/8tjhkP03HK7zidM+oF0k1AKVS3gq6T2X58NEnX
HtxznARH1MtoJMDo83eVIbb0fWhXI1YPTtIxbh1YR0Akj1jJK6bKLXnA6UaRtfzS
zchuw+amISPT5fmT2Yd20AcDRqpN9nB32gMwtn/QQvj3WoDnVtKdP3euI0NoXnwr
gmuzOotm9G5lzLjzfNK69zl4lW5VN2D2Y1DvZsqbP8khKT3ZjADkc7Itx1Ne30g7
0UXlLbR0B/eSvoob7Feb8xgKJ5arO80WZJaxzIGBqSXuzzeIZ8YQKoUkv6Pb4A27
Aad2B0+Ydac5brW8pdu+zgav2OEU4J8uz/NG2xaMWd2Jy21vNHgWLJ0boSTg9ODd
MrSbTCf5tpCcw3h8I/Zh9Q29A+JJVQrSuxK85LaSjY2DUsg6cP91plg6M70oj4pM
DHcPJ6xFidk8ZuEOt0HLAXLhrIC4mliZMX2MOXZ3VnWlGBZ0jpO9cOMUZmwB8FY8
I6rit03VqjrQX6e+czrq7XA2hvkanSA5cYB3vN2yxDatxF8G5cAkJANIpplyelDu
elorKKcg1n9jSn0oEgDoHS5e5pHNqPTRAAGWKwHQyPX6ecIaPU/3jVWV8jfpoa0U
A4GXsitCzxm18pR3XpakPMCT014nPWekcofp1wODip6l/YDReXwNdrCfN7x2K60H
pmkccrQT/p2j2y4cqHpXvbI72c4+Ecouo7E+CTLfwRFhA5p5Sia/jU75J2SwkK1b
qm51L5na4pMDqSxiYbezegkqTOJW3JuKB9abaSyZYpMdtzExlLXbvuLCnySk6MH1
60a7dBqRioHJHPK/J4RqgqR7DQ3+PpXxWYEpCxhTSj4KNmMH9sArVQNgdp4On833
FmfBw4cdGlWxqkMim4mLW/Rpkgp1PAJC+bZMJG0Cj7Gq2KyU+iZT8D67JjJ5f8PA
IpP1NtD0QLAlPL6l6vrbe9wtpzROCZ4x10/HWzNTJvDgOMR5Fz+ZFojH4Wv2hYXv
UdmOkq9O/u5oJMVN1v55Z9RX4pUmpsgj2ScgGb0ZuEEsfLSdkIlW6nHu9AuVWL4M
UomIPninHcTkinSVjlIYaDM8QY2+RwB+7OSM6UO02PIgLcympBVIyZ8n0gaQWF60
0ZdfwXPvhTWRahXS2lbIG5GaLixRBaqkFsMvnyd2pZyTKhL0Qt0QIy6+rOg+H7Nf
sGYAlrDVbnF5WKiG93EW++tqz3gXnR+9vBHT/kTBuYuMQJV7DWk9uLzAWOAcf1ZN
ZyQpmncA3LJH4/tIcAncM9S/NM4lWKkZ3SD+f2UhiBl/Tg71BKZMfBWD9gxi0Ku7
10DN0t+OHdEuibFQW/VYeVaKwIKdOSrFmL9+6NsxvR+ViguBSmO4h7uiQYvX5WPo
RzyrWa2ZmckkClYtRstpbDFUUMupEMmsTJx34V1QG8Olpy2pSYEP45BHjxUiuRYN
1VXFact1N+d6/N9SsmXI6Gus3LzBDo4OMkWxv1HhVcNPee47KcmW1RRsvyCeqIKV
yvpSLq/XDQn4oFEfnRyuxdCUtNmu5jOPD4xoz8RFQPD32eGiZfmMxP1LxeohG75e
ht8kyFBPYYgpsmxdSGWxH7Oe09wDk6bMziSIi+jKSVTbyeqFKOLsEXpITMJtfvab
4hFBrQH8pURkxiT2RSxgZZ4WpNtvJn8f6423TBGsh5UJBpHoX6gWj9CK4khvRSv4
PsmX8xvEX/n/vzedFIMaWItGhQAnAzlLg1MZY4Ah1EfO1FSS0awXmsWAkxqMLY37
1xumJgt+7xGNsD0akPoEQYd3BKB9bnZV6606Ji4GWhgBWaBQr5BstbG7vp6fs4zd
+yCia+l5+ShrA8wiXyUzgBQ1r2ole6EsFPNNt6JT5weWzYNQVL0YT8Rw6yZvvrYg
NJEqzeejbdfbfJeEuLnZYiw3N+eXXtQ43Yuw2cEUa4tI2PJa0gk95cunYN6yfkd6
k//OezGMZDC7nolxwRJW/K1C1rz8UFvU08+RIRQj7+FFY3mmxi650WFjucQ6kjDT
BtPz5QKYnUne3/k2MRHRq+uDUqRIVrYsgP4mKMwPcxnqYogNpBr6g4QYhNFVVbT0
gl4AMuQZI88l5plQXxwVpI1Oc1n0Zus020RLLI3+aV25dxAMCpIBmXId/Rr5/8jW
CcEo7ao0C+/3CmmWZ0MrOjimg6owadMrP61c5tk63GUkaTUfWqnDDC2Mt1nHBsCU
xLcvGsoEJ5CUAu00fiFUJr8x0iddK7zeSehx7M+ynukIO/017y/AqMHmj/sgF1vr
YOBC1Fr+oLLvjICinrsaFrah8zqINgw1aaPLn1acF+Fxm1pxLDrmGkiNVInfN0tN
BGuJWsYXCTKmDzX10E+je2/5y3TaM6JjtMyg0ZGINmLR2UdWn/z7otnu3S1JqrqL
N7XLI8ZwjXiEDeppZ/QA5oiX5un/D7ebsK5NXRWSdpUMLsyNcR/SVfWbqUaiz3M7
fWCgEiMZbf+dlHkGYw2+GPEG9/CFR/joH1GHFYpgczaFRTc2KSEhuTh3+yuD29R0
7Pt1aqEV6RrfjbcbqoGtydAfe9NyNDTlbUpuzxUi8xkmaDewP1s/utIf8527GBAy
bhUdZ8TSlPqfTp20BFrIiaN/NXn6SXWxdKoxh8FMDqPoDoaFpmu/dO3vZuqqRDV+
0+j8OQ/gvzpA1BdT/ePx1mUu/I6qDu9JUnQWzMkV+lWfuo2G1B2V8l/dc7IMeIzj
yJ75nuJ4ue1jHJSanweQ+8Td10kiJh4Nb0DHw2FHbwsubbT1T9P++LT0todiRf/9
ALym3Z+nW3OOAbZ2V+gO0PGZr/hLxH4uYKo7y0Kl2WmIyIySgzafOC+KhKfExOCa
8SpXdjiaNN6y1z5hye97GmZrMyYAyB2wIfGQ6n+ZRcgzXcleVm3EodkBO7SZa93p
ke5M0RX6yLKTgmACnxoXpH65tPnLZyc48R4sqtIory+UDn9p5L4L1Rf/U4O6WXwz
Uef6UGjjT+ftwGLXJZqWakzLPUbm1F2TEUeq3n9p+s+PPu6jW6uFKU2+q8Pv3AVb
Lza43/P1p5m0OmWXv39HOrEoF9jsVo/MlvXbQ2AIlWm68SJCwyveogiTLruDGDp+
wJ0qocUq8aXSMGEsAhFLzbVo8NqPrXtOxCKgrcKEev+z54p8gsIcrtTUpRiwt8jb
+oHIRTWBGV1tYVtFyGLBpWPiMw+ChSl4wQeId8mi/5wK+j6X8TZdSBYlTVHFpgwu
IsQsaLPBA7aWlK/FwRfGxIDTewlm7hR5XZ5z74X3G0Lyp0METr14eKbmeRJMqFkB
0QXtwbypgXUhIVjFDChp0ATTnEQ0PVmnyKgif/TUuFRhk+cHJbVOnyhHp2FT/G+U
v8GQOJ2CxrMpb5xl4/2WFvpKXHdjkrenyWSigMZw0d7WVorhj2Xxv7g3CCsrZ7cp
mD0FpBPpt9Lz2SPdVl5uk1zzERaaAgwVibo5UDWL4kYc7/tOJ2Lmj8HY/fiPDD4v
SMrAureoUhWfqFvuqLHJTpfiswmUvQ1j94QISyhV8oFGnOw7kYEyLqMrUhmIu9qM
UwBaa/WKZQCcqgGOa7nh6u9ScOKwcLg8ANvvo/tQN5zGSrjDiJ3f+g2en4JCmRR2
JEM98GTZ7vlTmp78S5OAckthtLMaWQhRIWgKbvIi5yUdGtpLVNmVNsfTKhcd2JYU
qCNYlVXKdpgTVarMiUZKuFITBMtG7cMlg4OnK9g+99LvTOiARtCDrSx5+n0H+4Oh
hiUHHVqOERYgAQVpX7ql1t7zcddwxwe3/6Trq6zgFwhYLrbvQ/tvwX519z9TE+il
ZObyMUPZIkDJ5T903UMz81Ej+Vbc29fYZjcsK1iZopvR/hP6SPMNv1SkHTxnsNkU
50G6szO4PSN4k/0dIV0PY0ff3nM5CrJLC3ScUFOBZ3Q05iiQCWOEItRt3uPuwROy
SJHDytWvmmwwRa9/0vBnu02p88VLG8Df0moOJzbI7krjMlqSMFfA4BwUCt5Ow0YV
pSLzHuyP2Qld1ru0FLg3YHQhoX/tKm4bN1cL9g3uP165JPJRwvaYq1D3p1uej48C
0ZMvrCPBln6cREsxFD9DCNM3fjnnxoQNQ/KYCFSjdslncH8QQCYbdqg3iwafvrED
thTWTNLv0cJO1M+zHEMR8EbKeSruKl82JSCUTOt34pohofXF/nlOy2/g1jLKEQ7D
Rp8WB6bondNh5f29lDoM0YMzrFp7CN8YR3ydbjKdpzq66SKj4fmYZhT6f2NrYUZG
LoL3IdO1g4BGFdWmGmyQQjQWSm4v/19BKsOQhDmtfskXZDWca1lsMqcK5oWgh0gm
jXeYsA8AplQ4eXVAIZdo1MO3nR1+ASZNR6cConvC0IoOkHqGBYaY2o2cBfA8ivUl
Bh26tR4zVn0gFwCUJiH431dFHemutpmEF/DBctU5I43XVCvesSeppgMGX92/yuyj
zCdK1QusaJPRXxoCA2Aw3FcGd7vrlY2HR0QfFwhAeHXac6vaYxhOo7Tu9AE34+56
Zi3edsTYmE7EksfBox0hp/HwQIKnDhwSs8AQ41eulVAbeoIgSWE+WajHswQb1RIf
FMFxKUlAGO5mERbCslewAvo71KuvzkfemXAZddCAURUOWHZ+Itbk/uNhNcYIPdpd
rMkTj6P/jcbIvAC9Dg8mEQ9dUFJoM4luNjEBVdPXp6Yj+wWFH2hYXiSYXGYEqavm
SbNiOboWNJkxTCqOlTHRbX954tMxjgjtzgCN2iSawIbJaWfiHOf9ZMLAB0m5RHla
XnA2DIcDvDk3J3k8823hXzHy5OTbhW4eOn39d96wWXa0K9xU3jHZyWg8ekpnawvN
bRWuWOVlnjzDtX1NMOTbZpZAe6PUbZM373YcYa6gEJfjGfgZX3z/bn/ruSqmGFo8
3VUG3sVxbGjPxQbrpMGinuUI9gGuovaKhuhQGxldiYuG8TaD2l+5DJuPkaF+2aTe
HbGKlkHHZLR8nodg4xFj2+R43iKno5rGbzzsK8q6gHL62VmlAA5s/BKwkjD1v4ct
Ur6RsQfovBK9JcDhb13DxWo+T2oXgzhr70eS7ao47NM3b8YBx+HO8qmNsTWIf2q8
HIZ+SI/hPfDBG6Rzb7vS2IxXpd/gcA8BJvL2X6Le9EeSJvSZg6OQQvL1uJOaQxek
J7dX0nNyaGFAJXaexy2MU3dtmsm4OjXQOOc57ZRQZik94TusEyJhyvPYbS6g8vu4
G1GRAy/3pByh37j3FAKnneitv3dfGr8Xp5L/p8DDWp6G9acNKoaQXgnV34dxiY/7
woX431ojrUyRCamODXw/+8DYXmrJZn5EvSyGnpwH5mZpMV1K68BL+MybsShAw2eq
LZ6QOEv+gGsicT4T9CAKDkMNGrMO5b49pUnmyauT6rx9BwzNUBv6Bt+yvy9rxbkM
LOSoPCQ4qSc9GK4HaFLtNjZ7VlBLbro5Mgonj89Fh6KTMHeZ4LiCGKqlN7tuArJi
+3I0z7GXGWnL9Z906AhMgGnMu39t5Jz5Dj9yrP3OK5vKEzvVxaKheT7oV5t9Fmmn
aD+CCAR9o7a2WcdgrKw4D/ZI4HBXWAbwI3T/fTTe9kwe/CCywyfC2jCjothrQKYh
AYjzE8YRUMRkhmEwl1PLH9vGdSIgAJvErFPPjmgecHwteHmbj5s3Y4gH80iQrWiC
kbO9GFI0I+RqR+rG0PO/FdwsbpBcAuAFfryCgTdRIZs16BmDAPzlEdsDMluCW8xS
owMLwFSjbUwXV3blT6EP7CtgPguKLJYy9Jd/mV20oSFwa8VR+24KL74nFZDF3dlZ
R3mSFmLKkNGdok3ZRBA4/x5/NZG+TS9BrpZuc3u4CmaU95ayc66Inq9gdFPzfL0j
7nO5HfdoukqAQXn62lxbH+a0f481DLudzW0I5jlIohMdmer7uM8fjmPOl4gt3/9u
QrOUXHpyBvCSkiJV17pBFDzY8wNCGdlGBlQQw+i0yT/kT5UgXlZmWs5nR97pWVfx
i/p8EV9oFpw8MIfqY7jZG9JWhWt558/xW5lsds7Wm+sIZd0fiHlX2kGU03u/xMSx
+fejB1g/kwkG/IWmOw2qtX8/a7bhVKhjRDwru281I/hqdZ6p1th+CLCyVO390gkZ
9j/Qi85QHMFrpu+f0PruwAFYQ4dHP8T9EjhH3UPjx3ogIZq3+KBhtp1POKSwEyXd
gBJYps5uPW47+tb0FyrAf3rNwhELvw4jC05eS0PNlsiM0jwOuramErU73Dym+wAj
bWMUtJPw5+5NjK8gQWW9DAvFuj5b8VnV9hx00DO85Y4eDrRf8AMJaU1hXxxLWySg
d8NQTXpMODV5NWjCstR9FVY+FRAc69aVQNSALF0TtMq9fneDhBsWPtOYbgek14gy
Hxj+u3LAD218c0aCkeBgpqwBQ/0/z3j3h+9WmwqRSvwqSfBBFgXJTu8QQE0j2fWs
wxPhjzYKDCvpKCldPG3H0Jnxb1vV1fFxBoOb0GhaVjPTS7/3PzKpknvnoJa/P1bA
KOoJ5ANElqD8nYLnhaWKPGqVsygW8D50pbuOw+rSwAm+GpmGdIEQlJxUX125Qocq
kpJ1P5wJ8k9PNAslyUBfHs7i8fB344wSgjhZYHDp59Ow6WKv2Ncbloqm9y+teBQb
/h9vgCrO3SWzJJ47jrt+rwxXbZqgwjUjj3xmXtHH5nO77dSpuyB8H9yBjoIG2HJK
2esoy64yJCPF7BiNGbvjZXrwonUvGRpeyuwUwEWY/u5IJXwCTekSSgNuAawfspCF
astMhG1RJmx5TRbxOHVJLsab+B3SWb+NPwBG0H6jgsYz3+rtEJNgS6IPMI6akpf8
1yHTQZUW4pMOX+l3xMJ/59aeVgIyPR3nIO7ssZWg7y6woiWFIO5CJ5hbMy44gnm8
pxMRtQqUb9nbJJN+p4tZgxnce6ph8RCOA9Zv7MhYOf3IIueRSwK9zsvoL1U87wTA
TxrcyRpZ7WothchdbgBIUBi/CUnrfTwnCE6S/601D4DWi3bP8JFzEu7lIDvoJgkT
5Sp8SWNq8i1WrsEPfrgvDT0Zn/NNZjrfbgdljNQqz4wjdms9jrmVupiKdn2BMxvg
p1QTngPlCWNY+sBhx9WXi+ylaVXqw8fJaBQa/kJMphTm3JnirRJ9U7UKEJPwIVMP
8sQpHlpMslHd4FECcYOvR1vwumBj2/hoomCs+UB8/4gKOwDFeuy9ecVYqedpK3Ha
/aXJ6toJ+LC1DDjWJrs4TdImMKB+L44YHhvsuDDDAuH7JLtmttXyHRM6sI6xh1Mv
Hd8qlPAgQ2tReV3dc4qFepRXKkC3ku5otsYED385D+vA2LN3cP+P5wnnFessJt0Q
3ZwfsVG0pC8kWBBTXCPeV9CvFhyAAKM/kcfi5O214soWGKdCGNOGJ9P3Drc1UeYi
R0u+hwi4w5wCwdwPXlK95UpcBS8QkHKjGksuHh+5XUEV/I8HQ1YKuRX2RWtO+E45
ckveOwhNV7P/Rh0WO9ijdw75fkkUTRsyvqO/gCjJCjtsFtmQAZDoJyzkxi7bx+3o
FCbw0ucrTYt4C85/scPffE1HwKgCtDMTbfCeA6vleJnmEGIHZHPIRp66/CK2lPL4
ZTahLi+ubJZDmJF1N9sCvRuCJzoduwVkrV3Z0F93ESVP3jRx5XoKx0DvcrIU8b6m
0Jl8pkMVu6C/GXgFvM7SyHmmx7SrAdXQP8E1DP8dJoSFp0L+wE4/JoI8t6FVA3Mv
jANjMVir2Rfpmqo5lS0VnU2UZawwgS/nB6fSG1ghDIgjfIBkphUnTYGozHB83gCA
/YyTkoYTVk909jwd9Da7pQEiRC0h4bx11vd/UA5h8zDREzvKUJEB8HCFl5C6S0ZG
6h1C5AEIcrbjK2mOk4vtkPmFYPtzxGy9x9K0SlTcXdOO5RgzL8SZVnmSQ43h3wCC
HJMg5ZHJN0/JYydVhaZHRYPNiCjd+/xv/C5Yu0Ky9bFp3m5XAdfyiLLuLfK/xIxR
u1GsAothTKmoxUci+ESnkHEGN0dPJq6AMCminrEsMfgLems0IIesyhpcgaDxGvc3
wOnvY6Cxua5THVjsqrjzNRXauhJB4DGhE4iPJLbW+hNG84KwcDVzjx6JBdNOJZD1
JPV1lbMPaM/R4U3+N+7XeYqKEyiYDBegr4x7M7TOBDxTtbL6UyfLEITnZkvoDZr6
vn3rU5BZdHz95RwG7GTjztH3ztjePDsOQHm3mnXHrz7Glt2nc2sc93vQEEoGWvbl
O8M41/9ZwAqLTPfHcIcEbb9wn3u7vjKaYlHMtRr9YgOhHwCrs26TuRWc/pWQjy9O
VEnP/CAdOG7l0+rtcYlcUWaBV4RJ8InI5Cfi8Np4FKjrk2YTbENrR8Z7WUMaEEoM
AvtVxTNO2t8ox43p/gMtixD2CXP+r4484LujLGjR62HHjbJhXTFbukI6IkmjJgU/
9LWf7fMMwOcbG99iMiiv+oULcYJSspFqpZ1HTuMqZvlsLxK+Ri030z5qDvmE7V9R
Y0KGCXMBUbpGcmIBsW7nG5BnC1ww4B/bRxrDYbaylOZ7uH1GohLgvu3F0ZhCGpwD
4j2MCkRiivHnGEOZfIJbeEsDow6c9mf99ohO/oqlTf2/p8KIPFI4emD2ALts7rdk
/bfCLerfPaJayChGw8mQkcbsADexKao+9wBiC12BnrFgcFDYrlb4Ew6e8/lUlWmu
6oSEITpYZB/Jz6a7Y1TsWsw5JlKEWJUTKpik07C9T2hIUzJY6yQQUwtpAKnB3zkh
RcwlYziUhJbTvHL3B9l6tmfcwzFPKYvi6/c4s6JHhS3Ek0hnkSAV7j8U/URl4Wzf
IS2HAtKvb4gbtsgxcdV1rXHk7sbSOhwXrUhHS0/ID+zFAtb4NwsypHkehIfMtVlr
VrsmmVBkHtYBK5CH3udFRc7vf42C5XZZ5A8jCs/HnAzPNqPG+7yQ1XMMGYqCcFai
Ik4z9xuJ+VbnFLntLtPcJ1WW4VkY+3n7bZp0XKUKkALxGNnW5oGSMVXcv1FJkYJn
ls/uDmqK6wV8JH+3N0j93dJGtds909WDjcl5qJtjO4kX1AqN7fOuKwHvqINHSQ2o
GstV2KcLO661b3873n6qMdzTME9AM2itxjkhCq8/baW5QsblpLLbwVWV8cQuSWyj
h7Ru/VZjfgQLSX7f1EPkPXrxWx1mrn9RzR+g5h3iX9Mbvt0mT/Ta+84z26ncw8Ai
ev4CFyrs04gI2x23oWGXQ6HyAKSnZ/4Y+4anu4wSdLHuVaY2vIjAhK3062TQpMWb
hLfFEfbO5DOBAgHPaxL7ozGoR0VTqdqxwBr75e2EkBHGMk+gvsctSYcsUv1VdNyd
IKJb4NdK/nij8zwW7qtWvHHTqWjojFGRZV/5sjuRqh/1nhsreXDkSw4lPNGpCJhn
a98ZrwvIcIW/0KXHiW0DYfW5LSH5sUZzcELWoaUecngTBQLkh4akY6IxLY87iipG
KUbeqh8AKSuohm0WAKP8UbfNVHRKeI1lwDLv5hKff4APsgj4KXVZejufg3nnIeCH
IdMO6Lzqsv2YI9j0/37ew0bBed42vqTuGG91kh03ljyTrCax75Pi5I9c9LOcK66n
XdMw0/a8QgYgLjTHwfatGtw+nnQBHSDf6bPqlODLpTQQBKUDJJF0F4IxdW2rEQ/H
goFL0W8KANYINZWDKAgAtamRUNzi5IzLVfoHLYSAZlwjwHtNI7vhrreldh+b1zWv
iMqF04DddefyLiSbbUljOqbDOixXeosHYJq+0JHUcEfqrFJanHRVBssXqxDL3QW7
rZroMybBMUOyai60Y1uxPx/qrWsYPW1gQCGStdwWxYtKuUdLGQISwxncSGEqnTgo
9z2xYh+x96O/UM2N2d3nIu7B4rvzk2hDspjuOfileK2e4E1U84xgpgI8PS2DweyX
bp6vml8PfciRhGJc/JpAOSxjEIOAPT2cEs1gr/RtjynBsJeo0Nu9IVnoHGIhEG9D
+y1JbnKqcSMrYOboeXUZD+Dkl0ILCCsARQaD5lBd/C2rQQVcleZ3/CV4Oiv9pD/c
exFe66AMysi2shLMV2HbX3mr+HMJN3D8zvwEgyrOx4ht5WtSDaU3dwBhZLksJqSy
mY1TEbgk1R3lGQxiUOrhoGcd/AYl0unZ79LCTjWov+TuKpEKde8dJRmu5RqPpVEt
e9ZKC9WGXvBWci8rX7511GAtWPcjdBRfZerwy4Z9KUDe5OdTbiM9KoTzxQfjGkuG
CL3ShiwweQ/iuOK4fss0w0WuD0cXYmFwkDqB6Vsae5PWZ2Xr480EPtlNKUS+LD6o
Teg4L+dbGn2xpCYHIKC6bmE/kjay1OXI1ia6AKP0cODsTgCqmf7KZDOV/l1L9YrJ
Z+R8suvoDcR4nkomCDYXKjyEHlSQxzSOh+4v8ZK6ajCO+Uih3uqTDj2wmcu6adYw
G4C5/omOq8DT7Gf12N/ndw219t4rN5jl8NP4q6Ql5vSJCBSt/emj5tvQIplEXGYf
pBwlmT9YdX3DuXwZ0rHbyKJwg189uc1Pi2rllsd1TdyKXPQ+rbu0/iWMJodHd0Rf
LK0IOjgCpdLS8rH7oUGINChsQxlntNJvnhL/IF2VJA3jPmcJz11yCkUN4fkdm/Zb
lp4ZATwPuSrWpTJnopb/NFrJYBt04c3MQhQZbsa3ibJBa12HgMUApYNO171NFnXz
v6x6oN81YWXvMYpztMLRhEL7FRxT/FNE0Bgxft1zB09+FmGdeAg1cWG+Di1ol0VN
g/JWu6Mf71gNcj2PgTkquEnbLjn+9unsScUa563FytNSj1/vnabl89UtQjRwOlE5
XEND13lnjHEMZYsyPLUj/ECU4DZSftWvxPuSkvpvVgW23dLoinZCNzzOdh58DZ/F
jAk3Vsl3QKgzA0k/mFdnM72+QgED7AcNBb+YC5XpIAFYJwcxG7e6j67ZNTFMfLew
+yq/S0TpCaGROguF3YpxF1qX7VmQRno++ZEBGxu7lz3sI/SOWVIHTLar236kFJcm
tfpkQCaCKg7HGMFFzWvIaDMiO77q7LrlVbLgMn6PMtrRchc1R+hIMiWVuQ+Qdprm
0h1370J+o+kMcmeh3ZUQj43ky3Ce2MkoSL2Iipvp15jHkFvdb0kS6tT+XUjzlTgF
CEMBdAUD0YF3bHKePfL2FrnTLKUH1tY3WXvV51jIGz5gAd/gzZPtPHLXmNcZy7VA
LvkAPoxEBChmN8JpEXOLEUzD8R+GdK+M5FjFSA4KkMoPfpTeS1e3l9yuDn0kfZ0Q
yDCmMIyupGSAOm0arOIrR4GRYusHmDJUseR2P1acYlOWwGXFc7MwOnVymNLg5083
QFzVMJ4+xkvySlHVX2xGSPDwv5vYGSPuhiAi+eoRqYqJGV7/58NPmrw5G83mrzZV
jvhOHL168kl2u9Y3jHdd0JO8EnCEqXFJ4X6xnK+K4A/7xRrqH+8b5oS+k58LcabK
HYubf6MFkS3qTjc9Xj+FTtGJuJhc1BG3DiTbaCDbwtIXuzTpxbzCioeVINP0Qi2U
nN44z85xiUkkdRyZ8c3qVgGZqLuKe+XefK6mDX6zFCrbdaq6in4JdvH7a+bwrCGf
vki/c2QE6l1AeSjgfNeYlfC4Z7m9Yent6oQs1VXnAjY1GmQyB6uucd8WjlV2BBKN
lIaEYA8KH6z9gyebW202xt/Imeepzxi3UlAnpyHJGqTd095djZVSTynxyt1cAXJs
cGHRm+fVBP1lwdyrnwm3hRVuPDdSCFa0DWwXzdC2vp3bmvtMOlY4heqfkXlmtkpD
AuOq5Uv0AWCAFJOMeSNKMl7CBjTDnku2GQ1oRZpmPud0SIWjzvybkDIYjSLUQNhS
Y0S79v7z8ZttXg3k2tplslWW8S9F29oIdPGLCA3OqByGviR9l9X6WQt6WxFyb3Bf
r/rO7a5zJANKBj7ZcQpKMrhFn/ObEUnEYJ6rUWxN0DX2z/MCeo3AC9H3kr4ldDcN
sR+8K1j2+gfzpbgKv2E+PYly5bYBImrz1hGTiO3SChCa63WKXjRpahxkNEr1ovgM
DhXrik61UpdYrhFVhsnn4B35swCmmFSZPYdRwGfKhYOEZdo+ZlQL6y8SUQEOC5ZG
CBi5xeapOxCbcpG2k0pihgE+pZ2VHJLGjY4tBPv8z1Gtsmn0IjwXaqcPwzEitfef
ObdcSB0wESDgqPQjnXW3//lkPGB+DOW7BwU2AaD5u5POPw3qbmGKzLC3fEasLJv/
HUO6DK+A8UmqsAj7w/rP9MtnpvcmwSA1sqLHb4Abz7BdgX8JEYwMZ5vCSPiwuZV4
dv55YIsel096VxzthKwRglvFW7/7TKNAInahbRSZKaTpi/caJdAvoTDdGrag/q8u
ezSCdXvZFiLi961q0BQK6zXiu5hBwkz/pHfXAbuLNmolZQjG5FPiRdawEobJBMc3
njqb+V1pkpN5/7OMsKG9gADoo+90tUDr5wMEtJwC3vEWMEx2Aj9FzqzWckRoLQGs
it1vTf7Dlho9BBBUdYsJk7G106WbaXb86y7HdDLm5YrLO8RAFvZRUppv+RrmChRC
z7T1sOUefm9vMaBdvtKHTytTDPhSHdp+GmSzjD//7SmUOOoTrE75EOzNxUllNfgz
2RvPiD7tPtI/D80C8lP17AtuZzAO0xGCy6Ip+DTusans0TJNDbnhYH7UFe32jqdt
ud6wC3TZBKXCIoPVppKtp2447/WaSgRIOp1tvEaBxs0K/VrmO4jScBkWDo/1g+/6
LvDl2Cs8i8icU9ZyY8jmDhKP05idvqA7p/Fr2AExeA6OSxCbFosAwGEmoG4kcuWn
IU0LuFdwcWABPfn0/VcWaOdAB34c3OLCw+4l8Y/pyJe0okWh0ywmwMVibyofUEpL
gKP3HjyxgBxiUU6vEusoetzU2BBGG+OkrclnMyPVA5WjZVUHzsyzh7tN6nUJJ0ny
ZW+sCIjiRPGG2+ryMs/DCVybneg/r8YBTU+P/lbzwYdmCq/51pLCD5Kgmm3XJuYF
qZHKKyyTcQjfqbPZu0tTXxV9lxhXVZmO/Y7ssTxiOeVqcxM+U5TLSLCv4S65E0nE
2oQkUiht5NIjoRf5G/3Yi9NpwySCBrnhpI39OY8wg/omzXfY7OaLoy2SB6yFX01D
gH33ozeQBaicEgxTAPc14GB43EfsfGoG7tuDJSCKiifGzBCzg73QYPrYXvCeB/Kx
VR9RT7OtFjUkDgl82ATpRoIZCK5u0aO58zKu6oFCFtwdwAaNKJAm8drp+AVpZnSK
ADr8ILyBIjSHq4ZTT1Lx3xfkM2HZzGnomp3F9EbjLWpdpfxzAxiDxEsGYiX3OCz9
05aZAfOi40SPH6F95SWOvWue6E4fWAhzQL6jntthXeV+vysE+V8eq7Ajm1E3IhhN
/VkaIKI7kpUY2rBIyV2eHzrmBN5RQXnuAN7v5mMOd2pGgGGbr6vTLL7Ng7nD2TIX
L0biiF8luUoUW4aiJnSoQpH5TB3/jdbgyLwRA18my0MHJMah7bQcf/c7J66ikAEM
Gj1PwjsTU50BEfuIV7mU7DyCG3J8ApggLovJQJ10YKu/FGmjOjHXLez1Gqh7jE+u
zgvkPmnNnpOrdrrqiJxf5XLQJy6W1iKfNMDy1EXLEDGM1ybxoQEWqIhodgKHrKoN
sT2pYgejV7HLziHtpJ7YTmHvOrv1POLm8N2zp46mG8+y1Cs43gR2owDE8vmZ3z0I
X2wiKjeckiXTq2ZKTih+0dHip5X9wX1MKmJ/NXIAaETL2LIW4MN6Xg5TZwocWF0f
1PPjOvAWsv4f2SYqFgK7qmD0bIacnkqRB/q1Maolg2VyOCSxrwG93R0ueJ6kuWOl
u6bpzZcIaTcFYWP0siU2POV0SG/N/xgJ3QCb7sCc+jZaaWjtX3dYwZ3onvUALD4o
p7sCBFzjqTM9EhY2UILjYzLp+ym2LKRkzEy8SsmyyznSAf0LEaMK2ycjkCA1Rl0l
0KRumfm9buTDnjeOcmHRZvW4NF3DSTAT88ZhLVhN04ILM6UwgaMkDw8lytnjEov2
50r7Am5MQmH6vRSJp0kkWuE3znXJGf/Nf7/2rssfsFhboamUH44sq15UlKtkot3f
uT+8zk8oio3/IQT2pYroa0BQCsMn3F65V/+wYlF2z+9nrs3L53WSk+FiQp5SexBy
gPcR6JO8HNxM1ZxY1grmVx6zX7LlBVsJ5AFpaLB2qvxRnhBcsrdeOdyQI0n5BJyD
cdmATfpKOliLWvblbiaye8WNQ+ijWDRdfSbw4DQDAd71nP4lYyBYiZyNchtfQrU/
Pyj1lTRx6xAn/qb4DD90tGDhquMQzZ6GMRC8QfarsTJ6YAIqcqZ5frDH9+B5Bsu0
sSZvr3OCmBsACJ1Lf5QhmrJuIFDySDeF0JT3mp/3wFrKoyHkhcozNk5TuT0tKvCF
uVwAIrW50waF49fQfbRYjuxJu6mA/o8K84pBGuOng/kO4oRTXyFq80GA9Inf9GzU
/w2if5KMGPdIjcsQwGut2X9UoAC33YTOWPiBbU67aw6t1dzNfv/w6NnjzO/q/kKl
g+RwlrKYCOCdjGGs0THQbABN83FCvRS/YXFF9+KzlG4i1MN3FaK2SIR/orjPahUP
aeRKnBT0ydJGO8f+f3HgeKKaG7RaOuJe5SFPAUIu7xL8mkVQSgw52qxsRDCFppWG
0+W7DvCvHX6Oy0syYOGQlgNM0vo5hj1nJLWKQriUXZawJIabkdH7LYjYBnbUWf4I
UMXUiOYTbMaKve0hPnA8LqVvL/C7UQJ2wVpgopD0S9104+MOduq+4LcGcC8aQqdk
u34umjQ7N2F9Rh84nooLHGAYojLw3lnHOaNnVhw9GhTJSkhdREjnAkcEhyFav4Ly
7e+FL7DkTeb1jx13M8Trc+24lzWT2sYSol/n0MmwxokijKQA1vPjzwUMlccZT4NF
TupjiulDUBtkTgThBKvkBjMxsfl1psQj7PUnFeJBKj7A5RDnmC5nljg2BgLOSBfF
MIvh1sKpp35fiw0HMCZt4EIpEWvZmmF6BKVnwpP21YBpEf9HBAHcPM0Nl46FhAgm
kpImLk5LBA8boOoEOEhhJXFU+g1b6XCo1AfiZWtAyp9LL1yq0ijlaK0SnR+YXuVy
K2jeWpk7fTUWjptBGxqmAtmZhh0ewBe+olLEdiH4hqkiCpCzbK+2Gy24CevYCGjg
Cl+0hElapvt0PattcOPgNJzxATKLyymczCb9HmvEosecqGjNk8cfJYQkLknhMAHg
cM0161QDtUwnEKkHJ/DdjbbfJy0SeXF0HBr9fVDxxTSn6GmBLCUXCMbhSg9h5pva
1DM9Z88T9AbxPXaaiwEUO54atiRzRJQjIaTCA9lRxsO89sC+U1u4rpDeWyOWBfGP
sQZoCzQwghqbEAWUl0qoP14XakTkblfx8ejg/HI76RGBW+50hi+lFYVZchLn7+6+
z86sDQKcNqyaKc53EQMJlZ4Fwn3IdKI1bgMMb+p6Hid2SAbe2jINdRyfX+lZQLt1
1l3rL+w4/rrX8M+Wf7LslFotFv+94noW8dyzb3+rdR0/wAQj4nL4U8LMtUrbkLS9
2puC+i58WSaYgOyoPv8T5n0xhQl2vODaVNucrB8M4v/UDPuua13RBDH2PRiA4B19
r8xFgDWc4uPS4BtspgYQHLmHXX165ZnIgDpInrHRNgcb+mmTiEbMA9qGQEz0FvmA
E6gD003SOtM6uzQkpsJ6bmAxVPGO/SB0YeQgUusjkQdPCnBaw2BNUndH0zaFTUiz
pgmooP7kXR0Pt3QMC3oNNACVJmRLTX7m++xYpzCRugUASo+8QaO1VMT04gdorqVA
DxJpMTRPIWAk18G3iCNeX6e+HhWaQB1JTnhRd/glsBr2TR0gu+McSM+9N2svK3QX
FGTPNwgW72La9FMLmniOsHjzXaoGm6K9tPlKtcHfkOdGIHtdW8suAaa5wPqqcO2n
R95Y14lAe5nqUT0E3WXmARSUefWrDIDE8nza1Fb9sKJddpRn6TFU6IDys2WNYe5Q
acPpCUgxjhsV70tY+g42IswMcaydvqlFtMshrafD0zsAbVIxE4ZOMH4OManL0eDT
Vei84/3l4pSMkzpP7/WlD1HWlvxun5BianPZfU6DOuT7NNSDnlVvK48wvePoR0Tn
ymG1kIuy0v+Rq6DZvNIhM/g8QZU2/fZAnwCyW5LBcNi/VZsT6z5OwBHXif0BEmaC
ffxm3rcPEiBeSh0RhaPe6xsxFepvTOwmA8ced/O0YhxzYgs2fw4OgT9lL3cvD4Lh
LuKQoAJjadgL8aNUmg+jTkKdH+yG7FhPrePxxyB5W0Tai0zWM62ZHEqgvgqY/9xt
7dZ+WWIfqVAUSdUt2Py8DR2+Snw0WgWBOdUlAzyaV44hoBgIputX4CPlXaYxAMBC
Ag2TKqs5EK4MumNzm5VQ6hDXdnMwkrGOly9MVVA2qCS007M5AZ1D7nWpyMFHLBud
u7aZmN8Q08LWOoX6GIeZcdPjBYNnuq7UVeAdTyt/F/LoRiUnsr67JcAVXXUhzbim
KPQoRoaIKUcLcSNHn4l63CSgL2hqwnXAvB5YtVYxdSMW6J4FsjNF+w5K1pn9x0Bl
QEXUQHuBWKaE/5hey178Nzn3nRhELv4r/r4J7jU5+aYZA5AKeLL+hYSemIr8B3/0
at53xml87r3d+Jho5D1X0WRqZcVr4KPDxgyuY4u+7Q3fAQhJOt5h3P+rsafMVTnv
fqVKhSKAKIcRDyOUgHyOk1iHhjbGFg7QBbQTJRE6jwQbSzKsJhvHJAIqUQiOOJH3
sRzhg/xA8+gjhzpdFMWBu+C+CF7tdWdDGYL3BNP7CaTUurLVUncnBb32LycZFV1y
LjlDgJMJhJ9fT7puM3TEm2EHmMt23BU8bR+wPTq+Z4a2BTKCAp4E8NY03ANJZlMm
TDQzgRh1R7e3E4liUZxZAdzu146GMD2vF4QAe6vsOWO/RhIWGQPR8s/3u9pwyvCd
sG+2ox7r4f4MK8JHruvJH3nACUBl7kiGyLsF7aP2af50RfVzdjaGy0zSxGpwMZbY
9/wthblGJnregEZjHbxu3SQ7tcU1Je65C1Kafs4QaqIzAimc7OZeJ/ngRKH7vWay
NzQCSpJWfx5NdyHBf/UUIJW6ucgciQ3u5TYdkNhS6owobcxkiusJL4IEkp2muYbl
tDZTynNzLlp/Eqfs5MebCfvmJxbdLTQSwYGgZbHmiQC17FhhqG3aydN+NVAFpObg
cfHV8uCxPEaAhgYwgT+ZTaMfuLEygujOEMRUI24NgYMnBggMD3Tbi2Bd2YogApKw
ZWZjfOQs8lt6jIwWHBh23V5I+nXZe+7zYbhnbdzA3hThQkroLdBDKnaecZeJd5Xr
3OQ+ezGMHMMwsz/nlmO81go1I2SnGto0NpsPHrLqVQTwdv0My/PVHxUe4unfD/t0
0f29UdQYbEz9yTfrh9o5W7Z/crkx3Sb4zjNFVYqLLnxFY66I3pWWuM0abrifa1pE
U6AJBltPZSSayGuOo2NjPkulrpBTLxbasSyOAiXMscK373PvMQGVUCtINHTD6f2x
Wvzs64smqmW16yzMoQQ/DBLuiKwaI3ECoIkfb9yu+/23InbvOG2chVWmTTNyRrcw
kTZmpGitOSshdNDUYULmZOEYiG3Xrz6vVZ74yPwuIJdRDsvoMS8i2WYCKCxURIxt
t3Q9Kn8kc/S3C0oBo9zUbY/leliaAF3nFsREavA39VitrFY6EKYXFlz7UV3lGy+L
dVONtT53kI8vT/YoWHRTt9SID+ltCFLuFsXU4I4FDHyTTknMBkQdTNsnaVQRfniI
vpAqmW6L1PeYXfn6OwAaHURaKJTmm4JwZM7pgVrXLkUI0BOslZt6DFmDpasAJusY
6/WDbwOl6Shma3m6Y2yLEKuV/5KrdXBqqNXRZah9TR+/BfaE1X7bXBam3oka3BGt
htpernoEABWMopoBSVruJe4H5eYehcGBrccD5C6owDQTLRsMDKhepx/1xm2KKfwP
C+bZwVxtjPP/+bb1oyOa0fDoe4pVF4qa3WXMqIeVJajAHFLSAOOvMi1lth9KREaD
5MStOgVSbeYuM29ExBRhC+0lqIwzsiijgc5bKFqm400sjDmkGmzRnPsg5yxd8NM8
aJUjrxq+j9WvS+pTLEQgMrWzQS6w4F9qztw9tr1/cvSeMi4uYLx3KuaNE06Xzf03
4fItqgA0b7sad9zU7GPk3JZDjzXXoweRpcKyf42Gvtw2qs4sf3f3IQgeoco2W0SX
0tXdUfxfJwyClJ0TpJPngHuBU8MvAHvLyZTXotYQDfQJBdYEeZRyRDO78TNfWD1O
liiI61eC4vQndP0fngXB7JB0RoGq7Ply1O/BoxKjiTFr1hkM4ckNmHaUBYVv7W6V
2MU7+VhEDH0S5t+hLCOvzqWj4zuJJS0yS0j4aoavQaBsgKxXWBfJMn+Ko0+9/Q1E
bJZYwt110t4DOqEcuONrhbEoJE3DJFxh/9zUQIczjCK4WDGZVfb1g2ynibgWqCgK
63v2yBPU0wYMLPcO2r5khKZiRZkAFMNMpitC0vxYYiFy+Re8diiIL9E5CODTENUM
kLEGGfM/OAEkwiFJ5SLA1hboetiAloem5ni+CVyZVa5aL2ZATtyV/FjDq6lOKvwR
cEVBEWAR2NAcVSPyNMY/curVAZSX9fDVGREf6Rc0wC5a0iSevAHO3zipZp2sMYa5
2K93xk62DGf6q6b7Po0cdCXfzf3jaBfj1BV3VKLWj142UBkvobuI0zOew8fJUyFx
S8G8jFyXN0RU995Ag//VDkD+TqF849FTYpe0jd8qKUrMpKhgH4hs9BE0N6w9sF9h
78GNa/J3P/aK11NL0uQzwuWEig505ocEWtmaVvir1zaAZIAFL+DAkT6YOZxZ7bnQ
No6X9734aCFvyQM1+JxiYwUQfY5fJ7nzU6gevWvT6Yk9y7+RfDkrcEeZMigMQ0CB
AD6a5lJZvfKMpL8/qv0x4qHdN9LLspgKKkfoa7rFcybmOIx6RHLo4thhRO4T3tMp
tgLW0n59ZRKWOFt3CVK2R1AwF18xzhPWapw1QvKZFMBrRz3EE3JCzzCKoWOHiqNy
pxuhZIbouCBXD98UeuJ/ogPqwIrFQ4Hz0IBm0wsWp/fdeJLtiWjn4+xH6oihMkDk
jXs3EzGh20zwJfc4x0CSHw3ZAAHcgqe89A5whX5D0oC3o+LG5M2rSuU+kOme+EA7
aIoFD7ddwqw+nZrTPBn7pYZhPlZJN+jty9hwg3gdSfavn20HQrJELsM42elzD2kN
9Oa2cS0trYbkVdfHGGdgGS3hUjTgKUK1KTjVnC0wOjYSQmvrT0xbQzdZXS7gY2Uz
fEY7SNcbQmU4rFnrkKfKxtEhLaT0R0Ag2KOBWowZBneOdhRgZHls4nODZFN+B9On
YeQcvD60DxBKhP39b41+ypkBpWsM7e9Jxo+6xxUpoaVmB5sX6CvAzKnZeC6rAA6t
PVbXUtDo6E9k4DCcnPMne07FVoNMRVcLxXtm8bG5mVUv8ljOuwVtPkS25hR6vF7J
OGN06x+u/6QKTZXpK1B6vYqx5h1HWWESU+csSek7HOlHRBJ8s9/y7Go1vcPqMvjL
sywRK+J/H+B9EwbUZ5CUhUdAKjGLG5f1PjlhvmK6JfxV/ouJ2KZ5EIXIKlfgACUu
/uHYTsVXlrf/aJ7gV8BILMH/3LDS8P39m/eDeomVQnwxCfULijGWzRYaV1fa//cs
DlyCtHdZwCfAiHyZTz9wllHHSL8Bg25QqP6cjgfJlDwv9/v4c7a0h6fAoh5OYbFd
rn85cYz2Y39TACLLfr5zG5n1aViaIdNcL+tRxHHNXVwS1bIcnQi/U6F1KXLGg/St
PVtmCVtVL16kg53C0F3j11nHdx2XbGs4g2tPIwmnce9vsTI+ys4dOJ2ulHOGUM4M
fqtyGdS64T4hrdquH9BpqL+MmeWpJAQGXCzoijMy+vZSQ1zJfMa8x8aCA+2pwG+f
WMCZBPI0Lvw0hDI6C6YbbBzFypNWWeH/ABb5Iy3s3i9fauxFeLOlWX78yaInzcef
4O790XyBcMupgfZLEcqoWvRxhruJWiaV4nUKW5J5HWuO+NwwURqeeop43g40MW9j
VcluLEBsPyHHV1IJp377ZQAaI5PG1JD2wSSTkqQaqGrmWN9LdvDxr2iYgJjlZy9R
q2Ky7hUk1G7YEgW6Fo4RPIsfzg8DcrP9dkrR3rdQee1Lhf6F3QwJtCpLl9UYy970
8pr6ZE8AMMK+SWofUxWvXa+fD9DKUmbXgmMuzXVqaeP6SxgifSAZrq4uqNH38j1M
b/D6D9mXNPCqG84MHQidpSSAEQhbKF4OQSdZCUBGsnZYSSL15NIUApLRPRHpZLhv
Pmga2PrB66VizeTK+TL2CC6mAfgI5dt0m+4+Z0WcCvxxUjUFG6fao8H0dfaV7B9a
nxklKMFzmJdV2qcyl5ne84tFTEsR8kkMPBJM888bu5LKFWwSoOqhMEUz7I2cTrxi
uluGwj9iyL7sKSVm410i+rLb9uWgiXBr5hB4dlLQE0KZlwySCk/rk7zYOpguAwzj
cWBLu6hCuh+LwIVn6KTCgw1tFWopwXduYHO5M9gNeIv4xkcoLt9jKhrf360TGX65
SIs1qOqF/1P61ZYyKqLGXnY6g36kD+BE1Y07y4Jfnn2Om9Z16PyU+r71iyvKe51y
zEfuYYQSay32k3jAMQVGYPpEsZJ0rH/7gi3N1WepFZ/u6F5B7GwhzrJ8GL0wQzcC
sRJ50FePgfHIrWBdodHUTKe1oOIYULjhHsVuo9GzKFCPXKXuHxCK2hlw4URD91zO
u8LrUS6XGRl5U/u09XwOBK0JPzsRLs/Ig6+1NnfyuvXzf5WMWspQ25wE+ECENJEB
WUQHD4d1SN/M2N6gg1bRpM92U8PYmgfKv9Nc1XpXyQMyNIGlQLQDNkPezjh+sT0I
iW0LW/EH6sbkZEeIrCfIU61H7hM2Z+LXZ7JBGTZG7yyvM6W4M5cK8nDFWjavSwgd
vHS3aJ0cLM4fZ0JoidWNadGsXGLLKFk4vqLygK/FF/GTuF128YH3sqXFLuvJWih1
9VWYWK6aqyWUDWNP1DItSmyz6f8psb8iL20BGE53wzhKJktL/hPwhfknvXEoyLUO
+o0KDcHbLGtLskC68syUzvyR0U4Gb20akWPVJBLyZH8YNLOmDcjqt5oSzTz/iWom
SeWi+eOV25RCcBI1c943wA0m5VsrbetrdlXEGvLuAC/4Vl94o90hOdaVHUcpwHBO
fi25oqu+cHLZuKMCP/jRlKKVpKkmyeXe6nkcTbwROV1FK8SMNijczuO/DXgvRfqJ
ZjJpf5F+j8p4zKicv4l812fUgCEA4Tj1hgWLT7doO+X6iSRnZKzWdJnRhvnOUTrQ
xBP5f0LwIpDbs4FZW1lCn5vTBqPfbcJPRO2Tid5ph8K9e3mPhGdj1SeCFzimtQYo
LEeIjK3Q8vIxEw4/gpk6gnNjETjqkVC2Wurr0mJow685g2W7SjIkjhtJ8eL5luq9
q14DsR/7Orz+ECr04wRO7UysRWbU5T2Hhpkr4ndmyKei+1mtQJqtS6QwmiIBTCwc
6yncGbrFlXYgxvIqrmu+LZriPZ61JGKasrWAg6S2sn5ALs9XzdeuY2y4Gcpqb7lo
O0PoNlL2xAYs2MMGjb21HUdRuARn479Na3dHLj09Ah3/ZvrIWiUEiY2ixYkKEPVA
1knIli1+wtQ99IFRLNeYxCRvxj1aSUKUn8t8lK8dRgtRFwV6sMndMmsEiqJXF8xs
86SFru3d78eijk2EAm0/Bk1wIGPSYM2clUt+CXcVN0jlC1xql7aYQjIygUwIUWQr
9oe4rL+xWWfkXORmwAWZydVkzpbiwRMNgsXwzBpt0w3fuTv8FRewf55lpOc6Vhk1
3aN+sVobuGjr69R1Ram2mIcSd7iJAybjOE1lmwqmq0+2LAAl0ySPCaRH28WhLeV7
OK0+bKoHyzaaP6/cwzaBJ344xNgR5vlP6cuL/CmJKgofZ6rZ7JqdYSHisKnQjEN9
mgzHmMKWIaQdFi7Q6zr6StMfM5Ai2NhjtH/x7VUdp5zmCx6RvHLGJr+Pa0FQsyx5
ogR1hyruvYOeViOKPMrDFpCR2oGwY1h9/N65j03LtP0Y9Oo722hkwhNYOGWvsn65
mwse1U3DuAvxbavIxECS37hoDBLd3BHmEhc5WCHlt34y8GuRJR9DRSxa2cmlAJo9
j+DzJxQ+hRCYJrOhZUzjReN5cSJYnKuxwqGQDm6tys9neCqhyDB3PkKl8ALMIgfp
vzjtsEcKkpduNXd9dDIKu0jf/1CsQZBVXPbB5ygFZlen1SYRjQ7fbK8lNfawidiB
neaxgy3X0RVG767a2i0L6gq5GAzFk9yfVb6eGEd8gjHQGMHoQ4rwN4BlICJ5M0r2
+BtJOQnAhxAKGxEc1Ll3vhDxOowAMb2m0SKvKcQeXp+qwgUM0gP8sclc4wN5g0q5
AHtJrqJTP2sNoYqw8f8bMoZ9Qok5kx1kMkrjps+x8n8xxD2lvI1O1hs5McAx+XQN
/hLOfaQh3vC+1ap3CLM3AqRXrfuzs+TlinDB2wfMAqwMsxupEwmGLOuhhXr/r+rs
W1Vyrikoh9xVhJrs1SbJmo4Kgb5h4JGZx47fhzlvjytjWpKwlDwe4uVQ35sendD8
azkXN0/7PJ/Oc+EKaYQKFVYYHB5Yx6JXaWviyH0wjC+XD0BPBmD+uqJbqoNrt13J
Gg4chXB6Jv+DqH7bzztqLF6/UW3gzQFZZzG1V2qmIwM0bTUM0OqdPwAhsPn3jvSj
6aWzp4JYdFqBYfE8ESjQJKRrfdeEIrjuLRK+anwnP1dzFP3R928Dgqr1gNW1BSMr
2qQOhNRYZO6xRZ5EDgHi7N4usuj20xlbbOg59nPL09DJ8TFzqrX8clUsF8Mp6hCS
chTKISHtH7skwtoHJJA36vCRtjoaFWQ86M2iraWKN6TWDJ4SloltVyuzSyd+JtAP
/564thsPpSvxBlklTMWnEsQJlQPArTCyhIvzj7ga52my3htI612teVGJz9IGxDP4
DRMOu8A81ca/Lrcyly33fRruU0hWC1Vq230hJArz+rpkIxDdaiUD7M2TEttdCn9x
7vCeurlM+mGHNl99VFcLUrwvZUbeSXRPF2telnpAez0cRlZysr1oCDjPEimQT06v
dNgjyOvzNXRd2DVLNvHBtMW8aqoJEW0GxeMDQjgDYKJT3JBKOkLFt4F/yyKAVM9j
rMBQ6eJ3kqjni21eGMtI0+26BM+VDGZCnx4Uquiua5qkdSyIK0XtxtgMrS5a3unR
MTf4XbRfrCuMIjhZqh4frW25IFstDeOp/vaXV5SXzR92ggLb2n8lwHlz3csYWILD
VZtfCxs9b+TeS0a9IqJ4l7GtVB3CVXc5KDnGFOlMXLSrxm3S3DuSEkwCD4ET1exR
C3KvUEiVjUCpwBiw8k9Y5Nr37fkzN8UOV3JEENstHvaxld9WsHSp4WV3yfrAdBRi
VrgXsiG67aKlTMUXzPlIuEPC40IcvsR0dcTRtI4y6xI8d6m5azZcr7FkUJZcA/9H
hxtOw54Cfok1Af42i4Q8gSiNcSmRQUbe0BTbytLmvZY40/K0yLcrOwLvcdOYCEZb
PdQjdk5r36Hz+6tEMT1FW5H4RqK8NsvpCpeQOPVMSNCyCr3uBcpb0eOrVwluuDLx
j9mAmjtqT1C9fgb4e12bSWTCc3eYZWa/N972xcu3TNzm9g/eNjYMXlhN9GJ5tEF7
SHJ+U8IWUKk0kZqtByN0Mk++tQiLinl8GjEnM4rf7fm/EfH3Wp82BzjxPnu5KVm0
isjVvilvIE2pwRhzJbdNyjBUPsCUmVNUalqGJ2NCiMnk02qIEEy/jK7YHt1ON0kO
5MOKSs/R28xp8oLcdqus0HffabEmwe9p9Rn3eCC+62Z3OAL051JQ/79AA698GHiU
neHUuwtYSv96fRkZtzITNCKyU8BcK9O8bUqdJfHYf7sZMm29WMOoPwm3OZ6YOsla
0nKn5kcwte/CO65Drh3CFL1uzLmBFbT8ApD1hN9mhAVeuQYNpJa3cHReqD3QLNaB
IrZYvmttsGWHD3YIhDL3z9QOwLxFwbj/Ho8253nnbQlknrEelc8Pa6yGZ6Iyxclp
5zTd9xCZO6afuMPgeixTc/gSMjntpxPsY50ipH5QkyPrFLKfVYKbsy7BJomyXdDP
8aFCMwqqkjH65fMw1fm7vVaO/jpNHhjtFar1SP+i55qgbmF5iOyE+owV7CPfhFCX
UJnAyhmfBCGk53TDE2qoAvUvc+MGPVu+1qf83/KXFF4MQ0DlcTBy+U2RxkZVOVRn
du67blTdvHXPof/hFOiQ1AwU8oACNlNQ2bOj40glOwgFJSNbB+SREjsBW1NWdZ3n
qY43YLv3I5z6WcXIKnlub9uqDkjGMnahblGTn++FLJi722fi9Rnl9kj2tKLpK6q7
byNFgEADaj6CIPZsKC2BHXo508iwDgb6x5dHO+fZDB1vDCRHx3OP0cbZaHhNr799
rehXNxW2U8MW03UOCYzgrULEcCAzs8j610qyUrF9/WZnD8TM/XJikpmTjcfzRyxE
AX6DASAL1imAd4TcXe35yQovF3BrszV90xyPFM91jjQZ8DkdkWBdelCdN39x4SPb
Ml3rMKeI8V60ZHSHm8jm5Q/1eTcaVtjLbtgmFpVzFs9qFrLkDPIYNJ/6kPLJnIeE
AHZjkZU3AvlZj53F3FTwmFTpfHSjhrV+divQrcOrW7q5O3Y5gwBbp+ozx90ESHrR
Ew1Q90RAo5RYmtCPJytnKUqCJTG5WR4dW2gPUFc+OA3mghuQccPL/xAl0cKc51w/
sv6lYBvLp4Qg6sLQzmeg/ynpqisjgpj0aqIbA37ULoOcATkSVrzyyoZ+/TqJay6N
4tpjpVkZdSZVWxjHWG9oBxb/bhUqUMq1fLOE6pd6FYG9HBkW9gPiMFirF2AtcO12
l73nz66TkrNFZI5D7cE5snW5JEhe10EjuDk2l+kgsy0nZEwjrwQftHwTmcTRXKNV
KDu8qNXNMtCsazPIXq5z8308JK7Uk8QVqEQsJ8eqVwESS2+mxVj1IJ9ssPN7WDQd
Mo6cdIlOBpivzrt2B2twwt8cySKRujnx3uWOY8c11gKt1RXOwYDhZCwhvf2UqTVp
iBRunHjOu39WF1+BADKcXkUsxcxxO+O73fs/+Nt0dVljtIMCPVdH4zk1/WrBs34y
D8h4rhLZQHSA3LVYAuidQkbvaeUOMds+X+Y+TtUeTXt16I5/ryKqZzd/bVGyDOqm
Tq70i/fpWLEEuQOIYRgIRHP6Ug+pmALs6jBYLGeCv8o4VZYiqa6HmKDx5aee8D2v
xiCnWETL/SxcG05sb3SWPIg1BDB6+kQsoxJjxUXISC+v4aUp5t4Iu+P2t6byCZ/R
xKk0hiIiUfNhbwJK1zNcS5GLVdajcZm2lnzddQcobOxfRKWRY87g1AQn+IgqUaap
RxgBuCLOGRXEULoWfu0fuLhkJS2YOip0bsE/XzRJ1g4GfeW4xJwGQZTONaccmRO6
Sg9zEr+F43114PopsU4sTtYPQ8hc+bCsgfGbEqUtY1c1ERtbk5ZBCQ7OrZD89Pys
iPyr2HZtcNerrIq2JdNUoKjeVIfLivw+q1IAuk/nBwPrqRUOb/nVrKHszST3pC+F
8sHzDEUXVrxpe9bWod71ZKrgIeAA4DEj1AQtZ96On8kyy6MaK17zUmm7H0oZx34B
JmDK8RoO8ss8WGsyZpkJwrqAxayxpDbASA5iYyRN/VTV6m8N5PR/EV5dwKDknda4
CSR107ZYV5jtuiAe5cR7+fSo7zGAEwia7vwJRQnZJe1B+D/kqV66eiaAKbSTjohe
iJQDqyz69HnmIZprsv91Oe8yMcnXBIL0GLcAqUJHp1CUv9Df/Ta8N+KcOrgLCKV2
/xp4xxB1RKhYhNqitkdr5HZOH2Rl+nJP8eX3FoKc9M7uX8fdG8lrpf5scqOlu036
xc3j0FwYSS4VNCesgehajwmlhtn2fDTn2R1fiSXSlNQLCujMhZm6ErgFBba2+K5Q
D3nfHsmrn3V5VWooYF+xxfR0+k4ZsYolge2U9B1Bi/pVIB2hbCPKE98sKIwZYoik
vzP1KPUGBndrdgxeQhOK7q9mNbmCkFO80lk3hrfAnJZIn0ONHRU1OEFTQBUS0Fuz
UPmR9km85zAhferSgT7fYaJ0rsumfsrGGxaYNxkQYXKY/7SmsencUOQ8D+udAV0O
Jwa9XdTVGrj+zkdjY8fuFXHkQvFAfdtCloRI7yDElJrQ0+GOoeeZXSUhNkAFNNms
ISEx7TTt1o02PETojk/5wLgK4mvaS+qYr91DQVcz9cG77h+rww+YE36Mh2xAoq0f
cyFWvTGF6z3TwwDTP1XpkW9QnEZK63Odh0rtKxPYkIjD040mNL+qqT1yhP3T9Wy3
cuSCGRsr+3zK9n+vb1FXpk0r5QunxmZbSj7s1zhjncS7UbN01qOmEwoE6ueYlawm
z8V1NNGO9MVBXqqH3ozm2EQrGymDA68P+6saRrn+lgJ460AHLW8RvjF2+QjStTFl
UOw2ixzwshYKxSsPBuQdpAYurEFxLtWde8SCKnPH072AZ7dqr+pJccdHPnkHdNzC
4XwRz3EYYekP8KP6Tz+J18dgsc2KmKpCTuA7pFAeXZ1uNVlgFpiOfedqllLlsbZ9
8ovKvhHaAiQcBHm+Wkm/Hny52J7YYsbOrrtgk1urx8jBmRaCefMJEmB8ndpQNufs
sVjbmUal005FYNWPqK/DROsEtDhYlvmi7KcB7F/XuIDGH5tCoKM4kt0+wUIE38Bd
L8kTaiQKgW+XNj1XVyB/9jRcecPCvPowVRijoDFWaPnf297OlukMo6spdKln1jlU
mQmYkZEm0xp1e4Dek7MDp7+E/8iZW0uisJtlhQm+1mGy3eVAOQZgFpDPQmvHzl4Y
PoK8MY2zUryJa4P76qUQkWW+1doeTQIBhs/XSindSCS87+Jnj/DeWHPLwiCc/1yd
qfnsE+//hcxsUL7jP0ePjycvmRmZK47vttkMNuWMQWoykMri8tOADVdkNVDYBh4Y
zgbzNwxDndsKZWlUZfH8Rrwuqlemb2V8eQzX2L4qJjHj0QOu0iPIVsUUAt0dqI7D
95rndYLqJwQGIGKnDbcELGpewS9qJcZMN5H2LGgx8lCUQW30c7uANeSvi46FdHAp
JnuCxtPVj1Dqz5vXfsannUhyGPMups0biyMpIG1JFwLSpjqp1H/sEY8JlFGxIK1b
b/qGXv2gJxYc6nXh2JSHAuMhGYQjqi54uTS5B9KnD7UUyaMzTJvCPdico113sj3I
a+ZURVG2CX76hEIOmKxDaJHZVFraTCsMrLaQDs7FkB1yCtrn3R4jLqQF0OpL2iUV
MyHYU83Y9EnaoixVnd97mjT4jOkbSSAFe4pLu9r59Eoo/6lDkHDJLme6k5Sp1zLa
lN0xXgSvs/gXxcEF4c9GKhFrlE5fir15sgD2eCQu41cKdGS+5hsWFZL0sLXCJl5l
29cJLIkWaL3wICJRN38rYN9naFG1gqHfaH/buI3TPJzjQv/QjdSm2a5XCxPl7YK7
63xxF1/W+PV1nV0dhImp1keRo5mTol6rCX67XYRQc0Im7D+QlijEbTtw2DPbk76Q
uhl1bN8Hi0BMJhOEQqahzbo3EzDtuX9NzZlUiY/u7Plk6NME43nW1JuQioLHzCiI
rOc8RfHVsMo3bx9EYnAUpfRbWO2v5TYp4RvZ81yCrZW28OXpL/O+Vpmf0YUFbFXY
0xO5ZiogYxWwZ2Nt7jD8cgvi3kGd0i97dCvJAHt8EMsNrU5PJjsdaz/xOaWrcgWz
aqpnsyQnPmY73vTeItixTXligH90b3x3rMkZr0+ocxkvBJb4jAH6pCEyDnIsb8HW
x/7+oyOhWm8bWcnKP+SQZVEiSuKH3R/XF1tDkTmQ5gmytKkZgQyUVaJ5W1vpxLzN
jxnxiRcvWG+QtWPHTVZVL13k3lIhVoXo3AhCGXsTvBvjTAmgAeGa+jFQtX5r164G
9KP0axEXAc4LpBoD3IjZ8E4lKSL3zB04i6OWTxl25hkWiXn/KCRPsKG5aVU6CbKK
eUG60zBy60Ha/VqgON145J7qvMJeg24ks4tZrOfA5o1tdw/hA69Stf0GD4EigP4Q
FuPDAp43qQkEumoJqXZoxfTToWvSvwWexqGyfFa7RzoOkINrOs8aUQCoaBEknubN
AMkaUN2d3xeJpmcvoGbS0knjMB/hKeO5zxkevwwhoptSyMKvetefaYB/zMy6BmuE
4Hj224Z0wlF8p9jWHwAH1AyaNNtmKCe7UhOI1XgJCwUgiu5+JshBXHfAUBsqqIN6
QnbRHeicTDb4bNxy7zSgqEeCRk6yb/rkNbuMgPxIfn5h/zvqOLPEx4akKYEZO60+
qz62jaOK1rSbnPjR6KNxkVnS4Vc6BQnglHoZCI14LbTUBL9JbrWR+jHNfgx29YNo
FrW9t3IhHFpG/RJXIeFmmmwxyd7qjQrDdMwae1UCVsXVyYe0kNJGr/mw6MIH/YUb
V4jmTuAbbdsUCZtaCYoPWqo7QYfkYaa6XlK4WXc5ZfpHTOXRBevnoDcVLwNubmAN
p1gNMX8T9G+He9lgtGoF2kw2vpbEcerRjhj3QaW56v6FI/aER7Bs/UmI882pHq/e
0W+CpT+UnBwGr2vwdeW6b/dnR1Zn2wAUjFW2Rhk/bYz1sv+XDMv+odTmR4IEOzJ2
RD8UC5E/6j3VgthmX/ZldEZAbu9m5UjxhfIAZ8zbR1M9PO3hXy2s+r5RH7osl2vS
sYpL5ypRius0zt8Y4QsnRg4eTigv+AKksy/EXAamrqukElLAecXEuLCHkLCjYPB0
GQxNJoX73nKAAnGdUGEyU0gYqhHLihXSG0ZCSh60a0/QSfLPU0eYx9jhmHn1w4nw
g7shYy3JFVs4EfGBZd0tS/ki6zQY63+P7irF20bbo3CE0fdSfaIZ2MnUZ45fPdkc
M75xzxNgC8TAlJys/CB9i0DiyHf2BlIuIOGpHALWSs0MffM10LLG6ZYfmxynAkwF
YVhdFbxJNERCcEE5wX75wkEiBXKJqNFmcEigCkKNop/8FyFfskZnVTtw7OvLVngo
c14nr5fOjZ8gh6S2bdVlOA6AIomMx45MB3MQ4DRfrJn6+La+Ts2Zk1pL1OyhnrHQ
Yyv2KvXKXOARnoLwrCk2GmB2brhBBM+PEGaI4mmmrFdqMj4vct7zCwM9rLkbhV1M
DE67VORrOBfXLEa+zrOKvVLelJdkfQY2FfJoxJcwrT0JSdTsw6j/6l4QH+vV48B/
eIimH6KGNW0atGjEDOS0bRRbGjq0I6j4aZoZQGn3OmfUZ57zcsdmu6biy+MeaTPL
5fWK61d1Ese9Da04Scj43BpHGlZ8rrniC0M/6TKTAzpayMQb58vSsLAvbxF84zb7
NBcH5Z1q/mVDFMkUtKN6uEsek49gYDCXzjOSLAPpKMkRcTTIicX8B4oEmeUmN6E5
qh0ahCMRtJpbb4OcbODMiNiQM/qsZSk444UYF02gP3wwPvI6tnQexnes0otOjjug
9NuCKTt2kUhjCqjU0MGsaWOdYdlalY3PN6hPH1tMe8tDhFd1o2dgHBF+IvINjueW
3VpIxgGY0/PWpb+1bVx9JbOepc1NVGdyCQB0LKkJJGpBVzpbqUgtue2zJlEM7Aj4
AoBoxrjv89NP9WDXOzEFHQehceBaVvapzlKmlSBtWt211tiCUBFc6BMQ7la6mORh
F74EnCNjRkL1ioFJKSV4BijQx3DjqoR75mugP9yNea0bovLLPSb9bndRhqbTBaku
eHPA0RuTDapcPOMGBRcL3wpKi2kt4NV7hpc5CfkTPkuDNpQnf8/bRdu7aF6/SEa0
4QvMBi0/RCblYuvda+P7pEBQagNpA0YHZmlPipTcd/nCf+zjYP9A1mRaedJghJB4
6tzxHQ3SToz0iZKjIyO71cBEMMhyHt/d1BHUhCK5YYGaYcQ31IA6d5GQmrhOnSJ7
fg8oXw+A2lFazFuN5g58WCx9C+Pk2zDqfrmwEirCIjE95S2GII5vvEgjuBb8H9Oy
y5CuSyzSNUe2Rvc0xIpx4f8C3aXpUu9fiFssH01L+f7CzE2DkP7/tgoczT9qTtHP
Qk6H5GHRS0b7ZzP7L1kENFJZ39IlmKV7mvTb9lGePYf5enP0LmY0OALR7bpcOXM3
ss2crmHx6gHxyhNPlOFWPJEh8YG+fsS0Yxua+jGeDUKcdzGur3z5t5oWjDQbW6Xz
MjmWCtnnDgod3/RBY0skyLjzIjsm3ivoMo+dY+Lh8iOkY7upDiwf5JtPv3koynC9
evaR7UAQAENv9GTB3spp3CNMsvhgo0MwUoafXIo3Vjz7u8MT3eRO7L+EvrrcSYlJ
kXNR2DXTAegKUHqyLJhK9kwqwIelNGJb+cRP61TuYF/gxBDQjtLWN2z2UcyWrTq8
1IjQwCeIslSSFGSQE2gf5ExQFFbJEb6tmKGHtr5RkOhIUoevqZUeShbNjtso6ryE
HyRXyoFCGk7U/hrN04iHLtikx7ygjLiErgF2bbcZ1y+pSWRWqX3rS5jb/EPoqpSZ
PfqJPgXALmUwsjdPapM/o2Ge2ipRmS1vvWTtMXGevCq7YEFPqvfBEBmpmMlTaRYl
12sPwBpIPqeo/pQEzEUNHGPXLQisZEAk8UwejC92yO/tubLao9nPY22XWa2Hs+n0
5kkM9bOZA9P0//qlQPZ7ER5JXRjsgTh1QPV7p8k/r2JpF6atB8XA225vkf6y0Fa5
MuknIBC9gg6XW2+tQEC/rfJWde84ONpM3NSO+cAn41cB5dtz4QsbHcbYU6Z5ZQh9
p5GS77XRigY6D0+HsvNox3kPma5gUs7MJTeYwlsntQ2VA1IIntM8gFvJGYX7hRgj
Yg3wSY699yw3LqOybPRFM7Kkq1ODkE/XRMEE3SyBuqbNGxPYHNgYJxHWOfxSaL4D
uDQ0ivobYyFpA7poIqRZjx/PdK3aLnmls0q9IHJJK4kmHcl2Eg9vKw8iQt481Ayt
a6TddG+/EQgGJ4O5GZWFFd/Avb9XCcFaiT3cKt0teJ2TL72QmjTiBcAJ00nJOz5W
AnWS6HYQBOj4vmvKoiIMM6UJWmBymQewIn6IH56v+240wy9eEIh2rsYZsgdufOxg
ztL3Sf0kbaAdLhMbaep1hydpilnsWWtzDMbDpTv0CnRuKQyXG/zYsiV6zFijX2nj
GjsNxkGc12OYk9xpVKlhT2CLrPJ5Im3cpLwwmeEa8ClnN4SwzIPWP8+KkxdBiRVO
VDNYAtDxzAh5Pn9f0hgMSTI2vLVEbb5/OSNKQJD6yD9LOCEn48aAKcGlLZlowrOU
AMCYj6zqlpoHuNQVt4RZmgn7L1uM52i6NW2FS0OVtV4TmsDnLKlzywWnaMeVrBud
4miHTn5RGhAHJg+TB0wktSbxCWMwNb46DkXc5/tQH0u8FHpvlntUW0EeToTNKq0d
u0jZGB8U3ParBj2heOGaYSLwzMQzYmUB2S7Ia90fxc9s6P87kh/gol77SXB4onbm
vxec+Vn7G/Ag6wKLbhk20t9SjVKsmgTrteJNoXGS2jqmwY3NXBOCpHmzfbngK3Pu
oD9IZExzy+ntj8XU+lioAtWffg1wDDPHs02ATFRG4X9s/qqjx2ZY7hXl1PqijXjc
1YqqKOh0qwPeQDbFvlHPba6qQvzuqmC2PqlhqmE4+MceiED/krJ8SNKixmgnfSMW
QL2j5SUA/08kMBoS7Kj/Q1dXTNNlybfQOkTl1b5COageNhtav+GBVH6B3o7e344k
Msb4nWFHSOKIEIrp1g5cYJgf/bguuhBcIPBBGvXavqjPfguLavCrcmlg+0KY7Rfa
ktIyANeCNZBWZSgB7k6gGBPCRHnrTm1RM66StXw6k+mxi1E1SFuSYhNMbeNXK3xC
UsT5gn6SnyShrIz6bPCjpxN90imZH4snkHkkVBmN9Y8pTRzlQeZNgXne4KTtJEsv
EMmn3S0QOZrUsMHr0fMD0T0w5U1nmWv4QLLpFK1jf1SnRDueSI+EunAWH5ubkRLf
cqG40BzmR+2eeFo75diD+fyosLB5SNHQMr10E5UOI65YXhfI4eTYDwfHLsOiCRxg
nZo1+yuoa92e7w9zGabHyMNM1Cw2MzrizvHAsV8eE6Wk8+JkCIYq8RJiZosE9C3i
jQEcqrmG8FUc93Juqq6OU929pza41eafr52hgzNRtiCxkf3rHG4YrJNgM8Zqle+l
itxZiLEDZ8u4UP2U8d+NkR0pjrmW7lYVUNRtRYrR02A7mIsQmwVH2aYqbi5pxFVv
w4ORyDxVHha5c434QXDpY92DFrU6Tqkg6gW/YAG1AbHB51kOger0IdBZ2eqL0EQk
8cvGMb+2+jCP1CJWSc079i4WSs2eAYam+Z392EMYwy2z4uhEq4Yacjq9+89rOMGH
L2nrSIUi929RTXGf8/k40XrWkvDu5g1DqhqPPi3roMRKN1p0Y9Wdy4dY5mRXxa8L
DDyKSYBkHupwcxZmpLQJfLQ6sgQ1eL3ytwdtGd7Faea53iveZ6fPHrJLJNbFIqQP
RUkrxfXMg5RlfqVPZfqU380PhNi2QYpVSG4AZjtawoccml99iApFYBdee386st93
tpBN7iEixR1Djx1nsVosmHqpSG3opgWkTVJn8enqPTDVxftq3IAj+XjLGWbM3Sqk
T5FqWE5hrYpIrTTT9j9PePFlwMO3tkwwiKo3HaSc/bh4Q3Pdq3l0UeqfN3KejrtE
aTDebpjQfXJRe7FLJljkQhLgT6FWv6djpJRhRmj2aKo8sjuEd9eVXO+cZknFbANc
HwFC0+JnjxKFgHQzvb+0eS1N7hNTSWDLf/C0c1RdciqqPvlnfKaN+/5W3XXHlT0F
fuSU7WjTTi9V6f4q0bBZUn06TOV6z7qJDQu1Phm6Yi5xWCEGIcF9vtZez1EbF7j/
iTl8lRnZTchQX5bu/wzxvI04OK4Fp/gLYHITcvoo/DdJd/JRo7oRSDJkQdr3meZe
fckXWmgweFxIqZnHBRkplnw6ZhZbhmv92GpoqAff8mAzdVXa6vQWrmQ2fGi2TFfb
YuDD1WnkIEBHTwufiR4SjtzbntFU/Dc6jXtivrH4SzYewVYhsUUh1Wmnf/nojpnZ
W2dFM4gUfSysvV+ak4r/R/3m7xLzzgaZa8nbaSjP3ltkxF8FHSM0DEp1Tm9U9fp5
ka0ocimqi4t+Sq1GbHdMWV0bprVVog8vWYOzTrIV+j/05KylMmQPrXJAFyBIlDG3
TQbqIEMJi56le68bWMOrGswgDpFhWVffYDkdHAqfeVOXRQMtrGO63ib9OHV99j8+
HbbNiuUXEcY/ljRZ2QyCemFD0OzK5XE+3ZPArU5IZMK5O1Vw/e9ERbvTTovEx+Ox
QaCsF+bdFZeVoBF2OFftUSkTiMlQH11rHYx59uQslvyvo40r3xCfmPfpkuBTF4lv
akuSnjijjZ8O946eCF4RvvNi2wnbslE+BQJabyxm6fC4c6dmw6dTnSbh9pJdxgDy
uNKOzAvu+pTK/ZyiFqU2mh85meyBVA0k++Eev3TArp09n9oX5FmxEcdt+AzkXJAI
c4rV2sM91pmnb7mxZABp4Mm2ClCFqE0UXRCfp3wn1HTzVRH18RGzlOXDATWyI+xx
2FevaWayhyjYC1VFn8a3coHCoyLoY21M6r7rkto6xe9ePweVaTtaz9IrK+8l41c6
SUU/MmxcFVDNUiAWNnkZ0NXMLsx1b2kABf0GRIiuK3XSEW6vi6SFSQpqDH9B2M77
8H4wWtbURPkSaqofNmJwUWm4+5gPXDTwddr0YV2UtDnSeKbXP9UFI/yqlJeCZQSs
HIeJaK0eao47WEHi5VcjJcVF4PIjLdaiwsKiybbIFGVsdIY5d5TK0RHWCzbXlDxp
K2B8jGN9nfpvVY5RYVsjrfD4noUFZjULb78SkYMQy/JLu19wuhCt9++KJdqD9H6N
ZY+/n+fR1hmxjQC14OZqCfCM/NshxcJ+r77c/PYkxH/X0Zc6sKr+dvMJcKlLuBoi
AAhSOAsQs6UscKKljvRt0eZuxa0pTur0wbO9xyzmLscXRoaAF/bXYgAyi4cvkMHr
eX5D5U5Hz4vjwE0jt7DzVLWfRUXUNEbeNo+b2o3OYTsco8K1W69tYMkzg5HgRuTH
NBaAh/Ya/18lFyhzcH7dmab+JfCfOynxVdTrzt1zqM01jgUjLv5MarLwvxZqbeRr
xnL7ZI33TJ6ji6+ugQQr3zwpK3guk/6of4Sv2sIl60GM7b5HjFI//MZF+Ts5cvcN
2lgHUMc/MQK+60M3OtzgUD725FLxYm1+JJSPVWzbJ7CB9EjHazcVgCyIRhGCdAJs
kaFmkRiZ77vrJGLwjzQugqsLBdn0AbONvKlPzZhbLaby9NSXAe4JSYtFOtQwsm8c
ecep/cwm3uDImYt8sKNmlIcFVITPnaJX6mubTd99+s/h25iZwVuLTfHDYSzOp6eD
sCGUGWBA7aIInTD09abVtvIR04qr76fNBzeMQk3oLr+z2YpKDcGJdX8nb3i8q5Vz
gw98Q22TLhtQH1cr0gzTIkG2prjoI5tR846hpBFlQHZW1nX+JEJ3ErgUCw/iMxGg
+6HRKRrePWdyXs012QXO7vBUatfs8DtMK/MuFerIRwAG8bstDAJqIPuYbr25QWaU
VYzFSWmU/UlEJFq2/BrpHVlgR5rKbQW0RRTv0q8IMFPs5vSInlMa+ScpqIS4dLYi
FeCvR3MfvQPsyRUetkqJiFEtJrNZ3RDKQ34loDh/925pkuPYQPcFhAP2DKoD0Drk
HgxVHy1fD+m1KCq3PKk6+D6tSVL215F/7CsZvKSSeNAF41RtXjMLG6kNtEYBV4Wh
IsmmWjTmhpOVpo0fj+65CqWfi4qNpXEB+Vyq97vlDfQ5v2FF//n2qeNqLjQNT+iL
OyHIk1F8+HRqvwijhZzng6ISBPlkXnNqQYC1c4TycIbqt9EursK+SR+E9V9TD554
pcMWrX41civoqpo79Y7k4Y6N+aNR7YpUuYn4KFywex28D6z0pBRei+RbsP+ZyA37
O64sp/putXeyj4GRfaW+H8IJjJaPmLapOwSQSd1C4l37MK49rDuvI2NzE9+r26vO
+VhO2mS4PZvn/XkpmUnjNGt/vUQHJGrh7rcLL+FS90stBxmA0f0pgecAo5LjtIH8
3vg80rrLJNwAlCiDJ8fnsgczj3S67ss18KdhdP/xqJ6+mDzaELyjnTF7rXL6LyJC
3ordZ0vfwIgkcHT5MqTPzNGnRQNRA2dE79vq+HBF2dUxxW5ZnuXW2SKhPTj8YjHt
0J1ckbaaYlg1v5Dq4ewn5arkQohvFKom0Ct2bTkJwRwFIcg87mACRwD2U/Vb9Ul7
NBbPceQgHCl7j+nvpc5W3Ed2IfolyP1E6ssgcmByIc9KPfe5tXZvEg7ci5jZR/h2
KtoByEZR06k35ayZbKrL1PD/75qLF5kuDKyPbbOtJJ/kJy2WFsL7QQjORGTKaqOS
p2Rq4wvr4A9ncqGIKNuXPSKOLbketpanUi/tBgGVMxQIIVgMeYWBhmljXe3Aai+i
/AdyqMLPbt1xSQCwuqoSKMWUAGVkPxhIjd8xVbEF8QUIMIb3kkv+EmTCVzt035kV
wP/JJDsNAkziAAWMQ9bxuqf1K8xlUaLtn2EFkYjNkcugGWZbSmW+Fplo+HzVGhqf
T3BChYLuezyOBD9c2b/+a4vOfhA7kxDuAjC8fjAU0HXNs9Mfiv5CHvlCeAdrGEia
989+rsf/xfBHbjqtHzG/Z1+PMJrbW2al5zvtrXjeib6GoaucTVjTq33GXpK2dKwx
lkaTK90YOA1LXyQDff+Gjlv9I+0FSy9cEhdBclQ8bV9NvF32DsuVTtjv4kwuYxIK
kgbdUmXE5WmWvPWjFQZV3KBhtK150fAWNpdbdjAdFfgPAcHSKVu5nARSAd01ur61
/1N9bnpxLpVDIAMv/iIOye+iB+ROzlRJC4PCu8LtqPlHDll8hcusj+y6ru4Z7jM3
h2kLGQj/YSHBYOCVDeAnY7u0obx/ZclFSCU9pKzueuIpWFjC5arpnb+poYJyuaxJ
yHwjRFlPhiEwgTBoq8niRhT70ZGjN7Uwqx5VeoGe8jALMnjBW50sjD2ppgRvquz6
BNP8rJ9OhUG2nCLpgspI2+cXybt6hKBKFCDlTHvkgNLZPVGFSBD7qcF3idHDxFny
siyXFfy9fWs5EzRKEege83tSUW/ZB/qZGqOgPJV2RYulMOrMrEC10WFgzWPS/nlI
mtCjIYY4PbEcUMN7FgO/gicFqnYPFg4KturjXdmmQySEpkgfNrXLKAsji/iE062O
76nW7MS1CmJZgptYmuyraIzQhdOUMYts1jnT1Pp9piXzfxCWLMd+HOM/HTtYhcME
ge7RLfVPihN6N6GaDtinRGcgsVBrgXQ+ajI53s1oTpsrlU9m4Em8S1UeR/Lv0QmM
etL4HEfjL3bpSi+jhkVN736A2ntCEMpFAcbYFgoWhLByx4+PIG5lYl6aJS+kKLU9
ioYhMKpKpRhv+LLEYtCV6oDv0L2mhX17qBCCV86KvpkD4mpZ+uqhUjXWghXHC6sb
9S7YAroudamIHT47r04OUg2asYIi3QNyyBoref/SYdakEI8pbdbpm7z71EMmJyP2
nBm39+Tstafi9OpR+F97T/VT5nsQAeGISfw9E8JcRE9TuvE9rksnvd+iIoQFGRN9
+Y5Pk8RGzGZq9aBzbmDHSfdMECc4TxdONtsPASA6Aj5GQy4L/xBy86MC2zYvLA0Z
xYKTrPfyQdk5kvDd/6fe3S2jOU8S/veSD+GHNd94uWx1qhEuiHP2/Upf1jSteyFj
3hqNV7A8oBZi2xbBVvNSGJMxugyv0v5DVX8PN91OfyTYGE6g3CQR9GSmB0dGpmeq
NrAKsRB2ZBD54YjJrFKNtsv805ktsr3XEbLAQRNfxRN8vulYOb7O3qOJvQXDZeX5
RARpctuRPOIz9Qz/mHOSQfqyTs66EJ6zBBqW85UiDuCmmkEusNjYc1X10Tx1xNCR
8cumrCysKKZMCa93kUosgmbGHrqWT+lEEWNU5TMW/cVTFU6pusMNNOSCezFUBDbY
KOV3orVYew04mQlOSd5u/NHsSJNtkivKsXCzb2MXoW7oHL0B2h3EHa/2md6pROys
vSn8B15qWVVf0E3U5QNsCtVo0hY+0TszP7QpGhiuEMahGjscHlrrXALAHq92hg3/
tuLn9oczcHrgmKXVDdFZBs3uasGlbzOCHmWb2kuIVo477eJ/YbBq1Da6AkIRsPhD
MnEfdRDVpSgAUSZPZ+aT40mOt7cOYA3SKMyNCorVfnmHF9fLfTEhy3oF65mluT9h
elHYIUqJCGGpWF98LoU0t8RbPdDywdQ9mh3bjoyiw1pjSpTWN/c2gvTOsC+V9l0Q
/fpdfvnL3tNnmVCwYWdedr64fS0gvSWC+DvI1sUPJbiUMJcffhMhMgtR2p9dpvbZ
6/bUZpkG/ykBfjm400oEdNkY1IsnQa290EOjkAZYmf7vkwlA96tXEapuA6SIPxVZ
qX4+vUOotXurJhl1OAXyJOJFc2/yxSgDhp4p9AHNZonH6SWK/4U2HTN2x+bWNNRO
8GhTcd6bMEC6Awyx08RsF2KzKbem35YbZf8DmpPq82dQ1epL9W3uBEjaCPxs7V6M
KHDIBVgHUOGL3/Jc3dsChVxJsQMihcWKfWsmPz8uSlQzL4084PyC6440jKSX1t1F
EoBMcgdalo7Dagk5i/O7ylGMn9XufYa66HbNkNLVgDb2goqMhExSEjh+hEpkcbNL
DrNRlAByGUoZu0GxD0aXqC3nsDijerkdVvwj9WSxPQDL/onKpQbkWdMzxRRM9OqA
rTca1WrTIoDD0oLPwEHny2C3c2hTRWmyKEjg1FPZm0JzX6iE/fsZqHcD+/3hxHBQ
7ii1UDrbsxtr1+3To4RtPlSDPRkQR+26NBZqCnCvQb7A5l2rfTy6i5zRX3ywrW6Z
ee51vCEV4Pny2dT38au5ACkhwJQUamKTKr2KiB3HF2XwjqSt34+fXOa3SI4O0jYu
NPsLZGGgkv0t3qLgRjg31SwM+8OCK73w3S+JumsX0RV4YsUKHteEXYmBiDAi2r+Z
ASACizPKDbYdTASQ8mXkFxR2ekGPtOV1XzhelllQ4eOiaVv9GLh4FfefHK3JInY9
vpTcSpdVNVRqTcilbLgupTK6otmH6WdMlQaacivEDeY2pHPY888X9/eYjmD8k12/
vBjY8HwbcPtpNk7E85v2+q6WSXeO9XERO7pvo6HbqgzgT2d9tItR9MjAi9k3JQ7e
UOU7qlCTx+EyNLBEMfRslXcFZZR0Wi6twAUlqLMDwZGNItBI9gdT3Bg8Wet/byBi
TagSqr3gFR+Qo4/Fb/L+GhGDMr8memZCdsClEp+KZwxSHT1qs7MqLXQKb5xrZT8N
k1JassBj1bEYpaNtQJi77oHUrSbtW8qOdrHS+Xu31roexKQhmhCwOhmY56uVITfS
D0/IBFm7vbniu2NZe6zAb06swE5jRpxUhdfpfzm/qtLIFOhicACT9Dv+QUdsgwFf
D51ea0osDU/CFqVy/bpZwaj2UcstrstyLSjLe1OsDvXUQhMHzbhbfGU3vKrQYz9S
yvosgY23L+15MYDnJtqwj8VviRc5nDW91Ogr8tS9UaeuzEiLnh1Zn5z10qtTjRRy
lxmFeynvWeUKKIMjLDxzavFurK6Mj9cifGpbNSDVB/yiRBjjXdotQtj96JCocu33
XpbyblNzhw7hkfzQcFH1cZjwN7V7YBSa8WtFq/4Rm7YPM6MxoWp2p5pUCwtyjKH1
PD6pDmZAvd0u03EN69z53jVGR8xRVLGsl1fuzz+eBB9JHz6mylluDH8PUFL2DCok
8hI89JE+O7o/Dprm/Hgf/Od+bL9iXCMEh0xM4fwd9+a6E/eqH+WvR5hDRQYL9/BO
u+F82psYUDwzbk0mMBDf9QhTcnw6wR7mmyzxbNCfFTxyZrQWrdZ70E4B6Hh7Mf7Q
Ci896Rb0m2ZAwGB0pbgcSFWXLrpcXU6H7Z1N/fdwBla1nISm4rmYFp2Nuc6FE+nh
w2vbnsmRDLpeiii+s2dL7t9NW10SuXfGuENhQgpcXdKUkMJLyJz+UgwKAYy+cD5o
FhrvCOkDb1Vn4q4NT3p+WAEPDBQZcBZPGaM7OMYtQ5ghXFY9mTnmhJh6mP622IAX
EBsc4K3IJotw2DrVLSbTNExtF5yrme3tRYYMfnb6pWSo/eD0S6wFQhsciWDHSJgk
U8aygnOGQnF3sz0BYJhbtKZE67+X9wfVj67+ESk+aaytA5BYeFNT7a3AFbelm20E
WR4L9OV5Hn0pv0M7NjSfIUhEN63Yjs/PSTm/5pQ/1yPT47+yB5Vlr7YAFGSbNsgX
uN4tWHlzRMsENZRi20tf2gciVUNgjCK7KpmIR/rXDFwZZqarnKcq1aWUD1ci6NrP
iY8NyFgF/mkRX6jgeTlMLPvqzaqqb5uC1QBQp3VHqtNgb/wPbFEzcniAYuLclrgl
QLPcUO8VbzzdcCYMU1peRbjbpGE54peFZlc+UKuT9wJdiS/CVJwcd4TKvFqPFxrq
eFWIs7FXNHkaFS+SB2x1ePtyOC7vyVtTwJDhWTq5cuRkCxchyr4tNlX0idSrDlv4
YIo5G2nabU8g0id16EMDfKeSXKtUFxgdsSA9JpS4tfmNrfinRWBaU6MnGTip9dMY
AVmtmVhLEOf7N/+eLrOdd12rfpVAUQ9n3PnK5JRVEs3AtG0veS9febObzbzt/LAa
Nc5te88wT9ua1rDtDmhCjTxSGWkihKM9j4E+LBzduCm0TpgG53CE3i+Ns6kU/TdW
+SExzF01FEgjFyXeiKGqF4iHcLl9mBihtNcg/IDQtmOT9DPrYFOer44TVMXhlfpX
DJkLXQIw5yiIOzg4ii/eMWvMcHNtrsKyLPfFUpiaAIjY/5FKIx458CzBPU0AXQ1g
llFQFCFoIJ1IYA6Y78sWC+X3YgsdrnVMtpysJspY9UG81Y6KIpHWGEMuPzsxV93+
TovkWAgmg0YMXNKC9QEgZwW686yj9J17RXUWHuwAaJOPliyM9JrNex+9xsDaT6Y8
MI4z+OP8uJyvVa0W7QIFUhaZp2mbkesmx3mJTnBQOLiAE6kCsQrL12CWEGl7uowv
va221zdZendFjI6n7fA8AcxWLbs6Ei+/S7INe/g/6qeNz/mCWVwdKAKu25m0RA/n
as/cU2TKwa49LrjHRTeTtjJo5mcM2mgbiF5oc8JisELeGYUi+H008D/ufKsabrSb
VK2Cm2oTulYwET/ebr28YzlRM7fdIBvCRoj2iKZSXkI9yDPN7zLTpUgkDsCK3zlk
lNI924Qe8jciiNvfsZTVgYhZVehd+Lm0eNHw60f4bsItxjzYNmsb4cw1UZMCusHd
vvF4GJNMVs5pzL7I8hVcN9An+PSwl6c85L4TISaAaFW9VXxSsdXKo6GI+0IqZ1wR
41kVH4OQygBTqKztlJyJCBzq/ApxNDWQhYEj8fP69FWYhiisjB0Tk1RFLs8TG9Ll
GC3uanV++PJGmxkZ1Z/ygmHEOASU1RsHMZbQz5BpSu0TMqFJUjzk4idj95o22emj
7PQ96te6cX94GE61I9afbvieoov1NWEkrHq7lYRbnD4TJG3pIwXQ5+z+mfvZXSiD
z5EkT1iJo0r3Q/ayyEgB6+t+hW/7I6bUylril0Px1flqerTRhMpxMFYrra7/iO8N
UzDOurGM/IY8utuYxgbBzUAioIJWZcFX4judv8zpagrx3+AhONg0CsTGPpCaQGCu
hYyLKBkSsorxCVECtgR+ba0WN2xyB/Z1pSAGKmh+YF9iVanWZuGynbxT93kNJewl
rWKTLsYyvb0gY+vzIhcVMoSLa9dE+jw0h6qZtOS/OB/KwZlkrB82v1eBasn51ceK
gVRUgl6a89W3duwv21/p+O2jc9y391SGYly4g0QEXeLuK+FUzo0yveHoGtznZ2R3
awUHOCDFhSVn/leI0SrZCYL9Vcr84TJmVC0aJKmYcOqKq77/s5NgQQ7ka7gDMkiF
GE6kNg2P632ieas96uqg3+GQ8NhPrPagGCZxdLq/0mSwhFfrTbIjoOUE8K7D4WwF
QSUJKgATV42AaGQcR/FqyDAQF+db4YUTU50ak+7UZyPFqgB4Geq4qVfBIgb4r3YR
mtgGlVWpTcx4ty+A0v86poYsyIag5lkIcUby2iR38II8YTnRgjViFroeK/uZ6tQd
6vIXb/cUGsv2LvlCj0y1BmfIP5ioIoVVaesfuuEN0oZY6iE+BwqIdqw6jf8DlAib
FjOxHnXWy+wezanBLCRiSWHSK8KUlQ4hDyBVqVApquG3xTyrMuXTqitfQKmSkOKv
q/KQhrghxYK4fpdhJF2P2jFdViNxRzvBQ5pOXRHQQN8nLEv7cSw2LoMkwx7Z2oey
MLU+x/QjQn0SuLK4ndLt33GgW/yI17ZiLRhd+DnQN6CsnhgTwl7z0OTv5MkXA2mF
7GvHhr5GzYrN4V31YefZS5qQRT4qv5fg9rNXEgAPe6AYpT1gtiP6osMpK4a5hxyU
fBlgaMPuapPF7GVaZ1CLMOmEiBju8hNhcXKlp8c2v9SJiBR+0ROGLcnGBESwy0yh
ptmbSdD5DXhaWn2MqwyjtN25ud8TFwnyKHLXBGin2RFwWVSfuXnZdpXT6BRhg6Mv
KMtuoDmcI/PW9Xja4F/jn0SDeeT03CiG1pE+qr0OBNgBfEnGrZrojHQBasugp09U
jq289IMMDH7VTEAD2Zp9qxbR1Pq3xtG3vlUp16zRJC/+IICOdWsKJmhNc5Pgp2dU
OQ9yd47wKqxCZfjKZ2S1Y+YF08lQUKfAPdprBxoDVRsHOObVJ4mkStnXIUPgyumk
d2cl100TeI4knUuUBRErg+fcQrSsY7v9YLHlgKxT/mRXbV7BZhQA7cnRXrKr909t
IwlIXvzfQfOFTQQmxhH3RoAWAg4RkdY5ScgNtdXdPa+Grf7oM9T1DeX6qjPeFZ/3
vT9fbON5Xhy1fsx7yNHI1Nj0Z1nEdKS3Ub/ybY7TXfX2O9TxekdWUav2Mz3t7QAN
Z7KpKz/3CwsjKXRGr4Xl/DCcRWJj1kqiOq8Ph6d8FWRaX4fMjlMcPRe7JWzC9c0V
+Uonwk7drtLiLz+/jZjfbNURH2uKhiaEuAhXkKzdYGB4dn83f9IyvXUuR+DOQHnk
1cxNAnxk1LqNzFrpe5M+ukPlm5b1b4nHWa/y91PjSi92DCST4N1ACtRT899wyKbL
JesaiA+BNBOuPsGWgqgGf/KQe0DyBxVIYsVbGetu5IIAWpb+AgoV04A0ORN6ZOy5
z6vxmKck13sL0/kgvXJaDoAj96SsQtuNXdxuJVPpyMbJwm0R1MuLebgcYj55r0bN
DobJraxwRNcS5WdNUfU/IE+E7sibIORceoh2Tzra/ARQLBXmWHweEAUUCEQyT6oz
MCXA0iVXoUiFxdp8/Zl60KoQMbp8z+BEdqAYeyniP/fogSj3kHKLB4XzrVsmOoi1
EVyqCumJ1XmKMwlqBUwca7r0Pi7yJStad30IlssyQ/A5NUZ5w/KvUw/65e9ukNCi
iiWt15qYIW4kty4SbNDA2fnFgPiHdzt5vuSDrUrC2n2/3+8d5oCPIhR0kg6JaIrI
cmbyGb0jec1/fnnsRa1yUvvgIMi+SlWq4kI8viFLTp7zuUey2hOXQ2vB/IT4TGtG
o31/nZDB3F536rI7zpj1aRlyP1gucJ1ib1+o2WBJ0Flh4cttqaucTpMoxMUgPpvl
2jWxkSBdhPb/iXiO1R5AbPkak3TFnMppGBoiofoRGJql2jzAYOhrmeM3g6kSAHEp
nn+xUM7sMS1IP+NJ4PO1u7t/NoJIXIcz6F2ZsZKqImaze3sFvOgTFwvEbfke7gIF
aPQ7ukvjdrEvEIpdv9Hmh1ZBSMXLQfTS07EdwnXI5cdBqJiSbzXjtckJYMRZjau4
eWdSFm9sr/ZWb7tlkYnEBMzQG75RGIqkndV6ZaXzjFEiyHn1mx8MRgydCY+bjsvv
iNszdI+knkd08Q1nOwDgl4dXW4Ia0LtWZ4WZkvl4jkkWRI7pfy70Q5FZ+CtFpZ1l
JZm/p3EatC4c7+ORv4+fe6C/8VubSLc1TUTO90vdQSYdmxmCPK084FLKV1t+16iI
6/EJqU2f0LEXIS64Pa/RZoDHyF2+S3G7AMbazVKr9LPlTf0/kb7FXgJQLb64xEDt
faAGOxlAp06/TBLiLPaBfPKsBWn07enVsxsY2kW5s+4/3CnZtmj0PW803kIMV7hK
BCil8kaq+XdRnzka4baTYCBPmSqswuT+rbwtBg5H/hKrqPZFpwReQVxJxynFVAKU
IQ+fBNRkSPOFmMEfBlTZpR/vFK8Hv83tHW9A7707pK+LQiOd6i4J/IvSF9Em+Y6g
Es43WMIVp1DwjnAJ0e8Hj9nIsZg8I8i3aVgHRZU40gGRH57x2M93aNb1EaOCPi05
OlESN+3BYq/eOjg2UbIm3aT9hEa1ep/pA6gsPhGSXr40rvkizv9FEz1/ZSsPhst0
qwS+BtCyFF4oVsx+pBzHcIm0nk7Ew03fVgULa/zf6CC4bPOCGhGEr/mShn6z08x1
BoOPIN/q+s4hKT/4OejB/exrLXJnjoa0qA1q2dlD0vKREG3CStvMLfkHuSsLnHJS
1M4jCM4ezCvmNBMyR2ohWuNiDr3u82h+SCnPeGe4RlLZ/U+N+TwE3Ohgh7hXynab
QVE5TufO1j3CRd/dxYbZf+OaJVizBUDslPR+G4FJezWMrNIwmT7nlYXAhN6bnEIP
8kOzU/8otjzEV2D3myYdc4+I+KSx2yzaYw+3Fhjy/ThKtvNujJTAeHKuq16yvX81
LXOSUOLhZNMdTiqbXi7Xi54zGdYLk3uKEsM32O0C9CF88k99I82u3XRsDMbzsHnf
JYEYN2zgdhN+BkUKvJ3XIADi1EzFYd7r4hcj9yY3wCTG6/g2tc04V16XtPqv2BeV
PSkYySJwwsxavqdENhrU9H79iaDTJmSEM+OaCPwxjlTPYPCCihpZKnvZc4ln8ver
BXHsWeYHBEl53AX0ENO9SpY3e6j8hdLtFkQ4MTEYdX2CiW9Ak+piHcLbuKpRTGZP
Zo38d+oMXIaPlpPGgNx1JiSkBimbyc92SNpOpwD/diGZdiOYyHKddJ841HfldL9F
4chuOKnUy6OYT4gGaEeA0w2qluNsHQkvJiRMoRRRG/XBwyP1oZgnczGw4pdsizBU
SyCPF+ejpYEFodkONHEOJWmKpaDZmz8f7UAjbH5N2cuys0bxCJv6RVKuPPhdxtaj
do3oiEcGghaSjfuEnAuBBg+a21Ja3tZEiQeHlSGUui5YzBwg9nJbSduzAELgiz/1
7csd7L54ZRD3hamzAlwhS/rYUuWqmhRXK7yhiL02iWXiTj8pT47+3N5uft/308O4
qlIBKhP0Ku1cd4fcSxoXEBv4THmaaw64ahxawT21j/BQQ7yCWwUP+l9i7/ktYB40
XXsBY3uqgUTzjUEQvadZyJIkvUXGEcZaxMS6/ndMCoaxku7zcyDip3k6FiDDDMeT
deKF28KhiS7OP7sz0JTDrM30rJRVrRB7ueDzjKxWJYQnLQ+R8ehQwep4AqBHGkF5
l/+HYolunmwHgmwMGWZ8g5TzHnPP0YzuLbDzg5bByhEUTfQfLnk0mZFgYvd27ND5
kBXS9FqW7RL1LRwK8HJEw+bSo4FAdPlOQ4cmTFKzONhIHEy27T5KiHxBJ3SXPL6P
Vb+AnH3RWJ2M+jl/88qzxJmA/RSs4sMmEnmlpMwmBqBUDKX2QyxhZlMdkcLHi3NQ
QiKfbBUeEuWLttr/cZrulE/AyEDDshlJCrcvQlnGN+IagvaOOoZv6OECM9kdmTbn
9tZRh53w6RFud8mn38a7AshVGUuCvKUXo3XYGlHzcnDik1sCuk4hsd3qyhnZvu6d
gugUEvxiR3DsjojYoqRkD0gcYlMt5i453/irdlFKcBnbLMFmtZXM6crgJOZNal5B
liQzq7MWGGa4aRbdxQSd+YfJp1ppdWpmSAWG2hWETuZHdx8e8Jx7Q6In6F7VFd8P
6lxjUmgqBiBs4zzHKUqEfXSOnyJjZboL5drKHb8PPTYXydPLXZPjuGct9WSCwfao
+yAqkmI8PCKUml50sRenijBFQepxo6ehy8API7pM4ASOSikIbu5p2kOgSEAUCRTY
0Wz3ng3M8cnzMfqF+MKPeWNBdnDTF0tHobWmUD4+bO6FNN+KtPtvpHbnRylKCuqr
/Mz3Yxp6OI+qZM+7SPZBkj/vWyc+06JVPoh9p5gpftEZ1I/Hp4g3qRMEMpZ/wTQb
WfC5IPdYl4lEeUh7VYcm9Xuz1EPj4OmI4aWigHF8GlYmyMMo++X7q3Ef6yfVBXn+
0JWHvfuGSPDYLnTt/DW9PLPjs0ng6gfqPGggpiMhRod5SVD/LQsRIo/X0F9gcALX
i5sei8QqTD7Uf9JgZbJsI7dhVRGW821YQzIKgf9aGdNBpgdlN1jdQtPp6RG4Ukwn
ieAr3t41Np3WcQTmTH4wdZGuD65LvcGNmQ5NoVsuWWnQUOHn43svU3TE/onDrKF7
5zdf2514RSbiDvmdoT8SU4wpFaWxqklpAS5pSR0bsaiI8sOMgAolLpDCQcQer9pK
QEgJsXC5OQu9zyhy3nlBdT7W3ElkQWQLS5SW5jWUti2M6e4ifPA81PgygrxVigYN
J/jfyELEv2vjVBbWOR6XNws/tZthH5Fjcv6uJI8ElIsUU5/zaq5gMMTcSjmG8W2h
RnnBvFU1XCioO+Q3Nrl+LgJ1CDuMuZa81z+H/AcwgWTfgMKPT+pmAVCPTrwkkRlE
Ri7ctoR9iI5nYYG+wvpMSvMxqZDtKb46Ztk0Yv3XP6LaqBrUHfqdF6lp2BF2PwcD
sEYf+ZHsGGH+VhnZzbk98QHuVG9QQrRHvwAyWnGu9CldEvzA0NfzKHq6zE6vSlKJ
xHBmr9TBdWEpq1M1djBCcHUbbDr27A5YD2wbvdcQ5YEbRjzPJe+0L2PjGcs8nVqK
ikYtM7bARIR3ElEpvZfDKI7R2zNTkdoKaG5WK9e3p0+xUtyCqHhvNs42tdvGPQBC
h6Frcbe7PpvvoDjS8eRqh2OGcB1+btTirUDHexQDaM4HPUUuzWol3rco3Gyn3Vu5
IJFAHaWJYn8hefl6fwbTkQXc5d5msB/Hmco3xnypuhCYo3zz1O8uXkAL1MNlhy3t
ejqEodt9BvjXXqU6YjpJXIl7Rqwvlib3Sj23Ni1FknoQ8bZxjweuOJUrRZpgvHkB
1J2EPL/Z1NOpEhR97VUkn936pt+ofuzbLcVcQhlFzEB52EroY+GOLQZ2IEOp/dQV
KNA/43zO0Ej0uj1UlkrpBRLPq7Vi9Romq30BYobDgD0kfH+14xvVziqAncOktWUS
mRkp0u3t4gTGpIosTLZVWUJG53I9aJyD1oeECW/wzM0f/6ixyox5KTLJsB6r2FOw
/qWWzFp7RU9o66Mv1QujPyJbWf5Pd5iyzWGWl9dtCPe3WTPE6uli/6gBCsgCMbEY
c8bdavUWc38gtjfoKF5+OMZzmQpm6HasPzpG6SkWYnwAcTLRmRQzLhe2GeRJ8Ymy
8P638jxQe+6EZ7RwgJXoK6JZy32JyTG2iAXv7ZYxRx4CKTQkzbqBbDSc/b05cnmc
KvuGWeS+KdQRUcrvmILfo4gka6yDxSURtzqrxRRU0w/5mlgwev2i1k4g2s/HilT8
GmKs6PaUVQBlsL8bTxf/Jv9iujv9ZRH3VfPjvBxmJ6gIagX3VkeIfuPRU+PqpyQI
wabN9sJlDM0styXExEurz4gJMBLMeQv26uOiVqdRUztUhu2TcqO0Fv/Eo/Ax4/dy
G04u/+2FdLFBVEaPp2ogvfrQ5JpfB88ezoqI22rnufiUgT4LBOkiZCj0Z+BWEM4t
oL2H1RxVAtg4bT6I5mdoHPifrU4C/B1XSjfSVd/vbduJavxW/F0DBxB3dwCMsjZh
SmxbGrTdxw3NrFeZJMGEPx3zQ8WEZmDZnTWHeluj63ZxFJ3n0SUONE7lsgJ81/Q6
WVmm9yUez90JwlRN16fhg1hLE04AqnBOEruyfB8h/BB971nlXqIfX+f4qUxgVuzz
fY9wOGNatqZBaizgVHZCsloFy5uZ2Oa6uawSC20TbmYTHNJUK9EgMpVtbHVoqr4C
5XQaByOeFSpzVJ3J+EtAuuutcIDSxP9lp8qnaNQ3bhjhVd6uxFIzq7OOdUu2hyGB
m7BJI8XZNG8y3c8RrjVKJUafi7hETrCB6jc4vFD/P9mOQXYpRmwMXikPmCoT5O67
2Q4Dl7nRNiXlPnxdy1qt2iKPgsZ8koFgnvI550pH2sIFTRpcijvgSxoluxI3Cfl1
22q/DHt/IzUMNQ2uvhi7hcgEoJMUAMV4w9ENSmUE8RIgeL2350hk1I6HJHEQv7V3
LVKuNSurdA+CRxUBOv7gNYwGnMvoTvtJ6LTbilTqj9pMfTEpRs6hJ6+UxrNyP4J5
MG1J8tJZqnnxkK96lfjKeh9U4NLwzBLRW9Vc0conyzZSMzqpmPJoyXoVDFCA7T/v
13ArxUkPsL6uuqKCf33gtgKBqHDdvP1rtWuyppi27RsC9xHevvQBtyI0IpYVkSIT
Pvc6p0+6YLXhWk1fua47/J18MhM/y3KoTlQGh8dcfWLWhTXwiyE1PVgWixYjzQcf
wNDgOCTLI5KbEtsJX5m2NkU0Eq7osYor1cAff0L0vluZXJFu4xN935y+eLQRb8BE
3WTGhiF0zPYg7REIgOE+z5a4FraCyxMm3k9s/jX4q4b0YaW6H7XN/O1GX0+DrYrJ
BVF+j3zvNgiQPADpiM/xOPUktuy2/ziTVRIE10BnWnAQUk8aIMkWbiPfqcMjC3Oz
reZPOK6ZmB/1XtBiF+8AhXm0jWhKswN0mCmF2DpAuP9zA8eAVVnwH9+l72/YUXUm
kVFU33yV4McEQLE8XpJ8reXvhEDat2s34kSBwDMsI6wAJyFwS0CIicNDRqpBJPmE
lfmlSsUMyXhiBvz1P3KgH3RMKftkyGqa0UdenA86gUcbvmwSNDEbFcbvzLA/ysP4
xotMsRjWF21/BtAYoXdkv3P6jfMFbNX8CwTZ0BYzQ+hnoRA9ODAr9obO/vSLr3no
QO2ZOall7AGjoCTNvxBIwH94HgRnnkBeLBdKIwMrWrcbzzAGdHKR2uxUY/NjrDRW
S/xaZvvBbsJAzd3OLUDDeWtV5jRaHv4hjFJQrnyy8QCSIR5BzzpaqutO6AsvV3pt
BkCm3BhTcqX7UVCE/GTe9u9WpisYvNJnmsYHqrfxD4NHDLqgOlQdUJS7qlb4u7n0
TD7l5Bp/KuJzUSzShWvsNxLXdVHonWaA2h4spexNBovZwspTPcBaFynb8JdDgaP3
18pmUdyx0FWOROrKnVQp4cuypddP2VrNoodoaEr5aeEpGYpT4Mk1e78qXjIAWWgY
5EvxXbC7bzH1JZV+ZIbBZ2xbH7Ux9VEtnO0eU0gUjLCva4QUv7cVuJiphL4KS+uk
HN9BMnBgepcPfxVHR0JWGan60cTG7fuG3g9ewWvK/q09ylvJBPvXYBWXnYnp2L9j
KwDw2+Wlhk23gdAuswHVgiFJEf8uTpmq+KNdEgkEv/EcW5WSqk4l3cdnTlG4LGTC
ooK1AxlktFt6Jt4Zb7+nZt5q4VVrgfLd1sII2q8+Uj8S61jAXsv7kQT81waBPNpm
/aviNiL0QJcIj1QJJBm4MBnnbmXaEHPYKIKvePLD9iYQIs9sLkWzhVxt6zIGMDjR
2SqgNldIrLr+3o+B/wXk+rN5J6Vod5/tgyflorc7d+RFkjTzFrEJyJwlc+7v6dFS
EFLOSqVnxdSU/v/1SuYcTZ/dBVDL7f92285RnWfkIxki1uthtNCzopGvBI+50kzy
V6qESUtlpqKgtJH2NzfGOeNSyl4PZlfIk/pkXQVBYQXZLYfOhPNu46A1uc+yoJ/e
7CZJIi6t38h3toQUu23OhIZdXrILdPpjkjinqT+UBADo3o9MUxdwV1nOJp6D5cXw
SUmzkqyEuV/xV7li7WXaTtBLD9apCX0JJ2vPbQSiqKaAwYGdtL6iuorjgFb0wxsH
XStHhOmhRYAxhCsuygmBZyyVSr85sx6wgtjaGWCCKR4CsN9xFdVJY/imAWvGCXM4
dPirB8g2ML4QCXrouInyLV3YfbEo+R1v0I5AAkDJbQ08S+debOZEj9UihZLc/eRU
89FAJ/LWWGb+04p01zqe7FLpCCNbD70CeR3uUGGiLPrrTLKUxbdB4BH7oEkx+5dY
Jaru6csvlJBo7VwY1gvX0lJ2bQIK7dVbsmMhHoWQsMwjRybsjrCpYp7f0jIvsALJ
lg0VJKeNbVj8w7l2sMTTSVPb+rWCb67E4bVAps7Frp/17A//nCmOnpcXtYpb5H5s
T4+DPo7tDAUW6/krZ7fprOgX71BVkC3KIPevX+IAlOrWpPnuk13ngkxEpd7BhnKs
Mud7tFvbmNZvNcRF4s9QPh44vRd/Rq/lSSbq/cnu6Db2a7iG20CpjPEmHsOMm4eq
uhNyqH+zsdgpW0/LGaAPev80UTfE+LVASmGu6WBbZ52WOWu4X/HM/DWbytbEixba
BlqV4ae/anFYDAEO5WCpmjkgNT+2cu4egO1ZAYd+Tu9rTdQwQm0oUmqy8cT4FeqI
mb/cvdHYBw5aQ0NanN98w+wh6MDn/eBwb40t+MlH9COu52qtbhMLaqmKonrkAIgq
6veMT6aHGrmQOqu+uX6ylOOAx6dIpURgCOwBQ9RKRaTFUtBOmY94Il0DZJZ1fhm2
tBbSDtL62rkCI0xelaru3cnMMm2ApS1JxyPH0xUrtVcFsNk/2J3ngUuYEBErxv60
59ST4nBsNnjJ1LURIBlCMFg+OnLK9oewW1ro1AkHaLjLzGXgb0Nih6R/ZrhfUzhP
/zmApVPiBNU2KNp2+TZVANFVRiEPLc89/+CgXZOErhC7hsfeZuclJE77E5JIYSd0
L+7DKmpV7oBigxnAy54KAW+ioSyiXxjjVsEZfwENQYRHfL5zNCg1g+mEcxfAGmaF
R7NKVfsUBEVD1PYW2N5pACu6Nh+xel247H6JCNzoT6eWZC0QlS/Zs5MIHCFvqP5f
VAZepU9MMsV8KDcw67eXadqsZYmh49JYFb61qDoFzDbMeqcma6m+zx//x6nJd+se
9whjD627A7GF5Z2UCAiXo/1mH9yTSMAW9P0ryocpICx83/ukBDiS/cBTJa5GJvIw
OkzrJMiLobjNHiB7QvHQSQzbXdiRjlQImTR5AHQbkgoxVN6m6w6RHFQyxl/pZD57
TCjRFrQo8uYgXiy/mCOvnkCxbCL9ZgEEdeefgO3DoOQEwzUC3QCutPRXGe7NGbI+
HaIaeIt56vGj3nSgT6NXuXQklfWUL/x6YR/ZYB/AblHErnooWb7w27/smEFyfnvL
zkcWH1pQOFl3e5t1SqnmBcGJvZJXr2e/qLXACuAGoLnIlmGyj92mWJYOLquPUCzJ
9F6rtkwRlkGuDqwp9BuUKygo0GTldiDrpDIaNm5xkU+xbuY3cgOdpBh2L9kLLyUt
oEQhavloQZbs6Ki79Jyy4P7eIzGPkmumullwsEBInDexjLdQQdjnWSC9OAvsgsqp
Aiq6P1/SdZ0MrC3XePiNnekMj0HzRnkLIv3HrvC4+cgH1CjxE/PQ0jlNN+TXG2fT
7159SEXNQgAauky0TvLoRr+My/RqnSj3NAvpl66zrWoNGr1VGmuqblmkt7MgQH4e
C1Aliu29hFBFhgPabSYNdT47YtvMhkZ3t+/o0he2Evqb3ZF2llBUMgzTWYA0xDKB
ByZc04d0d72ur3+UGuymp//WIQPe6jredjYBtdDDnNECh7WIJl9i7FASCLnB2VdP
WcZXmVeNMOA3qDrYku/yTmghLxQvTUdD1Ohpdr9ZNAMR61jxVM4IYX9NuQiwthWl
ghvBXa6YK472bBds9r272ur08D+tJ6F19k4xM92LQ5uQA4oZepqKrIApCUSs1Xsm
0NZczEsYy85IGsieCAjr7yKwfan7s+9hoA84vDXIlJ5G5weH/1EWsU+wl/5sSftH
2OkVdDXp9sn9lxuhU+EaPWz5KXHXdZzmyx+as6PiDddxJ1/qMB7lOBCEsSoVUxIc
fA02lvF7p6bKll2IfmTBNU9Q+gfIRi3RvV+MAiBL6EK49C+GUmP7IyQJIs6lYtw2
222NNGRYY5+SPzr+hy97uq/9wz7ZzhswKefwmVniBobOl5LF5GdkBs5DaIIZ5/LB
TWAoCjhG1N/8NprmLXLs2CVmCKEOLrEVgwrtB5XU+VE+t333ECg2/IdMcp1UNhgf
/I3bIvj0CFfte7yWhP/37ziZAZZfSk18Pqkej9+18nFgrTUQjTsy6s5A2ebJr7qW
jvvvllvjfTdiaKePH49cdM0kl/VVnod3bZSgR2/yPgvQm0QadevYxWd5MRX5JA4G
MBNkazGlIDV3OETp2teqyBeeU/z2bj5qYE2Pln6YmFTAu8SxKuLspcxVVvUGqcVS
dxQl0qn6j0mB5upln/da9Y/sYWBOn8/RvoVC9XR3lqFI2JOkNOBS2yKTW+sq4Ra3
kZI4SRViQGXI3Xxgwb7fZYV7Dg3RFV9IgJEdiDGQ/uEUKkfSE+yOwDsWRGoLD4SG
B0H06/0NWH4UPiOLf8/uOp1TR98wnidUEVeaHvyKXnanlBgh+R1r92gPB6tAE4Ba
D6keak0mc3mC5sai2+RjFzjxXZ8q81ynxjIuhNZ3IQ0j1ShuPNreUhUZ1BKbSSp2
1ethS7FHUy3EzWiS41xHOgYs3wJ3XG3MLYLHYKMwSR9BsQuArZsTQ6EUEOy26bnL
GX8EqcPQijGJaefmKIHF2f/QIijbdc37p26HE8OtHmJjqcNWAaG5SZFaG+wx+IdW
Nxp//X/As425ijLeeS1cKc0Yc306Xt5Dmu7Ns1UXPYsqIiZQkfp589dvc7NaTnbM
6Y+JWOOWApM5DAkDmWMqhIggVVWIhtJROR9lq42pS68NuTpJGQAUDgvRQ5CbW4hR
3ay2Kvxrk+tuDlK6IDBBWAiONbuhPsRRDNWhX5/9NEaYhxS9zfidoVn/SA4+7iS7
2cmQzQxtMjQH3MDH/NMZ6mZpISY9jUUj3+/vyBj47khnqvWwxSYYSGawbbuns8zt
1EbFEaeEezQ7wEAD02Rupp25O4kbhyWNY39+ubqfYXSppjByqVKru42OnicA81n2
EDweNsUJWm/QwJhmx5iNEdVp2YZFlOeIlNf8cqhz7aOJDPFJxO6CScmXD+qYIMVb
FHXm6BLFDYgKs+UVlwa1ujO96DDxjHl39nfAmneserowCT08uI+Bx/jZ+GngnGwg
3+sWf0n5kUqgrUp9dBNwoMPyEsrVVs0h4dGaqxpgNgXvnB+85utgDcWuAviUpish
J//4CUl13qZNd/q8hiUeVw0UBGhmB/7IvsxGLGdoP4Ib7gygusS6HfEfHchp2kSh
drNVWz3IAwWkJ7TMZ2e+gQP6jSa9Jf9YWHWj1phmNDWKMZIrSRztLoJ1vtGbBxnI
mwNVpZ1fwX96F8djbP9m2p9kOK1ksfHJJlRf60axYk0hGbr3Q0QS58+DPWSL6koy
uFD9Wfw8Y1jYkwn2qe3sogzTANna4cwJ91qtJnMq4/pkXNr2lZf24q7bhHXz8cgk
VTyyFLOnGrmxVE1KqxhEJJZYPNAkNN/wYkzo8rX5tHW4NuettCmywtxWAhD5QonW
RhQ+iDYQabAiyhQBGwiI32iIUdkE4wweLVK40lja8h6TUwxyJBVUKnkaKqHFxSLx
joIxihVXNR+S53dU1reNZkfKsdmzUwhYuccvXV4NTQJn/u+eGms6y5g/kfpH7Z/P
Q+WPJBg3+zCDLVg/+Ae2iUWsPZYpyMRYZK2lZeBaJp9NNxgzxn3yB2br1OVnAlPl
oWVWzKJTfL0ssVBGo71ZohEuPZLOwfQ2n5nxvdeXWjji2UP57a+s/cOM89kq1up+
bYW8+YvmZHRPNuql4A0VHc9T7c2HR/fgH3FAfCYj29/DFJ7CKgh6KJM8CtltVJJa
EeisMHZiKhhquL3iORHLbxyGMfhfabTS2THo4knNrG4AD+6pklp1Hnp5Dyqrn+RN
cX9oy/zW7bxPHc+80pDogLZbtYM4+Noddlxoqso9ik+jL6H/cv33f/h2s1T0X0Nr
RfNOLtmVHlE74aWFwyFcnrV4TONWlB+V4pwEMZMxd+etcpEan270BEyYRQm+DyF/
Qlupv7cCYJH9+IVTEw9PA3ZACHb2HvN9XO8io16Fo/IgYRrVkOHeF0Tz86K9ZRcK
bz4vdY+NJGUdYMrb+tFOeZkcCsMDGTp6O4V3xcntd+Es1VEBIt4KneQ/YKNcRm+4
j5E6EYUBeFOtAFhO+4ys6zIIBmVoxkDFEeZ6Npv12zGKnrE6HrnJvROBXHKPJzO0
UaUdQlX5ZeOiL5GC2yGHcCgu1cFBadziLj6owTGE2x3W81OdahghNNSEqoY6NfRY
gjT8DYTI4GKuqYqVWqjNaRROQ/VHlrpH/KuUOLBs0FNAeUyeKKgCmzX50dd5qzoO
VhdoRFyPHaBl6qKDBQdXitk6tG5RHO/80pJHPQJdZN8ppe8CAGQtNyN4xN3YmEKe
4zE6z0r475nQix9QiwZ0fZTTsq2WxC3vH6uOItvZUkvpWIT6QpQMFrmZvst57kK9
TgC0vKiOluyjI8nM5BJ5yVysd0q2ZMQFKqecXPaCXtVDw4Xra9/KTyBVtd6ViLc7
JLcgZSvHF7iycV4dUJrMOHKqfvQ++fqOVevsLWZqIT98hJ82p49kFFisAAThzj+/
sNjHGRG7+l/ir+qEyDtT5115HuFdYbKy3YohlJtnVnTWLNqj2leO4huJcQMC6Iio
NqS7kzvFX8FGm/6MO7k5WajanfgZ+v46dTDZOwTqq6qzYTzWLBLg3/bNIv1pKHta
aPxOfUDRaTvFfQxUNYnzTWZvwWfXFnsjzYHm99RFa3Yz1sv0VFzBuywOb4TptEv8
rFY6QdttEafj28q/Mk85+CpOA5NcZbwrfAK3KSor4VnOkfRYySpgPKKRY17o3EFo
Dr5o5Vs7RNJcGnY/VGHgP1FTj5Mvcfs7BDXARHUAXAh9o3eLfj2WHLxELWakEOrU
dCGG9kp0YZmOc4Fs0rY8UqXpwEAh9iMZ7Z3w6tKGHBTCqVGE8YxL99gbdntDweYu
I/iUBc8UseZUo3fqBGLY4C3kzWtgRIpOh11fqECJOaCD0em2A7YKI7Zr5LrQD6Bw
AESYod6hF1okUD74AETfM4AVS5gdy1XnpPxlubud1HGbeCnUoK54FQ7VFEpQnkwa
O9GZz9aDpAaKMni3uHQ8vr8ACScuqX8KDS6o9oiAns6Qm+T90TZ0krGQ5zQUp8CG
5ulHRTeHCnNeABwwfftjVtHiRU4y3nrmmTYiS8rYZAn/XpspQeWNZ4H37CL+ZrAn
M1OzVrABQrdfmiurtLVrPrkYU4R6AD35fKY/VJql4pX5yO6sa3PCOneNJwSiXzRR
0BHSJuvWuWcbg51DpeKeIvcmQQQJRqD9iHc/SXLmY+vyX7j8eMiMxtWX/9/7HUJo
PNhAAMNsWHCtoKrtH8EQCzIFoaP5yt3tBajgcOoaX5gJVQ/TVUaoV81UiRv0cdg4
UaG8Xd+YQwlxs+hXqlRtvsZUtIcXzTJpssgK+XkWVbAdk978DR9Ttw/VtA3CiuD1
UYifKX/oJJsLCdYhawc0BW8wLMb2eR2gBoZ2yyPZA2j8Up8uTVU5409jb+q146Zc
IoIrMfpG6HqE6kDWSDVGRaVK9rFpM4wB9pBiSvyBywgk/ev82VvrkjHJYpS23CRS
fBAu/+E3TXkPkjUJOnCyj8OIRF4rgRMb9UeYLjvqg2DnYOFTYDyW8DkTG8zhno86
AikYc+sbnuiCsKKBWQJ9yvHYqcLfQ+I7EwMQ/rkUSDINPem8mEXLdKKej76ktmDG
1ShwdSj2/Urz6cSKTIpidihJmW2UyyS3/csASwOi5oIjahdqoM/PRRzpoK5ea7ka
WVOawr/1YcnLIoqLhXJo/icoKirYy99iY0zFUL0T5jHZsFA/P8d012mXS7qQQtHv
JYtwwpoMGLF0RHJ6A5PDMobB0ZO/I3K8EaYPdYVvDbxZoNdyJAOaZn7oa0+8PE9O
xsHYdhp2ZssPjzqKZmRMiRI1/wkfRoNNUuLjo9BLaErlnJkUGb8OrLjWcx0FFaTj
F45XtI2iW2MXnnEsTakIeTElEhLoD6eJRj2Wt+MJfv67pFlcheQ0w2KpYKiHuyIG
HxOLOinQS5Oh5b8P3tmZauPPPqig9vSq0yMb1wr56DOMKlGoShD58FdEf9TxR96O
HdDwUcHGOLSynjmLb6VnQZmvLCg7wNQ3WjpKb2UuK/rZeD7VuwWCFtCwj349rmIX
tzKhBDSLXHq6WrFj92jMTgGa+SVzaOzUO4W3e1zYCzg1/mQgvr/nhag7K6p/hBuQ
tKPnCGBtGlweWfF8iNBFZNZsDSinAcciLRYaB1H+KvddnEvs3pcDz+L/Nk7SFld5
oxRhOVkwaOqS7AIxIQmyllJOCHEloF9HcHvFXnDmtnXPgnFDOJ3XIDSoBatwxCSR
tj3qUK7vDBo8+FuX3wiNaBZNKDYGPWpn0W1zRgkVvrWhc4tJ2Dedzxk01gtpoIW/
Igw5Cf+ZuzDF+G52H0I1fWhE8NY8YSfm1ructG+78hcBdTR5aRSxsPMaSFZJ3WQw
HIvkrw6Rr9VPQarCh25qb7YmQsoOu0KoEKPee7c3I8hG21YAlMgvwwBFneOFXVQk
B+8hZimnj8AFIaui24qhivffneWr3xjgRnKwr5ZaGbDxPxqGF6Q0Ehgyt3XD9Ol0
gYvvOjNp256RHG8mcdWjJdRatDPxCK3IymP4qcr/JIszRHzt4VaQYSLgMajCiiE0
EaPyTReJcpS2b2Vv88Ife6aDZU+jj8dESXRsFcFsw2xgVyYhci/ejpUhZxs3SRsb
lLyI9sEf8IolfBUvuxmG0N65dRpiZ69SjgAO0962Myv+Q62dWFYyzhYbVDphJIul
DQefcv2i14Gt5kAqDLWbO/o7krmFfu26SHFy+FRQ98Bgu1kv3tDPo8jjAfPMLOv2
a5231sbKesf+WRkzqMcl53Hb6aszHlPdWTSNMS97rWISdRzgB2pq2Ko/Rc6kug3Z
V5v/Dw5r/5Jg32iv9vwHr4Rxm5QmESpMCV6HTwotVOfiIuDNbBE0cwbqryLjbwh6
d5e5QMmjzy25iayds9z8lPNMTXVsif7A92Ycyp+xIgU2JI8vCDRWOv2XBCVGpw7P
iqpyDzIMlCkoe3lpC8+xjVW+hjlrsheRckKNg0oRSaZ5SNkRd/S9/oL+GDwfh7Tm
ImNqlF5tO1zGS4dj2vcQu+VSndybtnLFhagdiUY3NHyG3Tz9rDs0RrThq3F0NrBK
H+kLWRXRuTYzpzUJViQh5mnuvaPtkpxGvb9m+piImZbm6qbbwnVNdU1ViHJJ4Ywy
JjgCDGaJmtKCYIx29cZNtoa/E5mGVCaIpUR647lUBe9W2Z/XZBpIA+YPGSvfCLGm
SqU1D+0o5nMJpizsFY3C0Zyestj4FcKwhizd/CIfGTlmatKnEwYpxMqILK8sR/pU
4y8pvi4GVMugeDn+b/84JlpCIzABmEv9ST1DgrA1Kq3oZYqGwNe039qO1y0AGThJ
5oZqlsLr2DokfDtvOJriX8X56/hQ1+jqMRT4tV7/nc/l4kEDWV8RgT43vhkM9vpq
3hSoTQiu6KQbEZjJCG6wQWIM2qLY13vRwHmnWwio57DPw7xSX4nECvUz6v8+OVbc
kaX0V99rz7uQsZOfB5ZddcQOvswBH3LL/diGDROw/miYSy3IdWAxe6O9G/E8Wseb
FQNWwhWcrDzG/+yggXdPy7/zlzZGsJk8YropblVFTh3QuIhnqHErj46E5FJqrebj
DntYlGExpU1RUmvqPJtvcxZvXnA39IRo6o0nI/7fEOL+LIbRb6T0qwWABb/wqsZC
e/VtsTHd4SBY0ICtmliTXVe1WXGtjCIp+mYaIt5j76Zy17UHN3nKM8dvqDaq402t
t7C4jD06VIhv2ygBEYMA75PxImrotnF9D9tQyTNL0E7RStNnxjQydg0I8GYrLMSe
GJEkAORxUCRRP9o+VKYKhCv1Fwo6Bh7AN7UxTg5SST7yywzWJeASa+eyMcxxQMT/
T4N2ZZLerQOTCWgltalGtBlR7QVetNJe8tXMB/bUzvzxtGqa1Mpl/+QOR8C6acSO
qEjO4RWTF3ueCzueXFicQJs+rJ7qn6gIzmMoGl0qfwJCs5sMW8xUbA89pAzh4HJQ
lagedMs/Hy99i1HSOTeLdvXi3JSBUm20BJFArkKw788/Etm/1FSFfMsD4abiOfNf
WN+L8z5Rgq/7QMeg7d7duSdpk7Iqaogz0SQcxXlhwaamG8ZYW0N+8mG4qYKIwb59
KCATxjK+VZrRTDWAMdB0Iip/3WcKENS0hX+k/0wtpFC2D3PeOP/cO6KMk0fg9Uhd
7SxRvR1wbErCHLNLmFbPdJD8MQ/EEFe0bQJqba9JUzFDJZK/oqDTiCWcSUWLwgme
V5B8zp7BEyeY0C6/U/M1NWID2lksB9uOIScGzotQxi5AYyzbc5yK76LoZnKAzmCX
3iDYSL1BdHN1/KC9AtjcaR0xEOnd6LLdvg9oKWbCqpHIRvNmfW+frpHTvN5Dvjgp
A1tnnY4Aae+FRFzAfdRf7stwAPP1wr3tF69zXgR7D4ySKusZTNhQBpamYUPf/yTk
Q0vqmyloMhZuOd3a2lqoXUI6TIuj6grDiVDLMkFyvm9c1a3JmRpxKsjFxUncKeCp
lJGouHRL00laNWMKhT1V8c1KeOXcAeW1YuYzFVvry1JMy0PrNwPsawzgTnc1oeN8
zg2u/XVNOYdmalOQwBtQ7CKTPVTqnzzBi9g5jQjl1jK6ezrnmx1c6zwsDsT92V5O
t5ua4BO7D8Ljs4sFskZyx8loxqX8ciVpI6C1/qgwrirkxBFPsrCFAOSlfatAXLXo
M709TMGbILp1dPw6o8GqeF04TZDOHkRmCuR1JaidVvDRZ5e6HR7tAYUUasMhMrZi
70UbJWMDUOxsAZjeguIshji5XXfvHvF5+mGDErE44axI/7DVjWkW7XVjzj1O5sIh
dJqvY+MEihenXRruv0MFucuEX8EEYoEccyq+5GkbLLU4JvC62fhzzR7WkqKiowqf
rz/IS8Ccf6qe9FsgZWJb2sXiaXqL3f66HIf0uaQR+z+zWZ2W01PTbvUU0XAZdRMt
bFbrKEfGiDuMAKbbhoG7j4mjZovQKbz2LRGjlvlM3Ek/MVggGsOOdFKPg+E3SBji
L11BEOnrlE3vaocG74I4vlyUCI0uuJaYgUYbhPRdeY0gjCEPfdRXCvzh6MKcSjf1
d66w78k+BKQuViNfGBniqb8csdAPlefLKcTuF8SK8DWKjrvwiBJ4N3t5NqdsWMBS
fqY0aPNE9WtJy4tHNRc7Q3sWapF0qo/VFotDgkPB3Be+NhZg+VDaW//J+d6Kxyrp
33UC1Pnq4CEb+mqhzQJZRAePFKm2Ogq9RP64tIBqz5nJQarjLhzgaFA6iXsQK/5e
loy7rTlpYArMsgHjj8AbCsbLt649bzvnI+8t6xvn3BLfx89OZ4hcv3krgNS5JlZD
g3wxwahITQt8R9y+IUjG0DLJcd5V0GMgQI1hVsuwnTadv4tr/zI7pHM59K3lhebw
DEBw7tFhCh8/+4fs3qwI0opSXS82INLT9eWUL4CnLKMrzHCciEA6f2SyYSx/7ozk
GYsd50zEk1hPj2CYIVZ9N4t7h8B0RGnnucH9XaIecFcSxHOkd9tDXgr8qTNo2RYn
PRVpBUwxAEq3Aidec6ERW6N/GeQqSLa9hWeELeTJYGNjYLQsLaFANBqlARzwedda
vNFFTrZnKy699zqxrpE2lc9BJtljgV2tHJz8853HgvJwv5ZsnbRZKS1F0+omjFrL
COrT6v2SuxMS2hZN41XIdUBFl+2wPd9j/09TD6CfkDA5UOUagyxHY1acWQ5PXFih
lUaCz6xgjng49eIIWcVn1qTJqj4Q5YQULs2nHrXpp/0G5MSMgiyMwMLGl+BZgHtb
Q80ardNz9K9JtObPNRF9aiL6JJi+DPdf3r9O+QB696MKuLSekxXfjlPhvU6s4mAF
GvlkVwbCKpam/FGHg0u0K+FS7eNdsKa+dF5iykgCw3yw7DM7mVrc55PggC1jp+nV
J4OxTfZ5xriagLRtP3Zm8InGIJ9Y5YK9fiJPAsjWuVn/nZVyJ5wbpTqzJmnHf4NR
A746QRlW4PvqonM8t6GCSH5o0pOZME/Pcs2GYup+TjbHBLE/mj4fq8A6bJMPFdkg
FbaHqTmtiidFPi+DEHPe+JluKRWhHfuEZcB5cy+zzQMFeLLN+Nqfif4EtCKN9TD3
gblT4IiiJkjYxFg2EYCKMHnvyiSrDcJt56vyCzU3vRbCOhF6U6XS0Ai029ab6JfT
tzMyQFHwnW2ZPsRLyyat6TpcaQWb47Ukqznf8DltK2mgh3G70FIY6TTkAmF9pkuj
MI9tgWWuuARjHVX68NuRokXSmmtaQv31m9iFk4cJShmNpFNYjA/wKzXnSiiNmE8W
p4K5ONELb+NkqTULffVD/OWrwd2PXJkpXcU1sdhS9BWJmUEFzVO4NtBUmlvFzFh9
mnhxJGhCU1+U3WxnNwPU4C3YCV3QeyIaTmPfGuKLvt2fYRfmJFhwB0sr5Lh9S6b+
yGqQ43345bnvWyE/lH4+sMwyWDwwfbX7DndoyX3bA9GmtGck3EeAvGyFevXnCxky
Sl+QpOlAgQJCEKV1kyjx4OxpTvTqX5WOyIjd1PTfwXk8WY2RkHkoSeCqZckEEw4I
FjK+kmYDoAX64ZjeLW6mhx25pPrk/P8LRnLF7bDhCs7piyiqab5S5wNZPZDzHWEC
YCQM9g8zGeCiyrgDl+sZ0h9dY22GNcApBjZsAnVeVaQBfO91PJClZjO3IFceNg37
nBrmbL4C6fRXNoOxrfFX1UvguI+FHKSjv126/Y0tR+EwVYokYRgBnggSYRLCyJoM
stXO5bmfyoTor4+MIxt5dksa9is6kCSvnX+XNGtFw1skT0+EsVwgpFCP2Xl489xt
OAgKzTfSXeJr7iTdSa/qEEDpHsZfY38xTZk/HTRSgYSyJ9Ay6g1Wyp1QnhW8k+6p
YDbR94a7eFRAHuJIDjdVknt1Fqh4iX5YWE14vwiBifbJHyUSz5F5ZY91SKRChzLy
TWud4cVjbdo6mRnk2UcCW2YkxM119u1vmPy+IyCSIFTEw++jwhN8eZIiFgxPsvHG
i0CV/fTMZZZ2hhdmIXsxxntBHdiICVYbyoC3WRVql2TggCk8tWUomNVelPDMQdyw
wxfoDkM9c2gLYviHk77WmQaUcdiRHkTf7YJE9x/TP0nJQ5+SOY3xxwiwyl8dijE7
N3pJwSXAIfD6hCOOWQmtC9PLJK1sfuCAzgsipDLS5ETBSawzTuJtD3Hpx/nMOL5F
SiRAqoCgWJ2AG5xXKc4lmXe3DadvT4y2z3//JEEONfjobsx0OZ5tmHWIiiny71o2
kZFjoA7VnaRHkfzd+7QRPoj7TLgmPnm3IRcv/lh6fHrZF5VQnFQrTfxFP4LAKSe4
J3niwl4DTk5nf/ldprTh31rT5troDMDqWSwo6X/SqHX48UjhypTbzDBW5SktmZ/R
RNEuaWBdfpAwIAvbwzO6gne+eVEqz3ECpNg7SjsSuzYWKIFCXIRhvFuqVauY1BZu
S2SAxaZUOEewbVviiqegjZUyJV3XOSZyaLf6nVHYx1lcrYFMC4ib48VDqIYlujKN
mdTy8wbk7WCl28LV1pjUytXtLx6QyZ5F/NXWuGs13/dZHU6qQ4y3vpWokF8VugnW
3+FqyX5MTfKJzqCvPuaX4vrnEi5Cjb4PieKsExXE+UO3a06IC44IosM8CHY0BrTq
9hnrpn3aKPsRWrPNtndpzUWNjEMJA7h+ft4qrYGckYR0jBMYWc+CynzWDKXw11TT
q1JNTE8XMb82snmnYtj80bvC5GXAvqqImhIcFxXtA5JFiI7pdGybeTnbWuZnbiH5
6EPlC51RLYLF0DUGUKpbytgWsTcKbXBNXs2sK5LMU4gPsXq4RZXkd4kzqGen/vL8
YR4DAFDQ7e9ulMQU8NpkKQdwavJus6CCsYQ4o/I8HYqP/SXQnPhWpY/dzGQvxFXn
lc55U2WeN5kktYw7CiMMD0HYVKtHV7igGALZBQFQSOKN2FsqMfRvro0jqiMMp/cW
DRtUyjCKn4RPJsJ5vhBuZb5Mg0cTet3Ed1lhri+FfhrVI8QevVv00/up9qITdpGG
ggDW3dJmsDAkl8wfL725bDTsotEhS24cUIJiZl4NGEOldB71JxwqX2PS69VncSfn
md/QZ+EVHSuGyeWXbSjKXx8rNYg5qc7asoj2MjZt0PMYK48L392kdNHGb2MRKub7
CvelBWPsB8jasAk7teed8mXGSnbwgAsOQExvHDZ/9TPwJdHI5YB2K+yL856xcyJq
Aq+FrJg8g4zD5pjfO4awrdXfqc+lZW0Xc7RQvKBQ2Dz279EQ05EbmkNlzILi2rPw
iZMrSN2L5EWIVLiJovRLaLt0PUp451LBWWCsdcvCG2zc5lVXIM8ZiD8xVt+zthGM
n9sIJGkP9cRBQJQOOmdAwtwjN7iIfKICQrENIwaSbWixMQQRtpOjPZBrhbMbaHK8
vPFKa+r8TxjCsKvw04bPk2X/0MvRyQi89Tsqb0WmkejuHPd1ooLTCekIVQFwpGB0
qdM6iibeikFRwXhZ1L5ny44t9tTs3J/d/Kd2W9rMhNFVO7JoKC+kKF5mErShHzF3
CAZBgr2gWNsZYSVQdKmQXxptlG9gXD78BKdsHXjnrL0N68qPIth/WlagEknPR+Oe
cMJOy3XgAumtO0TIsnZWiS6jfmyILs9ulHOEKlVpcu55IggTSanFvDRMYCMHF2ph
97jLBg6UK9aDGJYz5f9BR/OpgqE8fKIHb0bEP0H5mufgeIUtjpciXXDhRfOcMJRw
RN6T9sMwDLiJey1NZo1JoDPrjWacRePO/FfUaV9obxHkrDii9oOfNpXTykaHp6Yu
lGpnObPeTeRdWZFKJNIM44jlwMDA330LJDFIEKFxFT40Gx+aymruVeuyE/5Yi27t
tKNhO7TRN6iyTvSPLfuhLvKmvQ8FqoBODafVDVtpkch2Hulz7wuNndBnYTDRFz8f
8E9O9w74HWooHrLusfxdRz/vWXtCftrVrC0+fYcnivf6buvX/fS94UgMVaQpYbnR
1Kv8hMF1Y6S6QAbz8eQ1vg+ZviaV8Lx8YwtaaMYhmLkKTZYbb2SLrSioefb2YN+l
jxcZ6dPLRiMfeDI6UDgLgxOaekiQVpYGPWeXl35TeQ2pxnCURlsoX0VmZPeMAz7E
KtC1K2CKsGXBod2pdcY969AQyeYlXAFA6r989owYcAdj2hLh206b9S8ZdYZdz93f
7uDunmwf4kt4IldglY5QdJ2tmM/osQFFiV88zsKkpNFi40ueEEWEWlfbGK/CvnNe
X9BKBZbeRHfIGx7bwUCzwmrOkqPsTlV8Vr78Ccz3pYvmEJ5OZRooYCB6hXdtMitz
USy462QH+7xkpG4Hf4XIpUCUYLZMCfN53FKsIwFZMjTkUUd+UvkwSBIHeLQ5ne7F
QQwpOv9eWjzfNNZNkU1XCbxW9GK3uZpVyCxqSWMC+IyzO7hDlXZTNEV0TNWGoZqi
c8qBBI7FJjQtGukRySRkHkSoxJ3dzNPwyC4cTGB2HhvzI24uMkeG6MiyjCCJNDg2
J9X5dBEKBu+c6ZQyOCM9kLQU3TrlQWYLHzMbOmKy/J7cSYUrwmCI3un01JEVtkSx
E5t1PdrLqtyhXk6xpUfHNtj0U1y9oGCdLQYCfx5w97HKnha3ssKqXokVj04YbNm/
ELYYilmtoi1YmlQKiIAe0FtUTrh+wdzJq7ANR7mosjR++AxgfxRSMPeqT9S0emvq
YxIs06BWlCqlmWSCQKs13GT73kmSEbCeSOvdWnTlWp0YzXcx/VgzI3wQUfI6Qxso
OxbncrKWw8apubCTRBYgg5xuPR6iVFCEhikjR4FCCYlF8bsyK2TGQCD9oM9hRrQw
YjzblPM0Yk/RyASXwA8OXaff3dsIeJsNnlh+sn0/zZT/0ID0Osd+VVwufmZjai6v
W6V3lqXphd6ovdKyX+rt2t+hPskpTLQMAYK6790meeEzHOb89GdZJzO+rsvqcUXP
05bGWY0mSxuieRFYzG/C+XTcMD8ks9WtP9tNYBUwKwSUgoasK78PKrvutsXRyNRC
3oLqu/hS4o9BZbGK+gGs5LETFApFBBLaSbZe4U8AHijFlSiN849MMEn5HZLl2tG0
xTuHlZgq+lSSaNltR3SYVSzs4SQdKzNy72xisFxvHWgXb2KUCxprggLsrTcktJIT
P+vspPTK2JDe1tt9YMNuMV9B6Shd8AinyCb+g5IX1BOjB8NIDYevdGcVLwtWZbUm
tqh3232FLGHARGfmpCEH4GiJ0l9SFEA1DKI1PlXKo7zcm1RHvpogoZOmwXE3xjHG
otv4SWgN98BlprgCM+w+KePxe26jkk7BNkpdSHCEua1/7fK2Sg6nw9fx9SdrRCvM
R5RTx70HmUxmlamGwKGjaH8cQoAg4Vr1wfHqiaRPUKAh0MgceNsVtc0EU5KMXeo2
Iy1YwxrTYlPuZm5MN97DMfuL8YJRmm2FkhXR5zy0oBAxnTpONsJoZPGqYvcrk0iT
6ksL6yGm5uHJajkR2aGtlpPZfN+AB4zigd2UGVYoRMh0DS2SLpofxgiCPCZQkG9M
kLE1q7iBNnigEy6VfaPKMZYaUOBWFiXJVW89MI7/bojr23VfoLM7xkmj2hDXY09X
l/LjT2TU34tokyBn/Wq9EBkf9wOKff6Uq7tXctW5y6SEgEhyiMUmaq1zKUzVa3pb
e+5L1z+s9DxOeBzB3wlHb/W2RldRdWD4ltU8lFOeo4TNg8gAze1mUvq0eG3yDEhJ
GEOayKnbmK4N1zsjvLix17DM5pbDnFfHDxtWx5ymYBAdX8IYzAVAEBdWaH3Ve+77
MwR7qMWN6BzfDrbbk6Jnm7RAk2G8tr+M8W0yxS4rCIQsHarzFOfvXXjydbr0B2+5
OgIHEMZRMla36VnLE+YRmKeFSAhovqNf9r0WfIjzHi+aAViOtP3UEt7ix41B6Wxh
N+gfc3rMi9imoHmzbxmEJGKebPtLm23YUSfZoti6Dvvhv0lpMApql9uNYH0JwsH6
JUs2VCv2dxeAwgiZ6/ZwvlbmvldcKqHjqJU1bKeM2YjzEi+iXRbKWmqDFfEeyRyt
shPKXYMzbUNCnH3/h3VZt5KVXmRo+vXbCOWmaKv2Zp20q8gxWqI3XSTFvKtJrJUG
YyN2zuGyBgoRzoSN88c8gctb0JiTtGnRooOY2yTI25Gx48AnFCej6S16iIL0Gb5g
JQYFKIhP3hvJ1FX3UN5FXwWgcAaLgaUGILdyex8egJPjA7m4KgE+7WyAauApUhfj
zdj7n0m/52yW126OJjmGJSf0hrwaXYquTmharCFq8lRkkwxMoV5GJ8DkY63r9G4j
hUYKpGADcrHDDHLxhUfelQZZfVc8Xz213+RVE7ancaA6JYvtp0IuoykrM4C9IVLk
iaff+GFPnFyFIUFAid9OGaxIYBk1gbph4fuo5lIhxlnXj/vb2oCksaKuT+YAwJzo
r/DgzvEUIBa7SPy32b6EUlDMvjriaMkNxyKeXX+N3UWH1TDEGFgHZHVmv+FZXMgW
rZH9aFCLoobMjLcQfHrq4yP/iphSOvsodJWXcDCL5oinzabJ4fRIFxcKOTCkdVgN
7eCSUoqxuN7mkrB5K95kqCvbTyXLMHEeg+OVs17h+7b8ICzsEBzRwIUUYUmUhjLU
oOgtzziG+CJJHuG9QcuioKQVZmBpceUU3++VrOEawtGT8RttXqS38wTwA/Ua0NeH
y5VYdFjnNcmfUDvbNwDn/bkZQKa56c1RDSc7ExTDlfW/Sy8iOSCy8qccfym0OTGt
nYMVNXSgJwkl8YG9RyMyZMkcojW0vg9n4QZbF5/ch90avYZL+HsyLjrWeuUhLIft
+NyLQCxpe8JGagRm1ridbWksu4bNTLIoDvcY4i66f1FyMZAtiTP5LJ3drRzg/nOg
CXQdwgZvvAtSgd3NL50r/GEwbRDp3ah+fdsoBMtpV73XX3sVKgVJSsdnczSO4dqr
ma7nvUncQWbI3xSuV+BrqaqvexEddQCL877px1mkDwQSyakAAzwz8av9xscxaWdW
ELRO9XnB0PPBGqpX02In5LKAwBGu2+EaM5X8NUZPLJ8IfAOkLxpNumJ6o3HOd8YO
pRs7gkoSqSwIUMwyNjiiWhMOVkNchweVS6A/AUAIHtv+UzB2qUTIRcNcgAwnRVHL
VGB1dxP8TNR/HbqDr9Hoe0/Qk6VenuRHXF2/uOHBGxZWuqk5l/0JwmrVNqZ6Aa4A
zvTPulVp5HhZ3DabsL9BX3+zjGgd3xBisGD6dHCbLs04cpfieSS/gtNi7lAFL3mS
Q6YQ2aih4wsO0fvYmhTgOO8ffBVppzqXIX2EkR93QpuXooJMYbEX/Ii/lIqy1twI
yLV/2AYQoEJJbaLU5iUR3Exrm047sjh2YFSJ3qyXT5z7Cnj19Rj2wC2JF+LXsOqi
N364KRhG/m3wvFNd8cx79pTkbv3s6/6942GI4ohl3l5KmZKgOWsUp6bkcEivRc77
mpHKgOZ9JNwQuuPgW/LotVik4RrtqZpGEHii0AYtQoruyP8E1bghqaDMzYZWjrpA
Hhlxh3eqgApxiXMj3TATnZWIAkWudko8e/2RMQzMFiSK1xCIZCoNsHTo03BsLaEL
9UIbC0vsHFd3FPqZscOEXBTTQ5kJoLQEwNdzp8CP2XD+oHIlYinVSGIORm6sw0bF
+J2KpAiqtotIBvq1/sbwUDs9U2CTX2tRrOG5p/jHqUknjn9/XwHgAeM2r3sHMf3r
56V+KgT7Dfjp27tITN8TfL7hmvrkvHtqCZYybBWyhN869e2CJJrerDzWaraybSsh
Ai3uQcRxt+cYwrD00CYAnOfQSLlgZNNhDdsF57H2ScP7fAfWb8815H/J1xlSam5H
TQuFXpy0LVQGiGZ4i/3mDRZcVrEjs2A+ra/++WVJ5ZINe753xi+E/O3ZjaVnmNPW
h8AYWsvtMPqKsPgOm/tl0O4LpqizQoGzOE+pn2Lp1EMy5USLYZnsBp/fpwSaxbsK
8nPl64SDN7epRsQFP2ij5B//y7xUYcge+j2kADHgy5GT9Gv1KewCI/Bh5quSz42z
Sah/pkxQfetjsqJpPGX2sGnE9sWdqiZMJvx+O4kpoavRtfe6B4MpJ2HosP1LizNf
uS3oqA/VXxCW2NTe4M9kBTCi2qYNUR69K6H8QmBLCQnFvbhsxiUuYWiKNpYe8uWe
XFK3mEt8pDekQF1tWmGFxtMjAbgruOdu4g0F+bFMvRC7hHkPomeGKH3YD1K19xWT
9WCQjshjHeW6A2gDcgPmAkKcaLBhrh9P79I+KJLkiTHAa3NjjoNLPcpULcpu23GR
1CnLno5TChxb77XrhTu6V1CsoWP1ATbr9xefHPc2gH4rYVphr5GeFF5NubVhnlZf
+X8cns7DzUhZ2/jBlG+gzrFfLoRIIKxcUEVVZrzkyE+tGMPD3LDyVMQskb3dCJYh
oIQNqtQ5gJrsXFEDaY1FNE0f/cSnioAZS608QvjDPSEKj3szyXR9Lpv1/M+siq3i
JXYwH7gY2t2iNGV3Gzx1EDVtiWaZX2Lb8mTuFOKdtT3lKb0yDf9aEgkQCnSLOcZx
N6oZMHvlXDvbHMzl5CbmSlcprpOSNZuBByewdtTlQe7xnb8X9rWmVPR8Dc7mOyRK
S5n2LySaZ0V15MuyUvEAaxBqAjBeSQkQ9h2CfOhjD5aLGW8qKkyCUPAnMbYwRJ3N
RtXIknUcs3sPzSLfAA3+NT6AN5WPacItZau9BNnQOt0tYvqIzuba57WE0jNX8RGx
520cw5Qeu+hPs6jCV/SWl94RrDzu1+D4JkLXkZa/z0231XNtwANgsA607/duT4kc
gFhz0wb0Yus0G7mNUkkA1jS+QilAk5Avt5kjVdkRT7bPf8wTmulj/4I1GlW+KRmE
5PIwjmHIeD7dzTt+hcDiAkk3UqTOOQe4B999HecYu5w3+daFGJr1unxaUdhmdkr/
beXF1/6ofEnQJK9w6554r6y52zb0e7vSej/tfdJ4ZWPfv0aGCd6qSOMjndoYIyG/
t7yqCtKtQ/Zage/P38NUZ19IASo18Mfot1Ejf3gtmPZNwV3m4AKfsD3GygG6EUdP
WwJMjdyxPSStU7H4d7I0AxmJCheGO+pS99CLkTEC0yNFHP8DLFubAhEsBdAQyhwq
5e9o0bc8JCUAZ3CZQIlgdNVP1azHYE7K+Be/CUlrjYpSABgWBUzVgWY7dEDWTs3V
q1pfK6GVP4spqc09Zu6ehs+XbfLqyYcvqfPEEYeGUjAfmjrc+ewUAbGkMubo+Kkk
+Cg0YNXi1tSuvWe/za1HeERe9SVCXYZVcykFOy6o6CLrJF8T4DkAahW9hyRSATDR
wD2PYuvrcmHoEp4Ljd2J7dGjTvaaBFKykDgiQcSoNnBQ0OCLYMYlq9Rkvcz5GJdw
qcqg/bLGV2PdfESiQ2wtr3AId1DhIfefRWlDyjPI4V/g2LEocqeoEqwrnxbH1FxE
QvWLf3I7zeBTXLMtMzZDtcefHtrxXC/FjTOsDhorPOwrSLSOi/xJuTFgs83lKZaI
P8gRhQ07cJBzxsBTgCDaiCRVb6E6iOCA1VIJRuYsSqRaLIgRYfPSTFh42bXS7h6Q
8oFQkIQPwOdzHf29vI+G6uEvE1dp66rEymlGjChajygCbAYTKGkawG0soM9CY5Ik
gZiT/+XljKhUk9ovEN4S26wb8r3vG8bIVk3dGRDfJqF+dAW/N82wrGUYPOs/G0rB
KLOgx746sYQwvlWEmI23OS6x8IncpMMimOJY+L0hVdvV2i0uHnhNUpm4+N4FQBSG
4+osg7rmhvQG7OF3uIlPiWz0v6SJ4Za8vXzLZ3IKwm21h/KA9KGcrU8/xVsQB4OA
pjq8baRPJdDFOaWcBBd0up47lu8y594v2F/aHbrn6bG2qhjTFYTfYpuai3dkgsh6
ItpurKPQ+1t7NFhONh6WbiIPQR5k1gPkR+409F3pxCGEGoO1rqPm4F6S/YDDW1RP
2FM1ulRKYIQIiJoNA4a+eCTsiuE5yEp/Ugw/0IVuR/gr33zzFLlTkNVO35Wsy74K
2VbT3W24SMPHfoXCr0aBpXBS2A05EpuO4UsW2OO2NPF25GqY0Zx7X8XFX8KrzaSu
HTSg66rZ+WG71VeBo/Pri8dWT0Bxa/mU7eKuNz8SknB8yCkh0YnvWp/NYZMAnEKe
xZI4QlpnIZbiDeT2yRUTGfuBGef7QK2B5JcmbHVM6hOl9tZaDzDeK0D1bDeAygyA
WXX6WRvf2G5SzCCvU5gOsJRXNAd4INfkRlhxexP0Tms9dj65RmQB6Dr9VPsPwhZ8
f36qYwvA/Q+tPB3fKslqP8B5zEHpOjiw8pApvsSqKRGHVz9Brz8ShtNjl/VCvhtw
kzuVX1lNB6eRb6pI1HbbwQArzqZZ/AfuDsG3oqEDBVXDxtfUtjEvNow2pzDKe/KJ
uHYccthwxKtqWM0QVxAWiCeBg2qiyz+WxPnK3CnHsIr47Agt+ehXBTeXN8SY6Phd
Ce/+t7cEiHphTICIvbO9Xf13XYJmr+oYrn79Yr84NVvxR5c53tledQsyN+Ie9DGj
OTvwrjT39vlu6ou5aDsSfHyuIdMpQgqMnP2G7jywxmFbE7s9DXDPrZZ5FEwM1hXZ
nPpb89MFkdv5K02zOcfyLl4IRwGvHqfDrFdaTRVRS0kmIYp8x/+pGXR0Wcdb5p1D
wLM9nYGD9VnY8zE6tHHAdqgVVr29xcRTQkzsV5mVKmtsPP8MMYCV6i1xTk6qiwAO
Hmieyx36oidbhSk9iHBN1UdZPHgOCUZdyfiZAaNGJGLIIZxyhFrh6udDc9sIUpIN
kErsN6RV1FrNm0+dmzvwLHU/dKdp1aUp53L7dITGoeUrde9bYGiS/wibRWkgWT/T
FZWzMw35kJwGjDVAIGsbvGtnuNEJS1X4MAVG3ReSSAbjlJIGDYKe3mifjfmKX6Ao
UuYlNSdlWRNjUd/hzbfsKtpmcD+lr7O9rqGdavxM9m465sz54n2D+9MLfPLaWMfS
Azn7nfcCk8IYru3rLhqcfITRrSwscsIy7nafNLkx1lQGLeaY+oDQqsCp5G57rNOA
ag5KfJ8Uc3BK1hAMpO03q3BxBvaissAhya43bEBaobnfNUcbcjhhLY3iae+2bJkK
mExCTZUFiCuKpw8i/Rg71hkY9kVNqOG96s0EdXU8MEjUzSQ29tOIDuiPh+jE8JLm
aGwwq2WE3KRRLFW4RuzQ62Oh9Zcyy77jtmXjA6HD35/+tIjADj+6Ii7jcY5wP8W5
1t4CwGTgWBa2BSoqdO6jTmNkAhvkv8lLSAsJQNHYXY2zqysiHM3oL+7qFYCQabSI
K8xyxTIKhQHHDGVXYfcJt3/BNTzBn0RgZah2GHrUbIaI4wL44bw4l6tbyrACCN6A
BgglmmZiAItf/56CRd+/dn8vTa+lV9VqZ0H7ENQgGgXmdBeu4VaIiTOdFRpCKCZ5
BKPx5/8wIzQOlW2c69AZ0N6lptlixy5v1aady6IoHsyeYuzp3qH7LHaSR2su8Zuq
3NTQGSjXeaS45iAHvST2Qje1USWOg6LCbIysV9TvMvFD8D1Hq+4aqDOrsd5cmbYy
tIfIX0zlQwgseZZKiesE5sa4QbI14MRKKeEc4EVBV75a0S9jW5v8dBHRi4NwhKu1
7PAbNtSr9HY9OSjBcv2ZFgll7UiZ1e6cmhrCploxlCEMwhzxYN12xUaFv2OP14ou
e4elsqCx3Pq5AVx2fXH0/To9K7sF9iL+p8GG3mndnebvUW3WDA3LwdMk3fwGH60f
KDaDvp8bFmRDckIxgLy+I5p+sR31JxrYpkNPg9vTNtUguKytORCbnSZGRsQVo9Qi
/OBpoYmEhZ4KY/R9QKJI1p6qb7ouejQ3dnO/fGjh1pWm3//JacD4nu4Dv1bqaIWn
w2lZ6WRZMs8sbPbD/5QrV/soZKFb4NHkIqWPTJO8TJBkGPcKG8GPH4Lef0b/mBHv
AWl/YGnGKioTsqmJE88hXwa+WYANBNJ1tfC31bTW3aO6pLsy/45BsjbZ7e/Dv1+3
N4g/1g4HI7wPKhWdhtUaAqcSHR97Lr9kv4ng7OBuLGQ9y5EfUWJRlL+SR2h8aKHd
YAPsE1fVzQpVeIkPaHnPAnuiIWiPwrS7qaXWF97XNgDYdcQ+0YfB+AOi5LEBrsc2
ZtQ2ArcKVY7znNNOOm88Fi0FFruKp8wChUYQktN1sRpWg/39u9caLgktDg7bdVOm
Bo5lU2H/Nr91Z8XWVSCpZOuKa6Tt85GiiKNyouEIwd2XKdFPbDFcnpC6RYorYL/v
goumVGjZsHL6jJscNIWmqepbIlZBCzucQEECpsSZnLJbRBRkamnymYztczu5E6nI
oyNflq458NhtBswoAqXcT1UUdrvddfPl5F3efkrRDM45fHVj6d2Iki7ERpx1+5ZQ
hhOWPXwbBBuUmtCY5lRtgxy5sW3aiLgqH4hz4Mo+DX9n4aat9QsRFz1Ng+c/ffO1
xJ29eOPIvXPen7ujbkQTA82luzXfWx7z1qj63gVvbt8xfX4A5obdIO486zYwHx2m
12HP2JIRVqsRV3kQcVVtJdr8LbLklrA9+i/0oja9LXnT2HqqDuVPfDrrTYaKEPHh
slj05RrzeRKVNL0N7gfVOe7vI0+QTcNIxxooqBffxUCoiRTENb5FOafsGVRrN44Y
IjIm1dnsfSP+VyoU70XWUaI/sxy7SbH51fPVYPwbhnjCLmqiGxM6IRdEF2AfuGeh
8gtjXBGrF2XAV+rrO7qysNhObPUqM9sxmtlyHX3XHrmtlYlbvNpcSiylzhtq9DGs
kCGqJDRGfCZ70AAk5g+EqGx7Ww0X9XD7XptEQ1xh/Sp5nnWFeAH6WxOFHiuOzXKS
TD4ecnyTcbvB8rOE1YC/vj2EkD9vvxE2O9ADodQY5PVB5AMbIMhOTh3VlDnutknY
Tor6YJGEHt6bdjsqAT6fZ6IdgMGrJ35Ln+uf1u7ioJEUyGVngDYP0pmhro5/wC1D
AAvn/qBL5+oShu8AVnJt3y1aI60746jK07QImDYSQkvaXs+WHmehPob3Zb3UcJ02
8xTEoM+KU5yxJlgR+kuzkQlyYUvauvcJJPXJqP0JSvTHbwW19GjPgo14K06JVYTH
112QJLnG92tdOqDxFwYdFcp/IofN/mB+V9qzdqZVO3q8AHmQg04JanN5h4XQJ8Zl
4W3jilVWzXNNDLc2VR48Kp1knFFPMJ4j5HPUcrQkh7/YoXWy18OUhL+oHkzoqC+P
IbgUbBOKqHry8qNtTeGqnYeYXrqZMrYsHnbhvGPhml4+exSUmWfkuFseOWBV51jC
HZrFw/2/4/hyJzoFeVgBIvpi00ffLeVjKV87gXBNW2tmWsb+mjXagt+xcibtyx3l
R0ANMZYuyqk0DYpA56W61BooveMKU/0K/6VlksyV7cjUomRlGdvK7P1PJuoImzc3
cTYZDrtYXIsOdaRMo2fDfqWZOa8taNlJ8MUCPFd71a3Mw83HtM7LlhAHekAsPuw9
rqcQIOvJqNXlo5N/SluXI43aSJn60HT54PGQSUHSzkv8MbMV0VJWgPWw9Vs4cRhw
YFeZkE8rzTnAH3YI2FmXJ0XQ7eVPxN8LMSvKyhEwMTVdeLk3DYRMqpsMry9HJCng
wYSJQh9FLo3mhxQThOGKpNknFoMT+iIoZmnE7y4u+cgg7/JieNIrORrdPZ0jaN30
l26tqiuDuIG43aNdXG118gRMK7Gp7vW0TPqpWaR6ePdyfUJNEIzq2sXwpzi+oAp6
mHGq6F0bG0SiGnNbf9N1veH6QJ+v+etyjQRw38D1XraNQme4zNvWkKXXP5dEIlWu
23/28ObXNE/kKYJOuINkhlzwv8zcTduevUZ18EUuPXfxAJcG6HIhA1FCOa6ceE07
32LqCq6On9ylCpGg12ZQR5tTKIqPkenCI8zoNbdso/1NBLjLgdVpBa8xA360NV0P
ixQZQTM/i+Pc5KSdzn+rXt1gyaOibYJonfqOONQt7AVdktGIkYj0HS2jwoOL/pfy
ivMtauvkw/57PtWN3d8KMAAgCTkpvevVirkAdbcje1DnKzWpkr/srkTl9lhNIo7j
RaZBdc/szNGy4dEONGV3uorsWZHtBYGk4pLsEucYmh7BroaYOx4o964u6EIbr8Aa
QRt4z6zEcRFddW/d9Lc/RVQ0WK8ARr78cpms889UYfTxBVaTGr79MTgJRR40U20w
DbNQKmE+pvzNR8H3oP3xPGYaRpe4mleGNVz/zK0Wck44bIVQa1IJ5Q37CAKKAbXB
YtqWfMsApK+mxUkMB3DBmUvwUuT8GB0jRzlqQ7lFJas+kIV7Wc5y9Pq8dduRPpOY
VOfCgjjUlN81Emt7NRTuHzFi1lIhw/nAMv7C+Vj5qFU/YCaDx2onlK3ht6lJU7qA
xECbd8o2v1SBvcdRkWU1Rx7UkCDxDOYFpqLqxOLkBVvg+wB/lAmBI+MVN/VHzdLn
As4X86f1XlIyJRlKpy+KaFAJO9OqovPfphB7Py3XtxvXSe6juMUGLA4pUk2KzFQR
SMQS34rwEQehIuWJgAwYrRQ6YCC9RXN2WRfM0q20serT73q2+uGZESnhjoiOUAys
zBCXSouEkY1puT0RZGuDdGYk71TtCClSc11c2ZZ/2FdRUn1ho7ZAyqG7IYO2Q7bH
K21VsiqSJu+aKiWi0LVdc06EUWlr1u750PZY8UZ0X8EzgjILe0BHp/o3EP1YBIa0
FVN1R9AZUwzUxK0C5OzXMdHCi0iIL51uqh6WpOYpED/uT+0AHaTmOI9GOGm7OR4Z
2z6eyN2lRVikQzLBf5BaFsm9WNeObCP/oZ8X7f5czR5Ju9xtXfr4+n4dGRmLpI0p
Mbudnv6r+LPFeTG7V0LeNFgttD+25XRJT240iM39Btixu7T2BWnvb4mwilMun2Zj
DtxVxM5cHAC0a6OyV5vMZ4gpksWBlUQzYGSvXEm4Iyo5tVpI3uQ6ayDQulUVSTlI
u5fOXsb15xF5Kg2gv9sW8PJ70t/5iECtjvZon4yYtfZfzOeyGLk8Erdu9O4qXZhn
gEd4cPjFtpqYmFvVzjoCUE1e9U0X0WEe0FOg2qk7JsQP9ITmsc6TYqafYu/sxbmR
Bx8WMQbxlGVJ+mLGBc+pU1OgYBresD0iey9xpdjJnK17t1mffGoinXavWT5EyaSJ
w6VJh0EAjxB/vas9zd2xyLrIgLPfw4fv3ggQmq988RQfr9WM8bg3tSbZE5eCHFkA
L1cPRSdt8Nsjv4WHbnrGjoS27tUDnaibmcxdXUU7ItgTQMVXARjedj/iZA+4tB++
GT8UPLWIodzEJkE3PpICjqkiJKvfEcFOgNc4KDroMG3Hr2lWOeAGUWePDUNnRgeU
GCaRF6tWRIifjfCqgU68jZAnUSWwYGtirySUB82J3/DPhugiDGTv2vFKJA/f+KDZ
LZi48rm6lVw5xIIqtP2KTJRR6mpts8M90jCrNGV1N06u6sX+hpUcmG+hk4zjXjS8
udThpwRqf9+cx2plIRfcAvhKd2Uak0ZPSlF4/DyNjgWNfKQopjw+5vP9f9Oe3vTY
6iiTr9v3ibWLGjNSTLEp2yRrwuKTOrRc/XgxT/vnrUJYHsQC7nyTPHy2LmWEQb50
/XYV/CH2LUbne/ZvinH9Y1cZjVkxFfAkDKAiAe7hpwEVzuAF4BqJDAoIn3eUAR18
wiTEbjFNagUrQtbJqZ0HvOGWofijbbEVcCamgzhHbM+BSSHdQafaSpE1kObeTDWL
c1ieyJTVsqF3gS4Kgph+IUL+ObeulI6pxBnueWMdwz47OTxRQBZ4dDZEP6D6xNpC
HX9800bl7ISFVKx5/r72BDi1fafWeCz8mdXk/SIjLr9fpsrGaRwIIZbVCCmDZPGE
awk6n8OEAp66yWo8eYCM4HKd/lW65TJXHFYe2ICJPKqAwQYg69q6pmry/k9Dley2
mObf+q2ZxnU5iqZNEX+R5RsueQu1KYb28mwccfmZ4xPBXbtQcF8pmDm0P7yAP2bO
2o+mofnsrEgFgbXLreQnO3J3pV35GD84q9ftyI5OAI32HRrhdkyqmYpGcaibBUYu
rRPIDoxHByGJMYGf8yS3R5A+tM2UmdHdIbvU3WbBuMEwrtdeZVcOmVFsVEuuD+U1
bj1OKwHP7xsgST76JmvC98VHCX7zpJxAumxDO7JKEy76wfIQa7Cp1jpKRtsDeP28
K1aOfZ4X3T+tyGwfu3gS1LO5Bxdmr4c+1H1p6sRk38Wsx09L+0+OK20RIJpyn3dI
nB4bWwBr5IOH1Kcovu4mGicnoqnKNS1+0znQ0LeQs5rWjnVBH0SlKooQSQZV9Qxt
FO7zA875h79U3tAzXP3Cwc7X1oC2BESrgx6nBgRu4HNL5LI+GP5gdROZBY0Ay/Vj
PWkmbSqVyRgsNz4OJXAj14BRsn3MW242tgCUZWMdzbxB4d9Bm1ieapITaiAJ0Ua9
6a9Z2PeCZbARcIyx0C36JS0sLg7+6X1vaMKRBChKTWPavW8FAuZOmT2cfttGif0+
P+41zh+pDwONSU8d65bzBSyo3UCZbPxFGzsiKkpYat07JaNl74REov5TAX/S7Gne
VZDupoDpvkbl51Hw0FGQBvEoiZO6Ii75CI71W+ijG3BKmYLYnf5mbggP0WLMWy6O
Nm9esBw7SJJcQkqw2T/0ugX+DTa3kwKCcRqN8uC5kUAQA8dEQyaf+GRd/6+Ount4
dQ/tYM8iUZ9wJ/9d0DF8y+xdAvBfz7JpvZswRMcIjnZ6wND63B7bfOcaaMvoCRfz
acOgUyCQc4N9yXajJzzP/b3u1SG+GIUdOGF1CpXhzV+oQlm8ZeRYVM8G5/fQUfNA
2RpTSGAt0g9qeqeKoG9TjY9IGwEKi8wXwDS77gzAYlTYobFkBw2Of3BPJFRhgbjN
dedH2JkatB9l4HtF6qTdywgzrqST6u4JdiKeunsZgQPcw+uf/zwl3gJ2/xbv5L7A
Df6dKbN/m1FkV2nCL37k2ecQITpumOyh3sFvxgIlsce/cXda1xwbo81I2t/en7nW
pd+HlF+JUCb0LIunu2THPNvj3rJ7v2HyrY4O2m/s+4fe+IDjgLfbiW7oeMsPZ8cK
DQ8QSoIlAR+N4l+tDWOCOKwfRQQ8C8dkx7oPZooxGrAf9Wu65pPyV6oz7Yk0dhfw
95MQMcneNWiccLzjKHlW8Q8U5RqXcbc4+7sNSVWk06450Cb29wZIa6sXuqNg4FPY
Z7HgCUG2IJ+LXVLeaLXjVflLIbCSJCUd3RZ9Ue/yOt1UaVuLm76PldCmzXQqaQZQ
hg2Cs2WD4ZxId8nna+OzFpV8Y0hpdlSZ5810DyXw1gd5jPU7BBZTyE4PGLQZdBON
1gg8dl7Vcw7/HuQr6z2bz1R5cQerqubSszVwOJfninRgmZSgILP2DnSTRcM8uT6V
UkBYw9L4wLVpFU0HbZrpXsRYlBuudxtiGpg0X/CkYuT11aijDhM2YJZyt00956DL
zkjm2DwBFwZBUSOKoICu/hyOH240I40glZqvU/2qRpTP5cb5wxlalyP8xyr1UOVm
sZnz5zQXqLT2CWh0DgqtoJysF4XE2MFXdfKrUZBoWtBJ35aV6pqnHqSK4wnBaO+T
SIARgD/a6THaTH8AAiLrcacKl0vyozuMxtTb4YXLIRIsR+Gf7B2ddAvaXLVXaIAB
P1ErsSoZnJW8t9e4X+6XYaXZx6rhNvcexr6JOMt1MrMZVPbtYtprDFAyxazlmhXA
9nADq0kd2cj4Pld29hjii86t4R4cmc2N9t/dlIqB0WvGkDOFMJBciUnk/MECHh2m
bEGz2KDtokK3FlChgD2FnQTd5oeEbcTThrI0cc8533s93VWLK1UD6lu42nxqyoa5
suCH+SVV5UbNEeJ8k7MGclq+RB3nSNLOszeWlv/QQMGXnQNQ5+UHdoxLvS7BEOtw
MLoTb2TP+WHLwYt+cYWvVnJS7O/ux9FCT2fTnIKvoZfjLyNfuRJ6qWd5iuwqGkQU
sg3R7cmbZno/N5pvf2PG7q+tVu1QSGtD5/rP0hMnqjQ9FLbVBV7Q64cmT1K/4uCM
a3ZIie7ttjOw4Y3AzH1ExmGyy6BUax12GciW5RHaoAiUm9muYQt0EX7UmL/aaQJr
w13HY/Ig/+xU1QJCy2Y/ZivuJCPkI1tst3JECfjMVaHNUQLDlcUNrSe4ZD5bJXFg
BD5nJJUFhxZ3sx4Zgrq/7rCCiqhwT8LdLmF4NYujV4AKTYJlQsgRX6ACwQFVXj8M
Jtka47B8PIGR/uSET/oC2ycZLyd2MlSKuvHokm6ghzi2EQFnPG9PyOKuSHC1zVLm
8uyP+prNpDOm13U66BDEkt9nYxJ5te0PjS6xUEM+9eBy1+DOUP39cw4+cAJe02tR
HbvQKc5gMLRJke8/qcEANUrfhqrmNGDwiXymESqh0Rwq4aQgC0tYtiHdX90QnRB/
6eZ117zSoixBbq8vW7B4yH5Exa1oH8eyr2kjmWgQBMTuai1SjQiH1oOLbd+tYaKk
y1ZQfPrzfDVQa0vzZ+jsv7Rsu7kx5JaasBYWhiYUVRmtxP0s4ZFh46zYisjD6ypV
xarVqBFTaArQX9nnttzLdpdob1cLaQAp/YVjheqKpvfJWceFulgH+POhfS13w4rI
RUPBh7jc7vPzxMVq3GFI48zPS6XQdFy8kO0vFT2oSBxu7oxzGPn0WJjTXqtj7bCE
Ppq+MlWhS8RsXeJOArKLmWfhc3zOrb2JyXc5z57cr2+JZ8XjorJ/hWGjfpdOQPGI
zPZDCasSVWbnLysMauXykcyCz1MiGKwl95OsJgmaojREFBLrAlucyGDieB5+qGf9
mNPr6Pgar0tXWPgnstwC/9W9PXffArVJciCpzR4h+DRoTP+Y32SeKNKgFEPypnDX
7B6SAZe2qdFylrS01XtovjN9shFKO8dOUCzxYbVC+QzWI47ErsQVdfCGG6lG11xg
O1+I0i3Sf90RIY42b0P/7adIFvsdcHcN8Ap+haESWhLLmmiqHFGEpfcjZiworTZH
IBUP0PYz/hCf8jXxTliE/OIONCbDYvnQAQDK76KuZXwN3rPfHG6pdjnk+bLmHp01
5GdXid6RhInaWHasCBfZ7a6NX8eJcU41r/lVoaCcbDWggIpwY+lLzBKr6puC3/st
ywg6tWQXarokERSZvGPstvD5562/df7EC9F+2zaUaqPPYUhtzdFb/Kd3yUWXj9TH
5Nv6uzlfOWyjasIesIuWVL4NISW+5Yb5V1SGPa7XddIfxIU4kNNojJRwVB+lFZ6T
sYbv5uu0Hd2Pl700LCwEmbdsV/JJQSmQyAGVOkzRKJsN9jB0UE5N/tvW/HW/YBPr
m6T0p9oLpskSystGkXYRwHdahaAP4KpXAkTGUkA41PdeCwmD/NV7VGlq0a6OQVMY
5Q6KqACz730MEnDaL1l2Bk3UwGKQifz4i8hkM2hZwq9/z86Pjd1p/reYhseBWEYj
JxYWY7UQOGntN7Wam1lIIAqCWh0AsxNQCF7iLGOfoVQLBD6OLczpkm9hASmTmdA9
NnSNALCSumUitAnsck2Qdew0/XKDTeaxiaDZV/WvEJOLOafaFx6XqOEs/U1ok6Db
mVF1R5hKroJ+psQTjV/IbDp4WFHKhKSbYwXhH+likn1FQj49TM1EoUJapAQkW4P0
5Mcb89FTPhk0CCLwhD/Rbl32J11oCsKUurnQzrMUVpiusez6UqTlMrtANddccH1a
CQq4dESB10cIG/q7bRSAW4VXk+2SkATLixMPvzNCoNE6y0EikETZyyJ/2YSvH6+t
+Tb01BPUlBJxKJFj3wtK1n/D2KNeyyJicSv9/s50r3TUKdgvA4CNlMvhqCyEofz5
rgUnqGeMi4FbB7ERF5dzSR6NSe5MU7fjVSZj3k+a7vR1tVq0A0aLNxVS4Q41WC9T
sX9JTjEjUiVtNjEyXrvZ+LrPYIerqlyTt/qAn5qDxS6R0+JEiBvKpzDMb9CH0nqm
/ZrfbalxsXz71dzK6IfaFC0u/2NhhrHiLB3heE9DxnULOawV/fyrie9i7yPdN5x2
Hus9pVWlL4CBvKXycJBvlRnAZ6cmbbJ6xrz9xu3x8GzJ40FuPaIsAhWqUldohvw4
Tv2NM9Ebi2l3qBO+cj9hPTWXye3/zJbc4hqkctu3El21vVubToPATls0iZpEIKBh
C4Q1kloQvuBz0zp5o15QPgEPCD120meB6AdfxLXtbr0y/pryS7IwGVpFA7RvBM01
RfGj81gfPNhcbvkeN0SthlCciOy5V1yID2kCSx8CaMcOq3rXPzMAJ+ipX6Qz9t6l
N1K1IRJxzTbR6SfGAIPF+LJGPCz06xgfqHSrurRz4NB6U3zOBaNFRFc07SCovKRl
jqran8N1nw0ZbPSFh8RUsDs8+gkZ88npyfktLU5AI8chbSaxn8Kt15v48XxP2Rnp
5mS4CPmuwr34WO2Dm0u9lg9jXh4SKVMuFDJuwzU9qzvM+MLJEvQrLxSA2MH+EYbf
Komjw96coYwVVrg/gem/jSfPuhWDvNDeOVdUAK18S6BOiuvTJ3uQj4ImyfZo8ztg
ODVDpjdFB5Fp9voM+KZf069ysTlBfD3ubEl0gQKgAiM5r9BUfCMIFW3SRKGSmt5+
wdO9tju6DRnK2MygALgce9RpSZQFbbTlHeJOQaMAJrysD2JmhMtnOzJgU+zdnZPk
LHTULTfJHuzpFmUq4JCC5JAve9+6mWCU8Cx73GGVprbyNWRCVFNvupxkYaBCoe4n
FNi18q3dWH8qgFFnYCde+0bcXBKPTigcrruV7UXinRBjJFN+7oFmYI9zcdY2Nl5F
YMqps9l/l2MCxpISGT0isWbNFdbAuVEzips0z7kCIdMogtt5x3VfE/+a7tpQ6jNq
vCMvZzcfh2JvrLbhbMd71CXb/K7LMGXd/cu2ZXQTtAVkMArk5QE8MpEXHx44aTaW
VX3EY3zMZht7FpHsakZzvWF0eZZtQ/mJxICDl7/LWQANyBX2rV+idsj1gSvvk3ce
Xnus/moHiwPS1hBidQyvjjMrGShQihAxsYcAed2z3ickjsfScaYitYteNhgiKiwW
ZXGs006/NKLF5hirySNaEwTl0ivh8/yvadm6yrTENXd9CoLQErlTEH5UhJEjfH0/
BavVYnWKx4tG+7MzaZ8ToLuhdQEujXpBrVmOI4MROOMtFcJSVlOT8B1qu9VXeUMD
7RNWCu7rhqiSb83KE94/bcplGkInlvZm/1nShn0KO9r42lMw5p0PY+O78DwLQJyI
HJevJO5QmRlAIg7fELvGEljAISJB+QTjZlLj3ydK2nBOMyNn26AxjojkdBJwBsDV
N0zCFie/nKcHRE8JUg8T8yQfZ7o9U6Crfdvc3bzOz6pQ1xlDPqkOkiwGiIc5SJAa
3H7GlCxlH/HBPUTLgDl5sUjuwyyj1/n2OhRHvkTjahgDK9+9V+HcO1vUwRjNhjDB
0g5HiLW5zr7OA1c5drTGBl86dWwSThoH5kDTT9wHaUBNPAz8wy/zKslplosiOh08
j3Pjf3Hn76NZHRQVbOj9JIuGyCWlkSOuL2ucDEwbc6TbBf+/g+2QqCfkm++B4UCj
JG6yTHEfJJ4ge+BFTi8iajQXF/U0upZtRWIspcyasfFRejY7aV4d91h/nnftNa2F
Chrb0bjBjTs9hiLAeR7g31Obo49n7+Eto2sTp2uBO1gZ4c0QwJHC1tj66qyQGQHs
a0WE6Ye5FcPhWLbBfrGdFLpWwNvsrBCiQVbvkpFYRaVBS6y0pSFrNI7OQzoKKdGX
lcIu0+l+6F2yU+jiJnqlDssftNvW6oI4JDCluSUYGMyzqPaJ3+o5eefE+lecF401
TNgHNrsPOfjtK9DBqjysqeDrfY0A5slIswkUr5TEOcv4bsd0wKdGzUg32x/bKEUq
jd/gzFFmDqJCKZxukUHxxlqEihm4N4lyC9SleWwA+9jVsY6CbXRwzL35403zefEt
pp6BDc71CCUn5VFL7dGETN4FTmY9Fp5rxXRRc06X96stZVfbU1bsKn2ew5ET2eQA
XSJMtSTOjkqb3vrNGptgBrjQ20+wheCl8HbDTR2vrz8WQQVNio4ZN2tdBMP0JU9D
8B7ofe63zRJjCzbxDONIsfavms/JVgPcYAT0ZurHMPfl2YJZzPlE1gT2RwvUBQKR
AlznJ+0tWdrSRra51M0XzokzN0EUE8XQ2DucyS4c4MqBAi4RHwzJ7Px4DI4YCGBF
UgB55fZmyAo3rJ+VtVtKDzxQ8j9783QZbAf9LsNnDfO8lT5yGCoZtLlKSCoN2r74
Mu/vCSMW62jH8esc5hGDN7qNcnS9RDh3c9w37Tv26TTE23V9VyTzkZrjFwZjA6yy
NCCRWxWggZso9DQV9rr6/1C8o0+6Dn7wf3KgvkBAZGAWKdsX9kfPLFmLUFONafBa
9VJjJv5Ogfg/YZZfBsP0kEEVjFSixscr3cKjFmCxmTmCtVNbrjj7N5SiKDsErx6i
5s5PYuHlko2aPZ3GQnZihoBa/8xce5qjhsvroxQ+200cIbj0n5qeO9k3roO9dI+U
T/F3iart9dzreyMxn+z4701p30sYqehEI5GLPysAF+mBwegzU4IFGKE6GH12PhEv
7N0IpKmoLtsJ35feZni70rLMA2om01JVy/8YaxKfNaiuk/XTTlphUzvy4QEWxTRo
qmX7YDHkviBTw+hZu2q5MqrjqBlkCBDTScisWhzNZ5p9Xy4yth/xWs03GoAAfMvR
QdgDsmBfptJB5fo+h8B3l7bsishTf61HU4eIddkF506uyHDXlT1dXj2a5qpwvaJo
CN/rEqj9jMWlxUfy7eVn5+VjNjPwDT5z55Zkk4eF/OjkBO05jiSSszWqPPrWFU/W
p99oXq9AE7OlD+PBmfKNG8QCAm1fvaCMajilLw0C+wc+FHTsyqvmYlEerR/LdKCO
vDjwDyui7Cj3LulcZQDJ/kQh37GG5oac0dAyjFTbnzi5REXimD6yrsPjw+Tmu+xP
6FIw4SPsBKn8rwkBYzJXRRdWg48CtqMMpeVH4nqCQh3ts/NfftdvD9bHWG6pJs7i
tDkzANc9Cxpz2nujabGckJsSQAeIwdeLrR6gHaCh7WKXOEy87EIM8ysIdTlVMc55
jhvYhyESVhAWlmWH3ES5otfED5ea8NFDG6xTQRBe2tCcFzJRMVJus1BNdUnfmgqd
WSkerV1s7WZpcazZzw9UvIkwIIu0JfHkni32o2W8sW9lKFlvKGb/RtdkRPFGwWPc
fEXty1Z5bQ6s7NQTM1lWzZY+sLKbJCwzg7G9fOWdC3fXrmtu/H0oiLRmmplFw6zf
CfDe17S/9QFKmiskOO9vaGpyq0L1pQyc+FQz0kwNrJ+xi4NKxM7KlopRMtwoeuFO
pPYspWlWKRQVt1/WyZWzKjlWLO1cvSkX5LHb3q1neMxH3Fu17S8HjIWU6nhAQJV5
J/yzCcFNCff5Aw6Cxyp5p/nm++kEgYmiPPEGpGwCebu8khofr1bXvChgqCt/TjYD
7ko/tRBdzVy+eEubr7U4t5Pbns9l9zNSZhIfOUOguKzxYPP00g2swVedHx602jQx
SQ9cmkJTwlpUsWmKWO1vM9y7CuNNcezJgU5bH3QslCJBMFJOT1ZCNq7m+3jvwxWB
zABoM8DpktWsmq49sSrYZH4XRJ69vhb4aFXCSyiwn30t1dx8siTT2RrIudVoufmq
k4xd4ubcjXReLD4I/QYYei3Uc4giW3dbH9pyUuBAS9AEagbNYxL4ARzRCySqyNck
iiPqYX7Lz5pt0CXJx/rr8nwIqy2ITjNy+O8/PeMZkqgFF2HHbaUgxi3N072Hds16
Gh30VyGNyb6qBTABIrCE/yfg0f8ErajAEj4X7xWK08SOXQHEAhwB3k8JzZS4AhDk
6uCuPWOPdyFABqItEmP/Q/58XIiaO7HyAIc56uNqVkD6Wl6NuCm30kquYJQdgBtA
9tmAfUU5reDnSE4jjonUm6M9Z6oHSv6Csxzpp8SWtBbO6U56l8sC6m/l8us40lCz
sM7+2ChipIbmMsntcrQFMDhh/ZJKO1ykLmZnJVJRXGRQ/UwI3iev1To0hcqtjkcS
IjcxnbrQzJmqiG58aRzDZDbyCGDeRD2NPRoIBjK4wQZ88t77p8iluqSgm0N4ZvfX
cpXnv5tbOQWVtV474yyDRagIMjUJMW/FcWXl3Ss+Zy60s6LBTn9+OwY1wRCv5YGx
2hIFvPzxjNKTrBmzl4VFz//+1YHseIMQ+YtucXL2sL5+/ot9Vlym7ZRCn/XzOXVm
dWUE+lquI1nrdixCg1dR8CxSG3qpBBVxdOvAi4EcVwou2l5gPmGgGMHUtRFPHtWo
XA9ex50+kyXO/lvoF5xb70nT08tMBWsxX3tKRehtTrws9IcU8stQtKgp1bPJ+1Vh
7GP2P8n0f6Qtmo4jYuBgjcZ4koJSOeHni+Y3ellMU5skHGQtHMgBTbyXPQyKv0ka
ufU82MrNJLKgUSbxJQPBregz+b/JEfGcly/lGlrB5AvJHmkUsx9BS3NhGZMCw+Wr
CoT4Us+AqPw85BgVDA1ytOy9ewcj23JtTut+K6Kq1qg9xa2bORAn4jDTx2I01I0J
njLDZHpMH5wsN7o9jTjRl/JIoczmP2arPUVEP02UY2rGBjsufsr/6S2uQSIJN10G
ygjLMxQZXXg96AVkehavHidfH+nMMhBgw+fb2+GGhDNXZdln9ox42Y52Qvc2jVJf
USD+LVTwdIIQEua98ibKTcVFOdk+uCGB6Nyn7zT96UvvyoerpqmKBUd1FTDgviGK
O86dP87WI+WF4Y+9Py5LxcBq8B4gJf88kbnBqXP2Duhssk5tSDQ0KeLCZjTM9Mks
jwwUtTK5GlB5tz6yLgV14EV3jsbiD62v4INA/JQkkRUlBqwN7BHDl5HqOPxOj02M
j+gDqqKYHohDyJtHjq+h48eiG3pUbXkF7+vbRYHmVZK1DwORpLcbXTxQ/u72SRPo
skOLvAIpkO+AWqJFWKC5uVrEpbXAl4cVamaK7e93WiUtzbosw3khfjShUaaTt6fG
wJc1eKpuyshgQyubXcQ3H5BZkGG4Rm08FQxEMsyHNhwzjPxbIixnFW4ZI+i580od
kZizTPwso2ILcntfhTfNS9eKamS2ShX8/5PFpIbgrh1Juyma1fkvI5n/OpK9naJ7
9UYmI5kuQHdtFXduqWt9Z1jMv7te0a60cqoDJ8iqcT2ajkStwD324l8tspODOSsH
wERDAkXpE+LEnY3pafI55UA+03NKCUoGRDA1Gb00l6YiTdxNU/QNxc7SUuzxFo8O
K22Z+k+oLJza6UNvbegE2oQFufQBnwvtcvmZiLkFEh9aPjk8nK2cqqU+vnVFPrwA
ldFF5a3mcP9Mj/qrIPVKQuHdpUzzt85h3OwnyTCNTRwiiut/+htMFTi25diEtBER
qpgw7ZWP7ZbeCbKcbfq32bSO4RGmUH5YQSCMMpPGVK/SbH+/tJjuQu0oJDxIKphv
M/6kuJSYcAlVnySstGqkf3YVpASLT89ZnSmh11NRjEpaas37RHGBRyhYZ7iVUa5r
CNd18tW3pjTrZiJ8xANU6XmG9hY/JsdiElRKIMZRuOZx0BNu+tvUE1MC/wUJDWo5
XSSThw6z+pc/ml45BurgFZ8TG93O428pZ2xpj1DHTeXlgpQaWgbqlLxxj6SHZ8W9
2xQavpLomWstMkRh6pMJZRewe6DhbTOMtdtSctT7n3AYFYTliiXEUc8RlYBpZUMh
ZOz0UWlOcfAi86OPKNxbR4IeA+8rfrTzeE3yae/lwN+ISp54LsXpIyKSzft0jtQy
bj+P/5XcqlPA4NEmo5f6jXVqNkeXf/1nLLwFS4F3F2+4fODJfZ9ZGSduT7gWlQJP
fpVBRUKFpyyYbVQm82ozjwlY6ZDwK02g1JGNEq0AWmhqcLZSlWeZGhrozanqO1Np
qx7a6yUy9y/M75kJIQnhFIfM9jQrlUHdXuWGaEMT8xxTte8XkFivk+gf4DiNPxAp
0B9X9DSolz5hz3a6On09Mf/qVobWVRQhag6gAjTDuksQYFF2Vh6IlQK/NEpDqseJ
2AtgtY5MUY/GXTVhUZfInTQW+BkVh8xaoJ1lI1jrU3oO4LVQAck7z2tPw6eKyCk7
5ir926bcT500qkYgVZY7x2kN/XDLlv7MK52uVLaGhpGAvdxLlhS3NEzQj+ig9LRP
vJGrzHiwrF5AlioTDd1bIgbys8yLHwHYj/P3KDvlM+aOpelINzGndtIUG2srRlhd
VZJen3raNGcDBxXrvxXaWSlZC/lWwX/bM5ZLCYNah8CVQhtNHEIdkNg4U+A2LWS9
kNyhEdn8BJ33lpWeS/t11LNA9hAPx4CcxA19c2B6uaSEbGDeP6CZmmY2xCWEHqJs
BBnW68vzKGqtvoiPaQQUbhGJ+jGQoi3Rvu2sTtsKEj1m3+tlwSEYW60rfsfSAm8M
EHHk0JpsPwMnqLQ+9zoVgbno7gAKjJIeTT7YWvLMQxWvYHJK+Q6m0Qfka3CyzJM8
L8afRaZBN4ayBfBP7CcHtTBvLObKqWu9sqrAFvtg1cfEjrVqA4FvR9Y6u4Fjhs5Y
AjhX5ei3rzl3n6p4nMxE8l3A4hj5PQRF+EXTxgFBXpv5fse3I5qp0JfPCX2uf+EA
Edrui4B8fp5zy8KLm/VWdsvG4k95PMA0yk+bHprBBRxrj23U3FkO0m7hdGHGp/dz
Sf6R4xBb2s+8LasGQmxZw+A059MmKPpsTeCGzuLjd4Rzf11wYI5xiud4MLhxbEDs
6sIeUA1HLAoQc6qXAldundzhNhsnw0AKF8esVHxCXc73lB63qtLueM4jeP7GuVtl
ObtECjnk7HWWInIpMBmvXUtq/j6XLRSlz+YKI5EtXNzcUlHhjrokSV3wHpdsi7Bg
SuMBib+Q5iP7/ubgdqwRkjNiU1wK/l5OuDV7/DlWQuThRWVAzoF1wOE9Z10uHPtF
3qV1okdbkpB9k4oWrmD/7xSuIMbZ6V1HztLV2y4zh9HtlUNJ99DcXlloYGmjiB3+
ibV9ygx0TwnpGjptE2dx0g0BW1KCNHr/7R8lb18rvSmFBp4KWqjFT00zJzcpRsza
GfX/zmAUQaLGP4wgBLpmwzaK5Vr8oXS7mqcLHQ9qS1a5ZFjeaWUhFOUb+7hMpIqN
0qg/PjNqktDbz4aqYI0RNvQUhlR9QZ5VGO9daLNliJvIbIK7Gtd0WO6K6YmUpabv
AqqFRauZjJfXyr97J80YB9QHTBQYtcQt8JjJ73hXm0oQgKsRSVtDc/8bQBhWpa3l
yv8ZXgI9AthsDZ5kPGcBmnZ56GxDtzl32jwRWlsTr9gkNHhbaT7t3Xra4FE1WqdS
+efCX2gHCma/g9m8tlCn+LhTickC7m6+P+1TnKE4+YhtENBA7nWvWrGjuY5yHxaV
jAKtucy9xOnxCmz2ZkRMRsxNG35PG11fXeIrlNx1xgykB1gWAHkA7IffPt90I4W+
uxyTm6k4J7QakUuFHO1Y8gWfSUmFVIC+5WN0diZkz5YlEcGVKrvrXPguWU+sKl/H
/fLQ0MZ3kFQ8y68yF1R6ITp3r//RPfl1hRqi2nWBp0MAhyDi4NgfsOZMjgz0F8M2
whKc2fJbuY1mCx6PyviWnrlRyJ8wZLwh/1lwiBQCOO98Q5por8JJOvHrnD6O+taO
rpzuhFFhow3LGAGU186gcbhDoVQ+vXUyhELF7n1gC1MSD5hNjdEFVPRradOMuMYJ
dIdmW3p09NrSq4vvHEuzjz1oYjiwt4fpoRYJe8wSiuEmK7B3nZotFbpXAOoU5xnu
EK5SGISqnD1IXZgjl+MXtThryhvZW67/D0Q8c+9dg4Rt3l6ltipj3Zn7r7Lj76dJ
o7V91qgEiY5QmU8VH1k4mxObs/97en6PxnR+ajHOFpF+Asde8NyUodHgh3fE+q8h
Z/bo8IwX5IRKlH1TEzGTB609JiYNxWD8yVuU0bWfJljwKnwplDQO4+i7tvUY5D5Y
m2J1GLSgPkXInA47eMOJlHhKB2hV7Q8lxUCV280xYUOcAyCZcFXONPD/EWRR4WX7
MJPLgnVLsJwg0k0bjZH21ohHopEMK8DyTD7nkP3yh3bEZpoos53zn03kKVV4Ikd5
e5u/cqSdhwnsWQQHNe7sMF0xl2DkLa0KKEpVXROamyox7c6dQGtyZJ1zEy+vOmh1
sgHdiINDBKFAtm2LnXlL6QQJaO0o3fQDCqRQKiM9/5zSkQVyA52v+GVDpd7A9Ys/
QbTuTdQLYHnM/kkqVJnHBlUVslwP5uNUvmsAPtAQ1Ur5FD7gZI3X2NoMEr1samZv
X895eP9LcygCRMHPkxFezZhBonUVwO6d+9ADo6OXTz7gAK1bQawfoELtvTmZavsC
RZT4YpdMqLaKptMWrKBz62745E2jtGhVSxqMn+hU8rRp2JRAeyTQ5RcMKa9dMoZc
ZAPpbl+fcVFkhGCLl68dMisjuuBuig0QmQyA6Ez5vctMr+pr/o88HRwmQ8xNSmQp
Bgu4LSy2oOtmq3kKZGoaxfY0VprlASfXvgrrRdDSfty9/1zPj+V5kJrNZXtooPOU
wIFhDpPI02rzZNTTpzUkFpRV5ew2zzwaitF5kQiZpsLOYPyO+2W4z40M0Zc+SHa/
Y/zqfJ4q42khLkcB6ZxrNysGjrXnjJaWuOEUtstg8UqxA3UQCPF0sJaONKYxxeMK
sAJb8WyNxqNS8wqbsyts84xfs9qitm+gUihpFRciY097KzurScEXge34gsaMNqzq
ap/mKVs4zkwvRgDK/J6AQnD8/h9yxUQz7Td4Qg/GugCahOOZFTRXfc2LHMMoutjq
5UqHxp6EMXjw8ts9Uh8iNUfVcaa5aSCqCAPWR+yPyhYByFmpJfivfwaS2+J2RxOi
DRzJhfKNciCWt5DyACs4Xhu8uL49lGAIDu0uBbFeI7NhSr7GGI+f8e7I2Jn6mfa5
LkMqj1bPqJXy9hVNTffX2P6WzoIWBqsqkaPoYoc0s2bbz0vWYSxVbs7fc0B8FCGP
YW0JHu1bE+a+0TFui1usJrmRHr8gLkNDY3RcDjdlK6wUatOPueb85cxx+JfkH3Uf
4me5kBweO4feLqEoJX+Pw1HnnKtvEn35X9ViP8+Bt5nRDMnpCqgzOxyyh1G0TP+4
tUyf4/gkkZb6ZaagMdAc3SHUT4SnrZdeaqzSb7jBgd6LQE2KiBtcbtVky4Yf92Qr
22QFdDTmUxNpznfvIFb64K/7jWw3Zpc9AHfnU2RNqPqE5cfU3EhWU0lfSs8X9aYu
+8aweE/Ul6srEsrAXThr+EZ78mpn3RHaYw7uzojqR9DFkHAQ4J152woddIzUSZba
MStIXF9ok4gWXdw9xuQ5Tpf7GHB+OIk+ZYZ+4FvlSggLR+tzBmiFU84VK9VXKroF
etN/TXs2a+b/h/ZMLvssTpg0Qp6HLyowaJ25M2SjItJ/v88w639bkNMYpF+d0ERw
ny//0pZB6GgG4+PIkhW2x9dogr6kNNR3wQgFRr+ESsFhULySOrV4wy0VwWIsxLSA
Q5txHCs54JqjsLzNsYUQT7LjTuxuqahZIbivG2fqzujGoqeIqGJuH+daAy+1oKla
8f/oVy4mf5uq8vEQnO3Us4HPiU3G+zd7nK/1Y0PqwgiIuom9e9H6Ohk4Nu9LxiIk
3QK24oXkrIerp4j340ScparRKkVhjd/m/wSMt0BXh12Rvc7aqWiHtuwPPXMV5TDS
mE2eH0yMIwlzqPP55qs6PuJtz0rRNH08yYPGfdYiO1F9MlKVlvvnjI5qvSzBrt44
+dyukCwIFiYWbfA1Ia/lMAIZQ30IvXU52Wl2lPnUtFfZX9MXn3Wn6CF8UG9qAMgc
wnRxbSo0wYzsFYj0mTLLeQegDVq0NxH5vdYS1qI0c4BYjGRr/J+6gf7bhMEJr5On
2DgnFF48vYD+l2jhzZDWSRSLSpDH7GLkD6XXawO3Wt2rxfj+EQ8CniDRDuyKZ4q+
PAfV/khIOxOli40ulRHFnoxxexbHBFKTasFYRFX0XQ1all3rNHRhRRaTeZ0ZK1Iu
ivUxV2vZA8xZN4q5DpsC7Ekd1WfgXMmHt+DNoBStDFtqN2e5hHngAbJ2sPD4g5IS
DmJs3g+NGHSuT8Zw16LtDTeMGOA1OOlvw0kYhP8OccDV3qzvjne85dVQOpCWcUXl
NUsn/Q2D4iVvRL2ejZZDn/cc9kZ8wH3gZJlbfmyjduJ32t5cd9SQMIW5vNpRYDkv
cQbgalXHzntf3mSXLFRPsHiwmg0eiZNdE6dnk/yUgN1/8onlOHlxg+hKF3Nkd4rf
Uen2j/f+hdvTIH8D3wQL4bz8LBbLR4ewfsdyDCrzOaAlbQ9+i8aA0K3CruV2btw4
JHd5ybH6liACOCu4cOoqM22DMFibpDq3arWgZYxGrZWeA/VHB34kucdZ8cn2lZMn
ZKCeGT1c2tXMdKJtNDYR6+Rkb6uoji5QnevructG6MwpMOCptSOSMg8Df5EqGtuA
CCybfHlMkskXVvodiJtOUk3DBjSlka0NxwDlw5+5p3VS3HK5fs4wyV7/P5cb6v/z
LbXaolR5xE8iF4ijcsImvDc4mXQ0QV41hf0y/LVF/NfS7o9c8jyLi0aSVgy/50qP
dIXvPu0oqjDUONosx1e67267WPWNgx5Sex6xaHHa44CQUmqxWWOQvIKGoV0dBwvh
aR+m3FIFlumt6Uk1csfgCwSttpGg4vAaUEZJUKZ6HLFMDSfOBQie08Uoqu3qYHYV
gbnaElX7KrB2qN2xmkOS0ufJh+YvUYFdk5LGuWXVXB7PkZ7ZcgIuKXrfZ1AbtPba
LFAdNXTCJ21OK206g2Y8H16qKqNshtFi5eJMgBGkJ8vblorl1CpR9QRwUzkpi/oo
MmH5R8GirmcHStJmbFdvhFmNezB7T8zmBhmF+wJIOUDJvF97bf0hXNAfg5F+yBSK
2lnbMjmMD0EeqtNHcc5gCG4T6PgMFWttl0dipL+SfFPttlF/uDHi8V8wDaCogJR8
bKYjudnK9/awa7ozrt0+yZz+Fj/fsUS29R1TfEwVYgsVmID0erKhIghWk2HSuRuh
oUt0ApIaSqgRYafydkd7z70DdB19apg1oM06eHkfDuEEj46dRHEfDi6nV/Lgw2TD
aWHGQSoOrye+RoznHb/whXFQu2MQjQ3GDk7z78+8kw/HCqeL9U1gUl7jhwDrpcBV
n8ftrBMPhCadqwlGrN90BPxmBRNiWxVT9idaKQgK4s1d25M8/oQjV/qavViBgI4N
BcWmJNAnBLSC70hqyA52MYfcl8AJSTW53TbZYd2oahlP3/hS7SK8cFQVRrNzNRMY
xlNrZBUoTWe4JYZ3cQ5Bap7mDE1Rxcgm4DhzotOdNs1DaNafdKWgVXIosJWRnF2Y
iNeQYmB72J983dIN1numY8aXTB84oYqGCZrlOi+1MsCDZ+wqy7dJZAe8Cf8LVWjS
qPqhlufcreyOcquPg3v04BOMJqY90LMPUF+dCALq8pDo9OwW1y9uAuoZt3W5p8C4
4o0upLBmZL7Rjdn96N8keuYA6dso9GoFm4sJY/w+IgxGRWKIIhYgizKIb5Nl+5F3
cu9EhJ1a48BsO6lDpP+oDyC22TrV7YpkHKMX9XJ7UAsM0MkjrM5RYlUOWGWBAPy5
kEGJYmD/7v8E1nIwbzHjiiKZzGQ/H45QdvCxugZBBjbYsm90WhuHjBBaGdVrIefm
1xPaQjOftCLG2+uM+8NdxnG6p5qjU2bAaub7BNAoG+W8qGH/WlYAfRUOFrXpwluX
RRETFpZtUF8IBRS8QhJFkW2PfEBNWdav/ZPoWst5A/Iopec/RN4wtdcUyFiJE6HP
kIqxZf49GFlMdPv/qARsX5rPq/MH7b8BjLVznOphKKhov93HNqtpoRKIMhYIDBRG
4UlhB6r9ZnspUd125dK1y02kN71VZ7AjtH0mB7JgqyEye/JKdNPPEjuxzakWkEHm
r1u17Jtwl64R32H2el50QZOtWkOlesqQ3xzFRB/mkDhf6hftkVg7hdTGWCFKiXKB
qzke96b1830PKg4f9RLhOGJcewaJqDQ6a/V2mQt3lRY23rbbBfev69KqH1yD6h/V
nY6rw4PjUmX+Q4oFBVOwQJmGXZz3UcCd6xX2y5FqOuTCTwABjEHS2VcVMy6r0otT
5lrVIpTBHxCmAt+Sc1vGVqXOwStvv+A0azHeOIl9cBSRskS7Bklvzkvcx5OpMMvM
nPXCnPAW1/eJbz8uIlVGyOk9yLvqO+Kjt3N6S6wixxoTNOLndE6UkZZNGUQlCD4f
dykU2jJqGMPwjJsQIAEFrGgeEiIAZZhTcFFNu9Y+fdBFLo2MOqFpEwfXZRAX6rt+
FafpJOS/6nHpIIY9Cq7oryuDgDrJl4LHQ4cW+3CF6ODqh++9+bkJIJUFL+BxKSba
fLmAwKgyDvInW9eRx6puOpR1omb1zVQxNAfN0Z8FqI8amInMJrAPK4UX/hf44xdp
w5spBReYKXc40u0QCW3CyleI6E78CO7WwsY300emmlgQ6ShcXqpCFXlrhY/Tzqay
7pr5J7BrmPc9t6dfHVSwg3LRIbboWk1xLqamozwk6gxjcx56YIKn4tvqQubSf52M
aEqR1kVlSbfrSmJ+AAhBLISPLHsppmzRllirQEaWq197pscAf0WiH3ofEtUeS0v8
MD9xKYgvk2oQWn5cvMp+vzAgEosQ1Nufw2NChzXEHnIAqqykCrk10saYuYEptOwV
JDF5Q62ga4hF7W0Po49LwE86PeNdHOw48Wt6FH9GEGJG45XGMWq18sLFWwy2oJpN
xy8/2iZpuwcD/RbIqA4//m8/tQK/vRmD3ZMVpxZIBjVvgRqDd23FBcj2q7fT+Z2f
Cy+8XFVxtRXJL1mg3Hj4jPnciPRlnGNTS3+F3F27YYJ8wFjmp/Hyrr1vAAbmV1Ax
dGOK163hXoyySw9I2MqfAeUAx+UFS/6u/Piq/Qr6sizSf2u7jddh9uI4bp/Ng+aq
fAY9s4ANPbcNGpmB1PKHeF3moDVTeb+9CDIBR5yIQ8A3zddviIEOpK78TN+IflHF
W68ErlnUaer34usT6+yqF7bKRVMJ+OCo5tPDE9CRWDHoS1ojVeDLLM6lx9FNMgDD
cIYhg+uJpYOgarv9EW32Ku6QwUrWDx9PJAnXU7gHTPBLl2PJbA7uhjnOiWdtquoa
mnYYm11e/VhOwnVybfntz3Ezgbhfov8WKgm8LjDPoyQ1b1Y0NuL1BX7Rr5pgC+LB
JAOiMxeihJ5JV1FAFp3Ri+GMsU6cl/WRomLiovPiWlIxSLp++TjFtxx6CxdHtQaA
Vt5PAe+lBXDBcswNuGKu8MyaOhKYaITxwFWYiA/NaBSyKcW6PLryQKEPReVuvVyH
J7aJ30oYsyAIH34Q1+lkTJOfzyfEf6w1c5cTsVcrN+kzMQps6hxOWqESEYOb+9xR
XoIj8Vcex7yOzVNONZfnEfwIs8cNF5bAg3lcL014DAMCOCuT+GccLy3jHTG48OqU
HEaHRoBF8WEkMnLTW5Jxo81dM0xFcjTYNTE2SH78e8amvjQo+tiBFxmudxTJJBA8
qRlcorC5S4ZFmJ1uvkaFzGxxAS5JokoS8l+ALWzMxMsDNdnIhhI4kBUZQGiEAnZz
0Eo7cpb6r5QM27h3Ja/tK6M7I9gomkmS2bUqR1g7bs0l09S1YX31+cks2DvWileR
LLCsOOaOwsGs6Y2GNNRpzgUS4n6A8fvRCrdUWiFUrpilZw9JvBKG1LW5av/Ts6E/
PKbdQ/uDqDkYt9OUMDQhGVs4k+0s9kahGvvbcMgrWOXae8+6izR7SEP/frw5JUOV
yvtaV5gq2JzRDfRbviRVXIj3ihRlBRMd0ryjzShXAIvxIN+iewRNpohHAJkBQa9L
guih0cmx3RPvOqAJ8TkckFbh6l7tiE8Hr82AbiRMJlL5BETNPBV4ivKQDhSJtnwy
uzy599KfeppGrLx3QLYqHqE3zddePmnWv8u8pVpNU6PbJQY2s1NG3hnl3SImOKlW
62lKTJkmcsD80FCfNkv9Y2k9GBtp7Os4iA1oKW36z1c7lRZ2ynjbbgHK9JVY4H/K
3Jb/6tPd09jQphRGr6UXwilIfsjKpnqSVa0zH+w9X1vWxW7JWJQTrOl3NCYGi+ZX
htU+M5nc406vldcd7y/JlzzbDyKwTJZuCVssEzdJ3UVqh00TRP/efn/F9RoviMjl
yRWCkVd1Bw1JqjIbAvE91JEL7R2XvN2IY97efoHB82t4L3sXnDVSDrRaIEGeKopz
Xi7tcHCFIlxg+iiNZGmG0mt5ajyQ/SI2Q0Z9maI6txhbL+DWyiFC5kMkGO+9M4os
hJTmIIrXdT9hq/6ntpXdp4aYftp9SUc+RJ3QNhD8czN04jkts18tnB3VmDUKvMzD
AvFTQjZphygeZWr3TqZKQKCaebaQIrEIm8Vfm20xXf6UNDRfPB1XCE8/davjAvaA
7Mf5Ff+8dPe+ljsV6tMDy5Mf0u6iSjYlJIjT2jecO8WMn/vy0yIrtZgWAumiW24/
nSjRjiDJYN7QsEyg2vQcGdSIW5F92CNQZNmwX/bwNkUF55n95n622mEjrq2+vyOv
OBxuvJqb9D+2FjwIOo6i7rBTinE09bcqQ9+s4usqHaCjNAQQDuIO/ZAam1P/EuCk
utQX9qd+yBFi/VeCKzl8tC6lAH/z1kkyQEbH7purJVPj79KFLgLzG+aOWSUiR9oQ
+cp9v75wrO1fBWbZ6Ad9EsUMrlfwXenC6g2vfECnSJh+rRkxHSz3Tjf1I+WR/LAE
XoZMJeX2XmRPAhktuYC0wmU7oVc7OZvoOnjY+G7ZqWbigsLbDaMcmnrBdgDBke0W
DBaU5k7y0O1iUENzK1xIqFaTyRrwCYfvCg3NEu+YvVI+tnAzd+HTTnbQfh4zbdB4
e7LnrawKz0TDF5/QAAJg2TjZJxuuNihAVlm06jcHjSMFN5+mg7XWnz7CbIv8VMMi
KF7FLKf5nLlUHSXrFhic3ujKj/4uygNXCvn9LOY59+wuxsq4MJt1n/y4jvBaa06D
S+Sy9/HuOpNHJxLdMM6XrOz6fw80wtIAf2S+/4jcukJk9PacwsLoUui4vzcpSnQP
47wBq6lD1YmHoCgQ+Sj6SVxSRrDsC6Kya10RLCZfYRoiNm/BrK6i8cIDAIdhcbdd
XNV7iOFgOJSdrSJnlViizRyIKCY7WsGpkPHpr/DZcuaeuWpeFJgjVEgP5naJAzt4
eUB6klLziK5olu4AACVsuUkbl0ehWdQZDYzPhwqbv+xL27j+PuDnpLoHSNMESwb4
F4vAM4ofDS8WsBT4ZcvSWA1Acbg92gTDQleCf/xJnqkomhi/wrJwDM7a5ONvvWOm
XV43iERclFmXWPop0afrxfmoBLXmqcxP3UoFsU0cAg/e6UulHwxJwse983M2p5MW
3C6z7RTIxiAmBygm6CXyDT7/OPIWBAxJsgr2iNvLqhmrIYiyfqXs+DJ9Y2Gf/Xes
YA1vHUF5Kivss+lUPJV/R8NyPhbYi4XzkNRtXaN8BBa7fQzzgtcAQ2HQq57/lZpn
vrFdqi8nqKArDyPhGGHYxtvxrH5or4uUZ8YkZ4p+EWvtoKqirU+T9NcX+hFV+dIM
cyLjbLrTPBCbFOlMGtjVDHgg3QBXv4UdOgB5SwTeGeoiLWgtn1Uo8QOF5uHiNuK9
t/uAFi9ZB0ct9UjS9b3t/DAo2DMiQuyrhUD352PF1Yh2zulUpm7Yo3YG3Ojgqre3
jK3huOBHHmUAPQWW+aNvRhC7bml0fiV/lgMZqLM49jKvqje+YZO6DGe33nrcyEXl
fL713Lmp64Yq3NHlH6a4u5dtQSrXpnzgvm4bntAvdHMZQJ8VQrCAV3svIupi1bYs
YLqcrRmFljG39S3gMRNKG71laufbCVMpOA7cN23r+nTSCfR40pLEaCd3wa1/x896
eT38F9bHi8TpKfx1m4jXpJwJ1lhjMe6DxJlsPfCMI/E7HaWenaPzYtUuSAvtJIas
hfqA33JNGc6WqVxyJuxjN7WY7kJIfck9py2MuvGvnzoGPjn6oV41kSQVRkbgTSq4
+k/6xZ7o+QcbKkUZHDYFTFW+NKRIjOy8ecUktHIr5BJ18vw39x5YATnwGmCg57W/
o4d7JT6Du7jEQeZbzfgwdGE9dWMnUSOUmYmZkt9ICVgxVNyv0uPJvMsX0BM5+fLc
zbq+YLygsjlLDthVcK7fqNyBIk+RBj4FffXf0e9xQvm8r6iVMwW6mv+6OAE/c9dG
DuX180poQZ+0t5ylxq7oM0Q9+HGDmJGJDK+3KCcGfBwGBoEMC07kc/+7QhwCr9N6
6USnx/syxskB+v+NtsxSR5g2vlNZEeWKTiq6xboJY7iSzzzBeubc0U3XJttNBWKo
Q6C1wiWBK7acDNWmhPQ82quWwj+X71hMhQu3cFTpI3/0K01Cm/ecVCdwyaGbUR5Q
K5+qHpLFsWACnmW2veAAY6SApk+Uwbtfc0hIQCtG4S1zqm81/wGdkuGXFq/ss/QY
7BRzwilC4pXWjumdtQjsoEbD0AAhsjfTwfpc5QBlGNL8+nQgCsMoplEVcEAh7OUk
lJlis1Izp2L/ISfhvdYcDY2VkS1APhVRywN+kdMcZ1d749UIWqUbsY1YkAS7eTY5
t+FwWIJDUYk+UUmoj7kMOfF7/qJa6zCb+gYmmpUPQug4HuCn8CSkOvn0cjfdZdBl
Jc8IXhBGsIRMmxnQyxQmLVVRq/pxJKvRw6Ht2esMBzKKIqHLwzEFlGk6Kw057vLa
xFC1fV10qSOnKZ0CEkexGvGwjeTpEL9yc2HVXdSMbAwlBocvEaKfCOy0ccJlM7xJ
S/u7bXToS9MeYR04wyMggWdkmgVDMMsRaJt2fjCYJKZb4Swf5jYXC/I15MdcUs0P
IWheMh23XyZZBQqYs3SVu9+H5fRR0vFSiKGwWfjfO/EnY/eOM8Qmz8qowc+0xsfE
HwFXkBXbe91KiqBiCdAjDv4mMlpR3I0EWDnd+YJDBSEP3hPZgRc4UuJxQEvZpnFK
Yg2Ar7GMUwXPuINE+G6+VmAHGzr0bK/TWGuKIB6eC/Jz/t/OUTgJZjW7/4235SzG
j4PlY5sCJ2LfBoedvUgGoAKUpdOZMpStSRhmfYMb71WbgnpjZ2U6qC/Kyw1y+VxV
pqtLd2+RyV0b+kAWVS9g/uaPuafXxCVSW6LNPuunxz0QNsaKEQwbF1N2/cE8HKqs
Fi0k8ugJAFwhbF0TQdT09WhnPF0gb/GfKpT27YakUN8xKB1vYFeT7TXFAakqz9ln
DOmPtjugebCzkS1WYVV9pnNbcNGqbWzkdP9koxpE2EPzNKCAfifAz1KtOEEQiaGh
0wPWmfobi6nroO3bYM9O/af4+jBFmWJDOCzfr92q7MCeu3wxqnas1+KaXJ+u7QVQ
eZ+2TjQPwvFagb+qgpsTdePFhQvhw1AaoPitGZua2T2J3e/0PTALDXQqrVDTILWI
UFMPotzavWTkTeMMvgJREUN0uK0BKeJ7XNHzEjNQKrDwQVg9Wm8ygDRB5MfjR4j+
pGXPriFdB5Bjr5ytMmmKJc0WxiCu+X6NsRZth15E+CLkw5nkhb2vjoReupj6/UgL
DoDEHAjTHT5I44LILpWrxZEolc9LPFrYmOL/9vREYWKxRQTQIoOZ5auKE7hCPANv
B1sQXAfpOePKzXe5d0FYkk1TQc3YPMntI+xkx7uY90FMHJVOlKwIyAlYFMRpK4qY
mi+2D0+W4BxwsKOf657wJK8jMK0Qz3A5mbfVlR5AGF0t6cLJBSX1oRc3QzmUfQ+6
78ndIc1idMl4aXvfDc5rC57oZozd9qu0dqxr/4BmhDjuiCV3wnJiNZhYf1NGCWFJ
VX1T6dzw51xPUsvuAVq8AW//d6qyHuOQAqyqodFuKULxUZbttl8K6HM4FBDUexxK
onUpVc7oNlfEDdKC0wISFBSrMFftIBle+i/eXWTR8t9YVadOHpmh3WXuwie1Rxwg
9uenfEykPcF/1Bw9QbCc2Xm0K3QH1qeBRkptd8iJcN6D+R0Fs/jYyAvk1Zsj4EKl
pODSKDMH9kOIcKrQbWDz0sw11YrmtWJxsZIfdLRnh48ZKpRFgirx4ZiMED5xOc9A
Jv3mrKEZxZ9aN0rUOhozNxi52DWwAcbAwFWgSH+6M8uZFRFcdoJpEuy1oNQgblrn
4yXXYDqnscLnHPGFRsWAgzFcpybHN0t35CGesxu6U4+lteu8onnvqx63wGnTByxg
BaSLEi8T23lzxi9xoBbvZhRU5bOg3gHz8+VeH+qNXi25zCULm15ZTSfnsfQTJ7Dh
2AeazY34EwaL8+1V4951HKTPBA11adrWZqCs1NiEKLpp0jTkIRKSbEMPJ66miWoz
6Y3juJihblORzWKZ82244Ef+YDQjwnWg+KSnvt+Ou3pkbhW3P35Og8ybSDUNO8db
z3Qzo0ahVY2WsiH79kXNjBYu+NispuxDc3ut1R0baR9hyCkMtBoTer/v4s26PZn+
TzknzqaAlDD9Q35jRpG2PhbR7c2oR921jLVfc51exoU6UieOgTykeMVXDt1kSU9Z
JbsbCj3umwomOYLEMuEeObJ3SRWoNEKIwUdeKgIAfJBl2Q3s9Wk3SYmHe100uC6H
5BKl5lmguMjRKwA8K1Hgc7X6hi09HtR7vrlPeX0y/XM4oH8p/o9deJFl5jC6XQkA
3q/Hg40p7om1LuF0WdGK157tQb0FnXyneQ2peln284NuvWdceNAIzJ1WjTM0u0fB
K8Y8EAZuB4vIIl1VX7IcAORH8IhhfzKwi9Dd25YHZuEPl3RHpniiCm7r+0hBeMi5
ljHhcSbt/WFFrGLofQ2ApW9VEfCWtJifYDkrQFhcXsCrhJEGtIXxGRfxijrJLtNn
sfirk0q3dYv9GBhe+QSDiNmriNgUTLF+vKKlGZGqyY5Cior5UKXuGGk+lnCRYc9y
8nqfYyCISg1MIkpCc9YZRd2YtsNgsskACBJPqvCxmSdrSNECAMhD2/gG8gZ+440k
u6hYbDpQMv7/KQZYnY0fBBLoV8/DAicGsC/vWEEzj4ByK2b/qFRNzoMrpJ/T3Gey
0J08FXPCofN9Ngt4hGiIvFumU4KuwagCf3uZgQnaS7I4E/Ez54MDhYatPick+rpI
uTsO9hd09w/xFFQ9HC0HQldexAdGS8y1r9ADJ17iOhpGAVnOhLpiLn1vOgTNo2wf
7KXeEmXi14pET+yX1WN+CKgQaG6qypEYO/vn47kmZzIMNiRQ5NkuH71f1BqLEI1L
EUyeRdDSsy94s/DSRbRXZ6xlbBGQWiGRzrYZYiORv2zo2pfzCvsiKwNChbxY82Be
WvYUB9XbIvcQ+tQHig7EU8mGhrHE/Rb0/w61IXr6VYPhbGclOH53c7HYPeEyEZCK
Xo1E3E23trIST5/gO09d1nqBlaZMjROUhGlTrNofQVayUj7sDny1N+VfjtoW+WAX
48Y9JlUJsUyv8uYNNxnLR2dTo7MyaTYYKzEVr7IyA6tr/VmRaFHOQiaectzQLaQi
WR8bBrGq2eT6wP9fShanxkKWoBlIXGAkLlwvRtexTBMpLrn8a6ccGUpFFjjX83TK
CMRy7RsDAnoZi8K+c1i4q47q+J2AHZXGcBej1Am3o+Yx+HgYASt9Xw9dHB8qH5Br
b2AgBvt2I5lMUCkkN6aiyklBHWtQCPOUHZrZblHyE7zLiDX7YbpdS5aibo2b7MWL
M6fXH2RHiFoMe9x15nRA/+yWevq0pW6UZQzB/yBy+ohnV5gRh5l0p2DQCE5GFhAw
RJH43PtV/EujlVIby8S6wgLSILkqeTl96wd5TLJmduMrj0+Nmt4LYTKtC4f5B92D
zPCuvqLnnnEshvQjiCgPWOikvSSvmQo+aOaRzZxRIZ1ftFGpCLD18RRLIHBBw412
TAbWcmxHCQajNw+6cCFbffCgxTxoWlYtynEoEkSnWC7MYv0Zph7YtAoa26TPDWKa
oKpeAQuRb3GiNXzuKlR2eccItoRHpjxI1DMQ7ItdPhDOUTsZABPEIEgp0PePQQeH
1zwIQwN4Qi2QeYHDcWujhPiu8BTufReUym55B2HLTltzEw4c4GKXtDra+krWG5KM
LJvPhqzDJV8IuiTTNj/6PjO5vFIolIAq3gV3krkD6GedEF2xCaZtEtXe6KUqK6Rm
+PBNvQnaBbd6iOQV72b0qJcHEHYxTNVs0+n+tR7XfBqT7/GvRCYHzd18d5Ldsemo
JuTHhn57QD13zhc2GOqL3FR1/nD++yJHDW+YYMo+m2skrUH6IqWbIHX8mEra/g8B
jpjTgtvctogPkOKNK3gc30elLuI3TVdEP1Xjhhq67AESt9hbQx6XfYZ8RKpwdkl1
hGulI3LmfJ9DlQeZNnVq9MjF8SthtPB0YMizTVqA749g6WxGaz/c6hLFHpnu/Kpy
BfwbCCsCYU6Q6Ca0cufxvGzEDQUsmQqF7sNAMj+vh8sHe4AWi+8Q6zWI/lWffv1u
kCdK50iKDbLsMEO/768nv2tc+i7u8atJZnNhzSKpFKkuqIPNNKYMnN0M88HlEESH
AwYanKGT7gPW1BWt/d2FjjmPwV4+OICmDxteCf5snz5TPaqAjnMOBYEImJyuNuF9
GWAcbg1d8N6SSi/LMbAfju2bLrRkx3cGcBPQvRs2ZhMidwMCXqmeUl1TrW0+taRo
9ERc1Z0JEg4KyKPaDRAunJtZYzVG89N06RcI3aXjDcwg8t1JSEGINlFss8jfF+E3
19ddHrg/UPRDn0oS5cKkz6GvblP/iFY7S1uI/PZ+zZqRq2zShSaM6imgU2g3Wkrf
fIOTnl/TuiJtr1eI8dXc+5X1UvpcrhQ6yAKy/DeaXAa0mm7J9MP26xNs2MO245C4
2o2S/5h+U7wyrVd4BZEkBsWsbrRhKoz0JWBGo89M3tTOzGjkHucH2D4G4Pm3o3eS
Fns2E/BWfKcyQ0EFlKx79W5A2eNxUVdZgOebpRveY1+XAXn5jjJ53Dlq6b+IkCwJ
nDCdQSij9uPsiXyjO4b11/4aN0ezDg/dHReJSdlw/odo2fIw+Z3kCSWp/PJqlv8X
+tAEPIzutRbgNgd2hkTDV/ZpzPnDQjUucJrDR0iIT6MZUL7LvBnAneTVPNdUcFTn
cm37vk49SVTL7v/rKdl5mu184KhNMrYWTICrrRgpg9VcyrWblg0kB5+D8ZJM3wel
DYUJvGEJCoIZLDTwdkRfPRZNUoacfuGzpdQprVEAnm5VCZldO/wYyRlRn9MTfrnk
+5ALaB7lT4p9cwoZooZyluaEDi9wKZDQDFreIcE/8hbnjDFI0Xcth89UMvJTswhq
NJ4r0iZA7mqpKhhp0NMABMvy8CwWn65NzeswC9qpmCqS61FqreRjmp1qHgqxMNZn
xr2FoVUr8Nev6pmhlMev4EeyJkhz5HAnxKChEU4Gt4dUQxYDrlv+/JJj1+3AUbZm
sY5dzpEtsDcb3pDB4hViJoTBCA1irmQubiVkXmtTyFyDqVtYDxP9u4enxVeP5hRO
exHQs7S5G0XmdQmOoB9M0dgfPqni5w/AYLeBhkbU2h8q03kvVTQPao0lUNv/NPDq
eo/GXg6kf/HP6aRWWbINebQyFuEyf5y/Gai7YcHFaEB9l19Padk+9RCOjucg5ID4
V0TjDbzcwU1aPPXZuM8QiWoyCcFdcY14nU7fMvIxWBaZCq3edmI9s9fqI5L+qGcX
IlH0463JKXvyJqUO77p2OgNE7Oav/8vHwSobrFYCSimICYwMkH0dooBak9rxRqAC
w1S3HoX7Z1LwZFffMcuIvtg3aC6zfCwxQab8yyBI+0BakZEgpJl7QOyNiMNNpV1D
4SHRYNWqrsyxF7pAdVILGpnOoQrpkdnprnCVWLDyVNoMQKd1N84WKsQAZ3vfZJiA
O3D062L8gbqQ07MSZzol3Z6CfUc6h3tLSjN974T5yGKvOBPo4nLDxwnSkTWsa7w0
gOJRYUZaJ0s85myI/+UMdMOFEUMUEU7CAYIvISrxrWgowQDd6V0eoFFYR8hTuuRL
lPdE/4DsSXKyCRWnVbgPpeBZeKYtxsJR2xw8UbocjNiEnN7YMVf76J+gRaKWBihF
5XFHnu4WKk9RuyIo3rVFwFr2zw6zuCMbjYoOZWUv3KADFjKDdwUHD3IFWZmwwL7t
zjHsraKdv1gPe6dobL46Js6Dugf1zvbBllgjwFvOO6QX6ozXqSvjp5Bxgfa+/bxF
MWk+r4r/JtW2MkcddQW60lLC09levKDNHDol3TjfGVJjyni10gMrKWey11Txl5TO
zwj+zCMeG4mkhGmtIHObAkIvdGAlihIsydmT9SYzBDGh0gI49I9KgvMeGWA3NQUL
8aOll/mqiBJzQa/h6Hc/1LKIFT8CoeTrWlh74bBVSq41jkYN/RANxoGjGp4b1V/F
+Y/A2OKHj1bX5OCfv2IL4pany13qAZxqc9KW2ATWNkdER4o0bS0N0v3C6uUVb2Fb
SIH6QJByzrJIm9fNrD90AW/VQPX2DwyBsiVIyVPTDBgNBZU9j8afv0n8THx7HXFq
G2Drwx3Emawqou24yYIJV2ErK2R+SjMct0oNLyY9/44dXfKBwyx/hBqMY/9lYRM5
e4w44j+5SSEk9VsEewvBrnSDHxASFbqj/64/rFBqxbFhWxnNMX7qH08GmEwZ6UbA
v0hj0YUEQCUM2S5I8lFtPo/FND2+9ZwTf0fqgqQO/nOHsi7LEaRzEiKsBJTCs6r/
EzioEYIwklDav/mcZIRJnxpYsjVjOEtzJF/K0Fb/5zJ03nMp+H33pR4OSNeCWx+5
tscZtLp1pUy3F9gAG7xh2VCcUxuEVfINhbit/Gx5WVB8Dmgc8ihH2sv4bGBmITN9
P0SEL07R5N77mb9zo0vId32uxwCQZklwM+rd+M8r1/cGg7dufjhzrhRkEnGSHmL2
YIVCY1ZV7hHP0FwRCUbWExx/5VqaucwLikiKkzQhXKY44YD5EQfhotAggJQmHLCU
KF/LpWcjWcPf/Y2rqWcNWEb8mjykCKs2k9OmlSJfrQE05JJk44TyrJ7d5MnTMqHN
ewYAWeMtUU8KUrAy2wqkfWqBgj09Ui4iViUWAyQDHcO+82LdE1qr4zBcB+Fx2Ca0
/+WAanCPrEwXGFWdOUUcXAvlIRJGcMh/+/+hu8H82PLioHV8u6pK24QkHXTZmPU/
eDF0ujuvLaO7tF9XVW1h9/QLQ9qrtREnes/YiLHX+eR7rZ6PC5yCj39gkluJ0I9+
VHoR52XD4b0H2Fy8nfIh92EjW5rcwCSfdCspSLyePVE7ZlTfBBBDjKWq0xZ27hlF
0ILLl6Z99nBASjQLRQEVvUYsstHQOTcLgEF/0IwlDkCE8QNQ/KagsV9Eg93KBcQk
EKNsPsGJZge7X6mLschssDES4CdHigvigJh5UnUR/gB+dDWdaaIX3j+A4iP/Ny7S
bhpfBz7iI5CwMhmgBlfUqm7G/6uoYJ7jKOMU8mdIxaX5HnnDwrpUtoOEWYvQWLyj
DxQiRVEMxj68walvXbhkZmTgGFW6LFmZUOyFYD+XT/t27I776A/EDd5yCUaKHBiz
G8l3mNtOZRU8wg0ur3C3J0Lrw2zDIAjqGJe+U2mFRBrwM5Zzz8HLfp30bl5/cf91
/sK2GfvMSBy5/ra35U5k7RNTFpBTGJct4EjyJTLcV608jKDgwP0FyEF3vISsGhEW
l89h+DWlIgrdd5I0xUSgtz1eEbjTzSrAF29B+e5EQUNbLUZc7BtnZTIvXfZJFDNd
3oi+wXOKLlZqDq85AUjFep8pjXIm1IFUz5HekMRcmmfaEHqjFxZnQsbQghxyQwJR
sTe5LZZpYFYbvMCeBTrDok26+SIhfjv0Td3zCy5zqC05DmpPcnmmxGNYugHnYRBn
l/k28Eqv+7zqyZhkZeJLr6S7lVlOZBIJB3PeYArkOKozRpzyTXyuzvXvPoXw6bRA
FS2HQ4SbQY5dDgvuenqMZmypiGOHmu3BPPqBfhWYsOyY/6WcxoRsr6ro/2Km9ozr
cH1A1CVI3q7+wR75JXVKMWqi2L50uQuJQ07Ht6AWi4itfPahUXHaq9ODDVH9J1jq
WDNMY5L1ZAMwH/Z3LByr77D//GXTBt2ycTkTkZ6rL5XrIqmqV9HD6vW/rKMSNCtw
txygbQvmfxdKMd+ynEWa03H37a+DpVCJhqlo8753fSmmoeLw43Nak+D+cCG15bqF
vt7xhbAk4SCc79W9Ds8ElMZ8VidVwYO3FYDnwere6E/gAeJKyet+Qw8HgxrERZU6
cb/SCIsQd3X4jH8Y7ZkFITeCs9yRLa1K+x7r5txCgVm53e1QLARScaQzu5fHKndN
dErhWd57sXTYnAdLY2pB3brp+3kvk9JW/DfuOoEgrjyJlEPxQ41SyCFD2TFPbd8L
OjDNRnYaD05nkragcM5l2SJ2H7GOxwk2r87+UyJS+HqdbkWebCgV4Aate2VqHiIL
q4KNePCddZwkIn2kZX3BWOMUmtKVAKQHmK5f0B8sAU/MRXlCX3SC8sbVI/KlbHBD
Sn3V82cyIAe3mRJ1KUg67auCqFx9ygnCvO3EQdmoLjtGZOpT6NK0Ag3r+/qldTey
uWPkW/7Tvx3/zG3GZj/NHRgXeyN0+jiuB8RFPdIKZoN3mk0ko1KXOnoRLVMOTNL4
4do2tR6smn31GHJYKuQ/wSLuFcYeQ1rOeJJYMpEg0xggmzpznVvUofxf0njP5C/l
pvxKisK+4h0YdezRwpFuj5d/wv/FUkr0HnTUF4dWG+NWqwSZ05XqW6uB2jSlBIY0
0+s821TyrBDG8gSg8aeAmnT0cyfLntx0CDtf3AJxl2APhOK/X7LOCBdo+toj2xgr
idgve2cQHlbZq/jlaO5OO1fPtPWb/64zzUPsDg4fWm89MJriy6lFxdRK4c1xZXHy
VI7VTZ9Aon+XH7NwVRRGP1wPpmZ4MOk9BXv2mUDIyVKjCq1atYL+o9pRKsgrsOtP
m96JFYEn6tvUxdh6IieRzm51h2WSdYD41cXbIID4NuiN9Kb8lpRNHDRf9WP66lu+
e/U4jBCT3PGFwGbeTQuxWWX6JlG3FigBXrP+HGij2fkaAw2ZSIYj+dolBrw9W6A0
mVAzvhBYRALTXptrkY4uwI1EdshRZc4ir7NBY+RzHUoDxjBkx33UJ4xNPPF6GU/9
4Zsp5M9q2vBm07R4UKTGZEZ/MyjAsdU634pRKTje8zkyXFNvqTNfkgYI3T19MJmC
mWs1wvZPcN1Phckl7bcmCcA4OEKACJfJ/LOo1Opc07jw4zRpVG68KDMSlbsjVXpR
z2m54C1HmvvjFPYx/fgXZdqMeqO0C679OYBKLUwW7phnN1EG21iuuJ7ZrmiZLDx2
1Yv4pioR404T9rFIYoakCHnAYvBQVuOOYuNiOQCWc9NGGN3K7pw6aQTXj8Nm/r7F
9Em8CTLSMLNF0kAqbwsrdV8bz4ue8kh+Y4cBvHVLVgbLVrTSHowMy1aEVYPmMhVL
IsU85/r4fOLNHRWuBcRCjpafAMIPAfVP5lLPMIdAR6QDIjACM1sgfNq5e9Hr/fJj
pOHCZP2SNtRMuEXt1QKFfoAKGk1/AnagDGTSd+JutprW5ERnnxYSTz5dpmPqK2R4
g6n4dy0RZEMC2BkbXizoI6CN+mN6JxA9+7W53fnPr/FX+im3HiBq+JuER95KrT43
jVXoMnCAJoXfAvewy0BxUyA7yf5Sp2F01wV0iML7WNHf8KdUhb0X1QGXA8cSV4aU
G7biAf+bnoRGUiD5fyTg+aO0DR/hcObicwgwHaqZdMlGK1YJFUOoQLYWk7ozB2z7
sUW9UC0gJ2JnEvuk2+49dhRWP+WV+WVYdkFp0weZg2mTYZ8tR0M/pSJi6NxHzPXJ
S0uaUrp6SHDfAkEsZeN6qkRyPpAOErqRG9athEkxcaSH09maRTG9gkJwZh0YsR5P
uuK6xTVwvWOPJhDEEypW+PGEN9UuOEAxa7V3zw6syQEEYSe6wB973rEzuJSAE5gC
EsKrlBL3d/I8G1YKtARiO9I+rHr74af3ASvTjvE/NynXHc99N76AVPgOb7UhhXvQ
CKjWJFR2TlvQ77fqU20L5Ho53i2AmfOK7iRElFrJchGV963w9DlUOdOLBOG5wBwP
1m/RPtielBM4UEOyhKtkOwmtkkA+gJqoRQzIaDUFk2iHvfLxm/zy8OuMDApS7JCr
4gJgA2EmXm+87NqYiGhZVsfFEYmModglrYrvAWxiIbNFahLXhaL2f9MzDHcKl2Z9
Ozp8Y8jIntBftgvw+9GEcyrD2QucvCsJMZkt+xxRyjofDQWWkugSP2fmQG9RJfAX
DPtHFepEIQ4zY/TOFVA2PWDe2esFyj9Uqu4QkkJkmTe8dOs82H37L0ULN1AENAj2
hvrxpS4sXizSR8rkMbLJQbRznNWK304NEKRIJQZJQ4BcwvP/LxCzwdonadFXPWeT
sP3A5A/7IbwXEwor6W3tNY7eg/XuwDrkH8x5OIRDfsbOAm/tXMCRp8yp/EuFtFwF
1XWJK05Wl3YMAdP+ui+ZyvMuMBg4E+guW14FmK83+km8qinhwNmJSmOvs2df3dPC
ApFvVnkiqHRjIK88YS3a4dVTlBNmsz6LgRHcYGurm5vD/xrRdDfVn42+JisJ33gK
L/QfpX0OVFfZ2U6XN+NsBXSLikEnbe+nR/fKk1vpRsbvTdX8NcG35uFFIXuiVavR
MiUQqV9UnYIrXs7rrDnEtgo+pFEaGARfOAlE7l5eHni9PMNK3flpgJ/jjwPF9HPq
Ox+oy0HyDgyAhKNQKWMgCxGpzmH9ilmOr1KjuX2i40xSQwBY41aL0Uu+xTMRm0TQ
FpO76Jcvpqm4xxR3KknY3aOEOzvLVTR0/n498tSxW/Wvc6xSIt3idmApD2hE/CMX
hzxrF8DuJUlr1GmMR2h1EIl2xPg6xQPr0qs6Wd6XnMM3VHqwWQx1F3qqzcQG++GU
+aXe1LYjcj0BzRW+9M3d+Yq/yT7h2CQOtIU0BTlVP6X+W8bFr2IqGwh0rYmhNXoW
lIDJ+nK65CSh0yGTZDrOjlXai1SP0GHwjFvVkB4ICp68Qh7hCy6o5nMf2ezL3ooQ
2S9V/3OLXHvlCssgAqjBwvGn08RugbwInHqv7vJUL9q6k0+aV8nIdhdzbevMfKM7
L9g+0ABFpLnWS6+5UJqz9jwIONks/xrAw0ne3tj5oEQB70+mnAEyw+eRBZ0fINbq
ymmV9alzydnusoQAmP6fQZSB0F0dJgeylFWQSpiyiZ6e3sNLtQsJOtJldhkiFFG2
A8ZLovMhyXijxDjUarFVA3qGFaWyrueuUuj/jgOeTSovrjJMbOc8s5vo11FvmENN
WQC5Ayg0V4IWVCY1sCQohEWXwn9C6d3YFA4D1j/RsBYTBxNFUyLWaCLo0ZD6Al7a
FmoRKVIbHuhr475Yz83AZVbGbu+Uob3P2iAUHfvE74ZbEYUd3sncdEUexYmut7lB
b7EhNpDzx3RdMnbcGDfWw94YRBLJ1io9lXV96uVaLStpoSh/atITSMWrpHfL0cID
qyGWxdQ/9+okQoEOobIIejvPvFr7CyXYBqxRksV2bZE3wvpkoXPghQ7oAizLB8HY
sbHdiIHCq3Zg9bpABDFbh9AD4snNUlhrGWdNRK078++m/t99uIGBtmVMKw7pICtp
TO81r3ceMTxbrFoYD+QX4SgkQQKfsGEv6wDTEyFf47qQxEexn0gOCJX5lJWyDk2T
CRIFFKnS+/FOaoro8T/nFBNT2X5smE1URYSLOeInxNTsNbEj/I4i6j833ekcVDB5
KcwrEq1LY95n2D2WWQIOZyTRkf7StNTB8yTRUfk7uS3U2d5DcSN/gHxblz8Wvk6Q
EhvHibcW53zyhaZH6vkElMK7CjrVYqoGMX+PTuGU00OsRDwRmOWcFTrTmSdz2Ob+
TfhJswqP0eUEGgnlKTDPkKilCkEejzZZDhzMIpR5DA5hQ7VQ/O0ILTvvg+PB2EQB
Dg8PsfyBQPI5Xh+tzFvlM8YLa7LBb9AKW2mqbjosvjlwQ2svH1vegSBz5RD/qfac
Wxvs/lNLg+m6dkRyYixwMKETX4rUWOI24wfMacmK0p23ViMpw9Er0+HlwtWZs+VJ
GT6JMymG9FVqhj98eXJTl/GiNLUuD+7OS9fsNWL+qOi06N4WPMyjFGdfJVuvIIhP
aFhnXrq6T3Faa0g+Hs5ytIs3D3sX9LWAkibbwpwdb2QuDRZKo8A0ssqYpR8VWoOG
YoVhzC5mp5MHf511dF3DrpgTDlRVTLUzXJoyyormKkd/8kIFRgENAx7qtJpm2P9e
nv0wHvYZSJ2byZ8aIRlOvGI+QvQhpg5y4FIYS3sYIIffXsx3Bzj3moZlgWUaydAl
e1bNEOTstuk0g7C7JfXm+n+YXkO9fqXHZiqz1hspq7Mp69/CwWbHDtNXxOyFtre+
eDtyMo3X284Z35RW7TbwDgiN9WqtCPEcrEmZVha3KlVoqcAFEYeZK1ZjBsrI4ZOF
fYCLmdxe5MmLddB9+82twUDzx6GE9vuueChqTd5lf0sK3VNuHK1fFOYrGEpvPUZ3
qPfmtt5iPMRwCyMeBCScH8ycUQ6Q+25Rm0FtH8xyva5GVBmDTniidpdiIpujKAmO
puaE4oYZAq9K4aMHti/riwuYqrDMBLgi+RZoJTj4itqndPfZerKlrSKHe3arslf1
yBIFebIXxW1SmxjT6ULiKtIK2YY8PwHfpqhK35HxZojolFokd4fSrHdYAU2JCx/Z
42cHeKzm/Q8Qbf2ZKn4YgO5gmSvNuerL7Jgzvb2HGZ/7kGbiLSM0RfxHV3qp+WYK
5hThF59YTSqc8Kw3+z9vE6RztNPf32rktt3WuPsQ6afHcbzt5FPvyPFDrrkR0++t
9O3msOIuiggNYls4qNlio+px/kPXQdRRGn+QpuPnA+eg+99lYehVD9MgbPH1xhe2
OIml6QdddCeGVIyZZWFTK8xEk7AH3YrcJYIDn64CFc7ixt26QRNCEu57zDjCRaS/
XP3cGMqrV6dqXP3CVAkoIdidbO1DRU9Vwul2VEwaeeqY43nK3WTlCW5N5qnSUwoR
keEJYWer/EQQaUjclsrt2MliS/8J+UfPZyEV/PyRoUjGbeWHQ3ze5Mf+06WvmsMz
RdQ94IuIOfPpcbDmkzG6jpPp5oOJZ/YW2tNtERvq4hXKgU4asPjDcP8GFZyeNsOH
qE6VshG6Rm7qO0QGQExQ3C9W64lxznUHWg5I/LqCP5OmbnA7hJhjmS1l8QE+uWMK
5qCSYV1blDvBdKttokczYShLMnc2xk+TEh2ukmnAxumX/M7CDoqmAbg/VKEIu0UA
3oT5LzvlNb2HPRX6XVABRsSHXkbXmna/NZL8pUXVUf0dlAlwTh9h9gS6F7zAMR1j
7QDwqR0cikmpWbSdJO0+3LMmOVBEMv3kudOPEpH+wmA95EuTHJAn0wMqeGgneThK
HYm0tmaTcLoTEaUcA3Gh8oKF+sljCJgu/JPNV6eHPVjhI57/1323mI3MIuo29QZo
LjnJWCyjXzLZp82dugnXaTiWtFITDKFTRx/J5pIVgtxBxmnLRN9l9SvdMbaRJoyQ
IAy9iGwqyBJGSOLVIqeRJT4uRgl5UewHoeslcqv/ln4RILEe4Po5yO4Rq/0Wg/a1
4h8JGcvj3rPaw4/mAkM2ie8fBrpx6nzhnfYVNK55DHXySiCaF/+qqWDdWCWj4pl6
Uu5UqonwuuqE2KUwlC2AHVTgn9iPD6EppN/k4+SDuD/ngkyjZO4eUFNZUNNdjk6F
hTmxLV752WbjFR1kr7OdgBWvdmbpdwn3vo9bkD8B7+7Sy6wDwx3uX6svbBP9ehIh
xD3Siu26+Ui5qExIsS2/3FGqP1r6xXN2oZVG8M4V3hIRH0kAfreOXEBk7L2z58JE
2JgqqEZ0NSHrkcLLK389uKF0ygUEz8D1uWWtKcJ45uGqDw0im3z+6WX2xMaCg60v
pl7lQUoVMcYdQHmU8YZG87/dJaOtwdNoIVylEiMmrhpcvHeGvu8Hi/qETlnLd/7o
/ZaJkPO1QKMBEGmYz3QUllIokdlTSsqR9P03zPc2kqUsO31v8qitqZZdEsWKeEk1
q9YVV1VBimFbRXFiKtzbh8WXcnFq9BeHBDgcg0YxfnvimRxQ/XFGMrjtEZPhaFZl
e8AT5ikamQcpYKL9o7W72BQIwDvTGh1nuvpGmlTQ0rCTo6cyPc2zWXcGGhD+xgk6
Crd1CDZtBBHMxF1lvd4ddq0o4oQZftZdyXziaXjsKcOZBj+OrDuv1jUP68e2iO33
v2PDZ4Y2UrAvPTZ1pR7AlJC6SioE/+EqtaVr6F6rjWji+C4Hp5Zh9z3v13OvEBBg
VRuw8pgVrLBirMNnIBxZr2VFG/cKTgi3yARyfMa1HNaLyKPO8xXLanT642FThbZn
wwpYgqm4Y5tZd7cn4LjiyXZCMG4qhb9TqB6h+ZNwW47WYIiC+ct3eoxItkDhgxfI
7gp3jcQXD1Bbkzf1/JSqN+SHWx77l/9600YubErhqasi8Eld0hyIj9ndH6MJK6af
B4c8EqvOHhb0AI0sCgM6dgBUug8c8YVXqTsWJugXY4SvhpEl6TAt3w4g8Hb+xcpD
9lFYy8GInkSaoRYGtQJO0r4iGY7Gge/trq6JVjJF9q4Tg782aoMIt79f/A4nqlls
mbcnMWr6HJYWpJVgiUmazZm8d9KvtzV+fneB3HvOejPPdkqlJWrJu3HNPcfvRydR
kQcBh7NIkNo12+ZrPyXFwwzGEUQS8OQgmRIkKF4orFGkHvR3vGynxCOOPOHD5QmP
YSkc+MTk5u57IQg4/zYPo0PGTpOGg8jEHxAJl1QodxVWb2ZZPl8RV7qpzpzWdbIs
UQMyt3PaCMoXf2U/ibw648kXtH1lE/sAwngQQw5OhMVY/ri3PhxTwh/9J16KWaFC
qXny4cgVHIjG2XE0QoCcBvH76BnsCWkoxaJCQjEqZ9drZXsn+dMl5XjjPXXk4aJO
ROTjaxrkUwegEMWR5MnNgpHf7afvzJe2fL5ZzomG8j21Zt6j3Idh8oyPotldrbIA
btay+goqB2PWsebmUDOm985n3RUwzZjwCPyMjnQ+8wFm6Dvig3M56UyL2Ok+njuN
coL8jD3aKQafIS3wob32RTnMaUZVXs4l/8G2p4jrxJDuY8SxmVILuczKvDFeAzuO
TRclRZS5Qek/JgDw+QwxWuS12f6EORxoA6Z/H/G/pzlEKB3dAgMYvshIYm+E/Q34
wf8L6AX8gHfLXM57cpVZZ5AqTqtJyLvAZ+p48PZSfbMxnpRaOepGlz8P005Eyjt8
rK3pkvHVlmuOdq5Ht2Vx2H6uFLNGwJrEn6wrYn6LOuUqzkzCwEUqAmfgGQOqx0WO
hKAqGdP4v6kAP4pKJGti6T1kBi61m7oH86bfIuDrmSqiL5+cf9i7uX9j1S710ClO
ykzHyG+lCM0bc29ndutfVPWhMq1ZvlgevKExkwqLZ7+dRkdwLBY69V87F5k8Qmf9
liGWTpcod+DvPgsQn97iyc5AKi01P5xiFXhi0Wr4RdEMvTPYlEVh5fEsTeVHCMnA
AZ/R00QGsMD70Cl6xBXrRf17yjHABXWKsBm3kYJmscTS9NHcjXjcuy/coBBA57oZ
QvJIEYMhk0tN4MomJPylKyUyl5bjk4NnZ46U6L4mP0BG6zxZIx0igdrmCKMpCgV5
k2tcZwD9TO3/NNZ0feBkC7d+n7DCcjunERkluQAdZF7jY5DQJtWtgqUyxwgYSlVS
zi/8qEPXDVgzL6mifFW6K63QQwvIX/ngO9iGHxZkK23QDYmgpjjILCUAU16PV9wz
+F2BsfNzCFDXb0CIj7u0lruHYeq7i3/y57cTQx19p/JJdfAXZqxn0YqSHfqElyHs
djlZLNQjBzk8bchT1U5S6jDATgnpwKXAq17nIgdo2ZRhMfPazb623hidPEfN8VAT
RPPt4ogAmhN8WL3EiOJFV5WDKLV0PCu/dezutA4M6Hc9uDkgesf041iDz/YoX8W3
zCue+NJYHYUEXLCxtiCIqL3Hlsi3jugYTV9jkCEtA89is5xB5yXGubzizmhmI/dA
RR1qxHMOMkTU1VXQG+6PRsb5rvsH+wwNK/KJWdEIpzR6DRKSZAtK++uVGhbEpO/i
SMTag6EeKZAxD6PvwmLdsle24lnzE0g1YSRcEy9ceibLtX9xwgxF1BygAPaVDgMQ
oR0rnh2MgDBbxQ7XEKodGDzphQWjDOXywQ9VWBp5UThCv+U4kQ68BnXMIP0RtRMb
X44lxrwTE7AKERH0RlIpmo1ifyoe/8URko/0h+ISqmDfmR8kC87K9i6npBTn3ffY
nb3bi+nfFgMda40ciuMKLMhH2KDtsmH2UCijn5wd/vMvD+ebN2qqkpjC6CIRT9Jq
SAYQrWC2tpxi18U7m/sApMM32k1Ae4FOQhGzfwq8D0aDKtiGgjaHfTx3EJNkXIcX
3Tk/K74gVLTxvKnEOxc+Ys96We79ieC1JapMSAw1C7Ng2CpKnKGbNW4MLf5huUoQ
szA+McDQ7jRLVYCvvabGdAstikgTFHErSPeqlfw77cqB9i9NBGTBLrOHcakyBRGu
ymzLF66nkdtHQWUI/tcq5Lw8GXjGOY2RCBGepSD1AvpUikYcU/4WOU1K8JqtKcuY
0UV+kpyHkG75rU6MHq8aH1TaXfaE7qF50y4+AIvLEHZ9xItkEh7M6AsWYCrt16ce
NVj5r6ddqtYJL4Rx875GPICdxCIqpZB7cHCRNnQH6VH6ZGXNYWOByE0xUn9THZ/D
g+8eGur1maPvZO6iPaKapcyK+1EdwqzcEn+PLx0uNtpwvzkQTHwAQIaq7F+Vg/2Z
5+cTwNWqKtxwPGzT+lmi8Db7YTs5bIbFEfZHBaAx1NYA/+nF+y8rXUdfzms+9aoQ
2FLuAODRJUskLP/+v2Ej+pPYlc6rqF+9WuH25eLLrJjZTIF1Wzhk1iUhqeZ7YFgL
ZcBlYWhr4oUQk7oYxXFb2dA26Dz0ZH+5eZcTPdsJyKOZRWj/O9cbqKuymeevgnPp
UhFhRKVzgcGplWQazGzJPfdE70MWHHYPl+sJHY1JXuG38q7aPHY7ZrUGuxArbXir
J6j7LeqcC+Dy4Z38WJs33QObgNSlWSNHD3S735giVHJ/qSUmESsWYENxldFO7JRY
CrXstXwWpIas2g4hq9ED45ySndSSudEOBn+26JGADBX06VGbdNfZY+4bdsQ/O1eB
uPb92P2IwgHDa/WZACUbJ5A6e3GTvwk/rsNTG+Jvh8hllleqFMzv5ldkQAJs43Vr
w11Za0hYeXQKgoWzUb52feHtjThJxENoxEVwTckH23HNj/8MoZlt+TxXCtAZ3B8x
dCs6/2+MvEACDGjJwHyKbtIaTK9zwXCnl22Cl8KNYIgZqh4udmvK8jmDw7aKQ+fC
/FBt1BFWC2ZumP9vynx029mFntJgDvb5eOYal5IqTls+4h5Ebs3wLsDFGN1j94kr
7AkMFQ1uD9fbtNJYlOz1UBl71v+SAQ1X5POehurq/kU+kF/ZzkGrsbIPcjwV7x1m
H2aN1Mzj6Gvh42+GeKmcp7HywaUE5G+gUrxXm7ETklrW3Pro/SgM3QIvoUAd+ftP
IyZk9LXYjvFRMPda9iMnYm9KFZEj+FrXjh4J++x9oJEJL4u554GgKe50+NeSJrwH
3APHpM3dpaWu7ziUOhdtKAhRYlLs0W3coN6MfTTKrO5asr+ZnHBn+0RN4XUqrKLh
vNmPdVcO/2WSFJFAoGWjxeBNxwaWU+8tTuEpbyx3S/c9Ng/vJCpsRhcP8B09r8r8
uI+HhtKWN5sueoXFOTB0nGHSTmEkgOs+Eso91fVi54xj5eivzE4yqZsdN+G6r6bi
8ovSbUfyxOCTeyRLvL0ltJtpPXiXKIS+khPJWQ3a2Z/VkBdDl3r66EMZZNoCZAg3
iOrtF/aSFcQ5JvGlmWBov0noYDIZuoe/dF5MK1jaER36lwIKv5VLecGSIN0Z/Q9S
IUQWWLOWd6+8/uzFWmVHsh5FSAbd11IAz46eemg73xNAAa9SbQoRddL/MZOvZ4wK
dlHGQUsRaMeSPR1HjznYfLNTey4W+/glEkIdZabMf264niBzWSOExPYFcftinUQ+
iwaW8RI3C25KyKVhHwoXqSK2ijU+ivu9/UnACxzafLh41d0xp/MwAQNjBz6KAiBH
sEtdbZ4GimwP8RyxYEF1uYLPOWb+FIUMccfbUeEwXylzDknogLjMPRH8Gdjr4v8s
mpTn96c+2udmps9qs6CQsi5A8MJufsOAJRpPWNb5Ws0Mc3IWkvTmZDQ+nwPpvuNU
ize2ZiPEQIfJ4WkaSR3wC6whey7mtGALBhCfWJ2WpW1769bJ2trA8fmBWbpR4MBR
94FoZ0QjwT6Ex/XdrhsWCY31d9RgJxgiXOiVs13+e6P0GNNaHMm8kuTtgtLAu93e
UhvrXfa2byZolP3I35aVl8xg0Ii2ulzkBrqZiUpEbNRMRp/qp2PS2ETUVcaVObaA
ZWO1KIFm2O5hUhpdGcD3UmM6FpbDTNnvyE1Nbt6zXhyQGE613JWaLcIjITztO9RC
TjDsUNL2bQ7YAQ74heEmc85+ODEzlNVtNqGF/9EF+yNABkl7Uv8QAfmXkPxkVD+5
fuwCamFjs3hH8dmIB9tiuVuyAnxduW7usvPNa6GorPgLZV/1tRNjAULCpe5BCHqI
WYNO1Ud/AT3QmnLWR+8HKGCfd/Q6oGjyd7VgbYd9zJ3pEPhKCzxn79yoU8qit/dP
WfRZ1OWzIP+IeNqumrvXT1eZODpkWqx6VyANqMDHjQUiCYY4CrSUma0Xai8Rzy4o
hNfIMa/mfF3aoE4OpECVYjS3YnrLFbQYdij4eITtu/tDCXYunMqUDVfIV7AFFd+n
s1TKmi712RTWzoF11QDVau82yXOIks+F0ulLc19ADnhDt+NFOojeQ+1Rap1a1CfS
KYi9Y6p9QpLlXad3OQFc9D24gKbIGI8adYqrlALxsCjac95NpeirUvUJf/Us+1BO
xZuVJzr2fDDQ5xLUETP/RhpbqfVuekeC0kQyu9D+pBadUjayV9tZdBDgcOCnlGj7
PiGJEeVXIXNz0GErBKmILRYxEfyrASWovxGSsz+o1ZCOa3h7xy7dM9QpW3s6C1PH
My+KXLexnQMIt0X6EHP7tPoW0KLlytG4de3F/5ltB+ajC4HIVcvI8Gvy7hlGPNcR
Xj9zvTRBc0pikkC5VDuhB7StfnaAga1lF//QYk9cKQKAxyByrAWyS4CYdhI0X+th
ooiE5mSEGgwe4h41cNWxsuROU+sf3ZZroszNy2oSLxx8paug844qOOK6d31MzsYZ
mcQDGXWMJOCewUcR2b6hxaQgQaIZEaEK69eqqJ0kJ7/S0UEjyHxLM38cwVdogkwa
h7V7AgLihY6AWn16rh2G1/dcy2kF8Kdzq3mOiw7QEj59XGztTXU9vBeUBezkQYPZ
Fi/OhVP9dzxL5S4ETRax9/OUD7+muVBFRmxXs0NTik39B92GTnqD2Oj+aixy1PG0
oVmXC9+lJwzxLpjY0o/1nwPOVxdQgsFWFOS7Q7oVHNOW5U8xr8549jdiIzXt0ev2
a1pBEkkeSOhmtir9/O37MUAwseSWQvu5DJexTQYeuadbyrzSZL2LUF4Wz8a0QwEn
//Q5N9qVToKcdbJ71xMx4z2wODwQXpAimLeqrkMlGSXmORrtKR+pqyF99m8GG8of
dXNb9iopgn7PX3yX4HgYOqJfSbcKnP7xPESGsTjfHsARqgHW4pKQfKLK1pZyh/Gw
Ni657FZH5aNw6pr5KYSvcS0Lslu6pd0K8ouY75vo5Vb/12fQTHDBHBJCvtMeq8Ia
AZ1UIgbbxseQIHVzSr5OQqLh22cw4hxRfYsHh0/O4Bi57OxYhopTMPm4JDY3LD4t
wHy6IPqA7GSDHv3RnbqYqAbN97QdEkof+ZpXWFC6wkIJts7wsw2W3V2TJni78BOO
olzqEqf12j8TjgE2f0E0E+zpD3TXxyOmUt3watkml9C+cRBHiDwyYsS7tSkBLHlW
fuB/ecJ1/WpBd/CRXSmxIYQFZHq7IOBr+tkIo18TDLzaRK4pmGGUQjSdRsygT/vw
6ahtwGo4QR+oJXyYCzDFuC1d9dzVYFKBXm1wH5frpFIhjWn0PWuuW3NNGz+vMLy3
445OrrFRTEXkDYJ6+Me3g8DGAsomX6ShLeJdJZw1GMjIMRhGdrCYCPQLvgRRoslg
eqh/M4bfNT2dfNU8ryFP3TeHLGxNVZJ7UHhWY0W3RdT1L9/O6nN9CvcDuA0HX2Sy
gXFebnoHQ4fxX3zYkIFKoMv57D/BK2vqT8jwV93+IPWm1z3aEANZDa8dELiBDrkc
wxVHhPakIr1DZChjC1HkJ8XuaroBvGEuUptvU901AVsfVpQt+A021KpVTawmIVcG
Ma6Ma66x7T1WWa+aPEqRYHlFzIf373I2SUv5iMGemwaG+MpSAklbHXoA1/UbhMYA
QOilwwF/6e/1ltDqKcoHeb7hVeJ+3zqRYe2ifgqUM9dzmzi4YHtQFI0XfSMzqqVl
qZNslUxdLSBhTkHrAdJAF1evkd7j9Aqc2y5a+guIED5Dse873VBqi1tZZan+wdX5
JIyHhiPR7ED17QHSZkRisAKLKcSqbeuDL3kHGYpuxm9L5ttxDsCjA1w0zcvuwUL6
QidD6GInCkcQbIu5hUdeqRJXEL58W0NUGhE6lZUsV6wbI9CFI74NwO5q9m6BF0Fw
Ym5JQW7Efo4qXmouNPyhTfg/+bs4vpYn5Kvt9x153rognb3Ucg3UYZl1oJUZ2NKw
hETTrRWV30fQGX0b/jKkVOxV/iykx5eCGQp8Xe2D4jTR3/BqGLiAy4memAL1Y6SN
uBaZsD4iU7CjAL2rmTOoo8K3+UTVfDAkvk5rqPBATiEd/VylwE6l/2KM0/NOEilQ
IDF9cFAI9hr0KargYRs8Fv2OoKWaP6v97heIDKicfq4wM8z/vqdfcYl2dlyYnvjn
kbB93Qo9ixMhtVtEv7VbuHUbt9O4BkCO72UA1M5wYmLXuj2etNsuli40evNVYSO4
YeAHvH2bNtV8EM7Hf6euqURZDj+2CQdT6uknO1lAXRc7ltclrLfhhAYtvD9Eg0Wz
8YmijAq5M1yKSr127Ep5403QrV45Vo+Y3ujwY/F2axeWWv4l3aYsuQwRvno2Cdfu
HgLXwxyWgonw7DfK+mhiPceS1bXZQI+enCIU0GvMf01DsLNpV9Fg7zLE35oewZTS
V7TPJAPwBpcH+wH8gxvs7JBVKS4ld/SsXZj5MlZsc9ifbOZ2JZg7Zw7hEgt3c8v/
sa7aO3qULJ6MJxeSl9+cp7rf9iObxEGPUiay9mp0OL8Ye2Xb6Qux+W0Kauj+0KHI
IKuPl+RSrUqiOrD21UsrvALjJBsIWVHpHhEKraSDmTLDxztMP4GOHdxYJBRok1cx
eCKlLzZOtcdzqni9xT1EeClESAlD85fZuaj4xT4bb2lnOs8n69RQBa55hfpL0EJ6
I4nVS5+bxOevCh5YJCY/LkXUyljfslurvgOfn6YrDobrV9GJbolJ5pHhtaUTv+UZ
xpRXb5yZ9Qlk6UKUsOSyWE7WDCEFxgKPR0FXLWha3bwtte8dlrZAT/jv1caeQk5x
BXqusMaszI+tw7hmR+3ugKuk553Tit8805+e7QSje7ZduboXM7SghwngBeDJwkgP
Kn6WLCT1OHKhJyFwKx80rV4S9dvHPo6rxJLad/bWLkIepk0KLCPw0GRmND8qXDWu
S9UN28PScMhbgEZ0efJ1MASRN42ChLJeCrPZMYQZm4IuwJ1TJmt3746vvvn3Ayuv
h/9KVRZZtJihZHShZizsO1TP+Q0wl/QWCAcq4LrT2IA8WhSQQqzTXubakezMWCPN
SGtlz+9r0tWR0SGKdjNVLX5o0ZUHukqtPxpQRsF7DWA+03LX10hqgQn+JgHhgg0g
6kqm0LodvHAXJiuM+cNLPrHdwLpl4rQVkGkJAinr+7rE17OFuDtf/uf+jyjxC2uA
KYs5/eR5mRbcDD0v9WW0P9cJ1+ksdJ8sZqsk+Jh1LnRpTZPBRNNFCGpB0UP2s7c0
a9SgX3lG3TMJWLM64rDyVnOm/N+lpFweU2iyhttfJDnmZ5gqRvBXXPjEACW/TK2e
lTFwdaUlcZRxdolLl83/2lTtVl5FXqszrT2bILAXVnD4S4L9HdMa3irElkxPLCPv
vuPMXii0cHi9lh9b6MLYnbg/8kCzLb//LdexMwSb9FyXNxGzD++AN7c99jAQT+wy
QcQFFZ6B7PXo5IzQ5IhYtpGgqEE0anmGy652fS26hwq5P3YiecK3iRKtr/rTMbi/
BKscfQjwB1hmXxomQQdwB+azbKdo2GVCAq+Rf2NUrC7nmWJ8uKu3SP2IlQlfd41y
Y9JgdVL47AhyrUl0nqRtq5ik/99kNjrDr7ORpF2BSOI6CZRDP1oYNBf7JSaZnvOg
rWSz/esurj6bKkqHMmiNoKPRKAQn2qwORWueFPU0N5celbo15LAhVIFCg2qiEiwO
0FOKGoh1xZPRVBi5Z9nfjnq1tyAonhpTo9NzjTfLh/iwpI0T11ISbrPZZ03fcH4S
52Tg6RO7E2IeCEMUcZdUHabkZ2Dy4ielqCyqiEJcPAMH8evZTp9qDLDtHGkPODio
weT8rxB2ca1zEudxu3aevBlhV/6AxeH2+o59412EfRCq16wZqnfntF2oCOCqt5Hq
upknHDlDs5hKCCRI0Rne6m6Trn8AefTMMAgBSWiXnsJMc31y8hg+etkYblT4fXUF
Zex2Grk1iRhlJZqolC0oJuiXFL4MIgp3oO5k+yh3PYVS4Vl7jZtga8Rf8V/EggoW
WaUyLjZQZtbcDDhHEydtnFNVsk7aDWwL1zujI7Z8qcLi3dNRjFMY/in6U14YO5V7
x59Llb3VLcUyGTHTMrLIKkzF7o7aXqHvom9VQTjllboV4iWqj4fs9hriWoJN839v
XtaeAca0anSSqSop5E+EkAZUsOQVqGn52jIOVlBV4BdoUDbQvvO4nP8yGSaFARCM
Z/GNrCalVkm8lg2G90qNsP9D5rgt8EcW1qH3QXkiF7NgJt2ICckUbtJoOxnggyT3
lGoJ92+xAit4NGN01WZB9d78TIQVG5XSjHfj+lU1xraCQtNnCccqYU2elZkNjB0a
m87Tdaj2gSqJEjhVeC4DhNCebNRk4ooqQNXHho1XSc/5N5zO9zsiCDuBPY0OjR83
KzRIOf8Qq4XpYRr4jIvaifhKS5SZRdEuOfH/CWAi5/gsVlhZIeGV33ajr1z6491e
enY6hWuaaNw6+UHPIkXi0NG0P8+GAapY3Yqf1KDXZ+hD9IY5+1NIwjH/eLr1YJgf
0LePL0WF3f9NHQx8Ilo+I/LkgZs9TJgMTq/eRW9goRbuYvdc6Yh73jFl1PyymqYc
Rf9lYufqJAog1eJ7A09grs7Oj3NcQJT9oKF7UyeGcY41vJfJVqkR07Gl3LSbXEcd
PVXp1VEYON4FwldWZxVWZnp5ZlihFnArDKiAAlr/jOifRhFDU8QDxbhm5O6gSD3Q
WwOKNDL6bdqL6VJHtAf7Y7C4DRtMdVDmp+Kf7JuJFBQQpri0Im3ZAY0lAXv7GN28
ZYK7bJaKedf+VilazUsuiIKrYdOeg5OM/qs64v+++StRRihTEQp4q8Zw4VXvCPyN
25+XsnVMhW6lQvfYXQDwrj2ZjkxBaghixf3v7jYYclnF+FlbuRRRdd7+HoApbPO2
pLb8gTWBoNdrC0QWfkM06SWROdItxAkhImwp8+SHgf0iWr2bFbef64dU4RSOOg5X
S2IHdyGsReTPE6qtQGtGJVzXFE9HKgifyRRBujlQmeIQ/Qk/1LRW4Wpw6gXK5G78
75Wv/R0HJBd4bTg2DKQjnFq1kbj7ay9ZkIb5EfQGGmhKbIttR+36HMoTh0pxs/wT
WqQfYMYpEc7BVZ9aMM9U6UZy+Pl+BXzZGgBjKXnd1UONIyjfMPvUyOs/xf57/+Fq
HRerSGupoROxvDvHrm/rYc9gSP3AAxdDjjShsXjw08ekLMLxKxkW3lEOwRjzt5zI
EV2O7UL3kqVoIRk9YTiOHnNkVbC81GWUrgl29JEErJ7NBBYFFJ+DWRPD3YEYfeXG
lNB4dxPlJoeAwJ1sdG4+/SgiPVmrUYdDHWQIswKmwKXRKFX0IWS8KIpcRvN2svws
Y8Re2QV1Ssr/wJVLsoImeGXZWQb9g1RzEJLeApL7EsIC8Ahv+IcP9Nhc+nLeCyZ7
p4JaO58nOXkLCXJMziRPjTcYdLk1uXRdBVz6C/JuLOngo5aNWUuN5Q313BNh8Z0v
nRx+0uN0b2pCGG+GeYtv6zn1v2DSUoaVDlBhSKtFZ7eCxAVGcM971lnlI3uStPer
yy1jiHH38Ty/hFeyXvH3Vli7A1fHlED+sBurmmf03RYXlqMEjMhbPLe2qmN1pMux
o6r3NXKSiMMdlIZDsAtbg4lXgwGvoz9GvmFrH3KcwgtWITPL2rb2naknNww5HAW3
pWrso3/E2zAScU1m2nb4WrZYWv5aotY1tWbF1LVBw289yWFdo+6Z4LHMvktpQT49
ktU6viiD2M6lGmgmvGannlOmm0J9h/PUdAvBi8Sjc7m/CS6PhbxeoPAwXpnEatsk
mdBL0HEyCzFLH5oR4dtw+Mb8X0OBW+rTs1nkjbNm89jUvdwWK8leGhFyGvUYqP9L
QAWSCs8qv4r8RACZpDQPgpJGL131OA64wcwdvobhz0/Z2al0UhSedsy/HbEk2rXj
Tu4R6FxBnRdW8Thh7UFDJa/A9/cmrZp8yy50uctXTwCsjvq/RTzMXC9kZFUpkYYv
iLVmbv0Ig3rUk+M3W0zhCH/E93pZ6j0iHt1uI4OqAfwQMgb5THh+RTq9++NrhAYy
YtMkm9MXUt6U0T0pkIjBxbU4EV8EcThjK+wkGKftdAVvx5htgOdTGChHQePz2u60
2+4s687JToEgu1IuNDggbPqXAA303bxj2relGCRqkLs1CU5ONW/eddwJxkggLxeO
oEcZLOHUEk+/jxLMSWAIa0ZSO86qRU9Z7iB+Zo6tES8ZnGBwMOpkxbV374nn0MV5
3K+u6kDnZEvdPF/xwrXvN8JS2+DykeLc3FJkNDQjvH+8Xn7/yRhj+rDVEpuK03Hh
ydYxXTDYTtdChjx9eRUn5Iai6RBxxLJOFJqiw8MLw8UyjKtIIT8ePgcMKkMC5Vqi
Us+waQjs/aDv2DDZlOFjzp3j8FMMf+4JeVvWJKMgnAyaOLsOaKkQu92QxWH3YVLN
Y88vZto5xhzZJnJczHdibtnPBo44/xPkZIEWlLxYxZ6qwC/9Xw6BxfdHTIXvZX8b
2UVixeaYAQEI95etbKPKGMJLTjv1/0WaHk61cQD/JCFjHeAkqcCOWy5GUTu+bUWf
4qC5h1WIMk5UBB8mgz31P+66qBalGZfpBEsxR3yOXmcnt7d4vGnopjt25t+yP7nb
zDscZKMgCT/mSbMsgREsYBeX9WT6jcgHhwdOIFK++UKZWOmFXESNu6CdN24DGNaP
L4YMlDHi0uVIme/UWHIUirCT5ViKdW9rFmBvaZH9n9S6VppdkMNCI7Zx3FoDz9pS
2mujcYs47ELNSFsLgmKN+QJDsD6jKHOoGoeKtJjyhQuHpxYE9fBnUP0XWdTW9dyA
irlTdZ98K3q/tP5iodwrmhHU1n1RM6E10CYENQP3kByoTCGXRS6sLykEIbOfOTeR
A0bt0ldQvvSU7+noEVs8HZGSgXfWCSKwnZgNzx7bDiyJ+giIwtIhxR1svhkODIoc
5v2Nwmwq2P3zccAOYfS29mC8OBmzzZ6Xkw9RICRdlcdEU/rHKj9MiA84blMU7cjo
MW791jx5OjmaXt85FIEvgBoFelGyGNys9BVWUYtsJWvb6PTbf9GNxkrukssFuo0L
CXPDkO/6buVj5jbQV58YFOt8zT0tpFZDXkmqI9BOaz8IYr7ThSPNXG4Mq21MYwaG
gMXVicaEoIf8FgoPuSTRx8e5hB7DFegaorekEVBHzWusOUMlcwuypzRnER2ba6bo
QPH31lVcBgzzm/PRbxes9Jw0FNTFrQ+4aeGfjnau86JWNc7JjxBbT7/PAkiNQSFs
EntIC6GtyBdTAH6BenqCwYLTaxK6rPridqcIIaeSbnGMdCcbJaMvylmMD2+f1No3
CXolVyWEp42tKvrNvgz+sWEk7zOD/hT5wbSWKrsBRRIIKW7UFD29JiFpaXybLMo4
mrm1y4K8eCDb7bKBbKWay5pDNl/sWJ2+8Hsjy4tXf89XAL5Ru+1dYL1j7QP9jlkI
qfPqIIqi76c+fCjAAbWcTj1wqaHYrp0FiHM+FXfbuyasvq18xFjaFgNFjx3h3ilW
feKz8+VgMrOYuMLp2G5izX7NM6X6UQmfZ52R/GevYGYxnTxkUioNzfExFITakXnv
KcL4x9muQTv1uXRI2FarXPSPf6a9cYWjOwuCS1MegBf0vfR+9cDTZk46X4f2pwCB
Rga7E7CCzpLSXqh4gCXDbzR6J3gwJRYpED3HYmayflyL9T721Uupt72gJujfMkWX
IHQyeIMZGJ2jq2k7SDydVp6Efl1jw13GQgVakMogpB6ylAuWuwrSlFqrhJuJeyc7
25+lfsvSOIED/mBsAqf6eFqKhHkWr4G5rx0i2oeNNjzBZ83KsHgMTJE/0fvw1jKQ
0uRXPdR3PXoqx/g/mZglsaQ5Zvcl/afU+BXDkb0sUdnSSROQ4QdA0cQhN3bMHVft
WoIKyTxKrJwi7odR3eD69SUHzP/2ebml881vLCut/WKBK3Kfxc4ZttuFmDJNHEXO
oliP/Br3iK2fKlEiaYPNkqukreuJFjUkw/0xOva91UmBH/Cg9vyw8a8fsqvpRDaH
DQzNrt+4WYRom3gTFki9Il95PjE9z0vaZKHxXcbWUbrfOs9nPY04khmQK9G8Ngi6
puWim8E0x88vlDI/f9qswE2pr5VEr2HjUH7lCupN7Gof1/Cz11CEMKsAXlRjPsKk
SFc/9PzXttM+PGOiFp/2JCcOHwd9XbNM8AUTnsXhZIgXT5JRmLk7ovbDV+AHOVdp
wJU7vRKnnW41jaKvMboyn3uLJ1FgtdxvRZFpotlfL0ktriDKXq1ENcdh9pfWtoZP
ynEgo9H/Z0koiKuabcbpjn4nj0zEuiV3WmvLYxX3y9m3EjgPQLi3ITY09CSv27Nr
4v/nPY+dOE2Mg+cDU2eYeyicSUexEAA0V4RUJ6g9LqwnsBR1L4dPlZC+jAzW7c6a
DELC64Z7GMtEmSohOcwqJhUUj205xPvLPnMtdWJvaoetlaoe4q+pZJhur0GpdelV
RDNUSK5Pam3LB/FA1K3Os0jazrXUgnHwOIkQrjPfBcMTV5VLCZuZPt7nQ0M15DzU
I3Vwf58V5RW64fwsjHCHR/4fzZhBEvgRbolAdKMy8wPWzIg1fEvqlSDiG5SloMl4
hsfEm2Xan9eQ+QzBVlSc9rQ1DR5c1dvzdfQZkFskEfG4MHwVQSNVSfDtG1RpODyk
vBA/XsbkUeaymbTgr3jy6ug/T3QKe21z0ARDfsGxsOBnFHl7Nruo2HeEa5A346oQ
JTg5N7yju9JsLKJ8rlsRFp2k6nPNKBt/dVJhclPBdzTikm/Db5uFKkMzL3cp19oJ
NC8QsUnqQcIRVNl/x0bwbCukGRzhFKHpflITQz3oEllVOIIWUtK1ABrob11K5kZ4
sr+aGv5mu8BuluSPtcoHfDnM1qKuKRgdS8r/AnT1+BOFs0QL68deWiIJQkfA717V
6rc3imj+Y18WvbBErwmmj6vrKL5P3SeOVjfXg1p1vPxAcszPoWhGg77t36JxqOHl
hurumMOEAJVpiSE984TpyV6eOT6hP/ZPRDtZaV7HZm8ppqwlUYyQ8k2Qa+203yXX
cMbZyQdzHhG7jQQC3g5eFNP1tOQ0l87fCdVUBICwKPtXDkz0P8aUxp+FrWupI6lN
gkjIaY6nw9vY7IKvKbwRbxtXZQhm6werBf9+Jsk7VYtlNEJ/XS1umTJrBIYE7mrs
p9BbnH+QM8dEP5SHQ0e4s2qnHzbwwP26orRiURDnqhxYLoS/llxFc/d5cBHVrBEm
PmYVBqBrCm+PQyomi9CaMjqNzJh6QBvePQDEiB1/rFTbgpkjwuDsMkfuMcK/44WB
4m++qNKPNw2hmNauAhV3Y9XLZaTGn/qFem0aPpSBWfPQNDNPDfcp5rNn52BIitli
lfXhjB1Eszxj9+HdXPNktZb28OAidH0w3/bjUb08eLUhmQa4QupMNB3LqwifLUwl
xEGS9QrL4Dpund3Um0Tjz9+X2GzkItfK1jf/iM8mULVp3SGo05sl3vB2DrYKkmSH
vQpgxuAtqXhJwZK+Zrz203QUklj9RwdKcpvAxC12DvXTUMtuMu560nTGtGNdcyB2
OAOyb3efgkHAiD1jFPU9gi+YvbwTZJMOQoKE8ZxMKCVlyG3bCg4KYVoqJ+WkmGhj
dQDR4r+Cbd9imtePSowlcHYKBUc8ht0LaPN9CKgnFDAK8Wj+XTIRyaMgh9DFUBBA
7XIetKxbDXb7snuRqSiUWFK5FsQdKJK42nSg2qdjjtOWBM1lz1Yg55e1xpeYaySF
VQhPZF5nLHY5Y9ZythQD2sjLA9xRmLhb46X/xijTelJ0E7tDQw8aEVmtMt+94iJ3
YPEF0D7SHecc7Xb74Pty6E/cyjVl3Jw0/cLvYhS2/DIEP5wHMq5HxnogiCnJ0Te+
jg8pYyCy253PE39eV7+w02dklJ2HSMrgUXfSbLfmb1p63MV8qza/bdsfiKrlfY63
yjt075diQq7q0xwSgzV1iaOJBWhyXexWBrMYZNzz4TyD7qEghrC33LFsH6+xnboP
DuezVAYUo8RJhv/SJi5B20TltKT8OVt9TF/PDoxY0rvLHhkTmjN+FhRYoSgJIX8x
mFbBPsbjHNzC6itXj5+qaFCF7wtd6VbpxJbFgyWrzGV9lQjYm0b0DUAjW2htwwhP
+UvVIs/Pe0GN3KfrQnHAZZtAf81e/mm1ZgN+5/BX5elDyBQYqps6GliawmogC3I5
WsWfLHL7wQbF/91zIjNogvtFxIALOlgJviRhsZgWvVM0GUkYY6aCDZ2yQ2BBo6g+
rbCUtBNOv0xORjaRU1hThPT4FF3TMI0rEIQHYoOVYLil5JXKL53kenbR66MRlvuH
gqD/HhwUCfacu/sLbH1ZGhbClMjUjmpL4wC43Oa+nPtDrrGafFaYioVpAhEJ1+zq
upGIqKUsy9Dy7ICQ59ev4lM/2B1BtpNXA2xMwa9bbmKoJHLE+vtt827RrATwBzwC
4XAS57F+1n/BlaTdd4oU0e931GuuxGVjZUeGNbC8hDhDPixJ5ZHgCzn4jOyKDUOr
2m4cmuPicZ7/jCxETBxBeoGAwItySbaxlVn/d8qAUGXcZFAs/CDY6AxDvavJ4tq7
dCHdPmO3c57Iy/M3PnQ6ASTFxezfSXOWCdzc2mO41tGej+hGuA1tQpdhZ3B7i+LH
63CpxSeYMepqKWx4FS6ww/fFKpAbt0nEpe+yprXDH/zjHgPWtjGjRTUZtKXYiWvl
BmEJ3k+auOnrMhXEAOoom1/4TVUqAJdhm7D4Fo2GpXuNHTfHpTa1skGjfGowrHGI
MNw563EEKogTEwY9MCEB6b1q5W9p3K1WhVQiInPIaCaAj5T4ubRl+KTqcguM/gky
0m6l0EBwPLlSSBDgRU1MLaG/bDUCYBK9UA7Wx4S5vEdel6NuuIfYpFBsM1QywF18
mLKoc4Weq/QYNgpHBN/ig/Z1jPw4LmGhjw55S4p7lfNmoEtvbqY9bfsJ8kIVv9SF
vTE0eFCSnJBBAqlZrCPyIqs90Hb3A9eUfyA79zOUobsrU6TMpg0fwfWmRQbaVMIC
AJ9hDqAbmmiA1KMUKDZSmbmrMbIdAnYaxhSAhKhMc0T4udZe7C356DDb2rXXqlG7
18LxWFQJny4DnbiJQ7r5uKs+x2eEfcVGMD8SIXQWbIl2Uea3hH1DUDBBPF4rxKbR
EO2TWmgzOYD4ELGZBtG5cmG9r+rKTqMb0PRAPejydTsi6g7yHMjm9+kMKh9xg7B/
9WG3L5vH3blIhDrhjU9W69QVckmpMT+t5cMZGiSnscqOJvxA1GAbi3Hz9yH/onYU
dIO6TSS7zAiPpsiHYXz4rKdWp1lvtLziCLx3qb1buc+YsbIZZDgDHH6vpG/1KYEs
KyQztFB1bc4KyQ4m/5EIDlxodW/BIhvlQc+rhwUX88Fw1D9n1CzIs4bMrW7XJwwb
peYbNcn2umfPeZxlTSa8QVcTDuPC80dhhO17nmZLDcP6VJ4Ouq7e/R1RXt9ZBmDh
rky8CluBYOY6b0xpA/KCI5dmBGNa1yE2VOMpzAeEYlyL2LzPAkkSO0qoOKw7IXes
0Rqrl/q5Xbw3kuyBFcDl2jBHy/SoVYzWPOh+RPZUZUdaGiscGYLteKrDeHpK2aJo
eCBiylO74WEvdzyoOqvnfvHRgIN9LNkSF4Y0QKgDhJeBjUpZmpTvxw8XGy1awGzh
W14Px4A2Ox85kPSPKC6tF1hWCJavtR0h684C6gC/Wy+HlIdOiJCAuLJQV8AUkyDf
bnvIt0BJnAW984fvM2bqwfoYOpPFgW33prAP3KBdhwvFTmxEpFlZUe+8h3ZpPhMZ
uXXKpYpVVr9gxzzhygn+4OQJoqsnqbdIr5cEVyZdsQ2efS900cTBp11K9K3I4mAt
7QbEc2AD+iWD4aRgVDTUaCFd2Kk92VG4K3etJgeNSylOLZvuFzGZTgGjKlY5f8N5
NhTKvBmQ2TaMFgJ+EsFf1SIq299vjWUHLIJ/zjWysRJmTEKcW/xorFww2TJcwvUI
3uNqSvauQlxzsKWrtRrQ7zJPdeOwV4sfawOhnRLXBN98Ld/GJjQeeRy0FubK01Vg
YSBdsJGlgo2E+FGhxogcyrqVhcwI2paH6X5/l5x9FQ3u9XrMhP3ZS9mP1xZcArLW
9kgZGh7AOB1Bf9Bu19mv01g+DFr0wT1m53drwS4pRs/ABG730AEQk7EuOZQolKQF
ZItNreTtHXbdTB4wsgc1gqgIXVVgACAGiVc9SA/QkHO0mCF2x46ZNGIWTJ7eHyrI
w8GAJD9wzX5KKJGA/xPnOj/kJmSdkpraOKXJ4VmW002+W8UE6BWIrcAJ3q+oXdVo
472gmF2d8W4A9+k1KjyXAUCcRI11y35KbXgmlcUeNTczL7SamESvcBKaAEls8Zqk
h9/hqmVyfNgJ0rKgCTNR6w92bayJS6v86ELCYPNgEbJEbjtnWbXPuFzh8ztfMddi
7ChLyhLwLXqcfQ5vJfyT6iOCH6wVaFZqhLwjX412Ato39rkR27p08XVQwrnzk/XS
Yhi17DfvTqqNoBfBwKBx7DombZG448n9JxmPFv2bplNQqCiniBRuElFR47L7+f5I
HgF2bSd3LYBuxX0Yah63YXIhXA6tukAgcBHS3adwIFjwcKH+QHI2j3uX3Ku0T/eu
nS0jUQcVWZunch4k59Fz6J+hIdv+XSy4VFEJUF6oWK/AP+ApFSarXhUVgERsDHew
6n4jjhdg18vw1WPZAuP+m4LmItVgZO1h+oemmlhFr4FfOQ18mX5hVmA3Axkyb4I8
esO5CNKCUGdZcby8bzbetzxP8Rz2hWWugvofKe2dx46Jq5GxSlD9wkCw5LfpAfwL
jejuB0pQz8h9Zycdw+xIcIK9Uus3HPCoSUc5Hc5+7NJX4D3yJxe8ie0Xd6TEo/6l
rcetF3hu39kwz6UzIOm0TfkL1BJGIUgfW1e6qcUUxnLMm/CgQ/Y1/VQm+e9W5Hya
C3vqRzK9gmXph9EjFGbw3chFpWCfa4kzhzimsmoeCzM/9cZe7EP1ietf0WOugR3B
l8to9UYcGgF9cZa6fRLqcV64VUCJsEg1591sJcR5rJP/zKeqsNL86kLDzkJ1PA4Z
/1LI5shtwSBdvbjpdakbUtig1vktV8tcudJy4QVlmzJdrAAgv0zsRrJ/WPRDW+Xm
Kz9t83otETeFlOS7af1Yn5JCobzJbn7lan9pEQeoKOfvXo6ieiTyw6TwoXbEQYwt
wXj6CbKIO2pQfTWanuxFpRQlZj0BB65lu3LXbTZfowyBpw1slsp/KV7xu6c5g++g
bOXCSOQAbk8AFtS7k6aqzN9cndkui2vlff+Bjht8hluYE4ADlPvdD/yTeqJ0Y2rL
7P7r0yHgBv6pq2MPzgkJHkshY3lQwSWWP0u8dve7Y+buznKV1MPYdcAZ10KIj1Ia
GHhctW264OaKABB1zYyuPNghWYcs4+RcJeILZP2+ZmJyIE+WuLIXEFdGuAbIzCWD
dezSfxjDSHPxLKc/ca97mju2CI2Y2K1FQKryRYh32TfLVlWVu2GRqNQrfhWzYdzU
S77ENtn5CF9PF3txuApCUdt9TfyOMp2qOmR7cm3UDct4Dne/wfVp2DNDjWE8zvHK
6Ng81dWqaa+RnDoSE5FiQYulFJJyqH41J08ft5jQLkfUBahYJloG8g426Q0jriOI
XhP40/sSN0f5VmU20dGYaKutIUrv08XpAQ+CqRpfwAlY648J6IzbyB6XjrQ7QUoC
t3h8lAqD6jkIfiKmQ8nh+65M8Bv3E9z8rhqSx8mHHqfIIrXA9+RbsnW05CzSFwUg
Eli04C6QZFcCfEUT7gaYwFmtrQFtbbLO//CADPAYWIai4PntxlJDBlUTAl9IwjrU
O3xGRGc5csm0vJgV4w+oEX6JUoPxnF++Zg3PU68wHWE5d8CgALuqj/aF8y69RkES
Z+15Uv7XbEdfSINekLrnbCZ4gTA1hd0JXCUtDV73bRd4YLDvXgvoZDY5HRbmFsEm
lcLeKnloWWKEEQQr5LGtWgbpJmcC6YN6D+GbuirNDFL8vnAcu/QkSZD/ndk+0gfW
lgfgYblm3aBREHwghulpD+nYh8wZBxhx2CDz8V0New/X0KtLCopB/VZCXO5G4Oux
bpRqqfoWtZXZwLGC5dCSZMphrfTrkzOK/k9VP4nhoOqWppY/9z0AbQYjlqVnySJC
7v6/JTiqnNumvw4/OHX432rcI9jce1kxPklaEw4jJrymErW8m7h3cMbTSNvwfLfl
8uCYeucpAWSCKt9xWVpb5xnuDzOHuDiXiPTaKczkqlT5mbl2bMuszJGBw1kzt8gn
tzHAcBSrzzsFXAN4NtMh1KTuBRjIBDNUrenvgOx7VtNeNGnVpXMg9VXaCa7yitjY
dLidpnOoTelcKBsf6q7rUnNAFBWqQvd7VzFxT/mMqsqfqsR5Rnk8KbM07Ofgv/t5
zdni9KiZu51QRbZH7Gc7GbaQ+Yygn9ah8io6Q6KZCVb8VYFvaY54RTMe/+9+S0A8
D2rPELOiz1ltqQXrbmYwiPm+NwAPFkEK855jCjoVXU37iIVpze/fpGASYizXr3uQ
23/Uerv6CbFZXX/JKjKM9WebSfOcWOm6SOYrhrwcZbBVPMUWX3W73bqnh6Ua6Jhs
80lDDqFSKYKjQ0PFIT8Z2Y3zKXSYgvMdi5bToNPznhfbGzC+UCR3VdsDT6T+UDZt
zj0Q6uyoECnv6o8y+qE//PUVOPqrEFjcpg8aGT/TjcqqSQVRoPyy0teps3U7m+yN
yiIRXyPxvQ//Yl4nrRRiNjLVVDLuX0ls6kPqRZjzfUAsBJ9vhn5uOdfsP0qGKgkd
lOAX0q/fijEf9GRNGRxrN0I1YlK2a5gjxlV3Jg8D/UfjT9MjacY20EL5r1zL/eHS
Lr6zBAMW/PPF8xFZouAWC1CBQgJsS+ntlUx3YfrLOHwkomx7gOc5voBWplsjtPxh
R6a7ES/6jUVm4CBkCptgdu0pnZKOPSynJwlB/ruhQ1Wybqj0RI2d1T9c6PMZ7jAB
wiSDUReWm4YNgbaIxWhnXOcSD00cGn/AZl3c2JcL2I7s2pYnsPaFA2l2OSfc+udI
HNfTIGKN+s+P+3lNi0FLVKx5foX+EwIholUWF/YddA2F3TZnMXXAGuC/bMzleUsv
p0JJD8Ca1AuYKuiTSeFHmStxnJEtivUoy56+xiGIwt7Q7hhIjEPNiPOQjY26wzc4
0lsb24kHUfFewrjb6yemam8JKmPVerUO+QJuPIIJ1DUM+UBuo/olCMkiQYUX2DbE
+mxo9YiW6ylaiTvNI9Q8V4DAgH1m4T929W3BiJ4fu7a2HUZwHum0M0lm2haAb+Cb
GRENv5O8DuDssm6a39ohkdLt/MdORrG4P56++4PZpobAs8PI5NWchFaNhiDT2N0Y
ybosY3OHlRWqHeuTprf2VUTpaq46tbFvI6YPmf6hK9QGV6FzvqxXmc3TH2x7DJ46
2o7NUB//mZ669QDMYK5lJdjAl/xYzDeXK6YF/Pi9VT4IPz75szEN2xtb0kGcB9Ic
TneM9ZRrNFRL3QOpMXd3+SgVrbmpWHmXJNGGWdTBgoQTmLR6E2/usqv6ncamfNlz
eQbd3OmNu99nQ1eOgB6p39C1KrqkyyRkatA4mfK4JkYI+lmPIZzo/YnGDxahuAKt
yce4PiESDflOb02ZxEH5LSNRPV3CqNFQ/s1hXc07wP7+pi2sOQtlMmyVrRpEE1nu
SUGJRM8yHBrm3CA6VRXq+w78xcp4+aHvIidfQfPlGRsSPrbv7Dq9sAoR1IYZ/MVK
aysiWbTXg2Oz60Abwr55bqZp2mQ8nqRCe4kU1qtdn1NnrH6mqAxhQzAiRhMYRbuL
2fdq8ZMNsIz/f9peROcX1ciug4u7uQCdXu3F3HGa68os+q8n2A2rSsmNVxZB8DHS
0OwCr2sigj5Vozwzq7yNLiMf/pqYYzb/3X478E15JUF9u03PDsLntG0RjY2ACcf3
V1fCXF7faUGy+qbdBbqTTh1QluAdEd8c6K4uvJ/qUtBR1hOp5a2cz4PV9RGe0BsH
YSmnBOmxe8ga2bHnUNC8NFKKODfa0lynknTzVF6/o7Ys9jYl9+EPr4hARsTuB0uk
KMJJxSM6Yj6pgN+1pHhVsoqWd/fH9+f1MDTZpM0MQiKnY5vFrfRNJirHuXv7ksOJ
RucD59OZGBn1vvWK1T/IuSQI201ZEptsEtzsYhMsHi7rRzu/TQzSK6vyurI7joxh
vv3PJdjee2dZ2UvbJl4nHwfgMslgLwveWgfaIMgSNB5gABcoj3108Xpg23AU/ipb
NjkCbJbX/vKIE+OSyQjqCF+rJAkMKg+5elcLMJe/bp+IwDiUI54zJ+BaChMsTp77
EG5w8fC4rH5xzf5WxFPfNA4euGKw9f86X/LFEwobGTAZqgCvM6mcUZYgTuUfmcU8
Gkm9a9w28v222ZYJDeWGdJ/guz6DyBr14wa2Ug+TXHWjI8twuFd3Egh7raJk+dml
I2S9W7oFICe2feXZqgE3NQKs26IGFrbeDpbuTqmiin7SVoGTIfXjaNSM0yh6UXUx
58PBoarDlK5sdWIf3QqQn3uUDutxA4XWGDRkF/8wzebJ7jLdoI1QC+BHZYD06kxm
KdhwAOieT0K3W6grxndJ6Zerltr04h38Dp3NVlDkULCh68gdQCHtCMShuFk+VpZ7
LYnW0r2vZMrN6nbHj85JAadqbZhefmgXelutSO7x2hFhZwh3qtjUchvjyLPgwi1P
/cF1hcaAn2qeEs7+YN6wEjHBnZBBKylfEFR8C6WmPPmJFemViLcJ1W67/S5bBMwL
UGGN8H+5jRo63uViaXKjIrwI4C2dLf1+wGjlnBKiGNwFeOZV1kV6o+sjIjNPGgsr
g4Ud4BLyN8eqJ+dlCD8F6UOpTIwDRYfdQR7DZW1wx4OJJ2YKFElcKOqr/FkydoWF
TDGn2TzkmvvlV6yjOIxJk0KMV5Ckbc36pEPFlxNxJfsCKc58E9RDJDy5cB0UfByg
34j1lx7JzGnsFk+95VUIcYFHCMjHbLZdtYUzbm8++i4P7fAJ5/hefPxyJRhq3vWA
msdHiy8VZ9H650vnatI/VzhVo4xnzTBBVjoQgtnQ1WW1evnxImyJh3MFapqAB1vo
ed5jXGBh9NXPM25LUEc1p4UIOfn1g0ZGRgZ3fpNlm5d7YOmI5kHsRwQ1THEt442b
xIGkd8Y2lC3OHPdT7+Py+mxhjj7AbPCyDm6CqIOTNUY2C2aUg4iJA9ydWMk8QnuY
m+ohsLurwgs7DPJScYD6/b0Ao362S6qf8rfqvNHL9c6zkMfMFht4vKvSoeh95ryQ
Sux66kdyXe5NuQU1R6vihid4tP/IXOZ184HUoXCfPa2IYlXUX+QRvrR1zMNni77s
v2IPym3IJisuGzXzAAs5LIR0c4KY2pBFasKnXm8MTTM+lP4pLSYZEkqYuJmN6LDS
5OdM7gQ4Hg+3GHS4MtD9SmA38GRYKSPMMYC3lWi3ST2YnAltZuaRGizPulC/qXVW
SOFUiOZ5suYizqotg+Eh00wipwNNkHdVHiffkCjSIFTutBlC+SEKUMMBmYOo0s4g
gKcuVpWkp3an4HafieqHZxjoZEU0Ju5iClEIHLWBpPsG8NnoZlCoTNluQ8qH4T4S
768wrsAtY4sNuMuMC+cUZ6EopX3cypYBxplwknIZLsZtuKLGbWjFqBhV2VAc6RYl
WE43iPLlGhVYsjn0fVdli491VWAtLKVdpoxTQ86X6rx/z9uVKCDaOY8MsYD6RJBC
0SyoS/jo0EoScFNIkQWQUiNtAYudG93CbQAtRekrTl/jPjudisM8Ub/5NrZ97mIC
qNKqTrdIjlurvLRyo4jBizaNPh7MKq65fC9iP5F23zK+C77h3dS1tOpZ69KARY5D
cpJp2PsEaRuHXTUMmnN1BFS/3p+N+ZAd+fMK1/GFG6SJQIZLK35bE3bcKP6XfS7v
pnCYJLIrVTziEb4c/sQnrGEHcbtaOPsyFzmsufBFAw8pbugolF4V0AxopPcg8JIl
QaPrlg4fKr+JKIeATFmXH9IH0FAfWCUTlly8BnmEqk7JBQicIygx4JhVyCxZui4a
jPeeVwMlKe5Hx16Yb7CgER4GlkuOvtJQCQ7daF9YN5tgvU+OQvt4VBmBfl3dQcne
IbrI9wzmK9NWToiKkKQwfvx0peONfpmtDVbP6G1ssM+oqT7V8Nw/Dqs0SH8znaRm
A2OmMgwZUmsPZ9zVDclwvSMK34KfB26v5iX8IprUyTJ7aYZBdBx6FlCHiaCR6c08
2/co573FKhFfF2HkV9ua5A2LcD1fUg43t0Png6nAMNaU57egpTF63ShLxg3JFm0/
uCmv87Ad4bvmKT6sU1pypU+Mx1gVjxJjHArqlfZy7xUohFcCBCa1pSQC5s7gvBLJ
ebR/kURVGeF85DnVN0w4Y70BZt2iB/ovmHetReFqDCQA8++wRUbF3ThSmSYEL1ma
dg8IXFjqw9OWJej+fdPKhPZLSpWgqRAI/NbO3Xd80LQjIN4jwjjgPFcIL1XLoUw2
sNCK5klmKaWr+9ETj8ETZPNjuaWpjlNwQE5HbBBXwNpWPuivtU7ecEdi1v2bPf7o
2Uu+9/mN48FRKJsmCPcsixQiBwSKQbqK8T+31asCywBnbCWuHeLtKw61W5+NEJxi
BizpYsEuQTIP0LCUvKRSypLJHdDkApiBXMmmtoAmSEFRfz6+vO3z5Bpo8gALO7sF
Gm/nSkk5XC/84v+xDE5HIRaXrIRXQO2Qm5SQryn3UQmtincRN8ga5A33Mgu+gBEw
g4dRaVM3lFwSuOWhorr7L8OsrZmq6EgJaVqfHYNsW7pE4gnNoede7gC6LMbii5WT
1OvgomWcOsBgxw92AQlbWdWCsAy60rByZGIcY09n0ZRpAdOcuAKPbvsXpH8JfnaK
JsWDjBtJGN6ndEaVSmugkJeQGOlvKmwcAbsh+g2ZcWxpJnRBbqd0io8J9cnsWXug
iHoO0wO6ufjY0B9VasAMJ8QE1VwJEYeBPWqAuozMWsn8HZjNJb5BgCKrG6N3HNzX
WBtn/bCp8pTemZrTNe4Oa8KlqzmN/AxKFeK662jheSBHd/CnQedOEz85zlaMat1k
Xd+rnSVTgeIQmVyHNkYgByZkTxNSbTmElw24ek/jH7j0CBSrIV5UgZukYDUUT26X
vpi/9ia7ky2Xi7Bk5th2v0iJTT7Fp42Nq5ukKSLE6hBrWI8/Pv2Taq17PQWjWw1Y
ssHPBevyZLXg8/azqc/nX0PWh7xJmBar+wbnjFNbOcLHvErEUHm6LR57wQLjYLAg
ravfHVKSbWgvKQu/Jru/+02WiRsHQa1eCtAOLjiSv+kUSzXt4h91oBBmYNGCCxWJ
0lvwd2rsz/LDENjOfqQj7kEZZh2pCUIIAGATWcwMNr2Gsa5OXOdPP2yRLVHa4dEa
pbOBbf9/O/2BrBaeD0NULk8+tx51BBjt4KpLkf/Rz1pgX9m7HM+0cXTH06OcMicL
5VE4nLM3Qh9dFPQD819P7/GX8fgldDjO1piPKDYZaF2n8SRc9ZKwSRGuBTMyHrR6
lZR/2Zw9s8sOni4aS4O1NpQg7zxAGuXngPq5usVHz6DrLwGx6vz9h4VXpMQraPXj
Wr8b6hqLyyH/OJjKYZZOFwi+pHie52lHIaCcVWoUuu8AbO6rGv//YxAbDVAuyg4B
zkd29uWHdUeizunJCXZP1O8BZpYVMVo5WV8DcMXUyXtimuu/kbKxNPscOZVH+7hX
ZpQbU7AAkpzn8ci1wIVYnkLG/1QzSZXqT95DS5AQT5d5F2ChKcDBkJK+QaxmPfBy
gb5PUITzXs1J6D6ktzMsNUZYboCV2JfkrA48gEqlrt/JMTMqUGHPya0ginumhK8o
jetaRgNqRRz2YP/G+9pFp3KLtOomPN1rMnDmu99FO2pNb1aeEu7fo7RyYB9t8Ohb
/eBUWSpFr/Y98zLv11BC8fGBlJUfhjQ2Uh0SiB2kQqEzTR0WohpZdJPxexTOgIAs
PqOWbNyWIMsABmqOABM28yW8dPjE4pB8RBC36BS3UphNhsHEROV1ydUjt34EYwGY
Tzo+pDGbiiFEg6Pd7tr4ltjht26ehd8ihF/IludS6TtaD+o/rpXPqY/EeVHGYUIE
4c0RZlSYp6wgG9msJklnp7nImhxQmiMPp7LTlQluBo+UlHvuCk3SUFrj+RDmnlj8
QwJMAP9Ndfc55k5zbPN1O8F3iYZdJ9+4FCGBqPKCun7p1eZWxB6c2/GAJTIH5Qb9
xMeVNQQpXLhKVnpe1ZM9vLOyQh3aAxRBLh4JAQ6UxJYLQ+fGAbY85mqEqprus5we
0JnVnZCErDAibR/Eqktd+i9ROoXKw4AIAtQbrlBLVMpzPqN+EqDZuSY7qRI2I2tV
/RrUNo6tbvMa6rZlqMaqTwtWj3N+Fk+69CqqsggZzZNYlPpfy2MqYejy8ZidZRkv
/dJK/0uym8bUd4OrJ3wPXoHq22UZP9Aw6k8mJxUr6JiTlOFCJn2wTiAaDQcLOHp6
dkeywd6EcJCcsqd163GpYoAnSc7VJvxdOpsorKJme/hpAd2GoPDxrTTfZL1ga8n1
NUkwXeIlAno3NjsAEP0+t0MYrK/12nu+A93zDAQQpglRUqZ+kOWT8vmAsngr+7OJ
X1uE1dgegffzkGg9K2OxKKBsKhD6o6ExDSjDWkQ/C8vs/3Y3NcitUjXZYxBg781o
He/6hHcvRWXZDeHVo+PLt0iQ1RUA7k0GHCt6qWu2rcFPGJ62mNlVXtTGLw1UDUrl
iF+lyhivOHXPIThf0lKXitGZrjodjSoRRvZxlC0iUuKgaw+pWv+ITGF7e8OLtxaB
0C9YlCIcftEMuMkOaVYamatJrycLVQGfQe+oAgPJw1dNHGm2IJMc8yhFrI3xqNLW
BggTRvyPS53zangvZxABF1n5+egCu6x9e93YZLenbufjek9QmnEN1y2RjS9w7XCF
sOnbwR0OXxWEqPawK/MgejRsV1fF53pn6p0lpUIEYImk4xscP+YVgwVAQ1laZwm2
GkPLbUcgrWUvWmBzgaTUOjjNEblkDH+2cTtfclsliiH7rZ7CvRizk4vSrtWhgPJf
6z8eR1InePBuO6hvkCIJDTFqEN+bdRKbFIBKgiDMWwpyPnj+NIz9iZucCL+FFek4
GJ66qSwV7MMi6F2N7ef+A1+wTvvCcZ1eRmyCjWxmC8sHCdZhKMvbuuZAzg8Jw2W+
ze2urIdoyIpinun0qVGtf2SqHsLK2zdYKHu4zA/Bm0A/DD/Ii7ZGv0QrVzDJy49n
/2yWBwPLhUtOAb+KHmlkUSHNDPIUEapey+d7W/Xoo8R0kDjm42QpuCjP2h3/BR++
Fw0yqL5Y8Wp29FCzGxMjYZSVUrkZdYRd+g2dX+hM6UBHyx+m/3BOH0LHdhqb1bkB
QysRJuh7IdOvQ6TYX1lK5AJoDY7eqooRxFtfGs63f1Vedi9IbvMqK6EMuUyABwZs
97MEp6bMl89x67KAWXyLe36RYqtzXHA9Dljev0SV4NV6s+udZSdSXd89XyqJb3nu
/aayYf/FbO+pl7KYMXwBg9BEEE5HFnryPj5lLcOHT3VmoRL1xv4+rLFccbUM/+yk
GDoH5fn+EbzEkTBnjGKBa57F6AaH0+Fe5ty2FqQpMG1ukzqGhiiADnhnaRDVYlbS
YdxQGhsBOAj2oG4u0fTVdPHKv0Q6GXuHVVdJbf43FmRomd3mzNUUnYwJlrpsPW//
kg6/q18s3OCe++iJ0budY71nZGPy2rZ7crrDtUbbRfeJjCv4JiPzrevhYBHFlmHQ
wpnusfY/S3fjdQ+UVD3F7NiWcr77Gg3bXZBpR2AgNxtZf5zeHEzWlBWSgRKb1gC0
8j7GATqKuBNo/JL3uZCdVTRp/Gw6MpXoQ4SxcNgBYkEj9An5vLfQ3xLaE+SRpQTU
DPhwkdykRh2AQlgZ9wlnmMulKoBE6BsmJ8CZXsH0H+SmjkeclJ5sU9TLT83/BlKr
5jDQJAJ8TfwyG+64DcBLceuVu2PWpqdtb8IkAKDeF6Yd45DDOIB5XtJEi1CQt3ZV
AYr9+PGhrsNN6Ko2qwwvB7iQlJSOn/Jeo4zSChqyomLthFBVJPpcFhljM/oaQjRQ
txM2P7MEOST48BTaXQIyfHf1partrSF5s1C1JdhKteFAfOVKY327sV6Kbl6EnPY4
inhzTIEoEboSz/h9p4TMSe8MEaolkZYCWW98KSKInWIHZPswaJDoTQrylkG3JLO+
tXKn5JAbVB8YgTlORy3X4YdymwYVqcKKOvxEMVQnYkplFN2HQksfHtQh/kO/FToC
4L9j3pHlXqw7WO+XltXF0/VAVSZQBjP/Gv4X2Bx2rhn9lcTVLCx3xFFd4JmWM2YW
InPbr81ZTyU15wyCqu51/WJpSFJn3s9554XedrO2VLUsQPsPVh/Kc7oRGqbJsKxy
Cw/2cFTUxGMd+Oo1lYuJhEB75vMIyjc7HNh+pP3WyPQwS75Ht/X6eN9pifwvBIaJ
u7Ol7mIiDbuB5yiuUvac14AQ278k/bSCkMCwD4nVOy37WPk04QUcwiU6COmBcJoD
dFCIFImsN4rLsjRs8gS9an7XqDXHmOvNh/ITYXn9g5Wafa8vIsuluFbh0pDOyLCm
kPKcEujKZtu4y5v29QdsWXx7h35f9MARzurTH8ZD79SBPjuo+cwdLzJ+XMeLyr7m
KYa6c0b24hkmvTjNcXJI58jzkEWEOm+g0s6QstVNcPkccC1i3mtbdK84JBwWiLy2
vflfpsgRhXiL4l9Tisn0BuBwFpNDIqWo+8T+dBSsydB6m+NxsMenDqkzsKm8HA1s
6ghq3wvoCNTiGMCEqlaWfQ1i00TnuFHLitv6su4UPopA9neofIgAJqUybhx0HqSE
+3ivzrYpLKsxNdXFQXTo2C/jc2N57VtrA6hZkZR13qwHvq/X+fNOgZjSguHBeAhg
DiSN5auqavz2PyxZaaUC6xjctexLVK6NtzZkG7c/yDJWfZ/qZTCtChZ37CIHWFjP
wXg9N3I3HwQ8mAwVeDNTde9RdQt2/H/3lAzceOA5runLvSj/dfaSrfY+Divi9Ydh
uwzBihLcJGPS8T9DLXvRLAyI3LYe1D+P/W8b9ADMOzleD+Q9r9Sh3UDcyho/Xkd1
CJ/JuFU8kgmJirj5V6NWhJwgWETkBQ9Bubji2rBIB/MtBtCLpd6WRqfujl/HI2UY
KW3Va8frUw1jq3THTFkjjYwEtuOh9INydcQOwZ77IyIrPy+GhZ7rAQVNT4141Bph
EO2mWGExZ/B75WxX+9smPR/sZ2+orgNwsAwN1zlFcbhisBFwl45vBr3w9fACMeNL
9Tj59wSD8Rjzx2pToSM03rQi08qt64FX1ggyF5Riargv4dB6Y+cgmX4st1C82vto
uLiGrYRXXLdfwoj/gD1H6+YMP8650j2DTpinNnLRXX3aA4Lty3c+bBCSY1PN7BC1
rzuL1Zi86Vaf1WyYUYhg9d21WL0kvOLGGX14rHpxsrrWRrmCXuBpqsy1Y9pkQpfe
Czo7CYqsvBBtjoxl5v0OxRXOTeX4TwwJkeZLxzvPJZKcdwRkD4qDdJKWE3cg/pmd
+x10AHebVALznXK7+6XEDkauKA2xi1zhvl/OIXkfobigufx/j40be7nsG/1H6BHr
nLk/83qMw0r3BUyrqkTnK7idd3tjc4PRAmz+9n6i5Bq8Xfea0TzTi5h1dfVpKvTC
aasaOKtw2owikBRNtbW7S7/xzm6RCIf1mBmql7DEFOnHUyZfAwf8em/E6jT7jN/x
ps+zXg4oAXQVNIUGYzHqJ5g82W4xqkLN43fagdLckeSqj/4hbJ3gqFkqoKgrRzcT
cMYiR6wteQQX0N+nJ9/5Dfhy5UWKFWM/K3tx564T6xHswmS2YRpOKWerVtee3856
+tDCjQ4HUQlcroENpMn3xTbfDVVF8JBWjbJZKVlTqO3GUc0YdBl/gtFsMM1tVdzF
SFbdaLfsbURGx+cHNZ0pCs3xMZ4cgqdnELqmIjsZ3Cov72+GikElM6rkboEkJfHt
qXfV89ep7VlirzAg+Z7l5qyjrwvRpetWGDXL02wXlt4PvgNhrqGpiFOxT/gqLuIr
lOeOSDIeTTnC47FDQ949ZkqM4qLmovq0ajVVGwC8wYdaPd5s82kbA+mbMCBwjX5q
ZfbkoDe1+TGUyXSnhfYfvW0syQouuxjbF6CT1mj/CS4PfEHlPGG70eUth+KgKS4q
tEp4qy9FHA1WYIPxhMTDy6Gy3mSC5g6ixnXGTHad2zOtGxeSU+bU04RqW+Y4mEUZ
87ThqvcHZ8t5qiaupriMf/VTiq0nwwLniq41dYUQSWqpOmLBb0LAwswAP4J/5GMs
Eup1zCW912UUwF5MYoMo30wLJG7alGLPsUHLx8weAq1cA52+fXN74jExEeXPnTrE
ZdqIMv12GATxRppF35JKtqTw4fDnVTqB0Qbc0MoKCEInkPPzP+U5KQ5lvgOL2ctl
MW3Wm5LXGp9ViWCRj8+IBPWBPN3WaDlGI8en5jfqZK0iQuKUzY/DkGbDpcySJetZ
+fiu+knUkkbf62VhTvL3BHoPc+4VlU52VK64np65+n7Z01U0Ev3/tc5IizD4moMi
0SOZ9wre8o/rU1Q7p3NPnooM4+kpfpk3EUo9yWE0xw+Ej77Juhd/ldLO/veFOk75
KkixfChdB95cGQ9xRUDtkW8T3lLCAuvXdEdPtYjbt+IBdGnHfwjLrVOPaGkNbUbF
NdZ77Zyvzk+YzLBEN0j0uB8LA5mWQ6MfdqFoNdMQwXM1yFYZi7z5gZ/JyJSDZZQE
BK3vofbANgSNOS0pBCMcc898WdZ5JlPmES0F6OBOyydjtRsTLU9FFNFCT6WTU3KW
wpcihP90FumSiFbWz+d/alrHKcwK650oHIuCPL3eidh9EwNaZ6fvdq6BHlrGn9px
qVmWj+iekk0tmfoY+5uMvo3Q68geeW0dn+g7r7fyKJBStidX6XTTn0sw8mcGwhZf
kDvVKRWZAx5RwiTXHNZiZxoYvSOjd7tT+pL3kKL6nw/mILvpYuYRgwV1zCS5Wwbu
IJYQ97OuGUFhnCcV0uW278Hf8E9ZU31pLeI/idIMEPykY+QOJgf7wpDnCYQrNDfl
NkDl5JphXrjXoQIL4Q/WNH8kStlCAANTiIVN5w6eOS9obqMI3LHkE7eoGQeUij4h
8Z5CSsoTf2YLBzFS/HX6O4W6A5gY6goBvqJ88yFMdmYb1aE4bk75kupJEX1zNsFt
HvoyqRsxptnoyqrNNINuNhIqKd6o05iJKxzgzHw9Gh8RIDf+LN4EHLJBBBhb0yJ3
D3g2/QPhlmFxyyvxF3RY3BtsGljOZqR6LkooXFbilBWlFAmNcG6NGKfTvnwfLpRX
OVrih49NEbN+j8rgMb3epzEGzI/j7FshEGLGLUoyhCgONiF5jIkC4DhdQUb5eDZq
P29luiwaoiNGyvc7Uuy3nGNBrjvCoAYnDCxei0drCx99wUk/08BSwANfGromPb2u
UhAdO+/SY7GfMhQVnPBwlBeMiUmK1ILn0UmZCOus6qCQSBckQzWOYzqKycJ6CIg+
BrTjMo3kZK9ydlqTi4WRw5M81KEq2NyuNVexiyLkuakBqvsV4AAs/8wfdMhRucUv
ptz6Sok+hPIRk0M6LJ+Trw5Pqe/vRHTGdpHfP6T23D+LRay4bh8k3+VZ0BW395Ia
83B9z5xMlCFfxhyE5gPgmiVnIdjbXFIi5aYcv2yhwoe5e4as50XCcJ+7+qkjK9gH
spIIGop8KVn3P+BJtb7IH+9Wb3c3OT1I06ZeG7b2Ma0f795sTdNFxy36lXG1iLrL
vis5xpp773GtC93GWCaHcKqwlO5y4e++xtu8qp63SPIFRoLF1J4PmrVZRuPNFwDC
PnuYOayjsMcwZ6gVd9e8WoXWuBgpD5W+HVncdULaR4Y8lK059zHj7v83CQFThmLQ
Py6NKCUQ4ssCANlT8Y979Az8dYj+dRnMIQOa9QKLwTjWbzZ2gM+TZv1ezi/gCzX4
OiatnHt0vp6MTP180MXDdcRpVQEpE6eQMrNE8hSKLcnFNFiItVNqb2iSD4ytaVLg
fk1u3YZkt28ZShNAi2bCGUeIgRd/S5FIzEqCzTkN4gT/ZsWpBGAuuxLA536/o6Fi
TWVq+cIpXyDbmfUvqijn+24voO0NiV6FwY/kt44BnXtpNeqmOtEWte9VQ+4iUxc6
3rY4sZCnFZu25R/VBntVANf+AzpIGBtcBZir5lJeansaVYgisE2fSGQ+tynN9GQZ
3ZLgG0xDcBg9KEB1TI0UstQbs236dBh3JXNhaPJBiCeqa1fZtQS2BKgj0G1OPpFQ
389in/6iJqT6WKwrfUYtLgzMpNbUHo4rPV5Sm8cZl/E+cxZymAPPhrIfA5Vf4VPJ
kfvoLuPlfaVjN7ZwKVGNedfFFRFUeuN/r8g1ev1lDeOlmn1+sn1uaD5g9EBdS8pJ
aRRUkJ0exZw/glxU5sD5h5b1v05MUBO6/pErFZPftdu+CnVFjDKVUi3QPd0QU3o3
w4DzMd+UJS60KhgMCq742xV4L8DEMDmkHYcJ90BHmQTqb7gp7nGrC/rwCXVdY5V6
KmA1KVr9ZAobRtr4ce4tczahv3cZCrEf3byP2nZJSk79feYB9V95CZLA27bXJusw
CuhyztHjqOJKlXvoG3g93BO3w9WZibSAJZxfFYV+G/PXLql8EewopSQzw3XcA4cT
IxP7eSH8+ZTdOXfYP1ynAgVphjLuwu9pUTw+p9Q8e4pxIYEt1HxM/Uc/CWuRMDZR
CosWTCJDKuvU0fp8mmoP4De+Jz3gRksjrP74y8VUQR6NiFiuWrJ/KOFzp73JHfko
oIo/usBT/AVtaoYSR7JqHIs6L+i+D4JRtHf/h6x0BvMPdmt/SJ8hnJ9/U1C5cpkV
+2KHqGVDcTPI1vFBnkSYqGtDo3j46v1wZrlkNiWLSwAbfioo1jdsvZq31SjjBCei
QzKnVvMCJTDTFZsR8TZJeLhJc/SP9/0SskJsS3VEknhZhQFqtqJYL+IDW4yEAQWu
GANYC5dBXFBgMe2aqWm3td33IkAlvmw5rAiUtQqsqCv6FPx6bpZKOCKYd3jOqJPN
aUrnLp2vYNI8xvIGxUqD3dCYl8vOGvgqiK0z6d5l7caYd68PcZCCe+MQDkGek0Zn
lxn0qZmxNC4QjAQZJLrG9xKVORtdRDVWgVsNwUrGntZeF5lA7pV3/Gz6cEug0Nas
pId5NLIHody4BN6KdbIu8n1jL2c4tc+vBGYLhtOYFKLX+T+z7IDX/+hlvKx1xmkI
12c9GObLHPWHA2uMIQzIyPNO2ZXOiFB9SuScNI8ZYUeCom3oUNQN3uBoTqoA0zRg
aY9AIWjl8+10DabZ3tKtoXNLY/CaxHt2Dlgm4TdWVfe1MutJEeAH5jh4Apvg2yyi
jtUarS7qpPgbMTfF8tb1AGoMyCsGCgCdtA9uvZhlxHFb9AiRfi2lGNNtGMa3Rskq
jRTapQdisp20E2PX+6RHHD28H1WnZLouSpj7HqLpyOQHmlINVLSCkqzIJCYeh1TM
5NdDVGMtmOV9ZYogeruhlB6oqtO2WXHtv0V4TPglnRWs9TzI9GGAobjyJQV5tu/G
shPu9r5dSjZ2GZBZL0hAUWiby8Qtr4OvgZspfPUVpMAP3O/UoAimQJKT0bMM5kcu
4b35viuHYE53vJqjfh41VkwjFXhYldq+BE+apJJ8dqb2PpH8yBp5yYKaGsyqCPFl
taGQzSvvDcrPKN+COq6/l3whtUQML0XaS35ueJ9Z4e3fJoPaCviPSrhHlq9nXpmR
E+pQ9AtzcUah7ovPT8VYCicUciES88jiFJ+uSnS6XQxVIOd+P/LZxFibDyytQQx/
0EXVA79kbXGhodmtcyp2Boy3E+3hq8JeWRY8nWSR3h7IYer9GnMdi/4cNjq8P21U
9ULjF+n3F3pLm279D9lQMJCVDkkQhgkunDt/ZLXQlq+1pDUUyFxJLiuQ4cK9ZtiO
wYcLrjcHg2PSEfA5vqu9Y9onxebCfd6HBZrJC4kqIITYeSAei3JDq4XCNvJ5dgwI
mpSdimyH3E5lu3PcR+r6T+ikn06L41VudP+BoeyyRGZaFa+tcO8VZ6SELbe8FKmI
bflq8kazw4g7ruFBow/jywYSoMmvHBk7G8bfCLts+4Iu0D2Jn0Ha6ju+QuCcUXjF
MlOMdvVsD4QZCnYEh6iCua+Ab1eusVhF3or/2AJkecHScZ9ll1HGQ6+b8QG6h9Wn
kOq9cwQ/5V4noDDNQAwd34iDE+rDuwN/qhiWHPjBXk87jK1Hu7LxNQb6bOTmSxRv
KVXWDiNJTBhUJgUd6ylRAZhefdX9wYHp4LoqAylnOAkmtVuEEv1n468MXnQgnlUd
qEB+dyO2VXf0caGjFkxifRgL4IsRz6t0nmBUcyj3ITQwGT3h5pLoTBSWkmgMRZNp
gSjNfqjdYte/Ylpj2VAqb7GSvqnbkByjBL6r/olMB79K8K6S2zEWStdSGd/m1WLU
sRqVjFRxveAnOsiNRsoeihgxn45vUjvEiplUgTz9arjNc109jlD9bv0bLQvxwW0p
b5Ru3gVptpqcxF9sX/uW6nwa27M3YT9RXis4Wkx0MHB31KrA9am+4/80Hf50g6Ux
av93Tr97zOLsEClzG5w2gknRrp65+smzw0opphWhscf7ysmk8A4EcmbMz0EcHVzL
kd+OOqnnvEA7HlXt00cROj4m6+mplZKWgVaJUPtA35AsOwRVhCwkxHNpb+R1LY0r
jr67yxBrUsCrs3OxTRg3H1RBe/HTYMQ+HTMmSsWj9BShAiURTD4JOwuEj/JsXCRK
x6dVbIoWgitrK0KJJOo9H9avLq+8HgKrZuHTfiKK/5pEWkYd0D0FNZ70ksSLJtbD
Tj8NMRAmd1P8De5cQ1YAWrSPKhbvhate/q332mpGenSaGDTGXJOdqb8XatVS71qS
jxgFN6eGc2bVl20Dg+L/pgLIeiXEIf1gNfj/SnGuK9uUqtSUYyEjeWmyI6KAgpUr
jZyOd6UQ872mAeHKQs+QKtWxNnEpxcBRQipYsJYv528zbEqd81UY4SlkyPqNV9EQ
+ruCJeXBhRc6FFfwFHSZoSmk88sjibg7bUZcvlzNK1PGNaBXkS2gn089dQ8IUZEa
FA04pUN6zcz+CVXTkzD69N8PNUgdP++b/0PCy1mSN4+jfyPfXRWgfcEk3eaakEnH
YDOyE9praserNhSdQUG1bTG6fbxBdIlH/P8dvLvl6l6uI/+4yX3OqCrFIJ50wM3W
yr0yh8JxTymB1tPfhjNZMPqn6JdVGJ93jwcus7AUPgOlLEt6sDO+A1g8Vhk4dkyb
qjQA9qSzX0wVBvdXBAmEfi7bDcDMQM2Gy3FMDZ8QE7xEWwzVJuFECtXFMQWTsFqI
Qr1+sPDBFCFrczC/C/rSgUy08+u9BIoFW0AEjCOGY+2cfCPmffqoHhao0+ADuQCT
vCxUlDdWjzFxn0x+PY84f4NhD/sV/zt64dDY64lXt8BiBqdavDgK28dJaAS8JhY7
Ew7hjF0sRBpitR0CVUkK04aHPnsBeqciOnsRJ4WcOixMv8qwpMLFAJ0/aJkyMT2c
lWSUIFGiLKL1imV+s1s0kVGv+LmkRenXhW5t8nBhqtN9L71YggXHWsYViwj7JsjT
9vyKITHMdN8K1BDICwGNF75goeOdEviHjgqQnbvIrDmG5ZXvGsAWPZlYYJE9RCoD
RHVJfap/IvdYI0Nd+B+c6NaakdvwpC4Od49haIvvmGuo/PsfoDw6cWWPXc/++arv
FP1Q/bpUhfecOO2/GAsTS5mcqGkAiNk5yGanFoHpIDhHYZkVggkA56/AaIluAEod
PcXO0Ftspk6mAIIJACXjFVO0Lw2Iva8bnR9Vie/rvG76KBvp4WgTOmIIJ76tD6H5
viEeCYaYHIguCF2t/oiiX5cGnOh7720krcWAbSTsA5ptCPj+w+Tpdgvqh0v6dC5V
I02MHnVq9sU+1ouXWICpOwjXK9r+S3ZrU7EquZwAFJGoT0DOPOgv6D261MuEew+U
dtivogojqwsk0GbjchXCKXklhGbQ6pzy0kYksFaPM14YPnazkrv4cr5xjAyeH3fI
oKuLk181sE+E+kRYaPcQQ9miXv2Xb2qkJI30GF2KJTnAffrYsoZ4d/3eRM5EfdiG
U0ifPvqxlB3s/S8TZIxZfNfDOWfdZD4l4hzqWp5DtnzMKvYbERjNJkiPnfX7BVVC
A+Fsau377hgcFABor0/n8fBeo2La3nJCBMO2/67n7NG4pOAzZ1g6JZuMPmIW7SXp
qv5ODRnXdyJGmR/fluV1SdAfwdUyq/glpw+Q18JIhpD+mr2wKdRk0b0i3VwnJv5D
H42bF+L5o4ydvFekRCU/tPFx2PnTxRuhEmLVPRuiGRZi5lbA8jNev01JEwDUoygJ
um1fNp7bu5peG5V8uB7BWW3tCfJGFYfHSfkoVv2U+KuJ/KhBpMmlPP+UXW+DU/59
3noB0Q1FMdDoptZkGGkfaByw//vdlPFJ4YuKtc0KPAZtmefb1oIbXtQJRq1Hii61
JlaSuwFk1NetiH56riZ4xfyKrCAZ7yrYK5JZbUQIwkRo8SW85lQD1Fc3pfhVlz/b
rkLaByEBWmPB21wGg9K9qZxIAoxG2fOsDCmRce8Qeoi+Pf1TU5pzvzCSNAyCyBOk
cCyX8VG770gOgZUEVkIZuo+KcHa4g2MQw/2GI3/vJs0+v4yfFqm1u75fgpcJqGOr
2N0M/uMqburfjUWB+Oi1pwam//hGq+1Y6vb42mc/WwJTeM9t/S4eu6aps8s9iTnT
DptGmjOyJadAYA4yXxPwa2YfgdR6xQ1LTcJ0TEkDlhYCAZ9wGpnkkl66aWlTKVUx
X1EdrASk1i+cQQ058YK+NBhwOeMV+33OjeY4M++zkLSI08XrHQBNFo6B4qIQpijo
7ggk6XihCDqzK5tZPShKLHv4KPctdexWeiai8gs3hv53zrCwHKjjNB4Y2E34xp4E
Ll9QmJ3Mq+j6zklbEl9AR3aZTX0EAqr4z80tSiH2kYS/h/xsrrNeaMfSnHjgRgZn
Bf5cAIAprzz+6zAW63sUqV0j600fQmPo2eM5zaZLnpl95YKt2qhAkxmZ7S2XD7Xf
vqcQwTmu0h02LUaFMDRlq9lcq+tqD2zftThMLf7oEfZxaAFTYjcWgBdG4zkrLxR1
m4OKBbK3EZylgWU0EUVYbGBq3g5uiq24biOHLBLyM//6MJ95zFRFmzbyyDk+3Aj4
GAeWvZns8NZT4+QTjrTMTwTtsuZGT9C9TyW8Sb+4KD6tzkgmHGZELytZiqq2ix+2
xHdA+fam4vFGSrOfAn9c919rjpyLd3xEvc6IJBV0Cf2Gakm3gJEuNtck7bdR1G94
BMm3XgxMutPBM0pMJdN1RJjVJnKUyKbv8VUewv0Ue2H+uxKv3n3TdjZz9jjyt9Y0
0kPPtoBwdtweNqHJcSPB5Gc32SfviQoCHxtIJAaPBXZpJGWxE/p5NYF5j6xOX90N
Ge7hTA6p8t6UnKKgovIFcuTtQUiRkpDZpzN15SfF8CIaaqY/UZjBE2xUJVP6yeUP
xqDjrJ9r6YgSb0C/KTpfFlzaGLsY1AkoXrQ93Q36zUoKjze+yMRNdddFjJXF+eL7
ePlROt8vqXBLE+kadIIgFwJ7Tg3McUAjVy1F1GydSwuMOEZnxHvI+tPJC1K3nNwx
srfizYtASbxrvKFY/pMa2uQC/6EwuU+BXmP7N6sAo7i5lecJf/nHaqxI8oLG6nYc
w3p4dCNOfC18Jelvy8jlDzZ3eDxMCEMtWuFdC5/43e0ol2N1nSKjpAwKkXFhKD+g
XUD5ILacIX/iPd8kvZ51eWxiW3Qpj+NiS3V57ZBmbVMq8sgMvQ6qIVcERrbLwfTV
6VnaAgr0OVh838tU3JqXzsePkJEY1oWFoJeACvrjH0MJN/Xpsy5oSKIzDzRYQoUj
h0QAnEBuMwxjiPhJMH3WO8zOrgw3kyd+Cb8nVjyMSEnVnnWs/thQBFGNrD5XwnEb
mQJugnGbyvaKJeoswqs95d1ugR7Su6SkXaVZgBjBIaJbFHhAnVLKY2IVqZ9LdWs+
zK3tp/D8h2JdIgXHFj134XdSxG7yyIT9kPExMUIuKp6E5uui87ZYmwXEafG9UMX+
GKj1XAPpDykjwQ0x9t8oqY7Tca4j8YHKm+ZFV68W+LO43HlZk1ls9sK5Z5u5pPlj
lJUODM1UnW02oXZ945m8D+crXRUWgok+wXgZT57PefZoGf4S2Ey1TOTWsvNf2XsB
creODHf3V4yDxrD7X59E7FYVnuBXKVULX8NTMuPOt/J0Bhbe/4RrfakW7w/MzChP
do+EBAPbwRkDOmtYgUShIC2qfieW1Qf1tui7nTVvX2Dc0l8QllA16r9zfBJsY5V+
RGn0XJh7lMMAj94laVaShHYUk00+1i5514uPJ4gMqJTf6mzFLjjOQTUSzBqu9Ou8
oDqr0BCsRW3lWpaeg2uZOd7oaavja1RyjuKOJzK1s+fVEBp0Yu/NrB/TW5g5MJcU
185Auuqk3vT1p+j4pXZvqjsz17R1ev679xsNMD/0onl+BirrmVQHhEtADf7GaYC8
FhrShQvVe6HQ/a2wpFnqdaMvCkH4qRiL4YsoskBbPAzcgWWcEotRYwSCneVPZWyD
2nUK4RUe+YRV5Cc9845p1KXIstkeZvVldFgs0/jsFrhjlWqG65GDkfdQS5gNA0+5
iih1f8HY+Z9DWl8Pen4Lu0D4IufnuZi7QQWxfq8aEARNhRtiva3SY3QvDk+qaogP
YJcI4yyJPc4SeJUxHUixsEiyCVU8reXVWMaOqGZN0Dy3pO0emFoD3d0gsDb4MGdD
7WiX2XQXK+si2pGTVUo4Nyifk2H23HAYdTctjLc+zViJefo7wPxI+qU1SZGh3IpA
DIXa2ah6fiic39ugfpbGAcQrLkNzjleOE77qKMM0PRU1xXPGwLBcj7K8fWZArB/p
rfahdDupDtyg9Cj+gHTfjdQ2wXp2ipTOx+/aixMjADPtdaO/xcjiYoSzSxsW5IUy
aiofkPDC5lhfc/i9jQO/x18MLVpb59hMNCbLv90SI7PXxtc8IQlebsQsgWwmRHuD
fT6A3mH/O1Py8GTts7MSOigbvBk84MpH3J1jOapZ3IeQxCOeMyZn+GpENcW/zwyi
E718uEok49D9jrKSHJH2WFqmCIVJ3ho2UcYjx8/kApWdvrStaEmWdKnn7lTYTg/I
eBYVy8J4UCrUMoB+xJwGek+CwMy/KvBalGTxMUBlQ5b3xr1I6c+3MVYe7Vf9gQbD
kuZdv4N+UuygmjnVk23IWQ3YfZErBYF4yf2hxuE7kcoRs6CdYCwYHeoT7UF/sZv+
hYrY3PU0lOGKSQhqzrJwvJNgHIJLk1WixedQ9D3lOuXWaIGpn8lYBUeCsP3bM3Xe
bdRJrk1n+PnCF4u6Sd1IIqN2+kRXhNR52t9dgQPAm/xO/zZ38QoyiquonRbUV/hS
1zMmuCbuVjuVIQttabRhm2g/IBD82zN0DnTdeB5b5VSmTGctHzuvSTa5vZPyaa9j
kViJUGOVAM/IYI5KNV/lJ5cilYgfs3M4vvDsjvvt2YrJS6KBjvE2V/TZw1ovTdIB
+NKhFb0R0zYLi+Bt7Fe9w6Gk6Fwuj6XZvCFAZT78KNeUhTvcDHhZZDpjl8UvhUub
UTG2uOpOI8Dg9TqrSbH81Rqp0Zj5W85Oqs9poqE7BoSVXqfcK+G+QYoZLWLsKz4J
G9f2jo3FzNlJvhs0wjtR7SawyCHYT6rO0IaJEv+szwOWLRF2xuWC17VJzwvdqhb3
DYnayzfPdEFngbEzW8upQseb0ajbPKudZkaorzG2vmgMEzHoW9c0jUH3lbIqhyuY
xvJg8wI19vCKYmQ3XdFgJHfUMhy2tdHTLl51qKtySwxsfhzcKbCue8Wj9r9eKBBD
je2I8Iy+WUPNgAKzPfgJZHfAKr87T+heSehIxbS75ZYDt7k4v1GLL3vPfBQO9eE8
2T1dK7tjm909/+3qlZL2Xj01Qbw00RRcBYrLxJAnguq3jITyPHgqKVOKwgFJEIvi
O5uU89S8gEumMS0gXvV6rF2adwJhFXViE3js4W1l2GaTMblsIUbElcsW/J/vtir/
Zeh6wbPAVHwV8kkXoZeP654373xhRMiWnI9ieVyJxRhJRKwbKsx1nliYKtoInCbp
r6IwQ6QpPQqi3ZAUOc909abFSXj7UaSd4RevvHLLARKJjJQW6hEyhBRBKHzsbUcn
QgXwvEPobjnWeMeiv3lVbce4aITNj93v1lF4t5YlgbsJbDTlLIhzd82uxrjKWKvf
SUWaME6QVMPu1Wc6UBSPKNQrFechLDwBF0v7cf6Hl5jF6n59tvayO/6jM+blc+Mm
INjGzux2gXX2mkYKJG83sDwg3sMvCgMk3EMwS0ttqHFHBQRPUTLDURxr1Y8ZjDxO
3VkW3OwAYcZqELPeGb52EvuRc9H+8CY00l18toifEp2VpX+u6zQo7waClhMBdljf
2qkvmXsfieMEiTqKI/x3lBeOcrDt32HArX6VnObaJs5gcA6YohwIJOBU8z2PWF8Q
vuOwekFSfdqI2/+rtvSsAmfIVQ/jslpXf4DXcWfIacwSTbBSMR4wQngZlVv420rQ
LrXjMnmCBduTfegLnTwyEr+TeVTmsdgZZ4fKz3GKeTT+2EwJtMAsytT/Cy2AgzOK
tYYjXnzokZ0TfUoxGVJlbivRxXseYEzzDCsMSplwRcXQb9SFTQx1q0b1xcCfb2EA
eLZ3LEywb3RWSpGqoqYQ+9tJRvSTBr1yEo6UFCdQOtfOjA0EFoe/i/K/NVEUn4Jj
R0gd/WuvWj70U98z2FiEBL7ObmWjdl3jZBaPAbgdheb6goCEu/VVN3CgYYgd48Qa
EdGEJnu3h019cYeAxtWlN2w1oI3zGrGVeZes6zvO0ETBRcMnMxZkIS7HAPtvUMtJ
i5Ua/hHKMpB5xPPM9G9ZVVxEWpK+qGAsiQHfBV18h5W6BBjmZrjM2en4mvhHfGqa
HrLF57xvXj3I402P1oIaN/AXIV2SVl4DIAaZjxVd89So6lp74E+LVYuvK3HAsdRT
biH3rZXoid5rSozz8SrdajxzAYJ4L4TsAOvaA5feYL2GO44gl0nzwTzTbRawAK8s
WRNJ1k/SeiorocjKF8MDJbgZb5bkwsv2xIN+YXFuQTrGk+iACljOUoc/GfOw9mKM
jv8yS8kxNF9iHJCHRmm7Qn2MS30/Gx9+w1bjLH4bDAFaFHr7TLTs8o+oYsF3Zd+K
XaZR7JhlPc8yeN+kumvmM44dXyALFykMrx5ab/jdS4OsA0JsSuTColglhvlME3Bz
HE876uloKhrBTiBf3zZ4JJTvWSYIUM1z3JsxRRA6qAlD4L3ZDilmMs9ZiUtuIc1N
xLnf4CpldjSs+7NfJT+sVKbGeV0zbIx2ZlGbEDb7hLRCRF2WvjYlXT1XjcPm9NzY
C5IFR9qnQ87T2Xhc/yB2Cpuc6SKlx86ra2JyYf6lUtYB6qs7+dG16wzL53z4mlKw
ISzjmdVNVAOJICm9wY6va+Zyv5NHO/W+mMDZQ7V3dN8khK6fqAc9yqwzF0f36Fe1
qItSQqqT0/BCFtphuFTijcymw5TzDcv98sVHtsRuFn6xaWM8Y+wEzPwZnK3DogrC
XP36j0JkypF9wS2HZ/bb34NfP4jTbm75syFuugKhK9MEEkWIvFqNSVrSN6HFs4T0
elMGKLgspK3af63zJpbU6+wa5E2veTCclDdlNEIRb5NEZsdljWZ3te4RcOlfDRD3
jMy/oP6/OW23Yi0f1tW3ryWaDYegSalZxQ4dwPgpWboVaH3/5+qHJDSQmIUGXO8G
W1mZQjRot4kNRWcbpPrrzCboQTVXFL9foudVDpTBn0HPl3Xlj24yoMkMsmrvXHNx
7h3RwKYTGm+zdIYmBEzAr8Y1TfoJ9bJ9llIg6m7UKB1hdFhEDCSJyRlduMiZ9uNC
s/5MlNiJZ3JjoAg59qZy4B+uY5LbLhGLg7EIGKKzsOzEB471JmQSgTiGMkeY+YB+
RyAJUg0Boi6ipNi8XMt8cgCVC29BlJfATI4w9JTWUxFzGvfF0vilTCb3g0b6aUUz
y+jcHMdL4WRAWPd4itcnFYEEQbg6M0VhraBS8R/27k0iZsSdc3RxWVc9lQKBonbU
40FiwjElJ0PYKcxizdvCZkojG+GpHyUwe5ZCu736vW9+9icqR+c39VBMcGHNG9rW
2/m3zGlf+thtb6vXWiIfiSOFAEwmDWBnJr/nTdowMciJMQSJkRG6eXYY51yfB4Z8
f9dgu67luVrEz75cgrb6kQoiEOBH8fGfpdKWrsfkK2ziC9ZBtwcKBhqmlkit9bMy
tEir6p3dS/R7qyV1fBWx5A/InsiwZLv+PYa4p7dx8qY/0pLgO+kXB2z5fsH4Pswy
WCo0OhcKnykoNKhv3JKd3/bKeFbPFFDC3NzKuKG2MkWGYERAoJnHNcFFz3dsAohV
wtA+l30cu5eD2jmIRjoalpvFOvd+oejUFa+l6KR4QErWYsR4C0O760vSj4kwomyF
KMQ+NvXNdMxaYMBhkcwF8tcffX9/dw3vaGjo2+bnpgXVZ4ROQjtC9n9jgmswbHUr
hr5yayKpgjO6hCpyoigsZS5TnFI8NzMzXzMK5GMMvjj+651ZxlEg2WXMf0YlZ5pY
KxZPGNcHeD+qtgO354MBrh0UN4sGlxY5MJ1gmsIukpgUyKPrHZjly8aBnsHAC4VI
QVDjAwMY05KUBJdBs8FI/eDrFVyiU6oLFdgkyrE5U/ZgYBdbX6KG1iEYYaF3I7NB
GYF/LC2phbx6ODdqOAoQuAe//A/8Xb9oa/MnHXV8ByzlLq5GQAAm33edCrjV4pnp
IAwBZ2r70Oxi7KF3s0uIEd+rcuA9I6MyizghrlVE60D9B14AyYVBhQ3gyFuYhtJF
u6bCYnBU92X027+dl7yqZZ20Txu3cpeRgP5IV5Lzfb6I/EEnSqq7ifdT5HhiBda0
Tvhrt6exG3G2I50RssI/kz5thYowvhhU4xIBMOkMzlFK4AE1p8kDu7c3gL3mIT58
3x4k3Hajy3SC7NUapBYl+8cgzZsNMxmLN1/E9yAvxx+QkZEelBNc5uQRNfejntDA
PkII/GAWA1Mr6vWYw6aRyyw+bD7W2zXztJgytrGArGIf74vub+lSf3ba42A0903C
uUR+DJQa7LZcQJ7r/vC+7ZykqtGKOSXbPsxAni0cUxQNp6dumJzoCiHO8POpvYmi
SD1n4Uz+40Dy7yJRjF6xCAVA3lCmUU3PZrOJoIvstxTCG3PNJjHRASWC3m5ejMhl
5LwqaoraYLHeiRYFIDIWBSh2ZFqj2hWuItI0b/u7AY5e4qI1OcOJa6BUSxX47AYc
OU4xqRU2boyHxPUsnVrGs0Ily9MzqgN3/6h2ci8AfQbBmJz+RhcDRrJtqskUXQ+z
Tnz+7onYiZcj3B1L8SOn9Y4IQCK6ouof7Y2me/WFYtzF7nP3NRmIPWM3S+G8yJ4a
jHjB53GmOpUFcYUa46P0IBGsg8NSWtTY1lQLur6NUXKSc/sTDAo95189W4pMHVdR
iLb8+PXKLLAxNHKhK5cd2y/gg9hZinUtlYXzUDX/bu3Hp5so7xDfeYG64bfvt3rA
zIe+k9/CEoZFc/CvtgJRKlfikEbE0pQ7uqYoFqx4bpq0LEi3Op1awv6VslvX4Y4F
74B94npjc8CMppOCDHswetKyrCOdmruzH+oKaGhwlh+fJ1Ma7UYzqM2LgyOHDFQn
5oVEjDLaJexGXweN63Y4t3/iArbQVa0Y4JSiDsITakbSFs9gidcLd4Tmw1aCNRSy
Uphnfv3zsI3dhyPRzuvNm4Qr6eo1gitRpRQhCRlbyTJipZZYWwZPOQj9xwuMt2xj
CBWfrxr/KFvvbN5FygdYT99gNlH2W/AKYe/Fne8froOZsGpAR0KXFYL9oyVQyLaH
Um8PM4W7yCuK/2ACBj+2Y2o4PtbVqqCwTrZ4aw3U6N7DQa1TfY3uJrx9vuxv2nIG
uuyXPSyxuB3v46WsyqhI1LhmayBgW5WHSoDgFHE/XLve/ExErgRn8oxz4Owo1mdF
1FzC8O2RZ5DROpCvMXDtM0OVk6uNxw1J3OOePOgfY4WsjsGJO8QYs/InqVP3HzoX
gh4gqagRIkstkKIFimRSZAjNa7C0FaHl/rYICVcao+loi4KHnMHCDbmW6BJplPIs
ERLqZICilw0WSdJk2WU9pe9+1JpBQx9/HW/qmOHmAeshnjdlwHbkCMS2e8UCHcBW
bNOR9r+47/ayxzZOcfFOp60XjYUhyNB2ZyEUzXE20g7o5nT+W29A8HnqmMy3RmUx
ccyBzt1IJ0BsPP+mY3AbaUi0HdZgMtOId4nNRKHypajP/pOdz9dPsxDgGKmmox2f
I/yeZONiX1l/puPO9QS5jk+/aitBJ71H2zZAxbeeA2QNiweQ78QvtSEPdgeW8QuI
YgztE1pBh8dO/LNBjy18Ljl+l5ixQtCzCp+0GUdVX9tSbiqB9HhBZZDBWVND9Psp
+QVA3JiHF+Q4hoe2eCOGkkKm4unbGymVbxhl6aYdDea1SnzgZ9kD0mkbehngKAPS
nfsTMts9C9lw3b3ADQefYKFL9X4OnlgM4mA+Bv5iSdRG5Yzk2WZ9CGR4PwBVz3S8
1gblnOuXKZlz8wJghcslONDvSgVEj9c6F3kspna51EE0ABgzehuge5qWk+sbOFqn
bD1sDT1JVoRYuvSzCf5OiZk2JP2fomgTKJFX+Mt80+hD9B0hQ+I9eqW322/3KtvG
iOHNl2ROETxYas/vxKxcHujYUawePwcq7pp25jBaC9fQhnveCBDEj9H5JuI0VOby
HZXiueaYTw1aGMhzORxKslNtqND5ajYw3FV7ZX7QoQBZk+SHldYTZFc/9k2gWYN0
NaAy6sOASDZ8KS1f1KAGy1t6zQh8/LXabSjVYTqIcO61RN3CDfp6B9BMIVXqOqYv
Mhyz+Wc+2egRlc1sqp7tRPl9rwb/QbA6BlJCiIxgqxfWqz7chMyVadVAKGJ9/POW
kw44ahriu66OcbPkpQ9GyCEF6enTpwVAY5Y0YjPuwbNWtms7OeEPZvCDZ15E+bVj
b2czoFPd3YR4CevzZaevMMZvWty2lXldEBHpaZnNMIp02aj7etHvnwg55NyrlBir
gN3vgSGcJkFcYwIErDRUK3xIEd5pVRP1T0/y4IxU6lUj032fU/V+IbmcGoJm1key
wj5PZvDiFIKxijv9r7fCqW6jvqZm/r8MY7n8YG4lxTTWsA4JP3TR9CT5KIowZ4uQ
onFmVJ0M00o7hydql3Z6T6hYWdkPHdsO1flDa+BIyspDheFtL25IxjbWD2c0t5Xo
/G9vVh8WXlaC2Hr6AAj2Zqv/e0K4vsAr60efT2+p4D887kQmN40ZKGQ6KZs8XfkM
SoJhUaZQS0fafoFAUfl44vWCVN8GZ3c7FXiLALUabxv9Uxx+MjYj8+HUNmbKJpqO
sSYLFVDs0yDXxJviCmA65IoHeIg5ZdoR71jw93l1gEWhSffoUF2nLHrqmZaO4NOu
aFQOOgDZiev37DV8fIPBDc6BcTbGVEBXTzEXUn8MvN6+QWdTI16PzPM7EfxNRv9g
HonwmKaNRNOikn+L5l0FwKW7XDYlBKChUuC1+fFv3Xswxb4Oq5NaEXMat/IVUd2b
flj8TrqtWKROBITy7G0LHpUv5yQAr83bFoI++emB1jRXclMmCFRQ/p9tZ3UFvKgT
Y2cNqclTqejqkW+/uulYdEsXStybG5up8FDbOdBxsSI3qznprx9gLRXS0vzlWA8r
FBNCRshP4PEGIOc8mEH+wNqV1jKVfRHuIQ+eS/Ltnz3tC6Dw7K2tRM4Wbg39Y76S
87tV38ctK4D7eACzUQvaOE795N9/rSd7od+2G0RohYR6zUADThrdoldGoGqdOA3q
fFV/PGM+SjqmGfmeD9jrakwFpPIjjvqa2o9gvtiQn9969ifLopmoXlcBQAjV1JDd
r472A+QDtaqWGZ/VvnSUrR86cZ+S3C7LhbFqm5NzscwfLaFUGPhlcex8lLsKGpP0
6KgYLuAdvL6QQlcxxJgkXBvvVekXXakNfe892HhYn/2N0mUtuIKdOKoaDqEmM4pe
EUunive9f4eyy3SGXYEWwXgTNY+0fDAyixuIBzY8wny7D3axpgIR1C8w90MwpIO2
n7cvd8wYl/rfP8VPTzHtTxMT7aA2mO0bL2PkMfZMS4kbQD8Ocrjlqm0QmsWty9xd
ulqupUcnBhT4mfvyiZWcf5RglrgeexfFIWrT8nsFciFm+ZHsPMpUuojDQRDp5yM7
ZYuk25JZmEq9u8gjJkxv/GbWVmTkPAjXl34YJII4WcSZo/LVAmhvdQpCaOE69oHu
LXeUORqr25axK2drSbaBWlL54f0LSmnysQBtPRvJn1hbHtLIHCHjo8FGbhuL2Xkx
Iy+1Zad3a3IZQXUNDEtq8U3AuIIQ4e6ENwbfm6pX9J2uwBfrret37NtupeEl7Gp5
8rDg4uEmREJltI2lpF1SYLkSgLXGDlLib1Bm6Cn1vZ9gIHAMg6WW3aucmGb1MKDk
DVRFmINMt+6/6RmYPLZ+6KkSNVLRvnJ/fM4KbxbHpOCX2cE7p/KTgBYgnZZ+/Atp
vbOqjIBSyZ30OczgcWxZ7CdgJcYBJ2NBSLNZCB9mVLFBhHI1viWQLSQGN39gf/R+
j3VYMOQNOh6SvI65MioskGaj6YBnRRhRbnub70ig+HFg3veayDV5kMDi8JX3dQSn
uoceIPBVWOAhzW7z9OCeoT9bsUePIyFAHlhR7PEdUp9TC/B7JdyKxM2eBPA1uvo5
IgFAe+5zCbTfQyukFpRQzRTXlgncCaarAaNscB+pPJexcvDKxj3GmGHD6+fyKMNe
sRMAOaooyZzhy9QCN6eFhRuRMFfOCHeLg9nBypUNMIXbEmj8jjR1W0ckaVf2VuSX
4wNycfvn4m82Lts2BjSt1D1jJEjcg9oG1p8pqAVWP2aFuGW/jU85306Rh8uZbLWM
8SkQa19gL7ZYnZpe2li4g6xipBgsm9teHuwppiYE+aODUBmQlk91JFZunXGAokJh
Q1XssQ5J1rE6kroU2WSKJhY0Zf34Lo4oiKyZC92KFKNU2HCd1j8UYhcsTozFEFWi
sxAZ22AODwAnz3Hr+Xvwi8Dh7d4KerxGe0yI05eqqSxDj9vRZ4DZP4xYlJemO+qz
xChJdXUh8R6JVlG63hMRx3K3m7ktMlVwwCMAMRfyk9Tpxy42XBc8SE/EFpza1eYZ
GLT7CBneWu8dqZU1jtwfEjXAvDZ5DGxpLUMbZ3xrO/nRZt560h8KFmLJJrVVIJAy
gR4lqRlqzB6SFfmYI8X4phzm3FykAjQGDH6lG159tRPkwa83StKoJERNGPDCHOjn
3ML3sQLTufBjr1gwVmUnRUzyx1rHbWlJY7NsGexHwMr6oZCOL9yIWbUZu+EqREJl
ccl5wAvunIU21u2wBZmeDhHvPYhv1sLuCGUqhBAes+A4FZZEj6qs2Bjk05TmwYgd
MilOWDNyKUjw8EzX5KbeLSgn7K6xM/g48EIfRjBgfVKU1o9bGIRLLWV2ddig10MF
IBdk11iV/OjwjnWfr42dgvO6WHTJOxqwtHm2iUwk+ZMt40Zw0hRsqG0ZzK5mIQtI
Fu53WQPC5Y1SpBA0RIykao9mkba+KA0WF7gL1cvfuGHJ18zD5DHoCrjRB+Ig9rIP
VsOUvC+faS0P7fsUnxQqVBYPcITNWtm3ohA9DxG5uzHD2Gx/gHxUMTlRqivoOQCd
mD7rJ3Ws/g7uTVOeV/jof5hT6lhENrWEHKf/PTYfhhRrxgG46KixIviR1Vn2FLN2
ZunHju7h0XmhkdtbfFxTkYvQGrfDZl6RFfTbxaviCemaXn1/JNlNeABHXZhSVKL/
9E/YWV9cMtn+dVuo/isczSrMuPBm2DV2vta/sozTxXduy1gPl0WIGBH0IwUW3cF7
LwWuZCJXnFXKjbYSUGbrfHK38HMdMbxBzZhZyPo9goCemWi8CufCHOiD56zxKiBg
Ni5t/Q++bPf1/7I09NT+AYr3ddEhc3GZZWNdEmlz/W+CBqj/tu2FQ3gPzaDiXfQT
Ioolx2PBhadQ/mdE58l99aARRW81D2KvWwXdH+wCynzmenRmRX0bfFEagFxA8UDr
FlAUOgZ+ptqSurrhazOmiFMhn0hhrXaW2jacbjARUEEdr3Dp6zuRk7bvrnnJsFQV
dd5J8uSpA0HBstgnwbtcEhgJkQgrEDDLhjyooVW8z0BtzGJDT917TUG827wefbb/
rvEgenUEKgPIBWm6uTJiAkg8R0dvNniFnXzVvFFHSVvgVAmmapAD4nzld8jX1fyo
wJSQcRhJAWXrf51fkQBMPfLNr3bPSeySfCRjWYugO8jfobxON4ox9WC9vNL6cAJA
3/FV6tzVg3QUm0jC+9WyQA9IsY/dwk+8kA9fjOKDx/U9jXpFqNnt9Z4VDA3STUZS
KxVczWLLLgzSIwVP1MDMxSdM4/YsnDgJVCsN1BV3OLWCQ7ZMf3RRFL/dop47GTtZ
E/sDieFLKNYc31xBpkSWbNiWO2R44/CINONJfucTnnbw6yG4nTvtedWi6ZeQ/O6H
mp6chnPZEm13AZXCtdWNVDZQkQ8vf5Cu/Xfm6U5qSVeIjcSC4vU43iquREKxbzHh
YZPodbP3HRn6iXx7VUodDLS6c/6rTzCHqFeV1BIb/135RfddWRRbV/gmz09ig/Kq
zxQ1YYGiBboyNpQuh89Tbic1fYWEfriWPS5RIdfQ8WOGtRpEZtpNEN6XOKSoZ2+c
dakQDntVtCfYSS7EJw0BhDVpKx1t1nB2ZZgtPtk1UtE+aNkwbN/SUJtOJ18gmX9T
Z1+jr4vt8WqoOGV2UkYJwjNyhdvc6m9w9i9eI0bArJoU57mxNlfqvhMAsJ5CXcmd
Q3IupFIqmgywWyrl3I9pMn22mRL+lGMvdaF2c2KrIko0IKfWY4qK0njRyLWuN0Zm
u/8CfdutIFHSFwqw7MWuS8TprIwWd9C7XE7jekxp7Gh379BVElU1u9qCDztzHUaE
wFgyWv8WTf9ph9KXSnRIGjFTsXaVdxRSNiTYWEnkrXk804iQLWWHPkQ6qp7R2zUn
hIFFPHesE8B3w+NLDFiIMf3JcrCUQ/QEwnVXpzgaQzmJs2d1TNaFGEepib+byXFG
N1yyy2ObhEbvnm9WAZ2z1yCCJxpSJLAk5JQSvzPWk5S+OSeWtb9zVI676C9mnuSS
Rzqk6tPFczt9BOZJW+GT+LYYBTr/ameHm/FenM3gSVrTeVQK/vJMw4Ie64Y8CcSq
FmfKNFgnjOro8yR+qCAh7Ek5+ofgTQgT4LMq6kW5oEUvBvAB8YeoPVd7xNPrLBQ7
GIl1OL7OT+a5mJ4+4Yq6EPL3WUH7JReHiabRTprbCcudRLa5GI4N1D397ikD6xVy
OtRsK5ZCrnPQtoVmLorBZUH/CLJv4NhH1F+Zff3mMgNllxJlbjBqtctfL3+siD+Y
hb58feufPrmmvh5RGtT6ntwdXRPK2bzupJfkhQwhCuwZP+Njp6Dr/swaW2iByaUM
ZlGBAZjDBXjsS73G302gb2otWxzAKexdPvp4x01qX2ivvLPepKDNu0GVUlUzyUeT
1/5sTqb1mKD6PIRGbERHepz0aofHMd8bW2YYAzTdkVWecCfd3vYN9vrU59mtM6Ah
NgqFHBdCk/HAjg093LO/Vju9mi8fC5EEMMFoJCPN71SbM8Z5FOIVZxN1MK+JNeCE
9LW8OjMGyE1b5aZgY2OiLiy0XTcWQUB1JJvmWRPi6fnVkPyzq3PdrD/ZTuY8n+T2
FBqURhf2i4AJm7nM7w1y0liB1nTfqClVosmB2mq3iXZuAUXZDYzQawi+P0an5zHy
1xHwH5lEIg/BMyyFGZZzm0TEK/GP2fLh20611+pIJIEGCfonh2GhONk+uZUJeu9m
CJQasaSZjivgQ/CI5HFaN1fMKGPFGdLYNfkdw9W7bp1+dtV9zqylJ01zed+h0CKn
2Fjno8OLtcX5SceBGBwRMlWxEq2I7bs6yalJY2YVhsWhhl5bhVdxRsGDqhPfpEqI
Rp1B9DkCEOOpihBxqYdQ9FKvjOslVApYahwtcy3GRRzi5GCx//GoN3HdeE9vMV4P
pTin1ApFQ0eGKkbfjwycbO8QUW8n3oD4aldwuNxF97TYOfTxVdUD4ZyxpYUWHKhL
TUeAwZmLjMNLLs6gN2Jm1KH4FLgDuNQvvFXDH6SbUOyXpoiP/wbjPLgQv0Vm2ceB
Vv9BARmlUgLu9T86KSrylyQh8yWG4YfeYFzSUCjO8RLDU+fLya3LxQkRNsWJ3KAm
LiTGy8fT7bL1wsK/mYOYXvhM+BbXnW+fOsuTcwcN3WDAFqWkDhTGmacuOHnYIHsV
cIIIzv5A38pPyHmknU8Mdcs5TbL7L9WhX+BIPu9PAXJSYd+rfssmJJFXWWAYov3j
DVAL2KovtKzjPgqOfCIcD+0V30lBBCjzQK4XwE5sh6IPCZFhJjzivsADwbCdSPpe
MHCKM8ARGZoEIxD+0nlFstoZ8Zlv6i267qtJwEwbR444DjsgcpuRw1MsL5SU6Srl
2BPDwqustITkoq2AS0+6yYWsZ9B3jFXcR7p98s8n9lDvOrB0IxsF/Va+V9YjAqQU
2ddz/f/cknP8qRzUF+NvFx0taGMR1pAxsfLGOPKH0AfzIzf7GADkVjUsLCNuKOk7
CX6NpzVLftYLWTwNIO8I56FT+g9EvdVC/6taylESpFjj80Y36Z1Ijn6Jd7Irmjtf
QJm/SrSl8S3DjmUBSguU9IrHTiEaHVJ76LGjs8ZuP+z8OniGXFMQmB0M5qQNhxzw
ooOwe4XVu1/tL/0yE7E8ZFLXzWqkP3z3Fd8Sxi6v7DauQksYg1SiKhTv4E/MnsLo
u3R/X7/dr3eScpMA0UpuLFb5bhOTTYnE44PTMeGYoaQ668oOzLEev+p5vlGkk+oj
MritjcUBi2pCWQ/AnzT+cUiTkHk1tqmaW1kCD3vqZjqn11wZ4EeyDLA17JfY7U7r
0KLj4fYoYH+phzG8n8zoL2DvoMtj1U9bwP97wyay9uKfNLY/PnrmfY4hJZ8Dcg1E
EQjITZ3fsDfo32THCMnuJ9b0/jfHNJY1umOVEJ5C5c5/hpjJfT3op2ujH2K7pXS9
apY4QKIe/92E1vLmUIkJ722SrHFQv3moiXkeuXrP0Ee+5E89jyUEJ0R/KbkE15hy
Anqe11Zg4d5aGtUZTuLY+ujDjwoBf/+ZBJ/Aj2QSPAgdjBlwCB3SbecwOK/1ERx3
t3+WxIrXXrjvM5+IZmoronFLiAH4B2CTI5hxrBJGodLPpCPwm1BHdS8A5cSIPzXI
MD0OoVGsOvqjYZwdKZyjgLFOIhtcnwjQ9KN7huvZRVxYqUkHVFy40c2HkDSWZPfJ
mesyDZNuWf8lmV+yKB1n2Fb5fmwx2jTHYct37JSDm0sSUQNe1TDrms5s6h7akzSt
arjHlVhzAPcCIT2vu7KHnzLJAdtC7R76X6B6mDmlxGmI7xDYo3ZvGJfeKEgeDhRH
U/HmKWAjf5qpYty1G3RW6HciYiprDnGdpxwXdKn+vUy/OOqF4SEwImsL7XVmQzk3
R8bq3LR1N/TVJahbpO/hXkSxKN8AberuJ+7LVdMmgCCuWFaJtPxXVBOZlYyvNuZI
Hjs2XSW5ctLlmJkodRluUr7iCbau2Pc6mX4rRbY+ofpxqSsV6Rh2FUj7cTrZ/efd
lZ3B2vlAGUg86Uu3g1hPTf8EhGV0Ifc5YLx89YQfEwpaod8qkEi31ePapTulo+G+
Uo+qenOvJCDeYnvHxFOOKVoBzxidk/sXzCgcko5f+qEUaPgheizLBeuBb9AWFleV
+G4GNg1a4DBhMHsMTw91yjer2MJErAgJvMbBVXQLH30V2jZB+K1KYzx+S9vLffKT
ed4SkdMd2pW2MPiYloemICrkkaDA1dHHM691DSkXQ00vN5Ze8wcIRJD5yieQJ36s
38N8TB7iGiEprqt2kdW/5s9LrUSgTfC531nUuCJQQfK7srz8VTxoy2cO1qgjTXXN
w98GgugGmG6ywkQNgLpZFrgM96RF29OmSfbTKdTKir6AJBlKBO3Z259sKcHL8i87
XvurL7lN7rQ34625gpSi4uDrIcdl3rBqFS5TNpUY7Fz+KcR4BYuNZHLHhrE3OrDx
WmOpHhsnv9S8bLnjlQaOLs7FDs24rkEvhnnCaqj82KyDShv4Mpyd7VJEFWN8oxjc
WKK3Dp8zwfnMlIfC4P3z62N4X/EdOTyWpwWo9FgN+SWCrvUPLG41rna1K6nXiswg
ltopK/eG6dkll+mFlkGaEcSj237USfGxvOn+gPOlOgs0RHgUlxrbFSzg9WgBXaKi
rDKvq1HnxJiYoGSRfTOzm49Mnv8Pi7pe10un6LWYCb6Kl3paqKvfgX+fHX4zhO/2
IOw+QLqHvul3/u58ER4pf3P/PBnK0xJMLQ9DICyqUOigTT5e27CPwcZ6unDhZUtI
unkIdJduH6pqon0XhPqokBTreV+rDM4wFS0ED3q8wgLo2lAwZMGPAakDu4onk/xV
rsGLl8mlpVubZ3UHgms6Rn1c0vQUxuyPgfY0SRv3WMbekGyr6ZfGjAo8b0m/xwJ5
KSTHwzLd0KQ6bnWP5byMOtmCeOPv3OR0SrRPLCdLWBZRp8jqbgmN/5Poei4LAZHV
bNC9YHJBru52EH6y7nQ+75bW7YZafe9CkQnmgnSlYnLVf8PZz1gXJY+xbnYb30Th
yuYM5jvF+a7SCjk4M+UIH2iKIWwb/ayg3hJ/5Ne/7t8CO3TFMjgX4p9vR+nlscB0
pkUY+mcCFFIbeKuOldk1aBP9l13xIOhYuL8lX2VkJV2Vf4r4cxnktCScsqreBfmA
SO+Dz0x0rz/O+DCUm8WLUU84bvGshxPlf3bo5KdztTUI9Z1aRnbsDsfX+eLeNOvN
NUBAVS+zpnRU6qHI1o/i+T01W4KFyVgzBbc6oQe7+prSePMQw4WDP0VWj9gaRRas
MUIldygkBYmdGI3vBi3A2bBCNCzlCP/1MHqK84nt20XV7LGOOkDFGQtd8+h9Ml4L
HurV/+VPyVsxvU4OSy8zS1NjxFtPK9CRt8tLcvbtE7iKK1xPOH8FHWGPEleh1/5W
x/qXF6XYCfhziRCl5nVRYUs/pIvJ+bVte1g06EESzzRBQi2wtAYB6Tu6BdoBSELr
yAirYJBZH+sa1oDeEQA/iHC0tWTlbqTUlHdArGdCV/R/pHRsT9QCCaFvCPs5qUF6
JXXWwcWtvU8qttDTp+imRLWyq2VC/wfGmNZeaeMP81zqRBqMKe5fRPgmMxtloxux
SxYvJtAyszfBRqpskl9t+Bh5LIhLy0q+ZVSruQzO5+VNDfHVHAgQDPtqeR2sP5Y7
w04PWMUtKLVr74/opzegIHtQSbBO6oTtqGO4Ahhu9pYVldm4E9CcWMuUBwXmQEv5
SyuAStWQFkvurGvtuWgFQ7VAc8LpFqhH1DDs77+T6e4UvR6CUJUeeaCRT7u/eFzW
ROoyCZN68PzeIkMy2skRtdbbifKVYD67O+qxKn53CfbWunoMZS0s4Y6fFUr5oiXS
RonNkOVFMpDW/WJmT1HDdQ8KtecJZCH6FexfR+5AzTNeHHUK5ujC9iC7ApeQjQvt
/Z6MmpxxCXZUJyIjgXyAGoELAwAj2UjEUyWjBIT2mzP1GXRz3d+EBL3SmkkhDiWF
m8ax+LioRsfsvgq58f+LtHcms/W8u4ul5BQgWf5QI6h2iDCTLKWgJ5OE2eQJbcvu
1ZucWVpU6MzwcLjYb8DpHJMGYfwe1wAdOfkbJE9c5r0ln+n4oTXmV38QbBByd9PB
wSqLcL5FOpfcYiiMgY1xow+hObI59Bg8NoCVZIZe+IRMWGw18/G83l4TZNJGjqxd
8tBeeFseDYFRWBOEG2yzJX0tduYAeA498noDKzpO5nCja6K+o+SlQIOqzO39TXqf
RFN0a+tx87tMdqr8jwejNpSHE3kRIPaNCoX+YeaMAvMBMEgjG0dCsuXzUSD0D/Pj
wrHcoyaCndly3y30qSmArycAhY0TYqZc8CRpc1X8FFzI3unJkl3toLC5eF1CUW5u
26YCYkDdK6Ds6jNyeAgUVQcCsx+oL3sKnpNxFvjqe36vLn/TXWtlOALMMJDu+BKs
jRLJZHVFNav4wScQuPJDFeM9kgevyhiQuatmMG3Hc6uH5figwZsPZLpNPOz2mXQT
1SmF7QQawhxO3a3plQof/b0dvwjAvG4rsMzF08tv74618/UDNkZQLvqLhRglp4hR
bBW8yyILjwf7M/X+AHkiV9oJzLdIUyLTTHsT7Jr+vAPc3wPFQSUL1DKe1nWKVxxM
M2/ZC3Z/mCzHqVqOVTRqNISGjyp2T5IBqOKjnbQ4j/xzZDpJfV2MF91tW49r1WNg
vH9+41hYqteFBRz/wq3J4Q++LGahDxV96wIo3GCQwmSPeULIbUT5SdQbIKQc9CR3
pYy1SvzkOOjlaXD0p9BwAwlRRq/fH+0KoOs2d6PMEkziB03R1a5xktFUy0khLPUk
3GU2yOwzA3rDpQCFZ2y8RwdlB6v2XCoJNhLP4A1lViBJybvZ3aeKoV/UGk8VOvDP
0fyCQJN4bfuXfDgnzRrZiFmVos00sZ1FtfR308ZEOlUM5wt+AUL7r4wUjEThyxsa
kvgQ9/7gnpUDpN0MPJbY/WI4LxdmAwViJzve3YpRu66YMs4NHiqnaDEx8xtrP/2F
Pa/ielZBP7YoTXOH8IEj+btIeX8mbdsqZ/l9aBcNTxk2yUFGcmHmStS3lE+zE1Gg
RpsjEmtaaS/2n7yu0OyEsrMh840rMhNDLzwvOf0CYSz66LiC/egKniyeH144udwc
ia6rrxDwaBGVxjno1B22KV2mtLfDTAx4mv32kOrL9Ev8/vJ8Tr4O6WPLODSoTqoP
kGiI52OloFKik3uiUiDuEkYQIE7MKY09qnq7uuNCVIiYNVMxPZuPEAW0aEFMJvtF
kC9LE27+C+ZVFiOwfTeArjk3rgggOnRxXq9NCEtCC4Hh5JJ6NSVnuiEVvXGPAoX7
U/a/1ah46wquN8pTnmXSnx0iyUbaB5nN+XluFQ6SdVq2hVROes9JNDHOWFQySKyq
c2yl7tJUVGDyoNp4/wv/dM+MCwJlr1CYzl1C+JIpwMkePag/2xv81ESFEHgULyzi
CKS2XwvMptt0IBH17GnqgKxCG4em/ZI/K/Q8v6bZLKEIPvMvPrnzJh5X7X/mt4cq
BmF5GH8ZCgPueOff4eIVcDrHRe9nOe0lGh+5DLMobPXBazxPEZMHUgB8sMT882Jp
0VEakUIp4et1QtyUfjqBUnDuvGkOUOW3FnI6Gi4/jG5Dj9U6BTjsy8Zz8q7IxCQB
wxW733xnbZlQJ/BYMSBn6N3aurGdWNukEs5sWdtkpHvFfDBJYKP41lE0ibxxhw63
0zBMlrju8gKwWGQ2tedFtQDLtx+JgwTNpUg7+vXxJXU8jMI5cyTCowp4Whbo3RUA
GxukF1MIllBRmeiGJU1lPjsUJo61cFBiT/AnXoVQADeIc+cDP+0VLs6nMmhEcM6P
YmPWkVXnzSRiE1Eh8K26gkZkrpncavuKE4WUMpv0hkSx7UIP/ysNBmzpTYesZG2J
D6VSkCRZOubvaM9kc8kLEEJN9i2F88yLC3le9UmhvkRuRhryx2sd2TgVWKzQWrVO
r/0DwK8Y67F1w3qGpw//PvuiMi2eIsrfgC62aya6GLPYGXEmDFJpJVtR55FiQ20h
FE4NJB73wFniljhuIDk1SBp9SDeF6reZexTC8j9584rPyJ8dJ91HmIr++m7ZENzC
b6xFYQ1KOz3N1CqO+GdBQ62Yf8O1mNkwfMMGkNGzzpIxWEgYSQiy8vPAxri96VJF
q/c7fuB3+0IerHu5/rW8EKlPnDjG+ry8XmBruWEPrWpsJiuOxUF1lnPAS1jQ9/FA
Q/mhA5PVst8yG9qThHXbariasJ4lB3gLD4Iy3Zc20gd/NmxxRr2CT3Hj61hCSeNP
nRPaWM6CzP5jlz916ephVLl9pdkbWi4Fx4UQXDGMkp7ombYRmnlTmR+vZ6nCf7ch
cnoWS3/DaODf98tkgtGOwbLn88Y0h0bEoNd+5SVsFJjtb+22sxANcEbhJKE4YB0Q
jM0ULhvXm0VjK8KOsAIr9ypU8r77QZzsJJ316Ez0X09vro6th2n9rfL7591lN1AF
aS8Yh6IREJIOU74fk4tGgfug90SG+mXnBLNJPmYiWx02mFVi7kot8hvP6w3C7U8g
uQiDLBrZySXG1bP9nBnQSkg3ZMBdzE1yT0oAbYgv+mOF4wWLM2+pE0VpzqtWi1Kx
99pHfmvopbOoTqeYLqXsMB+gJKMFZt2P9nUpnlpR90g9fa8H1iBttm1ZixduuD0o
wST/DRGWCdWcSdfWi8rBj+0JRS3lWHcPSDwY4gOfb9qw6Ac1KDFl3cqI/85KUkqC
qhcIsKTcqqwAMCsWh2sD/+8+XruBt3O4Oc5yV5h0eOYmPxmIHuzVDbdY5Hj8hb6Y
A9SccyiQKqqiTqX8p77vbB6jkjO2KFgrv1sQBAT1coNJ0tEJx/B46FRtr96TEsHI
G283qOYAu/DvRPJFFXW4FWmr9IWebaMtRQfl3YYo873Vf+dyk0g5kjPcbyRUlOXt
tfAB4Ps3HAncJtzjZCDIQ44CXozDCEmzWgtkBDgSmoAD+tLgiLRuej1IhPO8yI/M
PRS5i0HpbNGgIibEVRliz21nwNZZwb0XAkkMY9oK69F2geSL2QQHhIwzL50ZPYxD
CmGuaopxaAIC+ean5yk/UzUjtmmWo7SivUJoSAcviVYyraPcnu2dw+kj3t26w75C
+OWaX+HHfR6Y/0HInlIksgCBhX56eYk2PtQgr4ey8fpkgBf/qpeHNk3kLWDTMVPX
qcw26g42LC0WHABBggL3XbLIFpfsPG/RRkFeh0/5BkpDRW9zoGFbxEfX3J45uiMH
tfSEeSNp3qsR10gRM7OPON0+j3PzoAn6IBkRwfOeYit7EOcYNAoWQNDQWgsbCnSF
08o9yuubKXmHnc9o4Q8big9qSTRvWCZGjvBNFNINmmKTdRvVrcnfjneP/y2a29BY
i5hManCwnybTQyOnGZitRh6HlwierrYQhgKmNg1LSImwrsZaRnkErNBAULVUlel9
bgZcalUDn6WG8zHIG+KrmfmgNMgr1MIyxO3MqN0ooREtKGtZ31iR0skpqeiy8SDo
99IEDn1TVXUNXkP7z3nbDMoGlfkjGxW1Wtv1i8Z/KIL6jfWHIacf7YokU+kWtig9
f18bKkSjR0PzEZQXdCj3doPCJJ3MIJxIaLhauzjQvb9A3bE9RgYIXp3Db3tVfdCg
1KjQY+Giv6RgpYwx17fPwcjQth+EZlXj8WFdLqjLpjLCkVUvmBDNU1qss0uZxx48
VPF5HbOZ4yzqhn9u0VQC+U+IUDa+FcahyRIb00av+sFANLFz/OtVpruJtcS8NiQ/
AwTmtOqT84PDzHG74PQZxx5ggeRoWnKIcDojH4T3CIplLRyTH7ZImK74fttZg1lO
GzrsZ+7CayowU5YK/KLTavO2dWZ/shSWISzA4lU5B5pBZWovNlhh6NrcSHRJU+FD
Lb83Y4KDOMdDjTT4ABwMWYTC28Ad916XU0vZXR3O28rSk2xrH47p82iu56n5H8sc
psCs31KC7wvwEAQB9M6q2ydxJIcvfBFcWPUqz2QQVHB0XooysksNHB7pTDv7Vvik
YNAKok8puCRnQsOXBNl8JqJcVWUoZYCXxExX3qGWzyD1bpnap2dBKZER28HARYR1
6J/vLckM71RJh0h7jj0fwqT6OD1HXIn2ZNPSB+DZpIQSJ/ch7SD/5PL7jwnkfv80
GO2oX1WuZ87Mcz94f+suEh24FV44RGLisKFrnn32CXMvm1XgDWsNlzMBh3pDO/hZ
d1G5PbmJjDTJpjPtGZmpT/1IEkjwcnz2XuomMujT+iWH8sxrdhqoSsi4AZtOy853
xWevI7O8TN/CRm6pD1+89KtwVe9tfgN8ILW8MnSgV7+GK+4FRe4XYjv7xnQlVuAN
lqw3o+p8kJXamsDDdXN2A47vWIV67R5v8oBkcLS07DE50C4i5+M+eaRivkXOrSso
IiIBuxlePrzN4BQZXC6RtQRSXz67Lb5FItkxQ++RxloWRmOiwNBRsJhQQ3oGMBM5
w4SN323DtkGq9r99K6H+VfxvqJtgOBRURV/vzdmEGYeovKez7UmGYeT5tkf4nr5U
WTxTDmHJ16xLKHufLByAEbR/6/PzMa52dz6sSdU6SyfWMqzKSK+kMM6nzUxVCMCU
TgI1RfUSwGDzny5FquAxgbWUU3/A1JAQVyzF2nVMs0VXmUeujzs/APZBPGw8ipBA
tb+gsx0TlT92eTxjIB/4oQM8aZOuWqPE6G0CCU0Xd5g62rRWSyIVZw8HCyqhfXD9
JiS+LbZzxYFeL9kiYnhnrDTOfZ07ubfVONIVRArELnlmFY+si8ijtfqgzJnfo9r/
MJK1gX6w6A4Zk+ktHPEtS/CozS9lLFuwjDLLabij4AYxYCQxGNrZyZrT9suwI5LY
5/op0AO82RKVcPWr62ny1TvnCAhbuLcrueEoPqbdBMlizLdKU4+o8SoxSPBX9sXz
2+lom66Wb2Dg2AvDaj//mWTYqJUcwpSB1zekYCRw+O+bdqbGz0qpOnB3cXlGF5ZK
NIp1JwJxOSB/7pGNqV6SzjOKl8ZOzMQJPJi+GBO5tDmKhCpsbrTstWFl+86Ww0ps
G6PCRHiD2ZYdwTc0Ny2n6ZFPEHgVqq/sy1lkON834erQFHiTcEFxfqWdDHwf+c0+
YhCyeaUyd9HZdDvi96tuPQ4smu95BnOZ0UezDFZd3KgdaeJY+Y7av4TufGKfBPpa
1A8oNENUqt84ObeFgizNuIkGdvFOD4LffBOW6j0mlTbLkjtHuWHcacAP0Yb30fsi
ZW3kKy1tAm8f/QgQs+/jnOkgGmFobFh8i6ZjAUJF3Mq8opUge7lR5Yfy70AGzpwo
tAe8UZwWN7Wxdu92h5YTqOTJ+LoNT0XPkYXgUoA7XYT0yn/fSredeZklnjkotKtf
A13RYf0/BuS3PIma0i5K6EyYg/c18lFM2Go9ACJRBPRuMaEpAW8pg3KnOQpoQmzg
u+A+kaV/NvdrKrNi0/zaHJJUb2nsYLQDyww7Hjvl8AIdEJo2IcpTunvO2zsw3R5P
p2FHcNWzcPOuPkQ//2n1MCC11GScc+qobA5JczIrgyrVKZhmy5q0l+H7w9kUP/zN
XJMibDNFMMT5I9QdrWgFDtNlXyPeCrkEC4yAnitBCXXoD8WuexQk/9wwGWtPxLgC
14SiJd6teRROfFxtqI9KmBuAHzE439ovvz37iltOMn56qAYPAcm82sNN3abHlDby
svn9AaX6ePHz5R8fg0yVR75gkcDt9tinilt10OqfuyfXwcBb1AoPl5DigRxYYw/Q
UXAmB1FO8XBtm1WPZpbNMW3rVmVjMFn8MzSIJLA2Jbe0rbsikJ1cMFE2Xq6WV33s
pbeMv/L782nyM56iEjivNJZ6FCFTQsFSBT+Xt5yuMvjgW1xdoeEtCCVJMOYlmmgV
j0bZH8/bzMwhbUjpc+2hsiHM2kxb/yVwipR9JToiuMk9e7xHOrw7IGU5DEw521Ub
AEKQRUFbUB5PFgFzX07zv7aTDcFs1AztEHEWBoMF8xAZ+cE50nCakas60b5FwWqB
vcGjUNlz5pOJD5Y35SWzGZxPkjblOe6Aq8LEf3j++rmDt76L7PqEpruFg03I/OP2
VPyvUg8PskShWw9TQ4xqwUYIxhm/YW8Ovefz5JiaHbZ+lECXRHK2LcMl9mZocKJ8
CODY98iLCXoCrRrwAXRKnoV5j6rSo/J+jvOKFOpBHOiM0W1sduuMXW2JxxOM7nep
M4PQ6yaE742pt63m0WzBTAkz8rehRC7YcyWFKJwjmHiNFDN5jcWoM39zLHgleKrp
EAvBPqoh0qc0cgECA2DsUGJRPW8onSjFWXU+TAG2ldZUx/IOE9Tnr+a9C+/OW7Sa
NH5fBnbIRUsy3jDUHdWPhkQ85qHAgoyA/pYUEIUL8aTnCcDhTTX+a51SwFrVUZK6
KTEgv69TvjqFu9F1GVSeZ+zZNx9vdKYoC9ZrC51JAJdAEUxCCdadKDfIs1kMUAk9
lnfcRNjODMbQ1dzwz/E1QG7AbnJ1tYvsNfnNHQaZq6hq7nDTeYbhlNLJoAI5Zxi4
IJR1wUl8Grm/OWFOfTj+BKaA6QnVWxhGG3gqwIzhEh48V8AkQXoIdToMyp5KiO/0
Zdn2mUotNrpsIjXw4i2puwWOVzbMdrqXVxYuKvWXfR+OBhLbt3LxS6kii9Z1j/tj
1Gcz+az0v4usHQUBqkHqxQAdQPq/Y2TRoddeywU20B8i2j0l4fO1AdUPWHus2mOy
9wH2DTG19BEpRtKzljLuXdotE0fbLLxo5QHnMTqCVa7u0dykXynpCI5e8dcZr+fR
Nu9N4Dhqx6gsRLkDdnDJ6kPiuDRIXGbHVsd0ckxSrJxjI9BWVUVJqHha0k6H/8g1
B7EN6tSUcJ65PkLcgfDa52QuxKZEDnOm/IDDqS/xapvUCWMIvh1Q6xOMFmaKof0j
3pb/UJ/IfoA4f2rdvNh2H8AdL7Zq5E4YOV+xvqBsXkXWZRB6jIQ+SWIoHDADNUYm
wdlcOyCj+2fas/HlAR8WaujFAmlJ+b7sJO6EnKeDYDYV1Hxa+QWHdFE2pa4CIrpG
hiPjfwcEnWVWmRJsRZioyecunw1tb7KWe7uwGPDL9s4t2wrfFPTmUYVUmWl2LL5X
EVJ8sP1Zn8Wfxs+3mqxi/7We/wAweyWgAaYdUs1+hpus/Va+X/Qehwj5wkLQnf91
a8HGLG6Eyg/T0vs69qqzzW9jqSxWtVaEsnvSfgCWW4Xp2lYi+JvA1/9gNg636Dat
RVAVTlDQbNaxgYnJfpTggoPu/IDMMZnKWVGFKMouvKYmmj3H9kb3JhOfVGBtjMwk
xYfE+htY+cNe9Rh0V+YFNMlDyz1B/38XQ6yKkfptyBxg0yVzJHAb2T94j0Lx3z14
Wy2utBXeW+KJRMjFtGKoUIx2VZgYgH551in6jvmgJauee2cLn91Ojd2L1LuFFgQP
j2/buOhPm6X6miJqslYCclTip6XXEw7rAS3ydUegbbucoMfbmtTH5gSC1TN1DGHz
oKvr4+iA6JCGHI23h4avknsfTSAlzeAUhPMcdYVJbmT4UV72ZX58y/oYUU/6DZp/
p6FoUgiGNhse7Z/Y9yXV2gpkssyWJtJ+TdsxRT6F1R8toFPC+qK9eGcQQiFYIkhn
Sr+9LlEKnxFq8wyiocQXa0UKVPxJjopgZugNsdr8X2/PGQqRRtHT6PIDCHmWJOaZ
ZbKytyCF5UfqiDwaWN3tc8oVV+AMliycGUH61dAcRC2tbCDDfiNsvel767PHA6jF
H5up+WPolhvY4r5D9nEnb416ZZxCSyB6eN0oXKPLlo32dx608WbE1g/KMxfqPB/f
nqpfIjbEuXEI+8TRJnQZb0OWQ2R+xRfWK8Jthi0XxCuVff6KIEZ/ayCH7ejoEJdt
ADy6lkucT0mWFgJsAo3u+oCM+SQqyFmF9YpHSdLOLLA/vjOWbxps9EPCEONDzlz+
eUSqUIYOdEUUSfw8J8lMU+kWbBJpueJl7D7acRlXxtkYE5GrVR19vx2vsfS4QPqN
IlJntaG5p8qIW/uCNENWYzlbYhntwWB5oSphYusXoFbhG6RuNFl2Op5KCejvqnL6
MT7kMBJf5bxu74ZUiidzI1Y1WyMzTUbpSX0j8YTvjqHZSypvLVEumAOjpMW7axBW
GmJ2Cw8wTi6iqw4ZbBVqwYoRM4i0OWXpQx0bFFGZ/9LSxVIYMBYRFNqr9pSfOU64
YwDjP8CEO4JnlVYlmj84amu3/Yr3aUjebasj2Ctf7CiYKEKMV8XhnZEuaS58vOsB
sNE1d1tN9pB9seKMLghGg3Jia+EYGDidUhoqsIY0Lsx++lKmIIT18PTYLqamPk/l
piBoHZmEAcdlpEdwALVJscG9fK9PUAssX70Gs9jyYP75I3jmx4d34Qk3wjQcAdDQ
42R3uj6uYmlXYnPQmLKycs0ZY5ljGVhcTxUvVek4MBM8Xn9SCvM4mC7d2LtJWl+Q
/u28s1SVBosnksn2gf3b5GUzlwz3FPqBbJZmUy8ssD7P/XVX52jLtlvl30zirAGy
4I9Hk+ILnUq+c1FdUlSDmTQ5q7mKT1zNmjDdRuxqd3meslSAnPEHUJ2BENCEUHjG
Jl2CkNlchQ6PoK6pkVyg8Smv7VG1xC6zpgbOJmBDo9JKihmv1wqeQQKU5KzVP7RC
GrkLkt38YaoLm5lIKV7eZUv0AS6xPZpj1MzT3feNvfqS+oKr8RylGNkgpS7kvdNa
UOr0kn17EI6dqNhufDDanz5Hl3OzbRmn9djnkWOynUSoeF2ve16+cOKQ0JnPUHBt
sHMuM9aEyi0m3TeW9G2AytK/cJ+GAQa/043XPQAn/aVHOQbIziZKJIy9Qyr6HKbZ
a/Q3VQ/Z4EHApVZHQiw9936kN5O6BW6MTyEkGQFE3qjU76Rz1JoOLcqq0oDAXUUz
3eb/kdWQTphrUFWmIXSRomp9Zrdd4eu82hNY9IDDrCJuuTbFcMj04xRfCe6Ugf1i
AsVZ1hZZxXOYD8b6OtuBfWSYay4w1JOt5qU4+Ut0lm3pGmutyFsJ9e9wqEk7p4Fa
1R66jG+naIUx2S4VkWAi1aBrsXsg1Qkj1HPvcGyrE8b6sW300byGvK3yqK32xGJE
K2Q+lhgj7QEzOPQTRD21Sv8MIKK0G5kfJxfIIifkwEI7qvbdLmmgl6VFtUDpNlSf
KEUjUNsTmvtLSS/6+bkzIhIZCc+h4pWb5ZOA7XBA4r9zOLtxAN7CfqN4ekP9aP42
Ovr8ANSj/QqqVxbIuJun5gaCs8jZHRKkrpiEhrA223wr3wtNdqkTDiQH2grQQoV7
YGDW0GBeIXI32Gm2HIsEN6FigHBpwrirlwmLW3zL3Ovsz+x6H4SknYF31BLLLmv1
AB1MA3lYcBgNeM26Y/NFd//f1lcV/hnsb/7JBeAlYHeL6nXvLhdrufwTvrgL5Rov
nllCtCUuDWhQJqrOhCufTBCT1wnVee4ok+zKyI+SxsMXYg7QnRWPtVs3394W2PIL
1lKxMye1+71zQMkaCum4RQ5DVJ/YCTNZaHpVWuoCpU7vP2bqQKfpV9UXsfAOyNPO
LBmPhmT3IWYVI9Zo2JrbbGAZIIKUoO1xDEYpVIwq1SC9VCXfMOuEcWO8qT6CNGMx
FrzghYj1VWkx246pblDdCYZold/7RMybW2TTSNqmFd4ygnTY8tRNhFoR+wT1xg5z
9v+tTV27qIx2Sl+Kj4XfW0pDfnNLAEYDkdxpH/hep3iUi73ewMzf4+x5q3nIUnwT
Ih3iuHA7ldOEj5e5/8EH08WlrSEXUI40ugjcRQBKVIPT4mkS8x87rATcmIJ/dVuq
HcGf+eF86cCV3Ud+CLfDa5Y8SMBx9lynIHdvqt8vhao9RpTVg8n5cCoUkr5xcL9S
+SgBVVt/y1ZSEIy62cfT4wS8TpFYeg9Qi0tA3JAFrHz0JdoCDKYWcsdGvyAZIhuP
ZwP+Vz3yQk4DVwZ4Sh+rGcOP3obkPWGDgRauQ0Cb/M4oyhE6OlLKw7+bK4V8wBla
E24kzUU+EbSySz0Ow3jHfWOeQvgAhF0nVb3fXk5c0S7rBSm0+4IkLz38WnCCm4Fv
m0S63mAiKS6W6UrQ/5BG/2CmEiq0OIoUkM0YaTeVOVeyg0wA58Ovf2YfqrKNXdiP
ozmBkg+WLBQc8dhUxaytqjrcXGmiLFZbML3fwX2bgdQV4/IN66TzFqfJ5NpRb8mw
EDPxmy8PasTCewgzZ/nL6d1MELwdL8Pv1yv6MzOWP6AqVOmabqDw3MgXpF4vE2TR
F3/gV6YHaz++rzTrkvx4cyNnHA1S7/LJhkKQFc7c7xklcdtZ5EfNXbJzETZwJ7m/
EsNJa9fPoPfnekMuye0g710enp5jq8+DhH9pQN3F5GQ3fnZLdE04YrM78+Tfrp50
pod0o6kpYfgpecjEM0fIaIS2PwTcFEFz3oeZ5aDqpNqdpF2WIDTMWKJNtbmEYBld
pnGLhHPcvNIyTp6W6X7VbE2uDFgWBP9+bbJ8azX7fShaR9LIik4Kqq6IUaznLT0j
b7cTTH9jZzO00yfEfIpHEUPB1KRbG2CaeHJTQJjO4tIOqmdVpEaUaFiDF1BaJZJD
mYGmUvR46Jj75EFt+G5yElvApWzAjDPJIZ8y08SyFuVOFn1guyD4wyNP41+AHrlZ
hBhObEnmnBLjCD+Eagv+2b1fnPKUrm2+bnYh8m4aAF/2CZ2+I2SbDP1CLzVeNfSP
7ZwbgQVzt/S0g7673wmRBmTQt2BUjjUT9sOYA8Cx7RfJqReHdU4R5KvPw10/hJrg
5ia2hf0o7NDJVp2wced+I+GJusVG0VJM9FWwDwcSwoMPbO13MgmFwhN68XE9rWp6
vc507cbaKqMcXgpaLBWPSNoxH8Eo6FeSulUh9Q8VTpSRP4raLPzbBzzbZKe89B73
oUzcZ7n/0zvXmcZmo4nzluOLx0q8ocyxMhjoC0Z3MO4+MyLWvcnV+oYvkE6PbT6h
oAfuJ83xVEVYh284WedxyoHN6tyLIC3Lns528WuW2Aw9YdHRuwILdog4qiE7wh2/
9VVU5iVDWNxXvX/3jT4I2hImh46IS3Rgi5/RzAh0VmwTgl7lyrvFbfCEcQFq63LT
/f9ap1TELWy9kRtHletTE9AgnZrcOkOx3a0Ba9C9dkVXn/F1sEbIW4tjbWDlWxhO
cBj/QStWcKd4VrCABvQMpgDekpns9vFtJ1RbyXZQzlGms0mDOCOgIXoYlSAl3xke
JSdZxAD8Nts9Z0XYp7bBvU5jglGi2TFw5KoSdfkj2g+2gbaBImOAe8zAEIuV3uzu
/MtxyPlqqWDh0sm2v5Yhlsx0IRZFHrCd8u6MRYRpZ+SdeyhYiUt5DlFZj+Zv4fwd
2M+I1LJvsn3NMHAKt4VVlXzVRjEkkwdTHZ7Bs4R1GZXZ9zYJa0F3I+sxlayu+ZvS
aO+jULsj4X64VsHOjp4dscNq/YC1w+tRA32Y7b0sMPFLBBaI0IrmUJQC5jiwMayx
POxjAVYj60QhhLpXU4kPmzq7yhzSNEeo+ZJEAVPg8wnVEdk1O9boC2b2ra2kNwoj
0+A+BDZFmAgBdB9E6q/0oBLsuG7Q0SlnRN+rRd0n1pwotCe3uvTe3hXWDSf5WVBS
H29H16PyXFy+YVncJaDG5cD2utdrjA/dng5YjpL7Uk94aLMCzMT0E6V4pWZUyVMI
GK+j1k6DSQ3Uxijh+s4AuIzIE8dsCYHDpsKcF3sA0u1IrjG7qFPrfybM6alEsv7a
ha4hHWenLe436cUAnfOQocC+Qnfu4tpei2NIo7kKyZrLHy9CYpGxfS5jo491LJUs
bpZMtHyN/lRgDoKO45JVsJLxlbArsoXlzZI7PdYVRuRlhuTEEzX4ouse4Li+8L91
mvLB/xGupAenmavxMw/t/VXUITVitgoI2wovZE0CFJfBn7dod3NrqKH64U6MqfYL
TmXL1Dw7nAWm+VIsmttESROgkivAICw9btw7kC4wuVzRUWE24od6cS72NAAujxVL
1BIxi7jV+MNv0Q+LkdX8TTKfHa/iYKY2V/OPx4JlmzdbUr9lbMhmkJZSRh/IuSem
KXa8kBPg+0jwB2YXwaNQfak15TD4UbyR7B2cxa0ZsO3dUrn939Dq/Fa9411VncT4
PSEJOBD7qePrT0oq0fXoD2xTTiSIk4n+75WvLbLFggNtzLUwaiJA797jQS6+3cjD
Rctb6KhnxvzPZ4Y/KVvuWjHoM5lTDsHg84uorM3LRTxtYX5qz1SvO83tIBKdi2ac
07IdBad8JCYGt7Jdw+dql0K3WVsv4iG02vF8SpTNxuasziJIWZW9OlK0jJG3Ep1V
iJwSHpha7UkOoR68qPJb/vpvEarDQu8ft9g2IxDfl0KrCHsFts+5HvtxQnwg/5Sx
6BlZKHfnk4UfLIkwpNz0LA1Lv4twiE2voQKzKJc3su6Y4A2MUsYJUJuHCzeiTSZj
vHJYp/cpFPix/XhHP/kmYSZrFGwn8A4T8f8SFSd9F+owu7skzJkCYN0Y0Gselo6G
47F4vNDjy0HWpAOP6WLFPwGtgApv585SSSG8J/+Mgt3zUM67YO7kKn2b9fCW/6fq
4rwV+oEuD7TF6/4qAl4qiIqax9ieSU7vEeLx6USIm4ZtIof4p4vRiff1HP8KGyPr
lbm8Wucw3+gf88dsenAraOVy6XY+f3DtKTHiL8iDRCofJb5hhhLIovstkfMiSyrl
iAZiqSwEGjDGo6xBxd3374/c4/zVhlVTEtCQC9fLlQ9kAhvoHn6BhgxQuDKbG4Vu
kzRq+BF+TEmyT/gUNe5Okvi7ABaRDzr8uI4v8qbEtbYT8zwWXUs/sYLPZrWKbOpT
GbAkwuSCxhRQxIj+UL/RWTF5b51jZ2l/CXT3Ov4SyBOa4IUm83bVjdpYY503G7RR
M0QLWZdBIOYJYPwwPC0XH7jksnG6Pccp4rcaoYrSnv22T5vd2jLQFNWmEpF0ie9F
70ZA2vcxY9439wlW+LUxdLfBfIRqvxXbciJwlfdfy/+7bhmKbS+VpntcLwwq7JnH
IfBFPn3oDk6Z/2r3qHs+MeJNwv9JQ9fBD2zDY2oX7ojXz7HNAshKIkRAG7H0UN71
f4b2KA05Hv5p5cg5fhxt4WQCpwQqwLajNRxXQqQUvJEPJPm1+I3ax0YrFJ48Vz8j
guiAnVeXE0O+nPB0W7QxbyWUVqVfsXl7PpiZEK1CTAt6M4yiu/CTd7/giVCp+enx
iUHPct6DzhH4CV7c+KPUERlDYFJ2yv1docpMfe3jxHVKC95eioNPEK6FaP5jkDwj
IrPxOFGw/INS9KgfxowT3vvAQtR2b5n2FggD3y/zuiaAstckMppUxHT8L+VJE6Vy
Y+zQglirdS5gHX5KPqlFqHeCeg43inak8tzVIBUbD3durDherynS+DkFiVAx8jxo
mFaDBgik1NEbXBwrUCoDu1cvWLwAjfku82wTq2G1Qn/ip9OWUqDbHENmWQtMX4Qm
mpRIGkvwGi3m/AA8hzu8g+gzrfhbVLSzbdswtPoVCnSyRW1qM96x8EuJkmlJHOJX
D/dMSqaz9j9RqtUMjDOdOOXwy1XOb6N1Rg1qX4IQwlbos/wcLlKAxKRhivAmmceD
oZ+zbvI3Pb9N9lnIqP0bInFTrbc0sN8IWB4BnnLRanKcyxnrd7pnKYRJSS+Poq/Z
RF6N/wJ639sTN9xCPcB6osgczCVPNdvgRThcRloRFtDJJVFA0rdDpIj9Uq71YLNs
IO9wGEpvnixlDC0MXmPDgEovSsvJuyNFKULCuwVsvzKcD/KUT5MuxAcLbHfpS5we
BwPfdFzJzWpIK9cY6kb6FMHankce3wyV8Vtd3iuZPw3OUgBzyPcHv4JToqEYTEgL
i+Kw01JzbqgQk5emjPa6WdVpUTdfSlQt0RYBaiOCVcNO6GAFwqHJw9SShjOXwzEa
TW0SpApromMeDcj7UQEkxIu7iCyAmLqdwPuGUXc9V2/+WAg4Dz3vzojIk6ESfAFD
re03V5osUs7d/S8Pv6PyA+L5tFqaO1Mn+IJ2KGUD55iW1a2E1QFwfeE15yqMIjgj
kkBfmGo7p1UtItGTB5VzfGYz2/XTc9sewM5ElgBweP32Nj32N5CXVOVsFJwHCwqh
L4pMMD/xiO/vA0tuQ4qquJ3eHXJpVhswqslFwKH02x1HNrbzAIDtz6Vd0PUxGTV1
xu2WwPM4leXTI+xnLm27cR7sj/WHb8GiwgywiIj93le+Kp47lpCuvdSgQV3n0BDv
HRMQR7gWUJdh7ascvgzAyXKLbdYj6XJYHjVswoRbLNZfvMcAbP3FUUQZR1sJYMRK
dUwzMUyByu2wOY2WeRlSe1Xb5lLHgQDFkqbiq6ZSu7FnejYZCxAcEFxsuGaCTEwI
5nlQVEjXRMMEgBkFHFJlks15+L5GZYNyfj+4rQ0HopBuhIsI+wD7m3/y/HGX5ssB
V10TTlAaCWtw/+de1dvrXMgNGWnKTM9xiRZFpKKg6GvcMm2q56V2Kn1fRA479pNe
AgAGiGmoslRzUyYHGBd0uaabGs+raO1cwmewZIPq2zJWtXrIVDo3gKtXW+wAmxzZ
1nAT/S49UspE10rtzZ16JKF5nVc9E2nW2twEQJ3rsqg4WEk7+3ypUT3xnCeuVY/x
jGswRoq4l556kMVL1FjrQ8pKKOlNdM32hpsQZOsE2hff8UudEZOyuxrnfkgYrIrf
dJiUWjhsgJZL7EWjGnWZqoaXhVhj51YL1YTCFLuyfeRm1LzD8aXPudF2DsB0Q0v9
GC+PKnGPd36KG4gh0TCoDBdXKEbQ0DQklOCKrRwMYJcR8e7n0j+Hyb6cjuFsgwSF
PmQIGCVy8OyngZ5i8GE1U8twa7bah7bzqIlAZ7SXJXyEzRSrawCWcM8mHZ3gyplI
PM/MNWcHblTlQ6cPztpmIfxSo5XDxm+OIegaXlVxz+oNBmgOvlBW1Dsj5YyfUwc+
H3z959G3ZWgUlaNOJrSZgWh3Wonly3RTqGysN5Q2qAnxEkVYS48eaZ4W49R33Gch
LZhEluXJsGs8YWL/BcoCRO0pZpbzkZCwWgqi4GbBpAK6VKpnqysG7a1DZKQjox2I
weeCNpr52keQY2STGLsSJnPIrZMJG06vFUDCw0eyhYfX3jrG1v7j1r/kFDRUvdxJ
nmHAtfYRPQPQ7TCd0aTLXLDHE1YNwMubG3YW7nK2rDsceuJNUCHuchQZzs3yM1XI
npIYE+1mSwoC9rTpebrQhI7tRyO/P6Ns6xSEkjMNf+VErMVu6K29S44IEfWalF1W
16tExMC1y5E0lVZ8xd7CV1JLJw6/oPx44DCPJ0OnD7B0V7MbwQ6mHwBgvq3oapi7
7NKnxgnQEYZuOp0Pp7Tt3bYyHyuX/Es9QxoojJqUVs8hytRlUa1IbFOjGNE/BE46
6x7UDM/bEYG6zmQ3SU8gDfp+tPI2HvwTzQj7rxLyO4+8+KhypbkHDgq1awGOkylY
d5pW9tgbCy+joTLY2M6hxnboaigIbQGpROO+0eo5ssEMQdUYMqQ2Y0HIv/TW+CBW
UwGbOdPTU97EHMz5P+eQuaVuxvDvrWjp8YXfXT4WqaXcz2an21vTl1p7oCXn/ldu
NxlDHpsApHls6+gONrhqlkibIz1h65yxZDvTwdAVP0gLmbfhknWGysKTaWSQQfnr
MVCC/QL6XYHU2wdPlq0a3MDoMlR01xYn6hvr/1gf3kYWSXk1Lb8u2owTY83fHeQc
DE0uLx2adQbqusl2OueWudc2I+a9ZaqVUi4OGdcaXN7btzKqrUGvIglNxtD/KvTV
zZCaAcCGiUsZb7NGYO/ouhb2lFfhF8D+rZ1/zMIVmFpg6VJSP1vh/YZeNrtbqMOJ
S8SHsa7vSLTDmhX7ACrmd5H6Ww9mED1h7FSMwNtekMbSfquNedSGfAHmWZqg8Aol
4qQalWyiOd770r5EgxqVFv5PstR989D3lnYTTRhm5KAYdfqMzFLD9qMpgQwTCPBb
qlViAn+Tr+UxarmXA0MiF5nszSjJ+2TotCKMZ3uVRIckoPzClemexRjxsoPJ/gmQ
S9pDer6EXbi+c8BSAIVkb+1LIWtpigPQlcs414oNeMIGiwPmgHxfkYV2PNp5m1Ko
46QYpXjgCSnNr3nE6c0e8pG56wi8xBho0e9IG4noNZXPaomOgji1ZbyVmmfTvhvN
wfNZ43QV7hm/ezquCkTZR++RnVl+zJWZgJ6cKaJThZ04n2kEQAo88xLtmoOY9kHF
1hQ4DyP+5fiYLdu4Abqp1x3ujuJnok4yIAAVKMv4blU7dwZoN31TQAXarMVihCG9
whnXOqGcalbEeWWD7znKN3zcNFmoCxSUUQbbwx+T/mvJKmdxUhDuW7smX3JZpn7c
JCfUvzHoBRnqHeSgzyZ/y9PTzxSQ5767PhStku3rPzdisF8Zeu7GN64z6Udea1mm
Nt5NtRO7nVTyU/EXypHZ+GNe8Np43q0pzhE81+cwgG/cbTbEH5y/Xw74AHYxUkud
ediTHQEyTzjsL+dUKmFWyxTbugQXJyVUpjscNtUeQaghcZvrtFYWOsOw+flLAfHt
KaKhj3Nrv9OzNs8nUexVG/tVG0sTk96QGRdoIIUpHE838wJvpSFcxktRANJo7KF0
zwsQecvxdIDhKqN0ZI78hj76rI9bLkUWE7MFQpO1gpnb2Lx+Lb760klg4ud9M+O0
vvRJI9bPQLdCIg9/xWB54ySOEC3mG8+vWbSXavyihy0eCcv/JiB3eafHKIXpf/mf
O2/xR+B7079KfJi/+cktryRxd8OBNBJh/ATnGfNGBvKdcPvCa4emVhx4i/VFKhbW
iZLVuVlwS0ebepMeDbPmOkt4srU1uYDUAhvgZC6/XIEXxJhyg0tY5BSGI2n/Lz+6
n9E7/3ASgENxYUom9q4oZ54m6cRhKsO5BNj2EZI4NTmITKy7wfU2hHVdwP+7w5bU
cfJ3n3c6oIQFaIPyRcc4Y232pLbecWfxbAYGl1ktH48kYaioYtUw3iV0QV4ZBvYi
rj4tPPT4JshCYicPKqv+prymgCXXv/BG/NmJnSj5pDSfC/t/0dPtSD5Kce2+OwTr
vz6leaF3VG9bA1K6xVJMEx9M9UGcphRQNNKXCi308Fn1vYPUUJ6xG/eNAxzsnvpH
cKa/PCR1+VAHumAlmXupSq74ymgsYb/LKuu0XamGmZJCN5jCMQdpoRSP0UyKa84O
4/MfJwu6jgzMa6eRnbtg+oQEWHNC8Ok0Z407oxw4+E5vvRtMc/RgVcuPIjeUz9Kd
zpM7d0NrqNrk+IcZ2Uj8eVqwJExGZUL3CZ3TW3UTREvPHqZUfPeN/zsQ0TXzTtgu
NbcJMRLltUW8YUFaKTcOz5xg2Hban3MqnMSnhp/j7/38H2DVZE25aXiSX1HevGe2
2vJVNvlRITb0RQtkuQRMb03lELwc7Pp48Gv4sYEtuJpepTHn4riQlc7TCBE/9hww
7ELcBOkb4xD2RHj092fSP4v6XQ8OBpfhFCZG34j2y/CgU39wdJAMmB9ItrFI4/a6
BjP8k6i3EoRUG+2olwHmgwnDOXjPX1q9rslLfbpWpMubP1gBS33hlggfmiAqfwT6
PkNsx4JZDmLPw7SCsODHrMXBj82Fj5ynrr9/at/ogWaRQLH0qC2ljrrtDsqp+eXZ
D/Cw/bPj10PQ57SkqlgXXRv9Drm0TPFpi73GkzFePfAu6PhBexvTRJ+ZfFqE50kj
OGzEt+IJSS/MU+Go4W3I7rGs34jEqGXS/wQF9lWdNsujFxkqndUk0rBu9Bd3/eab
uymOnTLtszHIF56lVjPoYpVhJWbmj4j68gwPnYAIh5Qr547igu0MQsUCIlLVaQm/
4JfUeY4U9cnQ1CcUOpJP5OBxQPefsbMFCKWNH5RnBlWIKBvwf3fDM2rRPtuI0WYW
V30zx/+Kk3yLEouIU+tGjwLgVf4LUcyao8qf1zXxxCytTkxHmfhoapqK8EwbEI1E
+kjTcVpqCA1S4dx6RRRwFydc6KSwOnny2BBUo9XRd0ZZ70EMlxOyGLoWEpvgoiUW
RE+PFIC1YYrcAJ0c97Y11V3w5OZ2w0IZxqWG629aORnzpMdN3lpeA/gboSbh4Rk9
TDaxNwarMFKS80D583cu4egFZhXx6C+r7HUzeHPJ9y+/yTk/NnMu6sLi+HgIWVTC
LX0sZ5xUF0g83pT5WDBOl87LrNv680Y0rUoPsykOyhcD5XXF8DyAR7G5gpC7iPrT
gcKtYiYbixpcTNK2MikI7+SiJ1Rwn/cQZK5o8T/HxAjFnX4rW1ItuI7BX6cawxbu
uRrwExoQH7v/aWGu8N1+NciZi6UbJWX/XUr8UWFSsL54hwKaa+Kyh2lQoPdzkLDf
Sj6v4eXWEKgMr31nrX9/ZgOH4tP4p5ll4/VCwwe7Wj0NuGKm23mlLnCX3XGdQY2w
pAg2BO8O5RbxU6JHfqCZGGsCXOnB284l3STyh/7wlfeXI1pWfR6UI+M5l9nan99+
kw/jSTd/acfXr5Ybv/wXMLhi62KdM/jV7B6lFIsU4+zYI/WvYMBKWhvGKoLtC5rd
o/Tl9UagWvh6fM091lxMzQq3CvpmCHXu9hfnWxR8Z3kwf9u3PpUuGTz/Ac0om3tL
oYGv9Ph05gwTZJ9ieAI/FVUgyC4ZVfFaDzl5+NeIQ94f1lrFEoklG2C5xyw6U3RF
MpEe1Kq3M0cRKf7EFHY8ani2lBN4jqSf05YjMBnIgN+EWQAv18CIIlBnVJ5P3TaN
6+yKxURjjZH0todPf9wiAegCSR7LrGychZFsy2AV8ilsy0aDa1vD83o9Nd1FH05I
TztK2dr/laZkRnJ4SXdy4PrByDLv8Xx+kTdUsHQYHUWSGq/m6K/HVQpjkOyquU5D
EKpmvE65huzCDvCBzRk6J1gcF7fpJHg5svY+DQyuAI4u8glxFK8LjTvF/Q8NBy0u
webxxKnjkDzQT+jV7Q/3s7IVYf1aNqBpcayGZhcERcg53XmifZpjVBSszbQLHtC8
4TIZlMb8D8ZwkC68zn+BDt31mGMtZCNFCD1mgxiVTa4JsZY9M2P/1Kgg0ZfqGBdW
ilQfXnot8eBvyHV+MKk1cx4OqS/vr9ZDpLwNrNxrSpYDmeJKYWcUwb9UX5ZeZ4Kg
H+GU2BenIIE9vQaoZZajlI+vWZlAD0DIC6C0lgti/2vgkTtdeEykFBPnA1YpWTn2
o69EEZCYpcR61GzPZi0S40uxVrmCWSf2pvXIbcWsrVpd7/TFvS5bwfuS3Ny2W4EE
aB9ituob6Ws585gPm1jhqYOIBzXCn4k3tNnRUqiD15hUytDIvLJbbAs1knXZo2nP
kUyYXp0J/yn9O3pxZSAKWdsVEf9KkBwQauF/g0NYwRvY5HnYP0q/BSZe4qebzeg8
l43JMRDA/eME+6LO0J+7a7/XBydHFWGqS2S3cz2LUV36l58qIHIf57pg3Q75KRCQ
JbVqq27LD2YevCkhA+GiF+b6hmVC/fqdN8EC5lrPhS5HtOhN9ejRpC/jteh1MEW+
76EA94iUX6sKwbkRPF7l5qDYO2ebHu7CwgGuhZj4aEhwwQTZW2q6erR43/fIs8On
iu4XHyrbYXfLinLaHGxRQH0CUQPUPcd53jfN3yURpQLZhzSXrcOFNoMF8jmKvNgh
U2WxIekAat1g4XJ/bO1w/CLSLBrqHkHWaAAxQ1AlDwXy7tB7eqmXwZ/020xCLtdn
m+Ba/LGCNNxcbmEhRY3Toq346C0f8pzlgLQW99Y11oW/AeZ/8+gvEXHIRKrGM6Er
JYVaSofEb8WWdYrRq9cZvNL4d5GqvEVuyoySJVrWqxj2H7PNZ5N4qqm6e5Ji42DE
23eeEcJWNvzeoka9NXJ3Fb07xCB47U55iZEqwMKRiMAkDlCBS7MV8L39tBcV3z2I
IAQafLumeFX79l01DZM0JylabORJPpcp9XLidPsmbNj6CbsFUumMwO1Zt9MOQrzP
BC5W/We218hp80M8OT3xPZPZdwv0/uZcqtCjSFvgGFTQUjxhPUy00vZcBupQbKfq
3BVpnpencN55mzwwX1bDUb2GVIwnpk9fj7f3p8gZnzV3Fpl3GYG4Al0jYe1PqoJa
n6sSZd2aMH8X+pdFTL28yrqSfFcduH5269+U2N6lQncDc3D1/Vqk6ximD4t+nuNL
i8ok4uNRWnF+1Vw4GYj0ItxXNHWImai7pEogRIpqrChc4MUyGmFone7lP/Hx8I5Z
PHYgXqJYZIlsrHGgPAMk6U+cyPWY8+9PVOBDQUoy9r4Ga5p43shH7A1fwGgK3MdT
E1axSMDDTcnTBOOUCPdOawT/xAht7KkDLnomezkZvKlYB7mzKDM4UmB250p4PfM6
SUQuC4LcW+df3d9lAGd1hmuJqZ5BxKt4SjnWpl/At3JMJOjcsj6ky0GKnyIv+hlb
FP2Hz2S1ovqeKudIYl01C44jIeab/kr0DIEu2JW7CK5clSFv5wapXlSkbHXtes7N
5/1e8V+0pqg6XXHDdy2NldlaO8RWrO+j7IgOARiRloYfl6nvZUfTVDhoLbWZ9mbC
pZLoENbKSOrB2Pdsh9FTVws2Sl1ruKtnUbb94YRlvw08wdsxAaxi6xDGYbSlfeVR
cSJ7PobF13wka373yJZ3yHsVa5F4SuM/qn/URQpT2aaFiKHuftlijYxHXPoCc/i1
iodnJzoPU9q0QACeLe8elorHyNzHk4pBrEp8lPbAo1/2TtV14eVcpzqzhsC7wMO8
1BCH6tQl5zZW69tCalLBksXn0Ob00yqy5A+Oc1sU0EdtaWV7IyDkgrZcphJx1ais
ej2sLRhjsTEDAOopwetK0kKNhfkKxb6uiFrkPkgvk764l9ZjTGHksgjxCv/aj/qt
fwyyWW07vrYfyAMg/FNt3WuBdWmMG3Q1yXRUkNpse1FwVvVrERZDBPkBEFcI9xSI
F7KI7/ADhYYbpPYHb0woaPs8F8T+qNh1DYXxzQHBcSXamwBoC54QpmPsuD3jeOz5
IDw8kITYlTAU1HxC9GQIC+ffBFRZeCWIKtsyGGq/LS6a10pIaRcA7t5doRUduLkH
AWXfYPSNuOxgky5zUOgx9oBrE24302KiwUHdzNk4EkhaUUJHCFuPxNEeOIcaBlmX
KsX50WOraiqJa8fuczCFQTNfOmxF1vEbWgrKJQ2pkmx+YXyx/WpvCShcOMQ8dBo/
5904rha+nF2dmqwv7+TYBna9M+U6Se+vhyj36cRbwY8FX9DRmg14VG6CSu4Ku7fE
Dbqk103B4AmDOuyYC/a+nRMXGvYyzCQhVopGPHSpjc78j4CjKduGgqlxyvMy7cPj
ZD9kHZm1GP5TiMZ+k4ttH2JeGFW2sWdHqWixRwd+E1c5wKfFwvwyI5QSE8QWrIea
VE9WLvdDzrJavpR3dxttBL3uwzxm1v9xXlqn07DjP9/rQmEF3TQE+NLd+iefaMg+
bPcPqiT0JpMCdGphMDysBXtviqmQNvWa+EFnCbuikqw2Ng3chz8QI/gOq11qHlqE
XgoNC2Fizu5FmyLsCGQn8UJyVqGN6NBp/topz7H+RnJ2txuXXQEILE5nCvvfOo9c
xycgNBF2vsYYeKkmFzNfyonKAdm66zah9AJJqZoiQHa50eKp408RTCIL00ZMTsB7
1fsuj520kXAbh+x7z4hV1fCiIeXp0mxTdV4H/Vg0s8GDZ95sXj5DYnNTupzvCjq6
e5mXOwnXni0sIp+n+SH+3zINhSmya9/Lbl0pgaOUKv9lZeSyqIEVs45dQ9mY7zm3
5NpXSLRnMHBLAINBqpm8Hg+9z+zkeDMnKLz8aVQfUITz86t7ikbBXNgpyU9RKgF/
IFUIIhbyhPS1qcaAWo1zcbJDTqc6g2nCcB2+XEqLHUtbCeITWjpz9iif7yl6CIKV
s9ucRypnGe0WnNYz0ldyJ7TJOMMLuWH4l5HOPom77sWvWh8LYkAEOb2sESBOnoyo
UkgfSZ2HF5aC4ahyzMPqyUzMrnXLvwUXg8H2ycENpKV/gGbpuyYgFaxuxKnJRKrv
O3cJRqlrqPYUd3saZqRCgT8fcsmm/AkPG+PniF4i863OseVS0Y7IgqBC+GpzCE3P
9I/5PT3UEhvx1yii673AnKXMCkSQYkNWY0yWkliZqx+dSucJuCGNWq3wXaCDhcDe
8u9SzlGODf5aAiS+AZZjcM5Iq/ozNYUgmHNrnGXMdd+f6uH+gZO+dOjtLMWN5Lvv
c0VSAT8lSz/zO6W1gwD7f+3qOGCiX9IjMjkhsm/FZQrK0neuqsdyK/FK6hTM3Ogb
IGsFPsb8dbNNlM+XuVIFKHmLnbHlgYlcJbVNNGkslrbIPpXv9D5226KoeXyGkMTr
0/0NfdUM29aoLsrj0n/82ENZcHn+FBgEwBNPTF0KnBzEs+M7xB4DASB+4Dd8C0yk
w/bHCsR3jIkBz/Pq+Y1KstGIyu2LJcnYSqApxSA3ql4XuyVP/vtuCH4roOvI+kj6
hpbVoz3ZjzAhal1zi/Ciu5xrUqj7DLGthlHMl8JgzpEePPPjolXElUMhURL5YrzD
4yC8EKpZW+4OSEOY/cpRHzlaFHknbCbPhsQkJm8Kr0tCs66hQHhow+4buNtYlHLS
JTZgRbjkEbRUWVJwWOWEykUa9oWz8N/lr9p36MecEWF9i9ZlKbpTaEV+4SpX1WY5
kGu58gwFQQYyiUL7DvGp2zd/LRMUP2tGyv6q6RGPgO7R2MiKy0kw0niLhYlmc2Mc
fuK9nmbXC3nR4crSxUDQrYscyUHtNZyK0RAYGS1VkTZkhQ/HEHiE/gaTJ3bWJXyG
++PplQFCwAwtvsjAuO1ot6z5rQb+Q9Vl75xtDEJMZg7y9+9yjgIt/MeNRNs92dGX
N+HOJX8P01q9/qXV5RRT50nHFlT/IVvYXB+9PgN3Lv1HChEiysiW8V1E4QVBSdYm
mfeCzk206ZUUdSQBp7BgXe/1GpPUMItmIPhi/kLAqZSulhHfBHwuUUYZe0IoXzzq
wMufEIrl4hEAXfSHSTu5IQ+l6IDKJf+uN4+f4369GGnc3XnReGMuwsKMEdlt858y
quJzsC4A8621V9EXgr2+nZc1f0r1KljB377Jg6BjjOhhxLWlmnHUNKfZjrfvO4Rh
3cTaL8Fp5dcXQieiQGr6+K934nN00LplpsamjsRHjbh2cMnb4ShJoj+P4KFwlAeE
EKGVEEAGqHoMpAIQGapKu6zZDY1HAbfvk2UzyxcvDsKmnKNBXRFxHXi11fuQ5pEK
UXGsTw9BOIPOXq5UP62suudw8AH/TssZTgHzKK/FUhvXyGa/ZVljLTyt4JjojRMG
QOLsifzdvCAECeE7KwzwVRy7mrNEzk6WDbGtf/mxi1+IRGLHNQnU01Fkne1MaMca
o3i9yx/cavKpXQIRp3A8FoMnhCj/utxZdY8R4XMa4ZQ7MEMOl0RRRcoNVgi/0xdo
B6aUkEclldPw6SvnL7uUyqU7YjoII0kcbtuosZmJn8Sm++HpeVpdvAkQK2UmmN9w
w/P3mdv2ZfgmVihhu9a/68rl1bj5xop027CLZi7wKzVb8P4I38t2zxRyHgku7GNI
lO3WuFx8TBcU+dgVJqxUq5K8vb4mfSsHiQNpRy32SFSSQv0xsFuDdEWgoJxJKkR2
BJHaEsly3O5WoWCiLKkekoXoJBw40THCwb1+l3J41CfXgZvaWoITZUmyFzsVyrlA
Qdm4f0JBNeDAidY4BsShYlCPNEvDTE/9AzrPnbnysGX9NSNL8TTTOzyvGDQzSDKL
+Zm31Gh0ck5G4Tsh5YuZadTuhKsl3riQxW/QYosirdifFDMWylPiH202e2IrGEOH
vBnqkaZ6RK/H3c+hDWxkIul+NuTzmkkmLiwRGpCxh73heQt9Z7sohoeQ1GEPVeEg
1W/xsVY7g2UOUzgATV+9E/49QKz8QTQ4DTnykSfKgzygBNZ9eOAZ7gBqO/HWDJPN
0cxc7XOjtg8zlxpjY80V02KnZw5wDWD9+55Q5boXoAUp9LE5Zp4hKbZxCaFrbrOq
jFysGdMw+9R8BB2R23MIKmd5Re/+KC7g6YehlwEIktz49G8pX6JMbXZt2opkUZBQ
bJxyXGKf9qhPpsVbEYz0lcMtisKO0jQt0PAS7wcOc7XjTPqNQKwI3g95PD7zCnG3
/Qi9YvlJ8SBiiSjD2IibGIW/+F+EOADeSxSsm4kW8LYXhvSkoSbWopST2BFLgtIJ
bxVKFOdK0yglMnpWP5nejZNY/JHKs6RbMMC0vv00rpZ7idYQ7xuMit6Le/RdHK89
WgRGEhNtYWm2xjg2cYw0hHbsDh1oSBgtMskD4BA1S2EuBOfuTQ1/TyBC8NHO+DbI
9/FBf6rzUYi3+WHxD260AqDRTpdVlJ1tQVb2zg6XAkRWOcIph0z+5xgTMtoL0y9n
kdG4pZyXfpG18RUySdvndQqTWo/TXK1NrbWIJtH9JjWylzyE7pvUNk49KoS8408U
ZArff9OW311G6+xgIQMRc2YZe/AU668RhP5ovV47q0TCxzZhpJKEwfymh5DL5Kg8
G7PoMoRyrlXaQCIS1pXhtSAL85tO06dNwy8c805ZAsB2vbarhnNZHj7YDwP9SGbb
GMzw0WWbgatcimLcqQRWpOgphKSiudmJwcZMYeCzgO8CPI9aZXm7bLnOAih82jI3
QxrgkQRhw/94tyr73UCjhEBjy2kkZ6+sFNK0lnXHC7k4Bz2GpVDsWdqOKhXVDp2v
ILivaZ2dMVHdIX0jn5D2HmtPH3VTWqTRABLJKc5fm7SmV7FfnYFv/TQm2JCB1p4X
8n6sFeAYYxG1ZjfNjeA+uclCpZkOR6PF4VVUS1SPcGM+ZcQFPc7bWv4LfVrvknb0
MH6SsS4Xd8pywy/C67aSTi/FTmbfAs9PLgy3OA30QJwMkMJd+ILQrhlMLTmN8P3C
BGoFKhw9Ux/A3bchy6g7Om1e4Rpq0dVmkoJbhzlNzu9ZAgcZB1m6/6p3tEUYtasd
OTaiSKzs11Pz/r/jFlM0muZQ8GrVlCfHznIXaU4k9VgoS+IoUCpx03ez9znvh+n5
XVt7E4r4uGmCFgq9IL8DleiCgXHDLO20yOMxwI1GTj82bErgpLVDuSM7ckkT7YWW
GMFZJgrdYXZNLOgnXci8ffPwAzcB7l/wbtsLCSJKNvO3Z9rRChzxyWaTkubp1WkI
QcMbWTWrzS6BkAQmRjiDWR8Qh8bXdYn67UrWvLHDSWd1MvQC5MD90YSvmAFqKyhS
sjLGpPbg2eagLiPXoCTiua4C4j4rBQVIKIRfcnCayUmyi/c/XbnfL9VeaQ8bbd77
i8omKYqOEg1eh4gNOvgbSfzK9zfqFTN9jQukpVITrf3C2Km/go3/MFs0Gg5NfI46
NluhXXBoDjk7Ota37v28iiDpCDtimdiz/D2EwyhJnngtXAZUlv/NhAJoa5xBBltP
F4nSQ0D0h06u+0+8nbC+/VxSJiYmL5FM8iMREbN+1faZwJw6ovBxqynTvfIHoniq
bR9XxYJsgfKBYg5aLaHHhY/BVC7d/Cu6un1cPDgK2qqx7p25B0uwDa/M4XGv37nj
2WTgcNr4EFbi4VneuwagPBY8dfy6FkE99V1GlMqdvf5Ng0OXj06MR8d8EnmgcpXi
1xWeaCR5kzrUK2uUN/3wGMYOwz29UaYP02zPZURZTsq3H6geMDW21EpPZ16+mdYm
XZyp40I8BW/d0a87iYfez3kaSO/HnpkVMl4Whmy9zAcUmJt8sgCkYB8Cs3Xgd7//
j88cgw1sJcvIlvHxsBh2dUhhsOWNPhife+3vSgtlkEgJQs39LYGkdZrXt2WQVDXD
SESYeHFfyGCmoBovvr18cVHAPpM1U6H7hQ21bp8lOVp+l2FPnyVFje9GjltotO4Z
scnOTXaOomKgw1N5z67x1/w634wMdZiWzGXw2sQWBlTSyHL3ZdOCwjmyC1dJJdN/
fUH16PG3Ys7lJsNP8innV+jStSE7ueGnwPVCSmpMVtPT77WchVt5deXcyc1VT/i9
U3PZTne5qCy2lZ0a/p8m1UYhtcBgT7hFfcHhPtcaXTlcPqRWlrcYG1Vuc3UvKJ/m
VQq7QdKF6pTAhTbNPgMSO198h05K9r/zUsD8T/mpYndvXty5nn0EiET0vktbCE3M
R28pqcdWZpeO9YzLUxYrHeb3RO+iXxKtvxuPHm/3gYpP/u9CFExoIxygAjRvRZR7
xdxvkp3j9knWrbBziVilhM24f/HG/j0hryEmgOMZr3LEk0A5K21yDO2i/XR6+exk
I2p2zOhqUbCnx7LvkMX0SdNryob2yv6vk7RgqzW2ATSW83arG2J3wfWvkDrVP/ON
2OecKl1JKpdlPraS/OXCjn3rhFxN//ksrvQB+y2WQGqh0Anw3GSfe72VRSiakpYd
s1/l15tqIWe9tSYXoHF/eUcC6a8IMeeGiORNOfMpGjHr6dv5aZbQHD5q8xAai5H7
IK0TnV53S3YmqJUfvlc/kpk5VvQbbRSOqmdsJ8SyxQ0PFwlwFfXV1M15Cw+isxKE
CtJwBuLTACFrtK07iHbIExjHRogCrpHKEn/LmZCmYsmRrkxkaIKV2u+K7bL6k27i
Y/XJT9YyGLlGBbDqy0rhKHt6mchghCrQYoShihN63+1mpgFIoacF05QdR4R7L6q3
tbyRsHe2zYSm/RvldvGCzH5649EHRoA5ZaonTmP8BpvPV0mKOfQzNZXUf7i4QHVt
t0zTvwID++GCd8GGVA7AQYko41GZl3PUgxvypHlu/NOCtFoJT6lJqf/Gg9MNUiS9
GOkP0PIfsYKsqxA3DJEWuCWwJEcUvf5cI3e2xsI0lhwPZqNzDArXgjj+eigo/Tcf
/Yk+zvMCgBwx2Wl5O3cP3EEB6YaBDtbbcs/hEO9ITKJ84IKptZ6LXmDomGW+bISk
UUugigxZXLkS6P+VZxf0Kgh58Azuaa+Wv3yqcFc8sKZl1eg1HK/Nobb8oZAtyMBa
IN7W2cx9zmB8RzQbFnXdq9i+08LwxTQh+VEeCTwIqKDA7C9M2u6lHWKU98sFnH5w
sXFkoRDSF/0Gd59G0NYjA5HRyLWipB+CmBKvYkTjcKOpTBioWeInH33EurgQtjWl
eFRU9pPBi/2zcfZR9xMblXi36KmuhDsBfGEEgb0KVgAeChg+SQ5ZVuqAcYGRhd6I
+zLP4HHIXCP+euSUeZHnyZIyO5D8XJ/yNOknW0b/syG1SFTbRa+E8s80qX0uBLlo
9O0dqEr98OCSWWd8pOp8Gd+f2sMsdh+/2NlaDxqdNWTjl4D+xHurXgKYw4JXHWaI
OCNqjE6U2qjNvM3MmGnopxuDcY/ammvxufPwvFrZVG5T0zwE/YuFFMYYMrEKhXPj
FkidhLK4TSfYxpjky/RAr7dIE6WsSU9D8aCRvFCt9WNs+/3dBya715Vn0RDnhazx
d8GcHiXwrHHNWzU8oO0oEGyjsJttCTkxDIVGJNkcFHkJ6GdhtxaYOOuFGLSC+gK5
9gji3+JIcLoA+FzqL5PyygnBAr81yR6G1tNuIA6qyMO7yEYq/bRjmKN+5KgcPf0s
FLyXi6GOMGrJ8WMElpkI7RE5+OjuXiiHGJ0pVRkHOYUUzmwIduuvOU3fE1gumrEX
ewEh0d6iMkinhM5jGed3Uh5CynndLkkbvpwIJQdXIQZIeT6VR3yst415/A8ARxQK
stJ6z9Gt3xNHlkZ5vUJ1P1SDxYMNv1a2uW5pbtMnO5z9khi+clbfw1w/4rVjGpdl
YjXTx6v1B0rQK+sZ6D6H5qE3KS22w8XqregVz5sWWhEYlaIsBIIcSkiJph3qAOnk
CIoN2K80nfcdNsGV+1zrPGCQF0s6MgFCT+H6BefaOLM4dd18pQuO4d8bVDVS602E
/4ADquKL/3E5rCts3sMoSXRgJyF2OLqOeR1bwrlerh/AsWj/hrAYzdD+BOtiRlt0
EUIZoD5Ub4StN6Nk7Aki5G/2cEoP2aiCHh90HFBoyZ+u7SkAgvA2ActBw3vgzLom
kldb/WGFuc10QojRVFNiataEdG0TK7tCe/TRnBvxRROUPvTYNineV6rMlC3KUW3G
f3JduMPRxC51FZ7eno5FV9oNO3iwvgFrjywyNEJjKfMfaK2F93Q4AwAOw+is5Xqk
aZCAQy80qIWQ1YSdvyOHYu6HYvXGNx26JStK2FN6xy1R80FnhJuRNwxmTv02ZrLX
bfsvF04CT+DHYHFbAZc7jKGaZOvp/l+g18r3st+rTRLxhMGNkNB4UJLkeHsqfpl4
iuYBqgoOnJtiR3rUKWdfbUKA87SEa1wj/RAV2GtJPvIJjdahFu+wPBz08GzYHQh8
recJ6i9zeuCMiCpueYxylJoPp+xcgURykRgMjpc5DdIeBuQHHM4OfDGWvZOgLzQY
bvccjkkGcifw4Azbg1JTjtCwgaCmU6vvZhm6QMXn+kkRIUM3CzVX0dy3aceJQ1kB
9rg+/cT/Ve91hRdcve2frsquM92enbBWMS+w1POj32v/y/sWZraeGd/TXAe8EeEx
KmSZIulFViGVo/BMBdPOOZm7GuEZdiAhMoxX3MbGwUa3hwiUJuC2AL1YV1bFbtM7
7dzJxTWpPrkozu26eImJA2b6vSmrD8q/Blq/dxB0gMuMHBMBQGSe0+Ufqdhmx2XC
8Cuypft9PVTFYzNyA5Ce92lnncRyx6giorhQsrqiLqJNKGHSrmj5ttzShi0GxdGB
JeLYqwwV1sr/Byc7FIwZruzreBsr/47SxwUBBkKWtXQTQv8zpkrCyPxJ+C0O9RDC
IVwVIWy3Ha/9ZpwAz6TfqvAHLHMNNckGerTw95HT8CtQetAoHeaFp8jY2wE1ThGJ
72OVEYxctdXqj4lkyS+yd7bIYXviRMeAI9FFRI4Z8N0dRBR+KYVW4G9t4n2zw4rL
4z+mTy5iR4bmOhX8NVCJutYIBnZIxVE9ujBCme4iwKxzpJ/hFm8ZOwNZghEAgigH
9GEjLd8U+uhjUDLcIr/9QCqRkCx9RpYkJ3CHwbIxa+2mZY36JKsUEd4CBvqFa3t0
JXmGFBSTQhfSGol0JjbeY9nUIgiGzxkimpGSMPav/rr6IcXyXcxVFjTmB/k/mhQi
RoobDj32LX8OMItMFQx2i9iH5xmA1Q1AXZ+uBtvRkfzuif9wSBc1PVBJPPcCceJb
psgRn5NnpRneKU4FTcMh1G5CjBGoDRXRN6p/2ifmuHxrGG09RNwUk/eXHHlGHyvs
LVcQunTEjZqyiTNp+EXc/1A+YSZs6ulPsx10U1fnuwCFOiwCeSjSlDJzrEcX3HTP
13kwzDlvrK72OVUMNLFHSDWi/4DRyyBIXYU9c4zdGBt6xgZ+TON+HuH4FOidMfIk
gilUp/gT2LwebPdD+xcCWOdUV/geqaxuvNaiQVfIwtreJ4/eZvZouSb94a88mEA7
i9JpdwbpeFEs5PdM6YpasoGvU5dDhSEpSDpadUAJcE9FV/fm4+D0H8ZwZCSbPY0m
13VuWBsn0XguyZ5c/0Zfz0XTeDBxbLGKAlUtanxjstOpR4lM1XtMPeFogmS/IvTG
fGeLPE+AjwLDZxPN7KLAXjbppGNpDowylnzPi9ibXaCyXchpNQb1DGiUGVKnMqSX
qFwVPe5KxYyAs0aa7ayb5AI9nOUVPKId1u3FFsZaULRITn5hCIkCwugkFRPOR40B
OanlZXgnd7wPywzQRAC8l9gnIMySe3Zbc7mlggoq0knWY7kM0cgy+eFNHQetHyws
yX7ynpkt1+pC6ZGF9khqRQSRBZ5xu8k+R2gbNv5cE8VrylevgWpFgT8uyRmW+FFC
FINPViDzf0RDL+E3mXpAubi7E2PZhXUbBeNQF7brya2euL1+9n1zh6+Iode8okrb
21fb8Uh5N/tjph6tlvGsNLJ94u5ACeYIH+Zeflibq8cvyCXYwOXXXh2Y4pSQI4lb
bbLDRjsTpk0V+DsrwlmK72heTOBUy2NAGVIHUVTgtb3vVGQQcu83xhJsMLII38lb
noLokR6EdsyKQ/cndoH3Lnn82FwtnMwygzXH3yQth1dn2jZFhfuwAZN+KCzWlGba
Wi31OLezqHBGv2J7YHnztyg1urHtf52bbSsJvl2W3soxH6MrAnOwgBdVLd40drzZ
sbNkzkwjHB5oS0IXvVSUl0RYnJnJ9TfEednTyWuG4cHxbjLj7dxKlHVtU9QDetNf
eyuaqyoGH1SCrpMQFKv9GHc0AYvgmvtYIJ546RQmIrQKa6nni0+gcRFTXIJmQOC1
Qf215ZBD8/1rBe4Y7bUuSdt6mr1qTJogAlkxOOJPD1Sv8+2Eo/+xm7Bc8Mq1M3dW
Fm9Gon1L8DfenF7Anr1fcmOUGcrsYp5P9YtR73Z3LFr17k1UPDoieTevjhKTMjTB
TUaOpjsoLjFfBGPOW+NnD6o8Hg6dekV16dzrfqlPO1/DC/imO+h15/nh4Rip/MY8
V51LDVR0v2PAh1qtwOE5FwJUwNW5YorTA4QySdzCnkhcYpmu4tJp2XtbYJ+EbFIC
N5PYV+FGxTm5GsSFt0LmcCSXqVejRyjltg9O2omCbcL5HE1Uri4EuJJrQCHOmg8O
OGdrL+CH0TOKgviCNZA0VT1w2BNyeDSaq73Dh6zqwNheR2J1t1Bz+49p7ns/1xRb
vHk6NAu4aTH+jNDaws8ImewTkqiF1YKoaYUOPru8WUi/xPaUGK/UaRvc2HJshKri
kEBbjgmLA6RpToZa4R7RtGtMx79f1Oke+oXnevmzLsrTmbur9ZuVG2h4mnVX0UDE
2/HQ689Y7A3gvAj/qTOIGVKtnT+QuzdFmwEjAP1G6SGdddo2gKM4e1gZZK0rf4oY
UgzE2rN2dKcN4TQDTvrmP1nvqEa7VlPW6SabunHUgNgKADBNpyDKLrImSyISBNy1
1Lh+GcS1hRYPoYc3Sv2rhnUeYK+u8QEB30o5bNm5VYzPiIMzh344MLXbAcnIFtrm
22AJqpaSlM9/XJSwPe6VH4P/hXbcFN10iar9OWA3YW7pMVwjc0QAPXpwtDnOOcw5
j7KIOjmYTMxNylDCwXPYhz09Wq97+1RK19aXP2zKRVBCg5uRrsh9+WcBgExeLMN9
DAwxSFJjST0vnncsDgU+XWigIc5Ao2zv0wcXEmvWUM9D0Vg6bG9laHdiArL4GQNR
StrxGO4LtMLY0JY3ruhAQf0q/HCE4nDlYFh351fM6E17zI/6965jdXl6SxsyMRUM
/8RGsA4A63AzXlok8WqOaSwCJasXImyahJWCtLMXptRGrPT/pnrbYwCPuWmcwTz/
8FB1e9bURiV8emvYx+w7m/0pmhQl2xMCoGWjPsOb240BC1SaJA7J/LPecoaiFvf2
Ip0oR2lu8q+JzhbdCM/PRXpiUCPug1EmFYfJr9LDz9BQEkiD7chHqDlGC/lZIl//
kfeCRnixd0aBTtT70rWFcXYo7Sg4H3X5H4z8gi0Pr98Pj6cxs9SGu3oBlTCCgQ+G
Um89AV28qzw2ycQ9PVmFctZHYsaF+QEiShX+Ea1jEBTRJ0fyuFQeWAGjVULjlX5B
pl4zy+30iL075OsQmlGvlg95wb4479sn51xYBA1/5c+A7uLXsWrI9HkLXwiVL+sK
UIF6nhiNF9rnlkl81Zt6FgF3RF4AOrGetKQ16PmuhOoAoTBKKVRRaezuPA5eiXro
4IXixZNJ+rnFT63KL+f2HW3rAAWvcVmGKlbuIVeXhOFVHAHF6GbIckCUvRnbpkpr
qf4fD99H62yPJIQi24iBvPhbxxvRs3g/tDiFqKdbrNw1aI//2aTxmN3kpkVqY+Wu
77EBSgMQH7hM6GlD9F01owyTEt+GR3Kyy5FFw35aFQNXKi8YY7a5+6zI/qcQo2Pm
JDMWirdDm+egOcuOH8CAIPM5gpsFvTxES9dnY79oLI4xT0OYKdFwPei1lj1RRemy
I1IGjCV4dP4PIiRRNhTRkJ8QZAQzUIL6DhThOVflbtGNnX6uSLkK1sWOF/7aAgN2
D/vgihNrfdkRMYpvHJI+54JFru0+pKeV2i2f5PgKbEd3+NZ7S6TxwTIaoo4FDMqw
47eWjOp+7DInvrGNYFqMLKpDHunu9sP59xAPGPXrM5V3CwdLOmfikNLGPhCBzAGB
L3fu14VA8lV4wyd9z1tJ5ygXx5hZ8/sAeseAa0vW8kGc+V44Ojzz4bk/KQuefWX3
eH+VPbikRHNDvqMY0FGpPrH3l4I066V8EFrhj/2Ydh0wjn6IryUnscL7y9oeZvNb
HeLOrKuosSWq90jG88cP7wJOdwxUwjUJ39oMxZfWwu8KAV5scV+i5bj9LbOtTobz
xCaswNNWlquS/YwvJ2DVaxUOyougX9vQ6M8BZTm2nTZqC75A+UjxJApRY57lotXr
kYEpk3RIZrzFczVJFxbSUO2uZOOPw2gB0QPyhuhi3WB7lid4WzRuDMxttnwC1M1m
FjvtTYLfors50OHiuJE9htkEFoVENE0MQ9AF6UUBBY60dQqENw4CTFpwKO2YjbG8
6eaRW5nfarESPSo+92YJJMRhj5dCZ1hmr/J04yfNKTJeLUn2nf0ZNaRB5VDxAn46
QggQcqMxlDtPuLkiQ8cTXWX2zLlxkMaLCR+iXGlP6kGBy47ufPjdluvXBYBIK9D9
YOG1bpJcIXJF5wYPUaEINmKBMnHFU3DXEwK7pJIZLsC2+Xe4wjVWcuRKWIoOU7Ln
3/0vJ1qfxiu93K2rt2bwXVk2gax8qZH7KSJMqYh0Fn+LAVn3DH5b2FXy9lAcs7Hc
kDsR/WPTsiaSHd85MYE0jlyhOSMJMn7OpIZNpowaB2dHUsDI6kMyW1Cpf1cSVUdx
yzFh7RkoC2Lzfh0D89YBbBmQ91Gjh8CvcjlVSqpgygbd9ovyCY3UvJxf3VbJX78l
17/RAeCl2FAUe5UkdXYEJawjZ0Td97prJfiypkWnhjKHAAsyLDkPj/tarDOJo4V9
Xy0d0TrQjJawaZHvBpFv/R0p8w/5+2/WTsjWhArKDWUgCmuLq1aeyl0RHp+jfYkW
PwrhqiWrD03Hzyel0U7StK2D+nZ9eKgA/OxCxTGjCJYRX0/+QbTXptkoZFARVwye
fS7QexHfCaNRpUDWhlp/bpCTY+js4qH/x2E9697BVRc2berWaT5aW7szCSot94au
8xixOTldodKT2Hk3XKi7TlHaFvFNxTEq5f0eqkKmmnh0/RwahTmlRAUqTWsg5sW1
/LR/65udvaJCX0ZFEVFRwepg1FdCWdS9MyyllFWnABIV0EMG4ERQK8vLObDOzAsc
kxd7LDAsOLER1+Zg0s3RSM8PSxU/h2kz1LvOVvMeqJPagiOum4xYRsjc4Ajgfork
7v7Zf0w8i5xral+0fuGOMxomt4H0i8Z9oxavDoSsSz6LwmKohHGo4QkdhSyAJvKb
exJLBmwSVEGANBR7s8OYxyPt5QO5uI9oZ+FuBC+EybMNFjXdCALXL9YCEb2SOdXI
05SHuxl6NiLt+zERHhOHHfyQW9aJfGgrOGKKG43tN28dK/uGG0iULI41W7itVDUJ
USgPXvXnksMPRqQf/LgakjBuRiZys3URpsu+W7yG6r+gOp+IoK6wcGmR0CSHyEuu
XI87HhmnQSZJNZUCFpzaSQxBRP5H1VAcwtL3fMJ7KaYFlCtoj/HxuFdQ3ZWzIDTs
bzcLcr90F4sA6aPyFUw0WQQVqTs0M8JrNNtXAb+GKzM6qqx4vLZ4Srw7ZEqiZcaG
7/fdLLNV8YFDLSbUO4DArhg9lzhFwXHNF6IrVUzwF/IYZNLtqD9w7clafNJlT36w
9HmO7wsi2zAt72XjqEhE/gLjhnSNKwATkTEYa/keMrJ9HxA7vLVNCdl6lOC9d+bL
p6oYgZNIPZuNr3VARM/ineha3jHTZfb6P9FMNinyTJOPUFX0igFgiIOTqjJg0eq5
KUC5H+gn1ixwQ3UrO3X+4IHo/T+ofKeGliZNdQxaJqwFJYxvL46JVpQ4HW6GSTDm
854qne9O7caFO7SG8VJ1HFjZd4BSHb54kkvf5HHUDQiAYlL9JpQrcnQKaQSdsVgY
b4ONr1DVPrZNMcq9h3JwgyYx3Rn3rFaTTZLl1Tlrtdy9GAtFqqSeUIMIMpa2Bfoz
P4SDOroFcUe52fwcCxLAsE5SVL8eFRb9KF6A2hQH21PJvtZ2AqTgO51jhEgxzgpI
XhgTBkSMvLsVSJORMw03g5ZYai72dwCtCkPXUZ2xYiIyg8m7y/kdOIr/DAnYnUe9
lzkdt+GpmOijFQ5e4wxW5c9+BZNcizTioA6kCGPsYJjJXHaMyatiIXj+Ps68ndvx
PWk+k/vjo7gDjBUnj0S5v4t/lUiaI4OvqEOo9vvjKHJpx/ov4QP3g/Eo6GlDmrEq
XkHmTW7xbZR6Ub9AvDiOzpEMT4w7emB8s54dgZ0BX4/oaoXHflQj7RM41KEMwN3E
yv4kV7UiPW5nkVSMlPmDgDwszhXdaNMLIVIhWTe0iq2aR/tMwr4kSZsl+HSE+ui2
1NFlHvqAluEyBZ5Jvk51yJ6z7E9QD3+2ZxybYkbLZ40rITEdRVrmk0uZRZ2kcABp
SjwNL57sezMhzpnqck+wAftoVEH7Y6reZfYlke+cbnoFEi6Noao1nUYH76uEjimC
mNMnNAlYHtcEQJrs8pHVX257ssH99QTY9Gyljb6hy1lR1BNUcnQ18UHbQc2Yr88o
C3nxu0yPw7tSEU24sguGF5NsUEwE9sIHzNiMrF378W0wZEgwhePO/6K/+dJHKxMn
tfWxF10ubohYnZ0f5TRhktBM1qBTmRCBqeAowiBMsGLy1e/kJScosZi0FJT5SJ31
JcASUaD+zKQ4ns2xY1/CBrw9hc1bH6GVcSIDd9A1LisolX+hLm8mzJBBIXbi9Ndu
exnJSfVBF7Pw+cusf/9UOGNdysekLRluKsIUwcppaHmk+xkVAekatSiL3zk64nsi
c0bQ0snSR9i8QkbiycIRsShrx8oAqH3LvLO+/4bkvm51cSIxFK59BkaKQaHVli8s
LT18GsHv/mssBazaSBV3/XvBBpFynojmjuI8TEH7ms/85ff9kBM5pX7ohxnaws2K
Jq250H3Pw/FfC04QjcHtOBotZBsd5Q0WTPYeNgxyWHo8IqPGZonSqWc9N8zOGT+r
+qEmD/Mzme0Y0GNJ3B1jubNMHc+AOyeiJ+4uYA03rYvBiDCv3fxlLtl8F8S47HzS
GHfzKrC0tYUHtwVVW+pVJniCxKt6ri1SfDY8rnhvkGJrf5o1OjWr98LSPYFr6Ecg
Z2HaM1/cHxZamO7ENED995vBcrI2dJGsn5zNVeFRCF82OsFQWNrkDykH8UiAAF61
IFMKNq3oIM3D1vZoT2/vvdSbqbMl2MoP90KDsVp14/QZLonD9fRw0kBkx+IimVPT
KlXlBOBU246F40fGvE9OUIqlkkl3DcH3xndE+9gd/YxL3JFkkPe8lBOy2el1NlDQ
mowX1kawvbwe6/Ii7h8Bmx/5WdTf7Xb6sdUZCT6UYtRK5wnvGWuuDjwv2eUM4HBC
c9wK7F+Xe2NGEwsXKV33OPqi7A9QADhGrex5HvgSmFau8FZH/07FqAf/hVUGQOPi
JjhXGMXg45JrUUH7cKJc9ripxcpg/hl8UBrRxyeTHm8xCr66JfdH54f49HrTft//
1kQwFJP/mFI8eNu5AiKk/bOZXn9dBmclEOY282YjnZY1mSnJcrf23HCXkeF7YdJw
2f0QcTPEwx78pzigSE8H4//f53qoGCtB2RjhFHM0eW0cSrPVMbI6HS4FNKUew0iw
RaIjC7KkP7WSKlEgeARio+9a3+5QqbdWRDXjKFB7PKn/iTbjR+nob+o6cRw4xLmi
HBMVmCn28T/wotlEdhvv+fXwrgfOmmaeUJbhEsluvqmdwLvVGeQfvcKgZaZFp3Ri
BLz0ZZXrG1W7b3uH8C36HpWlqp7uMK/ZLA0VsPTt90JBn9jqPefowkLRxa2LfQz6
xzBlz7fls5lIAHgjIoxmFqx3g2Dl3EkdTmCRgo0lkzgNRZzbThkYOMMXYS5VCvHK
na0zeKnqOOs00HCIrFWBewAtQyP47zlFSJ9uJ6Bw3W6b+1qegfGgXPjd561GJ1vn
jqBBfyaUdBxTlJ9TEivNYvgeOf8zEZH03cnTSVjwHMvWj16evhdUcqI74DCgWSw9
0r7zSVgOgt5OctWwgIKHJAej5HNat0aWJQKs7tOtr0KbBO8IMmpm+pSAKGVEvfeS
G5p9IM3aLA1c+dHAcVAy38FDXvBMusrmifFjIId046tddT1uvpuh5eZaMbHHxQ9a
RpWSQnmm6chBNKgRnfQPzYjWytGzFyz6FrPum1YpiE1L2HaH5pB+9dVL7qBjEVll
XlZUTKGpAHjiMyVHMzkGF0NgQr7manhk8hVcj0PWZazAPQFrCu13zo204yM4jgBV
xzDeQ5ba7rPnXG+36vfa/og0cGAaNbOBxSdoQ1rPH6JzX6wU6seTYdkfzeEnXea3
oBPdu34J7H3zc8lwfQr4fWsnkBlcKcWfv7upKEGJNZBzMuO2LOXX19COpN/6y584
/DArfPv1V6rPkNmVuKWZ3908mU1P4xM9LuLJjoTxkFA4SsLwoeR/VWsoRvSW/EFy
z0lnwvuzGCpjJ1CgSfcn589JJaMTO5EqnzxDiGbFSLjeUTaRA9Xrs9oLNnuJktjy
yjOds8Zdcwkp/wseSGKABsUCZ/BHtwzKbQf1fJGk9A3w7SWQeCb2Y7Bn4PBmAEQr
UOyCTSXj4dzXCbOP49NWSitlT0faB/D5yZGBTIwrLBygUE8pKF+AXvaitAZ8qvG2
Ed5fMq0LmfVvnD0alKX7xT0pbK7sdoU1TOoGmCfVoZF7t1+pAaWmYl72P8uc3l/l
Q5/f4L5yUHdg5HBuxGXtRhOLPcFn5yi7gUarKWZnOYpcT1qDopWbZfTneutpJRbA
WFwG3yM2vmKSnCGYzcPwKqNJ3lwwIElu5oQzqXtymW529I2qVvrXbZ04e4vwZZvO
thfR57TnCfm3vCltjqADfAyGO6ZAkMvBE1fbIC3jysCzQqn+6WJF6sqs88Q0QM2T
aXEEmZjFJ0BB7qEqfc3dZcf6KY0biU9Zo1yRTH4vsMryQfj88LHHjzv/muwOWiS/
fKf3bHOtI1ZuzyQr8YBKUWYbkMfw1xQAFKaoGaFP/OKvDQ9GARL6nJBvr+7Pg6XH
Bq+xK/XfLtARFRmwUwrZyIOBA+IWkzkN+NqbGt7sKrlGroaR0IpUglp7JWwRVhkh
JVscFz7XOvv2sncSbDWx5ly4DQ2KwZ/KUfdgK7pibsHedMqbtZ9oXTnoSLHBZTi4
HsK58XLwTnlyooob/+weUvPMfaICiAc9/uiYERrSyBPyjCnGOhIp0AtOnDsFzdFp
xasOxcrw41RfvydXD33hB49wOe+oMwWBrmA9SEECEtXMBlW4Wu6JxM2ogsGUR4Gq
7MiTMQA11FgUhk+cjr4qJ/p4Br3UcAaPSNzhRSoLiCHMispsOzY0pOYEOd2cjfjJ
/HJcrLVX78NiziMsl0d2jiaodt4JrvdVNgX0ThXrVTswNzHQZJtZH0sZ5WwGye/O
Ns8RWRiQtdW9/NkOpOJJ45S2tGHJUq1YieNJ0iL3GPUq+vqV81ftH7EHmPNnlLbj
MB26vhCq3s4DLbYT4G6J7xWrQWdTkNcnRfyRYZJIyFlxZWfyqPxt+m043qMt+6WX
APnH96tXOr9gyL5LDmM8y+cMZQnNaArLPBv/CF48ztPiK+rfPTXky0ti9pVEvf0q
64Y/7AlxtXfBUTNB1Hv+nV7HaWbSkxEPVEXy+bTnGj40blOQlo1u/o0x17pnjzaP
VFJDdWr8sBooYmwV8RH3hbo8ojv8BiUZg5m0P1JLW+w4GtNNxpH3IIfm8SHENEgu
Rpu5CCBMpka2W0NK02wi8p7D3R2CgXS9dpOr3eCh3RoP1h2xH7FdsxtVSKZ/f7a1
NsBligeZT9oQvuGPucQn6S79quZ+p1+/692ho4pbOhzcGSjNYVs8bealgV7LhuCG
AH4k3ef6fS6+0WoaCjYEFeoXsONkMqLqyoqow033l469Sp5mUjS7YJuzTeASwgzP
w5PQB1LjKcplHv8pvM4HyFyYVvayFTM3hhZDoNyRjufIUba9PgTwXyky4J1LWGMJ
KE33UTaHCA+PIWEqDjUPaq9Rp0/kAPeVqLrXCv9x85ljwD5WIFB1c7C7EPce+9Sm
rBD0ciAp/cWt1s3szQ31iYgc1PiN7nmJ6GHwzOKgVtPHxA+1p7LU3aBDNnYlmmDP
RPB9Bf745ypg+DICRsntiyfDpVpOesXN75GTilVaz7ui+5bTN0CUScp7MPfFuuXN
zg5VDFykZakUGJGFGUko4d8kN77qcG+LZ/1I937Nh/r2jaoOrzd1dqfDTk1QsyLb
hNruTg55DHH1E6B2TdNLp0fdKysQVf6E4l7ZgNHgpmXvV74igrUCA+QI7AT0Kcut
V1Bq+i0ioBsCGMAG2PhaJ9AuWVNLUvRiweE1+i347MNoJ79VtjHwCD/dfkyAYWQN
vo4btTLcDlhPQrhvXYmNZYA7OvsYS9iIZr4Aa0uvkwyhm2Ea8RlHjw7XPpNtdlKE
rw7fgR88Cqg0QmlkLOdGt86VexXvmTf0QteYE7XBgxzod9sAAM/NGqidubUbri5v
uI3V/SmClI65l8g+XKL0iTU2znAecFGfNbVIf84NL41C6MRQ11+xVMrAyr0ZE3Wo
7NljoozMGyZXZzJuWyl5RkpaBl+WX88sxnDGUN/1Kyn07jJ+npkkBJXgoiwgZf6Z
eredkQDMUnjxQswo6/xWH5tW4TCSSTrWfiDfXKMe/TOGc1fmtXbX/CbS8Pv2i8lX
s+KdYJBtynDCGJ8a09OcYWrUBvpaYZu84Eqg8Y5NFNK11RkCaI3mWWeu7xoyVD/Z
54rt1bU5A0KkUDHhP1QIK3YNpPUahwkTKZXySBbB8Qs7zhkZUYcrlH234Nvzqh5n
PL4iEFphgz9nU9hLDzc6Oym4hVfpJdKOwQVm4KcWRXxiew4ROIMbp9qP4+D3GKus
66idUPcFiA5kD3tjHfBffrlyyza+bCtvX/lrk7yDNAQmExvmFcWUfMgqx+g0/BuE
jG5IGm8pWHFU1Z4g73bv7RZsJ4trXCS4YEA16CX83K51uOUapRiaJ1cMQS0ffHfP
va4VrO0715Zet8WrL6rlxOBoWIqTuJbOoerOVOeKHeeN402f0sGEbisQxrMhOiMd
+dgTlvaAL85e6dD7L2i457Ol/bLs1PgsyVlAVa69M2cW7cMxhM9CF9vf2uReWw0W
0lQNhMYKtHVogiTlLYzIjCOa/JGGfMZb27EYQpUI/nkFN7oykp4OW1Tq6bKgUZtP
XMVQdB0bY2QMknHg/AzDjNdG7/sSVQ4tBhewbhwX4OmaXNcQvJ2loJENfp4S0oC/
TgcDP/A9PatTvc4IYSYGinzljOV0g03ukDFIIB/v6WF5yW0qUbsX9reO2A3n9zOc
u6l1y59iTN4KF8aZMw7IIwfXPJQMTjU/4UIZsQEdZhFDpA83YP9DNKtDsUHFkNOp
0sE0KOwAYDOsoALJti8/SFy1IUGeawvTEShHRIuuqqxqZClBABYvsrv1CLBrw7db
xaGHqPoLJGSWkcd+rSygORLxDOpKzuS9229c0bOBo1IO5vJUBVfP6P90jOpjfzHc
D7UzlSSDHMEHWYyuawVTD6Fyl/AIliN1E6omtaYGfc0HQ+QD5hq7hisEzxP6RlRw
wFpenBHytinwdcmDTjqQ6W8muvW/vBKTyzsVq/TCdvrwH8KR+q6aiYdukt0f5mGD
ZRm/DCXDUiw6b2ILgya5aFe5GbgTsKS7LEG4UYPwFaZJuwF16PLrhOTt9aHWgadb
FI69zvVUi0Q0vd0rk5Yr1bJdTs82ii49NE+iU1PbVY70vuc/PjIPVz1Z3xc1esyU
1lVaRHkf8e8LhhC97M+q6aWS7kaAcShx1aZ/3aaGUn9A8CMBEAFDi52a4WpOSCe5
V9sZ2wAUusZqyeub5EV2MfWVDegI3ZoWFROtYkqL/+p+XOW+int/nPAqBFjeAo2r
evxGlbnqoYHIf4elZaQyK+NZymTAEVQozBZn+WMIOuI+vfiioeSsFbPy/VRHVHHC
+5LHOlOvwQ9dx1hWiqWegoxvqAyBLAbH8+FgNazVwiQ0pBjckFM48A8h8mREvBac
Lqj3g6fdgaqcL8yNFhNrknUYkOipmUpiE37P89UJSVOeWkAfuJg83sTBkLaKTC6Z
eXvg99qKMxsABD2eiXiKEWjw5XM8v8fljnzJUrkXLmo/I/n3bjDtHkeqxMYBoCCD
o1p5CVa1czTliIxh6qjkm/zlO3ePNKEcWlOg7QFgbToBQnxSnXUilqOhKdVJRFVK
y1EVpS0MBJYqciIIqNb12gp91K/d2wbEx4rabfW0N4sQs2Zg8PUUt3o4boxNxOBd
JnWJ0XwdE7r+0hTnfTi/qUyUOcHhXj5njfNwwsT0/4R2boMtp+HGdIfDfsEkUD8A
6MagMZ0uU+7VhlyMr+6A9VODhyaV8gVY+k4U0AAsnsXXwcgDWghQx/enJtjZUEoD
nJ9ffQMc+oJlvohye3h/21nG/ntQi90nuybOUa+4O7R4aeJFzCz/DqQSuL8OTqPs
VSqPUJ6it7eEngX7cRcwuj4sKpW1pYgIzJVqAJNmOs4RK/+QSSWFFqwNnDY+XX4I
rWny47xFZ1YzMIlshAh/E3B39XFA8yPhQAIzDNr8Sr5CE+qzKB+qBnKfQw2DUc8q
pCmaBH3xny3EiAsHnz0pQdPTOVGp/tRfcaE+lXaAVlt8CR0axeB5r0+CqRyEDll6
qa7SzKbXD1dId4L8wLEP1UuTMC2wtA66LYEl1JYiBbCUYjnOntxTA7M56Qpp+WsO
8YnBsMvULjSEE6B0kwbLEyYtoNcFV7RfhJKndWdP8ley0dgCaFNsv/ePjc+nCziq
T5vnQ4mBpXKjYOpHowk4KJe4euMzJwW4oJX7KNyC2c5NgK/+idBxwvQSftTZoGo1
UKdM1f1B6AvdcErcM4NRMqkG8u+erHc67tGNGDEqt7So9OJnR6+Ehhq/Ic1/V/I2
W9ZgeualY7zABTXf0guuPyADdpyZ6cDItIP57oej0YA8Zz8VK/oxkyS0M7LhQDxn
PyCD9bpclDaAClMSUhEkZ9cH6QxmBELSkHZKXeVHY4koMDYqr+MVBnWmCixBFgsT
E479P59WNcL1hTLifCydx/j16JLyJFJHbn8ICTQsTRU2y88T3Xp+IsBp9A9nSawT
R+Dd6RAh3j7vssbk96vKYv1pZzY/nSdBO2bcXXa33LhqV0W9qjf4U86oO2okfszn
t4F1zpKJKes/Q0fumqvHsP1/59sld5ZohJ8cTZB1bmqIENVWMpB3DZDaGqqQ8+z6
kZdO2F0VCGBPVNyvxEYivC5PQiGrWj7DAZ3hS3sM3DMhEcLYjXkm8c9oHPb01boU
a4itBel47a/DvSJbOtqhDYLvYGrGXbhn2tvHB4DJclNtjKX4+wQ4aaWU3u8ODmrX
9lbHWZawPpr1/fUpygYXISFVuJEy6+IyOCj+Ycijm/w40RpCqgB7CrQNC75b8G+u
4Pg8T3OIPre2caNsrRhShxock5EDZ/6VgS2WZBNwzyfLTOzjgZ+WFl6kG2+CuAkF
cDNFvzK73KU5wJrcsL+E6p+Cg9qipDe1ju/St+WzFWaOLk49B8pzltTSXY3D4Lyl
92VEYKBox16U7zIKKjGPvlxYvnqCLsK4Upvisih58aiSRpR4SPLLNxOm34BHgVFC
tOOv9Fdm+GJCZm0C0QJYJvPdi++k5ehrAsdjFf53t92COOrgH4GUMiUeIOMFfeRY
Z4zZE3wAYEsqVS494c47s6FkvdZRC5+kS3HrbmOpsq2xbBuWaOaILseAmmcV4A0G
meXsZPOvjxVlZmDYj4DP/YlQxHBQ6QmOh5185vkkGcQ+gwSNuumFQAl5nlvJXCbO
wcDRVhsMGCwpkikpK1v+LTbdBYVJTZ4jnoPs0YMbilD464BmpvZJX1QdPBxexlQq
iW3aHdPc8WyQMHXFvMOllXviFjhJZyX7xCTkdIh9HTbgToL6Gaj8M7jS9JrX1k/S
BnwkOxirsZ9XAKpdIX4VOxZ82WX6CisyxDAaVzYVp/vZA5yiCAEshnCLOum7u1CS
Am6xyFvyEBRwqUizz71EQisLNdcdc92ZdBEmydcIQi10cjAYJQli2t5AdcMJP6Yr
Mi+hBafWJlbC9/nhMjGStowS18vrA914q0bqOU/iEezEIK/LdRGvrp/vAGxQsma8
5zLvRK51nL0X2Sqi8T7Dbz5cecxBqpMJH2UMwOGrPGCV7hUyLQbTUk33xCOXxAIt
e9kdxdKOrMbcfOviepqYKetN7Vbb3kKWRDbo8zeumIEcpqmyNTWQc0I8ZKLBD4VY
25qjwzVJ/yfQN1JAUnfTDHepoiVPOrOrFrnGNVTkV0bJWPEAr/BVEIEjQul2HLuu
CaNwBRVmsY1NtmdSW/Qm32RVnDA0b0xhRP2tvLkQ4ArbtlfxCK35GhaW/5Sls+XY
5nHKtB4gIHsCFY4mH+pDr/kxY8Ivw6Qsv/wPq3b8Sq5+eViPS0i8+3nok0UXHJVk
oNOPJohJCnI/LIu84CPzKiiTb8gsypTPLr3ddGYqwkaUPUQKr5zGgFW8V6EnOjn1
ZxrHEySOYQYBW1Z/RbcFX4eP7iykKGcvWJ65pXO64HEP/ufXTDp5sws++tFJpfXS
F8qnOxtH2zMPeMiaQpXTwIDErN6XlU82XwcVtF+hd+wz4I2FxZeIRn91ScyZ97yo
KmUfY2G8OjevCV2XhXh4HKQW4zPXqYss1kjoIEF9jAyIJN5oLee6Vw87n8UAWAED
Lsu2ry9OlYbMaUAlDv+PoE6LsBKD3P05PyGHEwHE0G6YGDHUyJV/IF9Axu8Zb7ZT
pKKl0ySr4yvl6ZWp/jl6Lq8/qIJdjw6q4NBcuGqx9bRI/5M3BSkaAkVw9NGbjClC
HVO3TRXmLL/r3EwjfzIfV7VbLq3SOFPcC+RN8yOmcg0p8CRnWw7i8bmly0AhU5al
OETLqj4iUnR7rUb9VPIJLoPNB+iPPiYwTDFXoi9ZdlxYZ2QB9J+pmybVv6oPbUnU
5JVghNk3pQ1KoM+KeGrbJGbNHyp76/WKZeraHWcfT1NSCl8s2LBvsGJSBL0wvujE
a0Bg/u6j7TicgLMO6RtsjqTkA5w3KIgjQ9JIOygzbUzzDUTlh20nTt7+/puMPA3p
CenS1UhGWhgdg2E+vWeyu/iXFsMvWbOBPggOZwYZW+jNJIKyMUcYGm9cC1WyJAJN
lSDrEQU3QZUiJdOA066VZHy6Fqn4eQjyf8BA5nwvDc3xJRg4of9CPe21KIfmshsI
G9HQPH4R7tBz6HeOJHZ8IH0jOnTmM4uRHhZZXe/6Q0e7PuhFdXKl3KhftAzgfSHM
zy9Lcs85tadufCklfM6BqC8B66A38I47xaBMaFXdP5LDFwvMYgqYI5HDKO9sobEp
W9wOAKBSG5F541MlRAH9DvOf0PIKbKsl9LHzg4eBigto4m3MFCpsywe522h1ondD
XV6TGISwv08O6XxBWl428klvujgW93TtbdVtMFoEL0l5TWoLeyHsLph4S1o8vD9e
WHNQsn0SH15AZfocDskBEa4MMB2sM+TJ2fKgZWNCa4cPXSg84W5g1zwWy++SoY4+
JwrYV7h1lBK6iZ2IsyV5wrl/U23VmrvLFHIC+aR4enTN9NSmpbJGRR0uMnEeLsB2
fmGy5mNAU+d8z1y0/B+0Si0nTPNyz8Sajk9jSHpBt8Py4Ka0o4lGf8LIYL4x86NK
llgE9KrKpN4B3U2qGinuR9tF4qE8kH/w230H+lVBnCYDQTiGVqU7Moj3bcd1/zHM
rdHPY7O3HPOXKTT0kSbt4dSP1l2zgVoRgfxlqWhc3stVbdlybAHsD5OQhlFqgjfa
l+K2Y5xowgdQdIzSNEUi4FYvK2bgueQeLKqSeVKuh6pz8fxCyhtwC+R5cdzRN55b
z4IbnuO3f7/TfERAD6UnqTcbbmY3ZzHKX28um7giBvTK0lH30hpuDeBV3LNNnrz5
yKi8bHJ2xftcT8jw3WO6ff4QYgFENhaqFVFhIsXKpF3DyFwE453Y2G9QswIfrkPT
qdD5lLNfJ1D3022Ys36OEK4ZE4+7texzXYAOMIMMf2I++3NGToQb7u2GPYjkPJKG
OT33CMn18CTPS0BBmwI6pu4Fix/cERFLo4etJqHT20s13Lubp35vJQdjA+WVeeWB
FfQmfEEEC9CjB8/U2NC7ImwsT3H8p58r1QcUGBghxkG/+8J2pWl4eP1uXY4dza4j
WwbVBG7fI80of8EYvWM9YmprRMiweI6IFeAHlgLJpdNkRFjfWBkg78AwS6FDtV70
hiaO8FlGnnVX0klhiq4oxzJyuq38gFm3vMbBAnLzN4lcoEo84JS1R4NT/RUekus1
WJ6F7jSzjomLoMcoZ6oBi2kN4IXKB1B095fqd7mkcNCAsV3L6C4xrwYTY/zGpDL7
xUO5yzkZiA4bEtR3NuhQr6qzJWeM37sZnE/2GBAlDoWrJRYeYUCUQXt5h0VT5gPR
J69qX86mqSMl8RoTtkMtKm9akdYTAA5dKMmb6xw0DAeaqRwNSzVMp5MGsr31SoW9
f74vsM4iLRCyrnwsKStw8V36ELjonDJoblEXtAbUA/aTIJydOd0YjX63Uaorr5Kk
UHp0T9C85v94oBgkrCRl3yZo8Ta4AiMckZEr26bZtTLHc5Gb5UNUwjkzZT4g4VEq
gJHOYF5JkvqF3fRXhexi1o8mFgliNw++Ey3zgkkSFitD/kxfw9OhUxW51eQdq5aS
EnysvKDEj4tpluIXHWNSsWnIQWk1q/93FuwtrsKG5XhrU5c8nM292zUyu9XyAgtJ
v0tVWEs9pCNAeWMRsByTnwoGln2h5mDaRpdPqnSPoAV0wnDEXwecS27RaoaVqX2G
N63i7sjFipxEUyy5yt73Zlnu/PW8rEGWbPpMWcGBtOkYiSP0SzfuyA15nmu9oHaS
OLnVd35maAUZINaeR8R/haqPpQ8I/w6x5wkuz46xYyK+p9sWKkYt2HjG8uXFr2oD
PDsWuHWY4yII/hAkoc/EndlMYbwDILuLOMWxPlStgM2hYDEBMTyktIlTncpGR6Pz
n6ftUDwtcr3macO2A2nlc7Py3+V/flnomkW5CmMRB1faH1pq2otxPkwgeO7rdGeB
fMisYkAaRm9QWKUqqhYc64ExwjwkZye9jGnqUzx+6PtAgE17pCRbkAfsPUTwuzB8
DjP8+7isge3Bbm7dV9QRKBiXSRUv+1emd14g5Rs/6g7IMS1wp1JEw1TPsoQrAqKf
151UE1W/Sk8y5CbtNx+FKTv/7Y2WF3CIMf4JNja09C6a8bPRHnuybzgqqGwpM+mZ
4Z9OboLGdIx7hPUkF0neC8Ej6MpZbr89pPJUoRPb1tTOcss6+Do+vxj++Qs449u7
8QEWcRpGWXTwHKohw39+3pXv1o6wOOIs++tsZIBOMQnwNABJifAJI+9g6Z8ywB9h
NytBbKpbXaZ354i6pO3sZTCj4LYfcGeRckQKzaFGQGmghpowChhFlSmQkFb/G5Zk
oASP3tUKuEZcRWDN352Q2ke+grF39hD+RAnRzOiDerlyGqhqGPhzWY5Rsi07U3BI
EZfri/ii1Feixzs+fTl9Kb8uzlivhDBdauwaVqK0q5Xn/cPScXKFiQANIY+GoKnD
0EpQ5LtRv1scszGH23GdulkUy8Xh4iNURi2oTLvpzggjwOFgL2TCme0Fhcz99sUr
/zqcjJx5r4gcneVxHcyOrI7buGainHvQ8bednskzSOoJqM8OwuD++OYgkaqyhMA5
4mlZar7mDjQmXjruVQElVukiagihvEABMqDFjHKatZC0mbe8m1nSIc3Z4uBiMjeG
aLi+dykY1YIU8d3WmEpclSWiDUEJYS2XiT3m8XHQlM+H5AZzi2ECISUO+TePtb3f
M7iP+lbMObPeV7uRS2ylSy7He1SPY+TR3W5f1FLL1LG8lkbGizCi108JTNxD9mtA
e9Ug2pGNpq0Q0nhlRN5mX7jHBIKm//y49PRvJ4UbFCfzmvAUXMeawcHz9ZRnaY/G
5yC3vgzJb8kabZ7l07jupnSuoQYC2Vl59tpF1f4F7TUGhoIZ3E94OnDhTjVO+ah/
C4RgSoTmgrP+8POaKVzCY1/vJmImZZr4T4yhugx3VUDXX3Os5QuAcsv6HM6Nusj7
HDvTyPrIBLDcQWT9fLS8sp0UxrCOzRh32+lUkSfoXUibNCh3ZFMSRQ+6+Yzz6xEm
Ca60MoMzNJOsvoRjjt1VoV6E4O1z4yVBSI3hpM6uFS6TdJqBlNyGsn9981ebCWCM
56tBRGmHABDABBgFHdcOXoFRJNuVZKutj2UBtVMl1uaRhGSO+PRD+lLg8WQ2lvB2
IA2+luXd/xrIdQ7STSvxlue+C2t/E1GHcBItk+poQwKC73bUBlFKdbtOw3gMh9f0
Ao1aXYaex4ODVY4RFsghc0kUpMcvEFydCDaoS/6PzQxjKDD+aM7PAFL6iyV30tRP
/sZlPjmiH+2SI4XIKmukpygAAhkbJfJCzUYV5e14DJJ6WR1YuV2cCIRjc4gpf05R
wsR9pkoOlQJjYfr903ovw22wP3HrjG05t+HNpjiBGU0YkHGmdSvAYk9D5vbSUchk
tbSLM2aUyjI+BOxVfrCa+qqm8NVkhg4OpvjDAwB+zvXqYSfpsyPmpO++vPIfCBqe
MoKJtrvER5Ab7vHYz7JJI4d3PnFBqNDNWbLecujq0oqad7km9yIZRDEUdCqFmdeB
1SfjX8Wj1Wd9bEfZSaG44yiw+ZYGGXf8QxGla3TmlMojil6PRRj26QX1P53OfCto
ErGLmYchPZ/DQzTNjLNTzAG+e+8duj5+D2ZcEOyn/L9uIWaRV868Q63dxmi8mzhd
4gfJqIwLyIbjuJrJuJmompySLpKaEaOOp0gqo+6YSkbuevZFIwcyVM6LcKKzIC/D
cJb1TEwgYyMDdiod41dMbqYQJU446Wn6w6Omm5XSe9PMZidQqT6D8BCywsuB9iHI
pG1ZR9Q4K9Xh8gpIiGZgzhOj1sWGFmy4hqX2+eiKmW4Gz1XH0xpg6DL5LjWdUmVT
s6wNEIA5gCUsg2+6qwKpgwutrzvY3cdM3yIU6GTgITsuW8R0p6UmsRoei8S3H5c7
rzhayZM43XlsfmwumcDeq32mTbI2Ods2lwJQNhUTGPW9re+LKq6Ad113KyZ8iggQ
k5ggR2QrAeuLumIPKVowVtPdkJ1PXmE57CPLAl/Td+ElZ+OsRcabA3GfpnTMYtnz
cDu1qKdUb4Me7v3GPnruLM/u1u+RcVbF+YktLo5bIGQv9ZZeeFEl1Fmy0E+PT6Su
W2kv3H72qMFXZgtDkCHGReUz1aN3mU3EdaZkeOhRN5DmWcSsr9doNyEWPlAl4oCW
FOkojMV5tuv1gh4FmMSjKd6Kn6IR4KBNStJKcnvYoiJ8WIll4YXPl4hq84UbqUdo
MeV5zZodQ2d5Cf3+TuUkew0zFxAxnRpd1aj6ScsS2xpJw56QjL/a7SN3VqDypBOo
BmNhCF8F33/6aFbVhoEXark8UEyViwgl7qOvIBS4vRZDgVmvP9JSvtIr2YMDk05y
ueB60Pf31JEZ2V9BV17t5xKHhWt54ULAawMUd+Exskr/P25iaGMZrvYOrW8g2faQ
0zA7SEQ5RouzdB5AqKQAV5b/ceW9ra/d6u4IOYMOB6VeZuARICYTbvlq4ZsyoEXV
V8Wvwvc0oFR9TxLD4a+w1oN3KiZLRso4MhFL+KGV4JuK2YkcQHGTJeMq/GmO/aNY
F7w5GpiylmqC0ay+ai1W3J74uMJwteO45p6HCmGLVjjMcS39eLa80wFqiaEpx83X
QnW08y4+rY0OX3avArFJCTGJzE1sJW86gxvltdx4hDqLWp1BYYc+7Yw3TkEfF/x8
RvrUHOoTfGtiywcW5e2+BRHegBM0y6WQG0NgDUmJ5ZrXQC6ikO4WWE0Dbju6iiS4
0FXyZs2wnSIFGSOYEDr/O5c/9nncalcNq0qUknJNKf05F4Ehzu16SxhvNeLtS4Cw
AvpLSO5UbwM507UrciQHQ6uqCQy4LrcEUzrGVdHH20VUkRa6U5IjgmPIs9qS4UBG
uB6J7jXjADk/LPmHZelBH95hKVogrUZeMP2pYzaqI0opUU5BQgL+4X16BNs3kYvK
/obQfVD+TBtlikoSPuRdwoP09G7zOj5NrFps1aNOl4vyYlSj+lIO5T36D/8KWnw8
ShT3R5TBQMniKnZNzxZszrmao+WyC4vCbjVTz7r3AAs5CU6QGDuMNy3/eFWmxVsf
oZQYYbxNwgbbnR1t5tw9AKaytrXVuqjUPZPJNcLKNjopz89KT4A2IO88qN58NP/A
lVIDuqmJWY3QAFfH4N/X6zQBgxSEr1+Q+AElFgkkh28stf9xDqdpIhUMNGzpSUJf
NY7bt/89yAujIK7ZHXh827KlQ/SfPU5jelINm91/L4h1hYy2nx9vpcEV1vJ2qGt4
rHxabf6/ESx1JhlpmZW1tG3tLUf8q2LJC65t9hOqlnAyG9TNGFFH7dpRUo1kgXMm
nWHfIh1ZeR6lkGGRdFKSnx0k1zwIQeZcokCIKctYaOWABtPuiGrr+kSq1ZqhU40Y
svmcUHyeZQlZ1px9TsaN5SfGQuMAl9YKY0a4QTmTyz+Il1l3Nx6RHWNo7jwISlcV
VDs9rGCh31re2aWSnEmIn6sk+ilTCmbxBKDEMwqsRvasOumoLarCjCaCr2vC91K2
ZIHl7DwgYMil6ct7sj67izzT1hAW47Ihfs8R8GVebCWrvklzuCRtKGClnWZdSke1
6Je6wz/VHWFJE/rFHq2inrgUdNFRO94ohU3vu3UoIPYxtci0fbF0c/Yks6XaTihM
tIV0ss1ot8fZhHMJwiK7zfZwKy2a1k8gYS22JtvGl43xSZAS6LkXskreO3pZKGwc
7bL/OGmN+vlowWBz/2cO/Zn0fYahcO8fFrTbGOR2q/qXz0iDgQN8bfPhnGgI/4nj
SO19klwIj7qh/kH1stiE2DkIuGldo5FZNjPM/coQwPIlsGon9PCiIyIobRCnl2Ie
XIjuQ6YSECnJErmx6+3aJvfHh6+CDlP6K8ho+25vK21XgfMbj47DY3KY834sdtpk
ms4iDKrxVYCsYEs8F2PbGDXQuKs156XnM27uIALHgj4bPOw1DUuaQUXnvV2TiOoT
tSdiQmMcJAmlJWNsCBy2FK0tdWCyXQKLlfPbsPY+ML2wRFb0OV4eRxBIj5f0Nslr
WCIDaf2LcxkHGjBE51b78NIuV6hTXpePlFj0IhNSaKPwz4NkNCqa7+ecKZCLSfPQ
3PR/UQnbIAx3gPqvM9cZKhPJ9YV2S5OlvBTlY/xv4qS1yiM8XvsThBurlcq+0Woe
y823IFzxhuoy89QoksZYjnCY/kgrgSU9esIo/gJT4s8j1Zl/Z+wIH7FIMGt3XQMB
6UZ4djW2s8UTeNkAdVszyGTVL05WEBpfKl7siysJIx/BPSGQ4jG+SvFvFdFpc/X6
tLuCNADOozBrbZIrLd9XHHnjHh+KYjbqjQCikgBog+TrXLQmLo2GT1sSXx3+QcpN
Gh+H/Fsb4qJuiaytuI41WQuFh5N5NY+ez0ss2Pq2zYPIa7bEJ2Xhp5/JngxH7sEW
EzwQBPTLh06j9XtT8HrCvzGNR5XZVOTnuYLuKurI95ai2mp4mdMYkOnuovxpni7G
J/xoz9YYElKXjLRbuoHHcPU9t5R1jYNiWGyGnD97N9Zoqf/rq8kE9jRCCuQvMzJb
FDTf0BjcnTFzWK8xmns93rXZitqmOVY9++XPRYHEsfOpGFQGp7ezuaGKZ/VRLxXd
2JDGG1ghzg3gMa2kDXEApuL6fFiISjqj5agi7qiBNoiCRES0dFf7ZDp3DahTgKSA
vk85lyKvd41Dmi4MT6HbjeWer5pMYCCNT1QuXLgTlZvc7htLEoRjGTgIMUhJOlcp
gKUHGs1srl9Z3DwxZxfy0VWl3E7mr2J6V0qxSU7tM6l2WRf0ebwNkBKW0Xb6xcns
9f/+v0/i+FWMLJxQ5QTtGbknx9zS3kDTZ4sRGw/nxnUHQbT8y9rShAurrV22zr+U
AKEOTGTG0t5FKUm/zuYcD+pA0UX/r1B3N4gGrjQzgoZgY1Or2McRZ7vige/NJt5A
ITAdyHWOno0XskvAscvzPPimv94vMiTgjo74Y1ZU7p079Wx+fPe9PdZFNyPcTJfS
V4baWKdzufvSQKJ+tuY83PZtwS8zMYw5rORywMmAAKM+0vuWMEBDRG/Itbr4OAwJ
jTHQg8oJQNYgKXpLvXBSxwpuY+RtUMUD6lqXMGYWwASB83pxryg8MB9eKEyJVvTO
gniu3IOD5r1MbQZh0KMgZgHDdJRcXT+r7je8Ce2cpQ7IqIH1gxcFGqi18JDv6rXR
bjMPXbARU3J9AIMmIJp9dno5iE12yQTktobRc8U2NtWoQttBF3Fj3EUa2ZDdENtu
9HgiLHNxL9htv+5sN7uzHx0JIyjnCRP5E4jAw4VOx1MZr+yfXix0rtqpmTw6Up0x
r7f6gztQaoq7V0v7duCgKK6UCOvWvxlBgUUlSxe6pRstt6LLqeR7ZigUR9wk7rnJ
rVctHl2r5idGvZdDFbB3f10oPWkzfklWna60uV7SINxLrkoN+QBblPAOLlX9UAAx
31oWjBXaWkMbO1DM7em9ZiNsJiepwY6gsdXYYzxm6lWcr4EuB2XCJMQ65fUd/zJ5
7IvTZ21qywJOR8hVeouE3YUhXNmODWUhO8XkaNPLeZyXlEbwprk4Qg9YgAbFpRCd
mgBB+h3dy6AuOOP90E1ZQn2V7r26m14xtmcQk/F927ZP5rPdc5SpUIpL9AOpRIcT
B6Kc36WC5/N/D65j3GKCyviatvR0eRfNL1tRJQ50pTH8gK4YJCD5MWGmsLtxETLU
PwNuhz9I+KqwLg/qYZ05TglU/7lT53L7R7yAz2kvOSOkCdb6VeJD/7d+bIQTBYR8
JIwyXobEiEWciB0gbHwqa4oJKreyI0kjdwRMfCM4d6yBxqVSEH//lv5Zw/Se9dta
EqoTAtoQ1d9B5JFsuO055tVpa1B9N38yqzGQVVwJUaQHt6G3lVWZAqssgpx/eVHP
24FT2glmnSX8U1pJhr1aaoNaDFHUBVJOcLiU0S3IvIykYHAAzyleUXfBcFPfk0Yj
GbEO3Sca43q+dbG5CRk2LJHtfeIC41SNw1emF7+704nbFeTmhyMPSSNYc9/Bfd1w
vEc+hoyr9FJVVv+9WoduzR3cAMsZfsVVhlqnfTl5dG52lqCTV8cAvUyCiulO0r5m
8atSMwFe8tspIlQzGO9HC3eIzpAj1lvttek7ZA1XAD9bxCXm1RfrZGPW9tluRxPc
y2lgOQivZhm7PXfXaKFUJ9T5cHSntFZiT8NLyNogA6AIuak7acqNk9L5wE7vswrd
ani3AJXNKbqtOyNnggjxykOBFjdoCQbBYOlriu5EuUtCf+KbCGNa3+Ah0zjQgpKb
/GC1w2B34dq8sxAbvZGkDghavpD6x9ymTkKtsj+EQkz/Dt03xcRtAxzbNFh9kASZ
QHlZZajU99XFZG2Cm4WG46oe74DrhgZ/NzzTZhuvlO5Qa6rBWvHebEPPBkx+wna+
x2vge8OCejSWMKcFJQRUcBIYOnmgd3V5UTVAKDJVhMJtBi3YviTuCxEpp3knrtIH
p0XPeAwGibIoWL8CPON/D1lsMJbhc2nPKmNpJZR/HWHpInZcn20diwxtTlYUoxIZ
7hAxDKCywdpc2oyKuVETPn7ERNOrEVpReIuvWO+aW5asbQHCxlaBHtzYASl17Upz
4v9TjznUbUO6buKu5pHImKb0dk9J4vQPnI0VCc/BNfmUZbVFsKn9oDkP3IDHnwIg
3vcnQeSNRuogCM15sDr5jG85iMZmLqlqg/Dm0UH7uas55h+aotL5DbCF3/vhQBuE
dr8G/XQqs+anhB6NAdLO/veQlSCa0SNPGmX4Xk1cT64P2EUcKWSKpFlgx/PcoAJZ
IUv7XE3LwNBJ8us1kotq/t01pfK0MoXlzZ7Rsrz+UEZYX1+u+O5jY/08pJfV+GAe
Xz30Uktqa+pDvbuQcCEsYkPWIkM08RXIkOlLHMDcvqyMacagSDgZW1WoJt+sY8Zc
J3VmyVu0OrE57e+UYR8srgcmzzcdBOWJZeva9YWOPOtWF7LO6Hdi28elfuhksHUi
0i2UUz+ZaHkVZT3ybbWnUp27CuC/5lTmw9Q41ufjMI1r4x3l+1oWjU8YAxcD1deH
de8tgQ87HYzRLGZBle8oWIR7zoBGZuJYQaUpRb8U/MfCQ2Vd+k3yXxuC38q3XocL
my3flSINBCBhlRA+XHHPviFL4g5tEN/KANhEIPUsnnH8nZ5pY2gfx9Eo+YrjrgxP
tnNBqMZElo+qhEChHr6wpYv8jXFAKMPOeH8UIVsgQHAkJbTd0r1+dY26Xwax+wbh
a0REi2cX+dJqOkY5ORMQ3Z0mBZaI7t5QKdZyr7RukCUeyhXePvhT9GjhkipMlbGf
fvBJN7PPVrZp0wigopBQ/lOAImUhKwSrkq/TxzX7lXVli9qO7KWlMzhakOHMIsiX
6C9dEchf6PJlqePM5GokJbXbqzuc4ofAgBt85Z9jFh59J73ViGx61uV9LdKWUpkj
kYqhdQ6yGthl3kHLkwHRFHGDkrCZErRnwhq62XP2KMxVscpi8BV7dn4S1YYJfFkY
BHzt4w/bOzKhCp7jLcLYRkETuzGwNGm9NAc/WaGNJVlCroLFkVnPhNSMpBzM9Itg
YGFwewdejEVArDkgrD/4qB/81aRnLlYAXRBipVOqYj2NldsIMAla5czUdlL3MGX4
FwWIHRhvOZqpJcqWOHz31CJdzhy2vZ5wNsK+O15IfIiLnxcXVkptJ60bCCOQ46jb
dZfo+mhZxui6HcL7NHF0hd2R9o5J+tczzrS0gIE9QrzW95uS32+/PvsX+1dDUzhq
jqwRrFQPjPvF2VHsUU384Lq/XXPTGvtgE6BNkUb+1yoM+ouYG9WLy3XsuYPwcEAG
4BjpY0jKL1UkLO0NV6p4P0c9wY4sBLE9P5bS7uZ0Jg0Nls7KKBKQu+Wy3B5Ys3Fr
UQPix6Rt0yno/1OgQM2jnKOMgSCpXfMs6IgPVHL8s38XSMQczqzRAdX3ziQxDIuF
lNoI289vY3tzVaC2QnT4QyLifHZQxa8FxqsHjMka3GpYBoB/s0Vq2guNo6MV4TJ9
roswHdtyfWCZYFI6qNa0t98jMR3hsK32O9yqJ/wAADVhtKnZ3zCqbU9vK2R+upth
ojhryiE1eZrDKxkUklQm5Du6kug6mhqGgclY4cpJyYSy3QpGO8CEJv0a6HtOxUWi
WGX7dcBs6ojM2yk3Gk47muTKXFDsPTuNH9xWA7Ec3QZz1+vXBbpg51I7TgcX3iIU
PY867K20g7pfRsp83xA0bChWMMWrHGSXh+8IS/k0+AUK0W+b5zXYShlssa8puOaO
sUzgxlWxtk6xjb0gsDm1iJ9DtFSYnBxAjLyM6GMFD9N8CdGHFiWcVTV4QZvsopbz
Z8piL51ARbaOP0BMKRuB8De7qzNhmT4XrAB0UGI07FfgXZkZRplKwuYejtNy+WSN
cDCVOZ9ByA25Gt/q4wmr7SF+rVNY9NPIarsoRJtf4wbp4qIK6UsjceyBOMIEk0F2
miQXZxKa+gOt9ZbJQ0BMuPn9KeOxCemoj7H3M5n71ewo4/pAZtHBmnmSwk4oJ137
OS269pHdDhH6745IJHigICBEKmLztJ15YWtnyuLFDhIAVS5+9++3REl7UmXsiTds
DUnqjXJ8OaMbGe9WvQCu/QstPj90esj9xOKSWvSZZgW5FFb1i3ZTTO9VO1N3UgSm
Rwuwd/vV24FoaIIAZzgtootEgnAQPVMhI37sZ56lYW1VEqHyvR2pOwQZbQ8wtlmV
4pEI0k0B2fOcdVykStC32IgyPc1JfGsghpYUUvJZc3rzZRLF4Vg1oGPsC+/XXixF
0caBdJcV6gGgTzDNXO8xY/TrNvKQYei6rOph16LU2SWApCFt0/Yy9iobl5nn0+Pq
69XCSdPOlOZ9194zUFOpv9gQZ435C+XCJZWLWiGIPkfBfjmG5a5IwoTah+YX1O6W
/K1EH0fUE9WCHnIpZWHfQ3Tihxtic1sTLwS80N1WA3FKoPo4YWY+f2iDDhr+hA2n
KA16G0l+2a51EUrnRFxcYDBW/et31ulOKp3m3X29RA1g/uSzXrItE0q7rmyaIsE0
+OrIzVh6HNTri3uqj9Lxllpyo48ElgLkUTvxcF0uZ1KWolWJoHxbp5DarLesyt+3
27st4cxqtav7xxf33HFn5wPHBQ/dVSyAS2GTiW81E4e6UEQbyhymtcmBEpG1hxG+
Ts5jKdTm78fBddY3065+gj67nyBra9wW/JvprOUFYDSAfttBd9DAGzQJjGuN1HWH
tr2eSQSxwNVtDyt1xSCeWSfIHG3zTAtQ2HFmdzaP5zeXPpnlIx96tb1hRMLmmpKl
Y8DQI5JDE0A8S30QHbPW4QBg8m7Nx4LDEm8cdCqIKReYw7/YEj0hxpuw0bX//Baj
NTqFG2TojEko4RUq7K/4YVbBgVIXv8ijggwpH1yJRb5TIZt/BEVkkfYomwnQYn9G
03hAs8txG3l7TGc7OPbNONoW77Q/6mbfp7YEvJQJgJSkv9wMmPJ6h1tUkcABpkz2
KnrKI43EIWtVlHu5TgCBboGGvZV2bJUVeLzDSwKbYYb976NoyGmQMeZ6+hDjrcxD
yvxGPyOhq6tcXzU6bT1dH1+i9Kv4cljS9Tj2VTe+Q4CvG2loA+m002vfYF3iqn9R
lC45Qv88Z6ohFnzctv79g1cVNLPQUaqhDW400/+gox3vZzKnWTPNbiMnNKRrv5K7
3p54jbmb2Ip8uAU7RoKOltpbqWmGtMy3bX1lcgkiQAV/RpRfb+4ApZDC8T1H7kn1
dmiR6dQla0aUz3loCWokiecnj4WJkGdUODBHG/5hYW0tUbF3JW9rn7EUSSF4fkZA
r2TT4UCPZrYuIRd/VPzCMoG+2KNAhZUAfpYPfvHLUVM2BUyK21jSdSFCz1HbWhlJ
/UGBu7oNXcF2+ZvcPETuycuzHnAM11D76Qrr3/wQzZd5NVIaqTpwk4yA3z9u9vKX
k2sf3datZ4WT86byZNjh+4t3qlzul/CZfexx1GEuxn+w69+oHub+MgQv8E1xubfO
g6+bjECGCJQU7NBy1+ukAg3SWqh7j+XQAFC5IRXEW4EcbbzTYTUpgaMfyfpaPWp2
oCI+8u1uS8mFE7fzlrr+lDxbL/N1fA48lImqTxrucCk5gYbWq4bmecOSZ7riwXbP
+1EGmQSmgEeoDfqXnX/e0rlxDgGAVTo5x6sBRUBfdhAgoEUJhyWw6sB+NH/s3Fof
FEerAt/raNqhqwNrnQ8p1QulhTfGbc1f4P2n7x6qbWIgqmiKY0J/GFZH2cIII2Ky
XGr/kfHgOp0hq6dvTdFwtBN+1QiySbX+9gogvW/2VWtWvqyevcGIeQgLF1/NegyZ
ZVxE6KbdClzJ5Krms2/5yZVOLfp5uFcw4FdMF3DVeD2N2diV6lELK7sYKrnFW5bb
L0IfMNvB/P76flvzCma0fNfahldNR6DUknVT+fotzirEqcAROTdfKEopn8Lna8RX
oS+BIBSR7htHo9XYQgL1uEPK465Q3l9G6wSe98xwtCPLmPOxFUKAtQpp0s4Wq8Dk
wyuZwaE3CTKlS+TvKdH+pU6K+bzh2mZrZkoFq1nFvZ6YCxy4t8Dm3lPDpSEsJvU8
g4WuLLb25NtM7a7mpX4tfEuTr0k05XqwRoNe9aIouP1zQ1ZsB4ctMyzljoNAmNFw
6DGDu6+XQAWw9foJNJ7N6HkvjFpf3YA20mNVfJ2p2zojDNCuponn9FOxsjTi9wpS
IFDqIVCjUjwWx+B5aVPo0Y1PROvrWs8hrkDrkTl0ihapcxmOBAzHJbzVydwo9vhy
bAMWlPXPW0pLnwfRcq3wjjhGrMwwYYFgn1JwlY7DiFQSMbba/+DPXF6rfvF6PxUF
ATq/61PIKfmYY3N3oAHx6KwDTedL6QXkuXlGq9dO19JWKUBli2PKF145KALuJEnG
JvEL4gS0HF6hpk58kMkJpv9UR2TFJ98UxgLwrszSwDf9Oj9Y/O7l0fe3bpSWGwym
XtZTRQPnV92eoMEObMjJM47+EVeHgDeyEq+g4X7/lll4XMXKqHfaOJI2teNT59Rk
8Nasch/JSe4YP7ECAfgicqLwHLdGXruGQr+4Sfdqoc04drKNDh/is7TtX/dklcgM
W/eML1x9qro30mN2YyI6W1EtzWG+0HHar0j/YpExk/vDy7EUvQi0QCHIq2hBmsNp
DnemEhtMvv67BwIC0wuIl6geAXlgmKdeKRoAQ8Dae0uDCiWw9mW889H02VKKEXmN
j06Xz7Ykk0yLfkPhjCnAW4AFD0SQVp+4y91s0pWju2k+dMFejJjd+t856W3i8bdO
aHAxytqmmdAKK+s//TPrqTo3Hs5B8y+QuMv9PeJQEnfgCXsr6buJUXWLOgLp26Ha
I29n6flNG2w77tSeZnp+p9fem837PoP//Yp+q9OJ6VvsgCb7kbWOkVpOZSN8DJ1J
EHL6QZV6b4CV3F9sODKtMQ+G4cyi98jNChvXmy4gyc9g7jb6WVQ6EOm8FTphzU4C
mXpj4ICLlb6D6frzvVKV6NfncAtanwmK65f8PMKd1G0GXCfCEuG09UIH1lKdkxbL
rsSmfSjKFEZIhnvzIMKrJ+6emu7ONgjoOVfVjDjdUsu9Lg9wRnfX/4Edg9q02Y+M
lCh9SOPxzBz2EVaN40PKE86P6EgAIAHrKuX8EXR7I1Z0HsHH1Y1hVkYRDUDn5PoV
5xEj3PC7hC4Q1k9VbKglOoATquiA7lChdpjK1pHhNU0iH+X1r/fImXjtJiZvbaRE
iaUUgoAB3mJ3bNniXG3atxV4UQOF3F8QJu75a43ASkCGcc6yjBLrldQ5ucpoy4C6
hoS7wC/fIHa4Cj2UB3CXTF4JyFZtvmtFNHWgb6eXNcOlb2knJ0LuVZHAao/E3hZ8
uE6nR/9LkJ5+svsSsuX1mCleb8NrkzEb0t/lRk5j5kWUhONDYS+YpA719N00CWAu
KkVp2Hi9aXsOvSZonXwbSzfAnosPdFz9Tq/3Z61fPl2TdA8MDWV9wVX3qOtWOStw
2vE/lRUmwWDR+xw00j9jU6pCsksFYbSGWBzXEDGJKbWQBwiC7oYLIhQUaFG2jRrj
gYZ37wWMGgkmgxrjXkxp2QuL4mL1OFmtDZhssCWnRUlcVa0JIh9ewCvQTPvmO4bm
1HtshkzgZRwwkGW4HBgdojqFTIDSAQEZYQZsLvslzfFLiIA1/SvKQtHp8NldvtC7
gD5LcvsgYHEE7GZv4SNOh1G80DPyYCxv3/HujAoMmaY9BDPEigwkrNOdG2e8PHZD
LoG5/Izr+thllfuxhxSregWoVJDtf8FcVuQOyWMFbiGYsDsg76tQv0ZmDc5yDILt
k3nc7UhvdhvftZT2h0ILV6jPcZ+hpOrb8J1pFtiMsvs3v21OrChd1FOh8QEnep1W
nj0xRxZSpCw278znekdzbofMeTkL34yjSx3LQ1d2M1iixUUEc8RG3ZY1+vzinw4t
kp7hEqX0CimDje2EVqgQODitnXzJMBs1bGhKUIUOWVSdsnQptkRBMjao0DSuwk39
3SEAOKtn6aaqc9GekERvz84Mw7vhGtYDCiu1K+/oH8FmwXOmcp3/IPQ2WD0ER3dP
SVWLYPFS6g5PAvudvAD7QSasG0UzPY/NTJpygA9rRnB1k9HlusaYjw1XF4KS3Bpm
O7QvstPZKH2NXZ+8z4qvXtqc3aToKpv94PLleW1dM2DRU3zX9CUUyyWZLxZYqpzR
VboHB9U2Qwgm756Ke2LBWw2nA2r+DW2PzNakOtX72IL4EjGArONYeIFR4k5v4LJG
FKeRDnvvHzWorIMgt+atgew+xvzJya8Ok2UM/H0cX8I2DAfPcyUEU4C5SDYSqagm
vKJVtanjqx8HbfKD+DPihifoNtIHuz/xaK0J1iV0dahMxdIRcKx0hirdCiiuHyfa
lUfxvJ6cWly9FOYGvDQJQF2eG2rkEW3DCCdENrjRg6GYeGKQ31lOywlavFPJHerP
Aee9Jvyw4UTpWOLu+JV2yrux98r8l/oAc5hIKs3tsmV1ZVg5+vROrYkYeD5XdbzX
mZBF37D0yfL1xw29DhnatC1/6A418D34I4KzOvi+niiVZPQPRAr9rHhjEMPkW0Fq
ziLhwzBigTzjKhSDY6JlKoSkvJ8fLihGRXszDkGXHQLI8elOwj/ecBoQrD18NzZG
SscOUoq7yzxPHTJFMfCb/QE/O7avCjUy7D//Ixi9yfHb+c9soxloEzY67KsBleAd
l9e4QuD/hBQwdEiP5NOFsHbxYGGMktY7N3JD+1b+772oI1Jj9yotuGnfPVa+ZuP4
fj5iV7L8O6N8fECLkhqCcRepBHaA1ZVnBFaXnXi2VLWjIIIRPhTAYqymacAX2pYx
uG18d7vv59AIWfTIeOLJRb9KsaQ7PRSMbOGargf+xpZ6qQl/beGM2jvpt06aKBnH
bg9M8qPn9YjZyGNluH0VNqbWIDL24++m7csLTdShbPqKk8SemMI5KBoBckf1HIRS
jJq4LJ7RUr5ZXlrJeOISjBUuUrzexApgG9HLhEQEdhX4r2REwBUUnP2HdnfRaQ8q
7h765+MLmLB0DHlbf7Z05WPHMq2+V/CZ5GI/K+egym4UXxrruqBv+97ETk7AnvGs
M7vgItKMMnKWqKK3NMQd9CPSfvCX2SBJ78rc3XmeVKODmDxV4etJHjazeA39LcS2
b4jF2yCfhXS/Q/GpRWSiGlVsgaEeeaozIN7qEFbaprzjj9rACZDy9dKhpOQC785H
JtOTo//xUZg3hqW+lOVPK71jDej4Pzm0azq4yQX6Q9QzshrEiPFKrsuz+DCJBgKE
SfovM8NG25XLIKPSo14dtLCMFpAPkpivMXCdYTv24SRL5DRersSQHQaOnM6mbxF3
bqO1majlBCRV0j6r5CcFn2AhnFeBzE6C1C6/eXfB3R1/JgZIMZppCveFpj/z7N3K
xCL5DvhSIWqU1xclQdiLbWpna6KhDUMlX/rLh6MiiPe1S50weN73TgoQm52n+pud
bD3vADDS5HeGuMFMCr6CKSOA8MQ2983nFiK8P1R5CVDlpIJOXO75MW1tX9haI0RK
2sVMis3UPbb/Vq7d2/jYktGjWlLYikVHeSEOpYBOSpz6qALIO+BbobBb2m+Bo33c
yJeg8Z5gAWNNiMe2JFdD5zUEd6hltwKqSIUQsthBVFjvv3afobGIqkX1zC+Pn0hZ
efpWl6waQOJErHSHo15igLF5MKUhE9VPgid4PorJJoj3HXcsArGcN4oc7Bn5CS9m
AQMwbgf9CSitfrjYRAD33PJjpm7Xp9jww0/aGK0dlNQpG8NNTAGI9Pf2nPJ5c0bc
fg0L5PP6GOUojqrZsSlA6Qg5ouhT6yrd8CKa3PrcimAMqYKsRqocwvzuO6sePMBj
dpil1k4cy7A7n78kfW2ZSUIEXErWuK5plI0E5xOXHx98gAk3TObEqa0GP9OI2UGs
gL/mOACir5YIgPMbOFf3oMbnWWQ8SSaJlwvLvkQDb+xp6YypA2ZyHJfowh0XitTv
P3cp6+aV/AEotUFTV0BENKY3gBXIbIhdqx3gso5lk5p3DfGN20BcitmSH33llGBA
GOdgZMoka5FwamALlAHahrbOibYxYkvD5becC7DWCXitdeXnaOBthf6CrorqeTnR
gi/7dlLWC8BdgR7+WcvHpGuBbEIFGGpTnPO1cbN9+mFlqxExJuqbqlrynlj2CliC
gihmhESDsY1SFYoe8ndviEzLH2YrvELV1y98ZKTWP5HCwevcJBAjWkANEU913UIL
siq/9d3E5vy6ABPi9Iekfwm+2Qwb13jEeBeLxRo91wc1I4JKYGkQOs6VbP4h6rJ/
0qc/cw/mxbGoytfa/eX/wZMCeIb+TjmDkcH6dmKIYh34pe3ZDrtyKtnuXPh58+Vm
9cXwwyl8Yriu0/tbAWWCGM9kdPqZzqBLeF6b0MJvy6YPtb/YoM8pNzj6PvQIuw9r
CxXl01jr0Qr1JeuN4Gr3u6QWJgMT5fxKMDfoxUhwTN5LQ/wODBGfXnmaVSjvSs9O
HxrNiNBknm/wMPlh4fY7GaVoMqOHCsMaq2ujy3fg+R5K1NRHLbp7hE3wxhnX7XzD
OkkAW8CUEaq6XlkjuzMvEsPNHAd7seE/T09aTdE+OH2LOoaWS6id3mkehy9F1ZKq
lA2/YShMcQU9NYCQy8gy6V3xaahcDDbfXLjo2JgWPY0q1/eQR37paEB4cfDIw97W
XtlV/9COMk+Qw/VLRL8K0R22zJtpM6iNf4zUBe7ssZX+jjiWhCApmS7N+3drtmkP
GA3FNaN4TqvLaqrjPh4nlUh4nNUphgNdU6c6ZzZ9+3KwR5mKJsFRAHyONVPLbGPE
5ODwBfSEE4e1LDDpSKuZXG7CWaQkXNFPoPe1zLJ8hpJU0SxYrzw/GYU2eq2ksv0S
34WjsSsXF4g0rgQy5fCP1rv8zRgttNsB4BBcUjW7YrCtlUq/IxThPS+mgweYpTzB
RIJP41eiqmtjQWrgqt7HbSRPdh++PHHBCCZyp5zQ21+RZn0W/fIB5OTgwrKdio+D
HblaEtkhD6KH2/3zSFxP61SvZeVOG/zoitjrgijUlw8dagzxjZnoRh5L95exDNWz
2ZShJxhD5MU5ejgEPGokeC6xipb7XFBHuxAHfZ9xYxYmtckkJX3IELPEdplN+Kb6
pJaj2Q94xQNygGD2PZLvH21JW+qbTr2gsn7nDBB63LtC0//54dQkWH6zfrSFlzEl
ihodCk07OIJsLwlniYXvxDWpzub8gkLMimRp4LfhNgpxaboSplZuRulBxGBDgWW0
svu/rfeDhqDJRVLYaijyccvJexFMUrtjZIm8A5LhHKYhrTzhRviSqiSZJrf/k333
Yux2ZJ2ZP5JQ1s3YBBkCQk+NbeoO+k1fgrjuwd9jQwdT/1IzaTPKH/ls/L3X1hS1
9Db4eMlkjumbI1+5yn3SK9UfzLb4wH3yPjF3cE0uvh3ChY8HigPRxsX/IhhHuEtq
809EU36E0Mf+DZfQtWoda4TzwLpBA9LDfN+DSL4Fy8Hp0DpCsciK1FamUF8obJQx
wlYkgx+i6nukSOCM2JTj54VVw/8NxWAINEQTZpWOwFrl5NdYhDZjCn+0ZU2tWDbG
lyySyYiXYfUrRewJi/oVUNC3/NmKOwQ19elROUM4z5zfRu13n8qbLBzNC3/Cjv2h
bw/ZCw2vWBEGSzDUyj8+SAWLwaDn+bvFnxSt0AGKwz6KENDio0loDXoqNMwdpvT+
0hIIB+advAF30nKJT91jTS+0gAIg5YGxwIHvRz+LEqv1gGps6WpnX7eY7W5UkGXw
Y7sYo7rdichT8faVY58GaLUSDToJYU2G4atxviwpU/QRFRcdLJqWMveyqzvC8Lb4
DP0MZvReheBAH3F8wzsqLpnWRoSL/gjevRwiGMCp1g2l92UpDAcONBwt8SpfAAVo
0AuTeH8m+hLkuNaqPbKdUcFKTfhieD7LVE7MnwR3Wyg239RP4vb74QIYgfpWP3kF
kdKI8FhaB4GT6/RUXVTyEQXHl9yWG77iatloYS91zjk1lIuNt1Dt7kNKBrek7pb7
7En8dX3qMblkSlRXWJ7fKPPKc3hqUH6T6k/tQwBt+V3+5tQe4YPRviVvdyzBO3gG
NdM+wo9+vRG+DZBOaxv97jsXj2JF6yoelD82b1mfvw0Y2/foACQQ52AdybmabDaf
2N+fqfNpdprHZrT+MSUBQ9fm1L72u+EcMDEshkkUb7eUCaQ3CRYtzQ+zaM26lAK1
HrnOJ7OBRfKsphzukTF3R4XJsNr+rqUYs577yUEjfuclTEaMEr/ItZJhkZoRl9Iv
NF7Re6niJ2AOAR/Vzd356uqnvOSKAfDSTMo/ufHKBgpUkO1hy8xiwycoJ6etIIKz
2fY271ieCcvH6t/1NVgmTT9QGnwOBLQixoLe9e8v1F6GHn93unQqbd1+eoMbQ2c2
W8yTGQOUfGuklNmJX8/u6mDQAXn4n8L2FRS1FREmgp/tJVEo8HvAnwUULwKhQD6N
DKe2WnpLmo3rHeO5VbzMgw57AKHHq/KvqrWrJVtQXPPtHWYJYjM1RLqa23g+sxlQ
+93KksAswXX/yoNxJ6J0gZ7/8aWHUciM7DHesM00Ad0T7Mu4KxhLkQwL2DzQqUgg
LDUtKSYObuNEQA55xfuqgYng1vUQ+jJvlS11r2jjTwybn8PJhNjXj9ciTYhB58uZ
/dsPE9Yksrk3EStn1dKiEvoNeFpVZsKyGvynTnIPlivONHMsovRK9ygrPiuDBUdW
J0xb+ufx5EsDfelbDT64cK8w0xuI3LK5FdiOS96KOZdvZ2ZmihTjefOOKUA5IZ5h
+lQJyYO7oy8IFlZMKB9z29M8A9fdrZyWtindFjfskA9Ux1Tw+8fBw7V7u2y5diCz
ZEYVi8cXxBkUoNQvDfxf+vsY21ZlJfV+uAt5FEaLHQoHsC7LYM37qVir0mYeCKqQ
z2TBV3BlTbv42HUmiWY8RJQ4SSK1HmkuKKPgkhuX6o5fvly/GSoR5nuyvpcecLDM
sVzyeEsS6FPHvoMNcWJuoclqJdWrpv6PIKzBVHbCgNz6q48JC8pChklENkB5PrEy
gBkBVbylbEeFumpma3FUuB7rSjKXTRa/nASFjjInWW+P1+gLVRLjQRL59fubKz6o
JnwWx0tK0/OrvHujgcOsCbk+KhP784PMCNo+pNeiNJpok+IbMBPW23yA6S4hEo4I
6W/FJvCG94Dd20w5/Xexg1KlsKfoGq73x6P6tQaYS9SiiS0V3rZEGGBD714vcO/a
34PlT55cPaBjvJE6KtbKXyl0JEh0qtmDxJosmipGvUD+0qpaEZunZ3l+KA96+m7L
QjgHCGTOsKxUdec5FoENvOqnZ8X+8vh0X1mLKpE8Fm+P0V62yWs4G2wFv2mej6uG
bkWVSuN8mrOQKKX6h/GzKYhHzRWtlOMQZ5xgwbVOEpa2Kvh2SEgaa1BRorIn12vx
Hr1wbzCbq6RnY0MfSxYybe+GdV969qnLEG05ekeeH7nlM5LgzCmQtOQXzkHUCffC
aqplIgKqzTRVBWv6i0w3x9tg4VHgrGPIQLhKlNZZTRW2ctIirk99J/GH0/A0ymp3
+RjqBp27Mq4InG/PBuJ40ZEpPE84Nn5SRRjZRwFrHR7DWKW9e+TbCjjEaRTf0Z4v
zURO5AChEhF6HYTa4lXsEXFvHT4xiNyPd9YZlu4rQK4JBXoOkkxV/NJONHNWpVRR
Gxi6CHPOkdycgkytSj0ET6XG7uY5WBGyOg2jN/+3sc8/cLfJABXzMLYQ34L2OxjZ
iQQ034nJBBdIwg0NiHM8YfHV7SVK62oN0WQKwMP0PKSUbIg9Qfl1IID62z1JghAy
TFxOVoOAKy9Cl+EnLEq+d/I2TEhvw+1Y3zEoa80jtR7AUhkRtamf48tdXmYUT53T
qPiXHMPCiRHl/xfu4oQnUUez5VnyRZLYE88vCCSe/z/p8J2JX3yvPp4YPVIVNtwP
Z6WsN32LlOkWQAz7eO+LTetlZkXF1VqYkE/kJtYYhkXdtJjwS5QR/SpIDDlTO4iF
sLQuBy+cQOePp6GzjDgxbswfpMOxpnCDryGS8xTMNaHiFbRgeGXlzqvCSHy9jL+S
Y/VFYQbINZ+2TFFjjqmwCD8wxbdP6RV0SSCoW+FYb4dH1O12b61a0FkTcsBCzbDP
SYAf/BVleFcT67a7ldWlQa8v0No96EiAmjlYXgTSv5J3JNPgHbnFlVGv0YxaXN0k
9o7TU5FGtBmmJbIXSjKR0RKRK2yc5PXqkGiF526BhyY4Paons/tt9Ep0bAFkq33b
q4be421F9i5AeyTFJcaZCk1l716apMhTDtYHMJisO7MifN24ACRuZtWxZ1O0tUmQ
1N9CrSJ00EmqdteOEPZoL/qanlKwSODVmSlErJ+Y+FuX+kGtcwRKPd69MnacH9tY
w/Jf/es2Llez5mCsvfOLebkYfOxVaGq4LUuvb3qx/kEjlOliro/Vvl0urhryrsIU
tzA5ER7YDv1M8PpGR5zV/u/2uG3k9zWYMaKFN8datqLcpuDXh1Y0Z6cpsBRZ1hVm
vRKkL62pSG7sYEpHcHM9ZyC06+LzcyjjTug8zBoHU5Z7oUnxYItcakev1yw1QNyH
7ChgjRQKpbOhnCUdSHihWDQnp4IYMJonC/5rHtMZDlbbxRY3J/2r+QO7WB4Cd14h
4AuSxYd9K7+/rTE9uUkBgWm1MCvXo1rhDTpvUhBfLhPeGq3UN5dWBzSCOmaVqVpp
NaoR2fDB6WXJFnBcHJWm57xj3QoS7b5p6b3KVnC84oAO+YtYIbF/d5rWfRtJIZp9
g29DsIJq6ALa3+UwTXXRH6oRy47/J+Ay5vHE/hYcHQgaTazNufY76AHOUo5zzal7
QUqgce33M8SbTBwl7sISDODjsegtPBmlNne1xI56t4XMPBnJJ8Z3mPaCs/cgPNQp
cZ6Siv6OUf0T9kGpIPkzMc5RrQD96AGPvaQZIf5n3s+7pLl+bq8xkl9FovSAGLsy
ti5RcmkTdXbefAOosUkTyOwE162Jp109E8qcdnvrjq7W6ZvdxhUTxV9WJreswpnP
DVqpquma7pvSSMTGGZnRFB1TA9g8j4HCkQQ10oAeYGkP7bR1H3WcwbZAeqwYYOHG
bFdSJFNOzxIDk7zR7zH4+k6B4aQf8gw+LeGKzWeDN13OynDR349hntFr/TiOQr9K
dmszEvstrBtcoDe+OD1tewJp3lHikKkutJ15kpFAludyfWbUuOCAcZwrG/h6KYe4
cj//9pSBu1Nb9QXyE4GthTMBk4DZb1g8/60qPCS50wbGMLkHwFSvajDod7B1DVyq
tyyJINnQDrx/jFX14yeKbZ9Jqo4tp3EsUa2DxadACalkeZvplIz13bB8Kcaw52PM
DPzGaHfkppfG5MBj/HrMy30e1r7tYzUmf+F6CE4gL7VeuF0LMDSJuWmA/Njtcgpn
nCAQGD4zaUk+ONPnpW97nhh0aE8zW8JAsZDQKJzPSD3o3OPM2uZelPMITKVOB4rQ
A2aKWI7HlgmTII0ROQOpJWONr4nAU2QVvWcH5mv4nHSlpwN3SrFGWjJ6T91mfH9M
yb0TdsxRpV/cMc4IjnUVpzlpRDV2ne3UWW9HYsFtQts7+iFvMsUGva8bzZtYbB4J
A9qQvTakC3yOuzwtnDL0jukeHRM+kjYvrWE2+GAvxFn6heqHEaKBLlOouSumZonb
XSnX0wLVilnKn/T3QTEQ7zH+rXrDMGr0mU1zef91VV1xJfxYzgAD573g6l7dO4xd
FXJJrR4rnVk0G2dr+QQEISGe93I0lbDfdKThDYUwG/fly4cBNsGYOrt7p8+kNOmo
57cxx6ckCkw86PjoHF/hX8ciuzJW4ey+1HHPrKUmcXut90MgE2F8QLu4GDwFnypd
T2QWqDs2eRfw/wTKnDLl6yXSgIe0GRuVx/ew7/JIbULjGHaRsgjBjnflDCGmYyyO
sTZgkAkTrGryAsxsZQ+NBAvQ4c1wGBaXntqfhPnQn8VIsOgSsmuP9OEzfIUVMX2D
dFgpqGsliBUmBarmd/jlSagrO4h707x79/S/3ZSGxiWFcWCy/guCXBfl65oImUmK
aN+iYf5EFDoNE6cTqK9+ul5EETpXEqoJbHBGWe03Me8T34bS8H23v6da0ixjOy+A
nBKO7UZvQDRwN2sCvyVgMDyzvxmZnLR+zBitaLgmxKW5HKXVe1rwd5ht+nvYPG0G
4EulQjll2ziK25cw8KPl0ZcaYZb43uplkAXezonysKG6KgGYaMpWIE0QCgeM6KkJ
f8Ng2haf/lmCbkwwzerHvlsZnrQ5Z4Aq3GJWem1GYzUDfnOQNlm6aC4p8t8bHqOB
DaotYEqax2bpCtnBEASLeIr2o/mITxCfIv79oi55MTIxSxv/RopG9ZTzvKtWk1mX
otjW6iQJzj5nhfBT+PRfiUktqBaFY/14Kny81iNhh2mHmSR532kAO1XECpVJms3x
OP5rdCtUhRUm7OB15RaW4d/XSpQZem1PpgYvd/CMmFem22RoT0ZSZCF7Bp3cUPV2
F4WRfI/dIZDKohOLYTENC/tlUuz5ujCAEnqUlEGf8kqM4Orm+nQX0Yk3Q1XYBV2D
wh0txmjjb9QqJ+gODGRO3f4a/AwYsNkRBiVr1GjQ/MZ5I+2oc7RbRuNOpU9qB3V/
lzaqOHkvnZe0odAvNq3drxTIyIpKO2G9QGJoptw14wz9PLkrQ2irZF7SEVe6QBfu
iYvikwb4hjKQcNaXRomRsOlr0ELaI+qGHU3HsgZSYisgK3sSQR3qltGXPPqyr7qQ
1bNSmYbBjt3dliUSA3z0pNruzzgimMFfBUVnbsfgdmbblAkghXcr65pTkD+N++iP
HGwp669hxyxq8mq16lx/YWpdCGhinzzhZ3VjQStYtjXNJEVRmGqg9eqdHVDtTCN+
xxXzLdq6W4Bh8Z1+3m22utBxn4dHGz4BSrOOiNSWbc1yLAFco/m11a+yFcyLu2nQ
DYtn2viH88dkYWgDM+ULbtJN6isQYULWWJifJyWXZCzBlaYc4K3fhM6pVHVZgho8
CFFnvWIGQgpRj+BS09bMYSbHpFIlTS5T0X8fr8vlRP1jpSqkZjPnLuA4XCXfl+kR
HYpnkqwE1Uza0HLLZ22Y6+Y51BWspOAAG0qqvH4sh9tnrwSHs28CGLQA2fabYxtk
PcxKBIxupf+kaXY3Z9P18NmdiE5cAKt7bv4cpKERtKOS25Xqh0runtgNOzxS3ve4
tYJblWDFm3tj/MbOC23W6MSzGOQwgAoFRWPvUZZbuwtHQBx1qE9Af1DSiywTlgAz
+DtghhC2+XHTzulH1wwUMva3kxxzZdD/X0C6//LXSjUGzuNdTy42o6HsNVKCUVhR
b5VYCq4JIWWoiGc2Dxb/mA93O8QcNO/F8eCZX3jKz6oe0JzeNbUCjMmaIMVmI3s/
5PtoWpodbmtaRwusfvabyVxgkRF0sAxwQU8hqvHfH2CYZyKOugIeU30zeI32yQyT
2lguEYU1ZOonYs4Qzc5xDKBlPK283qYGYTU85mq9CjP/BzHWdaUz4PG2n3wpG2J4
Va3UyA/El1a/pFjbgr73u17YrcONlzT3u/fnHerdTj+8DSVZ4EbU2nG+o4o+zqKy
YsGbHNgnf40Tp+oLVEbWTA2y1spvUArbATbViR5eR1I49IX2v/MFIg3sJrt1HLBg
90PQub4TfsmNdx2ug2MV7G4NuT8B/bppBn+NYjdniDa1TxuzN+UNAJtvmgwCRRiX
sMCv0Zti30mPAj0Bim83JYszhGDIpKwNAYgnK/MaTf5NSYX6N0jPWr//9R1tRxOf
Nwh2p1vt6QBR4Hb3/AagV2iJsm7+rORN5jFgmAEdSY+221/a7o3IdjmDGX/zNmvH
GyQB42qg/ADSLH28qJwObtEB/9flSOGNhqVbRhCyeJvEIYSRiGCDyP5z2VOeApyj
T7JG0+5p6kfEH7Ykdn2iQoWIGPeDUcIVIlZufWS0ypQGqrhCH/hXYXCI1Fn8IZ3v
tJ0A5kU1RsOE5CEQWKXqXHYHY4K5yns4Jrr4/fQHR2XVpgp8Jt+vWinRGXPu3Ebz
l+Haj/TssErWSV9H+i9jSiJY3xFPiTyCOWfZ7wuiSLozB6eYunOu6cuw778sNvIa
xCmLqkHrRRMmNdOUFnaSPKLf9kBdwJCHt8LrIraMlag1SPOgalLXHGiMmWw5L57L
70R3M6SHDkXo9e6wObd69tQzfGh5VXrxGiaA3LLNY3as7PzS31Y1I4LaZ8/Z1Fab
h+DsUaH0KrHwytPk0igZ56a3/CkiHVOLbVedXW+91CZkOskc2u/jwoO1r5IJA3Oa
NYB7DMU3AL01jEE3NzSib21bRysmK/mJ0ZAbeMpNGB+nsICQYzInrkUBXbwdJm8u
PUhQCONILoYzj/a5CKB7reB/AimknciIZamSUtM4+W8Mm17VZ1fEZbXmcDAvO7dY
UwvWV8dQ0pTszFNu2JhCY4YdLRSlUDtjOWEk7AcMwga5njUWHIvSFQKFn/7iDfg7
YkuY/0Kj3KZXaD9EKVNYVqW3sZs5+7Wmi9YF4cqJqW6XYrZeGZbtT1PVqbAAca1J
YTo2c1CYy/FWpz/h0a5Y8ckYPFhdVZECNoXmQVUbgBUHufrCnJQA6Xfr4lxtsGzd
xHpKOpp8LClL8oohLODVnlcAEWuNMfoEO9v48cd853nXbxukXGF5ecOlUkW3371J
UsVPRbGHOhJoQjfuBCQ6G86DbmQbDnee+/LgRvDNDm+vYC6UiZf/ENXauFasDitY
Etq5/ku9rIomkB06HQjhUaOwkkvx3RbYYuj9/bup1DD2nLS+7Hbmo2h1rIZd2bd6
0N8oUFHsAhq/q8Xl9wpzJ3Oe6Ew3FvKsHPgq47kvQym9w0/ruS5iVUuWm8EFTDZg
AIFWv9Gi0GErIHuT79WuOK5SYzyk5yI6x940wUp9cmJBVN6h3FS492VtEuCCt9Rm
wKLnsFNoZtDtJJreD9YSkuUFRklMzPPOY8G33MNpFpHQTsXWnPDiPByjFRxfI4Vb
B5S3x0/2litUPYfpifUXXdPp1MxiiMCK1rWAGhGB9afAi+TQ4hDTKBRBJVlgjjQE
1ROa2XAXRkjVjkzKacbQppZ9jOQGl7WL69FhD60VURXkmUjp0WawyFOdxjGl+wiP
dXU56BHEdH0QIfGBy7kUvyOMBKjvGJjsVDh9ncK3C/evs4IyQDzBWmZJ9EPJaQVz
CfJ1GcLU7Ac+XmMy8kE+GzwffqC76CKQEvQ+C7C2b9sLhajB34um+buYNaWcUeLv
HoC3GTEDF6xBaVeWCDG4BExvIcWZRyvcukZBvwfZi3Xd3n1uHaND8EEX3KmwUIGl
xe9qFynx08zZbxmr0andepnvyMnakcJiRwr5We8WvI4MmAuyuTObrHGPPxUWpG0Y
+AKpVMEH77XkTGxMTPil8TUTZZ9AL3Zomw0iY7rivBd1m2UCvp1bEhqKg4gKqIAM
L6pWPMRzxBDrdBWFp6DDeAeHk/eoo0t20AtWfTv9/bBqi86RoydB19BzZLmH77Vb
SG5B3hnPJ4zMqgrCfm14I2PzHxQ8CG7dEAlOnBUjyRCfoDq4sVGUifYsthqVCtRg
EV8aJCgkuINgW3/DjEu38P0Yj8dccaK0KMeopPW3sQzbdwP25lepqCTMt6fk2RbB
CWx/IAJWTTywos+mvCQi+lVi6RiEYgl4DUfMxHoGNuJk0QW0JV1kEg1GbEVAD5r4
j6Fy1v5Aj8CZXYuGeleS30Nga3yGeW5/WYxSYLfasZj1mQAPkcTseSLo0sUsgTk8
zq8cKHaNN023pU4s1YFtpDsaCK7sQj/cHUHwW0TqppgXxAVg/GmuYEAnYBNofOJB
VQJFys2zu/oJW5jf93iVkImthaVnQluTWAFdbpBJA74i6IKVKx87mpP6S1q1tteg
UQVHnICT/fjCQ9Nf0dLHlYJ2t72aPVhkJF1dO8SU8oydnHWUjEgCRu3yfvvme9Oh
WKuybREN+gmajJhwVeFldhhJz0ZTdgV4g0p1pPHFxpRl0/XY6GZ2t9o0CjLg2JUR
YVybkepwWPz8qK/G5FGscolj/C026zJRd2n4ZkF8jbajBkKDBkpEr41g674Q//nC
LIQpBr5S7EOkR8RF+UuMPzWI8EeOlMqVnQTNX3j+gUY9qyxOIJkKQLyycbZ2WKNa
z5JtstdHB+2dSworxEN28l1y5CnIqq5I4baaX98N3jxeHGlYGqxI2CDqH5vivK+8
wac3qZpAcqiwNBR+4PVQL01ppZJjGBR/oVAaM/wb3RDJvDeixd+UCaxzgw4Cz39j
HK/9z1O9AHBraw0LGD0ij/xvPbofuFPR9Zj0/iZKloe+/Pv+5vuNhlT6wSPjjvl8
Fb5Z8wx52WHVp/diwxLuGdfMfh7oedZYRXA7HL6X+tM1Xv9z6t71wtHK9jswjre0
wArNzn9lYcHlI48f+atk6r1Qoa1hkSkOOucw1LEiUTWVN1ySoZJ+ikYDaSfaTQsh
yK3kqxNwnGD+YZJ6UfTPPc46Lg525RYqBln1NwHRmN63oKmagumF6aHp7/XUMbAp
ANCcrCVc79O2xcYmkcUK9ztyCimX9Ftj+QmxtoGUFfR3LqcbCqDGkGRpQV5gkBP8
rB4szTCZGJcX6EuWZu6WjOiK0M0TQJk0FIp5vACfTtS+Do8a2NxJQpWqXzEhoieg
OfcPeEWO9PKtSowk4vxjQALC00h2finHviqYqiqRl05utm+86b9UVIPpCMP3Zyee
JEnr/i4Bv2FxWF56wAg/DvGUAO5YjzUgX1zK7gRtR4rcM91pSuFYaQJ4Hmx0CEVW
NkLweDseXjYPqUOlTsexGcvDqizlfRFoo9IbXjswKCBwYTgr9te6YKztazi0qd4w
ndL3WI9fc6Ds8dNtwJd3Dul6uFLEx/IlId3kdLpxqoD0deeSMb1uCO5PG1IFz+G2
iEHXa1bxQgSnCYWqTZVXgVcrmIsAbs/OAep4bxxYxBg2WxtOsHkDRkgXT1det9t+
34mbzZoNOtd75mZNfOCdDi28JCdlHHmVukjexda9vNUnkQAVvUl6uM7hYxQ3kDtQ
Mp0h/yd6IR0qcyqvHAajwvOuJr4efDNvWXFKQt/QM3d1tZCPavrp790+JP/45aVt
6St3Gw9SbcNpxOsKIPvAiCmODQRrQWOtkZbNedjm8cW2hHnaqfySiENN/9CMnGvQ
/gg8ZGaAzaiV1dIXXTb9b5BWlqn2hZAOumIkQJHZV2DavjMjWi9eo3tEnAPMQs7t
3L9Mpq0XD1uIpduV1solgjB7ZZJlg5qEe5txVgsuD2kMWqPM6CkNnh0qlfhshbZZ
1+ZgOOA/M4Rld+xtslC7MzzzvUb+lO4KTiH9JzW/H4pn9GAxYPr/t2X+P9ftikHV
3i5ePGmYHgd4rglAFT4uhBd3QuKFrC8OOEX/tMgtx5Hf6Ymanxwn0JTtebr1c3bd
8yl2TZ4TIpOHrwRKXi3butKnI2e9BP4LhPHOgds3ZhHv9lh23UgcJ8fiiYA7aeR8
0Rn8yM58ZkY59q6mJJFentUccbFD9NAzBqalta8j6SNLSfheV+kPjZfN0TfIM0hR
IZYaf8WE+wmfhNv6B30DWcmP6m3Mhm/k5hmwYrsOKv3tfnRk4ItTSUUw4CAdajIh
rBT6ZnpBldSOmdEKT70jkVuQ7knOeVNYqr3uPurfRANzPTvP3ZtywE0ZsVzaQk1Y
Yo5MlT/BqHuYDJkSnp7Mni8SByfGGjbWAnHM06OLwMUJsOzk3VID7FL/sB6y2/1i
x+zxGl4wkN3BCyyFuENA3jRUvaFnRkqiowwdKTZjXa18O67jgHq6gBoXyoy/TzqF
ixRTOQKA6LGhHixM6OeK4OeYud0rYPFPNVHIcUF54wR2JYjLBVDyhV6flhiVPBND
F69roAXYDcdHnBrEc4CqnGpQs6uS8tzqIok7jC00dkoaEyAFPe1GiqcXX9HKQMCE
0fM5Lihbougq7R7yeZCscP4rP389H0ceLfgynphDVIFhwPrhizNGoiyAOgeCVPwS
H+JN/WHuD5mB6nGAxV6LVifU446RIHEqgkw+F1QA+fvA+TDH6rXCHg/FUfpphZHN
W2kb+2d8EwTYJ5q+hSG5V/QqJpit003ZPUCW95CLTx3KqMInSc8XP57KsvekIcb8
SvQKl3b8ze56vu6uAHsmOg6G+av9+eIccy1bmn4VYetFdGpvu31PXF49wZcfcr8M
IyUJO9yuNH6J6m0peUeGGCmmhmzK8uY6i3WeBpbsCEwndkREHLw1NBXLjXQNp5tP
p8Wkl8AgArZEx2V2Xc3IYo9UiOEx9+7EUUdOrA/8j4cxIDXDwR4GOSPo1y9WGwh8
nCATCVkqf4056LkDAAvH2IxiFPApazcdTj9LOlOKJTk7yI4wd8rAUC3xdBlc3ScL
Wad8iLgBtiEGTmtolxFUsUd7G5BEShiZUAo5zVr6yjiU9nZe5V/PjuRR1JD92slf
mHc8XCla592/RdIc1eRyxzHJfe9K8VIAV9B8N55P8gQbPS8VWFa0ohxh6SkjC9eJ
e0yldQDsWdWwgtdI2jBAYc0xoouj22m97e5JFBabi2F05EBLshzC2yHBKkpWgJMd
GBjqV7lofQBfGS9AwFYOACMkOUbSOdrILPuP+D1ypkpcI3JaHgWKCdJLJJybMsFD
aqHWLpa4FXEvt0KZR9JHaMQ7izYVpRCOV8qOp81q7evqOG5VFCU6pbBeSN3pQbtB
IM9GcpK1rYPxoXg4PHAJCl+8QiEyVPcqS0Rt4/1hMa69PnZv88JRrZ4DfYb52Oi/
jsWTsDenotl8MOiggOHnwJblg03eR+YeB+ikrUeHibpiiLIjcZ5TiV6+tFEy1Zt7
eNmpqDo8pRvHnWBHwSPnDm03BwmZGRnEW3P5jSx2D9ephwTIBV31wvr1NQamfh61
d71eKQGjm9OeGc2LuMjVxQgFIYWQPchfxUILaB2sTmQZ3nMGP4fZGcl/phcSDm0W
814Aw4TchLisWFjrSQq8wyy+XwOlmK8G1rAUj+0KzMR41Ktf3Q9TmittahB/JRve
U16hxTyB+OsvGZVKgTTbxiqFqxHMf4SZjGKqA/TvHePKWrEbFOqzppBUhlUartWa
aVxB1DoiGCpMUJeu6dcwoNUig155aKMckNurbGoSiL5qDHSxGb78dN5rHCkKNjWB
lqvrgF4qvTIZUkGGuwvJSB4zgkkXmpgiF/oEIDA4PlHacuxQ0HWIWxlLdjTgZGMv
Hrqe+hbrHAEYoabdbPnEG4ZmOuU5ifqFfokrknhXgb+aFeUdaKY6KiU8J7PSETtN
KB3ebXhppqYgoHOpIW0lAxDSmiOrsO6iINRWQHp6mDOqqlqLM98jb5AUpDxRppWb
rwmEzq5rOF8+LBINg9Ubr6alHBz96s3YHsEmUbScOWKnqXw4H3HJJTdsY9uEhMum
ieAwL+nfsNH3hg/s4pwWDSIpLxHnmLRa6EJjya/Ie68h+7wwYFqwPpGCy8tjoE4B
Bjw9b1BdGBWtkcUV/Itpi8IKNusqe6jACmM5SgOrSLS4iqBuJSmXAKLzdpo6ueFj
YmPBSalkQ/MhdY3wI19CZk5iTE+Gu+jFF44N+B3cqC7JnJBpHTj8yCk4LgL4CJ3X
H4erGorXdBNuG6J+9AcPohrQjpUYuTeR3Cl175wSIkyzQSEoO9eHkWUBCM8cOftz
kISJDd9/0jzD5XRHDEvFegKQZz2+e1QSGmmjEKIBFjp4Qa6uDLzhyRhLflU+T4Pe
6aIwFI/UuFjZXrMR1zW/izwx9y+GaJgR6kkCM1WDrIGQ4YDTDfCqUWHMxJNlOFi5
rVGLiezbO5UvoD8O9SVJjwngLOYq5AKGF/WQxUWiiNVEV4HZ0ZRI+iyrLNNXqetY
KyFhrnO/4Sp3blLlyYgGNvHK8hI3hZJgTY5rrVxCA5lZnECQhRTMWpRK25fL3OH6
3biKUbEPSnWK24tuiavdmX7+P6Z24e7RmpdVFxQqPBwjGZ7XvSFc8mKbrSAiK0BA
knkUrpu3qveYi5vTn31HRZlJTkfrRLONR3ZKvxrJsAQ47QbLj2Q4n0WL8GV1A3sz
CGw8arBzEMpCCk0KduZAcuZeHp3T926vKM/+MfuvIcW1C6w/UqX5H/dvQray9aTx
Ucc+v9fGweXKQyJmydp9hgfI0+OxLqOiieq6VGw2+cf7PKTSRzQ5R+XgjhJGZAvH
y52nEpC/CMgWIfYBLFwUeG6ak4iy36rKTpV45cqf6V6v6msnrgvXiFCu4y/r+dHW
unOKhLeQhqPPqbToyLIKq/hg9ESdoDiZnaoknwg4XE8EsBLuJ4tupLbYO6GfaYDX
2IXsF1Q1LdRd6n3zko6elwKX4894j+p6mIR0RKtMHMJz85u/BFsw6JY9xKEWTdDe
WYjqIWTf67+RL+Mq+Ajp+3J79vrp8scHnBgL/6ziTOV1qsRSYbfUNiinZa9V9Qkq
DyTlGF+zpTPGHgYj4gZsO2ZlN139AY1pjQDYCtJAYT4ej1jnmf2UcakQgukpOetl
sZT6us+o8w6Zy13IZdIdNWOXglpviNWGc8+pqtMER/yvMv3Oxjf99187cAHSnYtT
O70i17sgaFvJA6lvAQUXejzSRYIsGBr7Z5T81JfKZHqCitd8/+9o56q7VmxKbFhO
7HqIswzB8JYtdo/hE8tgdjmQO70skhexFkoa3qVe41aAsqoCqjUxRPhKQ591ebrX
kXxayvys0iu8KlNqO0w1RukQeITEILCGSlfHECk1SNLQXX0PphM3BFAehPGusGGN
JsRbDSRW5RGU3Hox1XuXQ7HAmVF4YpDfXDsuUEsvYrWerbt3cHIiT2kRDYxuzE5E
VodoYSfj3QmcYhOCdQzpuF/gSlkol5hfg5+zHb2w/FQ2XW1cUQgS9dHkmWtuR6V7
XLM5fmF+AGNNeKZPZuv+XhYFKut0Le0cMC669+4hlMRdwkikYpIcMtOr3J5gJGpf
DnjOsdjIo2rNh+QK4yNqSNH55NE1/6xZgfOeoR6beXdgzb6Jpq9VlV/6mcDhP7nn
91AVQ5NT5N3ezI4fTP6eHkRvKRmKpzxX7BqS9P+DEnqy51Jd2T3nDqkuCS7/sDP+
40jo7DQOANOuzXmLyBZWP47+BuM/e28uegVZcg9BRuaooGGGiUoXth11ygM5HF10
op4Qc8qAa/LnZaLZR+zDsV/WPmFVC4NDyc3lHctjSDiSrlEzP4XxgReng4GGtxFE
Sk3G268npelb2/BD7rzdnAiSn2NoT+7bLIV7lE7OQBFltKFK2dU2KpbSy1w1kNYP
ZayTR4tToEFkyhgYMV99owmI3K8SWduEHb/o3ARyw7pB+HUOv7/bayqZ/fClqzRg
b8xNjlby4Uuoajp6cKl/6bqvE0lSxvo04IGAQh5yErGmJ1XCSEJ8QdUf6/JfWYyE
7LeconDxruMghqi6p5G20Wz+YFTL7yvQoShjSIr5KaZkcJkhd0veWVuu59faygdy
Vhl0+7aF9JUALDvyWsljAdBW0kobP/mYTwn3iGEYLxZdfBa0yiwU04jtBBdflVpg
5ZO8wVnEukkO1+eL9rQlFGjvVyzaBkZFGuhi5CGFH3IWyi2tL+WV2KUk58w1VUOU
63M40RvgMCFVJQpu6u5hjX1exPyAxWyQQJJQdgfR5HCo/rB85XgWI5vDzUnPjg2L
1MWTnOv7nZVixr2PXVFRm9EMPmBO1hV2SZawaYLfqAORAB3YA9+bY9VtN/WDvpKT
jWm+wMub6W8X3pn+5j6etg6p4IzLmhccKBo+3pfi1X/NRruTHm23XLi4EjxKXX9+
e+jrq63fQa+LXhIm0GbM0Jw+hWQZ6mnFfPEGChSdm3JE6xwbCY2Iwy3Wcbakui9T
BkOvoR8bj/wSK3wqzzkrJf6buKAqjcR4p7N1eF/cMmfcX0odYd3sedRjIWdG7rGz
nkrItu2jTwDHhbFEDsQCKfB6iA3XEPK74dbbtPp2XwwVFkmQDII5X1B2h+96RHwy
tFNNQxMp9DfuKMzPpO+tEZaWGDBPt4O8bBp7FuShQwb+eCnzlVcY9n0FsrRsTzDP
LDIz/ZGXVGxC0dBoQM3Pfbqk3iLHD2WaxnSvtgxRKnqCnCKHgOC/gh4LDDiwtuF+
rMc5uL3QTu7X073Fed1f1XOwnsKxMtF8wpiQtCkiSt01IPmrmk6JmSO38yUcLkkd
s4qE+fviFItNtTfpaLPZt/1NRZd1oEuyXdyhCItqSyDujhPcGQAFcyJI9bUlQYcm
d6m+og0Fxn5+AhOMsig+shS9KFclniAVZ+EU+q9a+LPfzzUmWW3ZqcBaMDHfNBR3
BcEDonR8sCtfhDweHql6D9Q4TJ6UyVz9zOgJuG47nxOkRLnST4JWulcDZJdZX2Cm
UQtip+D45O9aRf2z7APr5InKabJ5vDIdZ5nTgSV6v5VPDfPA1PEeeJkCgp7cLP8m
0gfPwi+ORJ5tfv90F0ccnFE3i2JErkVm7YfGITxVma+bXJpgT3F8RZ8nFm02OMsE
cGzxDkJvC1617inJ7q0Ho7HSzcRpiV1zcaeHRWfYKDgmH4LnwqOUqFO1HVOkuT7p
luoiYHItAgX63Xwt1GJ9VQn8C5XjEEGP/RXDZZMXNYsrx20wdrJ4ujCrh+9M7jGc
hG/o9HSNFFEikZute/sCE131+FQk522Z+fvNmpEmtZITNe0WSDfDufM5M6uZjSEb
HUcvJjlJpKM9ysDEWm/D6Jz6aZnPMwCDlBMFm4mdiZSGEIbPtzsUPZZzf14z+wbg
+h/NtuG1yDFyaGVMizPlCh+8hrxsWcSubBegEd9kv7sJJGLmfWBAxabPMVDjtkKY
DqGflpY7tSHpArXqx+i2M8MxR0Ew1eztwnDi20qhY2ZQ2SZa/BZT273gJQGSQMWE
V7I8uApUruDAi5R0mrLVf8uwwnzb9xwsmKUUA1/KigAxyk/E0E9ZhRsYQmwvYcck
+lMVKZUsvKZ6aO14u5BUbzLSQNp2pD9f2ytf7Rt28lqqCGFnxKis0SNXcd6SJIb4
XrdfExxpq2JRW+OgoY4LGRzxGZnHWBQMpDuLOTJ5vYSumQGCX4lH0Bh1y/kKYeZ+
oyGdlN7xmZU/6LZLcxzipIgZPqFfOoOQIirbotNKSuQs3JxChAEkPexonAbpd/Is
fUk2R7jRnQHg8/taTBOOMIW/+F/k7LYBd6UDE6StwmJRrjzfTk7k+5DNgLQ20FI8
7fEtPcr0hS+IEa808z8JBhtDRDYAfrgod/KTrwpw9wO+PahvtvEH3hex/QC/Nbgm
aG1H5oIVtIPdcGFIF5ZXBwAdvKYVp528urbnO6YAdOfLBg9MOp9f7v+LUPjj43Ur
YNKA4FcD3MLvCHvCKzZfTEpuoBvKSKjUDVrOhgfEq2TgB08tA/H7ix7X3a2c2q+8
gTyKLlETW4sSBYamwGONA/bmj6Q8SS5Qu+LQbIfJL4j+QRKSEJfThT6RaAGVfqjq
NQr3zE9M4EBqRRBGJuq2iTFZqbiThbZxepSbk/a7C980Q8jhdjBiVZR7sVXx3EX8
+itDiSFfBgm38tlrVojlIbLqnxsVnDUr/mFdFW6JsmQK0CCwZWsFo5ikk8kpgLdu
6xE/Z+HDbbwKTldlHbd5A+44aQ0DiHDpH2vXbPSTDjt4PofpOrbei85Ywy1Wi3vh
qcgfUjkVZMdRPT+URe1muAntXCwSWYZJblg8WFfWTOJsRVraELssTulXerTDzFJK
Sm1oTGB8yc7prvk6GVaukslyDW2VryGloIs33G9HlWsR5y6SCSVMoPC/ADuvVG45
auLnNVd7Rao9AsinSrztPKtScCKPurJfCAPhmyqkJM9o/9VyBdh7+TpDubjN5AUT
BCZLS4rVwlYFAh4d17bLemG8NmAcI9NBkFpDXZJmrKpPTdFUeKRENYcq38XPG0w8
28BtnFh21O/XNTjQbOWs5F6iwjpq7ZLPULHqoQBhPJ4iEB/V5RHYsMG8zkxeEIZ5
/pHkheszWM+im6lLX+9YaIWCh7Vu5YEBNoMiUf4IM12vIcjttm15tvyQJ7mm07qA
nPTGYwBmqJPsdh4v8ZGtdU4VlDJUdRRAR33gBjecXCsqYCZxwV5Nrlqlxc+utIU8
srzRexfRSDfjx6cqgpOsDFtPRmYYQQa3+d6d2Z7eD+Ji9MAfQvjgaEv909ZvDzyu
6fyHyNOcEw/EE5QrHNMnMMYC5yvAewBc38hQOFLVTrTu1zMpfv+bZzCpUOmmwTEz
noix9jrLmTkX/FvDQKL7Kcb4CqEym8/4HO1bmPLcCFaHdvWmcDkEM4S3XA+UF4Ac
Cz/SVolggRlVioi/qnlCakCw7KXWdYv8cQN7qtZZgx/NCm4jaUzDsvRp73kezJfI
FFE+DSssIV4z5Bn5zRBBafrOEVFfPeMR+TwJcG3ILg8Lmh5C7vmoaKNc3dPtUYmv
T3Suc+csy6SXo9pcWGOqulD7dsmfueWdv+00QUWIDG1z+ofiEyzyzfclvvtCuU8O
MS7A0NflJTZ3N1NB7bs/nbBNCQTVcXjn/SetWUCCo2YPR8n2nNH4z+o2FQoG4oto
4VeNZdvb7tJFQapv59dYscc2oj0I/fYn6vQowUtRw+vX2IwMLA6nj4cF5lrciYaa
tjzc/mTx1SS0U67v5IX+aHDIFmJtpb6k8vcbYqh/h8+snl318fQVanbQomZcZF5n
lBKEZ7/Nm1emMjucDksE/kEmu+3LCFnCGKadVeD8hvtPpzxUXTa2x4NYhfkm3W4m
xJzqF1OwV82edDeO3HKixriOQTznSOXcdgYa+1tUdkn3eEL2KWr92cuMoCZ4MYxY
0eVrPtWTA3eg4fbKy/r8LTLzqNHgjmYJ1gWx75TTgapnrIpTe+0Tb9KLRbI7mLqn
EWEOSBR2HCP5v0JPOV8GgqMsZm1dY5FFUoqXxNzeQdqP25HUiw71zufdWzBZoyNo
Vae7i9ub7kAYH0DG6ISIq7z50BD/+3cwanJz3mRRecCFLAORhr1cLt1woW1CeCA4
mcU1qnoSDeWS+ezWOteyCr16zetl0Z4GQgd6l34J76QOHjsUfKNJkv8DoKaimGbT
bC0Nd5xYvWqrINeBH862+1OErQ7QY/kZBKyVbP+RIbQ7Ddi9kVnIysW+GquAiqvo
FNb4k2WolK2U0ITQzmYHM/a7Gs2ewaudSeru1D9k0i3fEp/ZUNM7hzY8I29SJEpS
c1UjOne7ADCXkb5FRXqzPEfJUyX5JUD/e0X4CeEYla1FuBefusA60bA4uBcmTBZK
TpIns5ltYTxj3VVFq01huBWK+ia+SqxJZRYogv3IZ+7aQv794kec9yjQG+TNpTSh
QpGOms2ATexEk2LS39WMitbDVHL15SSgD+Yry25SUvgASB9ymj/OOgvXbYn4rxRq
KxLn3YA5muEtmVvW7GP8udVmuwnUVkjH5pYvBpXugpFr78XYxUPQqYS8iZLQdqBN
ez3yODTCS7xQaf/f5ODJnQEN1sgBNMxPSE/xqjlQC3yLU7QaFAbAfvKE33BpNf1Y
Kg1OGZPwutWoAHFHPbIQO4xQXAqs6t0AN+fhLmdRu4w0bEMdCDdKyc9SOwo54zl8
hRAnMMNp/tzAWndG8bOJuomuoJuGRsMEB8K3O34YP/S0jKplUtbU+umdUBaGtY15
PoVsITGsD2qSo4vCyR0qhLuFi5iFJmiUAjej6iqCTMXttfEC4qU6L7nEP76miPQO
sicw4A/Ks70EaGo4ICItr95IGR7IlDlnlZEyvT6OwW2s5nkt1+VV/EY+FzL1foh0
lYtcB0oAGpfeGDR/xLFFuNGq6WingUaitqaTxmFw0o0GUqczXl/kiIRjt7TwU3ka
J6e+o0wA0d+CFvht9DJOZyly+mpW5dLY+woi+XR1cJpvjgySk7VTsw6xkmKpRRiY
TRACKCRp1NKNd6Kjf9jXbqB0gl7CGves8RNgZFb0cCUvPl0JoeCY+kgmaoI+cdDL
OATd5Q61h/EXK2tq1GYdUfbKnMOlgEZsj5ZqgpjmzVOVwXGkkXOMH4sRaiJDA/q7
W9tTm4J0E4M5J3ZcXsJhnqTCKuGaC97sci0bj/WTYx4e94+fhXuZJw2hM2duaEip
2D6Ef5J03bpezHLa9/0VbCjd75S+3YH2UO0znZfeD5wTN6Bcb7CTZRHDrWG1IjGn
FCZ+9HRfM0Mwn7yQynH4QIsywHmmUX33p+z3e9hjSE8EQ/AVvGzq2nQjHfYO6kgC
svwviqy4/N/UPgPjSdEPuDb5i/7d70UXPg70A1N7gHe5pynM8ZBMKwn8geYMKeqC
MyQp1q9XU0wEuu2MLjGMcXP6/paMCLtxJHeKGnsjmPPKNHy6MqyZVnCKWujfOvgo
TYae3zzZoIc2TQ1ezxsdQxImdNIziS/O6K/BBhf4lg2g6zBfDV/sTOxEwehUmc/f
VBCRxeQUy557m8KrzJ/uv6DAOH8pejjAtlJUjEAKOa6OtrinKolsTxQJNDBAxaxp
r+h5c+e1EL31kbWY11grS4F/rWU0Fz91+Pta1SDDLsPzJxlLCntc294koHugH6nN
ObxMc/6jsmzGY990/Z9mJg1dQ9+nMjLiC+8q+d2Fbs1QO4/QgBnLKgMOM41RSZnr
gcOxjIN5S1whMXpq7U5/7iqMVbEA7ufKGXXbcaGiGu/vbZWw4+/R+bign+HlUxZA
LfhtwSLBJBKAnMnGYyLIooZOL5YSO1VozAmo8v5pO3C3W+3VJe32wipTewqAedoN
g8aM7nWlb9EB0lAwAnUsz9xIbQdMPh7pmt1gmgHEwlm8S05w1KsOi/m4JB/x4wRj
7k2EYYbf2uWjKSWi+XA1NQFsErb/Mx+XAp/Y3VE6ROqZ9qaqB3Zk6eLhYrYdKXH2
USBRAsODgqwbtFGOfBecPV2aCGEcKmqNdfY4RHFbQfobedcdDiuRN4+I2ds0QCVg
ctzOuuh6xdm2Oz3oYYo02RzsppmqigfBu7SFXUNBLZlg6MAPkjs//4HM0a2mNtwI
NWdO5evt3cnawes9pZQRiM1m0z5A7woHHVGH4ysRGL9no0iHyrQRxY8UK8WBJZyD
iUbCZkDQfHIcalShzToO2ijHc5ZBRN3LmaB27i3CFWrCufsYeHMg/f0pdLt/EL1j
ZLbU48rETXrQEMj7fZaI2bYNTr4HVOVOAZaRSBPHeAaVKMSuzOr2X5ffUHn628qx
2k65SJkNJkl1KU0nrdyAo7PdjMaLR/pVzsyomz9npLq1KCVOxFlSxmkndxSAPOsy
CcOkdv7ZgKgWhNGvrxJMZNnjKZ9v4xFF0LsLcSuvvWrZwMUKUbXfvQ5aVBKUZc2v
03OOTZh2qxu6KfoGsd+CCbaJdKLBJoY/QaxDmBlNs6e71RGraCOnueVdK55A8rpA
uhcP8kDian3n3raVqScopFlghm5Ci8xPl5fAgSZxR9D37Nq4Nq+qn4KS2MQTr9R0
Gdw5x4250l0Mu7cV/Zv0PCCg7L2QUloW1oH1BsDFmmuply0xPhRBAO8XFmnunvD2
njz5xq5JdE7La9p13mPZs4GrsNzPNAvJwOcQi3oo7rPGZsRVLPhzKLxsNrqZRcC8
ylsnPYDMz82YdSgFR7fz3HnEfTm+MJ6GQ/U55G1VVdaOejHPZH37TlQoGEWQBCZl
NcDzIep7E1Zx7R/71WfV9k27XABJu4LQpoGmpIQhjsnc44QrNSr3pi6cSZevinxf
MJLeAwJOudCmv4GS1DZNYD9U/UqHe5zkEBhuW8sXjF2pEjk3WGK4KJCPitC7vpmz
dO+eaLNuVbfOqDjExjVspto8Jbfd4ZQFsw5amQzRmsQy0SVE4BUSBPkRatV33aup
GzIk9TAFRLxhZYke6X5Haie4tYXGkcyiryXD5LXY5fuBy/vqzhKgSCb2tNKQcAP4
x2+CWWSgi4GfNL+NPLXYj+kWSXP+numqqMoSY00aucBlUI4rRQnInYPeZLpR4ZKl
IgCVqtUC5ibDNAGdNDfCo6qBaXoenjUeidS5WbeH8Vjh9WA1jPODtxzzabt8Nx9z
qaLCS/FHz/N/saE1n9hA1DLphfGuSbaL/ehtu2Z8/kmtLLtSjLGBFEBWgSwiX8jM
f5u5/z/SMW+kk8nI2omkSXaQZPmAGhuNT6+FiQZhYgniOtDzH9s2i4+heYAPpkrS
vQpdnzW0RIwpKB+RA07jcejeV5UWS7WZkCjZmF+n8WhDqyZQHSK4zf+DIdBofDPP
Wsrjgv3GyMHJev9I5Y8cgwU4WeVLSiN+rXZqyu1W4jdtar34E211DT1TJZk3gXkl
rpfF+356XuS4hQ5XFa5gyR2AYWlaQkAd7aeni9Of7r7C7elqaHsbB9pWmU3OJn/S
PDw9qBhGTEgOnciZxx8BMTMYJy1WPp00dHteSBnoEjdXEY8Bqvsqi/uPn+uiohzs
mpe1HAT9M2hJYAmC4M0S2Q8gckFMuwZokYWxnsVtf8KvUCAU8YdgDOhnBWvIWA2d
t7ex7QES2SJCOZf8a43uUimraM7I4qX6W8Ryi2zMoy0OcfmFxMKlBfSxssqQIFdR
MjpoR8k9yjufKORZ17R2XXqcbIKcm/JYNeK98DZXw0RPldQ9fph2CSUVGDfwL+k1
j2d+1Rx6kEeI6C8AV0MRxgVnYZIdgn52XrMb84Ci+Q+fj5tzuN8PN/FWT6uyNybS
AfCrMvwq7Nm8sLhK3da0fY6fxfs0JQY7p94i6pMWftAeS+fL9pqLyyQco/mHjYZN
aa2rYlWFDxQtqG8/Xv4Zuy/wat+2pNlvrET1nPqLVUpgz7MuInAqq5nU9ePyeDFB
iCdGwEUmbyDwKathUqSScQZpXovrIoFMtGYD0ivf4hWz+aJHiIxni1Q9gG5aMeGF
cgDAIQOFukY+4XsEwJufdizn2nh/VD4NnN/15VbBMhTLOMkOw0eorsX16BRoqaZD
Dn29FTyHTd4O598if76X+1Mqy+SPSeeCYkHJLxRi9Q+2vI+/mayyZtWM3NxqPjCE
wVtKmeaEnHOBwC++DFxYN9Ma62RiuK56SjOdJ/HykZXrsmMlmjSPJbd0YBk49h75
IfqiDW3VZZDQWHJkvwM2f7IKCT0uz2yaO+a+vJKUIjQ1Mf9v6JvP8xgPb7FqiZ96
midRjug/N+TVSQV0axRWfsOdAk6YX3YY6I1LbjePG2s+PAMelDa1OlnwPBgWrIb3
ldaVSATxgupuhjo4U+Vw/Ax//yIBC6wyM4s937NWQzU7I8ID2vu54J17VeEoDgem
Nm0xyO3HdWygdTMotdd5p3WnUR6KzsgKJw0ObTK4aOc1sayYzMHej9nVhu42ib+p
rh+It8HG4w9ox9I8O5mGAFfaNWw20r2szOcC5iee+eYSCiqmVBBiKXtJJfYus2TY
WCnwEPxWe28T7g3a6/DpCuDUGNqPkC4MFWycYRAZHs6qAPMIGWAqcU3VjI19sLAR
gccS9VNxCsaalHJWzWHA00ENyA0+NSmHUxXf92RKHmz6f+jvl94S+iA4zrxB8apm
K8WLDvACp4Hl29Vsc+f75+96v/CfzzJPV7HZt7LlBbTZzdFoGjix213SZuE6YfUs
+NnAlgQCg8e5K1/UVNp2HxXvhuiwD8cwV69o482w8aOQY5g5K+LdZpi45C0GriM/
4KnLYxoGD98Mhh2O0ykL4Y1DrFC5/v0Db/4mPy32rPzhtPJq2Ir3bpwS05WEXfjd
LwuLLAfssnCwmenpMnBpq10RetzcWIRZyLc6my1ffxOaoX643fo8Dtqp+ciCpnJ2
jGOj9yXvrEVuXa77pPC7iFWtCQTTPpoQLbaRN1OCo+tJKgq2yimQWhkEW4WoAX83
H/gLfQv5Jrp8Ycsu+UaMP2lLZJqixLYRONtCFCKV89bDBxN6S7oHD4loHHxzc3zQ
qrXHqzyLiYnhS3qf7Z9ucBMZ1WtwrMhpkxFGmQHnAPPR8pzOatP8GjxejnbwWUC+
DlYQSTEmKHPGnu62zr97kkU+hBReaXGPRA9nBg6ysTRprl0/P8SsdEGpN9ZKKitR
YgGuvPJuBV5XWjiVEHqBNf9r1fvIGRCY1GfUtUJJltJTMpXHNiPCK+6v+YhFfl/w
IbY3SkK0A/A3wenSG8xGV84/HboGnz03lMyY7Dv+BlvUcyoejjfXOdAMoDFD9f5s
EDEj8GD57kchS+rENz44BPMAEc/STHzKOxUV1yQbdFsDB/w8Q4v8mW83wWR+kMJD
7fZeyM/WnOws4qETeEUDw5voiGHSE9dpPvSyjwjRkkWf4/wHGIr1IjEW2nla69SG
q01nr0QuRJXXaMeYNmYsi3mLWspK7aZWRB3dksfBitdrjx2zUJmUoucTKS+cJu9t
u27ZfFDfBcDiGEA0mfoYIV0InAHdwkO0w1rnd+UjP7GkaTmonG3t2yN3szCo2PBV
9Ik7GLEZfpWLowkGMfFDxLMUZ+Yggjj/sCS07BaJ+O90My+7jaYj8snF8Foyd1G/
Y5JU9mvcjOFklkIEgXV6iZNJsTqAwD/KtE4zUfDx3hDrNp6I0arZUfEs2t+iKvjR
natA/2BBv9UzOVnRPqRvQEnh7bsFHHqfbCyFTBawXItMtE/S8EoSbTdaJuuJnjYj
4cAToH+MBQvPCs81V1Ii9ZuAsCWoaWuhW9iPL+VM9GNSyS0IK5exIGNgObxbBY9T
Wpe2PhwE5axbCEqBNnOL8ekgkFeVVNLHi27CIXTS3SheRaTs9prAJxC0MJjUJHqE
eu6Jystz7DBWgYU+RRRvIH2GXba37vC1OI2EKFQETpLsUewI9Ll59T8SzJM6GdIC
2w58f7jWCvTuhhPICOvDIOlo4pDOvVTcrSDmKrhZvxFXUBq9XOn0uYl4sszIhkIa
ojfU0x3Y9Qb2Q0GAx5CPxbWj7PGxXLx/XLk6gOEMVoC3oHUbDnRjknCb52QLH/4+
pn6Rz6Da36pwLY3kvJQwrAoHDIQOkjoYjjS7iFMinKaoIfS/i0PDYcNAasK/553X
q9EhxJ0SRNwk++Y3Um/gETBtGWDaXNSYerukXyv9e4RzrRJjkIozyTiU9ICnDfvK
2fPOa8x0PDLFtlQa44TZK2vyh3nqx1py03dQfve8x0e5hXBoOEOjF93ZO9HroUvO
pu3+3q5yZ7WLcFkZ2SGYlX7/OpUi+StHWPKIWOF/g3KBf3ke0dKCTBW7EhXMATNn
iXM2balyzrTsNqhHpZ6POJgQ11IxwDWjpg98o7bqJb0CvUoQnEvKrYYfltPD1d2H
mDNzdVU5aEikyfIIeR//sP6dEzK/+EIeSJ5vXJ6yyqkT9M728eS9dCcNQliGqWub
+XIYYPU3NhMeYPNXogBZh+dBFxaW6GU/Wz1KkafQTRJwFFE1yA+g7IhAyTbeb8cn
fCu3P9OtxearIpL1fZqlGvcVPi6diAHiJIrLQ8qIXXeQ6IK6/xNaZpnmHPVx6ai7
MP1RsTCzvq+KavmxTrU5kBQsCKpWHYFfu1cLBvrOWNnmVIvmPmApjK+Ei4DWG5Nq
Id3lEescZHVkXQ+n6WMErBWoaXKntzjBlozXcTASybodVlK/nlSopNKZS9ZvOCvX
ONUW3JqShJXM+bC3r3K8aU6ioyWmGq3YP5zKpeUllmnTiCNPft4iSrNs3Dz/yecw
2/foJtmK7vdfGcCFtMUMIDQ64DC6ypimgaEw+ed9Arx4gKY4xskIrmbnHtWm4NxF
xQO4Wy9AglK+Dr996erHTl2mdTNPHoAXD4B5BjygQz3vXSP3I87UMpA6xg6ZpTQb
8cbZqov26Mo1yky5+7DYHCyA7+arO8E229bYafUmBnYFEnj37MonWf0ZVmiOLPA/
BouBgGqQ754s1GpKkhWKotXmBAipO9eo0PdhfTJHZ6e8Khe7p8vebtTBSX2u0Njj
Dg381jlpUP2+6VeSrGuC7rLGMX0KqCLcleOQbY+TqFyMTJX9vj43BCpYXE1mMjLZ
kgEKIv2hw6AU1H7pc3i173M990e2xADPrq/4ra1hovtEdbLoO7QlPVAhI2UBMCLJ
7AdJ3PVmtThtR0jsKzwjNuZVjYiRtYNgMRiV4gkpm3UZt9DZPgBeu/jBln4HhdFV
FbU/U3NYgRHUuVbLSx+COz7PJgRLB46DZmSph0bjtnLO4Fu6wr/jXQYzeQ97eup8
RxIYfzUm2iidqMkulZytLgn5oVkaKsMbJqA8aEk6nLYDy35mru1Er/ueB13khP7U
TixrV0vPxgT4qvcT5PbbkuNfEugXw5a2KOv3LlxQrJBVzm7uccrmQX7p3Q4yyE68
nknO1fmT4WIngaz/zsOmea2LdT9EGCiQMXEvURDwf339LAcszZ+teXDKUonCR7YQ
26P9Xd9RXCblf341Nc4GzggqodlcJs601Kuznct57OJtbf2cdgGj6vrGDKd7cfPW
Afi72a2NXhrwJvI9xtHqdAfIJ0xeXjFHbk11M06+lIuxLMqltuJVTr/fv6gr4ZKx
Il2AtajlIfuMmu6Jumi6AfH41rUkcsyRk4h0ICc3dgAw84tsAfzZfKD89TdHHKEV
MsIKULKscF80mOjZmZVjbEBqDuii9SoQlikUQQiadOcT+g3vJUsK04fAgQ7r9/D2
ei93LVYTowy2o5GbGRXSJtSkbFYItCB9cKlb+hunwJYi3WLnLlteTVXsHXro6WIP
5YcyJfXQFuW6KrCkYnd+EEXp3GlNAaphNDkYwlcFhroTnnG8MGpc8nLiHFDEPuok
fhFCO1KLBhlCRyvezw6wAXkFIRRWszojB9kwZc1LU9qERsNj0W+schQeHE91CLNR
F7rbkl9VLY4CW3MvOitwkhy2QQVTH0/iAv59mBpw3blvKroQn9BZfQ8zub48nCBZ
rGAVvmmAOqboOaOExPsuVl5BUYIUmTpviV4xoUFAMmqndgBF4Mnp0aENOxeZsRmw
Y2bc+WC6hwsFL820ZfVvHq0bEsIRZW/i44LxcWHytVk4FMl7X7b+uY4TeIytcv4F
9km60mENYfnSmO+NNVBEiB5j2w0I/OpI2kyoB+2cNWEwAJTQAyCTZ/M+GYheT5yX
v0fcHUKosvnynUo2kp4t+AGyFa9oAE1hCj4DxRyZzAOqWzFxisLbhLYf0ar77SFd
8sLZ7YJbLwWw76gbt3nBPsDVi9XRYJNCwgj8KnV4a1c1hNQGZ0iXYDaf+e8LCihV
I7aF7LaRvbFCUbFVg8LEkFTuaIfFweds6eio0PO2sTykTni9oqB8o7P/PUvoP3Za
eNVjA/V+FoSVIH4i18mBsWgMFXBIWFo3ucljTlIH25yQIljENEXU6Xpe48anu2eX
Zzf1dmm4FNIegXEBBHuX9Y9p4mb6eiA9ns57M0ty/4om4e+zCQpGqqQbmHRUpZsu
X92xyIgS+ZVIfIaOC6PbDYr0WMnb79kjzuRRH6+t0fEgbRAmHHy2ZehScLDpULym
IbxRXAcjFPJ15IuPEi9yU5ndfVDmvgRH1xqdc012HCWdSXt+Lf6F4yqxJqAN3q2x
jDevqNcRcGgf4hSe+jzKOljhiNK0NcUWb7uqZrp66TLS9t7uameFhZ2HYu26ALGj
woOrt8flSb3rxHd37UdmCD2f9ysjXfk8qlzIksx5Mzcdtba06JM5Rf9uMz8xyctM
YuhJ5nfQQ9nOnFGldv7/HaPJl8paKKxMvHhknWfYiaoPrvEz+ajH9UUxmmq0+2Ze
1Wi3fU4CViHw9jP134AUvmBDpUd7o5xzBWCpk6uPCvw9avI00Z3nqb89wygt3cJw
09nYyOSPwZKlzKQ7aYPaE0wk2cUiNGg+tx5FaSblgHLBQlz1RXs9qtBXf5nNhX6u
yNYK6lvoK0PfMDVTW/lMZm1BhzKa/C3Fcojh+ulnZ6H/C8qkJyTExHn/bLzpLDRq
kQYcpJxdEaplDtIDGxEBwa9ERxeuM4+mHQ9oKMWFmO4g41hJXT/nmkVJifjeumfr
FPTTJh0SxiOSyrl6MFilFeRwRsaaflq52gbhAdKFLlpWGj4Z5ClEhQ8tevOAQDa9
8urQKu7ZsCKM8Hn3B0ZGWcmkmXpFjLp7Lgbeb6DISxJwoKjStLFlbvJqCfWScvKB
DNA6Dsqmplgj5njF1Db1DJAm7/ri8GUZ43XKs9fsihidd0z6g8OdFDkUyefr8aFJ
cwXLpL3aT4Om015p11vwdjPV3irMvsoZT3sKyagHd3yaxcubAmtKS14504jfGeHh
rHCLqFjju4XxjuUvu8YVPiAYmz2zwfpbKTXqoHVjPLVH69yv5pltJbiaWciGo0GU
i/KmEwtl6M7c+Uc8YKeSn1bbJD0h5HX9tgZ7UcaeyWJmKS5iTakCaDaJVtKsdgE7
l6gWxf7uY49FycL7ds2z+yTKIyrPlAC0uE45GyyxQpr2e6n71c1RwcUP5itJ1659
qQLg9rcAYnQd17Wav+ji0o3vBUb1Q4G5qwXrhMfV7lpjLANZD4HpsnTuuHYLLDhX
DLUwOhnE+hzctDNhZ7jMKBS9ThitmdCIR+0Mk/a1XEdrqLN6rFcTtC6jVt+SLpz3
2e+ncvI67WTmfSAlgKddOgk8gIzkhy2mfcHPbPYWBINqgnfkLmE0jFpShqmFl+3u
Zj5SoCArQfLDVFnOzoEZ4c/00187zVPnft9l/hRyt3YRZw36HMGO4Ok3RLurCLGY
ylPxYbsH4Vi376m1nmBrvRyKSQZY2AFW5O//tJdSZbuQq4Hod3a1kUAvwOYNiXrs
k4KkOYd+r2DE54g3QsRKILWr7mW4X4JWz/jFuDmRyIZPoDuTzc1dYRIh8pHF1TDL
I97RJkSLpj93fVpO9dk2x3OV/wv7U1q4BgzAO6HkgufVnsrydUiUcimQN+v1ERPy
XH1ZOpuQ9xq4ESBkvrn1ui4oK8wRatofoHjHIm+oDghLXRKkjOBIlqyStE+/9CpQ
0aw+es177hDE7Mej9iMV0Twuz5Q95vL9sq4h9tZ1P+uxu0UDLWjP+J1u+CRfH2g7
Cr65Ribujd5TawgsGu4f4u/8r1vGxqsEUrDR+bWJ8ibIohG0etB7do0lyvNZN7Qi
DTKdqrYh2haFo8Fb6n02wkE0watCxHxOjeCqoWTatgIJ4LVI2XfpH++V+SLLlgDI
ExNRWY5YMZCUeV2Us2huSaXkOQWFRn9hMEJ12V2TN8TkTUfrjxalZHKA+ZZqhaCG
lqTOKSmysaBVZ9XLa1S1pXNY+0kBYerp2gatnN+7nrsgGvi3SxPyAehEgBhaaNzI
6VMt5X2lKm+hgbojimsPJmuXd9451jvz2huF12WLXbqky9bvy4Ec0JYmPYMWiKvw
26qVvP/0NGxKxy2XrNjKcMPhCogqNh1RKexXvDs3USWPL/EkXws5tqnzgpqXVcpc
PCZ+OPVVc5Y0NM9fAwVEaK4/SeakyHAurXizKZz+x+nFiedQGdoRY6N9DHM2pq0d
Bv4OxPXmWZdnqv0bHegkZtP+2fa2dxsSIEOB7VrOIAMcsDXjwfnEmMITtWLFmiGf
UO88zI22BPo0e9OM1vJcbd2wixnY3P0prPBmu2sdI6cyy1Jf6bENjIA0DuEN/7Au
kmUl5zXdCXTZz53i3WNt6VjtmsQXA73Qg7QMQgDC1lIVi2dV/7LcPUyWxcwKFKn+
LvjSEYddQ+rVMC9jXe1UH9rkxg5z01iuYb0n4deVRWkuVSoY2XxZ5ETew4CF8Hur
Im7yg342UPaQYxkiZl74wWwXdnrxOKYrOwpf2UhonOsMWA4Fg2le2iLa0DfggZHA
7/MvxhRibVXsjhjYXvFnQpwzmYLOOoOSp/QGMudh2y0k0BF9zEoI5AOP4wvivDYC
bYYtqqWadr4AUfk7+V/oRCfcHi5slq/S/mVxWukqNLSwKKROWv8q9WPp+ZljyIfM
zRetegnGsRUSkvJwApyQexSOHyYLeVVr4cYKHbSDYfc0QKlia+yJJzcFczb4p4r+
25h8O2sgANI9gFoZGGjzx1lOD1ga1btYKZXR3Dvk9LnH5U0AoePr8PJkP7yZ2ksZ
jCWv99WzeRFv8pwlQg0X+Brp/ypU2MmwrWiVeJEn/buiRPNfA1x69wn6VcCGu8ge
TIr+CuVPQKoQavNbehcPNh3HEIBN/yKMdN449u2USILgBLMinSjZnT5DWt9s/iDG
xu9VfY46dKl9PeyrsghKlvvqAMi96rQ8wtttGG0rjVznZfP46Y5l6DOkWKEIkibt
fisPeNZOzGldeqOKGDf4td9MhqsmCmZno+XK0RGo51jDmbSf832bGPQSWXhV62Lb
XGG+cdZCZdNyHzQHWGhGhIPZnBqV745rdwuUMAcMUj5pIEOL7CVwziLYV7dmH9ln
GN0IUwZNOt746cpgRNJajkuSwZ7yjMXzTw7ebN/ON1k5zghQcbTaih1bIJMD4XEy
6L3XC7xm++fUiEGBNopG01UcFRkHx32H6YeHwj51unvb7VPd/P5dtNzZP60vUwyr
5SujOCuf73Koklgn8BrRbswdXVPOiiitcIOMaIwv9ZhT03l+E48hDxqilNRhGbtG
kJkPxy9fUEkd7dS4be/Eay+IZuM1H2NaeJ54S1G7njGKSrBmfTPK9svipZ/AnKmw
nYKsPa0Rlc3QkHiLHF/JqUO0n7UB1aagsvFI2rX3seZkpN+OxlUxBEld8E3LWnpP
5oNP4JAtOdIGUUJGXEWtHt+1rvksu96h6tU88zEI9qzuXNd61VvO/bDklYm1JB3b
q+1QYLIdCVylS3+JkbBOjk5njCSOj1ke6/ibwhivglbHnyu8RCM1qogCOB2mAE+f
FURTQmGJo3PuCg8O0M2p90aiNhNHeDV/FBZz3qgGTQ/itCXoKsEUZxQa8uKvj6it
1zPNOVbUjYXQpZQCKT+HxVK/pM3HrLS0290QWUJ8SQ60kXkdrZ+uxS4OAYY/Di4s
SJwS9/if3k4YRFV70Repw2SPqQBVwVSjSTdbVgas9oPbtH4RI2NQpMoJZlMj1feA
0HjhDZ3VHHlNuMjnzZa7xnA4ZjraD632k1Njmp3nijdsCHz0sgG6D7udd47aQ2V+
k9Egq8dHRfNTNmsq01VyOUUB9d3e1V2CJr4glHsFnQxIZiHrIS266u++omiWl8Pg
uUTAh/mjMQBr2YXRfwN7MlZs8VvJnL7UguU4u7eXS2UxmT0n+X97LH5GoOpNMQzy
SRaSLZh3Ks1IpDmUya45TLWriyJI8DvQbRwJUIDzO1WGmNNykiU28XE+isPUf9nF
yDzEqf/yEzDgXROYfG5DDk92HIn8tEuv9R23fE6Okwz952IeBg/GDHuKNcBVKLe/
sRylb3p4dfEWumQJ4zHxq4vmVgy6wgjfpIYN+N7kOtHQvmwQ0aw5w7UFWjYWfkcN
zcKByUNPFf0n3HNM4IXo97DHUXeafaYeUF+Z+sHEnO8Nnr4aUP6hrnRYjR1+zRAb
M0uMJc9f8uY5IRCRBGy75d8JbNPVL9hgd+mTLFjCkX28r0KXoAoBju+DnxvbKGY4
S26p+24xMsX5zMroigIeqmNONYj8lWAApuY6eM6mWyDII6D+cYGUJ7wH+JCJn7Le
RrMG69QrigyYaS0Mz3HOzJ+julgRCsZNfFze8k1pKMEnuLtIjCExGayXEggviSFP
vAuO0pxQY5z0ldLuJsWLKSyKLitJHNYFXVs1mOj/Auvx3lZdoQLIy/C90jq9/Be5
TQ1YF+8SIbdtUmrqNyhSB0lD6/NjGCRt/GSKSU8ZRWQjOKRt8Aqisjk7tT8d1KE5
Ew0kWMAhD16ba5VfcqqJPl/4KSKzt38XSDr9wBkAlxljkEyNwr6ZQUA5TnZnIGhs
lEdPxcFeR1mxEFZwf6fL5rAcMgD6IaF5Q9QpcWfyNr/L45Kri+uAfaLHq0hLrlRU
kzwLIhW3hIrD9irYZDIYF2D/XKk4/E71J1Cs+tTCkR1Y0qivB7ReSosKWNSKiOx0
9HW41YwCLl86rXO0bsJhKMCq4i4L0ITJDVsy5heHb2wxKu+bC26+ap/O9b9n/jW9
CvghC4mRr7jZkoUesLIvmNXDu6DlLVOS6S9cUR9lLCtICneXJWd56bJNvkL6ZaAi
/EfnmrX5cTlQBvqMA/FE0yADxGO7Yky5DycNGYRzqtGw+H8XSKyInMUO+jQLDGCL
RGCZ9sO+I7/9STmUyjJ4wsxXh8PArZ1OAWWc76vSUbJ7O/89szS7NhwrNJePUEG7
+LQykKjznyLkTJFyKI58Xa/3f9MHW/Mq6HNkqHwmxdf4djm4JPtsz1bb6T+iYKIt
/Lq8nxFb/lKlykOyStUfjhCiZiYHJJkXROa6jEAR1GMj+55KkwMEg7WeHdIz3EnP
nDELoe4bLeC8Cy4oAHU5KTdWJAh/tbIUGN7AQn8Q4BFHYjxh7Ok+cuBdd3XoVhkW
FS2EG+eM7h7WpFj3qHyVP7I9lkg/ZeTq6Wlz2ykIbTMQeMRoNb1ubY3VF8PDig8J
XkPvUQbcXGVmOKKtW1AtBjlUqI7hX29A1FoUe9TM9sl2Ifz4EsNTsilApVpINyFC
QHJ4ILgkv6TXTBGZLGQvOb7h+g5AKKPv2mAX2lhXh1dKBt4vNfUXEcprDGm8UHVx
CIGQ0c7GBjQYr7P8uu2s1LTb5HrI6BXVUuuf2xM+yCvYRRpkTdjgspNAEEx32vis
zAWS3wJazdAK4r3j6JBcltc8zKcOzrJIxgdbUX11ND0HUjORL9u2KNHTrmeJ3t7j
DZgQkNKHddUMbBslmkOgIlod5hE60GMe8pnZKQ9C+VDD5C2zxIqA40wzIh0ocjaH
E0PbaoLVrfZF3CAAzQkkS0aa9VEcZiMKtINntYMo2z22KNnSGvMcXWsGN/iV0G/k
FRGpeaiJknCP9xuDongcriu35ifnwCPiN4XM/S9k+80XVtWzdD4tLUPbasrDyuet
oGc6Tc02y2JnOHMyqA23tgLWiuof4U97xOCdMcIpS7qE++KjAm2GDM5Mc7sZHLnp
JvTT+38xgTVKAkyiuUVhPDpKWaDvOmffoC5dV6aY5YfzLPCp8vyz2op47XH4flBS
N1rGfXtMjOu7vipl7jw4uhiy+jxs5KLpNUF1uqWSNBgnk0rrjWCtJ9OOocUuzoUu
mr6iSpDJ5bKsJ7WohygMzSFOJlLvN6FnKG/DwQK+e+cf8C+2TZ+kIpPEuYGlsnn+
pDUjzeBJ9yXoY2pGva16+dTX/UIULR4Ih9BW93mSxUWa7z5jEM1DafAPRQLRCrkp
cNsrpO94fjjJR7NsxNDR0dnr/VX4v+Wh/rXufmgY+LJsbQi3/z0X0/U5LjxYy1Vb
V8YWYrhZULXAlghXxOHk4/lKs44LtIAXrL4Z4Y1vi4T36+bbINGo/wycgHoNUkMn
XUaXUgTZV6SeQ9M87Dbly3Jh63gIHp+VI81h24S9EV736lWv7N8Snx1aXC+EewUC
oj4mxxnFi6OJQe6ifYh5LyFvcCRXTWzEtekWt1dPyw/pQPY++gpDUf9JJUtaJsPv
ThDc2+0dM+IsFMdBhcj30qV/d4UqArz8zX8tkwSvnYMlDano6n2lrD/Woh6IaRui
V+jsdcgEZMOy2cgCWisbGhzkHZbS+dsRG1Qx5qQ3kFpyxIMSgxFCTB8eU4kW7t5P
jlHgvCWCRSpNr6f2mQ/XVK9M4U24vqmvqvnE7UJWSAESjJ+1IvV9x/ylQf3egsa1
FSuVLjXRfXYsaYFgXl9xzFB0K7XDcc/RcmUj7HofRkeCxYWpm1drOi9rTBKBEltm
tZb3aYyfBDAkqWmm9i4B3BwaCSM4z6xd635IodZaTXuOcwcY0Z67QFAfq8ba9O8a
1SSEyzkEZrI/NZ1xPV+c8WVrW25A6VOMuAnolrGcOhRCtznxO9MlvxBeTHnOms01
nzuT7yTnyi1vPxeXwexknYZgrGiz5Il5O1hTVyalmg7R+MYi6xu7zoU88dkv+98d
hBafLWigv1QEex2bBrLn7nRDALHUVvwQ3UUo1TDb+nzISRF/et0/nri3iPjIFl34
mk9rRZa4E7t39eUicnUYFkY51mC672NNoFr/TitIt/CQnIF3iEwwm5yeWIpO4iPM
gqBiI1BXhlWJHnMrgsNeIZvTlJ7pEto7UTt738vWDGz//cOwfHveYL7oOM5g40/V
9m0TUhbVEkeJJALvCsC5QCgWa4dwNdia6JBh0VzNXRNZBzLRr1afgkItBaRAWaxL
Asq6bB7g7O0H19ZKB1ouoscc75mZ2Ny3ZOdXNX4GdsiRQZ4O7yW0Ebzpo3tzNHB2
wkRIO762Zni6/AaZaeRyuGxxJj5THM8oKACQXpL07BnwLNZWQZ4k/qcmavh9mTnf
hcYwdhSqx2ScZvJ5O6sCukCLBhgvfUw0p0JkPcRGmVq4fmQlieLj7ZJif1U5MZEU
73OtIA7LSAZqLIVbG8S4OooCF70BGMgOsOUjQCh2ZoYUNlP4eQqxlYHOCGuLbMRj
PMVl4I7JmnEUxuS9B2OD66sndE+7UETUBmZCKUQyatFsEulLWlDe1okNY1zD/D0D
plrZLCCajrzi6CVqEKBZixG4SQXqwtbtalri6/P7GkesgquyFqpIbs6zned+6qp1
mG12ug17uASCe3Thf335G/FmAqkUYINfLOqgrzlRISi+O+bhRwaTkUabXN10Jb/U
joOTza/xvbzB7XDcWJvbIaPbUxkyhb2mCPE2YMudJaHf6NuP5HN6GLdF9KJkr9pq
zjq3ZSLvfIom+GpqPc0RzufKbUBk8yh+X/uVWwfxBdy2U78Z5QE5+9mQ7kUQzHzb
VnC7ZBqsYbJCOsqxvvfLzld/rWZIn4A+7a6+t0ZlLWziE1p4Z7GCxKCgUPCzMGd8
vZm4526cR8CcUfESExhN9PDhM8k0I8kk/58Nwd1RmN+Bb02DtNqPiOypu/uXN2rt
F4v/8b9F0573YE6udtynUmRCWfiIlqn6cq+WXK2R4lUZ40qcwq29R09FQ5ybIZbM
fpt6ltkTtKQSoOaniTqNEIZimvnQrMGqg9/H60vYnPLp0mlfpAM9qDiwI401Bwrv
+Xk+pIviBD9vmA5t4aOw/lLGNwD+FgKqk0WJZGa9GH2WgAiDWFTld1s7+CUKzcQE
nvo5hfWljfcYQPfLCtmR9BOYkEBs+3HnYDTroq1Vd3GP5RZ2AJS617KzU9+OBYyf
MkFu8PpU6zJxZaMSfGHbQX1muOAwJ0b79zN+6TFqrYAbhkD11BpjjVptnO/Li5PM
GoUH1Exrke5s3C9oiyMni9bRvh5YSB0bCWFZtWiD6uOX28HI/U+RlySeS2jzG10Z
JBAKNllFLV5FwF04+JSlwzTFAHLhPdh1r64zE+Cnmp2W5YS2yqIhCDE5QWOP2i77
P5PmTx24b+z69UH2ufGGBpZR38lM1AVNryZ8iiQkIgMF1dvWk60YXy4PyE1YsJ52
uUcI2vO4x1bg6lrckQgklPlYORzIjYsRreZtuD3+98BnUgjvTCtRwI5iv+4m9xfC
qNuewr4KMHL3tTifPNgt5bgCeVOmMS7mYmvMqZygzgPTZtey7je6BOj7LrNEcC74
oUOizEdD7+I0gMoygA1AMRuRSGwTKqrp8PympZdfx70j1rC1QNvekCPt11PKmrv2
3n/s9lY/AhZB+Z2vzGIO/3UhNSzVZ5Hoh0OZWedMS7tTCzvsKI1tybJY01u/g4x7
vbImSGL7c+zTkHhRZGoPEkJK4GP5w1kIwr7dWX7X2CY+96Vjp6+DDpGDR/+qd8/+
zTik3eXKBr5djcA+CkmVNc5/2hpUipFr3i+2AEy2vvxx0muwNinOa97HsRU2OE6M
JEnXM/X437KpoHF5Vw/6p7LWI9V1DS0X9nPsgBSiyXWJ1ibxfiqhpXSL+kpHvVjK
+OPu4mtYN8CbhpX+tSnd8RRkG5+W+3cyCbVbLd/xrRHbvSFf2K7ognOOCnUR+y0G
ybDXfI42TfjD0/e/SJdnAjB9/Q3Pa1SAMKJ30X74lbpDsjmm9AezabxLCROkDJ0s
14TqHyJiF56/tCJTGuKqkNMjdBGVLDI3YvmQ0TlBkpFZ5Mr8j0TPFb6oUraz8FkZ
ZP9l4KfDIZTCHW2lIESTUNZG+F6pgqTQKcvE3GLo3l+2H4rbKBNbUNZbrfoxX3eZ
5WF/8r5wNlZvfWQ/NZ8tC9ATcIE4n5x4XcaUUeR4lrbF/Q1FtbrcQQVtT0VKWKvO
xKlOgi0G4gnmER1aejEdn66DMyCcjvH/2fvbiOxTJVtO8/wJsXrAhFkLB/YU1UX3
6dVu17ASR+X3gYENyxw6axsSOVdI1CPXXPZuvpL61tfq4Em54YEqG3uha97p22gE
jjP/SGb4/F2vVyUH1ZaY1Yit4Gt5L10fTraXN1/+xoeo4umjdvZY2T4KXncd3b33
nLmK9ypxvvnAfsTBxFziNUoijAJ3utERKDbKWuBM4dfOq/RqyMdK1SB1W1Q9NGBc
qRhnv0A6zBnDcxYoU812aw4jVwnCAFmFkLnCxuJdYd1m+FNmiyma5mxab70boOgU
gANE8I7zpoHu77qfV1CeVIdPJ8zWdQxmZkphIlUggTwSQEoMZLaSDBlOwIv2Otcj
DXXEV7kifbMG+UzIm4QDAc37tbO0Kv0/r2tvxI8FRCSkg5huSuWcA8sd5P7QRb88
eHBlJaYMJFY/QTOie2WJXUsWcL3aRr5fOH7TyJkCC1XJmUinwaPQMFkpBp1Bivn1
s12G0P5VSz+uCpLBWd+FXYnPH5G4iW/rASHVig77Q2j2FKfLpPmKzwBjG4RU1PQb
KmfkP4n67/gHzUR6PpM1/T3JStu2H+nBg6W7k4GNUsYljaRelRBf6DYezzdlU5eM
xljp3Teze/X3WL4Z1OGCSOCrzIQzEDT/fZ4BgCkNLtB4MIvhyZp8ahRuGDDpODre
JhHd/Zt0TGI4WAPNDVPFWJtCHeUJG1kFx/MMwlXiOm1Rqr6pPn5hWVQfutUj63ck
f2LicUQ3XVoBxy8TYJivr6V6qukgBl0iFCUFRDhhPdRxz438h+OlwZAa/sOfN3y9
DKl2YRV4DlrBHhp8nE3BP75co2d7FxljRfGe4BAEo+eJiIMypKnPP2qgUftFuHJh
X+MKiYwBWI4FpaaJeeBLDbhItMsld5nhMGZK7BK48lTgRyhRzUWM92uLTVYzxN4V
cv+WRVDbjqQe64f7BOimZ1USCqdlN1MXIOBcFiEeMjl/OmvIyYnGouN2YT/2MXjx
GfhZS8c3syJzZgWsgBAleeHKtpvo7iWLoJKPmsmpLUPU6UKF5QNUvumllVycyLPV
9aCuvcETB/igd7eNz9vlifs99e0MjkS0cc1xNtleo6C38SeFSRAb+BTMII6gabiQ
690nzOEQZyb/exOe4NluZ3zIxwD/8ECoNFBXAgbukpWa9mT+5v0mRV0Ck77Gyya0
wrG86oUQD0z1NXEA5QbCLhbyztD1LgyqyPy9sT6juk/603a9yT3GNcjTdVHNknmL
hwZCG4DrhZhAyt40VgkLWOy6g6rCZUYesOo3yN/58cuLzeQ0hqSAsfTakdaUqGlC
As5RLLifnqjz48NzikxWe3tbZRQqnEyQzkZmbNpgH4aGqQE2KwLXPUlnfFnM1SzM
7URCevneX/KHk3bBLf8qPC/2hI+rGub3Nmy6/NL9Z7tpWGdEhhvE6v6BWWHh+MQk
gxtp5tAY2P5HSLkbx7LADeO3lVP7UUcfdqDhBpq7gQ0j5WJ26GC6jcDr7zGyesx/
aCTnqe7u4YP5yAnoXNlFhRrjtb65efGTqJSAV6NDOXWRKo5Mm7HRwaXGPk+N8xqb
2luVXKyeiWNoX+gwcrTUqUBWDVo7bOLkKHUBijd+qJUGhTDicBYL435W5V3GkfXV
ykhuvQshfUiy3ADkAwuwx+bC6t+ZqrcL+XpgPIHsQUCnUvOaCIA1Kta0i6oCgSdZ
x4hSkxvWQu8C0pFVAz03wZH/PZeCfUk7ncCG7WjF74s++5F7MeOP1LF7XMj5HNIJ
5Z61arVn32Bi21gipowbwHYeLKW2sckTqwuQ30zWMfXR6zsurmCYGICixy3t9w1x
KBM7dU2x5Kuuyf+wbmjV3KsVy0dr3XvzLMYEJm2e/NLb4z+Eotg5lM2DCqoaMas1
j6/LkjXe85dW1D4SXotEeO6r61ogcoJL6KrZH940FOkM1MeP0JypJkzRcKkssKqO
0gdG2yywUI8zmd/di4QpSxR2UOZjucJiIwI5CrJJyGH74/Ek1c9jDDGK5ySrP+TA
S4BnXUXBsPR7sbFRCMnaq0wk+UoTymeC6grcYHARfFbROIuKm1z1aJTJCRq2Vxyz
EHgSrijFnMM8p8b1Rko44tOIcpKQCPu69Ry3z9mR/9WjLNavpdCheg6/+lZc3y1I
y4HhBQKTXvq8HzJe1hjCzg6tef9UniAOR+r5S40EMVsXq0bqu9Ie6w4BH73T2ku8
5ymFaUOrSc9ydvROL9zbGCQTm5KezhOUwDGuwKBVDAhrEVIMGhiOqvoB8B7antTQ
upQ1p4mb9ePRReEoCaTZy6wlOxotQgKYflSEfEDHcbY8Dta6A7lAlJTAPfB4XVQM
kZKZ+pJw3fhR0puW/B1FkMNKYfoHLgHn2CFuAq4LXvKgxMaByM7OSjRWZbppbv4k
Qp9VqCUO84Db2kgzvzDpBsoTfvtWSDcYCfh1By11C2Kk72S6oUTsn+CoFOHIzG4F
0ueJUlUaCDYkGbOG6aD2VqTuYImGtqbCm11JWeEc5KAF5p9+MRJmDrpwfo+npE4C
37jHZteR727xtBETsQjsLxLlEDWtUypfaUvrlmmjmtBjLdDkkbCWkVPlDgdJGRg5
U0N8vpAyY57AZiAoN6XvKu3KNqUEDvxeb8fBrOKhnXh0rvfG2PEXJQ4C8tSk0tel
xGr2pR8EIaEAhdzgMAzVjqDiN1r98BAQ+mkjd5YkurscB8I5He8gwHHinPek3wXv
wGuBBGmirxv5WARQQL5SP9gmLdCHui8QHYkDwMkh31oBHwKXg9Dsbu7goVTSpetx
R3/Cbphr0JRy/h/RoCzSpd0Rrd9GzY0kWKeSnrqyi0TBi5S1Ocxp8zvSf4y68LvY
guaURmdfzlSEKuFZtg6DmQZj+6NIHY9fVahRo49+m3WN0EzAeOTlMBNRUboVR1/O
wcjw2mTxSPGaGTfREumM9IjQ8P2jXLrrust+J3J+S0ivhK3utD6KhMT65RtjA9eZ
TRrPNzbz+TFE6ywtNus6GmlhZjrKSkoZTVjAE31sMGyC6Bd/fkaajscijjLhm3Ze
OBfPOTelZG7feCOQrUz2MJvcn6gGuS/AXV8l+BWB0zGcWai6i3yEJzpIdQNRJgFO
j7sLg17A6C1WmsjTFSps4kfMgUNmhF0ukTc1iYF9EdNXPmTDaLK2uMy/9LI/Fs24
7T4ArNFoQ5NinpJqNp6kVZk3KVF6jtsM2Boyexx8pNX82NleRmUtqzYpbHye//mJ
AZrix32ZiwTvVhXA+KRzfWxMNYxw3Ve1yIdybXBYySZ4L2Bk71ikoRjXvN0AFlgh
N2Z7XcBeMddfFZy05sRR984IJT5MpzgZMLxDsTuNGjvX+SPc2m6mjl4QqWNPNyxb
yNkH9qnLRS+vzx84UmqEYv8xmaZLiU03uJ0aama0dtNrL6HXY4XUu9+rUhcT57Zt
PS2ZazSewOkBtkjFcuWvErLM/ZnNZK0Qkb31Eojs4z7J0GVN0GKg/Lzu0fon3usB
xIm3o72GZFtUsGK2hmQLYPnf4J/TykMQRYrr1AVd3WkAYj1gaaGAUjDYlaPWkLat
lskRWi7fQFlENRMZjok6QMPTkceR/HzcineNsHqYWO/peQBZ+xiyezrVQ1cjDbVa
CZydBwir/pNtYp3QJMf2E+uTnUxU42DNaWR5+zO4olPAPMEs1OfXzEpxfe+Bn7Ur
b/FK3c87HhGodQ0KLWqEZdbvc22fvTdBw3kXOs/rd2WRy9myF7tFOhpmKmjYWwes
t3XXUHuaskkc+WnJggNtC/MLWF+1abMCbtqKVoQmFEGhjOcxArzVt69Skor/Ruxs
Kh/QF2TeE4O6WT7UgVS7117C+l9piYzVQFzsb2dMtJB7hVLwm2QpISUc+fRYTHTC
sBhpChjCj405Ba5g/bNszKIrBbqd9AZCkYns9sMWxahgXuHt076ZEgQWKKIHNuAk
WpnjnmFQ8boc2n495r50QJS6ciszlcEmmB5gOHWxsE7GyO3ekN1+3BFAeEJplZx1
49qhbtMJHwzXIFPQfwYOQXuVqE2BmUQPJs8rO57yFRugxx8gr409VRTGGH4UAnRS
ncwtou9jevZ3YyuBDqt4xEoY/tm9jylQOK+gzJ2i0yoLXQxaNvx1EZd62D7laIYu
JBroPyjea0PIDkfpZqDgX8U1uX/TnzkR5hS06kxzLJ9GCUP8QPa1kbSqb6LDSKrZ
D3hNjPswh5d1BbaFmcQk4H2JxFoyBgkXmaTy/eXBk3SezVgOdNpsPZrvDwBdiOUo
uGObPUspwLEB3CosvRnvTKEteG1fYL6m9bx4cbLypDMcuIP+/M47RSDChWYHiOiz
A3Oj/xiRw2rA5H7v4RjJld1/G2xsUL66LahqAE+SjJLyq8ZMUo3wRi3CZ+RwLatL
oshfENotZdwRgalBs44Vh1rm/tk4K0lHNZwm+D16pzb8wCWQ5HxVRLXyvhFHoHs9
IPeps/nA4pkSWNXZOKqkJR1cQAK5Ew8gW661fwtBMcF2+tBWzxbIppo+9KfeqBr5
x8wqLGPx3e3IsTyTTof//tJA68No740LBLITnGJkHrg0c5H8mNGSuPSidd8OUKx5
f3r9B4GTeO7KJPzTIuMk0FB+6FCbQUwhNWNFKW4eofRNYexBt0u640MkHYmgTOu6
YHbIbs8/lCsspKxMmLxlTZkfCDFjpj7zjB+fSgXnMZY7K616f6dnmNAR12c8s4YT
EDi1I6E74Tgk7JJ1/s8ZYJxo22+tvovIVdSDoQccgCcEwXZkcX6kGMzxADtpgdjJ
UQpo9Kig3llVFwwWZnnYX+X2nVT8W4qg3OnIGIw2xWH9mR4s48E4IGjhmYCOTXOe
rQ1nxKzIyPPRgzQaHzgA7ElVaktdk776v/ak4HTK8TUiz+ZwvLPjS9HggnklEWpc
CEwkoiTeerBaad4BS6W6YKSQLq4FZuLZquE5yF0RW4PZXxfIQ7r9bK/IuJmMoVbQ
lq5em07ASMOps5eztMEuEdIcE2efROrOctaLXtRyxLpAB0Rnq2+yqrZdXOklrY6a
OecS+ybWmTKH0LcAOOIJUDp1wOMt+ZqFhTKx9t1OAITlUlQ05P1oJphF6HdK8L/1
6iqnQBHxNCqSNxv8EFUd0X0ihmMDiRF/IPmCgyJJ0eTi1gQ0MgFTHKcrSINMJB9S
YYe0K5yvJBfxqldmOgAbKd1/Xh4h1tODEDIeiBDxflMAx/0UGmGaERF82AKtGodI
BjICBAT3iX6Ld23+tWIOJs3C3CBMcIel8acBwRuSLqRcxent2YJLZomMiVqvKghb
IoFPZTCD6AXCqjEeaRJPjWu81W/xJO/u/EFSZSrDfmxYKd61hs1UHf9L891JX9Q2
D0wmNwNYGiq8mQnaDAmTsbNDX52iCVSUoVcbJcx+0MHN/etuEoO8fZS9DH2Vs3tg
NGC8qmkaP+Ji9+2iSJvEbjeqwn5PoN4DJc/p3P+/8PKDrUD2zYNPhxteeErrH252
40fnRVghu5BOaxXcmMGbztbx2EHDHq7VpnaPa9CtcTd/8z9713EBA7VtJ8f7LdIk
uJEpkSkBmYoO1accFyHzKkk5tnj4TNeh0jNbxAwsHM8GqwrhU+rmoEPMELJALOWw
q/Y9Y4opa1VfDsmiymoCAT2oJXP0v61sH4hi9gCnjENInW+gTnrnxg8bYC4IsHx3
TVEnfViKWSvIPggGT/yzH5Grv1lT90yUeRcB2sdJVn3CELMTDZDQLN7gCJtdITLi
sHb/hIN6qXqUnm6zgRUxfzFbF5yWenDga35AzScAccpgCZSD0ijG17QCVOQiXreB
hFf4kwFImBoofchhfW9JkgAIlfhIlYMa9LWD+yFYIqBzU0ERueF1WOtN28TyrsAk
9kMcFbeYX8G+5pHzsG9Bskq6/+OI3srpbLJgOCADIku78+k6JZ6dzw73736FzuHa
0KdO26MyZYNq7BHsdzkNDx3EF7eUFBwxhdZQKO2+BSjAdZA1jmBAPjRtKRz+Cn5O
cbMAR1aQa2wA8YCg0o0xEWQ5E7d4/DPMYXtVT/fcDmOC5RyRQKt9/yJs7XN1oJwf
J8TaiLDkErC2dPT+aQfIuI104HGwtrKNE47jfBN6NrHzmv3y0gZoXQkzMOLHGyRr
3rbNaTRBGy0LaxcyXm61CC8LKbkGDDo3fC7DBkN8mSDBjI6KleApE0BhAnxtAopT
KkiBYSXHUVLlvnBKcgiQMsm+/X/jWCZChbxCEUuQ0pIcE0cYIbHJPOz9x9s80b3u
VjERryo3zEWp227629sjHuY0AjbpVPGuVe5kKb1n3jq5KES4xm18ymb5WjRDPpyy
leYPzCodLevdmbOqd9Sxc0MNRcrrrMhaOSK3SwOJAZIR8QfgLw9aah7TlJQVOUFT
KrkdzHQVl936A3bdszKotrYdtPOTWJfccaOd/aU6bS0j+VWv9BSmeFfamDuhc9Yo
nkXB4KejvZJVEtJ/BiiZJBGHnFbNDjNgF9WAM/oUiHoDTxciMZjWSFio+JVD8fR4
dNh/IPgtrOjzo63liz3yQ0mxG6caQbvS5h6+lro/aRGqeiRX5NwzUcIpyAIqGuyH
3gLjQRg5rPocS5SrboypCdcM7AXWol1+wOZrVTgN17IrRCxb4QHTFYTf8aeQmLMl
KWAoRJ7MtjWMm3Zjnnbfnhi0ti4PM/Ty2TmCDtp9cWkjefz9jPIP0OTko2v9BzFu
NZnPAwTX/V1URkRVpDhDAeAbPs+Fo3bVmAXpdRHAnvwk9wAcqNEq79YGR00k1vKm
THeS2Rort/kYKEc5/QrzpUrMG5r5GqeBvM8UnBpEEwitdqNls4RFbv59/SihuEQ0
1dF0gnuOdYTCgfcFBVwl1mFCxg+dJOBJGkbWd/foBm7eQlRWYMyAbKTUerBtsobs
fKMdz5bgP29JWvvIRE0TfZbjVAniTnQCyskXu8OGuGSArxbKCEA1tFGByKkQkxL/
zurx1WUgEg/A4dgwx+0drJn8q+N0DMldRj4+bcrl5Ft7zZ9+y3Hzax+Gl/HDGQ1A
f4v6FGJaFd1E6a1DII7V8HZGaVoQD5s0DZa6WTSD62p4GFHlzgAZCDN/0Q89QdNh
+SFfaRKqmS89WK3EZfxPfi/vpzeimd3ptcGe5Pdk1eFuy3EUVzfOMEYxH9QSjscD
NqsgpeXmhUXa4rkT5RDbXn5kwwar9Y/2b70g//tYsIkfxzD7oJNSKufTPapy9fp1
RcxX3KH7erPI29J3JsJDYRC84l6UVx+fCqoeanWyOn/R1hWMVI7j1B7wEDLya2wL
CBJretNlasNjrB7ViFv/sCIAmvMj0lF3k1uKfTzg4FSXEfJYlzUFG2n6/pJt4Zqb
E06MSu8mO9udaRZ0whqsWE3VoFe0zGxGlvktGqbBKAEbVQLF9nez9Gud83dBmcer
cqjcriizwDw1ZsS3IsY08wRrABuS5ZZRZiI7wFSps0cztTFQP1Uh3AEjpeifwITQ
7NNVQj2JpnqrZGuRxEmOfpIwlCvgnyvPEpwa0fJTptwFmOgBh4AlQOSo8gUUTjMT
C3TpQokH9u5Wwlyqn+9TeO1is9vNmUuF2Lidvfj3pvFdoHCR52TraMCwRS2/wXSd
sx7ZgUqYl3LSRiBbGdsuWbqzwz1ep5BtTUPNTLWcdD50XMjmT1vEfSuA0WP+xoxX
x6y9bc+jgVzN2DAAaSVlKTVv3LROJvBmChtstWMOjHg6D3ND4As8BauxYTRCCcnf
+xyJnEXoopb1N/Dg/gf6yK2+/lPZaBkOv5mtEclOuKFMRkhEiEZZRFeixnf/GW47
F+m7+68KNmBCItZEk6Dd0QkMOO+WdSJfvFJNnbaWNOqg3Ab+4b5+HfKD1oXPBkAF
cNg+09JbKoLfUM1OYaj18Es08bExyxoWfblDvrK3hQDJrLs24M6bjxivLNcUYvqm
wPI/r39xSAH6QOzTnPzZurPbKV4hsiE9WLa0eI5zvhsto3ecm51JZCU+6FM+nSvK
ACYpBu1x2FFIKvBP4FaG2AidP+9i4w+9OIcV8EEKH7popeEvN59erdUIVQOgUZNE
Ess8gdt4QQ3kK5p5hEpYQtuvE+lGJ/N9+5RJifv8BoKkCCGkKC9c1iBdB+9+fuXR
iKRxSiRgX5eMNgZ+pV5NZhxxTsiP4vemnWljYltoxFrRn4nTe3oCVcs9cgB8vExp
vWTd7tVYRY7cdCb+tn9KbKCnjxxLWlisKSO4U57cG58V2Vull/7sW7Lh2LebPoyZ
2Yj1DpQHFDnp8s8ptfvnyvPP0dcQLKQL9M/GlcGk6MXn5HPFUdYwQXQ11OXo2NGf
b3phDNyI89ynXg2BG4jvn11frF3/OzWnYrzJINZhAsSnR1gU4xqTjpGqiehL+Q0A
FYy2CLCY+kVSPs+oJFmXYqKmpaF4XdvmRQ5KfEuOSWzrkKtTtfpjjhW4RE5hZI4G
/JBD/RTK97Ws+LN5wiIaxnEW88UMKh3pqMIj9+gIa4gtiq/TgMZ/2NnVpzZzrKqv
lacDiOAR0kYtDg5MJasiaSQQv97nekzKxHfMQGmpRONWWQn6k+4cEmkAiWM5H9Ui
DnfazWP6HcvcvglCgd5qQvm67vVMls1AdmqeISvfmwa0GhOZbYuEMqTcmRzczWHk
SzjBN8Q1dAw6tmjTmBcBSeoGbo9MHRwVC9IaUrSJCGyGkCoJJVn1vKNRK0D8TeEg
GcrvnycsTxo0wy8SEjZWnRXJ6gAKlZUzrLUt2Yl9uXBWljPjAkFFmkOQamnRdhKo
rK5m3+pSXmUU367zPV8wABq6at7gyXHJXW8ageOOlQKt+1zjf5Ep8H7dAupU3hrq
cG0oNcmJlYJVUnzvGOkEjqjA9QKtFyuPwSklNw2H/fncmi1LlF4rOI/8IzLpp+BI
sJbq90gXCbgjeLm52ww88bmgEQQ/QYjjcE3pGwnl8XXQaiNMog9ACL1UTTiThSYV
Lg1KlGVO5wI+d0D3WnPIlKBOOlQUHtEWdpkoO+KKYF07MsPx7OA7nWuhf1HuuyPC
U+FRltBVw0r9pP7A2F+sN9oWibSfNa6yYZgtNlT9rSmtgg6rKiKrCEDeWaRbq4mK
BMJuqCkqPgeqBFbIutvXyL73Hv/9b8DpZc6PFyn7LjmZPiRcrK+HXZMJxW27nfS+
WZfcYEVGWbKykOCIRsTDBd+kVhX9obbrlbruTRqfiARGX1JW1AMoukBRo+DFaY2q
MU/cv+KNGNpZ9WrcXOJWcI2tWM1Sc+Og19jL2w0YFUOOUNRnans8H/SgzHDF3ptW
CU6O5h8X8LxGrDxQBkCm1eSgxiuKFSJY4xOj2M9tkBeydWNQyp85nMv8FJAKdCPT
bvUqBD1rSro/Vqydb9PywtfM1Ml6T7jWYL/52/VpDefqlVBjGtIQ6a4+fNGWCKrb
rlnPQWykJmkn6atyR0kHbOBckOSbSOndYk7+275pF9kVrzWR7HrYK54Gmbq9UnnF
g5vOyfS6w1K1x6tdVFVW3OoC0/8Ha5UIw7vpQ7tVQJOJbJZv2kVdrHFFDUPNAlHu
ksmNcZNEttEf4pYYRKAcqzB/qJ214QE48ZkSOQOjSWaJ1Ofz08yrMo7efr9VGMyn
tCysLg+MqBW9mIbDPdN1EPltPyS/b3fcgXc8uDpikcbe1ruZYbCG/cHCvdKPP/vF
PBFuNbwz2f6bHjVHwIbLqkjMsWGdfdGIlh+2yBp6JvORcEAIYRuTYzS5gsLmgKJ+
yaetGJrNVwtqu6NpnsBNF2cIUyaRWQYkcV6gDRIDLuY2gjM2Om3kofyyZ/zl3Cbe
aZ6H9GeGMfeygDjgHbu/puCajLzzpve1d+gq+TyZZU6yHj/lOyz6weTrRe0S8eBg
cbRwcLLS4JmmOu/Yt/s9JNImuajLpxWKhvJ54Kjt4CQ/3KMSuMgv/QvRk3lOAprH
vJGXN04IS3E2+CRujg64hPRGlAWnlw683N2V/Oh3EvRZvs8Nz55iyagbWUTWiu/r
tb9t4YEGcHlKbyBPV3wKvzDpfaVDWRZErY1YVugCUZhCIDlnEpNM6Qc5Sb3GoHyA
SH1gihHVQQhcBISMAU32fV1Dp6C5OxoQgK76J1CLanpNqhA8Ah7pr95ub8+XvDpu
lpAfWzRX9Nr8yuVBSIWEsqoJqU9Qj4eWTKO6JTBCkTvA5mU7c8eNIxBcbSNqkxrS
SuGQz2b+HVLClZeqMxlLEhyqLtFkw//zT+qdgn+kmXwaGDoL4E46gkKgc2X5D72k
eQdgSzJ9eUfq44poMBnuHHFd1l5K23tIr4hmcLZ1iLFTcehKJhrvPf5cqOGZND0K
13aM2JKHjkckPA56yRo7EQdbx5nPx05eaI6vTaBoAPx/WWuEtfxl+TyYSPvDX2xP
XsZ7zJ1B0Uty9Uuwtqf8Lyxm46BDOoCKWJ4NxuGI/WD+7q8rWIYnpbyODF61RhW7
XXGm8ZUi2MjrGXQIgvbZl4QepK9ymKZMACv99BHFRGSFMDff+iSlhkM+Cdo1G467
FQ+roBeTQqMramyb7hlIct6sdqixkmivKRJ71E5L5JLMq+3SGYKf+tD/CueOeY4e
k5oKTu9ksmyjSIXyDE/gMB3aedawwcXOtDnJCiOFwq/jXpgznKeymGDZ0fkB2ZO4
doHudikwhrUKVV3UPQh0+D6PLwa73/uy8keopvtVEd+DLXX5xwqsYnCYH662nnfb
Ae7m99kEfqc5PjVxb+YGkL49/pvJQy72S+pz+UvhY7wslW3cIGQ6yAKASA4eMHad
2zQUoaJ+RYPo7+FkigHKoem8APm4Rn9ogn9TsE1Wh5ZlB7/SQl7TqSYUzLTOMyyD
S82bJpul8fR5kfzf1+0vxE3yBF6Y7jZn37zEKCt99haWnIZMvk+bKhsTjVlQwDoI
vIfdxE3Bq9Gk/Ted1dPT0LUjA2RkdjomJfdslreocY8QW9L2Z5ES2zgBT9P2nbz/
+5S2IrY1HWexbTCCjDQoxVwEPHEqnePLZRCxBxhPnSwZ8pU7nEy/rv6oJ0YrRhDU
bl7p+jea4z/nIEKtA9izsB9P2XQNRLm63cUh58G/OiuElLvMVkrRV8oh9zPcX/U7
wZYGzeR9tMXE6fRzeKXGk3b0z3RvQZSAnbhpdYzurJ5g3Z+i15pHOSKVwOSMC6Yw
T8nvv5knictFv70kM4MQtL/xjQD4EkYS55nGJpmmOIW+EydUwsQgcQ+9baubi2Kr
35vP0nFvAElv53lU4PnqenGgRkIlrkc0Lj+A6AlbpuP40WZyy2vYwQQIZzLU+Hqq
o/WSreGiySf3k4oyWKRVAZ0mPEbVtqCAiQZcZx3ILwtvpqm9UXk/YK0o0B91Cw8h
9Cj4gAlf5FIIwqV/jDLZe9z5c6uRcWOyF3l8ekZZ1dVOKUzesN8/WQ/km83Wk2jf
CKR/oVNY8FXWHmHGOxA0ffEk/Mdufp94YGSwBaHcCucByUNwJ88JqDuil1CILGXS
GeZ+QH/9kVveuc23vZnLvqcsnEVjQUK3X24/EGViVlpqQQkIYQuW5wzU1P2Nt61+
gEtMfd/jTyiGvEp1aSlltoigF8jFRlRHeJO0URwqn0x0M+xOGSWI+LTQiDwtwMRZ
o+5wQiu/giXrODKgEJT0gm7lMODZtbAbAFgxiw8d/i7En4ze8HfS6CmvyXBeafq5
JTqCsXBmu0gs+RaheAohjv27fEVeXARkk942RaHJJ0EWkBn72koqGz8KQjhtYklu
GSZKfPUoO9GeXTjpu/w4lRKbN0rCBbX/ichWgUteQer05zVfxKs1suWMPU4fAxg4
hNlBTiFUS986ndJfQ976z6ufAnfExuT14n+7HhVNeeGWaEi13ApOwGAu65MBhZC9
jTE34d4AzJFOtBKFD5jXEbgWhqutzpdtt9W9CZreRa2Ii+f/fBtnuoBJstj3wrHu
3V1ABvO8YLP/SDTylrB/Iankwctur+2fLoJOlHTlBXOfjvbUD3ZzR+wxqqy97eC1
LqbRReaXPULw91WdmkzDRKIcjx0THsXAFJOPQuJRFeAZ8Hh0Q/R/dcivlPWbbzFI
q6huCrkM8uxf8dEzfKwX45laiHOZEIoVVXwaDFCAzbjvN7w9nzDw6swWVy4U4jxa
yWDl232HqHP8PNBSNYky9hvhVvtkUIzUOHdEUvGxuwviKGdjLGHzLCAjhp7vkiPX
KByHbe9P/AImdiCsEmnEuWumt+5XOi4BUaMsVN5LpqNchMXlfiOmQA8x7lZeh5oM
JZqDsO17trTq2IiCJdxOCk03VFf7jF1vU+O3zwNKyZTSnOdj3/oWcTIKWC04Qm0x
TxktGelEnvFsAHRTCm2Mh2IHPRQcXcce4oGt8JClSnvBQwc1KzDS+xF18GJra+Io
ucLMfN1KLNGJXbJOZFWc5a4QA+qvBXyHNltCSrtg82Vd/8EELTmzVKpguffOm5yB
eSge3YwyH3yRSgFggd8t0tjzHUGT4qLNq4jfKLW0ndw+Y5ag6umMPifuXzGDo6JG
P9zqGp9Q6nYd+wildfkPDvFj+PzMJezrv0niwnJf2MZj9NnyWzuL0HHNzrXwxVU+
LkN8boUQWKXxzeFWBPVeo/5CPbzdt9Z2xKE4i1ZaswhdAXsDCF/eopUbhktN/GDZ
MKPb7wEXHJevEg8DBtCv96EawL3H1djIWkiXgFFUGWVcznVbDCix+JrA8Sa9Ua3o
sl+fyHdTj3l4YXV/WxB9u2Bdfrp9YdmhfsiLy9IaxrMR+131tpQj8S+OdxxnOTvc
6xU60Xpg/iogo9woQPMuLymCnfmFUPpb/E1gRm8riR1a5KkWPycnADDJRaoqcFZh
BUbEyFOD2yDNsJDvHoAxGjVuj9yZJmsJ1foMvrl6bPiYF1Gek43YIijXBwH+Njh0
efiu6ZcMTlffzGMLi6SWns08eFFuXCQWeiGfKd68r4YmsEK1dxYY2+eW1kY7KYTZ
c393GoIxSrVVyCG0xt8xHuYXC7B1YBdMaavDYgtarBnae/YSwx83MbjEcaH0Zk7q
GGZu2MThhchKZIlFBRZa4oxTwkxrQ0TEGUk95+1MQC4u7mWwdWTqUl+boMuGMRDw
py83buutyjQAOqfZdZQZntPtMGJ3Pn+MwOiPcOrzyjFdZXAojyfst9r1Uozh9kBm
uNTkwjVVg0gFXad6vLIi5QLhE/ThZlDvJ6/66XqQh5SmNOO/8uQuwwh2yAe7WgpB
F1wXwN3ngOFjnixTonfeRfkr5LP0ePGG8Id0riRHuHH4Wxfqz+Y4n8J11uy4bQ3j
cQwwWScZuioJM068KdSSXDr39M8AoTA93pDSZNAsEBGsFwfo74ufKuxatZELLBh8
lRl2jDE9lujhZhzk/4LroOQ/1WrjosCgaTgNN/IcSymIwBO7qeSf2veTb9GtJEzn
fjTFBIoJaoSE/L/yV5kvWDFzt8sSrTTuA+5PwfpvzaHuM424s1yuwSrVqwnrfegy
W065IDl3JPbrVo4Tu+iNQfdHYBRD/9q5pVN9hnwqsVyIl0H1/ccbbKtpNVL5SrW3
n7PDVbOmhAz2xuFHITJY5G7GemXOFldfKK8qIcOhXSJy7zrBoE4zA5R+TdNYi9fv
XFBlunxLlTHrfDiDkKu4Su81rUI1vavPqv+P2sJ4p7nXpmXid4fiDWg4Lj+BUwzJ
1g1Dxbe4eqcuVT+doZbYmAxgQTvbfCnHH2rnArcrFaTO+XEuNPAr/h9n++vV241u
Y7tYyt8I7HYjvqoewzcs7vwUDlBXG0ohsxUSwpeowsygvE+rbOmZgxn4j6QW2aBv
R4K/ZKreacWizDlBeRQDpBfUcfG+GuRTbQT6juHx3G1wBzeBc7F8igQPbt46C9Mb
eaxIACUdVd0qxslB/w9LL2JsX3cQ1Ef3QrW4DVyMBH1UfrhFgIwf2YZ3XIGfuT2D
wGgPeNUlJg9+pxhSVt8/hUf98XzvKFKk+tf3T7re/5jLsXHaJOokCs4kQdTNk/Qe
AAdYxxf9IqQSV3cLqEZHm+53vxpa+JLeu9O6EnyV2+Noz8ME0qpS/lDtgC5lO9JB
Da3H4Y0h+WfGWo5YiR2wRHmsefI4lrqXpk/7zkV9aEp0VvWWJUlZFOVwpkcfvzGH
2LdsLg4AKVNQngCGyAHd53tncvAzsh6munXdhgkueVtQGBa2W8j7G+fV1fnyJ2SP
KnqCN2jLxNhoK1a2iI/ht+lkD5u04vP6SxvXvGxfpMhmXf73f7O33qXM2g8zT2lk
439sXIoDIuXfrXsEXqZClyNN8euuy9sPJz/tv1dr87uB1CbnJ3XffIajE6ioS+2w
yACQkhmL55/wrXXvNs53z2hwIGxkQel5renkT7FSe7I9nXUMO4Isv4KPGcWgB1vz
JpWm/FQJEUHHNs1+12sLjT32MMeTn/HfWCbzQl9i7wirQ3hAibbyf3Bkw5XnJYR6
y6FVjUEQbRGLp3uOjeXjjZHU+RoSwB5BGgjEtqsbRgYgJqcwwkp0zW6gn6mp5d28
yo12K1hUoNQToZk37nBVFumi8IWTHPi4SIesg+ee3R9ZpARrUTNMYLQNyiDSX81t
Qv4yYILzWYudB0djgqRFZhRwxYqtoe2oyj29l5EcymUxUisQfy+RuRiYd89lHjb8
g7IKZLEiodzFU5RQ4lTgtdun5QFd4gfyzaZDvMnfk+27Osu9BaX1B+qy6PvpHqbQ
FR3VhFZNMgF3juSUl2YU6w5gXWUk1BwbAqE80O9Zd6xLpzYVZm9gVPg5d3B1MbMt
wYVClIqe5U3nZ4ErXeiUpc+ihGSuceQLQopnt/AjXogCXMaEMW8H9JAQzDX5nm7x
Lzr6Bui8bP3TCuxtTXN2Tp5dMmFzZGdh2tYzEPMLTOYyWp47ThHZcVbiDQgKqNMU
zXe5mbdjvUtu+cfwt8yDrO4CuObckChyQuqizh9vyFDMiYGtDt7nS2vm3oXR9oJ+
4/9zju0itdJFm9m4/u8whlWU1wPb17AVl0zQ9mHU676KzOyYuULLkSymy6NjRbmC
/0U3zstkmnumkEfu9xqMSWYP5Y8R8LN/mL5H0dUfsXc37pjOEXAA+syAHXd8RUHq
02ORRvH1/quTs7416zDhlYxJL6KaGRldAK6m8HJe6Hi2B+oWlya7med6f3XOaQWy
jhfSHG3rmabU7McDmw4GPocoY+SnGvHpfCVj4jd5ou0EIUrEk/znT1Crhbmc1mQB
KNOK0p53dcrU7hfsK02QJyucNOdzKcl2DoHMkAYSqzbzyljGNtZQ8JFB1DKa07VS
tifa4YFMpR3HHIAw/He5rpnOujXtb27FxITh+ZnmBt7XtlksqXSJUSheXC6fhsIs
C5Rm3xN0GnB4kGLUE09oge+aQ9p02PgR2Fpy98RL86VuIBYuNYe+C5aVWJecuvAg
zpvywYnMQ/byIcPT7SEAaA47j96zMEYXPp02lYznPheWWliPPxU797AyOBMZNAWo
osc1pS6hdn//ug62yVfwPHvVcKWxRFgvJ/pa4HjtDrG3UY6z9ugTbGKfUJpP/WWG
b2VgnpSIPaslNe9c8hb2CfOZ+hk0Is2nX/8WoLxaUkAxmM6xW1AHRwVaUkgToY1Y
ynskZMiRj27Qg3qai9JTuy/LHJPqSkMTHBfCUMndn5UbmKEYGTfzhHD0X7pdu51f
OCh59PeH7/j3mqNVpljybg5R7ZzfgthphiPbeIi1TS82CUV0wMcdmxLpwxM3FGaW
MbcWpWmqZm8+DSQBAkywM4pNZhBm5NhoG1pth0iIYKE6IErj7ljPu/6GyZseUbPR
M2x6zX6Lmh7MyVPFX2GCtoZTJGGmkIu9OTw2xGv1Ligz11ASO8hkRSarCxe25Mfl
IdshARtLh76neBcf1O+dzPd+QjffqEb4ScuzzlQVKGwxCSTHt45L9bw8N36WSNg9
bsoHftcdPQR4NcavXkjf5Ko8XQt00Fn/4BrbjDFiRNaW/3E1PrW5rjm0pc+fm+2y
b7bFiKcx3MDq5+LA5MsNevXY6f6j7kaUMstkZUc+9bP/VH4npOLPq6077OBoGDmD
WCaYTmLbJhfBs+dt2J7DPjw9l98cOyqGEORUsN9PPX6KHg1VRNiHfvB58cZOtK2e
FxTtPZYY9EO6VhxYiEvf7TMSf0BmZF4C7TGBaEnaVN7Yxay37LgGR5fg/mxOoXeI
T7uyWYHjQUDTkwE0rnSxq2qlG5/SZrBZqrovtLkOK+kwbrqHp4/YsNYJ2c2upBkq
L3Yf++ZhcetJPIZdd+KErTxBLt6zkq/YbvhQydIsj904z3x4Q6AINSDyMs90fwJx
cVKkgyr3ipwfiMLBf+Vto6279OB516poIHAaxbJHv4e9kJndU1Bvr1SILeNoiFUu
KjlOFqygT6UaLMTGgwOKJBddsGbnBcDTwB2gE6wdjX29urBlI+3m+LHJjsgasFpS
yNPA2jeylMBs/G8+fPY7LUwufG++HHbEvHrJ4vfoSopwaJwBrHqZVyjrQbsepU0W
vPIdlx+xQmv/N7zykH9fHQYgIrFgV+5EMjPaM8V17+1twRGVdXvfMxutqNFXUaXr
/L3FYgOVWWI5z1k+Wup+U4OgMVwGLgdj/ymud2ha3yp+uKC//U1jogo2ifynJWhj
em3H627SEjqDEDvHMUstw6GTNU9Ay46QOUBFrlSas1kb7XdtIQ9385gi/s7fP5k5
wKeViPsRh6YrbDG2so8UUC3oJ/FdH2qdCIGAtlL902PnoYLsPgDwFGqCnAEkJdhH
d2qLBmnF6Je5MOOJq3gt0Pk6zKrgIRb3BrihC3R2+wKfxElrbSyPCSX3ahig0xwn
ek2FD3JgkQ1DMwHPLlCfOrCJRdG94mcnCz/WSgE7Pednq7OxXKWJs0kTnvtWTbXg
laR0oJXwRVSXSGI4/fK8hbbwNttYI8/sIwybZxIRSUpvDqOyAKYLx3oDOpPtFNZr
U2BFpdm9IHj/9gHXIX/n0FX0yU86S/3rILXXq/k31isRw8kE8tfc4qHTqfwBmKKQ
DF8pIivHI5ylH6UN13TtHuboTmy6ojAPxxzF1FK+zSRyH2eWhRuOCPaelfVx4kb/
NOPnjOwM8Vh1SjQdUAB1kIaSqbYVP6n9V9ALG40ukv2aH02oK3jUAVe4Y4O+1Lnl
JTzHa0Qed0mj+I1MoVBDyMPrjyYxkc6WQepw2/8rn6Ow+IEQ9ZGUI3bodMRIxXMJ
TMhsRVRbob2PK8x5DkhYArIBDssRSmxtIgtUCV5xJ4MH67ScAKaPUTu1qfUpRpUJ
6DKPgwSpBQ4VSylStYhKsBB8wx0lr3Neg8Ms+pSloI9SUtwqh52nTIQ4ObLMg8KT
2TjJkCC+aqg2jX8dmfm321JxQwFhf//z/YrbZTyv7vZBO+xZn48tlLK2DG0DaVzo
fWHYFgXA9a3wk5ebsXZZ293FNMyacPuZ06GZYr8eJdomkahOEwzFUfbMPfb9nLv8
tpgQY8bBV9AjFhkPQ07jRILwNWEd3L3SakGijXyBiTTSZC8Vv+3sHqGXTmakEUGh
afdkDZ9r7kt2MZjbaJ36Tw3l46lHjQYU1sQn6lfMJZLAaaGSnylwhs4OQ5TjDSIS
p969VlyV/vm4ypnXawt25MTOSUoyH8WbAdrFi3+F0AxVdQK/c54wD5PJAPQeSvNW
tI5ZnIvwg+1BDcAyVdPwUiVUrnuF2gECHL7Ly+I3BIiuLdJfMespDnOkfYUxjwwP
mkeinUmyhx+FxpyDKPCJZ0iCNLNUQ7+rakfx7tHGrZnxYDLOJ+IG/n4VcIwCNcwA
HmmfMcGNBX4lRiNqPidFpn/D2GXu7qk3OTq8aIII0jbE5w2oZ9jqWVz0wJvUh+LT
SX4apONidpQOQ3qW/iUFghLTmKy/wEKO256tbgP0ZiZLef0hNP4JkuxNBXAqHym6
bd/Se7HHOQMhFMhxX4jA/CrcdqgnKKYvfm4Y2VORC/sSTm05GO2V1UFW0IZPPwkc
h4F4ajXAIpIhVY9iOq5xlAF0ckMpa2z071MknLersMDFMsLe1gefPjdUw/NpBAdV
f5xklj+Bg7s+KDUwLOSi3pkjAdzeXiEil7kU9EAdtn0P5XvW9v8ZLYnurD755DPj
NG9/Bp0zDd5RHiIOoYBC/M7f8wFCI+U2HPDPSVg7DALJyviapJ+7nZ4QXDBXSngL
p4uUrkKERWzTDP9up1h5/WOcFGQvIewCUAoOCRwz3LQNZcl95YE19lhgH+g3mHC7
ga8JLGYuJdXhjeQrlwcyENW6BfkQgtmG5/Op2XYEOCPnJpwwHznEWyax6CjtlVF8
W607iGf+gtlbbAhXNKh0FXQSGrqzCC6CW7axtpLrJW9ootUH2S3BEEGvoGj/gIj1
6ltEyXFyjoASo56SFVtzyRqhpopmbXiyAfvkbFmd4Yi3SEIZw0QBoqM3P/ikb2ik
+iO9R18zTseVoLIJ+G7DhMvMNxakrwDkoE9K8fELxTr61JfMDK8+EHaAzfZ69Nqg
UH2WvYSxySRYoG3d3l2PB195twkXWBUm8EhTz7FeSi28NyJ28YDsQhL5jtO+TYWj
0JsIC7Eu9XGrM/GiGHLJhaYnDBhZrSTdxgOM9TmO7YWhjXwekkOk/2pPI1CUoZ/S
BCUBl3QoO8/5WlSkOLRjxXtEMbnVhKQ4fN+Tr30bpkSl9BkWxWAE2IakAy2jNyku
iD5F5uRZNQS90HtH+docpRTFEw6L8mJSRaFvBzPoNGbhjEYE2N1zHtEWQQdUqm4D
VGO4WCQhBgUDR0yqaQb+zqa/Qi4aeF/mt1rsFXCX694QFN3XV0J+H30YuTPX+wjY
GNUL6ugCFBTB0cnAV5ksooI4LRmz/ngBX6Kwn/elBIt2z5JwMtkgwvjcAXzh9teT
EDBCqcd0oBi/fUQoErlYYD9yIe7dTBLKqMSQGJw8XmJECdG0SVkb+LCKsjNsxYDu
uqLdwUeoSPIZxRtfFOvyoum2sG1QqSwmheK2kcXtTfmOjVHMD31NT4CdkCSoV/JZ
OmDwxnRo9gSf4vPrlSUNTJRWyNhOpP3uHvs7EpzeobbzFe/N6jOtAxnrZGtmvE57
8H+rjXUdixwJNXFTSDiKoNBa99tvP39WnTmShg4dAJHu9U/8LNuL9gvbv8BfL656
LTw1tFpyrgF3gvQT5SB39BlyisUFANaUbcw2yLQk+XD2ebHjGEhU0CSVXUq7T3Bg
cEeS/upTd/KSrouqyK/+zr4nct1sC5ILY33cob0PEoXVrptMpGAgu2ES5cClfJ8P
nEo/4Uy/9B3GPR328NYe5lqJUE8LVbx9uv36T+l9bomi8anNG1fGOU6HTCEPOZSV
gjlsQR48VhpEarsP5aRV2VeJ+NCIl51sAlEhxJxF/CIEYRh5YfPgBOaNuoHZPOm0
iqXcOA7qp/rdC30708FJNFozdYL3xaYsVzTFemo6FiEdya66hE7SHRl50GiiIElJ
eWbBEajtBi9URE+eOH8BwB8OcUsljdFiQN1oCs6y47odeILNKUCrhWfWe4sq7lMP
V/j64lYRk/BK6/Lz31t3Ru5o5OMOfTWRX5Wn2exS3ZYjIfagEiK3dfIKc1icWsEh
h4yKyGiCkMX8ycEPVqaGinxgcHUJCZY9zUxzdxaqB1X+IZnBH9pUaMAApc8wVduZ
aju3N8CoumMjoPWmI6c7Sj6y8gJxgjCHEr3ULPCyHvM2jgfqa5jMpe2/9nYXG4Ug
GId+C8FLgFOSAy+pO4zARTQQhGVqEY+x7ab+enYLxuv6G/rh3eGo3OvE3P+Nvz5Y
a4t6a0eldjQTJInzfLKLdUlRLTj5DqlwQX+6a8QSJjiu9K3NI9EVP5sqx01dliFg
BzEZTa3idNEjv4UwX/w2y9XkpC+4xWEwreOFa40BLeinXdx4MvOskbsxvy8BeCuC
u6b2ZpO15TEsRgAiBX83I3hx0EqvAFj4r6elX86h3ELiysZDvsRqFDM1B+ZQH9GG
olb1xwJ0u5beZxJ8uMghdTDZEK/BDguyurAlDXMhcbIOVrDsKmv/U8W7DA4+xKVb
f+3s0ELGXdKld0V+MIwF0j8QekvY5sNfYVMiFjC46+h69CzMICR4iXP3aaf/huj5
+lVagvelKETe21+Ap5/ynwBQxcxmqZEfL7FSU1xFDsu95LrmwlBhglEkGk+G+V9o
fctriMs4CSRTVjAppBlWSq6dEbZcie3DtF4n2fsY/wIPlFPuhgBF+E+dok8P7Bg9
Y7Cg31QxrbjbjBymeOGGNtGPszQj2c663YxXHDvsBVrXbwtMJ1V1BkGTZ8rXsvKa
VL779sseM0Ai74PaoydGLXFqJB+CtKE9LrpTcYIiEuL5GPWdx4O5N2XlAA0zQ7LS
JpBS/+yXGIk4/cMXHpCsNLZB4UmxQApjyETPFLYUJ2zcg/9jc5sD09Dt7fZPOrfY
ltvQc0DLnBgrB6AsuJzeraockyCbly0I3ceWBQG9kAeJzFpNMwoZbHWTMdRH/UhO
xktmrJwJjkJmE/Md/HJpAM0TlH1hFrcxhCl0Ed7CHp0nk4YuEk1BzcoS+qrY0nuH
uwvs7TfLrBJ/x31yMmrD99zn1FRZS6Bya/+gneCy2aDaf9D5ZiExYL5bRftYc1Ii
35mhvfq89QWEk6sloD0LU7pvkbLBrnxlSXdsp6nKw7TOZ0fRH8reQCmZ21b5Pi/K
UzSIZgGYT29dtNaBvfmyZtZ7DFxngPZQ+eamtB8zZoz/Nb5TndBxCGEbxGg+abPY
VW0O9WqM8R93acOjXbrHCyDUPRX0RcrP2DNNMjxp4GcZ7hb3jPKHaEERgr3FoMUH
OQ0mIVB8PXOsG279h6uaEiLSuNA4w9rC74FNNyiYIJYcBFZrWTdCg0FZkhiQAcf9
QGTIvXrRLVRZqK2C3r2c/WRcCjgcqbaWc/Wp0LxgLPY3baaKknkYSvd0hfOPJdw6
gl0Fft22kzwaJsngI66mSCXyN9gSnrinhb39vK2Q53B/X6s4DDggPWTR91kyKVoV
u3+Z7CvPW78Gj4yhj0U9Jsw6OYahYsu9aIxJ3fgoluXYjx0fmUD//UB/33EhfEEY
gS/h1W0C8XcUsy+vSv4dZqF8+bhQ7VLfme9EJUvUv2H2EtuHT1DsajfO3CAxQ+57
r0DjbbyDpblRrcnc7u0NJHIfWk1iiYA73rVQ9gIDNxvEXbbO2kk3CXiSPKWyN5PF
XImYsyCvP8ONFjXTH6mWq2v2Qwatu2MoguAV7QiAjdGWLMAFcfwkfWUsYlshOyEq
DV1uPuZohqOvZn+/4C9b9/95z/I7tyilBzxY+ZWkcoWPHDxYiSTPPHIwutLZDdYa
ND85PC6/Z1OyVlLLYJ4WUTnob10lbq4Fm/LbTDnoEvD8zcYlbb2K8Y0xoFw8DLuw
GKbtQesfYBSB6fr6aN6kgHx2AXbEVaXsRvWGAgMHvfbq9Irj62u/y+4c1T0W83/K
3dWphJUk+64rwoXTBqIvQBm++G6XfmtfScHJTzFasdjzx2dq3TYc+rWWiUv8qzHE
9RHcA0ya5V5Hl/hOyE4uN9yajzrHJL0P+HKVRyAhtkBinS301HAANE0LQ6v8unHo
+ihRezOjkIAFjyWxoHkZmPAe1la+mXR2EEfK3vhPh8qGUN2LKQLwJ2J8hYW0tSYL
QixvO2GSYOF/asaT7jycrKa+SpPXCtQ98VCjT4UBIWi3jnBXCNgQUqIKau4waj6/
DvKf7MxUvE75N94ZejBep6m7f4z4LN8W1ALJkgQ6bDRYOC+dnbDtbp4wDF95y4da
tTQQw9aSOq8nbKA2JrzLt40oBgmEzfPFGhg+qV3mYkRT5wEtU9V/GMLtk60Gu3QW
zzA2Yy/erzc5N4uY21jAsh7o9maaCH8yGkhkLTJEBqvhVjACLj3v28OkdAece708
v4B+9YGK3EmR50QIWT60xvjN5zu3rL29kKtiZceEMl4Pe8qgYi21tVwDT0w//gDj
qEmbArnHsE0TLVkSNwbeo1qbdiky9JkEraFs2f214YJhqTK+6bpYDT34d8+IwF+f
QcahyElY/gdPjcNBTMNtnIvLwkpHPwi4F6WQGotJSFiNpjlFIj5WkqVo0sg2Hszs
QNkvV7rLh0k9NXVAY+qgwAonCHd8RAwvvhFphg96DvwUddm7UTTBPb1foQzG8QnC
+MFVFt/Hma22vcOINLArqEWo4tfXl0a8ZgD1zEKPTKlQ7bU7/daMn/s/XymsieVC
rg6UHIvaAogaS3JsLlqm3sL4wn6mJCFqHMjFPLjP31KbT8HqcV69iIfQu9RSrzoE
GUizflcgdF/W5Lgv2yYFqW4wtTzQGKytAyHkXpGQVWrX3jgJ11SQoVU184PZb+y1
m84UgeV4+IkavMn9FP0thITrh+WQcfmLieP3O3aQK/XqWxYS/HINn6uOw+EdIVS8
QwVFTxSo+hSMLHb1rRR2P2vlfhbEimoBpd1IDMFqQKOwdyGrMMjjpJto5oCrd+5T
nVnFJtBXnnadQ/XUD8F1MYgGm/vSS4skdkjMPWSL6Ql7vq6wR3PFMFO/Bfp/HQIX
N0WUUChWJl4j6iMTtrfXUwogVYGUZYctAjTkAvestWn+15GOOXkfb8YBt6Voj9Dh
+QPH3XLTf9wvj4914zuVmOEtfg4rkexcFTQ2VvdjyjrS9xlJri2yjE1p95kvdoll
anq1wcBW4ihh5MZ2tpk4Tba6jDHeCGtbZax/vWYWWgnD+9z5fj0bs+/JHsXgYxnd
+TBQK6k0/iV0YcFus09Ir8Aq7YZrDTw3M7EdimZENgcSS7J/6j7G5b8OeuPiF7Rk
LNamXFcJbB9pfUXIveMb3wdqPXp/5YYwAXL39DOHZKovwcmEPA0KdlBmrSM/y1iN
PqAX6oNwMBwmnhrjuFILb8Z4Hip8nU3DUDijgEfwfWDEON86rX5kgHdnmRqJnf3k
l/6aLBzAhCuI8gPC4CbcZ8lwSd1UEgb/PON9S2UXItHFYIPGV3Nwobf6nXClpvh1
V+M/dISw5vjgdNJkbVMQF5M22bS1ixpDAXvAIr1TCuv2BfRbm7JtiM1OwExnIGY1
32VqkwmWrbpBGYHF8N6UwE4Y8COjISclty91UyDTidonNkfC9uMfI9bGHOLDu/5d
kENqYDZ9qFAg34f4F+YN4nmUo8g7lGBzwX393hPpsbJD6FPbvt2Ab6Puird18b7O
6r/+dolT6/GyNlxgKecx5qFU7z/YlZJTzTrsBWFjumRm+28FubBwvs4Bvumfxsf/
/IZ6NuA0TCwQbYXYlU6MeH0ORL6/Cd4z8k7N5lxiURXBRnLE9s4hgYxuzq/BeZMU
U12TwAEvKvrFKwuVjMFft19gPGjuNUXI2GNinrDTtmHVsqdyBsk2+jm8KXnxpgY7
+zUeRqU/F75YDnsPzc+bAe1Czzv6K/1dRz1EC8xF/DJuaOJhHidDSCLXQGK2sPqO
7HdxPnqAouSmni0ueo3fa22/euAz44NmOlft3ZeNVq3T7+ncqmQJurJWXibFFk8d
aUojkUW3un9kBcp1MRQOOZQE+p/XJ+dp2x0cOBxcVUDSGiy+jzCatdhGpfS4Ml5x
5XuPSS4FoTjg0AeduFFQlccl3qlsQX50cL0VW4/ICeLY1DiwLw3Yns8mxYX6oKMG
IifyHuUmuyj8eAWog4GsCx8WVPn7wTQFRiEBxVQOjP5DrmQxk/LErK/jyCWcBLLS
s1rK//YqyThXKA1Vt8xz2MzA6p4SjBbrdgBOG85c+SimnIjz4C99N9prDF7RsrNT
mwJl704Zf3W0l57UHGb5nn/B+GXI5RE12aieXSKFfW1aFa1Ah9JXPkOK7J8hW7h1
7YefgkA5mDHWgOw1HSwAubfDmTKWHg6YJgqp0N1EGTuYRlwc2QhZ1ISWUWR85mN5
GAFwh3hV8Ut4srbeDPXIj7hOa8aXPXup4l4fjQ8yfUkN7Jee8NDKVjWWiRdGSULr
sJ/fqb9W6JQ7TZirodEDPigI+lcYYSNjGlc2AQqDjY9xHTYzp9lecDwzeb9hZvKF
yFSf7wM0qzMsfNYskSiPhEolkwv+ujOKKAohl/i1MFiKkd5leOQj1PjNbrnTVWEH
4G1mL5MF1dbbWfAWVkkx4B67C/uV7fF5PtrKzhrRdzUcpo/Sd9UXTgEPVxDUoREp
jCyuBXutlc1zMPU7CkgtQhJHsoJnO9KYS8SQUDihMzf51kQC7m9U+92m3zLhmhhf
PJZx17Cz9BvaqnpcqRr5rM1DPpkp0WnVoYxyZVuwU8w8hB8Ysf09HUKyedq8WDJt
vpZMW1/BDkPzC6+8JpifbzkFzFaXp+J4uA5DPYUlVcEuhEj3GL+nYUnf28hZXWna
cs7683lsmjjDqGNBm+sIyqiwn9QdG1mPrP3wtVBan01eJ6pcQkmcij3Ef8TwmIUE
Ez1k8NjCKKK8uz/0Etf+W0LxIdEj6/rHNDjUzQTD0Bu0bIcTu4Gt0+cG9fgH0whC
Kx0vMRlOr8+fIxe53/ls5GUvdL42puDIZ1+snFj4dJqYPgwzHUjZMNDlYzAKhJSF
/lEZ5x6e934UG3Ywe2milm9dOGEczFhmxkxMd+KMGBRYFZLWgh/YYK+f/7nj3Wou
UfTP/I5eJ5RV/EVwKY0BdX3ZJxcrAJJIy5pr8l86rU7V9FSlT31rC+dnEMG0s3OP
2qQi9GdIAp7qwk0QHoMl8arimN3BrifgsXVNiv0fTcJm2vvqfxF+zYT5n5oxr+C9
Q1DzQNm50Ji+qQI05GijzAerzoRmCp9DVtNdnCSndpGtYDbC+QU/U65KRgwx0qu9
ODLXEqaj5HcWZmpIQq+xHEafIPR5TxTIysZICrgj6u1HM/zGlz0K75oi5R7qc8r2
8Oa1vhfDlHN5OO0b2n/nMNNH/ltusD3nlD4rSu9QgYucMQNRix8zRq/J2eWkTEDZ
vGtXW5qlv/ROrZI4EvpUky0bSvlY3SLCf857LS2BR7F14MoWhRDfPfkQOLm0ifPf
2eAJ8HgIlolilFy7dPK8UMk4gqEy+28bzdvD5noP983NtoKDXaQoxqeFeAeH5ZBQ
na+uvOTxoc+9g/5dWaj9ALitykeWCeq4FvKv9e+yIomoM6cVN9bE/lwNI8m/r0L7
Tlcei990pX+z7Xi7LTwctJSi4lSH9B4/+DEAWAnXEGGEifnT5Dcn+ihYINNwsRFS
NOrZkfpt5Sc1RLMwHO9hYqFPiGST6pkjhDFGm24YQCSPxjBVBPOa6Xa1WrxTYN3Y
AIWaY2m/Q5g51h1I3rS/7ldX6cRTRWBf9WYsiLgYdfw5L78qwKZnItK/tMfLrv5e
RJogSmCXHR9/NtIX/4sOXeSTDSV0Z02GRp2zTnBvSxoFEmQwJUG4t45WHTN3w5gB
mZnG0s9VZeVFkzUQ6Dzz+7uRhv/8dfruBcRkvqcL9eWuab7lAX7dtxDv8+LJUaG8
B5KztNo+QawuSg7fPgYZK7d8/RWQkXh87c3KP7tT6u/qqVpTXRpYUqQUvPo+MEH0
gzexfGLt4SsQtZ7mu/18dP2gnmSRpAjvBl/PDhQPEIi9lPkoXxjBq3ktaRGfBskz
9h+jGLZlfF6DacV0reLA83kFjhpRh/yZk/8xma0T1mRhr/0uvHUVbilZC7EICUwc
0NRATCplxqD76Z1ZcS4GJ/3N2GgV+uaEimnqENXK1pVsOyirsQZ379l1E9x0Y9mh
Hr1OAsVrEKc9O40OPHIgRyT/q9tg9xdIhLManXTILbN2mSS7nVEbYvJ+9QVuSgp0
I6/AfAxbs5VY7gjLoQPZm5iUjomLWByvVretnILd5aAD0cDtrS7F7WMnBX6a0O6Z
4nztuKxzutXg8MLFmZY8fFcd4JNSd77Tk8WMplByBcVMsYeqeci11woOdtUMmZNs
ct7aJSBsL7ja20Ncmz7K2wTJ1cMMDw9HMR9wAblZF1lKGQ36Losbc6aKAeZdfXr6
rQpbvin21BNAnZThs3U//HZndwWIylCSQLQRwkgAdRcAMRjJQiLRSw13RJm8s7XW
FBUxzZNezKSg/CUL3Q9CxsZHJa0zF8WJgyVNbPZ97i9TAlGIfD5x6tkG/cI+90Cu
ijdPR3lMKBAlgimaRn8Tv5nkqIjLxQQwoyhTHvlMj/3isEUnUbPgx+1JAGDZOuqM
zRf4bPGn5gzbYT4N+vIF0e5jAtRSRk0I40/uQa0NDylNRlygJnyKuy85SnKy2JPw
XaJYfYCnfUjjyFf41vaGmslaxPs08lTrQL2EFsuo7KCi0QX3O/BIEZlyDC81/bys
JEoXJiOjasmoezgpq6cAFvvD6aR0br9tv2ecu+euHkD9ONecSdumlQ5yBi1GkulB
9ejGIBZOUmPMzG1DdAsw5rldau+HvDd0zfY6nf6qPVg2JzQTghtKNxcIvNKk1+/V
kVz0WvnQCaEwG9xFYvj3kIJEj+heQEUH3GbugAZewRiQTLGXOp0z3aMDKfyXdqdQ
Nvsgo66XuDlZEyjHqNQUiV5wlzop4KyrkGoYO2n51/pNbhh+nCNcJSHgDDSCyx5a
ysSEjVgQQys67DCZfQItg6d48hqRNIXQMQxXB3roNlgUPO/BJO77D2w3YeTwABdv
GuohKf+dbYEL3cfSZooKSBD01xXI4mBBidr5VKBpCabguQ6C/1kKc7F6nGzV3mnQ
cc9CGZNTMk+thD2UvzjJpa2+YtHojClZlH07zN6ple9FDavOVz4/lh2SpmZwYx7C
y5hc+0mOHU5xzCsiaDDgoAmSlHG/pfeQn/eR+GjZCc1guQYYKnxI4wE6dsDxh+OS
aY5Ox12LbdwwwaZsyFggBeOoacvj8lkHQ8JWHDVxlEVy4Fi+okE2EXZFNl+USmRv
gOvvfCpSYAdSy91Q3aVbmcTd1OyCsIwImAAS+KephJci81Nn74khtwOYFf34Grnb
smDmeyShyXFHBln9/DISrOt0PjtFK4DfUI3EqeBKNYEnKsbnILlPCI7so+SAJihQ
L2IalW6e0ZPLxDdvG99wzP6HieKC18EwdSaopKqd86uTeRHexdkINtjEsCkZBdrU
QziNGNXUuf8mI4yCAdUN2mU6oXgA+V+Ifw1pZD94FqBFHSwHqun41Y2yyBxjOVAf
gxyEz1dV2aSbKAF2re55GzPtpDa7aaJ9s8lLzvF3cNK1hP5941WFkmhsrga0mHss
Rf8fEcdjEDLeVJdZTTN1uL157ioZunzQn3/P8iaVXYq5GZz8cv3NAMf773TpTNxb
oDa7ZaGbDqlqBXxpwnkJ3lr37PBHxvpsnvEwbMK0epjg44HFy3hBo3klgfvSOElK
vEzn8AAbC7h147PpCSfA6bdWkyybtEHbsW3oucZ9g6bTvRH6HTLD2MmT0kJAuMJW
8CEyupCJlgJxRdkw/ANAEK4voQRit2+C4Uq0NaPpIyBLF0TwRVFrMHi21ktd4+A/
YHsI4FzDC2GW2Q8bByCd64KgyHgQKRWhnhcP9HMCHWgbX6daBqO2afg8WL3OCS5S
onxSrSrI2nVCieuGkPkLPXmxCHc9kBInoa0tmalUvd2sT+/DE6nJ9Wg380vtTA2M
X3O0Mg3jaqSX/UCbxDALwdflOo/IFrkKrSDZ3y6rAqbLut6yiVlsjxjd8ymL+v/z
Shf8yrHZung7dA9c3WHQIaMIdpgPwKaoH9sHr8C+k7dw5UtoaxxPUduJ54VkANwk
q0kGeBI2ZDU2MLguq+IfL8B7fiyk2tXhRc7aNcfzZxYW4nSR7gjoFosTrj1NDPmx
YrOqwGcBsnC17SIAla+Fa17MI4TxEP1mZBkB9u4YJtuEMsA1XOd0lpXLZ71qeUu9
pwY5FpocsphGBBJTRog2BtW5PG+1oxhEZVvaxeE1d/zQbP/OdYqBxjHn9iuDoC4+
xINJI5dyCAxxEcUHOqK3F+dBUqKRbdN++6w8PnzH6nkEY0aSxTlf5IwsS6jE3M2k
Bv4+VL9V0IarlS4HCPxRtWh47EGCtTkit9abhZQYnk1EqCHNQAqHF9fYejn+EIeD
rzczy4zvRxL4Zm6IklI69+KcMbB1Ynu9rtuufh+B3QxosYMTK2fYylFbmKkRFQEA
5PM+EafKapkipqZOk3F24YThGFx+1FhFXL8X+BmNQ5Tb/+uInpb6Omgz1F1odUqE
kDnTBO7EN+OcU0kwD0qduKFyDm1ylYFCuHGyniv308U5b0/kUDboD5z2JOqYuZsp
J06LBE8UeP10/JlS12lqqo/ZLqSTMS2PEkB38up0FKLGUKLCKY9ga68XkzhV4gRq
8EocHyVhVFTyrU1vOtSZqa8mPK+KzPV5qhVVfAX75sfqm0+daucsxuRbQptZO+3I
oPPmP5dHNXvzNyB0t+vLyj9LyE2Rzpr+UX+WAzTV8iipn1zDU2isZkbQfNPJzdZr
NC+XHP1v4mLo3ze9Mrz+9F5Gxq9gesj/XBIZgOXeW4QyL0RQVeMIZvoXZ6mNbWLJ
Q2GvOlBtsdDa0uwHeZQ6/nb8fAvhmaKl1H2/O26LUfEWyOZmEvY71pHcEMBffxNM
pPewNDPPwIpc7PnR1evRppEVvydfRjpJBNTFGLyXejpMPCWHYBGzqkJNO4zCcebs
CLJP+np/8ldbxtOUm7gSxexi6Xc5k4NF+DcnSn6MchUEF7rrDjMmJxsrxND5/Fxh
QnX7vr8njaIb+QmMGlsqcAG+eGE9XV/NEvjkeYUDZRbmMDQUzqqoGvtqUIPnyXDX
tBbzeh0tWSLoRuvjMghQzciLKNy+kskA+pN6qHkhtaJP7sLp55qiqOy/bKXG/ziK
HqnvjQQSNNmoZzw2KHZgD7myFaWA9VhBMQCKpeARJVx6adIWlUCGMlRtWTmOOTh9
Kuhq7oT4IUAZ/kfzku+KMK43yN6cHLzlmKcO3rqjpO84VFJ4+5aE0gsTk64OErHM
Sk+uFIRjPvZgzuGm53mYLeUNQ0+cSBtyKjdOY+smatV8OMF7gNdFzDc/Ump1Z1g5
ngBORtVdPKzIobPUv/aWOQjsER4EerCpVslVnZ+sTaBxTFmNgQlaIlld/U6ym7Pq
2bhMxBXTlrdmrMkHVIUW5G8LivszfExNJaiY4lnl9C+wSGPN8YcN7gsNyHofs8+H
bwV0yajhPW5jQ7d9BjSADea8I837eCL9r8DJboHg+VXJv6+4AQxiwgLYSw4MYIRg
l3Ei+evcKDcehi7wVGUwl99ZZEjzAm2ULQA/k+GcvitaesXDHoJl3Lxq/zjtwMzc
U7mHIWBstRBX/+ZN0D3Gl/PR3N3HBEC7vsFATQou9KBuFBbh+3ZsylRJ0JJythiC
UKk/WCYF3GFbC+zsB7UmXiqXeKskfV81gFcM0/mW3mc2ZKMZaDoDaTtpDCN+0iue
2MJ2xppagpwXP8Es7iTg96o9TrgXv3GcvxU3CbXPpjAGZ0wImyDN8QG0N47TMv8D
o0F1Pekxef7emM4LBrXbU99TfPhEiP4Tn2kMt3lBb7SkMjU13KhQCDSbbJFXs8zS
fI9PJG6la4HjW6FQRLhuGdcfBCp140ZiCjBi+aBKfqj1v2ot4t6zoQBo0NnzvvIp
lJcA221y9dDS3DJGJSXeEztoTN77hVDRbykptVg1wb991VQuJ35LIJpYCmNaqgD/
NPXybJn+C7q+H3Jerxc3c+MuQ0qspF1f4RQrSA7xCkEZk5A06zH+WaG2ZUFcHYko
orP+pHt3pibFgHYianlyr13CPPA7BcqfmwRQOR1RwBNBgptbUj6MGRbPW5+Oe0FJ
iGTRThUP9csM5xzbPFbTfhRxuGshs9n1FeDyK3u4AnBA1pMgZqh1hqsqKJMlJeuZ
Wh1My93kyu/w7ukqwurbmm4F4Dm4hSgnvl/zCxddBDN6uePV4GQNB1lnC7w55CqP
XZi2rotLepyakmlA6+wcwA7ZZQSa/G1MMX3KYV/yvRaWbTEW9ru22GHkvnKGH2lc
2nzLb1u+Ydv8Hw74/tP83ApMNSHbEiDz4960f1BxkEPHlZTxO+dwDjRUA4Yz65kX
uAhdFI9AFcd7pgNH7X1RESxlvx+NtdDY8ojmA3Dc2GiD4bBEgON5nAqLVd7ZoxP+
pC4hZI8I9RM3tVv87XF9pVpVw19R17+8cbltbNAJePZ/RwFtY6ZxBgFIKwqwemez
JQxMbq0s+mD6++3LWQwYXul6Y2Kq5bW07yjKH3Q9b+zD0aO0d9LmD/1Mg8V6OX1l
/ZdEqAQMBouK6I1MEDxZ+yb/TNhqUGcinZP1apUQfCRRrF63SxbgjDAU8j8u33p4
hLoeGPA3l6EwDRuZ7GuOcr4Myz8yH4BGtKqQo8BY4AdaGJ2YEHJIPWXbsY6kwoAT
NReM74FguIbGqzGcHQNAzxbqXwEWcsxjDoFaS1zCalnjxCtYqr6GdIQBGdLbodVs
CcU0Z5B0PME8aYFOuSA1mPi79hce+yYPDhfms3yetqtOGL18rOGnxY+Gr9s/154A
k2VbSFgfmSdnFaILJ2dTHjRDr5oDiKWRZkwWoZIQ8XQZUvP63SGdI4SJNelLkamR
5XTHCKqt40UjzVxiKZCeyLyrJbMpRGCQkAYqouDhN8Xf4qFlrK7rbalJBr/jMsD9
sOqF++s6+2yfefUDsuK1JdQPV/l2skuB8vv8O/KAmfr50SV3DJAAExunPJ6zJnZG
8NryYdk05aQ2l7ylP9pYk6HQ6jIpdoK5kEISpnQkBt1+FVzpAYDqVjlVrLxVsLBb
j+Jiu+yPawim6siB1yqEuhmI/3vNocNMXdi1uatO5eyAl9LuhEEJHW/DeW/VqFzr
1FswxA1LMpY9s+pdL7vBvKlZjfDUlytaRaV1IY9fNEFIHBS37XogWYfQAXkX+6Kx
JhsF2YFN3RC0i6gEmzVTof4kZEODeM464uDtSAECV6nDxBcglB/ACTI+I2MuINBp
eJ4IOQVTzvS6C1VoAttdsDqCFJKG/IkpCUlbw1afLyHWRSWc4LhVEHd8myuQaSRD
nbvfgF04rgcAm9sgwE6isXkSygcaZzCizQYl3mUHxHhz+hmCtECAygkpHeHbOZXP
EsJioPqz+M/4zFPQUeH1Z3oB2CN/bQMxjIoFRlq6dxSdtB9vtpM1OfXc19ni/QnV
a42kE2rAGp7DgseaHd0OK52k8NwWDShVqQ2st0HKPOuWs635CJ8VAA4ZL1GJbKz/
6mhi9AyEurI16D+aSOPbAYdHR8RiT0DPYAc4hsqK9QU8fipXOe5OTBXB2dcmyX46
FxCuUP5Noah94ZYLFjXDUe1awiQyH8PwU4se9LpQAHQwYRAODB494Y+1SfE0tcF1
7jM/udUqc4/tHH2h805PpvIsopV6zTkZDSPxCvJuwZJuEq23swB/vQiDJcq4g1py
vdTl8CJBoC1ncPUYY4o1mMywbNE4jAMIfwEFRDJ0xnwA2pqgjEruMrCdXYfUPrH7
+QpayRuO1TuWZqmgGBBMah1CulhM2wYXsiZJNPf1tuDl25npF6RJgSVAeoDFNEqr
KxcKq8IhpoH5+HKCvEurbVb3cdyRqBxfzJ0qmW9YX+MecrAWwiXcNCp/tMcg4yox
9IYJFgtkAT5fZyjoNqAA4T4UCpWR+LMQ7l/X3XouwRtp5oz00lVbz1RumuARsrRK
hDLRtamkJ8ZQdwweOqX0hKTPDH95t0MwA0yd6aDRLv8yXnx+mD7Di8JDn1VERYXk
9S6b1Qc+VvOxIJJ1/Lg2qGVCK7xZp8xRGMdq22hwUVdzpAOtis+fVPhQGfn3NEWS
SzY/v7zfsmW40z6Ko9vEV3ySkbBNo5k1rAMtnPb1iTlVdLCa3N1xF0TQE1ufphKh
2oAcWcVv5osaRwu8NMcp8kRS47EvB7BojRLAkk/2M3zJwpTZ57INgdAEw5RPvP2j
HFhtb37Ro03djQkZoIv+eobWeY/M9/RsAFWk2th8bHUCcjrgXqKBwi28QlQlQBJu
9dsKSpK2/9FVaNodWJPkGR43l+ZwYyO9Fv0HJletrBnQ+Pz8Jhpex8Y0C1P1LWfs
+jmZ59wKI3gKIgsGo5MIdauri5ZdRHgx6Oz7fFQ2dGMSXwN/r/1FmV2hRNqyr0Gm
MwFicYg99pcsU4/TRj2/zLTaGsJGQNyTNwV+fHWxIgIWH4vXKg1O8yoQGr3vuxFK
s4FFZTw1IczAEByX4iu7u3+RvFfRHvZ7Y6VddXrOS8Bl66j5jcsxZ1EATrm4JQPO
ltwr01bzMLvr2Qsc8vQfEEe8sgJCdwi3lmFGezrXpX6kBaVJ2pqnne83KFPyiYWW
ooNF9TwRws4hJ8lIE/fNm+mIKRcATGEuTEyQXH2WNvBLNiqMyrmQCPFPWLcxw/Om
0L5TOTYUTE5t37P1BeCMHCVx6naOhT6yPhofXxQDZG5rm7UkpnF75ZGeCtAeg6JX
Iay6mVRr+LFq4FpkYVe/r4nSOq8FEIKLvzK2g6oX0cackpBOFuVSJyizFZQ8V0Lg
XjtT+qAIpblVZXE3qyrqhLqnDz7dEAgMvXrcjjkK9psTlGHBJFQXXeBnMhwW7QV6
tpyXVvZsMAQRPUjgyQFPANTcnrvuy5WWgk5mjQ/piZg42MMdCF/gucaeFzkLqw0G
WBY90EoLleFubVUPZldM1S9sycubwDF1F6EUp+zz/Xsmdj2n+lnomceftuJVlKbx
qUfbIeOjgiX1xYfldAAyKwzjyoBRxVYwVsj59RwaXyHvXWtP8HYHt252CB1e/qGm
+2ecSJb1AzcMhW3Ez3ppEaWYd3KK5gwz1zRchzJfaK/USUSvKcjr5AHoiy0ESyLs
/e8g57E16FTjc10Gz1eQ3tH3r0sYKznasX94E6YuZQzgnxNcELlUEeawN9L1FdgR
963Eq3Oa2coJh4Bjf5L0zRwk/C+PdiAjypCPF3yTQTxj1rd6hcKrzecseeBAeyBI
wruwvEy7RAzsK+L1BzLIWEl7dmQuzEornYn6pa4cF2i9FhOwpNJXr6IiloXWNVIm
oBasLVhJ7Zwf40fvZ6nJkIxb3PlU6H9jpj0wCiNANF1a3SyOKR4W9OPk97AVVSJP
J0LgQ73zflpO3rJwH74MWRI4KZgObE8HnBIgauBqsPd7KEH6Y+sg+KASd3Ha9cPu
2MTphDz9g0nOptrROF1TG3iWaHz8gpNcWlpsaRqhT7NRJ1DWdsr3oxsVQKZuj0+T
uEB8o4yBNzSqjuN9FZMWvZtTgb1T3Uvf8lsNsF/J7u438G69Iu1X3c9Ov9FLVTkP
nBVFduHPl129i6M7Nv4svIGF3y0u05PELvwZBZHpHPffnxnCUL9kpzYdEEt+7Zbi
do0EqIH2PuKkDm/FnWLx+m9brQGWwLyZE4HUeY7V1YScmFW9UxDReKuJOYGhOQj9
m43JhIy2BPKPfeStZI3Oupkan4yVMXI5O0aV7R0110bRHWnDSNqmhtm0ueIXN0dm
wdUSU7djNOiUhUBds6M6VberOzdDwSsBbrfBvUQNZFTRRWH8+XfbIoAJYUP7LBNN
GWv1sLSbCzQAjzdRTRySpnbB25FHQ9cGo25xukFwHDxzCOnXwZYhIJSBOLwl/uD1
EpDotvgEfAYTco/ef/JuKVPny7KMRdZLeFCYBOVmxYIdLdhDRdImtzOX2m2GeWmx
LG3+2z+i8clmneixHvkQ94c4dnI6gYAKtuSzUXP1XpzsmwMnIb+fRT7sJOr1aA1I
BXanx0P2TJY/KsGlgnqXZG5WrZXU2Z/tae6vSS7ddsMryBqwBZmoErjVi/6CZeCJ
Aa35ELg4RKLQSqIqiL/rUYbvq9rxFny4oBBN/7IJoZpTM6B45lqJXF/90ZnmZ4bH
9s4w5eqtE9l4HmUShzX1orFKz4cRklsyXk2WOE8+W9CuQpshI2cNXy/NylRQ4j5E
VyPb1STYoHAEdOD6np8g7fPOL7NhJJ6B95uykBtF2U1Yh4uAWMlaXF8jiD4PBenc
u1sMA1OZT/wOZB1JFqhgRpb9pi43K3sqKlgsxR8WwOFg08Z/o4KQnbsQd6ivNLDg
ybtEY2MI4eTP+n8SUyPbHynvxn7DTliXnrQMTysM2pkwIr2+xFtrLgnib7JmrM1a
x4cv5ev/r/SaVQjKcehpRPt5cdjhN6V5F6vgb3PHBx+QxLfux4n0A5YXs/lVUsv7
jL4TS9xDaPDyVZEupFWorvKWicIY5NiIYC6slAk1a9PwPp1XsbE/F7odK0jdedhv
opRpLCke5r4sV/V3Srs7DPy0jOWc0t5R9SeXfscfdur0jzHErPs3YJh+YpGRuBcA
Wv5/lNfGa9WbavEs4738bjx9+v8C+wG66jrNZy7hOj6T4Gsx4+yfkCUG8j+Va75w
cYNCOGuBqvYuIvHfvYZtVsa0rKRc4lcqq+wGvhEozF5YuLO6MWgrI1BqJPbb2Sb2
TT2nnG4sDozAABlzGzL6NQpJqwFPG7WXPINFmJUup0aRMLqLmxL053bX8JsbWNnc
bRebYrMSYBn7Uby4CJ6r0yG7XGcXj08ntTvjExtkPZzyp1Z4521kXzlCo/rOhH/M
JLkZ9vc480gRHkZOb//IKiCDMzvgZJboGeNA32ndPd/LHIR7kAHzn0lfu562YCwx
s8Z3Yyo9J/op+sFaDEplGbgIclGnwhHpFqyFKktfiNKyMa2RDJRR3vknIVWyJrog
4foWkRCPEUSg5H42rUXqzwUkzKttlSmhl0vQqRfHlQOrM/ymOo4CToH1jnbMtPxw
QqfSscenHa0v3lJ3GQ4I8kzz4aLxdzrvwMwAFGSILLCUnwpiA1iPmLts4wxcTYo6
aBgoHFoBvxyAok4rGPBrA3Gn8tHaxRNkD9X3wK7IlLYsJ+anNrdoimbLoK4JbtrI
O6SNRRYllTqTufMPwnkWX1tQhj8aAqvxHP0KfchjK8fypsCaEmuSImZBcUBOt8F3
mnWiXk79Zc2sxT/Dx603Nt0QrgEBKyQjOjw9IUnaC9R71xGHg+KW8BZV5BwN+O67
ShxP57+kmptna3ly7V/1RX2dnZ3FxsIzp83fUhPbdyCqlnOfQU6zVtFd7jcCcNtx
ixfFPpZdLczLC4DLRrUN3p/s2KHuxKoAKL5Wu8t8Lok62/WNJRcfteX+i4xM6lag
kZfyzTeS8i4QW2RsyDZV61NTbwUoHbwM4RRtxL+u3GJLO+9mEvaYcQMB5CAezDG8
J7PY1kK3MTV2wXShuZZYwO6z9Qm1PHZ2vyS69UF70Q7w1X+Uh25+85uplCxQK42S
PEPNgTPR+xqhaY9/L8crjLZDCOTYY0dp8n6y5hqAqrKdfcVW/rn161fdj1c5EPw8
+F4wghMQmneP7wMG6/BP+nilaSq4vw5ys2ipcsSQSsPtQ4p1c87E2mYVJGky1d2D
U6EI+C8yWEkBApRWz/J3rhRp3jCDDpFORzXd3HoqUuUfctqO0iKmdDFmQ8B2i2bF
uphovYMih/IjsLWghzqjo4AuGRvUmqAcN0KdqhL46h1dfmIrq1M/h1WZenuHq8cr
MlTM+blYfmyPwkicPu6i98RceAvbeQFPxlzuMyXvNul1mKqwNDuVMP7xqvGwWmJ8
Svj15d22LAoW3XrHJIPhz/c14CotpScCI1MFDg55BaXojCtIKF3p5nw8XWNEAnpa
1/Z8944SPrFdrkt42Tgf2OQXWmm+pD18lFYj7NVcVF8Nw2ei2Kil/LAG+ScBXbtq
eptPwgMigacGyHN5uHx335tak4farZC8QA9Mz5K0zlxbilzUtzUGNzcVuAWI8mrb
iTwAc5x8UmZ1m+Z3eE9/uMN4bS2dBjdOJ10B5rOq11NtGWISpQ7ruhQBzmIqofuK
F5ol/M68bD/JcHufDbCFfWIrBOBQOQ7doxiVJPo1fZ//HVnt9zsrTHtJp6vJ/zib
+kSrkQ+tUQNLE8u5+K+N7H1mK2r7+lHuC3hFxXpts37OylAk/Gg+ccCR4oLUQEH9
vlDS+cPMXZR15xnnPVUu62qoF2Pxt11+WV3h7s0cLsLsJPgnLCKKobPldeA1KR42
cphnRQrTMA4JfpEX7IcCrGLIRabDaHyfCR5gXX7zT6tRMT9fvaj9+U1zd5uhKnMd
t9pRbwy7P+2Q57YOjXu8FFBe28fIF5yrQKay1tTO5jNvN2AY/zMICOuKITu0yVp0
UtTdjDkHuTfmXEfJP86sOrF+dJX6QeyGNkBVvlSzvqR4d75R1r8WBkNHGwl17L5l
pC0xkW3mhkV1YR6Qrt9/xQehwna3uxm221fALhLwOUv8iS3/WZ4mcszrsAd0SuJm
BE0wM6wsbDLM74TCTSxaWT6z9wzew4OJ7mGOyoJnVdeZF1i4x/H+Y1TALmgHpH7w
GSG+/TlE5VOf+PZJ7PxLBSenYxg/gBM0hRHgdlMX8R1frbER2RM1a4Iaqe/Tx8ls
el0sIuyYaswGwqBSgaPwwi6WZQhOGwBQCTkGaf6jFiPZ77nZuE7Nbb+Z+lujeWKb
mMeIFHajm1SqIrqCnntU8BqrIHz41Bext47PwUu6iS5LKAt+JOayQC6tw7TuC6Ev
ZDb9p80DHuqy8VlwbL4Njkc/hJhLEQCK19ihQgG6R9H4NO7w3RZyvf9oJIAVRbYV
xTmYgwgvbC685aOu/NlVDDCUVqukdsYsrYH2gebqLHHygFhH3QE1FF8FX+Kld0/g
dhwja4QbmgX+yAHG6v+cEjObI6FDu0cAoVNYgDGAhAFwSKtPwjHm7HXkqiAuLsGf
fh3aj/m6yGSIFkd5q6RkBDnD+cX4Q1NKEHfnED91Bh+casnTX0wd+dcFQYuP3gNC
cKfRM1ivIXIUx9Zd1yRsMbxItr+o+ViYGRFre9EA2RQz02PESRnEdEEGDRVf7kms
FOf9U/lpfJDarTKchfPqYQzfK9byvPV5JGYrNo4U36WkMEKI/OjLMaLfVQ2FQiKp
mNrKD3jDIEt6M5JzeZeCYWsgWoRm3UZORLLa3flwJ2feVkky9x99bovkXYWHtYJz
dr6+Hf1WpOTDz6jas/lMkCXe3R/BlUOcHf7O3L91BkDU71+46bysqQbbjwkPiX5m
pKt7LMcc8QKLNFZDwH67UNu4i2QxH6mVux3otIulhig9xUziiGno1aP9CKIOhfRl
ey6DdoSjjIl9P1KHqFnR2zGmufcM2ISIl56OoBmdL+nLvsbW4pS2gNMJzEG9oSUS
2aboze54mvaLQSsIv4QOttR/kUImluNNDkjSB4Vfj1YFT9R/pWwzICGAln/il9Tl
ykZiUfhxGTlOXWR2Z6pqCMY1fBjH40WHEoW50CdeVkkyUkzcSGUboxDIo5T0DGup
XfmZdW6eZdKD0I7uZ+8LLN8uA8ECAfeBGUkqjQ5R2EB8Yx5a4hIEiRva/wTyPu1O
k0QyjfAzim8YO6DIsjP/dsRgMXBQ2JmOoNa6HXzBBoXOrgZLkkSBNUw8qboN9RVE
04Hb80y781BVsa/UfBb7Ye9suQdR0zkLEFFmWKQvYv1tywT9hF8EgNOympB0z7j8
QePjdfrvKx7Mw71uoab08EZXqYZT8YayQv/YQ4qpm+SiH3dpNf5KQUBW20LnT1fY
W8puBqRJCxTIj0FOhs+hVCoi5GxbP80eBD79Uli9C9iwp6x/rhhz95LPuTijtLKH
w1xqUyrPUc2wVZUU8wqN6stlsnwMES9Yx9amSdPSMDNcFPDL7vk395F/OZC/1oPj
qyRx9vNDWoGtfGQ594FrY5pj2ytTtRDvKTzkgd7S6/jGq7h8W+iR5noY2LX7Fjqm
Erqt7zShZ366rPBPDTuOQcd9zQhWP1WeGkNCiOkc6gUbUcL3ojCYSL1lTz4SjBpt
1zp4mtgGF3kEId8gXeKtMRYczuZJibzrm3Shag2+sgBxxygckQ6grpBnM4+fTOF+
wVkAcmXyGhHZQXCImluK/vXNhDZr9UxoxJc7qpZCs/7dQyao+AJDDmSkaLcu9Q/E
vk0a3zc1nJeIwBoiXTmgAirKd65uxxik1+CAoDtqRhcZMvg+Lvy/HL/2EEgECDi4
VNZt6LOejiPr1e0OsWx7e0RfzSwldc4wcTh3D7dDzf2gnRz6AWTn71gzbv9l89XD
P4v7wp7xpPGqq+fKEIgDT2WRQk+2QEDXYrlMCMWSN4iYDMCz+MFnxKfeyG4IZDwj
9g+vctvYJHwSt3i77Ye+PVT8yVl+NYTtVxzG+IL00ZnZSxqgzAi/6yUZBoE0k56u
oOa/vcCsKr75I+ZrInqTo49pvoUeLypVXp3SlxGMh+2XjrJg5ST6Y0IKbYrz+DLa
fIfiS7NoiQHkP8JEsqQ+CJ6FNIO7kuSiB9QNBdvCIxpPTDZbJF5RhFFyQTDBLRtD
tIDRTtN+YyfprOKjEjIenQ081LtjkUqC4C51Z+q5YyFqxEJBDl/+rpJO0EZOSqyo
SQRR0UQV+G5r+RD//ReaNcQOqh4rlzdCDUNl7JWZLY0mbpJjWzB7fzEgpYMNPkDr
a4FTKmE2XumCr1M2C3GvBKTEeZSp/6sT0PDLD404OCBk9tn08QFyq0keEBQb06IA
e50GisxOTcmzTQrmavJm+0q8MqnWwkxGhNA3cV4Rdt74dJd1y6wVwSYUluU1sL3h
OeJdzT6FPxqMbnzwccFiweTXxnmjQRd5mZTxQjXY2yOKtmFirKcWuXIz9ZodsAEM
Wp9/h/RjJ3BkKD+Won3+doKs5ejRIF/EPIkATM9f2fcjEazakdChz/DCi/4deZOD
7fGlFyK3uGEZtEPOH49XZCMjYyaGvkVuaV8b+nQbXqea81aytu18wZS0MYGquh3i
x5+UP3XOjSs1wetSR//ADq2XpjWuq3WebozT6Q/VtOhrYkTaZNNfEj7Srg2tNUDy
S3OXBzV4MzV/Br0AkDuVTSnjpPZK2iQ3E3nXja150PtIYPZ0PsKeFgDyKtM5BhiQ
oneUsd0oF4raP3egw1Tt4cG/jEOR7t8HkPfKdaQMUKFFScTNuvRq3w7Ix0xNlzFk
taezlCi7vWUxMCpmzi3cOMFpWKxB3DjMGeICU1Wns10ij80UFE3/q6F1MXm24/DG
nLgw1BhXKgzIwAEh+CSU7xSeDiA2VyNlfuceGmzcUaCsndCJClAX/6KzrZqpfhxT
mnTXeywtRBX4rIm1Zd0wRacnG/0Vtk/BDhKCy5QYpDlfBY5+cW9hN3I4o4Fn7h06
FBpEEjw1L31e5WjkxMW7rUpJ59HsxBDHzI7uk/VExnT+OwB+wgaqyFXfiILcpOYv
ylO1+11XnJvfAejsa22h6BCk9fGbKqFko3H00nuuYLPoxha+PKOPgzpz6QGz32Ki
SQiYEcfABwjhMYfdHwaA/KqH7Zk0Zlsfxl2ghq68LFUjE9KFp43uBEwcW+WR5EUd
biYzdTqIdKcz7OEY/OOp9+iTrI7QGwxQPsicW+xiYV6T+BrlEkvVEz9VkBRvTeCw
v4oZLOdxHoR8FHdhePR4ng3O8aib73iN2q+JiEu4qIzVV3Xt1XB/pnEaOulbB0eu
VgI68GrNx1QRzSWhlPlFZMphAzdyU4ar6FG21D+/ZsciskA9/U/JmISPw5S74Kz6
xGl+zuExuqagDlXkV/qOrxyndzBMKkI/YEkHdGXZLZX4hkscLxJ9FCCm9JPmI2+1
zfWc6tck6+BC6bUUqv0eP9HBIIpyZV1+pgnl+1JimWF7ZDEzA/Q/c32FDMRIIB3j
+590EuKjaG/nFvDQfsRsdo1r4NW6n6E5vVmA9tu33cySKgS3VeGYgp/JnnbdbQbC
KlTzJVejd8HgqhQ/sdYri/wOdnYK99XzLIKNGY6l9SxVNVoek9LPKrWwmCIN1rqz
wzNHBSTnDdL5/hNML5bPPXeMFpB+sSxMFbGgI4TBiSaH7holAZ9URXZQgWFqmnaJ
OtQSKanMy1SwORavUaRegt9rM+omxjwvhAwZegINm1eAYCt7o8GJjQ+BxHrdrUyi
NtpcAufkBwQSLi5nvTUI9Ta5WAZPlFlxsYPxvn0/xbF5Nrr2nEwRIqSr6cmwy0qQ
P4YQFna7xZUBzXprbxFkjTM+VU1iKkmg2IcWvaAJzrWS7fPBgNdjen1Ifg3oGcre
kMFsoeHJ5iOi62ZI1mQjjgUGiTV92usizPOk7PVG9XIc+vNBecXaHZbvz09Ro4m4
TqEk854GJ5jc1U4Ucla7dNC9SZXunwb9xrlrQpNJALWAFoXB9SS0zTH+eFvH7LAz
70rL5OFJuLMhebqvH9y0AB290hNL2SF3fqiuTunO9yEuxQUM7QqzXjJWdf/08BIN
9GqTpQgH8RGX9tZYSeWZL3U/6tpWyvv7uIPFb81mVnamuusX5oUdf6+ddyKMwBa8
CWxrNf09x2T1uNUlHLq09JgJKCD4Tfsbjm+IhCrOhIKF+zuckiEk31+YDZR9wvlx
ovJ5Yb9rbU5jez9PAywXKe4oMfxmzW9v/qxKwtO/F0NPpHvyvr4AMs5r1S68gKLQ
uarAH/+VK6RKF8SJ5lF3MO/ubI0abf3u6a0VFs9HOh999iLo0LhWbMGWbcpUp3Me
q2nKyG1afvvvtXy/FyqbD89YIDrTbFx2nBZdwDE8uilNBVksXfwUex8fJjFd0XwL
H1NNdVqy1uok5jR/mjt410CGJUgoMt4Utn7vf+VBBi4TdBfegT3mm7Qutay2rtw6
3SLo5YIixvTE6Hq9Pf2pbgs+OwWM3ZQfxtS8Y4U14SekiOcyXJtzXsVUyA0toZdH
bs1Jm5hM3WVgnp9Wmiq/hWNU4/b0zjJDvWX8dQ4yqAGqZY+olui1OcU8eiYFu3r6
3sdMpKb5JQgy7cRmH0nnVcdxCQICYpdGaLpqDShb86d3GeqUZ7TVeRXGKH4bC6qo
9AjICJaw6kxCU768kY5rfV/9W89qEP6uAPbWUTDiIn2Og8PrHDtQOVMUOr80E9ux
o2VqpttXrOHQ/59LqNXh3fJtpazH3mdRlZvnR5RnYvEWhUKBrk8XWYwjnpT9ddaR
cX7R5/Um3zh3d19c8OXv9PHGrUCh7fs1A5RfJEA6euKDbxoCoLh2RSizvU1iIQ9b
xvVY+TFJufrqQqDzaITkZ94E4ugIh9M/FQoE+vXysVsyVBXZ4z5aH7VaVpedkWTU
ZldDmgunPq5sdQA3koF7OJFwfVtdzBUoY+5TmbM+mWMNuTmwfkGXL0HSJ3OceijL
oWJr8KWlLROEBC1le64WQ2UpL4ahLs3JBstCQA0Km30tR8kq/CURpBpQaf9Nqw9K
5Qmw+monewt3zfjz/05xOdHuBvTTmc113aDfd7tRBJ1kjtGGlgIH+S6c21Y8snc+
p2OyeDBbsvg9kkZMZkqIZ7S4zDoda9Pey19fY6K6+IWGoeWvIVabnkuEpvWcaVXX
h4xjyGoMnpDS2mA0kALGlip1pxY4LQQ6OAJ9Jtk9dn0Rvny4ckwirK1Q3phjE5zy
tIItOu9WxTcp1Tj3il+BOabC0XJcXCZjVbQTNdE0b6e0PiiHuZ263Y8WSbZj2g0S
WUaX0NUq1CR1IY1xRleGNwpTzXJ6gXUfT0Qshp21b1XY1fpjlClE+1TMaBjnzLkU
OUUX5ahM7GpnsQ0xvcrWlmxJUGqy9PDMbZCqvRNi/jHD0xw0Hk6B9rFxQdzsvbE7
wXblrL3HeBgLBlK7Jy/3McwHc93HUlqRSIh/fhOxnsbep8K5Cqewyi9BPLCxNsu4
g8Qsjd//LhS7F4OVNQaUaj1cd8z+2A0e5T1YXwU/NsvP7Oj7JY2/njGZVUTXCf5S
McUKO/vOxVBTxpD/kqmG9nU+oYbXA3muwULtmYSLa/r8PPBgtplWNLaaM4DngAMK
3LdIVAd+ejyerJxeCxPduooadfn/ssAjk//hj9s0KFFiycG1Kp+KDSHj757XHKX3
A8X8ERwa38W3bf9W25QYp8sJkgUtVKl+nEcdfalT5lix8t/TpgDv8Hs4kyHW0uWk
5xOZHkditM282eDoJzTifbHDeGme/231csZCFA2vT8F3GgAf6Q81ePPRelZgAL1q
nN+yp29qdtkFEYoXY+ZHrgO/lL+rgYpupyf9pcjDM8uZP6AiqnwbBPIbIFAA6WlD
eeqhCW9mw/UxtPnH8ssgosa2UgsGE36rZ8cnATLvXHjU9AcnicOeudYdt4SPuG/m
7ZjBscKNhe8Yk/oeHNx7aW8TxT8u1Z9l6CSBQ5Xpdv70ue3K40mGdMUTgh6Q5ax9
3KrcJohVLvDtSXz9iTBAbrQc5SrQhMZmh9lJyCNwOcr9vdEWOjAr65P37duxNgoh
LRvizgAd9OWIV2H+x86TtWn88Avw323kMGxKaYVcDITHiszpL2WbDPV4/cacTDL0
f0eN52TLpqTj007PokawYv5QzWuhDS6Qd0iYJIMQcRWLtheulZvIonv9X2+bIDLo
P4X5oRBu2IVdsIaHZCnoq0WYvN/Facng1ORaFK8ibfcbBohQkWjKqq50v++//G+I
4jzbMyJZjDFauEmusVwQ5NVOMw36w1Fex5QNrMAngg12TQOKQnQgSTJ9t3a2yb0/
uiPiz82bhfaeh9mPTjmT22C0cAdfp0+zfLJOrhroYVFX+ZifGMa7OTHt2LDWOaGb
K3hTTmNAOTOgHbBYWlXQ8wXlpXpJRa/FV5FNiTqPf3qaOlIkz6ldzrV64ptu3xgf
28WVsvUza7zWz3xxXbKru3VMDqQid0rFDDh2vGA8bn65sUNTpugm+8pwqvsy8UfC
uQ0a0UNhrUeZiuEdWzbx7oYtK5f79PXfIJKgVLr8qgeho7j/WeYShX0SjkjuBuhV
GwDZRsFNz4zORVdlkmuDMVKBX7YUpJR5TZjwCblDferAA9xf3ucASEgSqVnBj3qD
xadT1/FembQbDckwq/7eVD5KADzPokQy4WFnFfZS9kpku+pjsKFN/kVd5fWLORDV
7uiS0UT+AvOX2Gk6ZKBBo/qr4iKATLbSMn5zu1mwZ7LkVnPcyhKdMi2YGQUIXY9c
ltdThf8KEONUS8l9vxhrKXCgmBbOl9zS9IrNMk0ztpxOoZvP3ANKPQJ5ulZVp1ma
1+R+caj907JADBtzc+XF6mNh8x23pPUeL5jr7TcUOYgBYzhIvvLlm7vU0uhbcpxy
drY4Zz8oBpe8yVux3/Vu3ATasZ3VJruqN21z3cfRgCnJV3/31bWwGYX8f2El/duM
mJfc/uQpi9zE2RmLNE5hStcT96IBRy/3N8RGhjT6dX6+8OPL4IIw8qPiE4iSqHlX
iftADQ75Cecsa4XRAvec3FLwDnucTHxmZhiLyZULlKlWgRoNIvAQ1NXBfZb0Gy1v
nGZJ8wMN6VS8/NhKJD5VQSwBo/OJnOpViDyhpI6u9baqH6wpXJdZybGT+2YQ9vob
c95WojERxVcmymrKYXxnlSBaQ7Mxg8mFBHeOBM1IAqnsNfpQF6Oo9z9dC9Xm3lgC
4FhrvFDLSDUaw4tEkCCjFFvEPHoiMI5TypQIik2yd1tm56t4hxxdEFVrHI2uc7T1
zoM0MDilK/lZQl1pBWjYYmJCgQ82jVwlWZqMSutiEMCIJbaEVLtpXYa2CInV6Dwm
oZLkUzC1MeobXGTd3LCSaEboQkNMrXvviQhZH9Be18qzhN+BhjZe3mfyu0NUnqBp
EVcNIm6DzHAzTb9lpKuiQ2+DAlKslnlMkfrBs3+CHt5u7TcymUlI/XSstpDa1uDH
d/7Bwl763wUif8c/pqAbYwPktvfCz0OUesadYr8CofSDg1yaph5IojdtIp7noe95
VAz9jy4Q1npQDMCAer7rzwu5e68pM2DFWfLhfj4tQUyOGW4LblYMXXk/R4WN/2ts
d/PTB4yeF/d2QEiPK97aZMEXWmTLh+HGM3G0HcG9rmjdvlK6xgDk2TWeobsArYgN
K/uDDN95Nvp1RvyGWrC3W8PppRQed2KWqhuQ7EfJpBYytV+y27Non42wicfG/Eu5
jJ/OlKeQu9fWMkLf53XwWqUZAL/Fp44VfR/UQIK5PjQMWdaCVlJQeLsG6B8IDsRW
PusWfoNLauXP14NBCeKcbA+lX8KtzktMZep25HpQgbd9QBwtnyKOmCg28vRVpAeB
fb4R8Rd21LItu6nS/MCydNBnSwr1M+LbYWJzN0NsqjU1ulqrtLPoPGgRu5UOjwdM
WKNnVM15/ihGGa7P26TIgHyjNc0uwcVPNqra2bywt8aGPX1+IbJneAXNXODl7uly
4oBde6v5SEkj+qkoZuGfLMkiLLb66+MEk6PZhPcqjg2iHpi+b5ICfbVaQ7eNDwMW
VsuTvalCM4sWnSmVVpbL7qarY5OwlkA2OE9ftuskUQBZ/JWxc1PwprMUuSV/4rgb
AfKdYccrw2FKkrRLxooEBuICVe8B6wZFPaTRo2mbFKQKJYLKEHcEp2NpkCKXfZQ1
Z1f2335gBW1WM8NgIiPl7SAsjW+2HHwmmGLQWC3HLEu/r5Y+zNEmbIilVKS4sBvS
llCwKi+OLl2o7DAzwHFlqYtOyfd3rwP0xymnT10Rs+NMTNR0OQcVGPRWmW0vDxeX
zZRBhuIDCHF5ceexiwA8mICjb/xZSQ4qdQ97G933PToSgc+9528jhgEs4YC+UDML
VHAkumI6zP9+XFhwc7xWewyw/tACtxisQPesvfxnkoUTikc9eN2QrXw2TdSct4v2
0kIucrg18DzO7JL0khn9zKELVf7b2al9LjI5TqIc5bIZMFV4J4RT0bnmQ22I9YV6
M9P0GzJPznsRPKz9iysE36Y9Fg2oKXmdUEVdATuq+YeRwsFR9QkgFGWJL5GJ8m1S
qXUtbYzqR6xXsF24IQbhFNud5dpB9qxpbarQu8cdCezKQwff8CmoMumFxfALr89K
O1hRrLuXXGbES170ok1r34F2LS7BMSsVopNH0dGRjUyUIJX//tuEsp8yPvHyO6o8
EooTFQiuhYiubBqqz8L7jQuw++0tOd9JdIIFi2r5A8BLlExrVMZ3Yq1/S1MxOYNl
e7fZvacfaeW4o4Pm7tWUMShv0NIgUy9DIWJop6KlXTLsc0GDk1kbvodZiPkOAAoQ
/NL4phZI6xPw1hZ8G6xg2bMaubeDf7OiypB1qxlsG+fZ2I2SsvQ4abOhnny1QIC8
rroYX4bQ603KGf/xuWv3+p7A/WS1Yl7bsixqabdHyrZRxePvEc0C0Qw4pA8MoK1c
qcK1jto1W6ev7lWuODFmb/d6Az0228AmCPUhM63S3klG3QDM2vYtFmcwwNkx5CDm
q9fnRUMJk5ksd73CiUzQxIfhdgUHPtkFtyV/VoTr8D1bvjizOeGp4JugpXc/X8l5
+NMQtq0FrmhlXGsTEBWJcGNxuLycy+KfrmuNZRi1YQ/wI+u9EtZdMI715KTMQFQ6
aIPpOhStRI0XUx/WDeO4pV1Ucb6gboBgXUsrungie6c4lxWidQUso/JdqXjQ4GIW
HC4olASgTbvuGd9CNHZYRkJ3i75pd1kWnxdp/RgzuGCca7bo1RFZEqD0d6rqBzRz
//dneYAe/ZdlXkhCE5HrOmJ8WWBywbhPrrjerGbLm3KmK0+f7WAazUnAgCEITE3E
+fNnP8Rn7pbdBGmdgL1ErtAzLy4sgKiGWNeituIeK9gNgthhhev2hxpKJtndjsOW
u3DFz7c+K6pGWl9jhsmAhmKXiPlxPFPl4YlOVtoIP6H7lkDNCt4jlcwxtiaEWx//
rG/0V4cff+MHCVAsSeFHhR0NV0YPVZUIxWO4uc5D6LDCLMpASfEPZUupw2TgiCim
OYt5XgDiL2FbZWxKTBOQDbri71JRLDyp2lHwBjXiJ8GxbqmAKV8B0ie8MV15aRPH
ufzcxKMqmlo653AzeP2ybEsvbVRClge0uCf4BC+5TfqQYfu8nX5jM6iyV07VhNDk
OOK8gE2Q6tFUkqmGp39E4FLFIhuyJes9NcloeOnH0r6kGolwWNXTA4vPBDjK3Wwo
1evgfIfSOmkssnxdq7HXxtawL+9716RSumTZmya4knkxXlst3j5AgKCJIWX1g9Kk
sE12F8yv+kL9rT6ucZPoHnKrwfMBUyF9cSZAb6woSQqjIhz2zacJNpQnto2JKdbX
znYSLbyAKZFdtvnWDdQjsdlus3+IL8L56xtmDZDUF0opAcTNuL4HJ/tIlEKvnLNM
iU8PKT6K1EDlykGwMUMAuqMd5kJCUhia55dvDRXEIl4AWlSLpl4I1+dREBw4q3uS
KRwVaNN8uTRdVQhoq3l9LwYF0IUZQcQ7OAvlLY4HXhD7HkM04RSnSaZCpECdXwO5
LqUBiZ2RuAdhMkN//pf83w50x/elqqp8hGP/NOSkdZkyUxsm6xcb+82Im/DpPFbz
a9R98+z4sV7X/pLo+YWJwUdzc1cRm2BShm1eHqiWmjTuFgmiWYxHAccRJMGFhmlW
6prV4BQ9uor0//Uftzc2lRTGM26U4OTnHDZ768XMn1vQ4glgZidwyqDVcV2Hzehs
ba9ffk7r3kGglRnYLZiVsP9Lu0lxViSDaqWuQzS+wq4Z2WTFmr7y7L+IkOgANSwa
TLBJd87QUF0qmTUOoyBdOoKwyPBiD0n5MrFrNMFMVGc6MR8doxOWr9tgmJtX9FnI
8njfCazarbcxsAwg5Kxco7uESYGz0khrFr+HwcQoZ/Cr52qHUKjPFpet7uycRne5
9yex5Kh5LAVZEzQYkLzPyDRlGTnwXdgHYwnFjam6CsuMSCKvfVN7xzflWBUJ46CC
GKXxn7ymFUAkRdxBKPQFuSt5xn4A5GM8YJ6Xapq1tWO14EQ9GWWEAa3PpkP2k+8g
SyS+6MhiEzjOt0DhG+6rroc+mSX7uclWrD8agOQDvOxhmaODu0Zz+C6VH8XL39uK
3T5ZVdDtPnuvqaYkTtDKTQMmKeg4+kIIBHgg4/MgrZH39ujbIRTwGTO/rHqC8H2y
/VchA0gr177TNiLKf2Brn4L+H62NSveecQG/EH7IXGyPNld4IRB+NG2UhMT/v6WV
0aLVfgjp6U2ohDlWpeom8nCyd1eg9XuIuUfsh93eQW8gWnIQqYZAeP0fsCFFTyeB
u/3H1ZvXIoq5orhZl0vRt2N3zNIQqxB3ai4y7bgKjxOWYxhB9E7ZyLPJHv5w+zHt
0U9qGpobdl7d7J5GpMTBMy4xqpYLya388TYgyu+ln+C7moKuRLhCvizybmdwg27Y
VE+WqTl9d4Ek5rC7L1bNuY7hqRoTj09QSIEJkiRBFVfmxZJfsgocXb6+tq4xSX9f
4dj9JT0qSUS//ugQqtHCWZFhZ2Npk93cgCF6OxzSdUeV2zUuhQo5zxqCv2rdF1fw
JTcZiyMMwVCuXdDuAiBCLi01Zsd3k+siiUYC3TWHUFLJI0K7MUxWosMrv84ST5bq
hdUOjD2JNb8eTEYobC0Y8E/8kwtve2ycYeVmgokgAnXvIE0kwH0q7FbBlFCN7KyI
zsiC3mAr2eHIgvpC5QTW2yBHsC6oC4V8nDPkBdQ8F9eBYDSKDzsZYD7ZDM3v1PwM
GiTX08+E3zs/w0QezkUircC+TbjsOCOorUCN7h9411i1Nk29ZExYyghxjBaHPG0O
i35+3or2oL/x0Oy+h141c+Z1l3w9YQdp5QQC7kvUToVRihK2Qmrn0CIgETGDdJqK
KfaJa1HC39Ef6uMbyMjKtLUMlK4bbjRnm7it2H8GSoNm4ndje2aHSLAeCj0Tku4z
QOA/2CvIgb6zdjGbRD1FIiKPAFxhAVQz5P/nCTfLtJ9jWdd0Ls6pwI/xmch4+4aq
t29TVASL61A8LPVcfZxtoJA3yfrr6XrjAIyV3o7UTPqtKsOHJu4naGu16/WH4S9r
6MSkypefcWiHZxe8q6t3zXtQBQuauJNSVd60vMapaxxaOcowWWeO7xylXafDVxTs
S0pA68YhrXxZsdBJa65vZnjLr3jbZDVk5CQgWQyx6hEI9rJSKlxTLeOoDcpYxkrf
TLCErpZjW+fM8TVB/I4ya9GNy3ua5V0J9iiong+JWHRNBlHvNKyNUu5cXOJRiSE1
BmIP4T9E9gpN/nkf7dVRB8LXMuNEP7ycKBeAzlc8mWHPgWsnDysqH7Ye118eikXd
HsEJTZfW7jvCpxD3Uz2B2EYAYFo6RwA9f3/xMgdf8L2FDR4DGxZzXZrxCCgFabP5
i7rIcZ26u3fVGdr76/b4gkFnuHC2veuUMntTFqzLfcSkFNzTu2Tda1ccrUGR0M8Q
GoPsvQGkKfFo/Ys6gWIN+MK355aUliop9aX8iq/vcyhUkgczdMeQKSsXqwz4L5g4
JgzAQlCBaJhH0N6PET/V3gUhudSVl9aPFpUZ8ovzznyDEq+UJtjVDjKDV5t95f2a
Ht4mTPWmXe3E6Ya7tGJYoyoMZ5BBTQ3gojKef8EcMwM5D+qN12Hv0CBDzuVuwtiC
nF1X1w/h1fzAqHmmsp4kjbbJUnFLvwjINx/cHCTb+KLUZiwvZrdhBUglZhNQmmjQ
HVWG3w6NjzM6VxXQwx4l36n0++vm3da6OFQDuAUJloOz5oXPX12TZfXzuyuB5NEf
dWK+hHwqTRn/LDoWWxUS7UMPqaihLJd/VLlPvUg4+XjDq9IVFGhUbc00OdseITy/
CM5Go8dy0m1ikoBOAm2+2pBvaA15HtV8BbHXC345IuTRFVX2iNzRfdCDYe2i7k2r
kfxUZVoVu0g2TrBol8HF4uwmVAtteAui8bZTIKrcAcnILAxPklqXQqAxTtJBwuf5
MqBKSj23cgqRapsOP2rD2KEwIG7VQGs6n13u4XfJn48Q8bD8Hu6nK9RA4vugMl+B
Ns3VccmE67qVW0fXllGgD+2mmRvTxfxHcdHJcW5fOq59d92ne9f3flsLIGt/5PF6
gw0pIOQEhyOBv8E3Csg41ZB2AHcBQ8DWEcFbWqcBc+ukFJo5W5qV7RtMiuWSv3Ss
3lJNt0RKFFSc1wLXO67CwQ2mFKbjrY2Hd3tSoX5P0JeMDLm1uApmfAg5w33ZaXUS
9dQt7bDLMTtAed4NM+j0fCOyYw3/jngDq7G5ccW+nKSUhKzmiSIvIlPpmfeiCrn8
oPzjFPGfLQ4DtiWOOUPxifH0jSFSaUdXPDxZfQlJT/aaUVCEBVYlvMkq4jg2CUW9
88z6IMjamOrHDSuAnNk2viu5u0mjSIOD3MEaoiHGEKh0g0SNMlfCDfrZ6l1U0UFy
rHSnhfBe5WO4NqrOMIP867tYxvJUA8JfmVT+Flq2WXhNq7JKDExRWP0fWBV9d6cw
XzPLmgcuqpFvZFnH1oR9QgW8RW7fJ7ISa9yALTdCxgAlTanQB0m/Wo3lpZUEW4Ei
27BM8MM13NUaO8sKHBivGR0MBqQF2j7jO62NWts76ER4fyUVeErp4swdEQxjstuM
bHxxdD7OFwOi8KwYarBtP9O+2EcPlpwDNfy/MPYyen4NZ3UBWem9nqik/FX0WkuH
yAoGVMCVQEW3kDMLQzCK6K2OLr3rHWVY5yRLsp9ZcNx9kuddCEtB82mraA/dYiNY
SB6diaiKfzr/8iCOmeqQvrbVzwNo04ANIX6AhQt7lU4dTZD7GDscgIukmXJJn2e/
1gCS4KK67MjfC5sMFHDOfZz+k7e0bbggWGKU05D6zHxOo7WEIkatw5l1hsYdMJ2F
XeLeOBGVpl5GKB2odsUYegtmIo/FK3WiTYfQLI+kymhJiTpKcYW4oC1rUlTstdL4
5Vj8OA4AoaPl+PGbNwZnm7+DpyzdnnRu8FflA2E7Im+qnoFahIBMqI7tGVm1IrQf
a7NgrP7qHfnPez9pf62w9ynNLJFYnfZLIXlOaVDDqnTm5rpJVnnpHgTDxL3eoWkA
R/2jfxYZI7FQSZ0J/yffbmTbRMjVXtUPPvplJM3iWD/qMAlpiE4QeHh/TcVTUOk0
uDSef1g2V5xWL12vUmmywYjXux3xbIlULHZwwokAMSeHMaz8PFEUXoKzSzK+Cpz/
PidxaYIMWDECES6Tfj2y55xtDDN0wrn3PXluPLs8MxybbAXLP0G4GbLESFd8BpuT
2njlFl+17RXwZIHKF/VTbAWlINMVGx2VDdhAKZ+PUw9lucu6nLTAu9jWV/l4eKn7
fBLEtEeNz+uplj8ezfm/+gUZrLEEtdqJiQ6vOJ4/xI3rHu1NDVF06B+pUY9pOlVO
b90EaNhgZCzAu9OLn4lRz/LV5+nbiCyNt7cW9vxxriIRxd9iN+3sPvQt9XSSr9mB
fySCl9aNNkN/bfx8ho5hbdcgfF52KVBAyTcu33GOAdLme+2yFnnbGZsVhaWDby6V
dd6EitB4rr/g1+2h+frYcyy9w30ceQYlsM6q717Tbo5PMbQaOruiPIl1AbQsNuaj
EjNmhQ7B1Ganffm8jDRLHNQJyYR8oeZTumc3XAk9OvcI17wsfqLQskyaWby9DeUC
nqT7rVh0XBG4S5ttDjRtWoYMSw76B7cPuFo5VGdX3b0Acsj1EkMHPwt0WMkBitDc
7hKuw8X9AbXOYsjQpW+3By/TDgiyhNTYW8LXIUSVgsnu40zI+TzySNjttZSzz9c9
hReTFonyDUtUZXAcReNfqhcFpA3nvNw7jq3mVE9lOX6O6x5RBsNV2oDehfJIE+Mw
tSu3DFHyn+uc+Gb4b8gYh3AIjyFYGlJS7IjNUmnFaLweT89Z/ResJzt/NKWORIap
dG+QR8LQfG0/xv7scjmv9sgg7Mb5urkrnhU57SrONBMWAvF5uzjC18J+wF7B6+fm
Ae9GRcjQ24XBedGNS7QwYNHSSfKJwLBPsNF6hU0uP1oaSbrcaffHTcq+gEYzR0qZ
NeU71Q40JqlwpXuWdJZmydGHZUy5F42IuBFBkahtx+WQ4VDh0C138IjO1nFv2+WN
J4f6uvgH3v3GAgPEo2L6h6oMHNuOFGU6qrRNnuLhu/U7Mu53YTZC+UVd08lMZWaT
4lHPxvOITfHYG9lkYpOfijFEb7KvbxLt7q10CEF4JD+8M5Tg5EPjCjQ55wisOJl0
GeeB0hztgc/P1SirEomB4c8YNLP4QrhiAylieukiSJDrDXUV1ojWob3aPqf0wt8F
Y7HPaH3nE0W8Jywjimm/Qj/hpJs/sc87gyAwEd0CRvq5Dg3QfxiyFwFtZHXQ+ks0
tVObXvnvWgNPzpCaTUh3GaqRATOWSI6aatCRHCOE+5Um98w+9qVMcQvvrFqzZQ/B
Dq0Fv+Nmuk6hWiKi3swltuYMp1hphX8zRTQ2HJwxEB7cVfOTHF3jrX6VfMQ6d+5Q
8S44gAp5slEHaf8/XPQxeRe6BbsNpXTx5jsrB6fBsGz6uofvO80aNM3iN4FwVE51
UhIEWTgOEJ3e8G1QPQMGi/meU0h3s9BuvXkh1IQ29nhfav2Vm7RzjLjUTqv0mqiR
U9ro3aYBFR0U/os0Ok/9gnocoTxPrMuHK1VMY9w5P5Fh2xkSzOeT8uQkF3LwRcz5
6AMaezQ6I2z4rbeD448md/xmDPav9NCVXe5+LRIJ9E312mrvsjreHNtLTFjC/dAI
8XoRWtsxc+/Yy90QAf4I7MQFfCAZoy3dQnMDKYXMb1MEYKETxdYagRiOfO0iP/P2
MzoD0PTN/vanQch+7WDraXqRr70lUPqx0Fr9EUZuyu0R9epfG423xhG5rTZkQbwX
4RuZxUnIY2B3jrsGqgzNOZ/3PL5bS4KBYLho7wG2TNBlFt8hXCb/lc3uQlOGSZyE
qOcZ+sI866FC2+oBrOTngDZdrcMmjcHL7/tdn1QFAsUDgRqh/NGuXClpGYttCcC/
lDmb6OfullVLHh+q/tDODit+eRNgOn8a8mM+ozuDk/fQ7eU0d8jbxcFEk3hfG5Tc
zlYfP/JC5h/oDQ3xLF+oP1J7ebJ2G5mdhLLUlBwUDkE0t/f1qG3bpNGEMTFpjrGB
bKuQsB0lJ7e4HwFL3ucfZrwHtC6Q4ExVpPwk9tNN4SP2hPe//+d/RL39Vwj3kT8Z
2Wj4vvG3G3ueRohVffGAUEd+aCULPuYOFlBWOqJ8Kgi9FsC3pX+RHqZYQCsogDRq
zOsUrBVF2YjZni/jwSazP6FZOG7tc8yybRvfmUAXmQjmzpofhi+PLDmFI6eXMIq5
wk6Yk1ePEzpv7g8QoLf/w/Naefv13ORQIdn6RCFLmNzDNxTGPQ2zgKCuTfFcfcVL
pzf4P4hY6NgWUxdq9OOnqTxYuoMqU8LObXqstxTV0VthsgzaNpVryb2p36xb8CON
FxUKFc0p8V2PXNJjdzFe9Ezp6xEctv7pOUhPIjMEu8G3AOt/6jnh4pFhSHOhJRGs
OUeC10cqkzd9qGrTq+pYDDSxdT4dCHZrTjCMeGSqZUgBQyGLvyDx25Nc9Ky3IR9Q
EQYz2sZub3idkHic5IYGgZDpCmKrSW8zMqtm1KE/w05HxjdlrjL5dI9IrTDNGFx2
Azomh9+Oy9RHPFS52a72tyHd5ugFUHTNJ3Jo3NzybrQuWTROR5EA8L/bIiwVrpuq
y+CogqpDNRcnnz7JbRJ+ZT3Ypf6rT7p5ZOfrRMbW0xMrFKRL4m+RIhFkmm9SBLrh
rDMU6rdUeaM2Gj4CxE56GsmjCX/EVQRfFYsJxjpvSvuyw11KxnGCJMTa7UvI/B8q
SnND3RUsxvGfYm62qKhmLB/yjlXgLp6Kxz7Cg/pYnJixqp4HTZU5BtiFkdH4Z16G
ZIuz424E1vlnEMTGhR4YFD9jdAbE/uHufqOx/kEQgIJv7x4uLZOzMS/GgFX2bQE4
ECZfEPbsMw60hc1XHF+dO8slRS15wdW5Jpiw3qFce9oFIipp6LoL4Fi9YGN7ExTU
lVfYgtCzib+7nQtYhYX5kRnEGRYm/pxByWz4V1ME8sM7xlLp7j+KeER0Da4d+CBG
3HxODRWHaxQt5HP/UUaTopbTt73qSoSsPdUQ5NpkvnNwSuFCMLHbe4Nzjf0qBjG8
eFTjdQnCDzh7thnVllaBbLQaSftASrf50B9Akp/dl0aKZc33cCrOt12OF1bIkN+i
j+ej5mVNVYmo56TIjmiXGCbtaMBbT3jtDCQPFKl1XQz1yWUiQH9etEY0WWcBLU5u
5JpuDYvkpuCt+sXYFShyi3iSx5qMyZFDoan4djFNmxXYZABqk6OSkUqQvMiwf/zz
66qZfsELLdbUv+C4IJ3icv9gERWnLRxkJtxsh1q9wOknnCBcZ6nSNDxzvx9VetHA
rVXSSb9BmXYPhWpbkKh551N4Jb5eGrL8MvgMH4WBjnmbGgP0ib6fEatQ4fNgynLJ
pVXr1DuX2qFhiGxsRl2G/fb0zrXbgFwGIpHtQEx2KM0bZ1MEU5yjbullUMux4131
YVw+0MrO/OHi385fG6bH19K2n+YoQhBB2m/bHXyGoPUAxF7iDOP20F9AaqJQHXjL
Iyp2o69Dq8pjLt5w3QMDHS3maWLcd0Q1jaqRDG+Y5pDFTFQWTN/MS5xlLvyvxeFk
wjMW5WgFvndFp10hqAHIBTMiQvdu6pDF1HIvdngVDxvJcjIIxaYI1KodhQ+oprSB
IdwhK73hwNxpztqSUTiTrYvcxHVtD1/xtb+07vMxpIOIj9Fnm37mI43oKmwgDkuI
rhb3SG1plM5pDpD2YBbWgOF4eR2uM+vX7t2ClEynoINF+qQrZDCa7YmgGTE3RZ3T
zDMFvevNBMFjx6doT4+yRUo6ypw8EerbH+0K23Y1C5cE/HteSx0COTODA93oKgG+
MSmzue9f4mBCW3j6hYlq9ZOHaFw8eYhBvOxUjmdzEGiHb4Ny8qW4Ru6sBD3jiChp
gBpclllYsvp/+nqdfvaPeCbCydY6N1+N91Cce5HcmPI8zFiCHJoPNuBuAVJqn+Cx
JVm5Bwen46EqQ35J/KWkeTE5g/Cr6Ez+Bwn8YxTqMFiwpDCYYH9MY71HzUN+iIr4
TaDaSs/AwoSTJqVzWpvw2y7Z+ABzIVdXmGE/27DBxFtjZSxGyjY8569XIT3aQFBW
xa/D2h5f08oqJoubu1nGYS1ntX7coZlsOOT1++H/LeuCOjSykkbjtbqyDzXuIpQv
jpZ0ggawto0H5512cLF3KsSe3IT1Og5WemmmhG6/wzO2uSy3J2QXG5zXkUu1l8gt
r7kMpNE8M8VQ8Ji75qjrPDNFsaruSZPLMZB34vsPBJkcgP2GoxI3jsOlu7flqm62
NS/x+xN5M6bwOaFaL4SzYR6/Hvd048fzLAsdnTjmCLI8BWSlqK+BMUyAsMO/Wbue
4gvnFj/yy0d+3n/I6jKIt/KqHvVS7ANzDH7JXd37cT0dLhaRvBn+IobFMYOW7nT1
+5E8bvkf9d4j23qK71l8BgLrliBy25Bf4TY2qIa2+ZduV7ceejZEAD1oeLafJ9OM
Qo0EPot7JqpcI9TAD9O0I1VYntttLrg7vuE1apXxEqqFg6McA4Wt1tdwVk8XyTn/
QBdFQ6OrfvWufmLwlYo787amLIHxnFbco596ziCh1wOYzDQq1xaMk9v/vJCkklH3
cNifTNPzYi7ELOn4g9dTY4u7NTKQN7LfjBYPDcSvIKDrQQhYaTjY2t0JusREE70c
PdPBHW0eJT5UkkD+/1wXHRFOyEmpkJSyMqNEGueqkIsmzwfXOlvmTx/31sUwCsCX
nA7Fq4TJXmg9wMn7UgqWr7gzWOIHos724uyf/oKrbLY2lnkfVdKLHz+dnkIy1ZLJ
wRahLOzz2E5/2N4jThaSjg3+H/cEa7yn97W3RUIEq252/K/zefVXryXP5zGiKfs3
0Y/LJ+z+xS9s/1UtqbO86DsiKCpF8j8RKbUw+pIRrGYaxNtWnR3jJ9yRxl/IOFdK
2qTOH2HRPljgex+f+Ok1OEoE8xEPoqUzGGVfZja2dyxyrbVFdyR0Bvfv7OJFzUVf
co1DtWYaKB6ydSlecAprZuqkBJiiTZa6UYesOWO8BmRwmi/RmkoxA/oavqNJ8nk1
95qgWDjd7HQAWGjBZ2N4xZn6rUWRud91TPD38kpEPlQVLCLMrvgCOKsoy55rE9P9
ss6Shau5iup3wkrGXxmP8gpNGCCVOAxisMt45DxqKAaVelKycvD9Ei0zHi6Ttk+X
Mz62zo4ZAumDHDRBHEZwLR0WvuLKsaHwI5zi6itAHVf7M7uXD4hFZZk2zvW26o0m
Eryt+7AZ5ch4tzrTq8sE7XIoNwFE1F1AHHVHT8qoHuWXq5NIcrrHmAFWDmwC0aDa
PIbVeqPU3q2xFW3+i+GO/PZy8ZryIjmqhDSVxdGPox5J629l879G1i6owIh/IdIO
+n031M+lEhT8QmCCCbuMS/Wwp8luRcssDj9BNf2c7ouPR7PLiThBJ5U58VAYVxl2
VPy7nelD/R2VchEuiVK6+FdpRxugvWbaWZXK0e7gZazkLCK4iWxEurWS2X1cefxw
e675uk1uvq9BhkLry1lDCFUoplUPBJX6qHyHXfPKJpIA4/8zWEHyaT4e0yDjkk+I
qLRg+ZhcEeIn+87VE/ZEYLzLHl607OkBO2908v0bATJ6x+omAJO9uQO8rMYBpcc7
E+3vdMtAvmQMf1LHB/c7VwJmtDJcoGSyWtHZ2X15wa+5TOsj2RrGYsnHawtSU4gQ
asz+t4O2ogMZ24nFr2GGNSavkzHiLnhtX8KkO8lkMxKLffgccEzjpNILukBU/34Z
liW1YKcXEvYWSsleY8eqRVgBIS9L7gF/EXJXvL2TYmr9yFvzDpwtDh76xOM33FOm
zTUVAF8zgWP0f+L5gntD5Xtal0qmiOFyL/imAh/rQQ9mXhvwqmnIiAcIWv8d/8L5
gZpjDUkOmDnbO3+UIEb6BzYgP68mw3bfHV6xIBnMCNULmOmgSxkaNcVlx7oP5phx
yrrN62qtywI3Z1GeQAn7peT+vUMiDMXaSYvGn/nXldSEjvnEOPpayhcmERzI+GJ2
FtP+PbQJmBlpjdt+vs2BTGO8aA8A0BSlYDu8QuItm0E3DREdy7ZZ4ODu1kDu130F
2eCiKiodrM5fBrqteAVZ//VsafEn46QifU+9Vg9stYQZzt67xXxt+ywm/rs006rc
l0nxWSoyNYJv8HO5jS7TYEmKGt6mL0nYkUkot61WNPB/KXCOudfHKqkBtbXxATfw
5JEvQTYz+M1o6tpBERIt4koK6oQW3zzedJBgSUdQfu/SNBmD4whUDj2qwilkqKnY
Pg/TuyUHX4qN5EgO2sO1aEacey7wK1jh1bDH6FIsZrbAslVSO+jaXevIMwCl6lh9
+NPVhIfmuBac75aV/8zwbWiFuJWOyhpjlbXaoL3lJFRe9uNKhejDkzJgSKXBfL+8
2f77eL6Wv2etFLfG7W9PpbMXGRexVMkE8LCQgOlK+KP9gAIALPAxNzR928GuIiNH
VtkCCvinvgGM8yrlnGUiCA02Oe9esQb9vMCF4Sxppaad7999z0CCRINDNpa/s4kt
U7USVl8YLwCPlvtYAqsxmpl4Ld3JjdSudmAOqNhSNjWzIo/PL4P9lulMobTneNwT
DOLUz3Z0r1qN8ymdEpnLD/VesPNlaOuE269RZACG251h6dfoaWk++GPfOnNLdRLF
1f4H6XauQjtqxBm0I+Jm96N8pDJs2ttm/srvrOlaAMmduNByYtMXeLr2pPrZTAT1
JPgH8hMg787XuWAB+GHVlE97LXkLE2ZqDYaCrljWUVz8v4K7NUoSgxlI7Sgaf3Ti
ZOSFQN2yy7E8ZdIy+P7q5DCZFsfBMYHyvt5gKUzGj/tL15Rfb1VsUf8SUcCJpUlL
Wr7unsUk8TJDdAUHCndIhgRgUIHtTGeXe3UoT4RcivlCKiTBEFEmR0SdOO9zvy7c
h6wnCLUreaTNyYWRGKOCnK+lZRqFGfXypAD818zAQKItDjr1/n+3w4P/y7BSf9j3
Ks+pbhRCVmHvKAJAfScz3XRpPjS22xJmfj4vIbtPFpWu4iKvzXM7Mv8q1cvbDD5k
DnsE2rJtchq1GA7JneSZcSP3I+1lcixtH4cJxoH8YOFp/AohseFiggz1pbJHRMP4
5fdCwYAbn7ZpkED7LC3SgBQ2TthtL6Fa2OsOBbCoSlmYVZ/na5FAqvUtHmv/HCXc
T785ri3coEK+4T3J13M+wyG7czhdgvyKOL2b5+CBEmIEdxdUs0ppPqMqTymgBinX
CIvU6zGtjjFaY51rDDdakZH81PhI5mTwG9gNS2VDN8m3YVXEWTDVdgIxpHnsEBHr
41DFfmOMso7Rtqu25gmRKv+TjPQIUPmEaVbVeaonEzC3y/7+sG3eoDe1JZfdYuxv
V7ZNXBSNIEnHEohZoZzF/t1I2q9BhV+k8UX4844GNt7yckytGclSezxj1glFkfkX
3sFdqbJQhflGB+85T+p/FqEjSJW1ZXxDrQYi74kDLU49rV78jO/0TffyKrTQW9cd
OaEdpgA3B72DCm09JZxWaf+03ZBwUta6jnxCB640DsERE7WbDG/LpR5Qyd8beiUq
gpTfFr34GHUR+fbo4TTnN+VoNG76kiqL7HxcBainPUyxysFKy4P2nhc/vuw1cJdH
ibQK1tCD92TTrUC5xCpxLhImTcTrofbHUNsEGUAtwFGt6zhABqvzDFki63pT9dSO
7++jzFMq5PwNIYLnkzBDRHnc4SYAhRG8Hb2MOBYA6rd0mG4YB+KseeWAkEpzNLgR
K8930ewo5jrh0kVnxnXB/NYWJw8Ei+hs09153/DV0dqFva6mtSbuxOFf1RKxuaP7
icyjy5i/VsNSWnrUH8W5z1sExPGtgFnET+EiSZa1oJCD6fsVeI8qPsJ4HGVK2dXM
mVYLOhqZt+pJ2Efq1dNSQDgxG9spyHXpYW+nA2GpXHkUXtHZir+oNg/nekAlWxgJ
hZwRYshZave29ZRDugXgLN1HeDHnGw6vZ/Qo0/rqjwpXxIYGbNnhb0NKyPVeOGFf
6xJoeBMBvVUaXSm9SA/eHsHpJeBmc5dHrcrVHkI2kHDC/HaDuqpS8uh3HDO1mVAn
kEfX71MX0M5hTNNP3weo6m+iXur312WXzO2o4e0BxBaCvjhTDXSzj1x9w5i272G+
tkzxffTHdmhxef4N4DXT+mCMlcGCoJIb/KsOh/ThHpD81jF2I/6F4qvT0Ceaev6Z
KNzaSa4VQsCNMoHDLZ2sHPK9uf3cH86CmGQs90WivWy1lMSKUVnsbqWmRTz3JauJ
HvPe/1rXpReaF/i7vi4ewCsg1O25wkdV4QKCPhK9k0D+KuPJoanH19FKcBGn7bEw
aoqvUrVvuaiEnNtcDITtJN00wp1Vj0Gb3FZ1vwvqRWqACqz0SZgLoqfF2FImCLnx
9UIaHdG+wCG7Fhx4BH1wUQJPjeNKClgwMnjMWyvykmXD5Ez7uLOcTOCeos2UTGPZ
r7NA2NI9jy24yrmBDIAPb1NQOadb7QG/60oPKND5a0u+KSbt5ksYlqthDU4TkYVq
RhcioDMOiVcoUktmUlMTNLgEnKgKgTwFfTiZwPBkI4zLvJm4tx3SC+honROejiI3
4iUHzqmiSWljXRIFhE0/ghNWJReRM+JUgSDdf3h8avapmRF6cRrrYXnljDtXVnsd
3k7EaIHFDe4GRmtdKXldaSardH+DcnVm9teu+xFdlbjEAsbGWIBZz/OcLJLxtDtY
foRuC0yvi072tHDTgH3cR8QM/Vw6iVPUGR0QSV72f3r6fZWZaClxwLAkIkz+G396
cUvMgfQI9+Z4daBsV8XM7kPZo1hng0/CkhRzLGsqV5sCJPO51oE6ufsx2x7gu/xl
ONue7qYrZ0X8g4bZZqbZgpF4yg/VLxMDLnHk100Uc+JiUnN56nhwf3QWG++Z8RyN
LxrYXI29LoT74N2Kdz8Nb7bv1AvbdR2iCoOK4sie05R71Bk+set4w0oZ16PClXgv
VySv4MFogqBRHTzpNff1I5UxyVvOVFhBPvznkpGXdp3uD4sT7akJvSmgan+kjCEP
jWi9JHiZwEeJR3kk04QeRE+6Ly3rGfsFVbzqmHAKKa8InL7HqSVoOsVSHXx3bmT/
A7tIY1L/3QZfGlJyowgbcEKnV46RP6JxWg2E+h/mTom0q7Q6/tVGrAyY4/xr1jBu
maTsSy8pprw+bXkqBf5O3e7+ht8FzSSNf5cVRyzRXrt/Ar4Bo4jKIhQIvg3vaee/
MN8TVUcgueos6TUZxpT5r4YyCQRkZipDMRSPqHm+2Sj2MSiFzzgNVGsIfQ9vviq1
v43yshjHnC8slBeIGlVM/prfBXpBkXiDjDvCHRP6e4YhsImE4IaCdWkyifwQqwZM
N52NKWLHj0CiHL4grXcIQQvE45+iDFrONoV/X+vW/Jfv4aArMxcc2I8gFfM/n57v
s3AgNRqwLMatNrBQxZ96pNjnDRvXJCKR6r4rGGdRlQN6uPa3fjlmW+EEgVE+eTE8
psx/FN+CZIlR1VWBGWiBpTRZ6B5fPynYQTgXwEf9y68tck0CROCvugH+Hmv7iWRZ
Q8GsaRDGGxiNmMAKewijYe/37FkJTC+RLu2JzJkqWN9G1mVA1a3H9DY1MEICc++x
pQUcjro7/xTij+P3jza8I7378nZkwz36ilNFqPdiUtij6MAjx9IPtwBZ1/gtVqR4
xjP+bJajsWM+YSNJivxS2WcF5ssyVx69chNMrmUCTUIordWSBTxLF/vEQY3w8+DU
FgbEmqZod8yFK96b01SwrZq366ffCKAP8IrrTTAzQ1hNCeWCQH8sA1YkH8gzOOhu
RSanxV+fl+twFV2Md1vxBTghxmkgcgxMhsRYyRRGu0vO6eiE9HGrXANNXrud1gwx
PV+fDWDqugvFUJQ5geSyX4jepBfsiL0VMFmO985jMAj851yfkuxezNLzx5pedU21
5FwJq84G29pu06oA2Z2gu2dnS72Ba5hTRfkoieuiPY0ME/7bQ7i+COxHgO4cqY14
HOVDGTHifF2JbEufq8ZJpX6XfSanAzpKYGI0iM8WYeiqaLgl+oacWlUgKdbkuts/
5q8Y6KkmAbANt9/Agiatw1X1YTAOInL1SDP+cMSu8hL9lnvZKZIhM/MqAkMnxQXC
q5gW+cjd9xiEh6ZEFn1pYSOSkkg4nQZieOedNLL/WcnfY4Etc37YGRfyf/2KP526
dxLxtmNlW+l4d4Ka+36JtUMtmbZgHLiQrUZ4NphD1oL8gqIwkRkc8FjNXBVTbsny
Lci+47+/KhXw6IfPFfJKVld7Bbdwk+s1zICkj3SC0/8mv7TkQeCziJGMbAx65zv/
DayMX9bRqP4ysFwD9NkJitlzNweM4CdZ83tpo69Hf54RRJhSMc55s3dpwPLaIl5C
T5DcJJQfCR7sBKCRJDidtVrElMSs832rUGiJTnEulc9zLqyQJhYmaqJqvf+De5n2
cvXjN8X98aGym5fKosMPIjJS+lrjkeLdlwTrPZ/tss5fPQddqbkA41ehm3DwD9nV
6qTuMO40qwkrmQFW6PZmBpWL1nC+VF/CyOItsulvN10vm7gDX9e3mHyC5nT7pqmu
eFLJ0TY1bh77rWOMThqQBmkZxVsGjIORwXolkXEVaLIsgbygZS47pZAvVG/bxQDH
grvsQpRQy+MNfI+w20/3b4zUu8YRDQXlOn0bx0OWDG1F8Qb7WXxHotMSqs2iyEgJ
5tHduZg/fY5nl5HwiAGaSKIUne8gnbZAEdhejH+1mYuFzZT+8mSLY0fSrF30EEsN
7XdICUTkyLb6pDKXUQCVtHoHj2sInmmJCCY+aK4JcR6L1daGzsGIcTJwhsEckIe/
2H0PlNTnXszh3OCG77Yf+vBs/bmMvfiUlLb0flei3Y8+nvUXQ47kJZta/shbxv1I
oOXyv8geP39ZVnlS+vHGAzrtfLvYBnmagorA3GubKlObqeLmCQj74p8LiqNxQwXv
C1T3T5UVjrbnlCH1Yr8B/7qoYcAK/VElUsPyXRjNDJw7rFBzl+CUiUke/8M/IGBH
HsQJrlgRLiDxOIEb7JCGZzvVzUxvPmSr2HJvbAaYXY6KGMR1CTLi9n/DI7SfcjDC
c5+TmkQug23LgzFiU0KV3Zl0HUq7iO83OGdgR7Nnd27pqyE0eLvMPscf8gxFPBF8
FiqliHEsS/KT4YWYInmKqrwUk5TzDniytsoGpR/on2IqkH46sbrjVnZM9RJiUup1
itcmj2i+XSTZpG1kHxUzMsUlsjEcqzMjDaEwFkZaDLK1z3Eu+xHuSDsr7KhN9zrw
P1as0uEZPTY9BV/ENNVaqXwkvxkBJLzqSXSOPNTLgxGnJZGoKRlq+XEcEePwz+ia
bxXyCLjjfOxAafhB3EUeK606wY4RbUzakmVKmiBtVEURtntpaWZ8E0ImlDAUpbjL
w0d8z9jClM5JaDIhRjWxp4CH0wUPzPtM8ZMcg7k+jdpgTXt1t5WUQ7zVEMoNQLB8
ycPNG12M1tAG6qC54JjbE/mu3pTHVdXWQt9A1d9qa6TfQTIYdzzw7b1FkroUumpg
4tsi1GA34C8EXuKSOmmLXd2+Re9frCWWjErD08mOh49LmIVaBrT1Ude9Q8jTQYAl
D6uLOlLGbuPP+dz2GcU/4C5dxRrDwWsYIhMhUCBN84GK4Nv5jokN+7NwXVjFd7iW
0DbXsmQ4Rw67uQt7W2RDeIKVwD3LTlMFr73bst1+0RLsj84eNOdS0TpCVoYdBQPe
GHyD9ad4ogluaCKzqnozBjq2gcvzDWMOXzmDjhXr8Qj3qw5jPWJ25pkXcOnidchA
QM4uYYC3ANJ8C0Bvx6MaoUEll68SyTlk+BlX1lKdVUX4+GM8CaEP0+RncW9V9YPx
F6i4x2AV/xuR+9niEnNMg/4ZFOGvnm4VL3uwxm4B3Bl+giW32iv4ISTO7aSLPSG3
pAtYndsDlXs/4vl0zkDwIs63TV2g3e3xTtnqqc9d85aBVE5RIDqu4qZewjVF0vw8
G7WeA9/HMrjRR5Vhu1yWxmrehEZBqbsxT8ntazkzpQNLNJYJ6rzUU3kx8U1F9C2k
zady99xlGXoj4b111KEBFiagr3g68yXTLRtIDRy90FHyK2VVRaMenPhVQR8dzQo3
GtJ7kRu6wnAA7r3CBRwXKavUvGT3U0XLHarrB76L2rD8jj9ED9eSypfiVLbSI7l6
ya7VqBNvgp7bcJPkFzWV8hfHiOjWyD02qC6EVmXCHktw3is9D08NPtTJC/WooUdq
i9Ew8haMI++Lyy9qLukrLY9RyT83tgt4Ptn/bVWkV9A8/UNk2WrppZ0tPaJ3gxIU
wj5Qq5I3O4tvmf0KUTNpadrrTUJ0QU5qdw0rygv51kOpMhOvJy4sm9VQPoDm5/sw
msWvtkIxyvyEJVEI8AS6c8E4lFxQW6eM80uxtPNni0N95STrtdParvWyxPuBuCOB
TH2Jp/yXeb23IKErn9HniJ2OLbQOVVTBcGnGmRedV73a5ua1t56M88kDyalhONRA
sEstFIfHTAaYFqWkXEQtkw2d1vhYeSyMBCxBUj3c/Zpos0O3csRSzE1yOULr+Mvn
wF5ktofVooz4evMwIMfgsrTUHKPKwzfyi4bugzam503ISNtPwh/pFWY6zwa6ic4x
KFFboRt0L2aY5Hny0iRqoHyaX03Tn8Q07/fOozKmseFFA6KsvpbbQbubeONb+jtl
NOYc/9Y1qYM9heDcCh9sh+D6h9oeHI/HfTP8OM9uChGfCalIB0OFcmCMo82rGbJE
fHA/EidX8fyyW1kH0ZaSTVrkY4aC7HPfQe2ncO+3i6X2/xvYQQAxIaEaELshnlJA
Vs59VCFO62jcGPzCPsATcxJhbFF+/twYBsP0ZypRwYVxtaoIiClOErwk3U1mvdaD
GIypnZ+GAP+cJAI9snaylCVs5coER7X7cg3RUXYBGl3Ywj6TfqBD3vvRd8PjVyb/
e+YW1OfsGiAMMozkRcnuA9ik7Q/aRzMFu80c4RAymGEnSSAql9OnDuawsTfOq3ZU
oK/PXL9V6MTirozlh5lDyWyeGZ5Sxd3pWLhKU+5RZLXqXgjpgESRXPvIeyZ8zlTJ
idcs2c/tTBslrizLi7visHBj1pZrwMx075xQsvWs7ltiFk/H9SheEnlNTLkDqD7J
eAM+qJgwB0ojOJcdAr/Eumgz+80zY/gRPKdTuYFz37tucLXG75Nnik6bbyWpdOGR
H6e1BK/s12hx6a8l8jYJPrMK2U5o4mdh6xXndDrAfGBjogWdoDqe/VNDGVZMnwQx
alVByXhwfuap/ZBJ0BSth8wNY0RebJFl3Gti1HDJRLOq3I3Nb+g7PwtHVaa2N5Fp
b4e08cDScO5gxccidG4V4gMNcy0tV3njkK529lRk3aYnM6bYbqqsNakmB2QI7AKc
g13eFQO5FqB3spr0SakCWFKRY5UCAoYUW89sxNdirDxmdwuqi7SzQL1fsTpOAIBe
HVtLE0655YVNJg4vI71SdThByCW0aP9oePkt1hethF7I22cCjYsOrq5b6doJYXQB
cBDOBzcGu1UatXdqKPsCjX+dAowKXAG7nqaZs9oXp1/xMBDb3ElkF0sRtzzPznCl
+HPrn8SQq8VsQAACfly7m0XKsLBtAHJhzaR1liMto7IFzE0sb0zwNT/sWsSxYleB
/Qk1XadLKYa0l/PzhJMd3IbHbJHw/pCfnBS7S+0d/et3/jKq3K5+NrJqb1oWC37p
bqr/jfuGhcEQuAmUFAT5RlUpagBTnSfHONGq53hroQLcijpwkdGyvXG/csIfiaO/
FDRl2QIelF/t5I7Mi2rvHPyDRaTYLsGPBcVeyZOeYekSnAEYFDPtegqplux9r6d5
5C5fesr6GU0+7SxCvV01k05FlCd3V0vWtTE8LX/RhN0Y5U5z71vNcy0e1VcBGyTA
OUQ53OXND1seAE1y6o/cjHy8f1m3vrE8/q8S0LO7NNEZ6OlqapSngnDydbZeW1Kr
qP0iKxU1a7/CDmuhVRe8Ctl90AoMBqLmuPHaM4QHTNu/jBPMZi2WzoezVvp+qyWg
/HsJokQ/zxfitMz+6qiK8g+qvsac7KRweCsgyv5QWNrkMTZ3YPeFnzkHEZQrizpF
IdYHfXNArVLa5LES8l2+1UYERCRpc2ND+xwFKSt5uDf8I4hElqFIBIJkYZzBHu6r
KMHCJhVul0MZpwzvC7Gfk68YThnMCB0cAyJkvRwzE8xFSubdVIOmqtIOR6fcz76L
5U4k6khTBtE5sSNoH5BvFvfje6QMzEwDlkiEJOECqDQUXDQsF0nMR+wTbK3tUEnD
S7U19FfOz0+TjyvUbU7muIO1Gdui+nYqbakyJ9VH1BgGVZ0XNW9OgpLJ7LsudSI7
G/wvjue7X1RGgnCi6NNOFtACBXP8IJ7xvo0Szrh2JPYHltPe93B7MHGxMxdV5pEv
Nd/th05AN3HMzak8t1g+34l1qatGJALibqhkG8hnTTGRsWw8KOZnAOOzYCkAZB+h
Kq8/vmQYj/3QyzFC8Xdop6EVfDYcDblB4t3/apBsAvK2MpIAla+ObRkX8bI1fdrB
A9u82CtDUyBeezCMp0dbbKkZo1qtox4+eGrHrgCQ0b2XGzRE3mnHwYOKcSaYF7sO
EYbiKXOaVp/YWcRPgR85dAKrt4Y1neEiXYigfpmom4sC5JN0FjwCpj4qlZ8i1O4l
zxWjDRskd2g6V0xINou/qdeKxwyX0dM3/3zAw1kjcslt57EPOMEKkWI2umDJ6yY7
sR7x/jBOuGeee0RoDedzFA6QwQJMtaKR9unzRk7rekByGv8HdIfn5ckkoWoTmwAb
i8tWe6S1pPhiQ8pbWhPbnm8qnVmLNndsrjT1A+jmPaqAW3oGnJFxnGtZt/0536LQ
S1ifwFAMBeXgjqD9Q8kvzW9RQVpgDZR5tQ7iL7dXFl5eM7rE4dDYkYP4TjsphNoL
o5+dVADU/bwWB/pR0+Xgbx+X1g94NnlLxH3O3ZSellzCtB9r2J8MP9QxI1Is1b62
x4gw1O84Psj+zsHP82+jFLB5Ppe2zZYC0jgak0BajRqQ03MJ/aEA2IPgV+i67r9N
Kw3Zfr4+HpY5BNt8hSH21RWdH4hxOzRYc+QLfcbsCC+8c088aJIHUCUOQ5j/QsAw
cOyYS0w2IRv/AoTWROQBnR7Rs/1hKnCA7I0xnYDxseJj7V4BQRFl1MjkIsTFd7rJ
XRwEMAZqtd/tt4bI+lRTxbhG9NgsrBxyp46Y+P5uN4J/zLeP4jI50RtbBVyFlqjc
W2cyMcC+0dgLETEzey+3UdyJpQZp5jBH1CUbKVj+/YR7+qht80Z0WrvX7NgrNdlu
Ro8fgEaSMSBQEgFO/kY/R53UTeXTef/076Cg5MCEkb1Fyh6F9KzHqC14TPVt0t/J
xDSPKvG0aU2EpHjEwaSU0h9b1Fzfkmejduh9PTWAm5wPZ/xIZGqywt33JFXDKee4
1Xaw28Fzq7/08TzganaQDWuos6RRNPtLtwTGMvR2c39fqZ2BsNmAyaNir3NAFWc3
C/cv+y3TAwQCiko4JRxFbNECaeOkoD+9cgGaz5Zoojc8Bp97cL4le29PgMzXTrXD
8BSL6F3QqSl94zxuvjsajtU3l5psLSsIx9Xh5th0W15pCofMFKaKDnyzst9Cq/tH
l/qktxu4mgy13gn2Iw32hUeBhp8wPKGuiX0kOZSgpduKJYpNBhHuIdZchyeKE4q3
Bs3kGrUot1AbW4jsA4h0+6ZroyOwy9cLJw/xfSi80RzFDB93H2MJVFZLgqgvTDUP
XbWw8bZqxqwySXvsJFkMRMPa9J/2P+9xnR8NDaZQwI5KqS57/061jBfSAt4P6uGR
JZoBX6fFAId/D6rMfhuyHF/+vqMS+ToiYq1yW+Vmva6gyYM36lhCSIxsjcXHK6yF
yIzTY7lCQYBSz5ctHXkYCGztFZqI2HKnpjmzDkJ/wFD85sos+pUOeBTZoP6f9ws9
j6foYG6GMVpcbo5gNIgmcRKuV7DjOG4zhnuqTdLdIHeZBPSpMYKH2yXstaOzInWN
nXzM7zk1OfRdx05UKRW5ScQGtBUQ4VgGotY8lR/p9XLHQScNyRlKJ9+bqoqQcKdU
ybDil/PixsjAB0vXJwHLxZ4kfS4EuuxngSBIANK3Al+BrwLxaSEkodlVlgPwEIE0
mSdQDYefMIQcPJBH8FVmWKeXL15hOeDF7WVWsv+aBmhfRJcZD5pLvmq9AcHJhEMv
DWSiSYJ1i9wS2SOOP3fBPtjnWYi2h+vX4cx5oieUWxz2Yr4++hZTvZz0OksBe+qu
aI8ZZYzGVQfrKW9hdLGUqm+lWW/4DT56akjWB3DNMKGipGRJ3KEa41vfxcQvL3RW
z074J4e86oV26//oTt7c+cZdSTG/PtLzLhGB8RUfbTiQkdV/NsGzqcJxDQeAigyj
MTAKGUn/jHJrYGcYAdy0yqvpKgKbbwed+bJ3wev16xbxd0YfGc9LFJtILzy0iCmL
xxePA7uCziVNkSTZxOUD/8i7ls89NsGfC3VcejWIRkMII5IciAKa9q3CK8iacgV5
cXwQAjGUuwxb8Vv05qd0Kezx6D6mnBQPAJ0TJVhBhBHeTdbK7RT67fjjcub+Os8h
66ECy4R5Ykr6xm1w35gnLuHJglGVz1ocLtMQVGystpBJdIZECR0zXb1EZa4bW3TN
Dau4UOCRCa8cN12iPNLf/aiajugyGuGnhPCH5Sd5VMYk3kke3Lh/HvcLJS2bJ9L+
vk/IzuLRyLcqLTqk1/vspbYYO8fFiibQ1nO3cSSDgyXyKQcV9V7OwqJvi+PuOFDT
1zE7EfZHtb66tBNtry/Ju13hobuVCZuDbQRg/mkIbXDygU2fm8rYhLrz9Ei6dx0i
xMaLhXWjbAKwHp0hSI5Dz1kp73c5PkoPZQwvFXf73lwoRrsS+fvR/VCKumNvljQ8
69h9t6BpUPrUnXZnAPI2z2p/U9UByd038Ha9krhEFJ2PqID1bCFc7i5N+SdTlhMU
qZcfH/kjitUXTdLDRMDF9paPXGK2j5wCzdSqTUntb71hnXHRiOwg0cU6YH30ALyZ
eRSJq3hjWfA/ANL6sHPxJyscRJOSWcn4YqSsdIiFcjr+LvUoChq74rzZxSte1pMD
HcNz3waz/VJskxsezI19ZUIpU11Cfz9EnG/fy42B+7r+2vQDdPxQJVY5GP62471n
SXz1HKHndAapbriMRsb6K3piR4FWGI+iCO13vt91RdHm05w2fiRxaBujWVipPuVD
iR3Md3MiuQIlqfQAL6eLCq/qKXfdNrA1cX5LfBplvQ+tcwYp8a4IHh24HoWjBuDu
eNenD1IhpbljukZ9cowgeTawy5UZ40Wt8fTSmtUR4+B7zQFTgRPztw2zzNcZpMg5
AS9iaW2X72MT7kazzbqrlIXr5cJEEkqL1aw+bAjiXJvG8Dl71xcBZITrJmdAN6tz
QP9WL2AlM+rlNSmAECZPCowZ0xoHFDJT2GOJvrr37FJlHxAD0MhNFal0+blWXH//
KRWBXRMybdswauClKbTeuLEJAVrox7IW5Oo4sMh9MjSNlzyGBWi3hpeNdoFMhQ/g
prbi3bVi4jk+mg9YLFLXgEFUv5Iz+9oL1O4oBfOUPQnMVq1B6fag4Lbr5L2FxsaQ
kIo6ffpuN2sfeLv8P+ZKXlYQwaDB8XLaAsn5u4D3LtsdZDvJng0MEZwKvq7IWehS
ll8m0D/ZhnyEOKZjrizBCpsC2vHshs0et7g3I0KYKCWyhGCF4iOFgOzpy8JIWBQI
VPmscrnVb2dIyVh7GcD/fVWain7nyPVptPeUFtWGiiY0RQhWC10I0wWnHBsEDgYW
OLQj83jSx3Zcf9xx2DVAwyOtVvtz/ZpMaEjidpuWR8/vl149PTmLFlttymINhaBy
F93XNJN35wI0Tj7vD9M+ruN9bl+0NAZbdwMGzNoZUPrGtljLPS0Gg0ajKaP/VnTH
sT78D5fu57S/RLPu0uxfyg9kRXbDh9WGCE3f8icmjyO/rdZ8NmwrjvuPhea3jJys
3YAh3NRkgOYlpaFysKoM1qOFy7IbVQP38DhQhMh3U5Z1dftyC7/mj0A9JYQLK8FO
QpFMh3W3T3oUwd85HfcnHA291LFfizjgIpaE2Z/Kd3u2ebEyloKhZWl6WHPc/xr9
Gw/zc/nQSTckimXGsxqnIGYHMnkka/EJ9UKLPdfQVJK7E5F8UgA79SaiwPJLuytV
LZahSXgIQclYt4Xi3aYSlpbbnF46pJuE7l0+L1heKB6WFavExaWwhD1KSZXRJfFw
SYpuNvUWNLyeT8XnzgNd3+B4ReenALng7t9cMLAyuYZsH3lqCXEejsAUFKGJjvWb
QWVap+8U4QzQRubVy15/KInrsWrVvpW1vxeBR8ypWugzBWcJwBuv7u7LnJC65Fb1
MPLvjmCaAF/72QFbbxg/Q9V5794Ka3s/TmNg268rw3Lo23je0gqC5B6bIHCoqQz+
g77NMl3BxosPSTSHMuyEi0/iQKWlXqlc76V/HZhOjOsNl+r7mbzrSYJTlEExGQzZ
xUQalqVLuoP1U1Aqj6Y5EckaRm3h3Fs/8wPcu7Ok+mN+okoI5dTwUlutA0lGDSHU
nvR4GcHfWcb0gJEcldRP3717yEw+kVF18R6XfZ2v5+eCMl6ndpil9mzLQKxLRGZQ
NkDdxX0eXvT1p3CtXLTkg/7x5bwGcqEb+sYtlEW8VOBEapuLcAkZf/JMb69lxSDS
Hh+3u4Rg1o73XEjkx5wXtsbnMyUhg8yY06cHcwwhgFU9GfDw/gGOp1yBLYzGfyqm
4V3lKh35KEkm7FaTgD+zDCSF3QSUEk9X7q+yVuJ2sjrQNYiutAVeOC5eqNV2cILI
Z8oKuNxwYD/ZtY+WWbRl7abobnOvUsyTZMN3FKwoMP1WjnLdy/dsW5/dAL6UFik9
m+rkcYrd+BfrdYIuJSCVWI4nitHC+TBynQo/njDAFCAJgK8L9y6iLGhyF6uYTrvI
5ubxmEYQP5P+VXr2P3UMrRHKmUR1bXYfWZDoe5TBGDrIDtthgu/mnT74236Mnjeu
9MISUaTjVzvAJLYBYHL9kFb7DQHEVHxpZw7AYH7t8Yp6cONmeOEKGFoeJTF5zHns
hjPTOX0P5s3K3/uQNIMmwwReM4lir6BNMx6fi4y3FZeqRb/xylNjklrSD2+g8XLZ
okoL7GJSmBFHKF1zETAYu9h3h3llhqSDHBMkOgtmhjw7ADfXYaMov3yFuMhJQ4if
JAaXNMEN1J8x/PKwuetKu3UI7eUmXckepQs7imi76z1e50s0ZYDaqqys5qOuE7kR
XyCMWkF0we59cy/7LcmP5Ek+5Z2PUG7H1fnzZZjsYeC0Ch1k0wcTTk5HU32Ws0g7
jN00FnDa6zODHnKqX80LvZR6VNmblxZBRt13gzmgp9mjB6a2xjesS7wYj1K/4VNQ
Bwr0rCPDWaSTnh/vcDf+vLUaoTi0swD5hArbuQ/vz7CCLROWkZlCnZuR+zS5mLAC
bY1zSGPoqYA+yMc3e3ETLHkSFsMpwWxpWai4o8jGzp3jdo3JL4xzO0GfswNoTNog
LRIbjCbdyvF03vfcAiiWEIO2RCwaRP7y+teVos35w4YG3BT74KE/mQYfXtrvMAX6
ZVc5UGQpIQRUzuwA6JxRXShTACW51pyzldFFfehfmd7ag1SJsN4fbf4VVQ80Sp9q
M18aaVLxqDl0lTNfRHDOrMKFg7RpCeQLCV89Z3f4wZrs4xzi+Hz71l5nzCz0vksN
68XCSGG1lTmenuxGU8jCayjvRPu6oKuedpZd8EXDnwi8dsNHEb6sLlD1d2HJ7D0k
+JzsT7lbPxTpsNaH8ySOK8X9QiKmVqYqjkpiFk4r72SMR8WZMbFWfujjKbZvdFyA
YNTkGyEBMaa0J6fKeOF4n7spfsWx5VNIONwRgT2JZcwKpaCKnZKj5ZCs4k3CAomL
ieUivi+cA0iIeMLTSmUNSUtz5nVlNXXMdMHdHUyTX2sSYTUmsp6YWAVOjiPgAPIU
KpRukgOpITOlbVolSSMmuLYTBux30GHtagl9+cuNUq/eEz6N9TEeWOGYbInmcwtZ
LZ0JPlNcONPWpIvAFtwDrqUZd2rQ9JEY9HZpi0AfjNyYVmo4uzKL5+4kbGTkiOGF
77mDpmXfe+3Gs+p084Eb5PJ27c6Mkqgb0XvXu9y57027CGzOr+6To7OijMyChqe+
8jIicP0vS3Upc5Pcpxu4QreKAKTfAv+j6L7TxrSEz+EMQ2KsfL43qzW/+8BC5tMb
Yo2AfSG3Awze+vdqk2vBuIDWPAWZiMjJ9mNsQ2Mg0v0Hq6g8sY+gpWvdWootjrh5
VW8ME74UUC8hN3zw6sYUlXQ2pSxPYfbLHGObTgkn5+SG+R+vso5lQMdD5nhClt/q
Jbg/GQptfW6GyZFeVHFArbzF5uL4pwN8OXJe5x0Rg2dVTy+MPoJeKZEP+aJc05xE
DPVVg9nG646aosUOrQBxtZD7KiPH3c+ktTCx9GafcS895+oH7yd0F1piuA91XHuu
dIW+KYAPAmscLB+fJ0NXAwsEkthLWg8tO3tsbCeqJB9VwkxTjP4ZfRW6ntdr6hqe
n7aoLetfmBdOOBhej3vC8cEWHzR1FuaVgTEntYLgO1krKXCuI1HLZt2USMpWX14D
8YA0xUsIGFFCbuQKifL10wAyut/pveU1A/IUChmIScwY1KZ0gZ3t+5SGnJtUCpnF
GY7ZmktRp+hXJGcg6yIWA4n4zq77lMXFKnkrzTWMIQdh+YRpiattGjUJICqrD504
LkU/opp2vFI54+8LAIarL7547RLZVdAaGIXUQhV9vdNj5fgAKCzjXYdUwciZcDqD
55r3N0uQStWmPSt8vSdD/bBzSSVzYZP+KqX1ZjdXtePAbsRkNGHqoEL4Z0xc5e2l
9Teef6/DhZUkatxpFqLR6c2iV1PU+jFJIry+peW/NA2/f4/+EGMPfsTQZvXMjA6o
rxxurCaiD38vLAWfJqoV1xIgpSB8wsOeNzzfNbMGX0XWeM59NgnUWevbn/BbgkhS
FezC54z3uGxmimrv6J6RvAYczjYfq/Ir0l8t/2dIjp6dxHwJy8+aeXaW0dx+0vFd
1al/sHEMwmfveJy0hWk5goiZ+YckBx4dGjX7zOmEPiWKHnjKriarSpCeLXvIJzBU
cQUHD1mOyIHM3zSJlMxtljtLBXA+wUx6V43TtFgs2QAlT42XKZOrQleIJw86JOiw
LZHdtuw8Y/Un8cUOFmZvHM93IGLvXclUQXbiLhJVxaIjiJtPfp5BAT4bKs6v83RE
XMPf8W/OIi115yKEC+mCvgTiSwiMQCmHHf+ME2rdighNMRrOSwJWUX6AP7K6GqC2
O8uon+Gg/30FsUB7E+grvOfBrvcmVZyH2zW4+qZ9i13I/l2fDcH/eb+jQPV05eEl
vk5iIq5874fH6FINM5QqCrRGclyQWjLRVziwBKgbdEtga+6Eab3K/dpnucAJYN9z
SZdW+0WUlzW23keTnyt3OgjzPIXqZ42AhuaQ7iwBmUdSGT+JK6r4igIvN1Yp5LyC
OrVCMEW1eyO31i4gqTSLOO4zm/s9uAjHVFInCitsnmjjYBS+J+7syeTvCH6L9jxs
+G1mthbAXrUBvTk032bUzYJXOAhn9EBYpl855z3maUAkPju1sB1qWPXw9yJUmnGg
xxrQD00W+1EYk8bfp0MU4vlbDPvzZq7eir+lAKbF7uHKQwrgo+bVwQiEjlLwTCxE
EQ86o0si/XGQq1bWRlUgyvhZabzsVK6tCSCyCD97ZCKw9Bqbqjm3mNYniFdHuhKF
LVgr/VnTKKl/PjgDuNUvhnhscLMSscczCtxBaGBHE86CN2ebp/auid6NdyuFMgoa
a7SvOBqTUPmYKWQFNkpONkSXlMEmQdJt8Lri7VywO+vTpRvDOI0XraGex/lHzbDF
yN29OElxIcdYBpe7QesFkcUhiOzZa1pXrocSnPFnbxm51OV8bx9+RIrrkgkZ1+40
De79FDlOnadbXAq8Li8bC8t5ToQ5qOfOQtqO43QWaFE+rHXgvqtRU34igdHHqzXL
1E3mdSeEBJiY4IGJdur8Du29nlyLbAo56xDMOV6rN0gYeUWSvl75nWviGevo2N9K
o/tnP8X1T07ADtgYrwNLtFGCxx7cPVZsgWKD36fSPIw0m6qqsfrvsRM+IWwyFM4c
fZNX9p57WMk1TzkO9eOclgD3TK8XyLYMlN4slCYm1p6kGF+oa9W/+YS7DAr6n8zY
Py2vCykqkZ3yUK7ipzMHt5x97B5EJxLElM3sHhbVQ11l4YUt1xgxFW0vIJ7QRkBA
4C3XUkCnUsC+vIGzLGCBit76w2s3OWjWtpo6Cx6INiG3SlpLh8T8aRVtARlqMROt
ZX8ovRrpaXOxVmjW7tLQz+NZUY9WFqQPBN+cvROLnI8uVKLdUMondlM3kXH1myde
XBCeyMAbDd9s1RWGnuwy40XAeEPYD1N3uwnwKuSRTfSlc5jFjPSSIcCwfYFWfqBx
KYp4ZrqxV0k2/6E/n0kwr1njglJynsvNpbHKFHN1X9k1tcEFs3fmbztKBi13zH8+
6bEtpU9ii2iNnprjOVqPSlrbJY6Me1XxD8kJEVT2kybZnXpi7t71JTwRX6L6+22m
sKmcNLvpgEmx0Or2H9M6r18ZtbGKoYtIMVIPrrxRcYl54Af2uZ8m80JHTGFmP2tZ
QlYRWs4s5XKQIyrt10t6QkGPq5yfMO4gNj4wU9ptEcKpUoVF8C6n5JSHGSlWKAdJ
SA3uvlBRi4DmJjqqK/EHTAdyQ/hLu2IgikxABiRO+p+O1+H/F/nWZMqmBEhDgUol
M4WW4/PZFSbHZ7F6iC6j2lxh88kEZrbn5NTidxfZV2b+s+6LJhkyrmJQBMc8eSD7
RZqk4rUt8BUIUJ1mHlDMHw7AjKxksLzvda41DKDdEC7l4FdzsZGpNQN5qZ7nVhoy
HXxcUSu4QtPQCgfgkCC88+cYvGH/NYjsYJ4yqpo37NVdhpvqWxYP9BipxU4bn4y3
7mIayx4Bh7rmQrUlLgTuTIcY/0ToH3JU1d7CUx0PnPHGWMVxAOHonsJs+VSHoDSs
M+ez99z/jJWhFISN1Y7IL8ZADZGDMjC53xPBB501dgasmKBtd0b6uZNlmrxs2PU/
hKztR36CXGL75zbz4DDq49vwUxGh+19W2dogMSlsrHRhTBCV/z51/2EPIgYJx9VL
azD97VyFHIIimeFrFhqKmT0JIbG9EhafhvzfLX7hqiJE7/VkppPVDmRGyE+Ivyw5
ZXFAGdq7uOYZydSQ3ryOwPhEThPxAistCxOEguzR4xkDir0Tj2s4drDtVYgx2dEv
4q93Firp9iiWX4j4H6TPZtc6opL0GqOrLmAm0DSm2OdDkxdFglb/ZaDRFJJz6mvX
4U6iGwwRXUYQDSYLWrDeCuDSBmct+qMcjg8OTyeKMu27JT6WA12IBDI9+2g3MHjx
NFN6Iz82qTDkqAHxqKoxMdKz5FrY4IZ7XI0XJKCdGpbD4vzHekjBbYbC/q+ym8WW
xj8TTm5gIzk4looNLQ8Enagyb8l/OnBgwQ9jrOwJC4qvuQ/SJ8opGBa2ZqNDHPKY
6ekqPnQMWQkxMkVlrJoTgwJcaIPAdyN+SZ9BupPMrxtNdXmPxoYjyxcT/irdyxK/
deNS58sDtLd46wOJleht/1THmOApECYULSNXLi/REox3IMZz7COdeWSlX7Ny1CoI
1ks1w9yW6XEOP5AeCxP31B0bFSDqp0Kt1yHd0U66f+4rS5zk3Dvr2ah0OXCWSYE4
LBipra0ifQ/2uuo+OkbFlHGMAi3qU8zd8ypBxnbzABMJ1ksqGWG2GCTA/oeX22Y3
HydS7AW1vmjqHj5s/Eg4s6l2ox+gE8IJN5pFykTyrvrBK0KrS1ct399WmHmo8ktI
McvBqZ++ImA5iEJbq/Qiz1POARggQJKVaAUu/GDcwmJQeBTP/uOS+lGEq3OlHsO3
6E20xCpi6nS5NjHFnmA5wj/IwVtcMboPdjq8DfF0ZIDkrVorrU85K7JopLyv9Gpr
eMsC/SdRBeq97/rjYXTFgZwC7A0TTUvuKwEYnoT9z85Qt1qz+FcC4B1Tm/5/Tnzs
c+5d774hHQVA7Cmh3TiJ7A9wLGDU3Cxxx99XbGGx5JcqBxn8BDK2C/QdGHaNIQpM
cyOobTz7AQTJGjhj8O4RlsFLfLmmDd8YO/2FLIRUs+j98sZgu6ivGBhyjNY+qMpL
AU+C7ALdSnETRTi1gatcdkPhCUeyVN9tMXNCS1QACQeMPnv/BYh3LBl1Ui5/oxM6
nnsahnIYof8a8WRbRa+3hAGdONusahJ4wlHMVIUHjERzqQ1pdoRb+X4KWKEAoM1O
LYANpS5yzWWXGK0UzO4lrY7WCFxejeAM7B0SKpsGEcD8gw/V3Fp7gS+zgzlKbIBp
6fTsqirhyEMRjvdjdMhrAnyTkgWSf0nZ4FJDGTyFdloCnbdnFYjHexZNctOBvlYl
JpNv6ArHlDUE0ZvH1Y1xAi1AwGqQptnuh+E7/KREr02xp4CFW+d6uoH9AzOWziDF
S9gPQXlYVKZsHB0glfpnkYo9HqwMNNRoK95LLQAVAKgI6v3kfiFKI7RzuXxDY9Y4
aqySafpzxXKLJePsB6uulz4c4OdqG9WojDexk2b6vgX6gw425W8nBvLUghvfZXLx
TI9sqMgX3Grefzc8uWLRSHOOc5tv85ddZl53NbJgBzpqzjAA2b3goBADeH+vB9Qu
S1Fi9sBOJatHlkyAEP29ZV2yPB8mFbd0TNIrwy2IL6TVWfQdixYOj4uZTVkZKe+x
xEes33J0BTljkFCYzaMvkC9shgIZlQUOyrSEpePuI5s55p1QHH37o1/lelUKNDhB
Z56j9F5xXrNCdR155fQjl2QcVg8IBW6Ld2bjP+7hR0IigSpA5/O9gf1gntLTihtj
6qPh5WjrQuM2ImksGotno/fT/iillCPMWpRvGJ3FKjpiwsYVDRq4goHDvd6YQCO9
Q1wx77oDmOjdJ1IkTyAy4ReUK3JxWnHeeqvRLbykoMTtJrRLpk4K4VNU/K901MMH
V1uvGiDLUjVg2yHX1+dSXOEfSN9UdcULKffd2MWOQNDNWtXNfrBFrzolwOTA6ctq
Sn/YCB9HZBr/Nwj5KeB+swSmxVnXGQulvrqFKB5igYIsDIShX4koxEfwJbh2Hpwd
MaYVa6Ipx/pAS+R7yX43eL5QkI6OPaZjnLVAsLaB7RY250AOQLuBRaKF7zgXHxMs
bs2th4Dx2dbX4AU/e6QJ7Xgows2apEXbkckzaKegLO727Rp3Gt9c60xkO8eI4rr0
gTJ0pOhAuaRvjP/MRNxQIAxg4GdQiK4AbCjFj9tmODOrxg3iUV8RAg+ABAg3XviQ
JFe8rvO5UpxaxgP4KbJBcLMaUlyQS6O/Yl+mUb9H9dtODspprpak4GztoUnIJupk
5cU5kQJAuu5DfIxBjxQ/ylzju1GorjYoiMWvK2YchtX5ICG6e737CQu9yp7yEVZv
/BtPJjNnOu8EYbX7pQXVW0tAbD2U+rs4ERq836xS12QXS3KM43RteJnlxC0aTBSe
En6aeKkb050A3Rlb3J6an83xiYo2NnPjdA4NV5mzdVAiin2PTQ+yD4PeY8KFfLfL
3hQX3AOCKuQBvMXSlsOuLai0EVrVnvkKjPIK7O8vdL260+VY6Vf5hPM6J+TTvnH2
vHNTBK/Yd4J7tqGUNXiG7FIRsfqkb7KNw74bYKq3Yv7/f6xiDciZ6R9vk++/2e6l
BqkYxhaf1fXZ+mb+xa1LBQicuROWS5EWEVC31ptluBZqtxc/cuNuXaHwf5WG6pZL
qFov2mErRcSAl9ffwhmyH0VzhJ1PsTpI9k6D3L974MvRggbMPF606eTNylEDEeIR
FM6en5JK/hnGoNR322imCcpHU9sD32if4EnvMOvkN5gPyw7r8b4FpLyxKzTDAw4E
gm30FnzC4IV/1vxaq78cfr53j9VsdIVG5Fb4tnjcseGRtMruLAJsffJ8+SYzOxdU
dXkAW5JT5b+g5IVPK1oZyJb0MhX4Ca+PPa7uc59E7lq2IvXHhrNt5RpXkBiZZiVL
mlKWy43rP8lDBMBnw5jVytIQO8HZg2wrrlrltWQEaR41A69NT1scaZmjRgv5iERm
vhpMhKRheVpgGbvU/TfA9PmvqBN808/xLIWb6LvTeDT2kKJfT08WcJ4eBl6bWWAv
CvWNI9FwO71vzjER5n9jGV4EYCqZ+NIl4yL6k/qYSQ9W5lZ32R5Prb78E9Ac/uJY
7wRAHMi3WHgoaZfmPi4CAov8aZe7zD3eJarlUokg1xAi1+hFjuvf8sEeNTzS+8rP
cnGpBMOaAVPpfxBHrSDNJkj9dkHUhrXJOnXd1TShyyV23ZDwxDA0in0oS346s5DY
lMqUVMrBKLbKQZiNJSwmnFvJzv1IQVyuAyF/9bseL/nY7MrfRmii5cuWAEZ9g9nB
uT18PBvxu2v0Djko1zXQcbQu8bDYHyFvKR7Xg1+eAFNwUCU4BcDdZern8n1AD7ru
libiCamelZa4emErfdPu8cvGCDYnVYZz9Rdhj4us8Y90xeEUe4s0sZ59bKDFULP5
hV69of78AN8v1ZcAMHwEHS/+D1j0WoFUe4NPCYGjmCkd/AUz8fySpHGFV+Jo1vB9
XpTDtxp8N1hfrY9nDRF4xnibKp/jxbFzn7cYr4tYZFeSME7sEUrQlhIZg6uqBDTq
8FIPCwYkXdh1rqTG81VKOLubvjidfst9McvQiPRaca5Q1WR6K63k5m9NO0ZjPOuH
w5NgxmpGOciOvB1+e+w25ZjMFol0Znyw+9pLGYk944e82PErEQ6stE/2pJSPIUCJ
JhC/cEqMg7e45uBVXOmXAD0quMkbwXmphMobSB2TxYpAdtebvysuEihnvK5F1n+S
CEPbRIyVhVrjvPdBEVoWUxmTBYXZtCxzFJyxsqh4pRlKbs+9qxSGWXdEaDyAipvX
MttlhYsWdLMwN8ocGNvoFSlKAOtDnUVXh8fE2aFTdOC9q/JqQ4kkUvU5dWKsINRK
bziBidhqj8ERWk2SaGisYGYXM3CjCPtD2dxYv3W15lc4QPrVZCUZl1+uJs5WMCTZ
D6amD2mpj9DxpyaHBnhk75gUjjZErg+cWbop88SdF/HVprYF6yjf1NniPfp6DsFB
IGBO+DphM5YJYCAHD9VUsVTSHUWCyHtRzxgzHSwrZ4Lhnx5gqSdzqcJ1lyE1EEYM
gwURs4gvTaklOG7VTE25xNO0jSZSlwtecRXQSnr7ivSI2jio9x89dvrKB3gsOnsp
qyk8UzjR6/9UefSi9ZNIoKO5ipIPGh0FhkPtxxGtw/+5pFHExF81hPaDEXuOHu09
6+kiCuW9zJZo4Ibl08+9Bho5SQDZDJW71TQy8ksDDK5F+umQSMRgHI+RxNb2LhWR
BHMMwnxVrPEx+F2bjJALTBXZ3U+FLHwQQm2Ky9Zq3l4J51gWY85M/SrWfgk0a/R0
9sPf1tpaW3a5SjctWJ+RNh3PoNhZaENRYpQWq9fxpQwGggHXtvPa+Dbx7ULTAuu0
xs2owBKk4F/Dg/7Hf60oqKZIGR8O27Y8dhxgmElvo6IZ5mNQcCEtI2v6os/lOPWT
1akrWreX1UWuJbxv8YJ2zHO+R6k+EN7d/uTEtVjIRAvQC5AVfPJW3lJ5T1ep4E6y
9kuUwVOAfaLkPrCTJRlSBmx1j3HC5qSv5SrakvPP1ngQQjqHDEe2J9NB7tohUL+z
T4ASkttHFsZC+apoU+AKvKO9I9JC7Z6pr6zd06T8h0wZLDN8+Wosl3P8q5ENCJfq
jy00GQfLnYXdOPIP7iec5E3hyAtPqR79EETEwUmPefpouOOrKSKp996LVsTu9pL2
fhq0AYESp9rdaogr9OIsGX3/+mcr815CkmO5CbO+EoXZuyOmXX4kyf08jh6E6nhD
sl6XIivpQWolgBsS7DTBsTj3eyPVDQVs1YcINxzfXUwUNi4YXL3tkPehsZC0cOoe
hbiceqF6BE76IcOG2TtmpCmhKwi5O8/s0sbE0IeRG/5oarlxL5zUtlMQDHcpkOlp
V2iAiW5SnDmADoZzuCGF6fKJ5uVXrqSNoOHz2fugIHbSBjDei8WH6wFoKLRYrwKd
2u9v1ng4E6YJh3PtSrnyZhpvXaMMzTA8+jSniiD5dIpBgAfy5E1/X7CwPK+Eb1CB
rXzXEQ0Jstn3LeBLb5QKbBpatF49Ap1yT6fFJ/2AyPF9U0yPesuUujimx6TT0TFD
ZHKdTeOfpBHFVGLUXMRiw7Fasw8DlwXShQYBYOSmA6ny9380e2A6gJu8ls39mBbD
nklcAd7bRfUZwBUIaTuSTf2UosP8593GKxzbB67TwmQmxHzfHm3hDlREo6aZcwc6
GByAMLeVnCZWToMKvq9bg9bYH4OsxoCG4wm/buw8ThTNihucXQWxdXZhqVQ8/ANE
H9uLP1MF633rIaChtrsIMWKscxltADHCZGq9AlcQGf7W34hCZf7+FSJnFhqmexQl
XQ+s9Wyx+jO7mFgIMNZqRvCPV4rJ3CFwgCm4rN4BwFQZ/9hy7/HlUw7JNTIDf3es
IX2KppRcDi0CmTJ/Agzo+EE5G8hD33TCbrnT/o2LsAr6QRvaHlgw3L2dXhNI05Cx
06DdvfNzRlooae8v/qYxTCvJBSivRJqnUTLwuYKdwWeCG3YjJXVN92U0bi5r3qzh
l8+K/qcpozkfLv5/V5xH+LXXMVFMhNIkXnwtGxWjdeF0PjMr/71lhEvKa5h7IroE
b7tZwXFRPr2wZINGzZzgHEdKMBTkudgiV6F+wKL0Kj+EXvGVIC/Fd6DzevV8Wpfg
z7YKnT3wuNhTcEAxs+JSMkVXq5/9coTJtQsKBQZk4GwVn1TfjSgUtnrIg/pwkwJo
8tu32QgWe6i6DDHpEi/TG0l8ic7E1dCkaOlkHfh1+d5n9wlkc0qdtRn8wfKCy0id
vQ/OJp9H/HwdXAPNyY/91atgakKrwDjij+WCK0GHg5fyiOMzBA0dCIwkxYQfNyfL
uuteTkg/vJJWZ6qQRXllA8E/iiBrOYk2mSoGbnLyv3mdLC1D+PP2osiIcu5jw38Y
w5rc5KjRbTqnDX5rHpHeemlIS9xUB8lpN+WQ97Hq5RL6x+8vATZu2Vai7Wn7wd5M
3vQesr1nUeHmYXMcXebb0Yh2zTBNe+9kfM63XD5XaV5uvwPU1sj39UKWbCRMFfZZ
ObyYjG8LCNRhSnFvOqgJL247rIE0V/EawQ3zAOIjDXEPExaFhmXpCjDLqh4ldZEI
fmISmlMTjBOWB9IGQolzte97R2aR/B0w+iutHBdgcP9nRndsBZyRCj7XflyNnZ/j
XS2XuYEeNa5+IN2LqyyN1ZAwH4pwfesOFaynA10phc9HdTgbMOOYtH2wpHxx2xo1
IlIMo+62dRxD8ufh99+EUgdllKZuh9Nad7bFrA2HKW9+EKrpjgFobnnypO21W3Ne
2CKvW5iHKa9jeuBUPqzlXbw2l80XL+7vA7UzOnt5kAkHt3dEkpV/Hom0Ak6yuy44
pmUCH9pTqJjXMZnSl9ry+6BloOjsoCkboDbyUU24UACMvqk0J3JkB+Jt1Y9DjRIT
MT7mjoHk0NocMzAIrvuN7BOaupo51TC3/GdqBWL4ua2RrehWxfnioir7Mr2IGSth
aSN24WzJLHVlb3adpou8mVUL3HhYQl2bbtIjT8z2pwSri3yeN8JPwb3uMZa05A54
TYc7UFyh7o08uRMsIuAM+X7c8wy9naRA5EQTiEBt0hcUhhj5KW2VYCPQuvoFSQGC
XNlNs0RJFJuf8Lig/VtcuoscGlGttt1CPsuaixNs7zuQJTuYvjsd31rI/vXWppU4
tb70H1Hmuv+ErZQwbf8OrvolS6ENyRhQuiCAXY0/z8oY1E3RSZMOPKo/kAPk5fYE
xCT+KoDmiqtYqajG3rHs96k5OySHJupAd7tHVmJF1P5n6VuuN3JsMbAkqZWgrilK
RHsanT1j649ywa2sk0CAHnb2hDwAAxzHBWGbdhYrV1rK1RVT2zjvdToRtP/AsUvs
acd9as6EuKuB6H3MarXxL6ce9a/JTTkESU/Alvcgo1wMb2Rc+9oVnbyPcYi3r/PE
A9JSDj2UMwh7CmqI/eC0aJZwzakDXdn1GuZjSiQ98lPP7UlU9OEEm7rzyWPQz/Vg
21E/FRAaJHZBEfeTRgJBO3K/Ztxjr9W+UGm/bp2geUMaEzyO48uLwWNVT5ZtycJn
QV/gwhkU8Sttk85feSz+KdhEYGGFo6deYn0vXclCw6m7o2HBL8otizNIfcthRReZ
aaTY1XOAV7ckr3Gnpen65mzbggbTpetURUa5aarl5+BQGspNGbiHh5an1cMdI5K3
o6DMZLlaw3lb4wbo0xzUBtK3k8kDpBy2QCCvhVg8P4HsIiIKJmriUa8/ata7Hb0g
kPf32CtquRV1Lrc5nZYojSWOU2XIIbb7IdUNeb7APNiPrh20kEWi4g8r1JFB8B7h
oEgFUBbxzdloUkrrSWYRyB/j/bHID6xCta9yjgr6vFJU/5Uwtw6xLHn8bauowJuv
aZn967Mkm1ZWUSnd8gURGsrMtLIeoKik/GFcoH0z6nH/XmJtyfx8RYDRTkZWrzl6
SqxNsWG/w8/1x+fdvDS/ibNryzKVLqNxTmaOy4S3FBvGS8VKD3g7K7ANZwEnlC7h
neEwTW8FUS2QRixqvOPvLrrDuvviix7LEUCSn+4o00rN9GVnH9tu+ed5yiQKhzG8
USf0pAE1EL9jTg3pfJ9VcnJG4HOdvTxBE81QhCPr+7sYm0uoHMzUSjeplqKg4D2u
zgXlW9J12Nd/U/rBTqVocqxQJP+DapLEDT3WUjC3mzfSBfrohDWnw6mhD59+sHAq
cwK3lAAU7GoSdQAAYOerO13Q+80h3rcGcsEj1Fh9wH72yDw/OhHcoyDo1JnynB+h
iuk1gOg1qnWrIoHMmLpv+Aa2fJZ3wgwZsUoOBMMsiZTlJfYqQ2WSZ+kd0IWKM8Ez
8dKgZzTedIZ9PcA7PvHcAtosoeGINfXb7JwDw2w4+Yp6RfJMCt2wl0cH08QygbZc
MxJOr3ah6qgdJ+giqv488TPqYrGkbSm2jePJvmDQZJTa9mztAvcimRLF2k3EL3w4
YzKzKOxp5d08lwQEguo7ZmGQTK1w2z06tRMQTCeFS4Rsctaag/NSddnCiRuZZP4f
C0pT6CE1MCP2mTLrY5fzf3EE/FxD6WFFJSU0HFix+x1rTBK/ztkcraBwtO4ryots
CN9JJV797CxzasP5WrjYoi+H3mSTyDK/+ceE/0T8gfD0WeRZv894Rkg5n9QLvi+P
EsCjsqUTYO6oICAlspd+cOOXMbaqyqfLRXOoocj5OSPqbJtYCdRJe5yNdogfpFHT
DTKKF6lPEV4Au7TnFkJhSNryeAV/rw5kZySfP8Y87P5jNmnnY9J74a4aqoiX3VEQ
WHsE42NTqQVdUqCGQf+VfqS0shGPipM3YLPVCguqpwB3DV6MsYZ9tzeNLh5dPQ+J
Tkmc5Y5H+e/QJxjE3qjuF7G3IF0tKWPO7yFl+muv/ozrrnxgbeeqPBOGXlPAsVzU
sFmSgVA4vJV6a+zsNCFvJhlK/hYQSoJ+Svm6ph53VPyh1fTzRgdsOTVTcIE0m1I4
CVS0oBI2AOTqrZ8dSAR7lq6R42ELG5OHPII+kLdm9bUtmiW5oJDJhpau82jBw20o
7lxkKmIdEAM4BPKCV/KuCXJu4/q7clC/lJWfKL4lPfxJu3eAMlUivnKF5rLNyEOx
A0rPU54zhKAaoc4pv9xrtTKotBpfTqcm4RDswlZ2Cm7V9SQ6muRtWtgjykBrPwr+
DCBxTpQ/3XkYfU6fszApo/d/3bO89SPfBwrY2ijH5944GheRQOJ0/UpSFBwBD8qX
vhzpvH9qkE2s4mViwWQyOBX3E3uxthU3/lQ4N3x0S4BHBJbiByOf+673tNgEW8mh
vyI/RPPtg50UW8FAU5WP4hV/hsxl1PFReiSGWcx2TTVqJb3At72WQeBxgkAlReTL
78nZzm7Ih5OiCtRP3GUEmO80jpLKwyDjp7lI+hmtEg2AHFPOMOs/lDSyG306SLR9
6fxde2enLhO+NEHoBANudMvOMbFUdwAK9+ZCm8EJzRuLvPL3kkCyc7Opa389Sx1S
Tj1997Lo9k+Yk9u/uwJRXQ9zyHOC90BdOLP7UhQwRj4MrSZkh2Ftw50+P/ce/RUv
ZRns9fIAApSZe+89+PlxGXUo618lvu6knoHgCn0Upb7GTbeFaihFhVFbahcX+tXV
hk5wzQZR/1sIdJgtiAlepY8k+XW8lrehnlkYKWk7Z7P/UNWW3u/W0KTNT8kJVmbf
LxVICVIUvn551yxkad9uV5605mY5/+QBXiyXl3kPUFm28R1CYXIA/33lksfUDCw3
9QRqSDGcM+orfNt7WPnDSEBruQgBjJ3OKVWWF+z0PcBtgQDleMnU1n34r3uTCiXo
EnI07aRKCNqNGOLbcOwRA7A01tQpLtzBSIAmJsjpale6P3yh+87pf1DtHCBLRo2J
ghyGFL56Zf5cuL3reWhGabWKUoBmzELN2R9kZ9DBVR8Zz1AcLTsvoJfu6SBSp/fK
lWLbdVTvVjnPydtAdP6JhTUh3jMtBRkh+HbIuyqzs3rVvwJoOJFmrJxRPu2BjqNT
xDY/11fn0NO1NIk5NejCLpdljaiKrq+jCsPOkcX3SZDgIqltB/j0heKuwa4iI1c5
qVXLcQ/wDPBds8qzs2tBOVId9MfJOQ3K7zF5kRIpOgV9HJdZa3NN//g1l2CRwv60
bRqJdAZTHDqfBYEl+MZOB9lOIS07goIS6KNydre3gtFMAZrCMfTLjv/rsOHOZl7I
1sRJyfdWb3iRmUW+nZT8/kXZvPk7eatypO8EiIgANj0o/ykGd4P8qFX+hPtfQNtZ
CSyWc3nOJuDtKrOlPrCc9wIuzBUIQdUDWokkeWPhvKpwKZgPW9nNJEezNGX+kuSm
Hy5to+eTgvlqQiXIriFyRdjzNzsvOeueOKDNABG4hx3BQuJdQAjPwS+l//nGaHaE
WAWoTOqnCCkvaii0LHiP4lS5s8QD3tkWk05fNIYoA09OSZMgfosmQ/eFTKLgrjwR
lBZQcHFODn3FopQgVaUMgv/cLDwTCEPOgNeeEoGgfpijHv3cAXh9d7mFfWT31wVw
p73HM4lbR/UbhXaiEbi68zaz0PVBO0jGmkriTyOvUWyEJ6wQWlpBDyd2FIeGe/3a
b5bP/bR0ZInX5hWu7XvGvzVQ7KroPGHtFMofw/s7NF5eBBH4AGEyS3nQOEiHBNcR
XrPql2DiyJBVTKg/QcxyCnYOJJP3km4lUWXlcEoexd5Dc8DPdYBDe/qSy9AMdYw/
lFCZDTW4ak0AHdbfbDxOhcixmWqsoGHHTkLzblU+UOFjhwgJicEwPQyQHflfNRRO
cn2qIlxq7NHzhAOpmcnEkrftO/KBptlRh/nZuJeBJ77IBrXT5Pq7rA4eS7XFKmCM
MUZu7hzRFWk75qh8F3IGSGcY+Xh0/An4hZtG3cUwNSMhl+GUvEzGFlvDdTSZWDm+
tpesXx03tSd7d504DEliDcn/QpZSOW5tUVp16FYlIT+DjqZ0dnutmDh7qaTjgWE2
AcdUuX7PFtLP8cWdlb65Q+K2H/9z8ee5UKgbHrIzhWhTgZhH5+HAgD1NAdcOj9wZ
qN6RhzQp8Rk+ZVQgYcZLjw3iG4pQ80ZtXhoot/2GmB41xf+lhEttERHtSR7onKN5
n8diy+RcprjjXP3UImAhw1YP8bO5G1L8mqC/vDMxRZNEH1BJl6Q150e8IRmQXvXe
woTooy1EUg5LH7nJDMyCQfYE7JV97cu2JubmmZfY0/K7ovkb9+cnJwAFbdUYFx3i
aluKAR3NIGgeu+1NkiQhIijklG+o4Skrd8AO6J+dtFCd3XvCKAQTc3CM9FaPx66r
sBoNjVg9PoY4BgpgjvP0/zfPnkW/Lrb8mL/ne0EMfX83IzrwLzH+tY0DDRBq2lF8
45AkP/wBYLA558UEyWCVSDi2VFnkmWccDdtI6PYYT88v8Fuczj/ZCqFf7g9ePcsq
KLlPxmxQncwj4zGCcF2UxiWz/kt2sK9KAUQiOqbBJfP5HBU2BytU3xGv3vh3ai1f
zZ5pzS7lbM3gZ+T/9yid9pVabWkmcHxxYhTQb9+SZHWl2+2fD8elcfIPyVbao2Q3
WbKJTY7DBU6G/uxl4iya/+FcRfUQGhvX0a/UCqOeto2b4n+qc0DE3VpHS5kaJClu
3LPCrhMEAk2KLyCc9FQCHD73s19pT2JJtVLSNs10wRYbs3FFSG6Plpge9a0Mr0qN
i8kcC1oY3o6GwRh2YQtu4jJJ4MIj14xhuA7VCtN68hlY6mp0v4jhKu1QP7BdQC8l
erXLfFQ4AMfA4H7+ikQXSKJhz7hFFtreH18Z/1bT0lUjds9YCKo1lZoJbsBhs2b8
rfoXRP5R1wb97S9kn0p2w9xylEdW+7hkHfSFQEc1O1BWYV/MlyvtO1QPjSuAaA1f
CsbtrnD7L48YXZSOuMwcZmH5No52R2UkEZ9lBGFX2mIty3SJdQR6roTk33e8ObEd
u27g0GibvvZnJJZ5oHKIpX/w02YgQ9pYtYEbUwSTXnD9Y5fSGdyOd5g4xjz4lwzF
tPo8FVvCPSw/8XCMOpLNorHkZ6WUVUz8f3woGtvQpvwBV6jjf02M9xDuvtuHU+Re
dYdzAYgNHv7EbYIghtIpFZbURMUau+0Gw6U1JqHOLVU+0tlj+IBN5FS6UEPCaaig
k3dkEQ+/LV3fELsQ56YnPylPes8KgCWWn4vdv9XDCYJAE9OP0AbwDJDu3tl0+JLB
PXxZcrtm63ovq9y/akMZmOjCHLLXGgnDGxjrUiBdbJzV9+nCRiimedRNYiR8YXUP
HVnvNBVfEOuSI9eTLjIB0h22HOUTvAGdjcmsZaLta8CP7u62AnZdNEE/CJisy2OX
dIDlVPmjZrDUGJRHgzpm1dLt7jvZV4viuKBJfd5OLfhVZbuVQqAC859lJHRKbfwd
zBE/gn6uwVi/uRl0ytsgOFVMI2+qUfNm76RXSOvvaI9u3WMlBs890B3AQoYCa3mG
7nIkm6if/NNC3IiopTRzUc77upIVk0yDu41jNvCClNFQ0w6Q4QSPzbG85MnOxtTp
WGnWgqIKjgv54uBHtWfXcMJrmTKuT+pOFfLSFjFF6oayp4PQfSTKCPr7JJcV8qAf
3q6xS3AL29GcXYz4MtepOcOTQq8NCFdBtbv0tS2S/NjVrOVql35MINr3aicOKWBZ
0YUxOUZxCiTQU3BgsWZ5e5xVU34mXD/RxvMWeTrrd9DZzyqkSTuPR/T0lQz2JZj9
2PwCY1SYzbEqIK5tPbS7rdyjda/nzDH2NeYH9eJqkX2+0Meyu8beTKbZAyN/Ec/t
BYBUfl+j39OSNZOcPJo7SRPnYmvGsqOKJni0TlT5yaqjcNoQU2pZbKQqKY3EHpOE
R52lh1ti0ul8EjxwsjBRoyudn+F16IVFMm2k/VF4/cyx4g7qfCVjY7cAqtzWcM3d
aZMjlmm+/i+P+7m+OJtRSkag88teLQ5ksb/GYKikw1fvt+AVYUwSNBlubkb2dvdZ
YihYO9b7pAKEm4T85g7lq3Yvg2utFBmZIbOtSvupw7rWOR2R+qfyqjtV2ZRxy9wz
2otMABsR5tniQeVdX1TIojQSNXu7GULuZEzSmww0oCGzR7/CGXRSxFfT7pX0Us0V
ucUQIiKwJjUJ8WY0YDegB8Xr2aMdI0dVarUkxxdDES4+lSeq17LvWummOiA1HVBU
Eg5srQh8R3ldSGfx8eNmnsP07+QQIQV72JkhUPb0yGp2jl1sFD59u/bMdLXbiIYK
xu5xiXGheb+6MgFNL8z5x1kQhFgKyDvXm8Cgixk6rLmwlsUSKfD8jOFsFtviCsm5
TtdAetoWjatw0AL1Bdn61c0GilFoxA0QtD/vDE6nIb8BLg8Q75u2VpGzF6S300VI
rFDsDKT0ERWySgGCOgAVFB9TqJbAmyQRpVvI30Gw9fNITJzJ0LVSmE0jFOq4qYea
rqVM9iehpOywr3e1z9l7hyyRvR7I8YwI0enIkLvAB7Edw+fN8jHW1dB9gPvjPxG3
1RHAKYKe5gjgmNTWF8teLtLgt2fMTCxpkV9iYqLXlDi8NTZ4Jd4C8OUMzt07tpiy
dNNXebx+fqJFeD+ZqlAPn4vgXB6IcJAlsaRx3eXcaQYWTmF4apj2Q6BiLmgoCRJv
mFjRDDp/PlOPB1XcqCGhsoruwhRpvJLODLuuhNoMooL7Esbvm9AUjOsOk0rIN2Az
EA4N7kU/5RR6tB+ZMHSX+Qf/XG6t8/dYP8ZbzpBNBX6KdBcWUHb8Mls3DffPz4nm
ONv0xJGJHiUxDca70LSveqQ3QWQgHX5V9mGUXkBsIEaqsAxiwZk/PCQqZY+1o1A6
eEfbUmgYj5/Ty3S2ypXj0kHuG/OA5J5Vhw23L+hvMVRRwqLSrimIo4eGxsjcd46M
xy2/ZTYiQyOfMxHR1jGxeNvZjk5oRaPTTjhD2XqHgq9vXdXiFR2iu0Uls/WisnhN
FgZS2MHjSPaqbEpRQx6L4bDLfy5FIGhZe1ghOig73W/XbiPsySqUaBIGqMHC+Rw3
2sgEWKHuL3UN99NsPF88cE73LSzSLJyBkUbjQWzipR0QWT/kPk65loS/GPnIBrtp
suyFmA/R1RjzwB18kTHDat/Gh/qFSf4sWLj+/Fz+ZWdHp0fnZe8qgWeVIAd6o8Sb
3KmOGN6v9p3/Ax+luCOq6/S9EceQp1LEfMjucSDyEx4otOm5IRuHrgflEPQkyVHQ
xammkhwsh89Yeazpl4qF6kLp5kvJ9PxD7X9jBq0Gr+1rKkyqqlTdybh69qEPhiH2
GuEtDldhjSasuIMFJlVSXKyXutHrUp1C+J3fnEqZRp8T8x+3zBrTTA1t6n9gKGoq
HgOQTQG7MX0U83e7FGA+pzoq1Asko5xIODUeO+4xN23R7OrUG7Ba+SP2ttRcsK6Z
gGG2OvHWPoys2SO8/Zo47R2jEsCbdn4dfuiA51yYo+sNPAaUZlfhJXy3d3O6Y/Os
8Aa7dhzNYkSv1922Evt2mlDC0w0C6K9w0NSrdGHHm5vRyp6ePgccjJal0E54ZSPi
UFzfMyT7hfhnMK1cB0plhp3iO1h5CMzIivXjA3eJAYo0emEY8mD5RqIpTKvTLuZl
FdPvAZ2/hlhTZKzmXjiuAWdG2WGh8SOZtCrKkj15MRKA83NDe788tUh1bNAN6BPV
32d1IEPfNECyrLZ0t/6T398J15F9jHyV3WvITV5l1Ra5c9zKkaoxN/0uKr1p2ILq
lXs2E+mnAKwu9RQRzlARD0VzA/4Co13fifw9U0iay0SxCCgTAlgBQfmMVipU8OLj
pPctSPoWnJ04KDyNg3d62BtjAipDEky2dnunDIBF3dd0g4n+0zXI1vzEtS3V5e9G
hXh4KTo+8zNGcrAb+EzlmimRDfEAfcbMh8YUbm8cfYRTQWZurduzsnVZCvCPOmcE
YeqIvGpoD1ebdOAHj16WZCx3WL+FJfttmNoWsU7cOchNvk7YGefzG7V8L1dPWnNI
bygS3I5uktph0ybP5pyw8BPomo09rY+qohWjHhzJbtDrxJQqssdrZyQlquQpBhiv
Fwy+P6xGlhKqWm4v2d4p3nIPS8G2bPD7PRTiCdbJ6EEEF+FKpPJyWB+kTsrkJJOE
TIQIhu9HeZPTKSPEqZyO4XmJmsj09mlMxZdejGsyccUM/01OHvt16TpcRPC0GvsI
IC1uYEfveNQ/A/5XaqsM3lTujitXaphOxbavsNP5pB2NTOlcguFQdjYS0EGW8OMd
aQngghbrjq7VZiioYejCXM7O+mju+zeNwWgC1I52L4aqvFYzwQXVqmKPPdac9CL8
3YWHJn9GHPNom3qI/MP4TF+I3kPPfpHdhZSDYHDlxLQXcww1Z4uBqt9k51aNuO/O
NaBSsx3AgjsWdxTYtRRxDbEFakTSwmNJF8/ypep2515GvyrDKtOalFiKJDbe9RU3
zWTdWXMeLVlHV8Y9Mq0fZBU+iMpsNdlL4F9kc6yZ9atIkoXCUO6Do0p8g5gcRbfM
tAzBqWO276xd2XuvnbqCwdGKBuA7dIYw31IiaJy9JVHq+ihNJoS6ch/7S7dEJKRL
lcZNail0InYCe/W0LW8kSTTcf+XKr7KvZwTk8LoAvm2o055AjLEaNSG9cNimr3vR
k/z2m2t5A2gzO6bdDxKA7wNoACVFDSmKqCPJwSIToLg011hN6EsPJU7exyziNkq1
uqSx6CS61K8JyWXWX624mb1WegMd325hYmIGsrVdYDkolZaNg5aBKgpk7K3U/QZi
Hpnd4DRkKK64nBLRq9hHninlPXWVZKMUUsXkUEWa/p6S2LQKQOQ7IISuA3AB1l+i
R0AJsga8XvnRAPOgLkx4u+UDW0+unS4Y5hBnVS5mnXBkuvsa49mdXvoAW4Lid8xM
DnuJJ8UGUrwrkjwLHnc9Fxi8scV6KccoDIteOzKBGL90vCqL96UfcDkmAkrt3FlP
WeZJ5iFwpmIjOEVE0pR9+BfIYBA/KsLkL4otBGbd4tilCwFYvwJhCphNEnyyENig
cbVc2AGWzjMWV2BaBFvQYrw7LzXjgkUATtBq2s2aeIdPHJ4ZPBpXio/MvBiKZ46I
akGZsaTqWBVVEm7bKC38q5bEP+SzJ5MtQ3yKI11hF/WzUu1AcOc0tRjHfuVgAazG
RNq7KFvRWhu2JPXJ+iKYTBfidCXprvpw0OFuKlIBkavft1HK4opeisUS070rNDmg
vabJZSTnow/njk9ixhclIvV2ezfbA6LpGJwfQWfMToZtGCd7ubljBasSFIm/WYvo
HVRSG8jb+Rj2Ucn5EUIGi52tRgjsBOYV2bdAVJfIDlx2JW9bLSZXjey+gFKdXtCj
d8k3qouPqj2oProWWUbg3mbbLcLtj2s62Yaw9F+67AGy1BYR4X4SB5gDtHNyXC0T
KIRFwYbwX0WotMni7Qoy6TTMx9dTedRcRhI5CPQegy6h/Zlu0IbmmzuRMZAUtas1
W/gto++nsEhWdnBGGn5901K03RZzjP0QXuvpYrFJKTA1gjUFreNiZvrBdPo8gJ9z
79SfaOh7bv+MSPYEqXLwdGaqo8HT6O0SxefRUnqF1JvwLa5errmo/eMvM5MVx2Cz
roKbazRcBunJRbOnSBnGJp8VCQflYp4jw4A+0xAK5cnz5h9Zwul3n3qKLDn0ziAM
CbmulptQEiNAw8MQJ96yTT2x7iVQHBPdxRE8jx8aEf0IALtX2CbNK1wLTiSSnn6k
ppjDaV7o/si29HSRBCx6sHvwXKsxty1UlhnQP3J85PZS08wHyQPRmQtJpMCyKZaO
5DlYZWEqZ1k+m74ZdfUWU1WuaJHQXSsLIrLE3STTewr25Wa6pK0NWyvctshcAmjL
lCHzviwkjFz72XmFrzVSwXrCpmIqSQ2qCfjSawPB1erUgEKpTUUj3MWScTVNs4p7
rTEDJ6Lveh/qYEIZ7+i4xHWLTo+vftQPUYuyEwiLTiFVTi1FicE1KC114HfQFWKO
7XIJhr/iOqTHGdiCQ2FpzE2ab9GhHpoDtghQxwyDIpT62WcD6T1lDQbISGqieGRR
mg6EU2R9O29DsMz2g/CoJGzDng0iavNhPVUN0lfjUTkOJFE/FQmdoUO/7ZQ5yuAN
EBG+cvxI6Kes/D3rvpH+m/U+17uA3d/N2213I/5c4i0QL68uxGL2b0FBm4U+65gB
XXJc4q6fkgsFdVwSeJIbKZ0tU0hHrFJoR4+3TsV7GxmhM6z7ztlAOT24h+V64hzu
YS/Bc9qvOgRuWNYgofzECf4T2WqILedsAOJ3Z2Nf07P6iBYsnyYSQTeCg8/T2UFl
1f1pzzeP4c3yzB1eM+bFZk9yxUadjrsFM5hy03ow+nuwQOGOc/pKpyUkbnbijjMW
GTjId84XrD91x4PxJwMmgVgj/QlXjyj2mUxaEYp6jOzICy1z0ACM3uNhlsj/hB1c
wK5iPXva1HnL0wMRnqKWesPm7+3dVoLQXJ0kEhMoihqzfjFqgTmmrnUBZ0FEj+Fo
tmuWi21GAazfCkLaiLbsJMcNMmo7g0Uu2Kla9PeWK1mPpDuVI9brc2qu63Ngp+on
PfmWZnOvrXtO7UK16NISWMcCxGkJMGHI0Fa5o/P+nu8Y8TnDM9t4j16mHL7Yy1+G
LWxaTsaX2f2H8AvEC0LGBLNCzcE0sUE2ebs9rM4UPc7OQMnxvoEXsyBg6xZtEOfz
FJ+KeAU3NkSzJjElstGjEkgxMjbMnfer6kwdGbGKZLqLP59ss/9HioWlpXJd1VUv
0bmEVPmgBD/jK04XbVkvhS3a6wDdO8mzoam0Q5gLc3o0t+Bsb0NmKj/cOyEZpf1C
Yygu/jUKWfP5jqklRuIV2bWhQGKjSdgkXBRjdMLJccI9lxxCa3oWfzBqM3s8Jpll
pnXOtq2M9nHWOx/bMoQj/DnWxW1enKFQ2VCoLXQx2NPWxsl+6TZwpnAlsiKOJG+r
KX5/zTEUwOmCjk16pgwPW940GKn30q2U2XDaP35ZQ9EnL/FnyB4jDn4r6JfOmM9+
vEIzz491K2sye/gMz/h+ZoQUMZX53jYYDNKGsvPImdCQ7uWYm0ieuyvVWydNRZ6S
Ui0F0JThxeiqri5R8yQAI3ynv1LWpdTSfQXfG4NLp1Izy4Ig77AIMvDvgLKJ4LI0
ZC67IjHHnsbY51proNw4e3fvVIWERXosRroBqA0iuE+OJkRqEgWllFB7tBS7r80o
Q6y8wGA4cDh7hQtq+GpXfRJpzvCss5GymYhRGgNNEPRzYE3eOcDlbXbDJQvPgBZV
oMpI5wNBcrYxJJKBRGtXDF4SIVweZDTHxAyq351BY+Md1rakpflhwvHRknhz1uSs
wdOE8rjxHQUQIIJUbG9hjqgdzjbK+Qf9ztF3q0iFMetR7eODyKtBBJWs2hbvlf6R
GaKrWRm2QX8BrYi0kKlq5LqZlo9qb2LMNFt4rUoPvn4n+twfNLvaBgfKXm7BjDTH
AHPT2GJXj9uOFf6hMY9fpNZWcN/+CXx0ybFGhn4wsrMrhWsnCnX3kz1jqE4hiMZK
EEtk9sNEgtEWxpejpMZNkkkZqIh2ssyrSj4DvU0nwW2GwJMZb/nXX5Waxaf2sPfh
r3I/eY51xMe/SE4xN3jtn7p85WeSEnHjU6faBlmAALb2/hoBL1JepDHTvQXhx4v/
H53M1PXqJQrtM+hv3O1J7r4DxPccr7Ey8mdnKFGb2obv+bmQ5PZ2KJfx3bEmdU6K
sw5+FO2CeflyKwXklAzCI4D2VhsnsehAlNTmb7ZBxbd3RjR83F9Xmq2QyZtjrN5c
WoMXIU1bgwasUW9B+WDqFV+a9NmWdoEBLKCBQMKAzF3vAh0gN5zK5QBL9bIZpGDY
KQjZRQtkoj+t0JOOCFqvwP+QTsMqZm82H0Il4ARzW6OOkB+/rYYhUtC1kJyX1eQb
d1CkYrKBhqwtjtcuy4tFl76epeLgAu1jpEFRLaOWTQY6QoJhDqcnwTyakJbKrkV+
poOHCG2oE/rYQwFu5TtmMcjHUgpLtyNkjq6UuJSLq8A9CL9r7EBpegQHmKqwTjH4
YtX2QQBUY5mD83qN96no/rDy+G8vYtQOML7pSDgjWYZMTwWmimDRUaVDO6DSAp27
cseH/AcMFAkEAkUPOSDcgue8EhMgKZRSNhkZ2b/d0B78XMevBk58WlONLUpgCetH
1gq8+wZIttLusA/BCcjjP4znir1rSwF8nj5lNmn69hMNPfb7BNXT8aWFLcrP/G72
YtbXmPfceG1njwiAXL+uWwW/O64jCwzEbTHqCr75cD4CLlbSlfhnNIVONpuA17HP
dxyW9k5N7dZk8dhylivqFDweKWWIJwhbE5VFiyd+ddLes5pCLu7mUeuSyRXZ0jOm
RDSY9d2LBhv08u/zkg51g4Hto9k4Iu5QVs+5I320M6Wue71uHdpajjHAqWKsYyyh
tm1+BFTPlLUonzIFiXMY3E1pMbW9a18WjSVLh9XixQD4rdxCbxZN51xYTS/zNT8E
5TwJfzmR1RN17THifQFKi/L/hVyQvUGEOHxpfoKACYMFdvt9ugUEGI5oy++J+Qjo
4gszyO3qfYhDJhX8lPdnNlM+k6kQKRGnwYTkZghMEbiMm0DOxLKzfs9ataPhpzfF
j3oRxowXrSy4N1qyMEA//aPnCaCvfbMR9V9yrw8h4IuWtyFYeG9SAAPP74PN4iil
1cztwlW4IDbRE2udfwyvoNoW/qmkgfjXaWOcyicxSMVttH07BKfJUlWyKHfA1miM
AybV3ZBUvG/7bi93IEBIXBjBADtGXvfP/CbS8V1/p8tk4VS1CeBwr6zdPLkm9ljJ
/oQDv8Hd7YjR1t+n7K4WHdRpsQyno8u5jxufIkSrjoS0jrFIe+0ljsHdRNexR6R1
g+7ZH2FLEj8ZHckaALOV7cfX6qc3gCMVT30t6rJUCYw11eF/2KMPLi3GYXezuGb+
uG30JcPgI7nMH7X6BZqI3Cxn4bDRsU7bcIosd8vfKAuXfVUNfhdfO/aio3Zi4btB
rvWsEP62WeeyaeGFxEEfBcPPukwoL/+ar3Fux+ibEmTNR1IVcBE1NVeNpXoZ2c3J
fBmIGoAUWMJKkTnOyhymQrW+DUhtusLu6RGJtX9ByX8B9y6/s4fJs24xNbslhSxW
buVQfbopLwC5WnGBdY2yADM9em4ow/45TgQPwTwthvBnGsbq2S6JtfrzJDzCjV+q
GiovYPtnwyv7hffNCViYraxuXS3Bc4nU3OcI06Jk+hhE9w7iA1ZowTC6kw457wKr
9uatpkuAVcupYuCSwX5CAbvURkvctKrmJnGwdC/XLNym9QzAQOjxXsiNUJlPFmG0
E9Tmh6jxt7IyZlyl3fJuC2se8hd/pEtvAxOsa86+u8UT6WrB9IS8QEJ9WKej5Haj
28kbkiqbQMfBi9sey7d55Xm1ymD6yvNiofnYuIsmgLOC+aAMsko5hTXPXCHsR93I
AjjxjHrT5fULMMuEhlg3e9HbRMENr8De68Khsyj4IgskI025fcCrSuMgDc7OV5En
alYJ2lnKyOLx9niMxpkTookcpr5e56y4gtcb28cV7zjSpv9KWTfQcrtsS7XbkJMb
6fOgACiVJovj2j0eUHAI2V4Y2ifQ1ZSnHJVfHzy5IhwUbTb/7a3qiFolQ3FBiQS9
x4YdoZeHpDomLPemwsFxaLHd8UH+efJUYZiPkINy4hS50grfrKAgopWMzQimpFqf
AnNYSrZhP6HZUCGGia3ThW/9blIsToqBI1mArCTuHnti5V7OUoXnjeV/P2u8bupx
rhYv3h/hABvkWBNM8YLQ5Mn0fUuDMFw4/WDhohDqCX1DO+hZPOqRobJHAHx6vY3L
Sobu26GYdYs8Ie/U+U5aTYUIdWT1rJNy3OwgtIlVqf8f0uj4dtF5KQmmcNiTiuYU
TyiSMhG9ih8tA1DmVLw0/Jb/mePJ0o2aSeQG4Sucg8tMrfdhqJicw2CPFBA2Mb5l
hO3ILhFDMQuOuU7yAxcAdenipAz+bx5DkC30TvqThWLryGY8MgQx6K7rtBUu5koE
H2m71v6F87iz7rcaDxJRE69dH4kohpDyYAbtk7P5frra6/iKaq2kb/SFuKzYPbOP
vZ/pGav0Nz/86HwtJNBp4wyPdxLGxj26XGVdVlkWAqF8kpwZvYpKvlh2qTg8mWgy
Hgx/T1ZTztXwV0I9saVsf01eqEvDmaxfP5jSeNvuPpP6jhBrjTGNplPlZtUMDpMf
NMtz/Hf9F/O7nvYO9SNoQivh2pVQGULYfXaz4mEW7JjUCiXCp+DnabQLRB3T5X0P
xVGf1ihQ3OZWX5g1Lkded76ZFskXfDoSLSx9WIJYCCSxYrqbpPyIz6uZNImDYn+V
Ws2tNInDnCGiboH5qXnjFc6W8bCkunmTXPgk8DyLZznPP2AVdV/RlZK5sU1IAikG
R1ZMBkN32uH8ZXsHDT53SbfT91lxwwXpjWQO1iOFzRSP8jVLsPBFVVnSGqGT/MP3
fKjW9LGf2dPW180E9/bAKmCXPqRTTNTkMN5xq3z6J8ayzzY3csgxdNcEJvLgRbGe
IaFp5maomjR1XVNmzLSaF1ssmMy6akUS3WwY/JYHx4X1VgCINcflQuLNAxKITo5v
KUoPH409JffjXcDIGJ9HL4ibS7h4f6ts7PHOvJCRS5+DqN58zUY6xRCV1nWGfxyY
9kKwO7HayjR8jQNBjZnq0TjrvO7oWSQ/Ob+IwexHpQS0Wehsloxk8PCR6hjjT/bK
Gwnhfa/mpMX4sHOZq1LCwBVLjVuVi5yZ4dteT3CVaVgFiw9eiJTvftZTF0XRB15m
UwnJ1kmHJoxGduInxbVCS9SIXhFvvBNEl0PFFq8QCSgLJBODUfWADlgdSZzIX4xN
jS9/+DqU3VYltabZ6BMywAzOHEBq35EOjz9+BhV2o/jU1V7Ki2I51DMypwSNUDRG
5IAZXIbH8ofYhBMMwRagG2RIsGH7AUemwmnl8jYl2VAl/dI01ttLkcux0X/Wyl32
pmULwEyH5Oc4BpE/W88lAWAzuJfQeIK32P2IBaTKJsclH38xc9lfYulpvPWFcdtA
wVHZVcJ0ZPcKb+22YdPkH8Ln3LHfJ/TPZdXDc0aMpo5Chg5wRZKzxyXFcuucrsh+
7Ph59NQmYhAeQ3HgxLKsBBTivJw8LiWUPP58tnkFBIbHxYOgHz371Z9eA3BLle4e
I+y/O2/shGw1yTXwIKDsCRefktU597APbd+XtX92z/NNwGfLWkk7+ERZXqNww61K
gIhRrFes/QSD+azsEaS2uG8kwziuHcnFhM4r/5y2vH+jzRFe3ZxKhtZM8WJM/z5/
xJcVjz2dy+ugxsM8A8OimgWoiq12etDMAFkDlijLRS39Ej2Eh2jUiGm24boHEeRk
qhKOo/45E9mKHDHkUO9/f9g+WZXxIK/nAPcS5yr2hh9l458vtJmJ1TNDnwNDhLb6
50b0VQ/Cd3rMbgIJFm5EZLu4LoH1/QarQVbJsMb5qudCx7Fxl7OQTET5GwEvGU2V
zVEViaXvEY6hBkJpM4QPQ6ntonic+gCoB6oBygXbdi0euBkLwOays823L2oOLwN7
5m4QfNuJxiTDFUVqdPfi32UNYkNuyVBcQ5e0Q2IMdwl4H7sbZFnZ/pNcwWvv9HLu
4bZDabbfaoDUGRljuye9mlshjAfcVF09rcz6i/bwbmYhwZohOWMf+GjEcTuKffj5
bgTlD4NJm6Mo+eIHgeOGF4/qIZMaXuBWybeCGSrcxrgchLuyBr+DLgOpTw7aZnBR
Na2ZSfgH3LBiVhO6T+qciRFj9V35QulvF9CCiVVhuKVYRHmsF8aMFyeB8MX7NfUC
idur0JZBY89ekg4J/OaR2BqkyxmJqOI5TNwKaTzTxERtZpW+uAftYLZPJ9BqyWaa
x2ujR4DJPn6naiwml82gUS7FKz2wVmsuGOcuEfwYMq3atonG718FNBP6AgI3ugFi
rvdg1XBLwoIt3EGqMwIG1Cz0sPPReWOGhylPLisirY6INYpg4cs37ZWbPL9kZEr2
vS8okwjF/GKnBuHlGS6EW1C8E/QMIJ+SI7dO4LcgpRJJbWOaXwvt4v2mxfIrQjie
ZVSmu+bV4EP1Rp5uCJ7lSpTa8hcBMjS9/xCXav9IYUB+PFDZ7FsJeow/+SQ5fjlv
WHL9o7PLDSDYfoa/q5mogY17C9HvEc9I7VWG6MjJfBDJfS9s7ksowF/ayNQnxnqW
4psTobQHKYrhhiY679GrjNbr2R5d/PTxVEKjWFMJC7k6hwZZBg6xkX4YYDR8utrs
/XWjyejbDTn8LeLmkYLZNVA9dCIbpNDX8qnei/tTGUkt38ACqvUC4if5GNJKyBEY
0C8AKvItgkaJGoYxvuD67EDhlPv8T+gsSKYLa3h+rBqx9oD2KBo62T/r5t+kXZrj
PNo0FGD559JELU1L/l+euD8nu1E5egTQnymoMRkGwBKnTqWfZEJwcwmxvlRXLBT/
zpwzHpyzc5vfo/VdVXKmkNCRvz4CWSWNZWdFsod3n6RBfxoECZYGb1NSSV4Ip8Pg
mwsqiKLDh11PA8S7myW9C+iUdDv2tXHqGF4NupvNOPs+OwmktL56QutwwD4rL3bd
LZEYzmncBJI/VzUHSTq4iapfnWDqjTRDTvJUyKfxHRiXubrIIfSHWygAL6yvAfWA
eMlYRB3Tm8DJvVvwgSyi8r95UwZaY2jFOAVUkf+/L1D9QdD4+5y8f8Bz1XjcPIJH
sMpfM0CzSs5+/jFV8CWftE3meZLb0neU67ghxgSf3O+KSWZYEvdpn2IsHOhjeO5H
F7S5PE0vUYB7hwZYQWfdn5KpSYbVvT3oN4QmLszLW58keAcnfGmMLizipwqjcZKf
5CoJwGIOtTJLzkhP+YeOM2yvF5kEl1NLL/D829qpuwvHLlKIFVuhBcINGBxRx45S
QhoE69XvJdHmiwkU6H6+OKuLVD/un4bIGjMBCEPbMoNPbhMECcpG8vZpPC7ATPr3
C4a31Xeg73gkDTHfW68J9HDYHop2+qbL+EDJ2g+A+R45Aw16nuESkHIL9aunyVdj
ISRZKn1uNdLT14hNkLKZJWoTbJPKxk3wnj3esnqQAda2bM6B/r6IvuUuLwOaj86N
5V0/yeA4uC+0OdLTsA2FW6miyfj465+m0hXS007dYZLgFXFSTd1v69V0UYWHHdg1
ajRncK8r51pNxS8EOZw6WEhO019hByLaMR9ROGPlaBUyO/XZ9uTpLITjfxG+tJnc
a62WAaHfyHWLNB0xj1s0dJ9B1VKs1d/9yr+FB8gVo4rzO21BUYo210hV8Beu5qbM
/J0ksdtkeUS6fCUATYgPUVd+yet8+Iid758g3kCkeHfJC7I04gkZ8E3hFUcl/bZb
eOpsWPjhF9tcDyXDNGotYUknEzRZ7YvoPPY1vnZ9IMeQCsFMEma2vfgwOjDdwZru
fsxGWoG6+up7GtD4CPegTpV0GWk3I+9AkkODXij/WM5hlL8YFgfRHk+dubADMMaf
CSkd1xAgy+NsR2eHeEl4NJAFZaPAqxX9OcMnTFjLttVsdafiYKR2Ihlb8SrdW8CH
YNdKNlAlJxOm9duCHA8D2KxncYz7/17yUG7Aj8WNMYvK/Ng5Zo8rFKzBuxx7+SWV
DBAPEx+O+dA5pUI8CfR2Hwe5UniF0UO66XrK1VUPv57VCJAgE49NvY7J8rJ1VH51
S3dYi/htek97A46IJF5jvg/qEYMV0hiSY3gqcLrJHBQqYbcp4/LhXI/Di+wN02mA
OYa8COOvcr+aS4K/P6JkV0ZebzRED+/Mi/8qApPNcXGViLiSLC3lfEoaNKijswe6
AndaK92tjeFMOJX5i41zn/5g1NUvSCwmn0s6Z6fjmg1hJDJcFNlXjsd6O1KAcYQH
WHLi5RH4EwotBHv/+JkrS272+aYVCuigX6RGw06PnEjt7bb6NTCKMKfyW8keDHpo
+HmwSrzgoASdyKn3dTDXeebba4v6LN379IvB5euOvCaW2ATRRYBUJe9PawgFWEHL
4zoYDoCTcNjIlg8y66aXPULxc5x2T5Hm3saOwklOCACnYgUNURn2E5LWUIUrnP4k
Stpfb8HxGSgDiRpjirT6m+v0hVFk1FJ+C0S8Pv1CWFFm7sVfU/+uoY/2A8t/JEZZ
1qUcuz/rB+ifgZtKlDmeLwa5vU5IDja02Rmkjd/DzpcvDZoKgXv1+qzKxXJJdjq+
Y9FtFIm2adYbf4r74kP9Lp73iZx+ddMW6d/ylPYrLevZejz9AphmIKk3lzwjbqGc
HVhtANfZaeeZJNeM4K/kCLDdCFywSbyX2lM9NP5vxqWyBAE3XjEOh4Mt4FuWCxrM
2vguIKMrAeNI8JP+9eEhtcNIROGxucj9cdijT+etYiY2zKMEjsBddcIkOcpoL74I
kYCyySNyTbq4y4nEEtjHA6BrM68SLMULjxcCZMeNWWr2/homOxweK2BppoNRl7xD
aZJesNBaHJuxwM4gJOlb7aR6FwCdeaHwpSRzwOux+vHCOucqREZ1mzdE84bGo4c9
rexB2q1+oPcGOzYc8uF5J+8DCtl49N7ZQ1JeaQVA8cOrAiOmMQUUEVEfLLOutNWZ
8haPUC3OsInT9H+O3Tg9gIkXpu3lG5uCE+KB63oR6iBwbev+qmO+1F6iAc3f81mV
97wb4UsCzrHN1p3UR4sZdBmn3EFjz6yB1wSarPxg7o01nXW9gurqyVN+j2Hb0G2R
t/XrV8QrdhGv0hgoGXXMbrNb8v6fEbG+bNHn9mt5oq0LJtaVldBf7nezjTfuxbaa
qQirF0ElWOqa4wPQA7LZI7CA33mqFvcTxbpJnnIS8RdULuYPW6+g3WTVUtmmKzhn
o8fu4Wa3UEaNQV4Wbv1IKq5YEKL2+eXSayDCLEzwUWzjE1Ah2q0AOorvkXorkUMb
MsJIFM6d5OMO0DPFzbWkz9NGffN1nn3+ZXxmIszxuvxlrVOB6OZcnOSR5CeyT3Lk
GKmp20uG5fjO+bZ5ivQ4Eucleu0CgWYG6EovTH2Gzd7dpJWsZWewRcxWQU6OyzRF
sS1iEDQZfqhsitydXH58vJhL4F+lxGHfGRcM+70C8V5CPHl/qwGeR8wwcKG2jGnC
nV4hoVtwcnypiL8gt4bc5Y4bbQ/60LMWB7sq9ANHLy2tD4HRuUsAkL4WC9Bp8UoO
b28mEUbUFyrnO6XfN85CcRcRv2OY3F/lwbVDZKDRxrXjtJa4PtFFasRlIsrsVo9u
WncGlTY0Rr9nuCZDhhRCn+E9W9RSHf5qzhQ+tGvgjOiZwPdObjjw8/gUg8Kw0xp2
ZbaFVTpG7Gv97KEGWU8PeDPzVftSuI3296lpbf08PeSRhmqsmD+G1Ap9LdeG8IaM
+Yri29acDo2zDa7LoAtrSd10z0lBJq8kp1RivdI9HCWb/7Et04C+E314B5HgsWS2
xLQqw+/nO9QM5U7TM+ytsLBXDc02lFz9Z0hJ8N/lwKw8+qPTYOAkHtVRTrSgeaj/
NoxA8bIx2tQ83Z9J17QhHOAZ2uj3muaulrvNpiNw6o1OwxU7E78dFt5Guc8p3mvT
fTxdDL+Qg57AGlK8pc0mWmUL8ErvyrfLgxK/N/SagSIKWDmImi377V06nVnJlhip
G9zoJV58skTMkY+aomJknPzb+dj2G17rVU0MRW49deKKvPxJlihseTISVyFdthkj
bsHXd2/20z1vL6wrIMHGdR7Vd/W+85BYHZT90YkZdmZ2yJbH9EkfVT+ppYKPocut
ytAQ9fFM+7RgG2SMpX7dGezVurk/vE5+Xblw7hMxi3ckTcQ1vZhgx9ElqmE2F0WB
AkJQqKb8+HXinR+WXPYxC1oG3qzwRKtvUCThfP7d4WHcZBSEHHoXiynmAafYRUfe
8deq54Dv+utTOnnOBa2h4i5bIFsjdnbo84kvXbCnbTCFrbLYXK7nEN6g6R64SFO9
GnhRxBDjKlpu5x/Baut8yn6OJUAh6muldM4PIRYXoiXBB4IqMA9bdXoRcoRgRIaW
1t7Oy09ODJ0/HXkMkc+AqH2kPQmmsA2cOtZKgwAntpItdDpPDG6fQG/rvicM/t7J
gxLwKZBTXNo8G9sJ2y5LGuHZta/bOQxGa0K7ubXPx6TnTcB1yaqkfJHQeQOiBdf7
ANqrdXhnKDXgy7cqCgjF7ONicVqNfZOwwWuOLygSBrqBllAPRc5z5zUcQ8xYYAlP
OQ9JrZ41fGYTHWxeL0xCYfa4YllNCWrwa+YuggoP1DXSTmj0jLqNZKmxDvsCIAy/
cfmX9p9jlxNWxDXCVe/mXVT9J5xlBsCGgzLdPS8rJikhFjVCJSBzMhLevde1s3N+
BK4Akw0BSXBJeLyWlnIbqhY6OrzAGL6fgoUBahfYpbnCerGzJZt4gu0ACyVaLDsK
EjVWVBaigR8OzFmIYpfITorsttpPawHQCTjCEuYaWf52t0XCG/9U+m6clzOS6U7U
ajTxIKBD4DAKjUkMnA0zWYeyz38WMNF3uJtGOp1krHCAHm4NvyjZGXHOIMUrpAnn
MDLvDBKaldSfR6CIjLhFSs8/ZKuGeNIcbFPGFnAYHRso0FnCfqW1sW8M+f6ZXy1C
EHfT2enQ73rGsgsAGIZR7FZZ5L1F7Hx/q2oDU0G9FzByZZNv8RzLnTRKG/bSgEQl
l+YfhOs3Xw0nLlYGH0Q3ol1z9qtsbER6/MCaTs7VvHVZxE/Ycr211AHFv9CT6bip
KTNAH+WbNrHe5fTwlIOecCcD6+2koAfqIZ3pPhVpF7UT2pq1d8IM7FQom1As+PLk
fo1Myqf+sRrqxFT+cvRHQBaWhKm33MWo15ekqkff+5iAJ72a7kQfVP9lb/CrFJFT
3XBdjhA7DE/uCKIf6MBHmw2J5OplZHmu+MbMNRMtI6GKiZM/7mlcSBjMN+k0WpkL
CpO8x6PZqx3FruZox5QU9xxopSCU1t4M7UTa/6VM91PnYNcEfqdwjbgslSmR+xi7
amyRqLA/U6+n+aDzqgg/rDQHNPvvYeXwDwgtyh/+pB0IWS5Xnvlp4SdcmpXt/tRg
FFBHfvD4PrZWafDUZJ4kH2a+UF87CFhPRWP3rRT+ov7moj7pT7XItiSuH+SQTR16
gpBpp0uSsE8VNsMSwL8/8Nv/frE8tBi5agle8TmetZHflUcIhBA1FNuwTaXgy1Xk
veabiKCguICJcrN2HHSuWDJ0IF3JnjIXmjuD9nVFmF9dPXSvf4/awKkwAJdpXzov
ZmwJRFf42eGAe+NmxLmwpyPtAsHLggsDq58D4xnRoPf78gz9+S9KHtTzX84bCtvs
NnWG9UiQmfvhw7OpzSvC2XWPm9B8xvkmVg0u+If8/GuWRFgSSZc3OlJ9qcJBk5HP
VoX9a/pGAdfkSXLlMsR0Am1DLHTTMk3Um+854YdhCmUMIQYiFn8u7IOeUIurQ3yq
OaRNsf7hx9u7lwgaTeAiz8NoBMhlpANw8NeQiA8TORnSsA16Yj8U2Zu5ycyg1T6A
HAFuNnVSqyWBZrcdO+oXdiksgd6hXQIqSJCKACNgG7pwD/cNgFFx3PSLM25/Yps4
mPmWq/ByMPAuPbBsjDWIGKaAyLl1tjdcItwkkn7m1U5Y/ZmPqfDXEpD/uMOY1jOD
+eRFODtSejxYPRw/6XjtnBwwXimyLlLfiWgWC9rJiV7f4haZYXYRdX6N4t5BhZsx
9qrOOTqwR0shFM5cgAEbGjHft84cVbWV4JERDdsHhfGs7xn08ZSKithP4Xfw7iBp
8B1RIWfRAwrI8aDhnJ7QNIo7gTY2xtRIMq67hZMQ+nbr6Po1J+oDlUbQvgFCl6sB
rWG3y4OsVo8DB9EjhiIkKreQUu/KMXyqSAlD8/u66VrG9SV3vVycZBkg36xV/aRG
xCzzojumMh2vGi3Zu25R4JfFwIal7tNZNxa1rOl1pmunZ6Kf/5OzZ8C48FltFSY5
Yjv+VR9uwT43OrO2mXSgtQknOPmP357qhR/9tUyaA7nie1ceapKPxheTypRPh5rw
3MLvafl74LkrcvFUeq6HDA1Obw2DomLE2OpswdbmAyBz6yNaYUaolwa53Cf2Q6ei
3reV4zeIpPthZP0NnFj16VmEOlKEbyqGEAOdeplzDAv8LkuYRGaP+M7aaTkTOphX
ndPKoVweg2Lu/Dy5ym8pB5asyIe2FL++5KJmINTjS0nwG//e2OzCJoaTyk/pAdxK
NJxOiAW8bNQQOr5ZbW/DN526WctmQczVb4hrMJ2WxZaupx7OVe6gJ66hMcSZQAqn
n05px3N6VwQYG+JMNX09r4R9Y7N8e3Xr8xzEUacnaV7x/17kkIw5ZdSJSMbF26Bj
V3whmoGSs+RAUQZ345EGuGo2QEf0BToqEd2GuxpSl7/0kAR2u6yCA82dm/7JH4Rt
gDIH4pLlKeOR0n2fHlVJtaQSmUargaEksQR4BfH6LEOe/U3P19tIn61tz+sXCG4h
UfbGu5zOp+xUKyYgtqjloOf6sYYfVUh8Ela4LMOfTDFOB4PmS9FZND+n6zLyyR6Y
XuX6Btf8/C620Q6i2jQi8AjXfsXiO/aMEFwqbA+kJofSbWbkGpowqTJ3e8p2yPz+
gzIlKCRomoqLXWscxd6bUsyuPlgINkQ4ChCytS7mVKGau5bflXt9NO04uYnZ03/+
hNt7UjezetYH+Ci6JzFZyjBxImky4YkaVNtkreAjNTHupq6QzMcuC/K5yRCVdbIp
xkvc7kwtMueUJsdt+mngkbbwPQKove0ZjnGEOcwqly6dayx94TWh+x8K5Sm9GSq+
tNyocJdLg5dRacUT/9FZPz6rD4uA+wbi/dy1uGsKr4vvslZsLC1yJuLLrk8xIph/
LfGeFo3DTQpXJzI0ffR9IOiX1aafpLpK8TPgKpThRY4p4aOlWrsBQVT5Yvg0V5Am
m/f4FAZyRPFgt09i5ayw0nVlPojU+mZ9xhA6dqhCT2kgxvFm/LWEUu5GjEPaoXDo
9HcHQNMLW+nzlStU2B4eba9GvImxJPiZKD39comhV0PJiTw2dIDhpNRtRCVMuQTP
/gLsml6n5gyGeS6I3Xx+ST8qmc5Vvdp7THoIofAv2f0+cvxVyKSxaSxea1QNr196
uKpJld0WNmexxf1bNnlhta725tMxZQ9RdlMj+dTFn2kbzfGlDJWh6qtjsFHHSEky
9EMVA4PFma9MwVBSm2BxW/VZZqkhofYcWI97JSRD8bOaLHEuAMcHZEtVQYaJT0bu
pECl77URHIPAAM/OMa4qX3GGeQuL8l5AQHe1lSYL1Vy5Juj6SY7VZDWmQJ5QK6wn
tI3MReTTKIknT2plOEuazRGWkd7e4GpHk3IwLucvgc3Q+ASS1wFio9nvJ5g9jCkg
RRknSwt98gd3y/VGfw/EnjWNVGevNacYTf4m+NBK43MHudmIfaO7RMIulZG2ZfC6
ebNWYvvSCtkoiEx5aVC3mQBLkZPZq9/RhbpciMskM5ITe18KY9xb/a10ZMFzfwMQ
cM7eMJGw3rLbh2iGsHGCLpODOtdp6z1VWyxFrKFyx1rxA3RRbdZMaLtFKYlHlH7y
9Z5JLFa4dIgrIdxDbkqYSxe33IRz2BcIFf3uRdvvWx2kHOSiF7AzaXAk/cayQulC
bKBojSU4Wz3B/xWi5oiIjx3Zhk2d2QviRfXL/U3PNQ+DnSJK/gqrWuBjjgqEqkOd
qP+uCxA1krwpT+FpmLLRqpCW3Xo1uu85hwvObvfRotD6F5NVd69mMX/8m/E9jqcD
bI1vDHooHVl1gszBoHy5KbndF2QKCoI/d9izaWo3JgVeqw5h+sJy1Wkxh8vQrEmv
ztCsl3lhHoL+Cei8fRncDtKfR/Ide0kbXjEmDHZFVLMmDsWoBQGiWzpgCOhr2ONB
dAYhOTDFVls6+Fnq9n0YWQwkWRLNylMNzJeEmNCoa68labz9W/t7NcyhXxy20wLK
Zxy3t0eZV/D6Li88qyxiApC6JdsgJzYbUWMgMTMAAgxnB9NdCRnmY5eo7Da/yM6n
jretc+W8Em592EAo1TDQfHtAf/zkJ6+5YGROZ0RWTOj5t+XyF1615sgN9NkY8XBb
3bw+1KH0TtC0bHFn2+5TFx2LW79b7OiLw2kZBVXZOKMHY5vEazmwyC4okeN12tBZ
j4TMflr+Mom8Q+UzyC/g5s4aZC3mNYOStpmRdM05vEq18viR8nRhkQi1X4Tmz/1/
0CZ4cOZezz3sTBaXWj9pMSuLv7EaQHS+JrVvq8I1OMgsZKp8HYDLoR7J7mjlTx9l
1H05CfKxtOiMhWm4AI5K4diIyxtFLq5jNcdJ+aZT0/Uu7Ilhndate1TkYHgvReuC
aMZFAaXOEu54Q09dF76lSlksvjoH/Q+YcQeIndSyDp0Fg8orKsmz9ztg4OVE913O
C4fVohlCNQfzcWojge6JcD7zjrFawoXjbWC8HWVxHII7jsaiV0amgaS8btaWFIoM
4olo2OSPjO3gELKCQZJTCrNOEKdEMy1BY0yI4cW6AWKRgUb0wZT6b+ODCcqqYs5j
yCNV3Z60DYEyYvpMVW8d4gyiIwT5Fb0O2D8f9vPlSXexgA3bg8W1yEFSfWZsfgHh
GmVFfiXDOCXJiRn5mk6vXto+oMED+0hNffERuuUya48jFRZRUhXkGjnxpZG+05Mm
ReVG/nf+tkUnMS38kaJo7J79PNOaCyRIQeP9SXFdzKzJuXTHM5rhtjGUmtXd6ViQ
HZreeVGMPxK7PZ27nAy1qx/cxINRpnUJfjWeuHQQP7/9UWeXQD67RciLPcd87pvW
ukwUW6sKCGyKeTjoy1ZRQdKPlgtIk1I63dVllR5fFG3I+iWqtdGcJKUE6pFmU8NL
Qsu6dQf3/IgYClPvRoY2QRx2Le34N5KKQ3d8aaGfjJr4w3K8hPG1l8GYUM5gPb9o
Kbjkae4XOmFOZkcTUtJTbN5X2sILqZyK/jP36NbpONn3IwOSIldCFFTf34rpcuuO
wCQHq5sKJJC9skliyf3IWoTn/PWASliOr8mdOaZQ6LqDV6eg+Ry3gNweSVHzTac4
kM6+qCzMgS/E5dgQ7x++iPeTZWSqNxeCeK//j1/H2v5X/FYxDAG+X2OwthF3OLoP
kmza5V9OUFO8FKtTtBotSYypvcdqzlcmJZswMjbBhmw0eCMRYPJKdEtATyoMbsf8
S3KzBjRw83q4aH47is4hfnvGLy4g83uD9FwRqnVR/bbqpqMiy1MRAvrPzuZxx+t0
0kPZG9/QwP8+/BIGOerHEOCtrbG+D+7DGIE6+YC0wNkz645cdJ6j9sftCRzqQLI/
dFht7BGq5XKfO+z4PHnVzpQWat69cOPCk8j5+GBmew+T7GTZJRctn9+vy0SH4ccA
tb9wevJgpdlilFTne7UTORsIOISXRz2vNYCT5C69Kt879iBkw89b+QwW60PEwydo
iJIBES+yrX2qFueyhSY2G4zj83Degedc1OFnYwDOOvQ3L+kFI/zDRVa1zmcoVLlm
GlbflwyxVVl0u4AE8VtSlQkO3xv/9kVO6WfpkD7v0oIkXChq7B718ky8LEcX3nnL
vC9yLNSRNb/VexjrzvtJW7nYj6VAeV4KHmjGReEcI38nAmNsbKTwSdpDIM7YyWFw
nZExLThU55gAspKTzMn/UU5iO+UFGWbM0a3qAZk7yI5OuY6ThteF5Zn+LbZZVpxp
PIlANzyYupoqBn7Fq1SNs+dei1khOPCchNR+lF9M0aH8AWllNqI6L8Dxh4Izxwme
b/byHLPpYUx0q3TPyCfoYF7FnfCQ+CoivI2yJfNjxa5Aq9SsHLkdq8Cy7G98inCC
X3tMWurb/d1A8jRqJtSTnaF1SKOoxNJYDQQp2bU6RYAhaovn8cxFAicZdnsDtAXl
hZ0eP2sQNWQ+X7+MynJrmwMdhLpYf3a1cIXobF+gJ2wBHtmKpP4mytEbgocS7aZF
8kbsbr34LVpWa19raGmc/FOsA+FVMpZTRSbi7AT5ku3vxHV6wzi7LJIkj2X9vKT2
/QKh/ruUfKV3AVxQbNPF4WbQ8rsMxDw54FZh6/y3cK6DK0wv3enC8fSMSeDv7EDU
DoZJC6bMULyeQINn0kEmVWkpBKJB3Okj7wGOLo7wDyvshk5Vb1xN54wrOzWPcAGI
YcxvsFfnRFfpLBDfhcgGN1hkuF+dSrqoAuL3pUAYLJAz2nVeR44oSpInBhwc323e
/B0tgUplyl3CRuMqm1cDnZLJ8leGnazvMHJ9zJO8GXjviv1zWSUGIHVN5B+ObgDj
KKMWDodVohea6rQCS/Vi13Vta5usDawzlcGscGjLb07R7f2/4ozESlrflDy4fovL
c5FY6orVaBkETRVZwsn8cp2URc7eaaq6C/1U9UAXlOgAjysVCv71TjxtStXKjh7f
3C9XlKathRoRZz09JRBQrjUv09k7/VJMgQF7RTFlE4RKg9E4vkiInWLJ4HVtSWwG
GBRNtBlcyH5hckdsaaNvpqVWa3oq+KMBreuu4JVmMd8KPsNIXULEwIba91AyH/tn
KIIHXlKKa1n1wU983nPmYv5sqNwBwlQ0KNUDGtnBBIL03nyks8iyMObuDymfUemi
Pt2VZ+YpCCbtu41sI5/kBpUpiZM7osMCUAMpnsq31e2Dx55Mx7wkGR4JXlZlAcow
Zk8XS7jJemvHGNn62MTiqjmNxYIZfz1sl5hhTgqudeGxxyKWUa1zxEGNF+NEzqyS
7iObrM8U7daE3DiJVCgruXdU+oD7J4Z2WJ6SsjIZe6lY/Zzc+Tsvy+x30OAkKJ76
a5CadDF7vN2WBtAARHx54p/VeCikqvUNQ+6fsQU4dadzFPnEaktzfDHT+DwBWnKg
35CZJRzX0t0XpkECHlDOTE3MbxEJjp8d6HHJYOkHdPYSaNDZInwmpEnUAG9lyXHb
rWBBYd5TpmcK0tnav2U9k98+ZaNmjZA6aeTkOh47XXqckguMbyzWC/xE5FRzyCAJ
2bgm5O4U3KCsyFQtFKKN/PCweVtkPGDCGz69oI2zmxlbqDZ4bxWoovbpnZoaXM+f
ADUqX6sghcXjMoFIUNiS9q4cq1SOrCvN1RFDtwNGQpPT++kvpVsrQokovQ+hGQPK
TJbS7F1YhNgUcdTJw+DtZSRvKQkqLyIEkP17UwV42mC+yvlWzcpKFIHzEJL8PAov
ULKfK6mbtAJFxfjaGW28bIpqq3hIwDPsSYwQwXtDfwrosTpXCKgttWS0UrUzc2FT
kI0OobTxwHid6pixZaiG5JQAXDm3sGMYQ8/01T3/w6eii5ysD6qNc6K+irkOWj3U
7Lon3YKT9xVF0BDfZqz1uLB9bKz0U2VEPmN8Npzlf/BIEJL6mBk4hN5rzSZvEAeJ
oyWwLlxyYDJIdU3qVxaVhQA8FbJ+F0oP/vHVe+U150mHraB+NON1Afl32JXpUY35
ocp4kvTMReiyzFrC7cuFq/QETaIUJ0S2nHT4oJKa4XYO7g894L+xM9XMtBKA16SS
L7JouQgJWlB2bPKfTDZWMGDwAw01pJgjqG8K4t2uO6E4In/BAul3i/77SwciDszY
grtF9kpSy1+YrhLO1NJ3yz4T99dhfWJu95B13EFYU47mY42RE0klU8ZFRP4S4c+u
Xm37avipCxdg1/uRG4p1WfCMNV1ZUNKcxUyB1HMx38jdXQFEvVgNrn7KBZYVoZGo
yjNmjIZzY3QwRNgGsrYauFBqdQv/cGNu0YmTU4yeOVGVtkR3nxfqP51sTszgvjVV
mF7GdCnaeMatxoZtBJhTNtCGTAKoRlg5mwCXow1a3K+ZTyJ6whgykpjYAan9+Nhc
sDuNUM2PLhmfp9mfeDQK6DfHDMZmNrHqnYVa2hTwfvOaU3MvNarBym1vFbRk4ezD
x0/3rsGt7qMeaQ8rXoHYw5HXd9UtE9fr38D12CKmHXE9nUxB8rxUsTCbtbSzPsmy
kbiNHebakdhHDSevcQ/R+/YX6fwN+Qb2pDeBetSvzjdbUGnxgYk7wz6E1WxXsHtn
LdW0B6gYg9TIDPR8ILKVffXZSAb1jrCp5QatAgVzcs/EA7wKJuOzaHkMsPrKV//M
2xqx6VRmVgIpZakS5MBMg3NFvVgqHGfZIVBzM8a7kWxcSDJ/EG25MLHYeVSDVEsF
xq1U0RENbcirWLSvuhFG5lBjEbi+FyvOcsVUnSi6Zob+XNVlLLbWUnkSCRaCr1Z5
qXl+plLJ7N3VXFWxtttL1WYy1j8w2gF6eBM0spBasR11eVgYV7fBO0JNG3gzulQ6
LPpvvm+VZ4Ucq25X8U8TLSp2FO6L5zCmBXnLU95JwzAwKahCbKKNxzTHP8wjE0O8
6/UhWRkRUwtTm2x51Oyk/ZiXZqmWCZv8IM/t9K8Z6NERIhZbaxeTtsUy0tqWyKZE
7j9kKJZTwCx/csemLVX2TLOTNF6PdpBmIduXm6hGy+KkUsl/KpJPEpUhCIluKe7I
m2YdHZiEZys8oFvRuO8SthcoNW2HtIzxvNlYTDgM2doW3g9/Ni4lmwtcu58NRR46
ELI9JlE1xouMRl40xNDZj4xR7sR/3sKNp5+s8sm8P0BZkv5bGgRBp9J65Ww0Z08F
ovQBBR5Me/f/XEouwP2WJKS8EiGNtLUT//XqjIcf/AvgAfWvdFMxqK5eWaoj7YPC
JUyfw4LdIvvT5LphxHwNNSFr8DWK39bRjHmSDqNEFdu14jI0PdEOPfcjfDXGdWJL
Ah4mkFYpccv73V9ECriEseOYRyhdeG/w7MDZUEIlefInGNROKegGveWNWSHbuhQT
t6j+5gGVmRsUoGyfYpmwNwQsKxeWq0jm7xrpzD/xejnigexqlOkjDyKh5BDQE2Ff
M0rLsGzaE98EgFsY+s8YKCfQgEKvMp/2ZZBNCRw98+pxQvXRlcJEXF7q7AM19yOu
33vfEIarfNlHqNBHVibf4qNE5N4s1QIzecGj2ELzii0I4Ug7KBEDbu1kKVTO5v2R
TkZEzNA2GJT+r6KF9D/PizYKh5ctB+UPS7i+Dp0Bqo77Dt4lYljG/YxC2tqu7DpP
xZL45l580uW4JLbC4bYsOhrtRr/jQ7kHfihw4Z2hpFZZpPgSAY0e7+cq+kqpJsoK
Xk5OTiVKZnAvtlXkxM/3R7I4EOSDJE+klWyAABWpb9HiMntjpsboXCec8rKW3p3r
4UOcpBimCVqsQuvUo1mGv1v5OXpvMKaowXe1gtVbySmhn98butoQ0CMGApUDsrOf
qwii4YlA7XAOzLzdR0VRZovjdSs6BIJT98XxdDdNmJvQ52X3yce9BJOi0WAgJmFr
C1ZoqyUbFHsHJ28VzvGgXU81l8JDfJZ5/hln4uasrnkGn3iCX2/byAN+/RQaiZXl
GkrMJayz3L+JKdz6jmGhxCbH+xx0FEr22wmJJaz2JcrVksn7d+zWYlx2wBxosOQF
NabZ2ROqQ2YOrhNHI20tRlXt6B02xG8fYsvFpqN9P5GlEIeLGV4qfcDVhtBVT1EJ
AwzAWHL00KMQ3zEqoxCyuZ0ZKVVWfyp7YLvGCE0WUmkEzG6bn+xs+nzr8mNkdAKb
VySUXAwCcK+xgZ8YlUvutm2uxYgxWXZJyMgnTJo3cwyS7IgzyHu3+P9BvbRfDuuU
Auqm/fCd4hMuGz9z/XWJ0R4PyxfSiqAxs85Cw5CgK+UDeIFUE57THN2nnWucDDhW
VFUruhGI5G+z1oPiWOJhY6Y8FtMpBFjerC6AC8LWDemwjTRXFAHxCYhf45TGAzsC
ySUnB2SoFJVuhDpl3DClGUCsDf22krJtdzGXL70EFE8LSqGh5YjUoZTQ8ZsZBZBx
Uq8L3eg3v/YB8/0+ADPro3orBNkhv3lP1qGjpmMPh0kZ/DIdv6av5+bmcJK6i1d8
eI1PKaoYKPWaJDwjMBNp/awu9NZ/+RIqNbjXgqiaqsNAw8eC+t4z3gxAhapoUVgX
YqbBIm65efGsvBNPKAgCKS7kT7TEWsQTMWSrFztFsY/xz7q5X0L7LJhqD+0p+85P
rwRcCbNS4UtJQXrcqxJdDeIqAUYih4R7hwocN8kqGE3NAavyFN3v6wpGd9ttU2vG
djLrvY+Rub3TvHQ2Iq/0wMkUR92dyTu0YWJQHa9cRTPSdemq0ku8To++ZF882nls
YnBpN1HTwgVm6Vr2wVo/hfmxOZ+sg9tu6S2Z0usf8S8DefR+Jc6MICHDNJvH1FCf
ziwc5tMEVNp+uhiR9Ak8PV8JiYm8NsRyzVneKeA4ejeWEmbwCm76MmgITv9Gte0J
D1jwoXz351l8usu52jgzsEuNlOIrx0EB7vyVkBRjyGvmSznRl82uWprImP2sJGGA
JgTpK+2Lo8on2LEu8XsxMHaue7RFp7kGanR3dDDls6JjqsrDWGwKszPTj/ukG90c
m35C0lC1MkSjSvlpMz1B3wS+q4De5av0saPbG8jc3WMR5aKNVCO7Ava1vMguVa/Y
4sPEyr5atPRBcc81oaSkhJ+m99vYqG6SvHmvGmDzOMFzqTjA+acpbzHp3qPN0x27
Hpr940y8cfqRowI+QfNm/UaYP/vY8krkhu003JTjSayJ7Isp56dOPIgaNTFXaArz
z5nWMZgg+If5IDTd3mnz2YqlwnlcJDlLg4WuoDofbPafRh346ZHCCcTvFpPH+Q7P
8+8Iu4H4IrgR4tEIj43PpN2wxNNoIIjPHn8B57Spci12l6q99lXxB/jRQPS6xBRC
Oj9WZmrVpxcGTrsd1XDcI0IZhzI86iGd/nLyShzx9tdr9H5vGOMpU+QxmKziJw3O
RGORriBWUEWX3Iva2wjNwKTaqmbPjBnLxQo2v6gAtKnSbmjbqKbNU/IZVN1RpRQP
wIcAYjAnz6QFfl46GPnCuFkETekYkIKdeNZ57sIVKXVxmGu4lXC8EC80Xygk8M/m
UhCTrOhWBOpaaMsXWqSlILglC2YqRYeg2ZuZq5q11v7Ws9tUP96qmbI6lS/vR4JB
/ynx7vJNJQazD2cYM96tTMeHlFwhgXVDhi8WZ+t7dF1qYeafRGhc35/q25HcG/OR
tuVjE8izsSbxO3dIpuPwYyqDlXABmlH6hOhIcGrgpldVCl4jpYsUuav0S6MK7ke1
n6QdZf6sHBfbcYpGvFuB8YQxzj48VL40Ytpk9GTB07Cf9mybwXVbulluuY8tLstH
iC5SfB1INGLFPkLaq/9R1DPBk2P+2VpNsZ/sk7T9wZ/DMcbaoIDKbJffAcVj+wdI
+e/cDXoPCl3pa0JsFj9UOpKeTQyboA2SZiVuh3sT5nBeUyofN68ObaCKtjI7UmnG
SzmilVH/crxvOGDEyEqVnOKGZmO3GDQn84J986pu6nMiD8V2OZ7WkafEzFoRne7v
w/yLjxGicf1slk2Et1xjrt/kH011HlLNguVcPFfnpHEth81UbVArp/oR9VZxemIf
ea6HVh+FmHlDnDlXaUe4piu4LP3M0ldgTXRtYQslQSgk+GlReY4BzI+/7foZqNgs
A3LOnRlxhuGRO6lGtoaVxQpgtSOWkljHS1reLcF+QILLLkObyMUh4G0297ZaiKuT
SrQMc3Wt8PB3YAzMx7zTseFMx8zHguX/PVe6//CuGRjEXTHT4jJpc7+GbgJ4Idce
rmxZUOEJM/hSGvWKc6kl9rpLloV4bMtSCA0ZGNB3HwxULK8RY7ezA1zZJ++fCbAw
6/IJGJUKoIl5fVx3lgldgnJYumLIepJL53dGxI4kCVwDoCRs19mKTfaSbEdsukUJ
whm4v8m6nV24u13MFU/n9gvfoJWIMzgRkn2+CAQCcipkmnyXOweNXH6q9U0EyVK1
9N1JsWxuDi7E6nIMbaTVqWEIoMpP6V0DYCroDWHB745SYvq+SnEZ6/csiuwtDCz9
YPAK8NwL1kJFcjMsG7HsPQnp2hwIaJMNIBwmB4Fag3ACttaY83sW4G5tbuNvmy1Y
B2ly9+PhKqpIh4sNSOUZGBq3ys9TCeYNyahbA8auGIGYewJs+mRKpq8CsUdiAKu1
bOnWgZW0tO1m9GzGTkOppeL+bJwIucgMwOKh8B1Ao3beZqHmbjEk1EiOCxVYEppg
7GvWtLErUVv5ED9YSjwwtmLN3RWAKL8FfOC1G7p4MP5jxtCR5AN8Dd0IPCuhUr4O
DtKMUvHK3sZ31a/l4nalIwg3kQreXwD8dgQZE3YBE5orT3Nez8xem6/1hWf9no4T
UEqdsX4vi/FMMU3c0q30KQ2GoUhKK5XPbKqpPNDUM1Kvecl4oHnk0SUynSJuYvU9
uBFvCdKP4h3mGL/Pn0h8Wi9d4tuysbuNM2KKeibzxFQqxayJSKVfMnALr63yhnaV
dXyXWakkGUsUREAUmXOZKOj8nsOdT4P/vDf1AyYrnVOmwWYuP1hAzyegFdeARmvG
Fcfi5iYtuwMuTMFhmMmcDkbsfnipvGsdNI/8puW/rewK3Ds9JzrBb63TlEHy7Y+c
5GedLw3xwtfGaGR69XDBave5Dqcy8YpKOtKMcqQ4FFWmFBZiI5o+p1Ja62haGvFJ
YGU/I6L7jS3GYoo9E/ZJcBMOUx9d4zt//SUEvgsUSGbBbLY4YT2Kf3s9W8p6y7GL
W5ZlymHqAxkXsoTI+mIIrxC7JlrHr6ROzChxDUYjZVhDsDSDP4WNUBkV6eXTD5cZ
OoS5QN4PI2P/OY2UmSlhsgbcpvVkPqII2aJXs/RyZZYYgBNW9fjYMt3Xhoe8ZMqH
ufkn9zB4oqC1C4DrtchrOsCsiq0Lqv0y287Irg4pdKUXj0mPsOzT8JD9qTvU5Xrp
9lV5v1AzPOThiL1cJho93AUiEhFYbHHtwWGbYm5l3KqMzLsDhDdv6kD1BusPAII7
Rg1BK+cfLwryjFTU74MynmRVYUUyHUK1prh6rpkuftpqOAvxi0ZEJAA3DiGHigOG
I+bd51EOVAFpes6bid1gpoQTBRi5DlzmHu/0FOszx3GZ/9IKEcuKS4qi9J/aD5Ao
cugdt3v0JLb2Ypv+7N2YcLNZgHfAW23RmEfDfaIT0QZTySts/z7L1Vmh8jgjhQDc
T/we/4Hm2NosOJcRLqXq/j/aKQBcHgSgGZhboyYEKT/1JrrrMqsh5nIGaOBep189
kq4EkRJZcnyLhwq5LCEfiqqFC1TwuSeNTIguJklSjaqYjuhbiG1WLJyL5qtMLQ/U
VantauLA8aCCJuWy/MQO0zg3RqWn2M7oVKRKm7EEemZTRa/L8xDGVJCQhFbOhiCQ
15u0HhqV7lH12vI+jrzDDgDK+gN8n9Cq/8z0EJhqHt1GWSK4Oh6OgUYQ3oUh9dE8
qiq4IBQyXFAut4pLeeXSf5oY2scpIH6pifgAlUf0R5NnZxRnikvl4ohoJuIJcIPm
DttOZlKSMy13gtdvpP7NYE4YhOu+Gmq7B7hA1O0tDsR+ljdD4Dy9h0/gqKvyIpyp
f8ENqjjocMn50OiZs4ZIXHpHUkHVjYyYZmB9gbMmmjBBfgz/ZEZ0Z4Q11xVSZMsh
pHXUDQ135PIRCPYwGrVtu1ofAcKbhsmIQpcxf+thkf0pu/P0YmnJUJvwIJbCJQgG
M4BVx3eNSuHBBH0PTj7ppEtZn25QiyGY3xp+bkOHbfR3MtKbaIE0NBfIjsfMguL+
m3kni9zmOfBFU438FsTsLvyzH3bvI+LJnuix8iITPgrXMd6fYhlr60VLnU/YbtEu
I78IGSLC217kozixJGnn5bwWSoZ42TPfg9vlyVF2r75sUM92f2zFKaC02/hwO0JL
rzMI9LqXOf6BztXnKVCMou0+xiFZjqa8xMZ+SC9x6ACoLzxhLrL4EXCmyJLTr6Vi
gv7jPsQPZUs0qaeyLvCEG3RQpe11d9w97fAJLiRBvegjGQ8D+bxtwtpgZKgJgofG
SWd7VtUBpE9L2qqb/sPZg9SbcYnx5fkC6jn8H+A0yI0T4V9tRYx9pshLhmZr+2fT
6+Fjv8EF+Egw5yJKLWO0GHoTPb/xMhS/JcmQotsoSWJir+5Eh653zOYGSvaTyL9O
fa2GxdoYtzAieTkSnry7jSDvcWqqbYr0XWbBWCTDdkec0MjMFYjqALn9Eb8AdUl2
mqV44yUwQ/bxp2QDHrvYbYbupCMx/9EZEu61HXaUQNXVwFDGMWaLMhxfZHvzZEZy
7B+9ugT+wuPz+LKq7hOCNKTGX5/LutTWfcm9zWTuMp/A08CIH3m/CW/T3yg1K/2a
WuouTec1T/s4JXZ7DZawVPVB0t3c9iGZBRgJYo/xPtA4Z595drZURq33DKiRignM
k60L0vM6Oe508VvOaZY7+L3ce4g7IU/5QsydgYU9LYSCofjYdmB08a9pU7rjIkeP
HRNVY2JCxRcyys4yPO0+I39byvSq0IaNYd8M7bpnQyfxMzv9H+zTRnr63zq78B6f
+w1XMO1wb8tN5wgKgOi/oD21X2Df4A8/3P6PwwUbjZIlA6rxj18imyTCQqQNMb0B
FWQCFdwqR/gNY5Xr6ns6t7+j8AEXSSV0Mq9myAoJujjAviW4iCOuabs9KjSviCBA
dFe2vrrGQWyemL9HInUVXn8+kZ+mWAY4VCJvzqNM0EP6YhfZyfJDfibXmaRBV4d6
yT1OUDMyNv/XkUxaVKNLJ4zcOXqlh6fFJdwmXgMDolP2S/tYW/gdD7w2C+3Ly+Yx
ZZnmbOieT0nxu2dJJd6OodFwI2oc8hLSrwvADI5mwI8iUYajpxi+xt+iw0l9E80s
nlG+Son9poZIIrVBH/kavFLpronfEdhiPKEbBYjxdG5tY75zWJ6mumif4+0yywZr
azj3tQplBBzcw5FjsMvO1/amlGB4o+t6xJ4vIirL5LwX9ES4rzzOf+YDkQUFCFfy
Tzs1EfWxYACGRMzG42MHoiarDpy3a4lBiu0a+gUI0ePRm4k0NIcOEtGnLl6bVpvh
XYT+ZmLq7In6J4gkGWMbED+L6FsQ1J7NwD6hK0wd6O001ZbzEsSjqmI9IOmtdzHu
WazsmzNPR39zXCNRq2ZoXGqZAJovdqt3L6CsOQ1VJnsK/gPwSzQtX5MFIlWQaXlm
4+4i6YmI+HWVPuR+B2HGD+i8sRdNZXGstq+oIVHUwDouFzIDfUaoTV0YdH4JphX8
mAif8baA8pHSpPwZPkmlhzj74T/0XTXTVDGQYVYeLp1hulCA+rLChL3Fp8Q2HQ85
bZhLG+hyBvlvu4SOzn1C6XYj3/BlPW9D/wDK2RDgcWQn78oRH2Pjdw0rHDsdmX+3
vOg34MjsExaSTh0DJcWIlhTrnvryz2tdl5d/dgrd2a7787BcTkqqYWJNmm5nOwI3
0gw+dhQ1Nq2UHA/vwl9/5dai9bHnyxN2t8akPstCvMAwJyJvjgcGxFJ2o0XOFjI+
6WGKJpuYV2VLFPlUDzSVnJOYNcn3Ras80OArTja5xXf66ieLBmYIQoPkdDiWOUSw
6RIJ6fJiUyEYMAwpBiAAYVzM5mDBb2wpOGrR/CUzpxh5PkSbTWpvVOn08BBbhzIv
ahARkEDjBCc5+o8cMP6zs0h4nOiWqS27nKSxD/n9dJ+qEWPPXQSA3m56Erpj8m6s
BTIQ2meFAkdpU2u2SzZhpFeYJRdJtUXbiOhEY5LytFv2oavKrIWGFIqZjj3mnC79
nMmEuWaaZk16EYKSp+XLgY7N8FpODsCPgjJnGtvbIHkiDI6WG2LP1bTXn9UG4tmO
v6s1m/0yjD54Ln0JcXCsV/8uyqNbfSku1PlO3tyIg3Y8Q4SSVL115fumW1Kd3KbR
lDXJtdr7HAtN7gwLHQ/dN+N3Lyfop3HB7kfCAvVWPlZiI3YfUgX4h90uoEHKgpAS
6uEL62m7iKwBAi57T8kqezfapSdnR8e0hl81N1CU2Xi9SW3Thh+YdRAiMqRhJJey
YtuzUpFln2a6k2avdPlDv/GILpEQ5sQM0ZOJWQDsrpY4WOA220SxdpVtb+Bz1w62
nap2nsgwHCd984YK+YtrAeUPWLDObLtHe+mKUlYzIhRISzy0DWwwq9m/LOrrLmc4
DdvsPsDekIQf1LU64XXdJNXFyJ0t1xuCS8u/eh8Hal1DWvTSsNrr1hXy2WC+u6CO
QrPSOD2Il8LURW64xTcv/Ohk26+Insnj5qifTWUl6jSD6uwrpR7zD/WCuNW4kYUG
seLstMFfsTHhx2yb5cVGAY2WSFOCjWf28H9TDugQvXsinvQj6sy7IV33DOPbmJLG
VwdwkCIUCSWmpfp/mi58ocGaaFkmWINMm5u7yD48pM9cna+aE6nfx3bqeeahfFAz
4IhG0FAqzQcvKCr7tLnxIhZJpf8fh6j3PFqL4pC/ccFEK50Q0IcP9P5zkOUnh8Lr
FV0718xa6I6KSzJ3/flJWVNYmleZjyK/DY6+/sOSx7q7XTq3tZTY9ExoEd32BGH6
qG7FVi1v0mUmKOUzo57mVmfJUFFyJ3ICkFYqONiAygXIxucWi+4Wssu7pcqWVppt
77Jx4ikjDqVJJb0ysEPHyu0BwE9K/79ZixcvHYYzM9inaAvQEJteovPq7zcBgl27
WE+8vBxRabUv3+rIYnm3IwUYkTKjCinZxipQ6C6NSweSOPgkbYXOEaQetmygRH0W
x4zAehm5B5ugXemi+N+cdYyMHmzFEURw64BugVLIAb2D/pBsmbJ5npGJSQozQvmX
n7Y72M7lE2DLivNqMb5gEM9aIWGfMkdYTrADv7If0kluN1G4vawjFjWIC3nWHnt/
bcNLbeRXRyM2fPg57UsqNphwe6qYjT0D7h4NRdFQSZG0wd9M4o7Fx8QW7jyL/CDA
G93dK7R7zaC1dAH/tUBK/hi5ptjFRZuyW6GqK74617qo4faqBRBdi//zOt8bwLUE
LI2ekMp3WZlaf338qdZVHylbPVJuj0R6iMi69tnBU0D7p7Wj6EIOlyv7oW+94sRP
8gP1Jb+J9Y1bgYL1z6It/i4xE4QPwOFvAYRj1HXE52H91TSckqqSqmr9OCZsK8AQ
+k9XwgeKERKyQf4NjbKPqWCcqCazo88vs5zTdCiilUqfym5weTgUWMeEs2dWyOWj
bAZZo6IwmfEO32jODPwrMLWeJ88OyTow461xHENS3Z2Ii6W/e+xgYCzOrQCaeCs4
QVnhMNRpJVO6ciq2hW6UEAhBFsrHROH0FfEAUm2ViAG9EUxC9vraPXREnK//rjDo
5jzQpZKJud36grxnHR/JIijdV5NThHPXUweHkEFAt+KTMTt1aXfS3D7rfFfaAqL/
iAwgfkAXz3r5rEoLA3iKnS/e4JiK45i5J/PgNkJ61dYP43McxvjPOdCw4hBFDMgT
6slx+wFPAfUer4OVxRF+w00Uy7VdvyhmfC3Ag65B6IYABZ2qRcr1QT1HtbrRca3j
4j3sjd7ZBe9UVkqvqNnoN9iy4u/RXbgeb2dZA7R8oVlkYvYRQaioXIS4t1+4LN0P
T9yIjKgI+ZwvFgcS5t8cauOKE1yEA9S0hESkCmaJ1Q6MuRBcMA3VuEzj3t1kLXRd
IXiL0xssQxDcaSIqMEfmmLhxCPBh9uF6phDSihHM4goofpR2G9GG9kQZ6ff8hcDd
CqyVh7S/GNxcTsabfXaPTM9euGVqG5GNapXBpq4omx/YsL4RqVv9y4ctKk2H4Vs0
WlfnB0KbQ2LqIPpakYF1B3VxENpOVvievvOxHEgYoeZnFPWMtjgtO+ZpYf82rd81
VwYfzkyl1YXKdLUIOR/rNRELPqcJL4oWROhncSB/Ioiow12u6yMcI9exFSLwH9X4
pOQzkkNQaXnxXtY7kH/oUw/lzTYO8BhtrQ5q0QnA426YeRBq9La1eBp+lxauRoCw
1Tw6z20N5r37AHkkHuVEL75KgXepdBhn19VPw0Yw1gte31rr7fDGGp8oi9jlIk2Y
7QxeGCGcmtdh+8FlKoDzaphwjZXlkqEQvrvrki6/MKnBXF78otvLItyHpUJxen1O
Pjh4XYn8d33ryPDGG66LAweArPzaf9jxI/BLitwIpxwBcLPaws7c+Dctn2ojUF5u
iX/VNcdoVytXGg2l3fcRO4v66nPtObHYGv2rt8FRae9UMDQs81dxLpR6qO2wyX80
SlsUi9IBOipL/tzDLNi7vbbamVKhWw5JXFLyWpFLoMt9pn8t/IEe3p9XhEpVH39m
0546ThUahijQH6obkDdyM06d1TRuuluLWQpEqyW/9+nrvRnw22BjpP+4w36jSnGE
umlyujt16W5GnLcQylA9yzqqw/6EBDFZDzMsMoDb69b9aId8rQuGSVlhP+qTiRAC
QX40IhcQ4dzxAv89NxIl9vPE8se5X0JlGQdUjTn03SCq9bLF03i7txjPQURiHXcA
dDhbZtM6YtaaNXeCOb3xgxbhNX1Aq7bBwpnfNY61q2uopMyeib6+QM8nT9o70TWw
xafe40hovbprbyjdU3mn6nPlnKJJYUglIU6VmbHYopdmx7rUx/y9FkJfR/DYSPtV
EbqOSvfNUfTvX2I1rR1JpoYMZGScY6qqefhke+uiX/2niBNWWOkQp3zSio3TZ0ZG
/q4olGK4Q+qxy/ZHPHYZqWUJBXulU2wZAFps+prZ0K1qT8kaL9y+lUBscxWIKGR/
na/sB27tu0fscxgZifgV3uZ2oTtSAc54NYkxVKOr8AR4iq1mBxX7SIHaduTqTNUl
ZndBfbifL1U8J7hFTP+Hsr0IINRkfK/r2kFKF2LCaEeB48HWrudkziuMbVcxeqAL
LGX2uA5ktiXsjprAkppK+zpypt1eejfjPXJ929gatYhQFDbxnjjkV1hDDPckNY4e
hhUvq1I/gZUn+bPDM4vsy4Z9PPOMWNreKfpmHEMn4Q+oyDAbUTbdJFNhfYmG2Pky
XBQxS3XchVkKxrJrsl6c0feXN6QsF4wu088pNizpjDViMF4I2YNmmUnL2y+4BMQk
kQgvnU1f5cn1NDBXfU/vsKIG4vTcsgBsjZNUDRpkZrywjWLl1n6Gvmf8w0pHoa2f
g/3zz22se1M8/SqjyvvmUK+FbrbyAt/bjr7gxs++ozPIhe2ZRS/DI54WQ/WScRS+
6IDZFyNAS2MqQpbUgMdtY46SiMFH3y4Iv7y9JGbGl9/aLE9EAyD25zWY9zi1NEnv
yBl4Ug63EEq7uO9XIcXAuy0KKjUyEjvtlKNKJK5eLrADZgOc28KwHEWBZiEM0nw5
tgupWlQerPbdL6XpVyV1a33XfSyDQ4ddNxpTIQKcRxx/KfbufvtbPXnFkUyb212p
B+nud098Qpkb+bossykth2pFWECoj4nkAcmOCu4q2cpd34tejy5LZTcied6zyZZD
aEzFl8MVdtd1QiGHKnBzo7lPhpiOBe4xl5YDVl5M82NFpAaMAJ/Tns/CVEKJiw/Q
usFmXbNrmINf9PnRiceW9Uw2G3PIQTDiVKgtat0lSAtLaJuLxRxOrv4oDKlhInTY
JwxKiTlpKRMEjwWPKj4DIJDQY6/jAycXwbCCwiy4HmxJaMpKiEtFixtyLpZbO5X5
oC57xU5td/DH0VCT70yi4c8OyEOgWZTF3kIiHOx8WPnLlFoVdmJrUk+hLDwULvWZ
ZQjn651rwJoF5qE/KyGNCE4I14diwufK0fKcek/CT6VvjB+obGQIO2l44r8biZuH
Ze6Y/4msqHQk1nc4PYXr6t5tFtYPaCWneGLJ3QEt45s+DLZJHtvcI/7phFUtuWaR
LgBIyTN637IVnhrgwwtdUhpnBlYfpkEgMm+LuEucvgoXbKKpTuCg5qpLmwZo1YAF
Axeczi/tQ7Ph6CElhMq4CUgl+upkiYBU9I/28iCoJJtYjYIwiHMlANokynrmW0zZ
Fq+aMCwpRiD8dpvafRhh1HyPjIgK/ohZZfq0LOGwvhAe6pTZdTilPcxqzm5Hhriv
esIObhZ+7qoWKoa004itceH1itcpQhWxXb6E+rVMjpyaVXYg1cHXBdlt2WGixvzE
A5rZPlOgbcYKmpI3CdtHUtXf7HuFzM8K6iyYsUXslPibEgS1M2Soniyjhe4pYwXf
7ssHTJeW6IQZOd0TLdLaJEJ4F2+SG0kVeQJDIcmdp8fFZeN2hVFEPT9lec0/edkP
zURTWKAFRYYBR1IzpbUV10Ukp9f/jMDqIc6VO97rjT5jfPNR5XxsH86UTCfxIBWc
Gkn0hNVvm2XbEYI6yuPHHislugS9eIj6fdkZ+U9ncC8qQK1dIA/BoFdX6y2D+qaf
igMwFRrlJBItGZCnJwEpQNaCO3PU+7SMxsSPGZ3eon6evNoVcVdyzf8r+J2vOMOf
xeegV8zQqs9ujQefdmV/E9tWCWQgOGiYvwG4YPSC1tRqtTAQdY4NgCcJ5SIe7WAj
bIxG26uZdvQeTl0R3OVK2J9zEq2W06M4ULtKRrTjngEpcHZ9Pnsz4lbtSfBUxXqV
SMdjkKIEqg1lt2K1iwO1a1E/cIzyTPSiWanhYO0M2/UUUDbW5Yza/6zlEYZIi72p
aUPCQhOC2V0KHKQ7Nfbex8JelkORO78b5uQgz6Ihw0NjcwQzqQ/E5OCZxt5cn/uO
fW/SvAFrXEyognAVyA1d9HQ0dffeKhrD4l8OBuynVyssuqUI4qpl+p2wDp/929vw
YLXiAsusq/o37Fb9MDB2vbhPGS0M5PBv5RCDMmv+Xid70AUeXbOuJXtS7bF6ZSCq
G3BNy2G09s67KKcf/LXOOsl19r4IH15/CxLHggttS4JVCnYrJNt8kinPHZjkJVEB
iMZHp14I1QE1m9BQ+PqaN6CzMuty+i+12rDkFx5VLufL4FAONdiYSlWt8LBcdj0h
Ri3GDWG2jj9wT+3vMbH+h5NbAvaMO9BG0+fRMsMutO3quneTjSBzWK093wvHpSa9
byVIMc3zu9I04m7jko5j/Sq8ktfFnN5fOZEmDo8ZCPUPv36y0iNehNBvRKV4Yn68
EsAQUgh+NGIHX2N0TeZTQCX3LgepRYR2/clLVVfycFKSIVknjzNRcg3WJaCq1y7l
VkjerUrgpCKjZqxaCZMB1tVIEO2epbJHHYW2J4RurYKu7VITRnq28CcpkKVDNc/m
XIkLXDc5HyyP28/If7/Nh/eExKZqUL4BGaWdJuEFeGFxApZSA1adxC009iCSWLVH
os1DMxI58CrQTNIhpYubwDef+Wx6C68Vj7PatQcP3Ot39XFvsfkp6yD3EP5mkNPz
gy4JLst4fwcZujNG+VYB8+34qjgNE1TWq/T+iTCwomenw1I6/Ybctg2OKg2cxfO9
NDkxoAuNVM40fnnS64xZWss0SYnCsUvmWlZZLRg+CJBj2Jl6epaVwbZjD1HIeJH9
q47qTpJRW27w27mu4zpBvVWDm8hOhahGoZeFVFhI4Zfelel6JGTWssDrAysMFtWr
bk83mts66FW8mEAbPWW1La/m0FOU473PLi9SilhLiIRoiwUg2lh8Ixj+FPX2S/yr
/Su8l9pb/jqEnavLjIGw8CupWOambTQR2AS7coc7SgvmDDhs5J8uz4MAwwa6nG8U
YUz4Cd3/ZVhkdHgMxE4aykq6mr0hRIiXVJkhYkijMqu/VaVmdnX3V4AkFuBbysZL
aZ4lUqceOUf9rvvu10JNsTYg/Mu4LQzARk4x1UsI1lCsLMNbX0XXGx3JxRM6iwv3
dphaCpmB91+0HgIhCykFH1iU1nbcW4V6yYpURw590ZjsJCHNptxh9L+s83j5Rkge
nri0JWfHX3s9ZYAO2IY1sOcfm6TjBR0Iaop4ImLG4i6ADFMTMXtWue0cyE4OUapn
2d+u9B6R69cNl4l/8e1L4BdjpllVx4fKrdQaafhtv0kpjrISxCPICXY2pdAKGMXP
chiT2PZ6SFXFNQomxwxIB6WY16dtQ7+lF0+zr7gZSilpWKZlGRJRaAQ3rbJlLmRJ
OQcwwLDYI6BQs7rgc03rMyw33AjiwZwGO+uxNli33Yt6wVwTcLI/Xef9jJUmnkwC
WIUx4CIfJBclHenyC6YT1Sf16rnea+A/rHOARX5vA3jhsPAwM2p0mhyq3qmMY/Af
8y9fZOo6M5XtC0FCzVxnnfSFEXVof0yQS9n+57uIEvNYCR1IudYx8G8Cj834KJzj
qkYvhnGNr8XlQchCVZAShyaAw8J6WQhU1q6kexajsGYRbQ8I7s+W604bNu8KH1YA
Ep/HIRiGR9uUZ6GUg6csAFYikF9lYitju53AEyR6Y8yvkz8bgVBTWN5a1Hltts2W
TACo6+0q3HsLwfHFfgJoiOkFS/8c9m6Yqnv4rv6JA9X65Q1SOhigOtLK+fK6dKml
PXEH+Szh8ibjLCusshCZJm58u+YDyBclz23bTQ1hLP0mh+UQW/mW7GYqoO8Pr73i
z5Zn2QddY7tHPqSe86DfjevNwRJ/Fn1V9aiUum7vFe81dGUKnrR+Vi0C8E/4VG6v
z9NmSUi4IURK5P9IPKQO+EB/h5ngTkJ6NbFKNMnrrdUReY7ye7buRUiTPdVx3e6d
vl7DY5qtf8vVH+3XF6SwTjRkmJJESNXKYddTmK6UhS4UkEJK6cUuGYlk9aVRO0/X
8dIM/r932MuC1iYh+2N8S2Mon2FKK0ccFgbSiGmB4ErJT35BSDVcR1Q4lFXgwCCQ
1QvNEUOMGBg/Ys6jmupYtCSlvHA4J6qva222ktSmc+nqm7jF5qDI/UXU9XfCDD7c
mIpoED6OtPTX5f+4AoRWV3eFaQ58SnS+7BBMYEdDh67/3k9ugK98ua4icrwqoQKP
ItM5NGT7e56asZnOkZVZ1m8+v7JSMON+xpMfERYNi7xkRFKPvFofxmBDjisqviRA
3H3ce1yY9zy/d1cPaPsuQ/OvGbCUmn34kh5C4XXgajnvntLKuDIyS3Q1r0dvCoQQ
QW2d8WoHViDyBNCywik+5YJ3d48IEGH2FL7+pAl76x3c2fHZ0ycI/49gfXkpVyS1
PiPM64eJDzZbbGn0AAkwjjamFZEdAO4HQn5EZHdbyTwvI602+UQlXTU9JQpGGNVA
VGjzKjeUZ5zGfK2wIo3Ihs8xExceAifO9K8FWgAu3A7yDhqUQyfm/pFXLfFWpoRE
Pvh8wQTgEjDjrXWpxv7rkQV6YOuYKl91XFmnJ3ABAppyrAXnYdklsA8DzZPoEm+X
2TvZOxmqk0vXhii8MPuaMKpPIBD/1a/JcishyLslz0jgjHNuRgkOEBuDvFZcZZLd
fszIp890vMYMTxtWprBk1U7PhzuccF7OKEB07qIGcxbOPPABt36LR5DW/QyxVzGg
8T07Jj5xzcDQZ3jMX0YoLj06lJfPXMFEdG9GZQrHrgtGD3pIVYn/4MCpAdmlpsN0
ywXGUgHme1ozHg+mSvC+7JqUDjh/HJj4cuKq135WfAMdk9VEcF2ExUdTD0d8QRTa
4WfwZmtoj86pRaIlvLBlpkdOkCSbu516NzsmS30iOIKC1XFG2EG6YtvNb9BoIP4s
W5+i6/h+cWi/V8pfA1qAgyb1R/nJHKi57IBPqwutsC0v3Q9rNMwjTkIAsUgi3zKB
u5tpVo1g8pmqLpBeUyrpm3Snz/v/+CHoHskpNaNlbFtRd2iUCj9zEk+qokF9MUnU
90wpyZut8cVudVnOWWXllh9S4b3Mrw9JpClWno0zUN20B6OkybebLB8Fezi7bMU3
Bv5P+/xh7cN7eLnIR5HxY5IUNwCnHiOY8U61MmnQprrPiGWkhQynJhCln/uAsTr/
nIcGBumPWBcxy44mkbZn5CHKLs5puZx9fYalsooaTaS+unvqipMjsPtmQTvMJYUh
kkbqFnE++dcObqdxRW07FX9ZIBH19RUFMcnziBRgAVK25girFi182kToO6kHI4Bq
BA82/+B200RH4YiyhAn0bXAbgKD++vqVZJBVDgWA2vSz53k97Uu9L8aHU+VDPq2p
6fQcrFYogYoXDJGzELjnZtHcnQKZJMUlDqE/LBKblZ833j3UaDoq58lCfEg9u666
35qA5BD+8KX8XwSrCbV+HVegbHWadXCWa6afKth3mevzFpL8Apgk+5XjaDsrd0CL
Pu4ufsJfVXns7r5ja1/EDEiNg5lbO6Vyf6ZoLvBy8NuZHbaDXxCNayfGoNw78srM
fIMjVTg3RERT+4KIaOw8dGylzsDJ64ZTqAI72IIGDbz6/wCvQGd9/+LWenyN+4lK
G7Ptx59T4p6vpGkL+1sf/RrlEi62TyNNA3ooMTl8cU/GR2oaiDbRZbIqaFhAEaKL
TN/Cijd3YTQ45AJlOVhthkbKCUgKZTXdGTcnnIbNhQaCjJwyD29udAwVMIJYxf6r
roREI6wbE1+0twvn3Mte50xgtiKppNgBi9tBjsRpoTCaVGQPGRjDwbEQCgW8ngdr
/IYg/ABeDvlzlmk8GIIjTOcjqPs88xaMhpo+uFZz65JU0ImuhsQOfz85nPkCCi8G
PqQXwo4Tl0l3HkCpVMIS7enNNMLEs90HuHvrlgi0wT2B8OjzLVSkKq8n/eN8sHd+
QQtyyaLUruLX5D7grms8llwn0PTZ3kXglT9rCRRpxU0rIw3SM1JEvB42Ed92n+Mi
RbgV0L7Mvq30HvzJO6as6E9xJRQr1pKKWfuXKsxWXqRFQhArTPBdGkcLLEHUivST
Sp1P4Ug93acxChE9bjM+H3hnx67v96zfXPT3aYsjPm9wuvx2I7+Dw+GXMJlqJzsS
cR6zdRtYD2vu3DefVvHxHeaOsDLBNPCLhkgMs3ztG2wvJkHuNZq89kewJu5glcz2
Hw2rupxxQdPUeUYvcgka3kam0EmKqKDuvGTN70YVEPPuQWrdONgmn6LaWVvbyGC9
EU7ZUEc5MIlAH/ZEpEgON9oEar1DBgzz0sxeqHWOseY1uyRsRTTDlD/YnXGG1QvM
TSnJ81HwAQNWUEF3G2cZIecMvKCpdonwi02DBVaWT/R0jfm5hvl83PspqVfyBRb/
/sOP6H7H7TkSBWh0GUyHQ+LWe9NDnDJ78bZNU0c+Dz/aP9aEOAiECeoE8misWd4b
q0xgnCQL00WmVtJLMBTvS37lUc/Tw1UD8Pqak/4NQ/GpAwOrhZY0T8vq0KsLeqIA
cA4suqO8evzyJk0ifpqX7xhXkjEGq36vRxa8Qe6/Mk9WxfTk2X2qe+b7q+chfYCB
cClbFbVv+xv32b+Q95SjG/O5ZDYUKKSFuKYppUxPAt9iPD/cSE3uQzkzVOsGQ5qq
yyBPDe5r/mIqUh0lR2bcnpsN7YYcJJMZn6SoDNsYS+OucYprIxtykvGYgQaAuA/B
6TJo0cQiPqhy4vRoyKD4oQ14SfeG+pOrZK3NrGpcOTO4UEkeQ59XgL8+QHylAFHO
94riEZSq7jPOGfGf2FlpVnWwRjGKtirWMsqux67EXVLVG4yajhXPwb3fB2imWFcU
+HSuOrC4S/5TLq3oHu5HgOFpbH5wtLAg2TGzGqTkGzedDLCIgz96lsAO9a3DCgoS
mOmkOXhtMbjORYI6oUMOEA+bE6ujOnmu2lnGVfYQvz+3RSKyfcmio+0ZNrgCCRR1
U6I4vE9p9ewKQzFw/bt6apuVyN/toBxYUKQyOZ0hCM0yQ+1kdSVaH4+jvllMcolu
GFpyxa/c8/QIyS6pBNtITMB0IEdl8NoI5unbWUqieJ44MyqSpskxv7e2iI1ocfSz
JiOmsE1EmpblRtEOWXgsyd2Nw+uTgQp+oPCLFn+Qfj4nx+i8S2+0xk5T+vIWPIjd
sE0RK+Zn3jTdWtmwgvapgpeIO6TkJ/XAjm8nMi0fwv1fB+iI9QUiIf0JIBoO39Xo
WD8bM+NvBB8OdIYMIH0DrkXSswlhIt0I2+ckBfihOnGJqb6yGnf1LFBAmRc04/GH
hdnNaJDaYGu73cPU7Nl89egZZSfT7QbdrOYSugn5T2Jfc3tdfXOv4tq8EiYDomJN
Pd2ft/47z3CIYgNatch4INIXtQ2g7ZrY7xpCq6uCHTjf4CvPM6Fv4WYRvYW1GRUa
PBNHZp8VWoxK3bX6in1S6Yl80ilut9aRxj6qliHfo5aOKPPc0KUMFvfba7HHgAyU
kkHS5laIrmoT9dLswvMnRycVukzkI5HIUJUaHdsGQunuRp/oNJogwIFXXq3b1V0R
QglMwmhCi6dxM9h6b6Gdb7Rv+97Ls1iqhRQ8v7ZZWSdFxhCS2zCxruQVGIBvJ4eF
FOZEL4xMWeIbzcxsRHI0OcQ2SlglWNrCb3oemuEfthhxwc7yjLHSpj/86hKseXVD
NzSgPqKsXrD2utXrYv7uNPZUv62HLKp3w/hMAbv2q8NlUpT5DshgowgJwZHL8FEO
BFjcjo+Okkzj7k5B9nNV6v2LX9aLLWd2WR3C02NQ6R5BELRkM9IbvQ0TvfUHfXB/
WQDKQmpGq1BzeQIVIA6YNYfn7iWK0IMkttNCn7vRB93MHMHuIoCFvXiQOs/MHNeA
npSyAPDVIyy1+F/gsjxbly7usrjIjKQEVjLDlyi1iqwJIO7Dh4ergqBJ99njluwm
LQvRBCUKriBKp3UVtUTZsxtSR7x3g2khARitKJ1A+v7Q8mH8A1HiLDXMlFJxB1Pp
SvhV3HWNM48TqoR4/MrEPERVF9UOVXhMGsEtxdSNFhn9DL4WEvJ1MT+6MfyIIODy
vmUllDTOudo+pAq9E1El60OlDwm1KXElGu29ACM09B3lw0XzLDecBGn53DZVcGWk
aGM0r0lK+F0uEOuvdSFR7R86Dtt71Z8/GLoa/Pv+JzTayT7Gj6y+wjRYqgxDA78i
0UmIhqDXJXTCwBzWGBDkp5UmL3TehtRohx1wLQId3M63yePbw3Einl09xJEN8abv
QtJJseJUEm0yZY2OvpaImDTx2Gvu7PzDmwnbBOyCJFvu4Svd2+f2M0n2OWwSHjKV
W8/2gslaBks0am8fkpdUmCBYkwmr3R23Mqae6DVm1zs226YWrv5wSiNYXVqIbEpX
TFv2AFJaznPf1u9r8hzRzX+Wh1b1/aLRXLjyU/6/Y8Zi2IMv0mcBaXp6NsZpC/od
EreQvctbnXfuD3iy6WOJh1gubMmIBIvc3Ta4z3sQfZ//RJ9bELQq91r5d2vfwlnp
tFFhXI7e2dHRjeD2bgzA6kDlDjeZZBlAXwTYi3z6vCGa8B/AF4tq7yv7hqnOq3ii
YMmnX/VLpU/w+rsWx3yRoJ4cB4li0+JEipr9MJcEL+yA+pkEjAP3DuY3qfqKYnXw
CpQJez4SqxpBEWksWuflG6AWJwtCYjiO2hlmfQXeyvh13cDfZzur/v/oC56fKy/D
guyHLEyYC51ZCrpCTOJOuPNSp8nW3Gjd/jKGbkXo1uSl0mUq2Wrquyn+cDm8eTM2
msJEwtl6DEkKxCUcjEbGs5Vb5+CduVQdSfkoII5Nldvlepcy2c0uMiB2UkXYpM0Z
sK4pE6GOm06DF1efDlNXhXARXUAa7va/u+a4RLblAdaYj4Q9vUeiKUv44oqhMQPb
elaIb5lkU0/gcQoXGV5/4FuDjde4c5B0kRWoLkMTm76veJTeJKRC04yXrZ99lxbE
m0sacSfgUQWddHOBJVp17fk3jwqF+iReehNxJ4jvSVPQ5VwLMhDdxVrKC/sdqsEj
NAXMczHCKvohfkuOns76AHpsDNn4j9d+lE3T0P4BH4mCIKZunRRXjsiJtO7PN5AT
2P60cp0FsVwa/ocyK3TTQtE2IKSZcufaSXb2GYwMCZAi2JwrMOfK1etoNafg8i3y
ibN5wdngeIVLBZyNBT2UH961HUKQSX/gTJHe60Y0ZgMZcwzWL1r6e8uk0auwQ09+
mV86RZPW+tTn65cihOr5gY47gMBGBuSLP5bvPFHXSzaOOoLHnpGMkU7e4PT3TFr6
Fp8bFinb+45Aaz/kUqGApb5Cv6Gvoc5ErngyIh3f3u51DvJNIVF/ieu/Fy3ZvRkG
sQWTKVzKVcLUL6EUdg/Q7l0KZTlDe1fA7byPeGWX2P1xdzLP8RuZ+BqW+kK+kbld
geq4AUUnlc3rmKcyMyqVIAGzwVwSbvP7vphGYHAkkRO+CkX3pBzUuWu8secDhYss
VB1W7j3dXGNsfmSNsMGIOB+wfhSY9Y+Gvr2TimRjbKGYzu5PMbtVFuN2mFLNBwkG
0mSHo4oelF4NNW26ISVfdhVA5XH6y74ue4knNfbvNVXmcN5dWPhkX0vT2iZIP1yP
nbs0BjQ6lCpS/1trT0uS8HjcG5iseWChd1nyIshJ6x1dJjyrgZHqt1JaKLCAWSCO
qnQnxJwly188bvK/HCY1amGu61TgZ6AtdbODSC/gp3NfCIrJ/Glj/E7qE1q61z26
V7WoIyuBFv49VfDKp9zMsULnCb+vZlApXLc4G6/yxazAt67xGiXvC3dC0rciKXhT
GYncxiXzj6fg/mSAJl207kQPOzmz+C18PJQZvlVA8hejup+sUjU663uRdf5ddQ12
P3+UahW3cZCK7Gs0bfDTycZk+WPKXwEocZUhTPJH7SXsgCioUx4+Kh8m4hOGsIo4
qHPkr8m64pfwe6HUE0BMPoTaDRem5v0kmS+4SgEPKO3swdRCRki5/N9CCazV6Luc
iy5wRQw7KqN7Y12jUzFlHkMRzJ68/5DHvZd5+ob4/W7PLj5mGNELOGe+bNilu4z9
5tWsYQZaaiE7X9LiBc70rwUCDLDx5I4q8Mhtyo60h5f6bAHh+8q32npWLwtrx+WZ
RCSsGejPhqAF+tgHS2URhnItgofNdmx3d/3PkQuT+NKmijvP9M4yzOd/g5oVCS61
I7ZXQlR/qCUtH8bN+kDBB63DfZlSGP/7Vx30/FQiHKLGe/C7a3Q79O1AbYgRpZ9x
B+myjHH30sJNVDOKrQfMxPYoCoSteSWuzyVmRscTuA1jEkVZmthfPDRI6/nfuWsS
PT4C3fVl/wtVsld/4MgF6mhJo2AYJNso9hBKKGG9dtmRJ1jHQxeSNwiXl1Aushew
fo1A9MdSqY0cnJwnMcHH89Ntsb9gSt4wxUWewjKpWX6QfQDYWT4ZBx3MKMJS7eHr
HmFTtrUsPQcuvIzNiai2PjxEfhLoPu/trmrf80HLjn2LOtPLSTJurTMcj7b3tmtn
CrMRRbaGOVDiK7AbBWLi87vejo0lDgL1/m6/pUVcLTh4TQc02ExVqIUktJq099c3
GHNF6hgRaUwbEQN40js9PTRSCtWdOkY7bh6QOWru2u0GnJBGxt0di6Iwyn4+4tZa
62W2+yCVHddcR19oZQbIme5TyZ+0Gv7OIRuSwSxyXZjI4BTsiDd6Hr/CewgKTRjk
DNtUgnkFhBuFD1ekugVtjzVBS3anZsPm8gmENvfgptc37XtAfBBnRebsjHngmBQq
aNEEGiv+GYKH2EsZsvvhUURAdv1deH7EZI8TK+8JS4f83fphhh5NNBWYx6UgYB7k
e3xgCkr0IS6Vmdam0gW3nzmH4CmzIHPgSNUTedrtWQY3VfofVgDP2dweU4wi+Vgw
RblfWggSlCOS2fUmQrIxoLU/iQunBnT0n1gYhGeLVk5g46+QpU6uSV2xHykMLojM
GSzfCTz43OymYPypsN10HX1OxziyRQZCzBjY9wHPjkJdkz3ZcN+MqpLpRPrpFvmv
TP5UYrNDQlv9QA3eipp8+Cv3X9iXrAZVzlelrBhi/1o+MeJUySnamhNqZk2FZPvi
dihh3J1HJdwVvaO6sBEJMbvDqFm+Nq3tdalZMrTpELCu2JmiuXX8TJ3G1O14sIbi
zAt50jAfmCXd4Co+XD9g0ezEeSgLGbacliCJEtOR5fIrP5NM3S5B+rqKEK4OWBus
k6SuorzdaPIcQn9yqqku7n5IT2tJkKtIkcW5MeCdZ0wWpZ9EMemAtzPKYrvfyDOY
24KX9eBJ4PAh0eTBrfI/RFYmdCw1d7gInUWi7bMRB5rmfaOEFIOKh87HEVqTxAr/
y4UDJ3LJ1WQcepk4mi0mPuCb0S0k4itwqFnEupQwube5ztGjgLcAqwqKYKCerBTy
ACJt5wAvHuvb+Q5YxSrHeB2WI7Jx7PNZhbsysbeukXBBHLfKttcGCaaucTUm1JUH
MqGt4PeBBK/ZDw2hh6yuMZgnZ6kZFWcNNP7CKD2iDr/m8nXMwhvcxjHTLJi+mr1P
7mOjD0gkyq0htM2auYo3LnrZrDZS9FKNFWN5gU7xrwvOVvCsOAyXCSlpxnmlVylj
tC2irxMU+eHfURvSfpjA4hxok0CVbNCblyyRqaK9RDpi7tC0Zr+KOdaBmEsPg8FO
4MDRRjGonvrAio2IRYibmMlVMgwl/VqAcfPFkKmc1Quu8p0/WhpovRmjbwgCx2pb
rQwMoMCnBDL/KbsLmwmla77aiOWTvhg9ZiXZ3GAL8psTlWqhXBFoiQKq1s/ZMOlu
WdSxSt9DLybUiOOwHx9gf5ag/FeXNSFFbRv9saATJdXJsHs07tik4cwhA8Y3e2xR
iW/3qtmce/3jehoGRuLZv4J+AZ1Q7LF39jWkIsQ/h1faSFyrCKK6BokuPnaFa+Nz
mREebBamhXL16Pj7/Q+Bkhde/xG1tcbOjWZz0vF92fB9qsBByMecKxTWBhz6/pEA
oNMpFfmowK3Fg98YxbqvariaJQMpYSw4QipcWeAcyY6sKyfJQsZmNkLdZljYZQ7M
FpS5uZFva5u/AiSaHXIL1a8RpSp10FC1Da/zQM371G1SknWSp9jePrVNGM5Ypb2n
+1b3aSP3bJs1a205EBzaxOQPoFKXGLzjcLzxVbwaXmlseAqqgU1cMwa8xTUNh54X
nNhJrSy2ZsKOUyr1oYODqIrjW3vBBaS8K/fkJ7F4OxC84ALU9e2OXEBjQxxfNJaA
DFvatmq7yqSKepGK6ROhKRJbjUPsjeHG5c0wnFRP9l2Pt1KTPs8FFOMxgisw8CyB
fclA+bSr8qvFnbIQm8sq3VZbF2FnyIT0qTl6di3JDoIMjPoA4USJM91FeWidOfTS
JlYS0D2nh7pRw/O68J4REJ6yxhBpyvjJgSpqSbdHBzWas3deNFc1y7zi7cXUsWs4
GdOsrjPzSMDI0OpHdPOuYQ44+b6MFicFGellNHqw4hlIlJo/strxPoC+XB2wD5M3
FzBVo4QK052n1LTtReuq3jp8cS2M3KG+vZfqDSxVl+HlncFxAin5g7sBQYYzvPBV
DMAIoB1ljoqvcC+cKll+vot2f91yBf6sJw+lisxjELr8e/NmsF/J6v4DSi8aAGfl
+iquI+v2Sl2Q36hz5z+3y5IkY08IeyE7fKzUdbUoVFvi7G9xs7C+kXACDvA5mPZD
FbNXbEsr4/f5nUkHscibvL+6G3YekereQJV3BGunzWsYbyj1qXCcYGsah35OVK+R
8XrBkQ9JS0eFGF4dFybGaDMMrTqAASJDP8EUG0AHhmSys6yfyHO7eqGEjRIPFdk4
aR1woGOEEFR6xhlg3zV1owhEYh93uFUNJTrjE31z00uslyRf9//cSiw+DUMXPrjo
4m1ZyFLPGUbsBr5MFDb88J0M0AaB8SHnERSPBZmrspKD9edm4Px059+dY17/8G5m
1nq1GOMow9hlvushhtv5W/Ej0lWPUUC4FFaNT7eaiJ5AfVJpirR6+hY06AmvnCwl
f6+ljiAy6kLEG7eJPNZWnV/k035kyairo68+zggDmdBK0SckrAmnquqjl2tIqEtq
YqZ+DJOIRBrK7m+RzbdGGuj3six4aYSqvbCBR1hQZIMH7eFQKit5xQVe3mu4UN/L
rZ5moR+ucPpDlKjce7F8Zh1dWsxZl5qDWR/VL1ZR1JGziFjUZ0ESPzBrD9A8GlVS
/ySYn/rpyt8Hw8Mk1V/cEMz5+Lxmd4ZSf2I5a/MIDUlVOLDRP6DrCsI+qhJjTYRk
UTQKxFv11ahW9k62tnqPy7Tk+T2c+Yst8f/vYUDjPVO0qzr7ItF8qLxa/rI3Rqm0
PlzEMJ0dgRn762s4cfHWT5Dc0/F1eYrwMobqFL27U1xvhcas8w+uO0oD4Gge5kEO
SGLq4NKBbewD9wO2/a72eATWnbNeylSkroVbXkOU2RQZ/qanZmuqxDwBZfVMhxsO
LWvegbo4kNfkIa595LC+Th5Sc6X19gRw70XCp1IRms58O4yr1zCVUfNo1nlgjntm
WN9hhvWJjU4C61ga2nYykTqp7JM2rgvaOXQbchl51YOK+HCQoddnv2HOq8ZFrVCL
HSdvO93Lw2yl3d+bN1+ZOPyvEn5G6u1oHHw4JAU7uXSOHGDk6xMeHJopiwOBHauO
qWHKFUbw+JGlkV9lZrTEvkjLPHHL6zfDDYdYAf8oc7RRTWWD2T8TzwNaQYwcF4Q7
ylCZ4a/pHsc9G/GFlxRzcDxcpiQR4NK5phmo4qjkWfaZKYRM/LhQU/sElodPA6s/
hL7cfquHdD1JLZCXTl795FaGMfjk7TjH2wS3ba7KGDr7hJ7aPpiF+2bVxtNu14B8
prpZjQrY3wLZ2fiA69kLJdf6JMXszWzf1N8W+y1cZevisAKALdr2KKhrzXWk3Nu3
Ga3KtcfB9Pa0ml3esLJhKx4qYVFyOpguuQbHXoTe44uennaVCR2EOFaHEzKPZmqC
Z83sJ2hy3gZ9RZtT437VHTTHkgKgrGXTRwU7v8a0hI/SO4UwyEKqdk2BglKwKUdh
3J6I0//iaYj2l+t3aieC04PePIuL4INSKdRX58oo/BuMV/3cYL12cJqe3TlQanur
NO32M9r2wz8o3eW4ZAxbHK+ewwTWtEQVJNk0X6y5sznIX0lrpBbsPh4FaX4j3mQr
JssWIMSDnKFe1If9wK8PlzR/JA3bdm6rYxv2V+gq0L9S9hnMZKgdLxZxQtUev7Ud
CayhaDZggFIjDG5HcCky9B9BD4jl0mxIQlMhyvdstLx4W34hJSY0nzb/+lyQ4Lof
Gj9ImY8kZgKA9M1N3UOD4gTw1PZTU8b7+TZPz8ekrKbPID/0wAnSGbpNRwArV6jl
ShIUEuod4fa5hyiPnBLairadYrELy0KqpJAangDM+wLuxp+h+bnmPWNDDuhPSnlQ
CTjKE1/F6+XmHVj0eQyntt9gid+D9Qvo+Hvj6XnQkIu4V9vmBhOKWty+104348wG
46VP5nxWhpjgo9ivMb8M2SQc0KaYHoSS3xDz9tKrl+JtQO8PYnJ26oaVTKjlwC7z
2PwfAmZvfXtwKr0ND6BGzwWtoUwgwp1yxUqxqgZVEWL7gCCm9YD4VakUL5k2tGQK
XPHLYI08MVbAR59AIPzjmv51i2Wj+7i16ow4ZLoN4WBUyx/9VS3Je+7Eedcocqgq
l2Iy4LbJDa1fKt3U3xYvzzgWaWmboL4PsU7WIwJ+DNyCNPI28WWuZsQ1ImgROM7l
wOLH4FElH5OUd0S9eZIs4XE3RUW5QExj3dTvt3xIHzkboYAuSwxeOJBAXpFEhQqd
cxjsWcbwkTgdCCIxRsF2ENoVPZDlH440Zjuk2965tQOuONHDmSUsC225IJdnBZJo
xfHE3wj7537Dv0cFsyO2COZzMFKirOHBtrGhz0QKBUWmbg43DnyeC/iSWQXzYFDB
FQhZ4aoIeiPu/i15jDARkdPOUcVz2viKjjh2vM4VEOlPsA+OTdiI2IarSpjEHPdg
MzQk1rRVeASXUrJif16QVPkGkNdBdPsVfFdLE0ZiLo2OLVMbEY+gzFAOwbA8rVy1
gKVDMbeskLaSZayMNoq9Ct1t1XQy2lwGHLCNCKwIqeODbHdODQ0aDQB9wGB4WBZd
UJ2P/8RhcVFL4V3wOfN8Fi7KiHkbb/TV88C3Eoz7qMCrzghe7GH6IyXDY/AbQizZ
QfUxrLeZLWL05hRKXpe6wbB3OuSyST0ZDoeXFd28uPH4en299MOH2Zlc4HD+qFck
zGBXOdqxxVrYrxy2LNILAPO1qnpI09xEy7+8HcRhQQFrjyN4DMtinuZhdPA/ccJf
1e+rw+UJ6xChkN2yO1AQJsbnQpQzOwLNLTUgg7/rM5sHeTe/cyhpMzZY7/ZHe4tP
WCxh6Ls7wwEMFDMNNOx7mYXU84quK2LYFEIvSVKYSJXoZU6ZQzAKPG7OLpTRvgze
r5QDetjGlPYesIMcwyRPHFrARcKvJlnJ8cU7U26vMLALttWpuvj7XIea/MPeClof
aiJov1WhMrqkht7Sb1Xr1aNgsVO47g2/iv4RSrlA64J/KkIPh0RMIiGzaapUQTwN
2DJXW7JkfgCplC7sryaJ1Eu+K8vc6eJIU7LkgVPMXAFQ3T6Nd72ZnLT0+Af+AYSc
Am8ucIr6RvNs/+BNQBL883AkQlVYV+CFMW2geWsp6g+rVY2WaTEMH4+12e/1iJLU
K/B94ihK14wVfR5UvsKiEnHLQqZMdGK2uzJvWR/0wtppqmX4O0/kbWo01ysw28ED
hFdg+akuowAq6UWWE6HAWbgC3RskInLy3T+ZJeSGSFLFpOMVqhkm27F3qGXjbZCs
jxQaYOeWi0S9vJG4b/UUAarlpJSmEnRMaQ/VaKvN54J0refcBCrclEko3DgD++uu
TVF0ntNVWAz8eKDfWeryrfyDsPPzEAxgPvdjQ5lr7aMxCtLwCPu/XgnON/AhpII7
WR2ehQv3gKDkP15VY6/RlUhldNf9W31PmQungP+5hAQyUhfQRtJH/tyFy4d1A5xu
nh0vSuWbk8z8xfGu+CoEO1qU1yoAk5BvKUr7gAHfH9CbIhVDPuJDipZITcng1vas
JDP+Vtra2GIN4/bClGyiOmvO0vl8lWBoTmtvlJPSzRG41cIRAibOzphT7TD8CljR
mRpeKawHRIXu3KWKf2QSOzc++mX8pkLGZ5o74C5NXT6T34amw+DvIWGA7tT2sn4F
mlDxXnpRU7o+jR8Vpf6Ft885rbFwu/qQ2Dn2pw2dbbFXU34ceNPhbUzEajYOV94Y
a/cEcMu70c+4BVC38deo48fOhdIUZS4uZPKibsHSiGBGh3LwfefVkFSLeC4iVfgX
Vg1qcKpPHGT3dTx+Jl2w/mTbYUJ7Jrp4VvEukfKldsqglKtjGqpBmbDuLOtVMhz/
baY88C4CuJfeNsbv8qtR9+64TzivZS4SDXnFart2HMufkaGkxobvLay2GailDrB0
3LI4RWM5oOhxlZPZSITfJfghvFUTL/DfdBGTQU16bpJGPKDgS3uZWy1GTS0O9UDS
QGQg1/gb5qQZi/lviDAMRTmqZ4/LfrKu9FoKePbWlkhTzzE1kdN991XClOrtpQFq
1ZMgAyHtzIJig1vHi9tUHyRMBK+8xZF2zHISOTFdevtUVnk2yOOr2qIXN3A48vDe
DYI6m3U3KvfqBR03zyMFahBmSrQA2w5J2GajzXL1FyhP09ATPRU2pmPA7RfoN0qe
bpnt6aukFuaglR5tokNQ5EeWYwQxjjl0x4PdCO6CGHG4PkPQkoboMGX3Pl65H5+R
MbaTDg06ERQQI/HyBKnZ1AL75xGfOnRbk0TlRH8YynlqgO2tMCBDZluk7Zwc3pc7
xE1kzQZ+eHHX1o1BxFDV9PYqG651PI5Yzv9SKNnFe+GG0K1HXTRpfDvoSlmY6CpB
P4e9N/hnGEW3BRsvANOSfKiXf5LdKwwOwfj9APZAAZJ2xEsQNv9FkSk7CFBvmkup
aGEOktOOIcFVEIj2XYEXBsNn3q8qV5hn4tnsIlT3oum6SVGMfVcCCcb/ch0kqOK0
LxC73GcQPjkwnT0wGc6qg73EbmqEsy24eCgIVrB48XiQ8YiLzo7/rDGgZrTd8hM0
w8CcWuUxQYJn7fvNeXnH0QmEU0CErrd/Da3Nc/tuXibihDzRVXbSrvvzNXr8f24w
N7HFQoIzOxELta3CNsG/lFvI/6Gwi7e6rfvguVrfGus9+rTWmhs8GVWsNbvWIpAk
npMQ6j9WDMZ08BK6RAzVwwPuHOTxGfIxHpyAbYy772SXJrVDUOdWDYXkdbg8jNlN
GCVgpaoTKZoSC+4E+SINTOTGJzlaxIFWSXDKPgNWHgCnIlmJi4J62/fA+yUtl793
EczmNPadkVNLy5ccgkz3yXilpxGhubakukryNfsKXMR3WPGc9XpjJmSVZpKbZiSC
yUnAc6igUm2ANXH0t5zPa/QBN1lYZEc21nhkZeUaaW/SYhOYtEYEptIe0ssE8qWu
op/CTGVLSy4MvGoDWlJOakgaQvYx7ckd6XQhsrEld661sLfwb0n1BXICfmwXYh3o
tqCfNE738uDVOEkgMPv+ZYVlBcUntJYAMy5EgsCsYVHnU6EiChw0IYRFV59GBpXy
tcD6JwwAoAGHRVWYBCcitf3ZDtDSF7ZdcgMJbGDM+6N7ewNgF/zNEyOkrcnot59x
lDbPfDm30qmslCiaPAO4Oaj6UHXvY6OzdS6WOoEYPYj6QRnqDrVncDOLRgGHuaoj
7cqKv5NHlLkM77XyEPI+yAro/HVvTWn5AWkeHNqZbO6FBseGXCOjJG2JLDirJmop
x1NOfVCy/CrbMjHJVlAUo0dAceXop+Xb/65DL0D9eUChgecW/xqueDkOuaa3dHfI
h7acMb1GJtQA6YVVVE2H+EW0ewHmnYIMHrI60cBUlSRkaXm15d2tDGeN3GN+Nvxn
tj7HM75ZvDuw9XG+ynlFGxoPb6vg+qOBO3g7YNEZYKy8EzrVMmHOIpSE+X3FsH3I
UfKA1hFE5zcKNPZ/UihSSIpNvA8cVgOtcBN/tn93ZiYP+AgYtj195s6lMa3XCO64
SRhIJU1grejSKm2mQKLGamdkcQGO4GOgmp0Wp2yJyRqEDm9yq+gF3DB8MbrUUT6f
+QpKoUYaAM93pIWqa0na0AMh8ao9sAXMvxV9xonYp+2niQlHh8rt6i7zo6WjbuCL
lHV/UOhO+9sRhQqm85DI9SlMSsR0G4bO0eye3R5leWmbAty4u4kUgtW5npUJ4Gnx
FDNkvjElCOkfScQ4Iv/gzThlDqecp8HYfPAimc0YSynq/1BoCyZXeKWjkIegITBV
5xZvLiga89wLDU+OP3NOykzSEvCbm2XLoOyoNsDCmpVvFawLfvPz93E9r67wOdBw
z2O02qKhM8khg19Si32Fe+B2YVNUu0pBpUeYnHK4gn4VtoX6MQNiFD94FTv6zEsG
aDINcF4pyaOI6h6aFBP/5afvKE6KyNt+cmNovQVYjquqm8xkxv6mWx4b1oZY0VOT
S89K5Zz7qLDpIuF3kSUfVhXOqv9VCnqiRRTbE3eNfJxLK+L89iA/Bhu3QDveXEgb
mFTGUmTx5tWA7LtKFtwN55RK0K6g7LrTfmzWDSdxurRvJukWelcb8r7twOPW3aGO
9MN1aUkuiC3Icro2b/V9zOkM8VFUPb2/DSRFSWYfy24DObH1x/TfDcegUeVdUCjv
nsvLOuTiBXPYEg6gqhzeQ04018kKiqQf4yftChxgVFsfbK6mUZAIBSbWyBAkh3+C
uWXxF77ADKheKvk4NkeQMNGBp/jdrqhRy4nTFoPuHeOhCQRCMJ43DypKVMTHfQJe
perDl8QR0RcMYm9fU3ZqsaR9iJFcuBVkRqOIj5CgUZiJAWLdLxqfdDkj6A/DfhJu
gINirQvvwj9tGm+23D8KyAkpP/scLxf4ZPs5Pi02buqsSmlVkRsUwe6LyWm64qVm
4HfXzHXeKHOHT1Ez4h/TJkBq9N7PTa83r/vTQ0b3WnWxorZDDkVGDY9j9nUurZtU
WeoMpTLySrHUq+ZjbpAGsevPuf1Wg57qexwg1FdWOFQl8bYfNHABnO3C5jRROFp+
Ei+97J+EGbi23bUoY0V39FrySOO3rRmcmen8zzbWcT/KRU7paI55f5oOLOXIInny
3PVF1H2m68gL8xTlsBtLVTA4UO8yLUZ1xOkR6ZaSFwiDxhwdJBY6AXHQwudtgCJz
jLfkI5iZgAdnDlW6pEo/CB5+lkZhdRxV6jK9qHFqj9M2wnORmUaZ7RyE6e3SXEhF
Jgs8YNAetPB2SJ5/Fp9sFNHrQKyEguuooIygPwlclmJtF5D2NPhm9s2BjScnz7nZ
Rkfn9ADrSI2Itjrs4f9t7oxefxkOtdqUm+IL8ANb7LVxDR/NwUIbkt9Y3rlP89Cl
Gl5mGRCTNpkRomU4El1RVB57cPgF43bpK+V6psH3Kdlj4M/BfFuEPL7oJzkuAEGf
uX0OoO4RYf6K2KEQw3RO7abQogxL2NnvYINkyPIszYM6WP58jzLOsI67Hmh0fHOp
re9UiOWuzSNpJ5sugErXDn6w018xGRNr3mN6e9FrSqrui5f1qU8N197C5mZtSEpP
x2lF+reI4UY9Sx71W8mKbj92hbeOSFpQW1CVUA66LSxhc4u9gGrVYVA24lnxC324
EFtrHJ+nRPwvWu3nD8r5zft/00fTDjvRuewF4t471vkUYVYOuLuoKDpfKP8sMcZK
JXWKKTItb7oNdMQx9UKoJ6mdoqqUTmMyaeHMHVxNHTQidfwoU+IumYD3gfm1UJke
B1UF1ecyuVvs/gToUOyLKU0bZmE4P/hxHLaKVgBQ7Q5f4HjFrUSqmlWE5vLpqrbf
91Bmh54M78KTwb7O/gpICPQjSsCQO3PmHMO1rOcvtnoUtGHa3QdepEFlnegoXdhJ
TitPo+34LJrj+dCNbRZcbBA8JThjxo1KPSN7Wxp37m+ygGUJ9xivMWx2Sm+W1+2s
7v7H8eAbxKngv5J3/MfShkF2LTE4xsVEJLznObU9fJ8ikpaV7TeUqO3ah8K8+trL
HpVvCkcToynAZAkHT8yRaAqYCBpW0hl6EHV6N4MyJfYiDbve0tv79oAPOIkEm0Db
CepVVG0BmLPE9wPrGjOB27BYFbmUN6tVZFWXBxQBg0ztff4ydYX2bxEP6DwqIUMB
Ra5WZH/Lgz1+X+LjVJMRGmjq5GqlK/yElpJ6RcKvgSA92z+ZjRsc9A8aKBDxkdxH
/R1A+CavUmB0HD0vzqkT3v+aU8tVZhnaZmLTSgf1FpB9utBXacb4G6tvMTQfOe5u
L2BQ79rVIH0hGkLoT334zcyYC7k2UvjndgCWwBFRMWaz5+KotL//J5Nm8DaSt4cX
vsD/haMiegmKFH8VQzOgLm35k1l7K+UZEBpKQAjuCCQ5I1m0lanMTHe/J4xyxh7o
OpWlBEsBEJUKRt0i3ITvHOvXX8N/dm2Aw5IrqHOdn3BaheTCNJZSYx/IGsoDBxgh
9PxA6dda5XVhNesWFMduGWbEGwMaOd0076YWJaqLXHkI+Crh/KlOETydoe1EFMsY
TbK2+l5dBFdMC+RSJFns58SGQNRPVJIDsg9HvUv5Z7l8a1Ew2tKBVf2AQ/JAFZdu
0YITzEff5wJABFAlzzsn3tlO15H8F/Sdk7EABOpWOLpjR926KpuM3lDqMZpfd7hH
SVG/nEvgnFnQxKuWl2aRahr8pOROQBXRmjTgCQpgzhrWnz8Dogygj6AzPW/CUUtv
P2keCxqkh7oNNsYaZoqjNnD6Xrgl5jQGoAWo6AlakKt+nTskgOI19spxUhpLVjMK
ZAjL/7UkFyYcsuaB7Nx/DkOBFQJsr/wPSr+iw3SHn46wpfchYyLbdtQJLbKnanoe
R1Mv92F40eEoea/ybB4SsI/nernlzPN5GLJA1Fkht4V69KB81zJE/R/Ixe7nKu/v
DdEZD8TDulew8Qbn/apP1oRNJPCQB7q3FZ9SjtRtLXrOdIYRUtk3DwohaC9rih8B
h3AOv6vGnJYDzj3HVXr7wBhnv8yns8LYQ8CcZmGvHbyfLfS6kxV3coNaMy16W3Nb
A74S1GMLb0nc5S/XBF+hme2GutsbrWN4R7iay6TgeTKl13EKNAEvt6gZ3g+XFf6Z
IYlKQ4QMZS0h0dFOsc44N30LgC+tp0P9iqsari75kOcnQN+B5BLTdMnoc36OMnJP
CT+FasDILGVdLFR32ep0O4gytVMq4wm0FWq8zB+bIYHLcyBXx5eVA1etcyiCiZjS
6NPhxgys6BylqTDNzciasUbev79OA1eZfmfz8axBu/hMCAKhTY7BdvGm3fsyq5NX
/Ta7FpSlGK41F53ChK2iICz9iSEpkycpv43RV8VwuVqwDo8Ss+0qtrLy0sIlk+Zs
gjm8Jo26MB2BKgsTKynxp/icyJwDlhW0WEkih2n9LzPu/4GieXNuInDSGpHt+qfY
7rfyOSYCH6VwkSjqB80Siwp7SdroO5tYSA5662ORm7Sed4P6t1VQ4vqv7WlDXfUR
65CQSd1D/1mW9YQtPtQhY3yt49A2ojgrvYhKBiuXqnLSQfjB078Ciq8PytLq3yjt
SreCICetSON+SGf26AAeygnQ0yk2XXc9PLqW8l8gtZqcu2SFWhxfNAdtlQY02mDm
APP0so7n+cYQ+NIes7HzDq4CkMQKV/ATxNdiOd0VlrGmXUc7THhQhaL3CWNDlzLz
78Cvl7FuOyHXMot18Hh0mgffOljPII7dLw16bL3+3Fho+gEkj4M40ukB2bxJTtM0
mZoe92OlYfs0w+tlUKYCsPdNDtqJ375XKr235sm8UavC6q1OPRH0w0gXJ1a0yyuI
8DIkOygKs9sO4lXfwLJuNSykT5Ko11zBb3EYYLGVXT8v6WLOCemqTcMg0aZgrdbA
AR2qlLyFs+HQVLvCr0rnrdo9vHoYXxL39w5L8Gwa1EYmktLrO7nHR9MWmkdNgOiq
3OR7xAdZYrgqlYbUEYEC18tA/XdlX7HrqQNVLujoW5yhehKWZj/A04zTXSGOciGa
Vz+qI10hCrdH0FydpG6kMstNtxxNmHo9F7wBVXB1NVtzVExYN+pkNwj5fGA0UyXQ
bjoqPOg1utnUPeW5D13gEpXnaTKTS1WXeNOrE+fZdVH/0rj0DVjOS/VOgrfQmh21
LzD+1CJr2ISps7LTYiAvuXuBSWeqAWBBvjmYoGBKbCEOl8jTwUYDAHzJBDQXuceU
U0JnMVsAwb0R9z7zLpsCCPLmSH4VpVGtzWOmRCR2/7LJl3MA5WdMViJYLJ0d720V
qhLlTsosB/4u0aZyQOpEkZ3YLQ7sSVVCApgwLX9LS3mid+k2wN20hQAPooEAGtWY
MMWPJKb609Y1lPWYGqZ3HYRZAfyYgMsvKXa5mWzEXSdVbqSjKXPTPMIdkEfBw7IX
aFJkO5DvQ6/t2KyZwTsfslWdEC05861RHrbNvWO01g+KOT6jKetyw718dO9SpgAk
w6mg38B2xbluXhpAj224coLJpoanBeI5sc4gJWTxnZU5OEbPbLcmYSl9PFo9KFZk
s4uFVCfFTRor9fcksRitGQ/rc9vzFgOO/PZATkglcNlsFk8MfZdTF0cMsT65as/j
Dj6cAiETCMb/eiJ/UyWHH59oXwWken+hj4Lg3kIZj80xlP1dzkq4aIV5iC34o52G
LguX47d1eiVJtpfSswKDpj0Sf4FnEHfO2GDI4kxrOQby49JWdkovTal4DcrmmBQS
1T9DripEZYUKU5CBP1WS3zMLKG4pHZ3Lv789VZnYreVeYwddMga7sjhpAIgV+9kI
3rzgZ79uXDNGbVZhvaypRAw1+GMTexIl+kn8OlEgHg3B1muAMTHpv8TtdcE4z2XZ
E0nN2fZbM4X0UWuktqp/3+dJF7U3jFepPzQE8dGXPBo17IilbPZUuR+Xh6G102II
9E7o+ZeVCIPtngyrsj0tS5+KIoDR5BkAtGOaLZ1AG4sv3fDH1lFfRriwTcqYXbiI
/altR0pMsk2nDu+qUmKygPzmWdO8wWjEAZWp5ggcRimSWjhXKutf+PSx1uU/kh9E
iF1tfKfE+/jv6GBJqEdc2TkxFZ0wNiI+1XGmfYt9cRYK3R5RoeR6Hxgby/S00Ce/
O78PnT2M20n+6G124eCYVHMZ7crjKw9K1I18rFxux/FAJqtFtouU+Oo8RjI53sVL
hp5zcBUtlw7txDebYyVEffDypedVl4xQhlwTGTpJXV46OMLosXm+cfwDK0+2YyWC
aDbYTMuwbu4xylpdonq9tp4hQhQK6cZxPnjLPYAYMeoizg+ePszwYdrK3whLoRpy
KLT4vGI/LTeMOurMUlmmOSyhDGSaaXEvaYu6v+RAjkGHT4kO4jUBcgweVPLUdMz1
2wfuf6v8Im5j/7ThvkGPGpj7+9WX/yJ8mnZhl9gH5F8GjSN9PuWS+DC8GOCpm8+m
Xydu+pfZPUcGaWlBZJAXrcQHIIIeqRDbYtdpKwdorEIJHaTmNdwKnM7Pbu8sX8tZ
me1ZQoSEG8piYipUMfAnXTSVERaDf61p8WOgsi27xurnBx0EFrIeg/OKhrjgTHqf
eTIjgj2htKcf0UAhvtUa/ANLs6y/zXvadlpCTb+ippG/dUqoiOdemKjrzUbZrAZM
qXYHZPcvQ6hpEEv12AcFwVyOrvSOPUXhCyluiyfIS6gvqVZYAMtfS4wU299bOvra
MtOspf24wPECl58C6npJXA59pP2oE5pzzyHnFGwI61g9Taw/LtBX4tDNYBX+RO3U
7ytJ16g5xBLIPmwW95qeNiri95ofwrgcUf9XMY0er4qdSF8YdmcIYhHbaTnnglgo
XryXXRnsDsOMBy5DeiM1tVtLQC+D4ce7KeR04V6qgfQjD4NOG3ha0ZF0aYgfXwBb
nNPAzrqTjmW6JwqaTKxwqsaKPq8KE1IH+o5d+WCPC7TvBzkTKtx5MikKw5fRXiSJ
gUvuDmnZUfIIsQwxuaNvCMULjsRIRKVbdXKqhuK2ntxOO49ACpyCU8sdxPSh+HvM
Doj0RHi/Azki8ozjLitgo9Ydsc8PHPrdelJ2L2DpABsRXLQ4vWrJWDO1QvLSB3Om
IdAaDoeTH0V47ZAi9sUYw7WeEpWB3DTBG0AqOkQEqKzeArUhcuCNZ1lpDZnFgphs
dH8naBcKc8bscnAWcssGsp15JqbWeEBjPA9ttgC0kd/m/2PMwaJtd7taaWRtYDRF
nKiRtBOQfcl55snrhyh4i+0f+XaVY6GUURIlmbscJ511Hja7tpue8aLpP0jKmodb
P2eXpRi3kyxb+JvtMMong2TvVZGDAF1O22Nplh3KX23dYprk+q/Oy3fSdMhIL139
yTIWx1iflG9TbUoX17RyTzG82/xP1M8QdIU5ECpGa3EMah+9iIeSa/2ZpHEhZrWS
Y0PWM0lbuzPS+Zl2bSBezsmmuUnxobsGgwsmZJhsv+6E0eFZK/GecICn01U/yCmH
aiEFhCFzp/jyZrqH2T1qUiRuOzePjdKamVp+EAkxtlB6+B1NcObg4yZRO/yA6DxP
jsvSzoPFiCzCnLywjsWvr9iiPkmrh+kVuva7hx1MDFTBT4SvJd+CiJqragjXcqSf
iWMyYG7dkCvhFeqXg1uf/74nHzz4C953saA2VvBLUkg+E7I5o1vOrDcxKJBkPbUN
PFK9vLvkSEN1URsPUOXhG0JJnHftBcpzZZlNG6roOYOd7KAT4Vscp9HZfZi4Jzgb
2EBRrQG0zS1EIK8Vguxf8y1b3SQweosBk3vNkw2htNAW0heiiL6bhmrKjfSWTONm
Q7ELDWStboAMFEUI3oM/cM4HS5f+hW+wNeaf9tJ8my/kPEDWAtU6mD9zSygZ04kE
3JDZDqbAhTd04HBqEaYfloZIEgCjAXRw6UzrOvl3Yg66gLxeHjzPtd6zgIkmix//
SgqaxX3yRDd4iAEK3XCtVf5pNC5ndb94iu2UfOJlZWXikVugdAhLWwkqnGNcgFNR
X8rkNKV5mfwFPgqce28rau6fiqpOpVn3TuEEXD+M/ZPopxcorKe75YYy7TBjdya/
4S8ZjOLmdjsrJ5wYVxc5bByABefY2or14s8+K+imyHr6ahND11jCP3StkqRs20xp
JSD6ePf0ZAKvmY+zN8QMg5rFXEeVK8kq1FSGgHBwnBIFGr9MJy7rRPhSWE4WpZKF
xRaCeHYBI7vz6OM2XHDo/dX9R8smQpYvfdvwh0Ec0f+VkfTY68dIe8WgA0wUMcTp
XI2qi75TmjdSY9cKo/iLjzeNgIbVb58JDhnblS9i86MGDVfhQgZanvTE/3xNoGGY
4DM4ETvY+coQ1Ym/wSkC/2QkqXOnhoU0oKzgNDlRoWvBNeej0fulwXUZ6RjqrrTI
W9KsX2pSWlIpDP/eI90B9PCKxOww5bXXYFpDZ6QYYK3M/rV/N8fiy4TkEzeZO7iQ
IHf3KUa+8efstEWCo3xAGgMuktKyy20e8s4S/LJlFV94Sz4VnCxii55bR3Ujb5X9
EDUrWXIBn8YY+mbPRVB63G8ztSdqKU8csgYjU6uEhHJ5/1/EZY9Yshqk5rmqyBIo
afpAm3HBwxN1P1gX+s689Ar1fozwOz5jmU+qOwirG/quwMaqs3z6eCpWrm4l5F2V
T2iksG7DICHgYjAo6vM1MDJzaB++0oDdSCej4qXhmOh+RHCGP68+vEmPAnHbt6mr
Qns3L9DKUNuLUqMY8yCF+oZXmjq8xr/n1kKXI28CVvvFNl9TdSg4batw4utQH6cK
nf3ypKlT+nfM/JkK/gk+iQPXchi9hG8wUxDQp2FlQ5xlD7kAthlxqwbE63QKYBuR
u9mIf4sj8x0c/GO9awNwToJAMQI8NUG4hWj44+q8k+Q+RuHBAU6FfC4k77+Bo0jg
DoBdbLXJ4V+xK6QZL8ZhLJKbi7WIL7eMH5NjjuL+g/lwipTDeT6xEJyPKsqN/+lP
jsJ9TjSZ5/nUc/2theCsUM4oDbqqgCyEJBtjWEWzH6e0aX94VXhWBLLSPjBNcFRc
Xws0lruL62os8pAKl4+DEHQmFJ5b8JbRZPE0G3PmEyddA0WCYfmd7y1vi+fkThiI
P8N253XWFw4zvA0ifWsVy8b5ZDUMH+MNykAothKGPtx7t5l0lfbOankf+iow63xZ
pAdTRFPEbo2Za2bzxzaaL1iXeFXiXJhQseGYIYmz1KfywIAUwrzGSvCTFKyOHspG
RzD46fgN+jUBNjYTqYWTFxZQdvHruBxdF8qxYfDiATcmC2hr+WnSai+7fJGhHLxW
Jdrd8UuuWtxgjwqzDF6LVntOaSHiswmZvD72MOPMm0YnLi+ebmAaTJSiuEp9toyT
rW7iBQR3ZnnVJ+sMboBC9kDgd3NldlGn24MME6B3ELSr3A40e97/idxmZvFSuz2v
F6jOohYlgu+wyxU8+suX19iRbVoJSfX/BTQfEmDr2HW8BjGE4K//+ngGl+oxKJR0
gqeXr9losWqFo+d1A2B5ezkX7p74O3aesWX+e+h0Gvj/rSJr2i4h77s1m4FrnnF2
wkzghHUar+W7fUCd23gL+vJimLEYk3gFlitjb4mqTEKH9tOOUjwBTuXiYcAS6RRv
PVnqq5J2HUVJbBZGqRHDpMAxY8b/FAQtp/nc97z61g/87Z+XqAWEq7abkKYxAymf
xXDq4SSgM1Jjm6C9mhzQ05lTkuYFpD5ySNutaYGwI3ik6EO89RKoM9D2C3zU+buX
07qtMFnAsLJvX1qtJRmnW2xLiShq7SBSHy0Ed501T0JO2Enk0WpvFk7weNa9m+l8
eiRM+xrKBsWH8TWiBP4OhEXKPWVc4MZdiMCYpvMhEJHAOrQN112C9keBBbaEdZPs
N5/UfT2RaScReRwRDDZzyaEfZ59VTDpoICHyJ2ZSdXH2CveowoYZtEpO610UPqdU
5afikhiJ/EisHWVIUlliyvOjwKhBUBEh2KaKOeO9F7k9EQ+SK/p8h2ZOFB6qm7s4
Fl6nEu9svCCd7Kxa9KE6UhcX5r0lm3W4qEbHSJ0sgDz9MZCJGupomrSVx439+7vB
ReNzL2zpZtsv4nOOFzMy67AHZdLQzE/+l4IH/ZhjW4muVR8ChO4pNY7D1Mv8wKee
c6CeYFp2GvIpYTrLkZ151gzXHtl9uGmSLAJyjF0qgwk++ksXYZD58mkI8oprDnu2
qEZX23G0y74Vv5mNs3wZEgkA2th5bxoy6ngHIWNaa70q3j9iZ/9h/Mzfh/FRzJyF
z/+f6NNuutRGWDV0oatXxOW9Ds6O8TpQwtXSw3JexpVrNnpHWfM+KNnwBRobH+tu
FEeWE37+vdp0DmlvBTRlIIZDgdbgfHwdddGQ69KWME/YV+EdVV1PYDR8zkcWU8Zz
4LO4DyzQueJFW7JaPv0Y4WwA0v9ymStABAAamrR5hWkBbpXje8rLzjkWu2sYEk6y
k1c6DO3AE1y0237p5hJmBqS3RrZNoeTRi9AKBeT1eT+swA7HR/7befvmiCElaRnU
sefiwGcEboivWHVLVyRPeAKs7Pjzib1Q1pR2kDRG6D0V+xRFTI/GbKuBGKKGyPcB
tdTWdnKCJABkdPKMCTMfdibasC/DKzFkVRNUqQ9cXX+7RwbGVM4oa4hQcQ9kpltc
BQzKZOQbWX5z9yRKwk+jU8g8FPJjhS0msx7UJgI6iQTjiqyyQmW65WORPA2Qpys4
gOECmrXbRrVHm+6K3ZJ/rFcbm5wWCks8chk/OTiauiAYlvKVSpfEK0w4OXc6IQIG
KZJ+80QWLD/8kAvyB695cdDD5xGv/LQc5LPLuykXHCqVke2mwylF9wHrSws1QctX
tCLq4U/g95pyTTUefKr8WnCaVFwH0gm8iP5uO8lfH6ePbNjJU1KysfNZIRvK3VXI
HxQQIu/r6xg4WBLgoE1EDuvP2woQweHIL6euBclRUCjntYKJZUo0AN7GinpXMCyJ
roFAbA1H8OKrRrsuhokWO0g8jVPBwBtUGNeyXpUeOFbY3ANodxE9LEEa+FDmtkyJ
q2E1N8wphP8dovTm+uySzbIpE5mp3hu2Z/yg+Wf0MO+LbpHs+rv7mgsNPhPJD9Ri
5S8VOxefLljD++AjnIYI5EC8ZKbFM2GeHDeJX8aaxEVi1U0oJdrDaZV+sFtZTHFk
sgHkMd2LXfxXGr5I1PpHDMrC3G3rBBzaNKlNeO0ANdFaLOLk/yfsdn0zAqleV52c
f6EQmytp5GcmQyePDTqks3jR8Y2I1ZYsl4u/sdshwA1Ctk+P83Xs5LPtEXfsfJN7
VyuSj8Ey8QomLrWAGuYBf3UFOG53pkvmYJ+S6A57YP3rfcdisVZfHrOSDn11864z
8XiaSyL16UTSl3tNwbBx/43eRls8f2drORGstMkWQXvdOLJ3y7qsyWhs+URHBr/Q
g6Om+ZKzFAq2IaWRFrSpReUzPs6mCmLJStWIja1Vn/h+k9wohZipFSKTJ/Pb9RIU
cCiso6w+dL7ITwUaTAV7jZJYpCqxlHiCeA5espE04iUwnoAHgBB8ndi8BDAHw8ME
0v0QDrTvrLzfj2IWqAAXko/EyfiFaZ4o+z32Ey6POroUbQTVvdHUCUTqCJ07I01U
F1B8aLOHd+AKsFu81jWgzu0yFLwC/CcSZ0hJRbh80de6pBCYaqoXKXb9X9HpEiiO
yHEjJkn4Yk5uV0gjR8WI63GMuOG3KBKszO9Ymv0v1U84LmQLNK8f4ItPgajoXS6Q
CiBF1enCmR5tpzvUzN9iKN7wGGWvSygqJfI6U0hsJ51IGMURS1zORfJX48wXVz7L
af3VqiBUGCT0LX+UYI0gtS2bYfu4inYHv4xMD1ZiBMT1XQ+WB1920rrfgPCgkOki
0PH95g0zydK0aI7xFTwyj3kKLNGty7v9pjuCYYtWkfjJyoL4GT1DlPXUJQbzHISU
wUdW3ae5O1Q1i68iHYmB1MGeEj+Vz0RFIDlVHvI6fkgbToQBTiXWme4ZQK0icaTy
l3ymYxNZAaHu0mGNahsOkfwEBqja4SM7F/Sh7REyj1m5e0DWiuQHLW3PhKu0yp9Z
C+/t5n0lmLADsUWMDXp7Zdz1blqU3UIJqkAEe1SYFQtDtBF3Wno/X5ocRSHj7Dp/
9EZ9H/nKxT8tPH3mUV1mm5Mw0pfaQbWOH/zWCEljsNZWS68vBgRQCzcu5rJYacPY
90cnWMLeziN82suQC+1d0TOTPbeU06s51RAc9TN+xyQN6DYItVzenuEFHGoDpcBb
dT9KJoYnaqr3aPbWPBidxiEo+dZbLdcnoewmLBCXlqg5qrVytnK10jy0qltqb6LE
w8WHZxzwukYQ5JqsOjEYSbPyAmGl2ImQid1CNg/NXXmz5UtC54eZRpK7Y8cCTAUy
oYUFSZclUWU8Z641BiBIFPaJCEzP/7JUKhfHrqUXHkFGYxUdvJO3GusTqfMa9WX8
ifiFB/BeCyqkHsq9FxC3GltHy9yKc7QhPr5/5cbITn53dCYVC40oUEZGfn5h9lOK
FV5uFfBgKRn6bK9MCxZtXrN0ev3vfn5s7Mb/JnEtPJ6PcoTGfowFoBqxS6ihVaMl
mE/PhMCeYIVVqO7U9AzqGmFL5090f34AiBHJQervHaNwGeYbia5hyEaQ4u1YdtGV
S5TGOopW5YH3AHymwTCGkGXakGtTkYB5QdAzAT7pGiju+I9t2NNxna/taJZL/6RB
ixIaOD+Gw5biEUJfO4EDtIzRA7LWqsDioVC5GUe8XlaK/JmTco59Ie+K3yvJnYjP
Kwd8LSgERegXWnqMzdhD4FAnCj5fBfPL4AFKfNf0jy/JSEEGoeyDIwRHP+RC1wQf
loYv1/fAY0rAJEQWPT9A01qEbP3BwOFOPxz3glCxj1PEdELQl2GGcuNWmialDkua
+eaPDPqplbFEBiRuWTwu+3tvyOPiJjxg1/HrvJTzKDsLtXOkbmFqXVRLjZC729tb
Fy0B/DU1usxXYn6/j+E2uzIFLHQSmEDz9yLSdoF2xDV8keAT1Z/aGHvirdoqPEvT
ZlLiFn0NGOelsGPFJPz51ViTVEQe1SdIn9rYO7PiREe5YmW0i012aTlzIaGXq2EE
dh6g3o6gBT2HhKxFtGrgC/w/y7oeZyhtBfcoze6yGRuKuXNC8JEFz1IP1pdAmb21
0Bd/ovk20ZARzoByK0lsPP5O8yPQpgGfW2AZVyj26fAEVmmLC8Uaut46ub3ll+dE
Ml/3g92Vc4upXsNvFgLB+CZdNpdfLI4PTahq/dE9wX+2rMeH+HoIvP9YBZPQ5Y3d
0ouDd9KgbUg+teHaYgoq2EkCHg/I9dGi4CBRKzyKvbkRUYcL4DqLYmQrGyNGCikd
lIGCHozx7XvzfPYGW+TUxLEvuEBS0p5RChZ+9RGAF+MO3fw70bcja1DYKl8dTAyt
+pChoWJ4mOYXFb7nzuHl/LAyhTJ3W/SGMEszlE62DEfWX0i1c9yBDYdHFRp5yPNr
LLcyxMODeguQAZqhFiEHpjG3gR24xR9+iLSw/2vE7CEGeyFRQmUokr2L1kPLM8ux
+Hy8AtCgQl+1cZ0IhmyQL7MRssU7z31QopZSbmhacnQz/7WrNGeuzYoHangJu0Cd
7HncoonWDpYYkzuhvX+xc+orlwbNpb1KIHozSBIDm7X8HTy0cWPWqepYZcynHbea
y6jZpR+Mlr0DAgACi20jIRdrbQ48KrnBzhcwCbXIJAoq2N9hYISKK/5uKmhru2qb
u7J433nipmA/05k6EDfiwliGu5of7AlzD4uPC09VRcJ9g25oXd/upJLd5RF+Ocs6
N5erlVxQ60lzMSPK5g7VMwHMTJ/9vuRN75ehYTVwRNKY5w93uuGJk8imykBZ8tVa
bHcpNJKJWfu+NPOzbQ4EbskeUWnQH3L0Stgy8ERhTugV5Re/KSnDuyeitRFiGmWv
ttxQGTFB3XNK3aXjRkon27OAetkmym3uOjRnMehuF7XWb5nAAhI8qmWmS3LzbwhC
1RkWM4FdP5mOODwdErNnr3zo6JhDpoSEA2k2cfP92BF+wAdqhvMAr4sLV425sB/H
uKQbNWgacHn1shT3yOBQbGC5IpH11f/18QVIhHNCSgcTdu5Y4l6H8Az6SWpHkWq3
d/lSnsEIAu96oxXc38T70o47FpyM39KsIkxBQr/mvR9lKHXr2QERDXZC3QD1kMtE
jow1ZBHxyOVF4WxGkh1r2xl4pUoTlDIwWr3ZusjapaTLxZ0EhvZOJQf0DzyrzF6n
kF/gS3TDAGxNgEyY31mUShQppAvflu5XBYYk6JwRv4QP3MHHukUwKnjkgIsUPQ5i
AEKEfqRVPeNu5c52WSus9+XND5GUZOSDsJIKoym0Q3NPUAj9xJSMsJNIABTMd75X
DiKpNADqgCPes05194onIaRFKOXcSkCXCrJkeSfxK953w/LOfW21CCuOo6Y0IRmG
DRCgaB5iqi+ObCQ8pver1kG+sEyU9vPnPqT/tgbg22+d54cSVQKru0lo7c0pnBbi
JTdbGf+/nB+ikuLb+h0gV120jj7VxWn5YBzEmJ0JLnNoDBh/X/lU/L3RfFAhobp/
gs6B3Pl0UXzH2SkOuuTA6ZsvUcj4fTvhqkT3MX+YIO5klNesrfeKGpIuu/WCZxlG
AIR96fhBiJOBH6Fbu2F/bGXYp+Pi7OtFWAWrEL9PNGok//KcKKDPxtzCKOKBNPD9
YhNyVxpq+IYiULDhvuHeIHg20oKC9F+GYbXNvoar3iOJbNmaWz8mAV7IAlca3pTt
KiIbnjz3MgXThys+n86lo/fCp3yBVCtfLIt4Euc9JiT8nLgSyvZNwtLS1d1PcABo
pDgr3o8FDon2K2wDDMx5UE/nA+5ltXw7Q50AFaSA8AzMSsCtDVRv8cS+ZUb96EUV
K93K67jbwghT15/pbxFjNCSxlqrqpO0Aj6g8Lv/Q3WoDtKAf/4oJK/0OynaBltNB
Jh5c6W25Os4d4TiDnsEx5te7WtJvttOxtOpCRCzOpKKuMulZFDUw0ulgMpoU5jnG
AVmq4dStPzsTO9yyBNiFcat2Pq79hm1JzjGH02FDLkEIFDF+B87mokpLgDWT6QJS
N2j674zlfjPQaemLFcuqU8Xx+vu1ssOJH1igBQTFn3e4Pky2CGBWz4OmE8dGKRRE
1jdfu4ZhabO8u266RhNPA/DtjIJ/i6XsyDk8OIMpQ+NCuNWeIMjHARNBh38mGH6n
Vpojg6Xc2qN5rogKUl1Mio79YnJ5yq15KLJHy+Ka/bJacf+gbQMwDDNzh3BE+MQc
kR/wsrYs+AGl61AKHQidRwiUp5E91KYtvmXSRMVgH/gYsIGkLJ2+yCU6EURZ1ag/
krX4Jj8rn2xwcWYS9jwymyPDHxt1q15ANt3mefIh6RnbQtiVzkFruN4l5w4U2OyW
gOtH8KqD7D1xUeh898x5hrbaz+zMiYA8ufny8puFjmhjbwqc7J8ouDymm29A3cup
OaRU0deC9TJN1SMRuyiuI2sYUwpsxnF5q4szie7Oq+ji+7ezEQRrSstIRlJWDLsI
ikF+axpEiPc4oWgtggTVrJRZ5cioo8IbxvuDstJHQUwajfowVammDZmAcdezq/nr
+kkYmyxbjQIPtKj6KKo3vGyF6BrnlzJJr37E1BeMiCSGdrYPlUQHDUVDy9cQelK/
7GOtFszdNg1WhtHeIHfJLnIKowQd0UBvu5SKuZB8fDNw2UUGs4PGbJ2rUHne2arP
Vdax1gT2VjpQ2LqO4zYb11FtFZ+TpLH/SHb8mXB2sf3q48Y7RYqF1V1DHBBs58gf
dem+CPPbgmvbBcwghhf6oEPJhkdj+8Y9UQotgD6TyB9jxlkWBvjcNpAr3GjFjBjl
31luJAaeUVqOh+1cEVRWoKRxv71E4Pvsc0uLLOHB2LNoJJFyxzFXrlEsMycu8EdM
cAem7r1j7NGgn6lgHAQnieFSXglUppHTQQHfpCR5WOa9GdAGq86JlVbarxeFw4bq
Vn8FpcUW4QHP4PVFL+c3W0sHGT/gkQIm3HXqcC0z5Q3cKu6ZXseud0dXwucxDQ8s
sLRapUVMxFApd2rYwPUE27hluiOMMr6K9JOobrn6MgFxz3Po9C+WzCk3T0DpCFQV
R2H75xLyPZJfXzB+seU0lEgePCHjxxxQS5i4I4HHxKYTYvdTcfcixd1WE6im9396
IKJGpgayGX52OnqwwM8P7SELpKFUTn5wQoOOmjb2aPn60ruKP5enPuLOfx7T4Hw0
kcfaig+9yfp8XsQ3mAy1d2XpN8r1vIPIQGXKDO3HtbZvUDiBU2gacne3gAUA6FzY
2E2WG//OOzA2yTDp/2QN4Dske35u6gM2TOaj+IIQObr0PaYUB+r5dEqmlzZdajRy
H6x1kRxLb79+t3nLf0IWQz0yWU6SYmxWNvDsppkwRwqRfaxbuThVWhI0yOWqQeUB
xQ7x4EQpa8yJOmONNF6Y7uQZ1Hei0IEPO1iJbngwoQIQttJgzO+/PLIvI6BnjaM2
2vQvUOCD4qaE3ikqUvByf104N4a7hvMYE4OLp2p0r2fEDwgTODa05HtsZovvRQzd
8D18EF0pqBKV3z9a9/1kofvFDsgCd+iQQPGqnA4UU0UahjQcAxcGxYWa/aHcUruY
Jmp+R8g+9OijdpO0k/ynwzdcSuWyGNdcbe/Ad/adQFDivFYJmQbKqaaKGenKDup1
ZgGPtSkaCnJiAb7fncDvCVlgGqgXpUR/CPoZxGEi0KPKEImY2zhRBUxmQdGT4CYm
3NCBR7xwx5eiDFOYmYo/lOibB5chpNJutfKv1eDvQWOTsh9cWlRrQUhTDAZtw3AI
11LASA7VtHEL+6TKONTJKlgQwZMULAipm24regvF7DIW7mwUAB2NptM+l86w4ByF
J5rmJnqI1eUsnAj9/FhgaXPWN2HDSBA130LMdTw/lfAE2fEHsqBM7E/E/Y6F8kQj
+JohYaeeaMSe5VDhapysxdIiW/rrB0HamnbDjcOav7zRDdrkgfFcolKLA6O51/pU
Xaw0fa8NpDJWH3Rr9reo3OWElzTAkUh4VRPsmJGSiD5lCVe7aUCM3Er9Ygx+pkHn
0qibPARvh0qqHLjwiybVzrpBtdQXJpiGH/uILJpr3mcB4FtBNaQ0r6/tY1S3fBGX
NgU72r+HtEojxdiB7lL3rJiBjo853UOh0VcQtn8ruFax4AOS/GoiQKITEov8Z+Ct
jmvy7jD8vrncX8n3NjGWmDo/I9ncsWHz9yjYfLAnn14KLTRBwYo5nyFrhKetj3Zh
/AR/4Cnh6RD7fqogdXjw5Q6DEF0me8qLbSverUHSH/xVmvfY369S1tueBMUaCGjY
28mQZ+OQnN5N9Wzm9eKjJJ5/k6jAS00EcCVOXHR2UyoST8EPvRtPjMgSTcHSeAzB
jyNAevTosm1ud9MkkJpI69OGfSUhaGi0oNJSdbsxqV453+M0xr7DcQxpjnIDXFuX
zHrcG2XrjhmQ1Ba/+qduLq2VGU8witS8Qi/sDWHlIJoANzBvFmwaRe6GEkh/S36e
VsJ7/36VaLUJE+jL0Lap0V95lcUbhbQ7N2vvzYM05wheoj60HJ86F/8ywQR56KFa
/2Q6XDI8YVbId11RIFMEGgs5eNElqn54nomCkQVMQ5eenhmctQz9HGiD2y3pF1Xx
YyHdju/R9bo6DNfC2Wc0fDcRvf453Kp6c1iM/gIMc/lsd/dQ2hrbsu34gBya3e8c
KlxisL22EQGvJqUF3CgpO32uv1fxsloWZUmH/IMZUvMYUAKe56gwwlBbsV+JOD9Y
ZkKeKQdOPHihCwW5jehfbAQsk3qDFuL5cD+KHXF0+Bp/NX39gaGn30Db1bCjuxVD
k7Aw1qNgxbaYSBOHnpciQnd58ikSw0+otqcxiAdB08bFUcnbPjiSt7kwNLgYU3wV
/XQDJnn/PbfImsjTPz6R122OECpYANjHRONAT7qgXArBlOiwNwCX9LSiW3eFn+B2
GZflQ8M7pL7Hav6veO46LZq1KeFOUlwmGnxCwOrIJsyS4qf5Mz7qoJuNitak9BOY
Ga1ZGjcivKtlp1MTUE9JaOnxfbk7F/ZlBI3CCJtQWCjgWdT/+AyJKIvEcDTmtbSd
JYetAYTKu2IUZHm5zK4xGiWE2unglQgkw7Nr9BFSBOkJezDEFqC6PXGGaUZtmlzy
2fxC64J/c12yex3AscdGNgvlVgYwbZ6Wi/hx7ELO2Ftwtls6kYg+wG+mzHt0iDPh
BaBFi930WC3EeNbCwAYgQ3z0WtSSOdb3kAim8Yu/4pEDgHZmNCNlHfRUrsWIl5Jo
Hrtd5AZ9VfGGqcbtJBoW/5eUari1Ly1n86wU9lYhWIukcyXB/RiTbCg4zsmwpBhV
wxxmPZloNvJpJ2luxWo3RmdFI+1ucakbACpXcsgl/2+nubNhE3ejUZ0UBes63CD9
grF4IeD6uYurezy072PjvcAksNkVc9CTxSvudEt4R6OzJluIEYOBce6oyvI8dt/+
fJNRxuZDSzf1o16mlq3NmTJmvVEhuKaoSFT0OTdeu3pDb9atAU5mCYNotwezRNlA
gDctjXiW1HjuoRLBN1+GLWB3tijL5PhRlMiE4zY44QWzWqfjDF7rrNd+Botg+M6+
3Z4uSszzO/ADt5RvOE52hruQ/p/mwrACb2NsEgWvPq+igQNaA96BpJnkIcdiEeGl
P2WKrFAUSpg6CqBggzEH/iiNzxk+RZMKq671j8vCR4oJvGYQZC9926NpbWnGZTvg
1tLNP+s+jXwHrDHVD/zntUIRU5V9kwqg/Zy+iCIX16X8kdbkIvTzKC7pVMeJuWXu
355iQz+h0jsD195bksTA+c97dopKPl2i/vzz09Gez7r/wIIoxQgVNNe9U3gMvlAI
BroEPAJIP0uOpn+9jf8v5MJuAKgWNpNwYp+kagv3XGs+cbubH7kRXgBQRy98OYIK
Msl7YKq2ym/wAMclyj67Q82vkGTN20o8qasV+NnlwlOUZblPmSGvwMpMANRT8Az2
0H9SaWniBjAbUSzQOmdG6CPP3NwniCP6D9P01Ef5RT2LQ+0a7sZQD6QgIcpRCK/w
PKX0KSpmswfk85xLtfKiYFQDdN/mMiqdtkn4iP9bZyEtTy15Y44jOEjcHn3EYicF
xTvk+aN9xrZkjMUnR18q9S/Twt/46QuReCvS64c5bMz55jMw5Qva4HgfQJFE8dWN
brNI6ua6rzqDCOP3wLoYyZvEIq4pkjuvN78bgD5n8oeGLAg9YXtt5TYGkwpBVchd
wuO5rpzMAszkOSUzlOa6B2JFM0HQQ9Si5/5oIsoElWtPu7kS8V5qnBJ2YjV+dVkz
Gep1MKYYsZf2gcc+L7L0RdTWTx70npwkf9qkczHVzgY9tv9vGDga/eKMlTwuwXUR
eKOKuBjdc85D8HKh05uR6Dg8/IomF1Igd6AZPkA46QDRtTRAU4TIp7bheZNyb1TZ
ftotRzTDIRc43S8q+waaOTz91aFYm5bVHyp/hkPfNK3ww960nUu/VVDa+W6BvvJI
+sZPDacSaY4l+aE1KOuXsMNJdtBuTpLly1qLlvG7yX0CUyNUHm6sP8gCTKIXp78/
h8iGzLgvKIzkLw1OGW8+AZFRPeecGIK7C33pJpqacDtRMYxX9wHeHTCl3F2ZhWg+
fF4RHduvzMmPgCWR/aPSMH0ydxDZG0Tp4xf7Y9a7XfsnQdx0YrENSZ9aKlkvdZ1q
H0rCSrMmcclx5n4cvzbnsPTcnYT5YQLVn0ptHRmKRv1P4DpdWScK1PDZ/6KBFLtI
daxNq/XsogpyMMNg7MuoVG5792t+WXEsAvEPUVq7GJ94p4PwrqR+/UcWKpPjZi1G
kN7bN/fb19Kv1x2mgKEPw6yAbp/QlKKGu6tMjIuYK4texFx2TAjgXpjB4+u9APsd
t7PW1/isvsMWjsROiL+qTddoND77tIdu7uR0oap0cE8ZBue8Ng40/Yxo9475BmET
fsvWspqFQc0n8wxmN8yDUpNNlpHsJfYawsWT90p+YDuIKQO2U15N/Bg7/7LKy1H6
UqJNvmDgFNoh8WkorMFNm6Vla/gz9vDhV3riftfcRZg4bZg7ZUI/kd1BxVvJ3M1K
gjOFwfgYZW4ZEWA6fuZEEsY8LnkZ5mE/gF4A4aPs6rmFDK+jdfD/r8cPma/ghrQ3
w3MeH2XbjEhsTHbHWXDOkzsY4pDI3IxWyHzMtYcBgtO/gMJZJxoy46xQdNazTfpw
fbx8BGE+Hj5ppUYHAyBpBQ5bgZYN3A/M4JulwDsZcXTqlvtp1/pCQ0kw2Cjx1StW
3Vzm/aiPPVWgIcQgpDMozPdYCCpXg8qFbrV4lz8HjWTewuLNIATjIuQo6GarbPqI
2ceDRTWWU5BbczmimrLG7vRVUkH1gCMdQuCS3wt6UGQ/CRpo3fSuAMpZN0p4CNgH
ZU1FFSC+fFOQCh/dw7Fk5flq9YPFyFkImRzIXOMKccj+zDSTAlCxbkiCbtGPPThM
bYfHYIvO1i0V3mjObN80rsDnmYtHm8gfSC/Vgc0OSLZZjoYKEmGCRjsUmyQ1b51M
HB9ADNpexPkYTZ8gF6hYRdKzkjZJUEIwUwjTy7foErc3cZ/5ueWa16gyuvQI8jFC
IiEThhwNWxfzq1SPuYKpF4SCvI0EA5tz9cwLOmJX8IYWxNttySf1BqF5RTPPh4yw
B49O3UMgUfRIQtf/vvpncM2T/LJzZgNKd3gsCOpiXXEkTmcs06TL/ltWDkOP7gOH
qbGqnT38mLwHhfO0Hrvq2qw9MtxoyxZDJUPdlwRIxk/EwtGexbSaLTpHlE9qoS/F
Q0fsBKuRZdpN5ZC+vtQvo3MofAo5L5Rf0tG+df1J1X7IMZ6RwTbKj19GjCDdEPvW
muPzDMXlO9sGsdmaPVqbC2uRHb1zDenzQjUehWXWyfZCh9eaD0n/gSWmJ+oHXoJB
Y9znkMiW39VoU2AbPd6ElcS4AAhXv3crCZf7RmxiT3BY6H2HPfkdk1kzZjIncVUi
CnB4vzfc1jGPE5fmiriI89m/J8ZnenFBsA5P8XT/O0wmoJynyoqkjfQoc0QH5QCV
zR8k6nnZYfzg4g6J258XrlgGY3SoppDO1V1W5IAJiK3ZTG+gOWdi88R6HewVR6du
4zqPsGMU4pi7BKSD6OmzeSKrvyjdrg24+GLi4StO/bCksaIl7G5yN3Qh2sRHsl7o
VriGWhSFMey912sYVihMTwUe9y0XohauXwJV/Tz5WU478wlgAeOBXILEvW9A4F4z
1Yp2rXK8CCXnpbw9OYf0BG57uOlwLKW0DDJWsxhSJUzdIaGa8fJPChupTsy+n4Op
ltO4LCtKib3ImPIuUh8Vi15H8BWr/2cepesNDThdhC8poyx/ZheEBo76Hyvw4DSj
2q+hRVwUXYA9dVvr2mFdcTeB5RToaT5H4ZlteGQ8Iv6G7I2Q+/HksNgDNDzSC+US
6Ru2GSp5flIQzmE5tzDwbtXkHKpksDN9vIRjNsB5glwxlcqvHZw9VcfYLTqn6eq1
3xM+30Tg/eYCSg5MknrCSLKq3GKp03QSaxpAC5J1QptAFfpkkNSn4fLGgjLwajeH
dfMqYY1xq3RqJ17l01M+AviQmdZxoJV5SfUu+mxzI3gWhP6RYDNgirx6XCsicXdw
P3t6FGyUcOJjp+bfWF6WjTz9vUxHo320McGjst+SeMpT3lNXgilOYRhZY7frbG5Q
uiV9eeQGWX/jEvPvgIhRq5vaGsCQIhTdQFQ6Qt0UhKky3TkEAQROpXqhIZp8Wu8l
dA3OPQQ/1a0LA2++kC3+oOuO9Ojok39K85Uraa/5/8W7EgCwFeClocCF/hdsvfGD
2iz040AVkboV1wy+P+1EAd6vEy9g5YxM+M8dhEPShgnBwlCCyxMOUK4DdRlkd5f0
oZdcGkVZ14nXfzQAzNZtadOoBbrRxvaEEkO3lKsr1PK+oVh/OlSd7R9xRaQqUTWi
9HRzarXDqTMcftVGB8hIgIeXnc9YnENZmnEDhY+Aujhki6OVN4wLBKkKvbjqpOch
wgwEQaMC8M2QUsQiL96nmE87Y0ObXV8ZYlXxRrVv5k3Gauc1O+zZjY4q48HprgVP
whUw7OCiHJ8Jemexg0FxvuJzdUl6N6rj4pzGbcOhq0IGp2dJFEGRevxDFPkAmvEC
tS93FKwP4+qxpYZ+TQ5bUUh5kU/AjPl5yJtn+eJk04i7SRDQUXnCbre1NXYWiH9q
UELK5g85wY8hQZ+y+n2IuDrIBOUoue7W7IPxVYDq4Su9pNINWDvaV9phqoXBXVW2
K4zku9YkMAa4/vNWEq9SwkN2ICtSjHoOPJEkuaTrw+YRnO/QT3b/wzEM7nU56izT
zq0SrtqWGa0U57MEcC2k11AYF6f7460LYa5ETGbS/uKsKfWVtQEO9vRgUpel+JzR
LDXLip1ZLuxRST1echHL1fWHdBcQS2PN3QqrUjJsELnX6RU1Otu+rfWmeUhCil9q
jMFQlVEOSbifHuWVZj+6ptDsrMBdNT3YkSYn3hErbkQAwdE4/EDTGMXAd3OpmYKJ
zx/4aB5gA1B6rFeKMGpXYkrDiYAakWKDuFVKKw+GT9WrS5Pq8tA0paofyuvSMm7e
HRQzYv5gOFeb6F1v4lwkDC65T5ya0+fzvy+b0c1zNqtR/v2OSVMcHUOZmti9v1j0
lFTQdwmEfpLWfANVD9xEfOBQUzV6bdnx+bzu3et7Ef+L9CUhtQJvawZ6+kO+9I+A
kh3DeuTgpGZ0ul8FTNmFSB+GnCSpm12FwYOo+64g/vzY1FsIE27pZiXbrUvEH7Mg
i+KifEygWfMT+WUVpJosSvb74IVytmiOXchJa2TlfI93YPPtsujWRIYXeAJo6y8m
8S6+uFWBQvDdcXWySPQ1UVyisESHSaHfwwVBkLfBRar7C1S7Aa7vkYqDZ0Cl9M24
3Yob1fYRy2XEhCdsJf6hCKsWbJh7rVGHawqXk4FtHTInO4p3NTwQzsl6DK8JqVo4
KFZ63qgzK9fb3g9+GgH9H/W2+x6BH4qKA4eDGhSXzSYWafCZdmaQvt/7GAv14H8p
GSx5sl90CjPUUmcbNoZTov5W7IRlNvMOqmkQog2nEFMNLe9vdsMfMRIQ9JKzax47
ZuGn7tg7A5RFZifupwl12eXiTLXwWG5QO/B5Q72ZMaR++YisuLPw1q74dZuoWSox
N+HpVqckcMuMvtrajLTCZd0Ipt6XiAKaDuanierH1CQxEKRdoEM7MbyyYADFyzXL
QnwWcLEWgEGmURZCC7aswDxFPWCGeXXNkeIJ+nxNxPblKqX8zpuHsSRKM70YJaA8
lTtX2nKIuoz4rkK+i3QkmHCNOsuF++XLbjYckBMIRpTcoOPcRwSbX5+APJ17420H
1esgcgV1sCqRR5foKSBDI3A3smP4RHItEtE5Us/JNG8ZlJ8HievFyxB1hAwar+AK
gsUO2302/559B+gn7ISpxtPYugLinS1iLsT21EOa/YoVDZw/GGHD+YqGOaC4UfaO
x43KoelpNvD6cpX37JnVmAFLN+udm0M+Y6otC9SRdwCTbKZRUC/ybLaPpT5+8MQD
OuZGZcncpjJf+Te9OkNlXL9Kcm+eDRgHrfChTe8JCEyKeeyGDF6RafZsMzDUj9EE
a8OJ/appXKewfRMbzdkZqPU0e30KT8g29bsBqpqWzzSG318EnRxifpfN4u/wz0v4
3AZbcYfwbSBzfbuHagm1crZG9kLmZG7ZxYoZG488/NlaRI9nTtCtEDjrt9K1+IHh
3laW/fyKoOvVM/aFkX9bl482hX6yVM8ZEFzKtvpSgkYgxDxrTvCZwwnkzRPQWBxM
tLGLOG9Rh/Ycm7ery5znqU/cu/7Uq/g5MHt5xo7gt4yKvirDSJLPosILRadGU2Sn
SCFXMWYVwsqdsh2h+ZZIlZmrKEkmKECLblHzSy8Luq6tFTUocAGcTDcCP/yFpWX4
1iSEA2gzCH0XGyvuvHqvPcFzrj3XxUEXyV6R/vOIS4PmI+1s8DjRLr0pjAHc2BDQ
HgtGqA0dPIqFZ9Cmsi0/fmgIPZM9KnlfjkxOblokkkA7zDoQxHNBIIeyeKw4bjzq
wyhCEBrVUdT5kLJ97vpoI83JPdIgk64lliQey6UbB5fAQMkM1hn7N+DtLdNadNjc
th0BLGetU8zJtijwwNU2Dy327PFejGbSlmomJsDJ6FQZWIyhb8KlQAoCoF+9Ri06
+hVgn5+OiFvieLa9MZ1OqjgfU6u3iwzUP3ST2/BiuACGYLhBTHOmf1dN90hhlzSj
S6k2MgSpClW6iYK5bI4MlHBP/xE+9Jeix3cWk+JpEUHhKdTdu0RO2DblwhY5pkpL
3RCY+5nqzPLNKqKINVaAsN3ybFuENitXouF1AaX77LYzbBavNDQg+VLqPjF0W21r
GO/5uPOQL8/n6mt++yR/Y4CoFcFoPVQcoY/AA8w0R8rKUAVy3GDas6jQ8y8XG5in
FM/GzdfSy7SGqnj4EGzg4goNlGO+aRWhZm3TDGmmn2KsidMH4ksAQqe2GUML9v99
OQN5Tp2AV6l/gx9M9u0qgnEoruB2iU0o306RteYfVLWOOzWlwwjsTAWbb0Gd9Zqt
xdCAcYGY1BFwqUIVISK2Vrvs+dgn/h2Zh2DCoB0eGXZGowFvZCWpWZF/19D4GAV/
C8NOzbyiyTqua2JYP5HWJYrl5iytDwgbawO5hYdDurYZHn4qtRsL/87lMNNoXMqm
wvlkiG5DVt0kdorOvwzwODFQlwd9i/x1musjcF+0VBNLJ5VVUFJnrop7lcIv7OQr
n4HobX6u4ijHWzC4wpThl2FolTi9MMt7Zuk17CjnpAlsRMrJaNhnIM9cfgVRCojn
5jobNwCVME5DYkL8+wOAHgfAS7zsMm7DD90L3hJXkjZamSlONmhFk1YJF0OYYw8v
S7gtPCMGd5ZO1bwDtW1TwCo+dW4+HwSpIwPJqxQBlUhODsFGGuwUrcHiH+8cknWs
dLWWya/S5NyYPtunnc9BE/EDTcQP1YwxZjgHev0/A8wNO1ayLS1joIMyNcPKgy3M
Ds8PvndGTuWWFF4tz4pl4Qc/5lkJG9kYvhfGHv+We+j+catYC9LguaUUHjJUkCzT
e35kMjyOfYA7inRZS/ido6ckS6393uEqerkgpZPFCcMl3JUBZauQzgbZk9Pn+euG
j2AxECPO+3JMVagYiucFGI/IcjsgP9fT8l44J5CDSRfCBfwobkK7uS8UdqXS4EC6
gVCIwvc+nlpgXA/5GboihINGo4pN3rXt3RXgXHLEK2Vlapy1oHJ3FSsbF69X28ci
ZOlPXL4aL2C0gEWq6U3d+/8UPtSYVShUHqfHw9zmIxo/orvaCpffCGzcrikXSD3w
2wQfPAhza8wQLbWrrf+59UQhxoyWgMn+lKaT8OUnZyCZxPSisDsvtqflrrzvgATg
D6qWvgw561lgHN/gmPg0NCG8ER/3l1A2fdn/G0qx+EyiMdqlcI8TI5o0D3kQZ2Zs
7JowJTIRP6l7Nnj0EZKesGA5gkdKSTjgFVMIQ2BAIKylRiF9FfcQUeRpXlDVjFw+
oo8kDhvA/cxhoDs5hETRmuMNCXI9BUQVRe3O4l/DrdIdOKV6AXQpw3j3tlTxtfLT
uChQczHdxxkAuYVgKpuBDlEAhMPtYjE1yqyjuOyMLwZ50kIou5L/hE+J2r6cyVCq
QN62TQBECqcd1XrQR5vO83Hat10LDxhyKN0xOluNhMp4QsGbDwGP08Kpke4iCyqf
rurMhbVUZIgvhST0gGBKhzq1yrRp+zjLKZScvNUKzij4CLVVfEyZZThNMCAZN4KC
KAjCJtTW4bO3LjA+U2V4inoG5YEUjbePuNlvu/QGx1JJVHkhN5RSOt26P0B+6zbm
XrjRjnYQQymXewIECCDoSZ5Xeq1jCzfaQW0h+a3IEwG2onXhuJWo/vnNa2utrLNu
zxP751EYm+CAFIhonXwhucAXgChtHa4vG9brm/tVJEtdL8nRlz9PvPfpEcGXQGDy
3yHicVF0oM6GmroCj5sUltIz7eTIalcBnLMwpWJXXeLfIP86kQsRw39U8jM98Gvu
QsR20ZMK5hkI14NFGTTr55n1Uf2GneaVlIrIuQGEngywVnZVxrKffT1ZHLcU4Pdj
Nsqg1VLjsXiWOqWrKKLBxT+mCVOYKPE31OvbjmKuqjE/J0waTl9z0XbddINB+RiD
tlzBK3BOOg19BOIsofRkWBRJM51BKCZC3ulCmddvYPqQLLiiU8hkn/L/WUXjKgMj
usV39AjUfONHjV+tFlYlo4fAg4meMOzOIvdobfKTeaqva5qXCYx5+4m70Ex14J2W
0k3VGwbw6EKIsuxHD3p2QqR9eNxO9M5WvQvLekNbIsGIbaXC8fRY8mekkfOEGtJ6
D1hBJoaLKtmD/I7a1mss7/DV7L5yBDLZPuL8cTbjCeAL8uA7g0Ec8jExxaqRB8/j
SBOQrIj2qRSicPWqGg1OAY54uOyt2YifdycZyBqy5Vb4xGDyj1ckHPhVQ4ZDc68V
ZTRgjQNvj57AfIL8kujPK98d1BwzroAnaaSb+KoT1HNuG/j+RcnO/YnJxEl06pr+
a/qp6p9H3vFqROtbuLlb4uldQ38ZGdWL4gHkwla8vG8O5HY5HVPns6aslwyIGYzK
VWW3fLhPKjPAeljWhXc7bNBH9zZGMR0F556Ah8cUWbmBNral+UU1sL9RkSfq10rg
sXETLTE3KRLH4IKQ/lVGp33G03pzzapKZrFItnNTM5GdP70p0JcrxexTpz/oXBRS
DcbkJEpRzZsvnAK3d7UhhsFD35xc3j9PcpKF8s4Tk6aOVujpQQH3K5WhhZ+b7B/b
9RtC3X0eh9v2mcjBkkTsUjDHqnfsJWvcp68bMc+UMjNc1BX2SMX8UW/8NYWQ8iFO
ZMsdeobfqMTIgztIDEWm1l3ShloNEhyCv8An1v6sd9jUGg2RvuUifWPPJPN44vg8
rFudsS04k6Di4XyHQq8dgX/e/akKGxbp3BLY9gZBJLShVRL7FLWES+fysMJruPFE
jZMGkXbQ2XE8fgvtOM+R0N7RZ7VZDh3uUwdkdIuLWB8uwOmLWX4Q1uqSZf8ComsC
V2HHYa8RQvlXLmsukvEArOMWDR1qqjzBlglS2ZhWiWNa3ubIviWv1faDSyuKytJ1
A6u7OscpQZ6sw8xQZSThuOsmVnDMg/zsdsKL76YwhglnIj6QX9iBGZtpxPbU3jeF
1/flfUtZB2SgHzlv4sna/itq9XR4vo2dlRkmaJrxHTDQqQXcrZAPfoeUFbvgk0Q+
w8HtbTzF7Ead6LEBZOfe7Vkp9F1+CZh1caAlzFsyPUP/p/zV2EPGIszekPvQQN4Q
0zmtCqckS/R0SrSKa5l2ERZF12VV+FqSeX2IRRm3l0cb9WdPmQCpTkmCeq1CgVt4
Xcfxo/kA/E/ZcuZZ6SvMHMiVCLDIte7fYZ0Jrdkf0/0gKw3VyOALz6oK+e+xyQ9w
/kKf+qwdpAWx1z6shCW71jq0f1sJTuHexxkLfWYwXxtoRcxLWRdYneQE0PF9WnrQ
GpRk/W6RDugNp2L0R6GfLgXgBvH989bnfjuZvCBTiaUWnVldO7JvV+x12NOC7diZ
8uljFR+HMFNvIbMo8Zqx2FGGcYf5nL/2Mh+UIgGPolUh0Ec2I8TXrLwjsEIdiL1j
Ngwn7AtAlmTYxh+RipUtPARcJtdoDh/f/Y9gKAvNgB/Sbxoe1nhgrTpMuQqm7av+
od4No+Jc8H8Z/BWWbxPFnpR3yL8C2RS5g6Gbkta4NGJ7DEf7S6uqkLUS4GqsA0Sf
Lw1wRWUexA/SPKysc8eoehl2U/iy14OBR+PcuntQwzEOIr8Sa1Cz/K52bTS5k7k2
3uRcSJdM73IC0L22UBFaPHtdk5JwGqpuPrvxAwSolEfug0QnEM/eqod5GrIHp+2O
noSKcJ3aNC9VxoF0RAPZ1+wAk06S/ZUMYL9NeZ/5jCEDjuDDrvPitD1uZMI+t2bd
UIJhGlpL66US5XspfVELBcqjUJ5atjFtzmbi/m5VJW4zoaUcl8LapZ1j+zVDl0J7
OtLPqrBvrp/SSQUwZy+YDUKdcou0BJLb84HeJ4WGyxBJLHJpo105UNXpwP7Y5Eux
Ppm+UjJO8lApZ4JcIoJTj9RAGCGVDDdva214moZ+7oUunMtcFsHz8Gd8T5cAW+Vf
50ozkd26Tts74gTGe+M5lJBNNHWYYWyZdLBCRCXG0W5tqjL0sGHzOjF5XIGZtKTZ
uROQr4dA51vw3wTBKYY8eBDJ+oGPWFs4yT1aaM4dPG6rykB8WY2NxUaRpK+BxP/P
2Fr00avGL2nA5xZmP4HDmB9pE2p2ReQEy+aNRwL9CejzRvhiTVrrFfeHkBDF+iG2
iacXvvlZGYni2uaxx/7P8glTcAV2g652BrJ5PWKn+uno36vabw8lkSkaiZWaIeBH
UbL9OAjg/oL7ueYhJQD8fS969eDKGBahe9k8C50O5OvTVCf4n4zPo0qfK4AKy92I
RQeI0c9yOtrxabExBvtCprY/2QULJretNqZtKUfeJImtHd4HARaQbQJrBTswEWMF
cL112tR6owG1SgRVSaLZ4HnGPeb85AdlV6In/gxWUWZ5IfUnuqAasC9OkucB5uzz
Be4bCOUubMIWEjO1KogkvOUTuo4jIYfETVmKEBXV/UCpo+ExLc5B9lPl4F52q9tO
9FB/CgF7PhRbCkGeD+tfA16mF/6zrZj4KyxPQzo5gqGiPBPtNRWCdAYywg4F4nvy
IQdQzl6NIs/6DaR6hpZToY0VqtDxgj2NRMFC6Us6FoA2H+s972xmLRIP1ZMLJ/Uo
ZWOrCCqjY9oda9vRlF+e/W8TBGQV6zVehsxNpRZVGJ9yJ2WFWoBGIy8Y6LF91p1M
+Xfpo7z+9ar2dIoMGmbH5ki7dKfdpqRnXv2S9IkfNH4lxsRsOQVwHhJAmGUn6957
1ioB6DnmBZy5Enx43D9uRyWbboeD84MCVVsWdFGqCTz7iHOwcowzBkX2yRFEE2j3
MrW8zQc0SwxgMeuSG5EoHGsT4IqY0+mOMKQRpa44XxfQAJeXOQCN20i2SBFdECPX
Llp0HIgIFKQqZeOutQ5erA6Y3QfequKxa3tekqgXCH/vIO6Q0q9AWkiLbpeGDBeQ
hc9hPVY9QctcxXuRxejWMxvXcVPf1GxxFS+ZFOWHuGSqdEiJvR03bqJe4NJ4LJ5o
9eIQjWu5RNb6Uq+/LF6tmSuRgf1UJSpTKhVXtvuELD+8+nWtN/aTjwl6Pfsoaw3I
OnVchZFVB115PW9QJ3jkNIRqI1FpGjNGkx4Nr8eZg4cBAeM6uqaH21SbtRpjEv7e
dyBpzFXDxXs1fYERFxkOpb5fGkSIyItI7EpiIx4hDp4EQhT2dvM6wBve8moJdlx2
3UtDV+usMNYqlL0Ey//UlgV/xQswOHmJ6u/Fm/5Bsjnla6Z8pA4KHuLcm/+qEPsK
Gk4Ba+RUR2bLjLKzSU52DDQdcJzNfRbiQGHhMFJ5fqequ2g8pj0uNIBedaWZmbnh
HlVg9eEsBBPUXG5N5LYJNGNIfdpg3hoeuGSZHTzNRFMdvry/yTo/zqb3R8Uf/pWx
ryOOInL1HRgZZyJBv4rkqnx+KHxU1k1edq1AC47TnYxHT8u6/t2Y674Tot7MWp9r
6Z/qcTr7db2PFGGmR0yZ+cd5/2ICF1I5ITi3nBR/YV/qJtMhMOL8ihj0RpucFdk8
01mvUiS88f5mEFzEg3BXe6xNgdvW8NB4hMLdu04x821b7WJmZnqUQCd+n56/ugOC
TfIQscwCamT1+GBEMCkMG2PDkNZm7JFT7Z5xIn5+261DtiDglCEgGFASpr9GahvS
qhdQAD7dZLblHJoJ55p2tkRmrI1jtDNCVr3GLS4pimveBwy3CiLBZr/w4Qjwy4Q3
nGIoYYzYDy9ruDDO7TRH851xLx8FS3yO309dFMwCbbbulxzZS74wow1r0dqUxLtB
BApLWCx3WVb+MDdmLb30YKS5UypKwEzIeyfXBNs1nCHohjMslqdX+zRVLuZhnhSB
A4Mnbes6w+V43cYZFujcT67eoUAF56o0x/yzMwWB5hKdAnyyqRZ6Yj12SGhIdr+A
uXHaxktBPRhW8aHbhFpjpQkNpnTVjXjn4cJ4UmO3uXUyoQJdY2nfm5H3jFv50t3k
eE858n63H6uMoIJX91vFoMQqTXQzn5nz/3eROj18ry+x/rGxu7FGtFqU+6scUIKt
p9qUeQr79W3uapfvZyGzOFvcpwCiOV6CnuKZfz0OI0oP3yQTMIncC858PBsX9Lg3
iklnLNyrkRNhnZIhNp6ekjp0Fc8Avh2cuGBEoxkGVb7LYGLQDYV1Bk3Ln8SbUBQ+
7yem/pGfPOwIWtXXzNXuXmkJHzHind8LGjXEpiC9RCfBNrvULJKFHmmJ9vvTpymW
KBn9DxG24TTDzaK6xjgf5GzprP3zaVXsBrHMw2tBhXLfjcBFPdajM/eSPRHXOOIx
Zx2zFjaXcntYaZOdZNaKQITQV++hsfw8nLdF0eiyrhuaWFqN2yuhEdue5LAqwyl6
Et1VJ8giBplm3AGNVapkN5VJ8OGZ/68TxDFqR/fIhipZsw96iXCAqsLFOkB4h4Fh
dNQi043wZdSnAZC0PCdI9cIUtGrYYWLKUUusfXb9N3M7NXrxbY9EIzaM9SHeFOMs
1t9AWfdzyGWmKozBQEIPmhi4TjhqdCDtGaRi9jy/BPJ7njyiyr4/7hBHBY3ulhj8
PGWoeDArY1uC1d8OYg0qk6I6GTg4/41k//trxzmmbjk8wMBgzYzAV3zQu5psDpHI
I6hpTUUR3p6hbtFV5cX52zC4iU0be611Sb9CLwmPlNN8zZgOwqRsIGSB5QkrFcVv
xZFm1v/1t/g++VGWYLNVPngQi/zvPcZrnPH9B15l08RNoScRpFDMqL4e/Z5Lp3e3
ORNkpTnY2BtftwSb9Nkl8bJtwJ7bwK40LlaQEXHuM69kAFL+W1lzECot5J7gDzCe
CJNBJZFMFzY8zpynlK8+nzWLFohjkytuticDkhMLIcHPbWq2VByNMlSFit2ZbcUi
ssMAoJ1mIdP/W2blGhvwDE4jd0ap6bEw9MgRnxMd7PiILivi+5N/zI3kWnwM1xog
4igrBQmIcK4Kcm8cJaC+tX6fIK6cAbgiebQ5JFxjDBRaOPcAW9CCzBoi4qAQ3cq3
NAlnJo9aEq89hid6/0F8aR06Iiaqg/NQhbtduN2y66MyH8YsqWyQYBQvbqGGleXM
RuPx2/cgcnzWARH+Ez9jdscLid7Pjgz2XTlY9vFdXI+g/wYa9KYkhvT1TczZPoei
bAf7M7DnKgO2wi6oy7xB/8+twScztVZomzdCpd/CTlBnyMnWnmSOmiHFnksHr1IP
EmPuPs/+DIaC8BsZ+NDqt+eNbYD+0W76oqLyGGFplv49fBM0/6qYKND/yYdLt6ij
BZ9t+a+Uk6YKUnZX/guIaOI6MMvbGZ7vIdkFaJCHDrvty7RwOlx0mZydAFWLCacy
fDm7W14NRxYOjOY3fXmC8Q7xajjVGk13IU3MM/8mTQshaqYFEQgKagHWccjINqKV
OSe1EWzUooyN3CU+rpiV7cLzhm0mrHrc6IdRfD2iml79zcM/ctNdryvsOzQHt0AF
E8HfeG2oTYC0MqFwKTeIR+dfZXGJWHnkdZyLmtlNQSNn7v6VyZxcVTK6JZVXSdOU
ahTRT4CKq+Loeq8rVA2+AhfzDIYjre3hrpR0/Pxz0n8vWh5pD9LcK+pqgYTMsYqf
bmzRIyABwn2yY1c7VL3kVNMG0MEPkRibWbQsDytTxXO0DithF7lrY9hJpXF+TyEx
3Hsrt4eolEqg5ay71xWa/Q8lmA/hqy+a4FGa3AK4OdYqyo149k4p955IMT7vhKzB
DM9NzzdZSONrAcyEMmFnbZJX27P6p2B0mNmgoDiLlMkcY3DxCjXK6NZJxOH2ticq
g9aaK73z7+5ybxgnyv5E0am+K/yBZFlCLtwcsSY8raYrOCDkDjh3PBPdR7KBuZNO
XG45TmBJc3gYgtb16fSs92Q2FvMhny9GcSI3wTMJRtqMEWijpyj3frXcaDmzDvbo
wkT2fdpVkO+0IVbhvMayYYVZoLVCPsW5AyfU7tbnm94j7RBsng0okfuZuIYE+p1e
GRlKFLyvkucWRYF0qw/5p7i231EpqIILG9+aNyUIZrI8qop0qwYqDSuME/kQUPXq
AFcUDs7i1JEaYAGia3h4ZMboP2hmrKaDWO9fo7YXTNFD8GoOCsHYENVMu9z6Zqal
7vsiKpaz/dTk4XSwfrtdCc3UOK6FS762uEopV4P7N9ftRKakRF6YnlGJiRVJG4+T
eZ5qlzCAdBu5CLJa2pVTu7fcmndIS0D1QTjtOvc0wiWw4QVW1/gmOKzvviblGgCZ
qQQNgWimWdFvaPFnbysBwyPRT4AJqxI9DdUjo7hRKLef06HOQbR28jJHQXkM6Vl1
/of+48rvCDqb1cEopR59tkxQFRGX+3XzvVjuHTAeCB5jien3zS2jvfSB2d/J0sA5
ot8Sh1mdDcJvuY1qYCN/cbIK/fYAq83pP2ZQYeJT6JbMqbiZYllnhvr5DrQ0MTdY
P0rtWiahrlUVxb23WToTpb/UbNPqub9h1f4AFpT0dXdflWYhyfsS+4V1oOShPc/w
d/2oYw6l0iGDeY3LpCJ6IK0dsE4z9BFt8QJH849Ju/VkHJEpe/RPDjuyyAvllq2r
clynGSiHq3xxmfjr7GQpllSD16gaqzUZZz5AeW8+MLYCBd/OeW/E7zkMb7f7CV28
gmMBcfG0HRTV4tJdZGVuOKqLrUrpLWXBnubF0MRjoID3Ui6KZNVz9o4uuUFzJ+iN
3ziocprjj91Ek+5XvHHyJzUY76SyIiYo8VKqbcRlL3r9bDal/r6AkJlaxh/4o48n
fRgntpdcaK+n4cf22xN+vc8BSlSvGQ3v3zqQX9VifH6XUyIDAvaXh+IEO/9YQQSb
6Nrtp6GLjc9iqNgJv+z7PH5MqBjJvANDAlTVwb8jB9WNMyaQJd+eiGC+cXskI+0k
ugmmHQOwopbmAP9AgKZWmUVQFezjV9le/vQAWextAZMvP+P52vJu7WjibIK0ehOT
Xzg81ROnjAhwklnOP96W7w2vpQ0hVD3NXanJWmJMEQ+2FK7XpZHR4yDN74dk1H0h
DCEhR7fL4yyHN1TSDfBpewcEDbpCDWe5K3DL1IzzHpz9Um2MczTD02sOKXvE6Sfm
UWzLFImegu4B5bdCQLBiQ1x1vRIX92Jz87YBsJIQn6Pf9pPmf1BSqDpdfP52ATtl
9fJKtmahN4ySHrO4OWYwUQbDNFYhQqTI/GGqrhxBfzjgogfUexUZRuTypob5nZh8
OTfIlFe2wL5fytuEPtv3ShcS37OQ9wQrHvhzD++xtbDSceb76kTYpstlGdcNDANf
A8MgXqVY8Dc90aX2uy5+VEQSdPCAbgr5DscpKwCzkRRuHXRhge4z4piCWUlNu4T6
NNU+h8YruYFVJ6lWLKnkzLBFlcnPylSNIl50BByT5Q+rXAJfPHXT+fLP8Nj08IWB
G0+Ei4HmzB1qZh/TXpEDysHTC9cwxDQ2V5zmFAsAQoE5g2zxKPMiVMc9+0ORCh+o
/f9UMSEgEUgpy/jQxBb+rJLfAbcAvbOlB4cDAjrEW+p9LaGNgPvTYUsky5mtsZ8L
tLuOir43F9psZEJs0hL7wkRKuwbFLtaganKRQGtIKjWpYGvV1cDokPs5aVaTdtZP
Je0y163y37PYJexN9JS3u0cV2J+WbJCwjbHC9/MIxWYZ9gdrZWbk+waPekVkPU2n
vfHWyga7wZeCVcYse9c7qeS0LgpxBdMHaYxQIIO2Xbsoac2i+nFZiRwulMSVH1s4
GjlxdgYAnxYzcADpoQfFNRGGf0JWBWhOsQMYPGYlEhNsiq8jFGuI7uVdZMLc0A5w
lJBCE2JHENmfR1an4EWl76TTl50y5mfsk+/LwV5+pV3uBQrkiCRDadcxn4f1q9RI
calPaZwVHaVdSiTXdY7LRRAbUFPPBdF8eO36s0VHApuvSxfMMSZDOnd6k4ArGiIT
I2enKFEeOS36QPQW3TwQ2naKnBTCyfLaa1Wp2DeikSpnVSHu9sC1T4pfyXBzYN2M
wQKoVt9hSAPMOs6Wg7rEaWdY/bWrqOF0fcIz3NFh8b4I8Nfj/oL0mpNdj5bZ9O6Q
bR395D3+y6A9BM7gCCjUFxFIFYFVHizxUQa5lc3RBYs6z+IrOg0KcngS+fXZ0cwH
A2r6ylPg3fydkPFm6tjueTKCaZgTLyN+46/LoQsjc4OMr9SPhdwSUm1VjEh+fO9z
iprPVguk9afH2CPUJRUG5WsA9Ig5n0PMR7NdDH+hKTYqT/+EDVl4BnXyZozkaXyG
XYec2Qi5/WX6yEbXw1ovA9OW4vU4Vae6Yma1rFiSt3CAnUKQi0wno7WP75sEv/j2
vyDAwprpqudnf5IXhrfBAkBqJd9epkufHbVGKpVjzb3zoLvYBHnQR5RwY/kXvz/o
L8bjhE6gnsho+uzaDh8wZnniltVJTwR9tlZhvKFht3axINi8p9p4vqTefD76BHVH
HaDPvb5o58+GTSJR6UkNrX6rknwCj+wbaNplrlaPWPYW/x/GgZZ9l/75rhgB14NO
3nVxpLZb4LGsmH1TwPTg049Gd+kd4wMEtpK/euZgK2/ZhzGJDvVGpQKH3wct+0rR
Ut9X4wQZSZcBX4y3+/xkki9lFo98RLKH/Gd4rleC5eE9Fqe4a6yMiIAgxCJoFdO1
52gxaCt2QGCcvB2TqMSgppkIUAZ9DMWpTSPlP9capc4nlVq1PalrfZlX5k36Kf04
qXKu+2d74yohEPhjqeeWZxszJ1168VDMa11jwmzbS4kRm0QiXgDGuxO6v50T6kHF
xGByBXKEeaCvGdBj9xDctSFSvCccIbTuElMa25Fhd4/rwUB9707edhE+ZlxCLB6n
N43y1lhClUTBdubgjJ+Tp3pbAb+geg8raYeP1P4DRBHgA81uKkSVsc9OjwJYJ74u
liDqzjv7GBbcsXgybe/OIL3UIw+mVsc1FRlCr0eLIPWkubPXAUauJbZu4np1akr7
/SbA7IKMxLpcenllueOl+vndW98KAHmyir8Be5BYM4cv5b3ROqG0SQ4/6Kjp8M8b
NJVkZzZMb4cbcqcCjbGka9O/FO61m/jQw4iozzzkbbTP/VA2zuoBzBiOb9XeaHJj
fp4UH/1zEEXX4VpuQT+yD5S/mWe+nOJNxzQKLyWuZh1kxhg/C9Ws/k+sF7cKhrY6
mld0OOaxyM3isuvQl/zvFS5RTgcLIIYyPvGTiNCh3r72HVGTDMIxU8deaoSTvnZ2
Ecq0Xs/7Ci5tyTaynu6vezmiuNF/IH4y1Q7koprFP8Qry1ez75xBpko5UQmmhIXk
ll5dyauZ6Ydqs6XsMQY9pTUZcHVLhT83+HqSrxtZcbnUwGIEWPKZ02rgozQddgP8
NI0R0Hpt4jWGIIekeGmf171DUivst6cnVJqGObnCTIW4jWjirMI58Q6M5oKPFzIB
Xz3qoTiNnYQ3BE7SfeNRGQ8YRtpbdvnZVgwDk9vcy20ep+yliHI0J3EmWmk6G08Y
n8JMziG37XX7RR5oKDU97Wh8Fn2iFgnTimStkmvhU8Mf9SlICPci4W27r+cspZwe
94553YPSAG+VWmGFMdgDe7rr+meaqVfXsOG9eMZqc4karwbD2PFqYDGfH7ABBZX/
Q7CZgisgiuvFd61XWUGoczCpCSrbwUtJ9aSXSu6pZ0hEl6pCRbOGg2YVlXDla5r1
4uREGSaULAHge+xEb/Qy5rNFQQfJExMjS4h83ksAWhHQjrzgdy5Ee2BzodaFjgpl
nFpo6iCbhObcQbcflpRbgMSZjz+7WpVtwvfyPIrMJb/wrNciG9i/R5IIE5uHkz/E
Caei/PIOtDTFel4bIy5xZCZflQbbmb4DCgLYEff38kwAJWdackYeKoAiDLjrw34C
6RzE6MXnHMXOUAKYFvohLZsGLkOUSq/jYhjBKlCAdrIiKW+WjKhtwf3gmopnsTEM
LwrLigmylMsp1EvAl9Ga+xcMzrHJGk77Ms4ue/CLyCwVHAGXkWqaZJt39TS4H+z6
ZP4hggnu6xJlXmzqylAOu1wxFNbZmC7OIDHXKVc0O6+C4j6RJ6rzSn1Nsxnw7+vF
DkSy63/eyaq7c6TrSfxtjCbqjEPUU6vjPNR9mXNHRJY8rwdNGr28ke33jHimBg/F
mVUpwZMi54niFA3s6AcnOB+J36ajrNJB10ujLjiyUyBS0a9MGeGfO9gCCHsm4CmC
fYxjnr5YWqBnC8mKs3UTA+YLTO6Q6ilSbjrwVcs8OWbpa4Jd1AsFU7i6P6wxfN7K
3zy1Ubho7BTNYC0mTsHxIH4nKaE1wR9M2Ssi2/ZBWzWvjFkkggbFuGGZbgzL7sMu
puC8VojjCf1RUZroxvkWCPTFt7luobf4cPK9KFXikoGB5YAWHIRb6i4QTsBdoDXq
A8TyWvqqowGcdJn6nqMM8rO4WKlW04toa/FA26nyvc6Xnr3wT2VDpePRDu7lEy3S
+0yYoLJATvhfvgLnUqJIGdC3MSoT4grJmdldX+QHVPddANp7R3GR6s/boTCGjKwV
Y3xmnbtrRVFwAIm+hey7wEoXS50HEGDIrRhNUc+roz9fQheQqs3QtlFVzAerOMx3
WK5XQSKLP0faKw4XEr30Hj1d9++/OS6SN98536poaz/eExCD9vgD/n7HQlz357qj
Kr9+0yviAClcsloocq5NYSGcYFrEHLvX8nlnSqq9dGT8y650OjgzP4+NF8Kf+OJM
VKx11L6XQgc2+KeUh7FL+SUurE9MfN3PrWI4lZBXQTiVLXMKsX+PThHd9AuJH2J9
rbfMpRN8WKXtR+2eVkz75npXKjGhHskvKKCFnC/tGYKz5sViZcBqRqy8Y1wdJe3U
ppKhJg/aYhFkkDf9cEQTrzbxlgzDURLRgDkm2wheHYo172glhJupx7P8PUnnBWtT
fzdr6+juU0p/nHSuTbT9LWl4XqxkKH0g4ER+yj8BGkzz2jeXWG/gr4gK4yJGpEiE
GGRkI5WjddYTN2UQffl7dnEG38cLuj7FQ51RsGeReR9y6yov/CBd53D/XyEEFDG4
gpC0D+vJTW5hQ5fnF14dGcmzHSLO80aC+tWFom66PyQ50zbzCX7sBQ9nf5ppG6fv
tAiSNxUH/yIVvrCQEkbGZjrAJOFZtZ96dS70yEqHSULIi7v5567x0blvHu47fx6h
+OhAQqmsF17OHgX+lQ1RP4zCYvQDCI2YXSG30KRNHySlGSvGrtGDhP7hC8z+MGIS
RSa2aoUDzRXRzOH75QIJetwzPln2DL0PjTKdXqpoL6tfAy2LYbHVtD51zOU8I5U5
YRvPiFqqQWtezn4la3OXJ4PovGOHjidDoyQ5QluwUxJJp4HJzwYq20e3pK1ncJIY
8dCYFPqAd1HVUHziFjBH/8wOn/V1rcEC7kj1CwJWukPwvf/OygmxLArlZPiZ/gYr
CnmrzlSGDbI9HRn24Cxr/bKNMX4aHf5yM4wIKwEixCxhF0teSv5uI+dQUgW4opJA
CEGq/yOIkuy+rm5P+IN1RM88g3dcK/P3pVXbIVP2zoMvCyphS2fk7zBeJ5PZc3pC
lWLOgui0gljOScHxi3erICRdSIkeo2nrrcUGHHNXcl5Dic2QbAJrkKmATVQEteEW
2jdnZd2P6aR+imxTOKuxp6uwwl+dvdVfkM+45dBu/HhXL5oNLLuHwlRg77ho90DN
IjMJgi/v4l/jZ25GT5JtIo1YkPiLTJhqZcyYTSyKIHkXMSuPhznRPoU0MRCaM7zU
WjksqVoP4W7rIxendtP0sl2T4VwubIDqdN7qG/XGl2IlHNgKp8dBD4BCIQhcUI46
0YGGE1TticfHWZjvGgd5yNwf31y0On/R0J0vAdG/jzyo/j2ELVzU8GhcthQcX5ra
RH15J1+aFRG46282J4goyPRAigOCuL8svq8KDvGjpedwj43g9Aez72fL1GUctQv4
keskeh9z30yhfhLYA8iiTXGJ4k6MHXRS9NopWI7CADR78yvoFiIM/aJWRdYdZxyB
/+wMamO1OCU5kNPaN96fGX8YoeAt5tEA1IpFrIJ07ee/vXbGx4MhbK5w+p3jLmnR
X/fGiMQtEqU9AEKxwW6IFmH64z5kRSvA1BtKAWM3bXSdflnG0XEDBBUL7W9sMH3N
T43SgBb0E0YmpsjRJEdonh/UrFT53l40SdgusHExXOluwumAwaSL7eJTVEY11eRU
XyetAfUKKmL6jFUysi1nRy/QmxS66nDeUik/4/ea8CjRfdUlbnGRXfTQP7U2vEhe
vuE57y46PWRuZnoSdm2YRKuNEr2ROCA2OT1UPuhMys60238YWAb7ArGpWzBFPS55
XMW3XOmqnlIQ+XvZfrDlkwbNtXXRCVSrxRcqrUtU83YtfRGVnO9YGKbLkyt/GowA
en0XlL9NzV/FU4d3iVzERsVly9L/VXYw9laoTes8nFnu/pE4Yg0sQ21TjsJUQbyb
S40t0APmYG0+bGzwZBVbCM8IpbfPTHDPN2UVT018pmh6qXfVpo5EwLj8iYJwgb0q
ZduHkRGrPW2AWJLHy2M4vuQhIKSq7jaHi+cUERGN3TAAH7BPAU6fQT1/tl/4QOaF
za383YZQZLrvHmsERza//HcBa/hj8gMijLij9w2jzjihYHcUQ6nx2hPB84/TjUzU
xia1iDCcK0H8eqs27ZMC8i2+8f+BAXU8tDtdAJ4wph7oXWr6D1+69nzARsOGmems
Zf6uKdlZ0N3KLcqmP71Eo/z7xlaDkEOih5cpyWAw/gXlV7ok3MWwHyVEDXiadiIo
V+rn0nvkAIqOa/HKe4pKXv7OVkKUrAkpQxq1P7qw70BiRZPMPZ/Y/gD7gCKKNGV9
oEiIKXWMpbKuWv44nEhoNQVe0w53uYNlzNYCuk8j86h6BdxczT6u936r+8p07VGZ
qJKxq0zV6gBi3Th8+bLwUMozTYCuZl5wpfBVVdbrVFl3fGNMEveglOqMi5EcaFuD
Bot6V4mxnik5aFPzoyDuqOPRsvWzfnRLRQdT4SmhX6Q2QxSwyBPdjdiDaj21DT44
CGayAxOADDkMx/T5n2Mlp4I1gUfdRK5p28W8fHrLsyzyiUQUfdBuQSwdUPtOzzTn
ttF9rbUcMX8FWGz2gmhT4l9jcBXZBrCtQzErAOWt9iK8mNK6qwFQP34sBnrItXXG
4VVhXsUlf6Z1/qTDx/pKdCbGb8tfd+gq2y13b1h4l+zTFHO5tXBWwo3x1Tl9gmPW
t3Pp08FBdjYEjJvC7qYf2LflFqKq8XtzGDxXwDuv2cEYCjGv3z3peET4jVnZwTYA
h/2tAYpuDXFmcZrztfNMKyojkdAWz0lTqC/D9VdAdeP6CPDHO0oE1kRltll1cBdk
iP64MWIZPCbOZqj77NN2gcH5dv1M8mIH2RhWheYcis+GWnMy0CEFaTUAWIl26uLA
SdgTV2W7oDfPLqs7m5JJvqDSDLQaY/ssNQKQzKxRCF0CP0R+SDvtHQytrdKvYUGR
ah7KHHKhpy17BOnu6eKqdR1lglaOl4fmV1CHkKc+4XHJ4Za3RXGcsJUVr8T5xyEK
0XiQNyi/V/rYyI5GgCmxxxf8ipyxQ5r42fO5NU56tyUARz7lvWglzcY6vw9wt7Jr
wOoomtNs23q6UyIL62XbYTnIa0AoUUOwYX98/uXHmF69aubCQEf0b25c7G6scSq4
gY21daDca/Ikja0NJqkTzqXVq7Vvy7RNE5jYdXtIN12vexrMMVm73eqamOObZ0uc
wquLkIMNmA0P3uf5SuGUsJVIgOZwu7b/vXwKKXg20iLhQ7uTLk+JBqegA04D/M3/
U03qZaBC8/JuNMxAoNZq6veQIR5bWklpprIxKKe6YJ4cFr3jiwia8Zo7X5rUPQmq
uZq0AzlcB8VPj+gjucDypp7+8CbXwvSEW4ZAEbhnTWdfjmaTOUVNP6g3LXXBRKFr
eQa3moBy06y0z2PbhoKrRM/Qw/GwXr7CqVBHxp7IwVglzMvCD09uiBFno7XqqYI0
K3QM+bvwEvG7u9trW4ywgkSNpbdh2XPcOp/jYuA9Z9MKu/DIBGYhcX2Xnj6Ct4oH
+qH2eRyEVCdK6e3n7ttBhfYpAVog3+jPNSX5rp0x2fnPCGYginxMDyDH22Nfxo4s
ncF2AoR39vO5kZaqF4HjYjreGYyq4CTJZYw218gVW/kr2q2hOhFUULCLOzwDKtFS
p5v4g68HP59lhOSgybZMMCoiqcJ8xAIWhDKtarW/+z/D8TR8MSjqM6WN9KSLOuPy
mwr8lKyI1kqsni9C0Nn/XR3VCzat8DwNDD7yqqsjPy+9Y7lJfAJzjLPYds60oVvW
BWKg3utuGS4kJOajHHIDIshUkvji660+UkKBDyySNBbAsXzZshzHOQLg5fq6r7oS
s/uyIk/y3SqGd+AOfClyJyNjY1kh48jiUItv8YWT8ECd3FqssRqBl0+n7FLuVomC
3+TssNNIcEOTpKSiX2Tn7bvd9i14bu8zsgFlW3WXhJRVV9XtnXsu7Oaa/EikfqqQ
xLKr3fd2K2r36CZh55BehhA15kqyWNWEmgEBjB4a72KaogRTgEdviT+f6jXCPBWh
Vn5vpDSZDCkLbQqM71anOxSLB1pU+E1ybLF0zyS9Xa8JuB5Py19wsIaW8n4dfFyD
tLGc7GIId3lzi31AYZwEN47IOAkEbYeqhc32j/DFggwRFdIUDndHFqZTm7lhWBu+
hf4LMADQRMXT+M2/fxFHppeB5x2drCfkLGsEndxnDWIbPvsMkd8284mhK1qhc9w0
F1RtmXCUV2rlcxfgeE9jAFhJfnG89T7GpMp6e6TXJ2IJ+dX5cJ1RNTNItJ6mlNbM
UKFX5Bq4PcKtU0DLAjO6oElTZqLqU8Ujd3Z8lIh8Ha16+Nk/PQqAa114UU/JsrP0
KBQW7FKbF0yvTioNJPg61wsQaF5WCpVmuKhBdis3WfSIQdvEoJ7HC+vsoA24h1BI
ufcRMYucOaZAwyI3edbpqvjn3H9EEb/M8ehv/k0AniC6sQeBj9OgkCDKBeRjaHe6
dEwWtRtPXLG6JhVT2p1d+XF6POVw6+aQQ5ePnvEcJBfoNHKuRwO6amv2CI6THpO2
ic1wHpmrH75qpECFjFSTYefRgV4pgFvRBjNU6E3wF9G7pdSJ53ejqnRFUTmXmOfB
COTQiFZ/an93ddDcfth5dfD7K3O2f4IGm3XIDSj3wMbEbkxozbrgDFohQ4l6cdy1
Ms0zjI56lrjQzAplO9vDUUZxSogQC58OqTzm5OUgTO3WdPMv4nPf4ZUzkdC39Cic
rzPUgbq0610a628O7fgFrkkHSsZDqp9KjxQ2y+db6kPF4uITaUyQMQX/R65zlygH
/wCuwaGf7GUoiyvHM7/rrMFnBbZEK+fXwYrLMnV/XH3Cqxk9qDWiHvkYK3Qle58E
kJQtD7J1bjgiIm5vou3+7WqYeFbJMEoU75otOZx44l1HcTYoa0ja+uFW/ksqSmLC
HEa78zgP0pnIbv1029LjVoQlmr3Qd4tu6dSz13//3Ecyaa+vHlaJi0fFlTZnqP2J
4Z4TC6XZbL++MN5y3l/1zs4RGzbEHlVlEllKxPHpHrj8N/C0MSD/obBLyPYjmu1r
jq0QN45e/TnGuj6WmeQyCNSg1Dt40mpVL9xuwKVbuT5E/JpVSdgcwNSM1lFx+HaP
+8VphYdLswI77m9oVSzAqu9eI8gBJtJx8OFZBMuQ+XEg+pZn4d/t0mrAp8cYfoJs
n7BRzV37pdspwHh7cpFi6cV6UqVzsYoEQvUkSGCYZys/e+fKdl9iNZNkWkk6sDVq
y1zhd6BXck332xRExyhZrgPst/gJp4y6pgk3Y4yhWUXnWcIOO2YrCnUIMhEfAlkR
+gk5fnAiaqmBE1eomAlVK22ZCZ7T/KB+B0BfBnPd3uF8W4Nm11tA/hUSEQnA82ia
oLv9baJymctdVNBfIYTiuLux0Ai+KYs5+osWmv19KzlYSMXZo5KQwNBzjLEb2lCO
YdLKYrPkz4SopqNfgZ0mbG4bKsjFHI4TxORXKTR4vvV1gsjt0pvKNc5Drn+CtSW9
r+P3sH+vViQ9O4+eq9low2U7IQLQQluVR6fiDFJxIJNJtcWrtaSdo31O9JkEvjOl
As1zLq11Rxs1w4PRuRlYHxRgv3dJc2wWSvLkdaiWDOOnF55oOv2XGQFe58tq8cwS
AIAzClaoOVPIEEgpqTG8MjvucPPKoCH45vulWV/HCm6UCZRKoqTRchd1OoDOr0PW
8b5BWXEjve6w1JIme4JHAFzZQXgnb2sjlJ89nAqUdoaqEDbzGxTSc4MqB+rixzoH
hZDWS4B4fFxzZcl5Ezbeqd3Zdi2PSN1nC4win92B4AsP+hkBkPbog9K2/dRZjhCg
ZlD8ATN/hwk1RXlURDXTb0JpHp9Sw30y7WNZmC3jnA7mttAP8UpdQumVzqioPS5u
MApOIw+G/Z8WGp3q02Lfa9qfzqvQ1wFvNoAikISErxRG42GZ4d7oG5NOOSf2XVbm
L73HH8GzmSdtITGQ1coz5w/h2UUAqj5NVjqwl8NVG/EBo9fSSTE+pAiXn8PUA6J7
E+bi7WRkhoyCy6rLQsk1J8iZY4hSF2VEl/6uO593drThCPMrL57ZmlJOL/twBbjE
H3zMIVdzwdU531XttMtiv582niCKEsIZSfp99Uj7TzUmqgokmbUQ+ZAv7VE0YqA4
jhnV0/QC4f2WpZnDkj2XGu4Av4zAtTJtAnaBwY6zl6tCKa1Gc9gOe2y5k2JJLubx
6iDioJZq4W1QEHCd7J82qMDvwjvLpbd1p61o4YE2T9yZQaNXOiQHKeECw5Thn9O7
YgQWayvl9rTvYxJlp1nHkRCBicPhH5pYDUM0C/aJA8LvkfEtnFfM2F1K0DZ8GJlf
yQs62XQkVRMtHkJYZV6Bm2I426YKuJn1FOkwt5atMZU1UvhLpB4kLo8Yrz9SVRcU
zwuP+qxgplIqs3YZ6U6aCumT6VLUzQh1tR/pOKxdeN8Z/OEhmmLCtyyNeYJn8WC5
cGthRkI6AynbuoZKuxqsD/ojqO7Fg18esbDFHiqHY6u9tfT1C8MkwX5VRmCovg+i
iFrNxwVXYkdoA4PPIbeh+umKeod6ozIaJjk2lgb77J2ApFxpI0DUWsXK3AUrI3I8
gydWf4HW1yhMtD2RHrQu8fuA1/VhGIYORgsKt134c88xoxm/C930wlvJ3n4Cp8Sb
980nYi6T9bfd9VGD+hGC+eGYs1aLcQhCl5pbUlaQ5KLZNpa6JCROCPj1ggJGvMd2
L+5kOlxciu3BlMnyN35xf3bRwuA5OSXj6vggWv0R76VHiKVTD84u35/XMO8VdQAY
uUqvk0Sjxy5eYnc/+OntBqoMw7ZVyL+SPAPnF8NIz/4y2DXt6+4LbuOYkZ+0rsOu
t2Of4dlKRrydBFa2iZ8ixW79ClUEEctPacm6Mh4AIH2lPMwmn5wTFdAe3w+bIVdw
MC57LVXxzJM5rfL9Q3GHU3hWFr4csMRzRTx3uMSjnYBZFWqjjuQoHKdZ4jDX8m70
LRHOGILNuzu2lgDf9EHm6ABHJa0go5oBgAxwD561UtkqeOnvyynmghr5iLxld4xK
Lgm8qzAcmab+OUjneUcKQYis3CtekkJ3gRS3O3m+qSRYHHC+vebqt5f3s3VgWmtZ
SHTUacpm0E3Shv129wca1lDSc8IO+QxZM8FrJUzG5dkcb8DQ2ksebNbMPzd23Ipo
9vw3aoficsV4QaWVYx+NHUrCNcwdmwZI5fSVbD45RxE9n4mmIsMteWOUnlEWCmiz
67G3DVNuw4gAkzf+cjptvNSkPCUgAvI5wo3ONbGFG/bzQi+rlMfc+nbs3CTVxWGY
p0AI5r0a0vbE8KFJAjA/T/dvgznTKPrdPOwUDZ+12frlHFJdv57my7+r3IFS/SRk
+cO8QyyZyQM1iuNkU9lFQSFnoNi0VHBisFDqn4LzeBBNEnIf7rCAMIKZhEkgO/hE
3S+wXT+i3ZmM6U66b25ifpdfAEYDwleydxTDNsf1sosqSuEH5JN+DNRwhGsGzNBF
lHHfxjtuBP2gI/nwJ+EYufpIQLQeC2+H/tfMbAcOtu1fDGk18v0dH/UNLN7JMjr0
EQn5pOaCG0T5JAnzbo9xCUOY1ulYcxwN6zcK5FRhDNrOzWrgxmtOQnVBghgNucTj
rrLHj/oQGEIx31sMOHGd85G7SjpH84IL7Aky0mNbbFnSql/Cy4rc355YcaIggoXz
GTynSPzFAAZcGUMPt8zCnja6SgRrCTOdriKmwL1gwYPzJOZmd2D5fYFTua68uqAr
eAnYdNWOkHcmrP+Bb/GSGgoTtA2mm92oYAvCAI1lbjRj0KxfTJt/fHSL0NhXts81
yOHbNzL+vLl7V6NvUm9VMu6XtRGCHeLhL+WhTvYyzO8MBCfDKRHUTa5hkX20WyJk
4/KjrrWfB1ScK4ay4L20EQVJKrM30dYE9F13sfSX046N3idaTHcbeYb/yNlxkwtU
z94G5llwDVk5bXji7du3PQXKQrspF6qUGxdNWWG5tGrK4ztcbp2cCpuowLPw2ptg
i+sk/Z8dLFtrsUJjPOu9YFHxn9U2eJdS6hDN3QM0Xc1V6MwLDfqlSgMjRx3L2oKR
AI0o9O/g0Kj4AbtYDOOJuZd1kRAeMwINYKlRNXZEcPSmQePHyKhCgoD3KsR0KUgm
6rIlxxnLpQZb161cIpPjGieTgGhRdrxbLpq9JIsZykaPUWbPWiT8ainqEJXtWKgq
lnBQhiKUKF7xI4W8fb7bxCFf6Bd/S1fn7ImoijQEY00dYkxelmZYUIZhcqfKuzQz
MFyrehNDZROQtBbe1VS5oCP0pAJO5pUeDttDaOcpz5Z6CmbRtKpKsoaJJ5jPgmXy
zf7jrhXaKJPnWInVVxDoxSGEEydFE+vn2WfdOZOnV6OlpZ2so/Dgq2gDR1Kpj9lY
WjbeauSNcrvo2gZAq4mhA3je4+qdtHdqGlIr7W9H16vssOl9cJ1h+qk96fDKz76d
mcrsyyYxoSmylvC5dGp0QyXMD68cnnLn1/FNzgaHI82vLjhyXQf9FfZOalApAIIH
sM2t/bcoXC60G3yZWUPIyv7c05CwTvekz/24jIkXd4M8TX2z8R1MToNzhBMKDkkJ
Rmcjtb0bBn1848v0YSof1UNXfZLy00jcNYdmfkx2IqWCgwGCMYozWlqQ1LtbwStS
T/9kzJ4Cf+KMStwLvi3IGM4blGqUiUJb/hGBBkcfyTMnHD6wa7e71JTIxoKBLFGq
CDQ/g5xEpBQPJcqYOryLy9bdgJDDyN+DnaTntN/Cz0lHkxOKzKbvUIn+CYtM5R+M
HVMRwqxpY7L0KchNyyYEZkMH9yVzrENXzy9TaJAFSuXrdoLBlUYlHHNhJFo14iFn
2ExEr2nXLtYO52ryFy6c0c6dXqDitKDcN9h9dd4rLSZbgnPGOYaV3xYAfadRi2Qm
KeCG5QOLAzi3hvpqTFwV9DQqYE064heukAtNJRM6QnE7YWTRszWi8MiEcvJkEIfF
vPDtcRrj2Zi+LmOv+UZTm/TdKnCc2oPUtYB02diG0Y8LIskm63hbcJejZv0H4QnK
11YBNtUvo57sVnfyBkKw+MEgTNTff15Pion5LbDGvq6NXqvkgn9TpPa3nwgvf26n
s2BchQtDd07odJFZyGMEGbPyf3Yb7MPU4gqdAUwNNDWCUdo02sRPt93586Rs8efK
06NFHUdo/3Yf8ZLvmKkexqMGI0i5+MbXWWYMX8eAgCU/F0VNqK3bFQxz0Evx1aAT
G7xzj4qmFdVeY5JfeFBg4nm4RZ+n1L11h9aQB+FYZH505d3rKXX+KwpEL/sH7uYK
1X7i+PrOTanc5QOHAwLeyYtTx/SI7vIaU/ll4FxxGkxU0hU9fmLq7tcHAXdqmE0D
jVYM5S0lzdBE++MjDUqwlnB8baEH7eeHpWgvfQnbxSBkLzAN0BVGQlBfwc9ab6CJ
l1pmkE55pYEDqvuJtZ81Jy0KegU9pEg0njPeDzV1iKjIibaBS9Isctybf2sbavXj
r9TGm1TREEp9djlR6FlVEfcHOJ1GnCpamLuA7L95VoVSkzCROmmClZo6fr3cwkUs
+pj2469KAoak4mXWd2W2yTc5lvFr4DjSOvuYVpcmUvpCMtAgFPICUyLhdr31XKTx
HVK9KvepNSpmQEXgZTJlwrCZ3TR7KRjLoU/Baf4+67BK4pVDdtL1QFZyVQgS8Pcd
VVCKeIBUXtrj33zmy1PSTYn1/PWTgvup5NT+cfMGwEnHQbCXe4c4G+4Ye9+bDOkh
j7Lbl/VO+j/Sc2JUzF7EmA0tQnV8Q8d3ve2lhNud2r0WVEoUfxV2p2OFRAw9PC0s
ugVR2butWW9gfn+Z7FeIF9QR9YtRoPuVHVAP56yMJKZJWXzQ4afk3gr81k+k7k1z
dNS8MH7DUE5ReswCU1NLgblNSGg2WNDXsrgUhN8tql/rD1GXkmiSFEljdnGcgjik
9GWTy6ph8dCnsu9jOF88SqLzZQJFd421NEMKDSCtgoLLjy9NynQdOq12QHwWw/pA
As1ZgfCHFGTMKnrnqz5BXKSacC5oYhm4cqa/qlGVqWBZxhbOtKhy56H4ew/wXBnP
ciCT26HjcjTuQJpWFyYYZvS338pdO9nkS95jDm9D7ujDATu+bpBvpyx/U91GLwlx
8/03C7pY9CKEhEP5lKOsJUyUgdngNcy3pdKeY01sgla1jFpTYBoMgGbm4yTG8k+p
4xy+FcC3XUgP2jCfRizT85aOev0BvJSCCnA6rIigjM4HKUYQZfv9+TznZHHrr7P2
MVwKpO4qs+XqzPmmLt3Phgi9jCvdZh/p/agyo4O4bT8dhcEfri9xkeDNmYMWTHj9
aJWaPTI5OCpWzP4wROAbgGTofxZxfOJxmtYtaMpSPidxBtYc6omopi+Oy8TkuIhK
pMl/oBzEcU32FiIzXPx5ys2/SopKj9Vm40414lGIw/t/krYKTrwDevYe2AGikSMX
wB8M7tqyrQiTWi78vvPe/Uk5ZMm8q49hsUdNlNmP+2hSFnpx30E30H6O9nzfWrda
SUdanQ5C+pB90UD7KLSm4/M5dNIi0gC9OrIZ8iW8LYuNAXfSgHvzuRDmQ+u71TVk
H9MWpujapslPSDykDJYqHA+6/EKbIwaqMI0cd+LlXoBkziK2EsDA91x2hcVJxlvo
3RlPWH7TIIf8VnyK8LMdTtfBsT9Jg6stjsCDEiGN9qgkOKzDHCfG7ZtUZbubZNPC
kqp1bGKLtpPkU2DiQZXlgjunn39cN2MxHTXQk9gqdkqzfs/tLOpqK0C117YZAbfU
p9h0udF128jTGeieW0M7bJGA3PSVCulLMPMrsbDnYDgAbmWt2RErUuzQgs0DRuK0
DmKB+cQNrX5jLid44GQvTrLfnLYp+/3606+rmUzwfKEWC6sBAjKTRi/HP5NphXkQ
x9m3prhG4uzvCuBdevLGpeoj0GRkPYDbBw0qbDZDBOGJFStHk4nP6cT3rLVOWDaq
0oOCA28Bn4ChTyMuJ1GcuidKvBEGlwRE46S0PTMgtra+jL6Bx7uPgXx8T2r38o+D
1hiq79qmfnM8Eclg5KtgChtv/zUpjyRA/fMBoxNuw7UQMmksRx7t/rSo28X0hLRX
bxSyV0fy7AVdKa21Phf0AJ4YNW1QnGnfCWUYf5XOI1BMkgcM1OTGalApyvbwaxyR
6HboI4WrlB9UCWewYnZuCvZCdMgqZ39upnRx/BB943bWl7cOLUYqDNy4v6vSOhGY
fQR4QQvoJokDZ8h7E2Eg31ugLA6ByqAXr1sewhMuFaChiEYJNSEr54s7uitvffSP
sG/GdO2GWVCDkHOxUpmH5fRWzGU6doFClZAQZytns2LS/QOdl2XLf/LAjRTzZNAC
HBAPdfOCzWt7Ganuh0bEY5rAEMNGJo/an0gPjQ1Ea7AdLHOhqgbIqmF684I+ytE5
YSxhkccW3gSfbPPpU5oM6xqjzWg4Cakzpv/05OvI3hG/sL0fNoHMPivJMf6VD0st
TWnVmFCEjOMII/SzpxVg8RiczuEZ3u55k9DzufyceJG5WuJyzGZVS1f+9yKwqt6U
3Stpm+0EouKw40YMgwY1jbrEcXGc/D8amrROJOBh3fN9d5MGuAmkv0xU0S3CJjdm
Imf5Sit+AQElCOR9alNgmjZP/PopvZc3tnC31GUiQj7eJudu66Oa1lh2E6WNNIyy
B+cxWsnvTW0r5zNG5OGJMLcMjgwUVPLdk+mALkMqbqCydENocE9qm2oFJ7au8HO9
ITXJWQIYAbQ5NqDOTYpMr6d720e4doQYWVZBnfTJNLLQJ/3Lmxzzo+3Qo1iU4S/+
Dh4aIjNa9OvLNhb+qcmfK/aScjQp59mGJT40IiJjDsa8GjSlYrll089xAxEa9ICI
WJD+24eLvsjo2KZ18cnNwl5J8qunnQhrpcFf6qnM6D6MtJy9+w2ffq4+SfpBudKC
x+K+wyPTgZUiBvgjVaD/nsRKJppHgUmOKZRkjmJB8rZVpCn5cL5R0Jf8wXXGWZU4
H7r0Iq5jODxqIWFdJImkWrIbOPgBeGKR9pHCmBx0SuuislSqjPNtNE4l3FFYDZH9
Iimp7jFyNZtQvaQFnZUQ88lsKc0Qviw5Kc7KIPuosyV8fnyT0TvTDNucSrO/QCV4
JqFSmYH/YbxwFMPH7JB87fqjd1Ebau6zd1c3OxGh+yIouQbNhHrS91VeQ8pdERtl
cD3fs+J2jDCUikaMFAgEN9PPdAMeT+IAhNT3WtTDzglOfSOQhrvAl93DLzfkKS+K
gZOTkkO/6j1vR47INBqjVBeO+IV6ZqE8eXlJMPBBsBDgnylTsQD80D7x4AGP9ypd
2dsS7jIMQayz2xTG7vm0TcVTkBTJXi6kcgXBT1GjT/IGO1I91N/A3hhxKAE9aoUd
FLQ2pm8cJ0gv9lTfc0fTJElT/Qr8HsrC87oQs3/zarbaDIujw+6EBewUw190mc8g
RwwmsXUKlo/oOY7LWXGgZahh15NQgHz7DPJBZodU5TPSaZYJ0DSH9RJ8RGeSqZqW
as9AVdEFvR8LWbqkcNyAkFmCndSXEXszGtrEqrNsgn8DnZq8B9szPWknXLGWm+J4
SL1GVw21WvAgdLXiRG0IGnti8to3Nqo0DQi+/+6UBXtG8pMj5htd1CgJJABxRQnq
jPkH56UmMbTPqLYFbsbtUDFxaNmETlHTOO9pVgCUq7pq8Pw6ajR+6z7f4fPQwBVE
fZAgzPGA87E3B0B1sWVv7gEwEH99HkLk/5xPUCvlbH0VAADzfKDhW7Xs7SKQ7f2w
rWH3BLdpfOYhPiIPXpasqcO6DjfVptv+g/zJUj4KOwZ76BFU9sBs6x8IVBM2G/tT
s/oRk8Pr6RtdLd4qIk6mNUhPqN1A+inRPZsCSkzIoEu0J0hfYEcr2CjmcMl6HOIJ
5xJZkxy2Dq2Xwq0RYEM5FRhWldCUpFFmplyA4JH5wmH0duYz9wQqaLw3ZDVCuM3P
NVCsfFyJnyzYmffsK7utfEhSUedpZpWWl3MUoywqfQLB+07uneNOeHquhHLp28ys
jwlFAcSzKyqSr1omppDkrnnwdpOhfer0EPaa7mTRpkXurApcrhlP+JdVrrvFRPOH
uubSMGK6MKog5Lx6HKGrQ2R6nyaQDQS9AO3IkMlFw0TT1mf1UEhG8Gfxr9xDNmZR
mN7ZPpjvNqJ8XQCaWMULEzo7NbFgKoRGfSde3Je2QVLTupKuUn8et8BuGqI3/+/Z
zhvgLFCJ/lDu438TXJIMs/UMmVtGQrcRro9Yw+mefVxxp8VQ2oElDvDXbHslwVxV
t9D7b3byazW8v9Bvbj0T7mB7Pm+S9T2p0ZFxjprQ2DHW1GMxyz0Yaf9DnQHWp2Uc
nOaIKaojnoNqQpuzZWSMY1rFsUbdktbkBumZkTTEEzUKWC3zr3AbUwfYnHoA4YLq
x0NnfAT8gsSkiAZ/eVIeCmILfQITlBf5fvQ31SiCRpWfbBgJFS6bRUBNVo9tdxHT
LVuGwuIu1au/NG7hopAEgmmeStfa2gZqf6zo8jdI6XjVmwLtFEQhbPrVt/hT/XY2
lpixmZMfI9uVC1Zu74xN+NF8gCC8R30tQKPLg0lnfgrFoPAlPzPcnq/voQIrRNrx
ovjE+z7KsfqJ9qRH0bb0pWk+v+eruLtrL6bI66Gwly+DeSzFbpHT/hEf+FtceRw4
BD58kgc3F52DuXQhdnzA7D9SHmus/wgQPDu+bqaR/Stn/SDSs6TxnVbCpW+J6XHn
46FAYJTh7KaZ0vZltXFcFmB3T+P8i/47NgW+RiXktbligu75OuyKQ+0zjX1E0eQ5
VenKS1YXphQehuDdiVPVzOEw8UC5oqBBBFimviH5g/Ad3szNdSFMKjl4WAFwUKdd
0puhzCqu/N7aC9Hjowyd8FoYm2a7+HIN8g3NlcSIlNN5infLjkD0UjTQTyHvARxa
KXZ5xs8uJsx4D2hK1HubxMpau9tUMXhrLWQSIXlTE+MCzWezDF5wTLITfNWp3thO
ZaYvtU6v8K81OrFWzWaU9AWGhmz4f2rTx/kqA55TqvzMnghkKAqojBLCW6d5uBHc
4r/GVk7TXvjrv6GVCHI1cr+Cdc9iIv1sM3p78OOT9qmRHim1+ZSwcBTFY1DDl0D5
1pwq8+BOUCzw53ckOLkPFwH+OXvJJW3k0XaJr5G/+V6Gwt3Ph4oNS/ErlAiH/Yxg
nLQKKC5RQz49Iw+lHBGBnWi4WjbnSqxY/ju2ciO0tcWavlpXW3sJNRQSZso+M/Wv
XXFBQsOH2U5MTZXPNgyku4HOW2TZ8Rdu30/r3MYTMmJz8VIYKqiyQw7IaSMSO3Qv
jIrjxPFq4kZRj7xE5wYzep0bUCeueU6a4+7dZ+K5UaeNeDyLyVZ+HEjCGVrDDvto
KOUVzY6RaNDWEVZXkSKFyaipgasnT3cBMCTfD6uQARoPVA4SRXxvdm+Snul3yyrm
I3tRzLh4ye10j0p1MiERkaQ9ajZsG0nebvWeNLWdmBgK/us+vEfS+GwPWomI7Ob9
b+vWrS8FO51yw6k1kfLobconGD+xYPOPp9+t+M3pGaEKvzNPAQCXs3+msnBdrfwr
tN8FNCvT7Abjri9stq6kXtxEaUYl902wVmUu9wm3chHRKHKbeq1+Ie7UlyqZFAW1
1PZ2Z24Vyn68TnuaHaq3tThrhkXZSuRy7H0zxknuaNkjGR3vnPd0ZPUTW06cWA0d
Wbk8XgN7Uk3iH/DZ83N8DTK///3dQSv+pLzH0D8rtrCtUnPJ0GNhDJDwIoAHi4Hb
8hKltMk+cRyFhz54wSarXlID9oqhpdknhhHwyVJ3nmbv22jMozOY2yWMIDfb2az5
f4em29GZpax5hCl3X8MBh05gXz24US6S3HkPjGMhvUc16j3Sg0N0UEI5zPBn3RhH
LQEJ1Iqs+j4hYEZbDDr4fkaKnSj5P6zZMoMwa6s2zNq9KZT0dng3rh+ijI02RLLx
Ty0+XYIaRG8dxwPYi+6MNldJH658JGtcbJuc5XczvWrhyb0Y3QQXQ9vB5LRTJwp2
PnC68xz2iob66CDIGPOa7yZrmyxXAq27lrDghxtbrCYwABQ5dFMcOOVg8/73PUeD
m8347sWMKKlkDp6EbDbw/seSMXmBXbN8gWwycf9iRxh8sSaxLVdF/rw0hSNM8RB7
Gwk6siKmjz0XoN0HQAYM7dDWqVmNRU4RJXhXz91xBVvhx55PHRU7C0CG1AG+nNT8
HiDLu3um7cB1Ol8EDfN+FqeLDaKizbrYtVUM2I6Pk+0jizSLz/gglfilwb2uMpw8
ir7wl8ouNHoKhoBNXBK/rLTohR15DjEUpaeHL9ZFYPVlHOs2UGNjOrQ5pCjmuSvx
ffJxipnhpETD3RwpDtVF7wSTIh/U8mLL8Zg2yBL2GKCY0D7jUsK4uNMV2BLTYasV
NDcvvm73bu8WyGhrx0WRsmdI1u+LNFUP/miX3U0h8Nx9ygm2Qj2+UDQsxfezPTBP
BaEz4OY0npV++XR0ctr9QCz3P4rTOMTYv0/s/j8YKYxrCrDVVM1bEXiJBqAjoBWn
rSOblPBUnZnQKFH66MvbDkqHnes2sRL4NyRIl7BRFLKPBY/rfzcByEDOaQIjvaAg
yVEJNPvDjycBdL9d669k4+hRnowGj13ZOJZHq8ByTr6K6FB+/pWTceOMIZICT+hh
Z7tthCRuOks7vu5tq3ZblrTzDFQEYaZ1hZqCXTZtx4xO2GAYbvvKUC77otB6SyHT
LZ4V2dM7IZMHRFRYc8gpqatWGsHr/TxP9UUeRWbvPFZ6VnxGaR9CtF9tdfgN8kgf
zR9pakKuZm8jdM4APlqbVfV6plMM8RDzhMkwOElsS2TMgG95Z3SwhvErrqPDeDv2
arYtdRKJl6js6i6DG1jzbZy0JKsYUurbDbU8JCamF2zbApm7APaK36H+aSfQFPAk
wCwztpgArvIMjcWJLnXuMx3Oi8eXw7fbS286PZq3cBnp6dcucRxy4srTXDbiT4bl
5SUsDkYPBGQ27OuhAe4GF2vu4zzFkTGEgrQX5R6AiP3YSXJgz6ex+1D5F7040O68
cz8ejLiTC0rbUFo8ew/Gp3BQksue73J5l8HoflmhRvOjD0aYFxw+QYLRhwY3fZSR
WIEAhM6KveFRo63PJ0r9eEsgIcMH1kW8l8Dje+1e/aR5QeEpcl05T5KndtPScZzS
jd//hORM4ER7QEdAX/FfJ9Hst6YiJ8cnmxP9O5HhGwulLZcndOWo2GJxcYYRnzTC
08ZawibXiE3ov+Km+I/oefeckeYtgWZT5vT3qmIFNW2Erkf+ifV9iVsseVrSBVl+
+AmgeoNnSX2SO5oW+MU3xVQ5FnFybd+ycyRGBU6SnMnDk9S+61rAR+7vHDiPnkXD
duT+xWFntsVjxeO/KNj6/zFOHARI/j97Xo5/xQNBwukyc3fKSXNUnbLr2Hh51Jdv
6VMf9+x8JBICC4sKqdaU6Nfc9xYyDIqGTLj49yHXB5acSTM4QoB7/Utsa3zaUh5x
4CBPz/tU8DFTOcvpBPR5NHO/6xaPVGKd5R4H6FHJgfrRSoXsuWOg8KXX89zwCVVK
wwu4z7KsUGAoeOEabIBscdAWQFrgIIDcHo7rTv+7ICAS3JBjg3zNvwmPqVmy5nGU
h66c9BYodpu9CaOiiyDYffzd5SfmHqbvi/LEKCwRMhXgCwV5grj27VN1apMj/O11
R66Xi6yjXi/Gm7yFvRsmSuX5kYOG2ez5ABcf8G2UhZTfmReYVGU4aczuK8KSh9UB
XA+gFWX98M2pz7tMyQL6A4R8jL0WyUjgJOZQkZ1W97OGbY7s/4s/7E/6f06cR7sf
6cM8EmfmlGXxam99nkb8rVWyqu4nWXwBqDFYff1rMy2l5dGpLEIbpvRacrf1XDSU
/hGvMKaI8QzRb8e6PahbRFif4l/31bUh4poebmBZHXHP9MA0xjsZfgJvgVCVlOSl
nh4NBkNB2hxtXgRogz8ZHB/BpPju+wolZDMlXqljIj+PqyloR3zlNq64+cVVYdP7
GU6mKE9s1MCd2NwkJ1RFtCddcGyCYjVZpjjKq2xSNY9GpN3YSfWZcrznmO0iLyf2
Hn6CgtS2ikw3o2ZVgU4pySLNyC7jWG77JWimTAwj3mBDu2HsQCC31g+juZROJG+k
cLl8KJcsnkGdpjJtvA1blbpXwCfaPSpgX4s5+JTeNPp9AU8irw13bG3ZaRqVGJaN
E9hu0umDxpEbBcvZ21p8UEYg+dcspWIqzeVGh17yNs2cvCVmRdqjZodM8BCXPsY9
WCPZ0NJqnlaiI6FbleQaDwpm8dI9WkbXdWeZTncYytMTvEhkCq0vkoc50SU5NFTq
aUWrdjUhHa31Ox0PbxxKsI7kp4oJ+tZ8WOxL6GOaSmNQ2jsaklL+cfhaKIzvvgre
Np+pAU+18kKT5BDdP+7uC1bi7vhdUyV+VwKhuFgyzj9ZGrK0r0Ww14CezohBREF1
3tvOou6wF1AmYfIqY8O5BqG5YURSwU74lebC1OyWc8sdXhENX03F6QYYLfYo1D9X
FbWCBTnCFcpQD9NgvKkEoKIAZQxOfVrR1245eiM+gL/bWkUYOB5hutLkW+tdgL24
tNVrfCQRRo33GywcZ4CoVNCzKT2OO+nU+/4AM8RB2IlukIt8W8tdc+yxTDi/BjkJ
+aQUbaHCnJKLAAJhaBgvfesTwPqlUSv7yvij8lbmpGf8AbTfu99tkjT5JsxQ3fx4
+qJRXpq9haghuoDrFwJU08Dxr1UDhr6luMJwPu2aXN+i7KOEk8eU7958IV7lyZ3c
bPkx4hCA2juezjoeXrbOYet5Yp7Erwc06o3gre6rEZOSbx6XHK+AXlDlW3ZuD8ML
dCueRNXnPtg1iF0wjq+6gsQOE4KGxmZolzXXjFsrHd6ENNK8FjB5wXG0iLEwfh8f
PHIFYH8AMOs7iArI9XvINhVTF8ETjxfuFeeIN7OE0a9/hAy7dB1SdrUS1clMitP0
TUxB9gJtmk8aEZDIc6MSPsyxXm4nYHBGA1H1EMt4M4ZM3Mr0IP7SCE4a2NALhYbi
EFOTlv4Z2N/1450I1Zurogi5eGnc/3J3tWAZEsvgg1RCg0Hp6a2qGKn2NCnsGPId
wD+Beah7i7IA5arF1GH6cRzPfRPYO6Mh8QEyrMOrZN4w9+Q3c9qVfXpQ6z2Qi74T
QBN3BqXfIUpW1uMxFPyU8a6sLnwaie/Az7sfJRX+qjuy6e6XFvHAeKDwYqpSlIGg
onJVVnZ6UiyvGeu1VXrj+kXWUi2Ij0QMNPYRnMlpTcSBWDM+LfdkC64YtMhxwb81
7+C55rhUWY2JgRfqk48WjszPn97NbcNRC0FYWkYeu2czZLMjQQPZdUp80S51A/3m
rP9bUwcm1SpDzIcgZXN2cmzk/gUPDVzHn9rBFKlQG4Vwqw9ez1hU1TFB049tEPoM
1F76xW4zWWYjhFQWFrWL2LUXzD1tTzhXxNWEm4R757Mu+XyoG+Ge452SvtgZgfRY
2YHiVD8epRykZLfrFgtwHMC2jvVwVbQjUMWtECejUArogcOOaz0fWj5T50rpu3nr
HpLRNh6/ifogt2m98VXZqDsdZ/UhQ8N+5jWPWvYTHd6kBYa278ypymNzP5lni/mN
FZRJOlCo7WOpI11AbHp3+wLZwoqEBVltGro6rT8n8/nasqjt1lqtEMELuzbiJ/c0
0UaMWqkaj1HHhzl9MVn20FXIy801Q1PWlIQXaRP6jZ1mtqhbQ13G4XL0ZCVCVMcG
+lrKGTV+r8aMo72V2gvNPqRPDW64CHFOFc0AWqOjKBpJrK0FNmpK/W1pzl3DKKao
KdWIQU5o8Z+oRzB0ru3kmqen1M90+CDWWAFIv37PRXwFiycWKj+bET8Q2HkBVTpQ
5Jgocguzu49wHFpHcv6I9fmfQelrmEvGfPp5UR0bzJCORbgqTPTbj1HL1ZVqMLo/
LN6JTFqWbZrtZ70tnJ+W5HplMlDvgs35ivQteMpGWCf0s7099oMn1I6h9mf+l8V9
/FooZHv9XLfaki8BKefMMgeYBqzrBMRupOJpr2sSxhUQLlEFw0C3EY7KK07qoVBs
hmvVXRd6roxCFV0Ud2IxenwffvbsWhwxBgvaW81ufRsD93izLu+rjUOHZtElAnRZ
0YCSJ6k0AGWYZf/sQrYF97HaCNOnApdforPRhpFvfNuluBBUIVSasUTFSWNlfnSJ
O/qLpOT4QHfR0cuUcUfcPCIiNXs6/fBAQvwtucMUJX5vU++JcSJPXaI2Y6Y8Hh9D
9BnTy/3TSTsE5NxfUMkWUSg9+xkwsYZhZ/LLfdfkAajBaBcTd1C0RHZNUvHJSTmM
p0XXdTQ1OVe7a6c4S6rfeYT/AiIuik/fXxf4ZnvdeYVty1rpVa14NcRuPncBj7En
9p9p2YwXNBMNrlEWNJOUX+ChyIdRV/JHhNz3QXnBQjgeHE5v+YyWG3KQLrB2ZHVD
VjrwTgYCCSxECFRu6HtWWhEkzeaZs4d1wMQKj4EkC9luRpKTfGrfnxnrrdRF6KCz
zZOS8v1/BD+6n03/50dZSD8E3Em6ErMcl1mahIffH3AKVE2Vls8L9UX+NcPONsnC
Gb5XqDuDpZv5vT5hqMC+iNFdgwLucEoDyi6tjGpIhaFbO31pAzH1JajcSvPh803H
vwUnn58xS8hqXp8ZP+UQJWvCglBKbOES/WN2LqHqrEp+t/qKs4y2M4yqjC8F6T5u
tSZrup1VptB7qqM8ckAyNTEZ7jFG3+QLvH/HIq/jHPVc5uQOJk+pKi2+I5l547dl
8kEGmCiXQ+PEpMoV6BF8vBoFV5sII43NmhLFXEjqLIiZ6H/1QbrUXfaRt2POxBkU
+aR8Y2lIy94+vvdBOvFGP3zNOT9iiEAgq0E4YPELHr07nIuqLhFm7Xm6LGdDGwzu
6IRrivaJdZsVgTD2pzYJsFmMC0JaSoZj82+ZzP1GlY69ye7vQoBb/3Go2Umfp9pT
JVB1Nv+1+xDpglXXLrpZpJNHiVzeIen7LDQlBWJNsSKszR5BpNipOJYx3d+CEq1m
EA+wwN3VoiJBmr+McyL1+noFsMArf8laCTIrrykJww2TaSAX2BnxF8dAYTgEPpzN
ZpgaVtl6X4HzfzfUNj8qLlT9sGcktsp2Z7P78lOGsYA/sISlDyp6agmS4yzvH2X5
zMu+44m1Ok04r/oui87dcjhRKGcdU7h5nyRmhwHL8eQJiCFM8q74Nlf9EN8BDAbV
N78/RnAS1vOxcqeIFDVycGk4+kUNuV/eCToZ52yjNwE3iIqgURDvUnu1H5MwZf4C
y4431bxNovdGimRmHqJsX2NMNZFh1a3xzqLvRfLIRqkr1Ya6F/bnr5qQR27m4AXd
tIOF7PgNuoLCrr4u+DLbl83VbenF3wVlj9aoleokz74GZz+g4pqiMbv5h2cT5uaw
+7vQEIjeIeRWVZKv8A3a58/j+vCU1I3xeNYDt1mckZGYfy24NEEa1ifpd0kOCkhc
xC/3YzzhO0pnnVfL8y3mv4J5oeLSOEhGOoFdLtGWl3gySpr7hdRsISbxgOA76fAg
IwnBOx7bRGSY7Ld6behtbIy2jR/EjJq4jQDfa4ip8EfLAQ0eWq5kOW4xGx3ArqxK
Gxy6MVhsHhKbPdep1/TXARlZvIdGN9UOzI4Z2H8aL6rtlFIf7z2AZeMgcGkUy8cy
ERmy0adsJLYnHThm7mRaqKWXYHr7LAZdb7OdjyrWKVHX2Lv2qY+ejnFVqCbAOvfi
QKWDIbVF4ff9/Bgf+1raeh6BXh5gcX+xsKdPVUf+Zwz8r6v/zg4ChFA4Z9vLGODC
P9gLOeU0WCzNK/IpNstLTEqHCPYpJghtqOW95YzRF1AVIcQZbrh6wj01kAMvdLCE
e+sdnWZANaQaCfhPlaw7mEyocfUF2mdR/XY5IgG57J7DFB7jvOYauP81bsjk1CTs
JZK8JyMK55NMObjpuofEthMuDrDc3rex+5MB08qQP81gvSzl0m2mwmvyd1DdbnxM
nZDon0R8o8HYhZRjUE5y0Ov//1DlZBP+Fu5UojoSOXz6tjWOOXcgOauv9LbF5RNQ
qNDUsvW39x3hHbMGebjOIlfkOZ4mq6k3LfTClIPUo6IVbN/vSQcuPYt+EAa2lMNN
rkO2TQxdgZrEwORkqJ9ecYLicZsRPSNblrCOEKNFyYDuqWW+mdWbN7GHbUAtdfax
DoTbsjlsGf4igaEDnyxf3jLLAbNRu/h18BqNzFQ04kcPeexlDQ/LgRj2+HEcEpyP
AdnhOGeCO6bLSKxX5KLmGDY8FrHOQzBd/auBB+OidD5bSQrLUPrhp59brlUxp4OB
nifSvur/TxkDl+BInXlhw6i/pYDLvNUe1CD72hUfdjwvT/iDDO5vu9whR/2QYRE+
Ob6gErr0AqaI4DDr5UxD/F1KWWVzvoxxNJ00PNcQ470cSZZZTJHOXMiPLzkBfSnb
h+VEi+JoqbuOzci4RxHPIMCeBpgzundDvwQRE6+QAfOBEqjEcDCFyL7lzmvdiVKG
204CJ1sJ3k261/SAUb8MKC/Rl9yAAxa+b4a1UFhe8kg5zQc3EFQRaYvov8uSwGSZ
stbgLwjNQC7oNHiX5T657gejf+g9Kn1VzRwfOBev+tW5yaleZky6ro7TI8snO8LN
ljzJaEsWtN4L26eJtKTXyyRB2meFJgYvGeLW1EfxRIIXIAPcq6OA2iFIdowQyVHV
8JZr0y0sfz94O7DIkaCObIn3sP7FiNokOkEXlymiPpkVJhqWI9PWKK9vIlGPjjsd
diV+OYcJ1P9lqlcVk1RUwzadSSn3rzrsloamWhP11/fkylPFh06sGoP7JYDdH+YZ
S+ZLHveH5N/FsFx2+bfwcnpILgD5Gn9I7FwVwdBftd9FAqFh9YHwEKrSg/r3uQlb
Ts6EsU3T/hcQCnqFL7O7Oa5p0CbOd0Nc2cYyNszspJV0fcdH0VmbOfKgmHtGSopv
qaALAok3V5keGvtdgo7LZLetc3WKV4T6pvB7uUajnCy/9MwmYabcWAHcBGcwxE+i
4vI8C+9TMQsgmO/yUuDBTQNmjOqHUsJYowAjivu8TS3XwaDIAfC0evG4YF5oSrCM
p2aUhpMJ7iLHMfAfrtdCTO8OPaZDGP/kLyA3hjzJT1NZABfTgoVod2Ab2VELsOP+
PHMOdV8L6QPSf0CmmUm8++TfF/5v04t64ZvWBsENoF2SqYVXcFVIHRhpiFK/mAqG
eB+G5mh+4hz/fOgNPFVg0C7RfmBmvmVkNsXGVISrMAVQAoGAGj2d2pcJXQIiPnau
D9890dlViwZUfSqsR3+UX66uleJtKY14kJ27sdjrSgN8nws/gQGM6d64H6iHwRZ3
TZhRVLXdzr8bX43QH3f6fo1kt2PIqsw6lsGmWni41g9eXg5E3pX6UYg8oI261bSq
YgPRD7aqdzERV+2Mw9O582h5r27OjTY+j4YmDFYczErSnNKep6gB/nKqTRWDqGA1
tuWWrWc5THFoSjoM7K8ksHOt+NLLgkbQhI7iGR2gDK+/5ohCUyMxxohOLEdtjbZy
hdiZUSpRBYMamRfH1o5WphEjYvtUMe+gRWAwfoV8AcM705LsXkPaxk8ypLkFV9Mz
WXAfjTbiMu5KCzgZIsk3/YI15Xp7BC7GbIeyI3RycU9BZTcbOrYI3pMAv/61mgww
6Si69ziJJcu1wHzj9D6r3Ojzu9w/+0I9d9XzbbK9TBYJgijBu6Aqn461xdPdbTkE
fX9WypBh6Qugi3DenlSy14MG/kNh/FiZT8eT0IYbJvvihhglVVHnIpp5wtImcdwJ
8qOneGk9pEKsx/3nUsj3zQ82k2L/yS//nyuEi65k8WM/FRwctnFOcJwQt0cFl7ZO
/wcWbSSGh38Bghc9TRJlMVOdMzw1pvzWQaYTVo7L/gdq3CR0i8zNRVIJ3xoVqexG
QLnFv2tTqF4k/P7Uwi9SA+J8MNUN7R7xHSdP4fqXAIEzAA1bvKkppf6Am3VjfFMV
7NOlAJ5Fdl6MQEbkBjKEduTREw0wXrHpvN6XjltqrRZO7jX7J4E0ur5wyYQUTIFG
RxTmqSehaQxa3ORDZAEz8/1qauiiy8feBJKUFujkk04FfVp4pOugl7GywW2PnKcd
M1G2kiCj14xaazj1zQyjweIkdDgeq3vKlfrpR3XvG4KlpAtGSGn5/EmjUr/CcJCg
2q31jWAn/rb8hEqi4th1k0g7uGFDK0vJaNm7G6X/rkX2su9uYsHu3Z6a9gO41ZpE
w38+IGGwThLoOBSscZo4frtyhPprqt6VrAYA3k8JlnCyqfj10l70381TSYEbeIrW
dKOkOeNSeYQen3ruYQY4f5EJ/Tv4yt2Dzhwy1pQxUYgGVj+l5AJQhDNxJOOK2CyB
5LaxFLrja4CQfE3D+LQ7wQor2ll4lfESR2CDpurlI6RiO9eeOzqeSc/I42v5jcbl
AoM8JvM1DHRQP/Kt2HgPveD1s3Srhdgly69m5bvEdN13F/Xof15pn8uuLHRzVOms
Eyu2j00pxaSaNSdqZOw0WcxrGSJJorQNcHy38i6ZzgZE1njOOa2acHCM/T5iEoQy
edFQ1NrVIDbVS8XZNGhJMWoZaVFf4sVC4XqBIxs48ckpO2S06NYHcOGiOyaPKrZ4
3DRsdCjGhHfHdmH6NQCmEVGWRWvITB0Huvom9BgERNqkJJ45fGEviUZ9lFN1tKRh
l1XZ8sul02zKBCgVB3rjnjF1LAtfXogxBC5PkDGrPWHW0nBb500Mv2BomVh60Oqu
rSnnO2n7yFiLsLq1rvCGrtwMbRbVYArgHsDbhqPZWhOlRO7ofjPc0aKUj4OMc7k/
mPn13iwpfGXUiJIqukxmhE/Q2/GXoIDF3q8pklnEqV4jh+vXYIh8bLBhvcOoLD2q
sPyhrTzIev+nmOVeSFcFXsEVTWTbhQix9vTXqn2NlZPzzlT/IPgB7IeWWF326C+m
zUuUmPELIe+xTI6EUNxVzfpk9puPvcEsUN+CvfV9kccl6+aRFbxPqLt5J/NwMQxT
Vnbc0lGr6CLZEjpD3bWGHfZp84/KQjlwOZuIWCtNa8b9IMLkTBiU6S8kGFiIVkuS
5kk8FP7dI/Q/GjwVdKUTCgQB2Exorgwit879tXFe6tMpssdOmJoG/p9e+Ns8GwRt
qOF/fOCRAu92C6/EZJSyRDT+HACQtcEcd5x/CyIPz8BiGyBChE7mG4JtfGxhh05I
iBTFeVlMTLxoiHIWZLn77tAQgA6JvGwehl4Bm5t6Clh2BKaePbrkobw+rfPXMjRQ
RS3PZXKz5Z557Mk5EFp2dPHoDYikR16ikQyGf0a3s+iZMrHkzK47LLgFb6e3rizV
o/VSeIMMh9l5LssuIPjABq8aYhBbQk8jVWEAmutrMOKe9umWDedIUbewVpjBPbUs
v06W7TkHdMMWDtDmDeSABSpLq/DnO6a68KhY39yRjXCCzDW4w9FEcerFZtguYCwB
DlEZAIyU2+CdA1Kiyb8BvfD4C3bCN/ri1ceJ4vQcU5eTzsFv+uAYR5ot4I77EkcI
QHk4UBrUpBVKnP5UWhKo1RWOUpyfT3jTrXs3f8MRCJJqlrZ38CgwAzAgVrGjQ7Ru
cKTuDl+0KNT6CZOOgMcPk+rY5wJAxCxa5DtgikWpLZP0x59o5fSPWS7UelZNXMSy
1+ytuXiGNNTGioQQEGqJhMCcDpTBCDc/wcKYujz/eOlhL6ghMrfaAfbvCV3mO9vG
MNlw2Ey+zubUw+QP7/Bs5sEUPT3fxoKeCMlf87E4GX2upJt35qT8CsmFA1QhNzNr
3P0DwUrhJI91/Da5cT+V8FKA6x8mChUEY9Jlk+BpjqDhXv8UhnMIiDpq6l/Sqk8D
XskawfezQH3w3zZnEXUfT9WHbA3mdGyVhdAI6/hFVF/VnQevR8wNwsenDpxRThow
im9HKQiJTknz6CedN9tAc6SSo16j17lUuTX8DbvGHkGy0FV3rBNoPzSA6RMPdzK9
fpNJI59Nj4vq1HT/0viZ21XHtWtYIsA/BXWkSfqUQCnM8D+CdNSlt0x3ma/zJ3xp
W3KWfjW7HwYAjYkNn/NWrMHcSXiDOhhhtKsYqoiLaDXlDa1mLqBgajEdGUXIIWSl
9e711fURTyXFLbjDmCYC7qj8XRsj134j94hV3cpsl0OQ3B8hVkijEjjO1fL9P5dh
T8cgZziRCusi0X03Sv3Tq6fSCP22+V1YyHcAwKkO87txpPuDPZbkg1tlWbQSUBQf
JjPhc0NYrZ8DVpZWStRtekghiWNZWhYcu8c4CBF5NxBU5ELC254p41ortDVgdrwp
pHV0iBInmYUVvrx+VvJfPyRjkhoUNy6MYdh+Xqx/ei2VqR9b/D/s+eeWqNtgHQgR
ZIg0qKStqq4yqcsRILmL4x+yESxgstVOqhYjWkVyEc/pz5ZEkgBv0bLayAJiMmr2
mPRRDuFuWRO00QbK8INnF2uFtY6gHv9tYyJb2luNArPGGwJ2ssy+0cE8c9EDJbK0
13GO67vgxvnJRNNqac6a014buHe8dftu65wJI8i2u3TiZVmkOf/3SXhReNz7QrtH
tDv3G8r+HtlSw5mrWuBnkuOdr6SitaYM9ZYsZdGjCOrtVu6dtKZlsioMPO/n2PJ4
uqiPYiJ72A/cARizm5moilwlxuLpv/VkMONK0/IOh9UXSsBHUldWtskutEms+8MH
sWbFIHEJPNBy4wWN4n4YP/XZCv+58qAFZ46X+RISN92UK4SJsq6eh7hKMbApA5XL
01Mea7bJlxz83w623002cDdjCzaQ2iyBAXXEhYfPDQrecKiVWQozOMgsoLVDtAxn
b5/t/u2Ff1xSLzqiCs81P7Hur+cCTM1g1uHUa0yHjFKlVUAbrKzxAlPeJ46iSz8H
muLtCfSwz1zV0XMyLaV7CBpphpZ0VSJ0ZIo7TpTEuPGE2TzKX5tPYZg4kdmKw4xU
3J+a0i859YtAuuwym8R/ahzoqrr24QzThZV4R3r8qXkvjCFau6K4nkaW8vcrm4UC
jShdirQaLf8ezyureCJ3kVHU0JPJCYojStwhfa9MYeXL8ZzJxCfJtCMnit5dcoO5
3xcVy3fabE9QK7EbKRkSeX+cx9xHXbzOav2w738+nmDlacpE3VrUzS+iBYaK1jNZ
Sann2EywJd6o90HnqMhq0W5MhFYwyMJXzdnLI1fP1s1Y/5OsjyZ74XmRpL/Wpaid
+S9ecR8R+UnCU9KqC0BeplQ4/DvnccAmA0kTQb7qrTAkxFANdA3c2HDTKUKeGAvp
m2brXne38yKh/GbWK3R+twQg1J9GZOlKMrcBkjFZNjRzHhscP+8gU5wciImUV1w9
OCHDOvQTRSgzdgKSreqZeomhHbM2BxWdwGV7AGtna5SDMA2gwz0qMjE5a9RTKrkj
FimhbT39epwfcVhuC004Sf0YUM+636cH0flGsxn3U3DN09ZmlgGawoMLSGi1lkD3
ubtUIqjOfP+PFhCGzuAmlpAKlrCIa1Y+dTPz8u3072kJQf21p+zycJ4wbt+zykVf
W2T0mI1Kppszd5xEEIIZf/fTqnLbYZ3L3UOsrWWH9YB0h4AaGrbYYodttEJMdXMm
9kZos8ghKpabXMLWEfKMf9liB5DjCWrKCa303K0D17j9EeU18n2bx8d14vcmH8tl
X6F3NQT2sNRBxkNlLBHtafKwTSUnWHQHjGwe+JE1FCGWqIcUDje+FG0RqlHzT3zg
QSf/sWNRK/b1wY4GNLGG6+3RKgyThYYBF1yAWlgFVPZ0GW7G6f0no3ukRS0ba4zS
wgrUWsCutLJqotUXglIwNqVtd0hS5yVb5MRzjqn0g4ahVA9clFO/xo9ztDAek7cw
R1PvkHOFZp92BITbB+sE7WW2MsTQ+mbbQyY0s1JFXQkYjiljZ/5BtQisJ/UVCHzh
RWNesIUlh9PgdQToJltYZa3RmKVzX0ioO5Qo2pxy0bp8Q9y6wrPd4dG0YDyb4I8z
/dooMRqdbpJs7s8GM4pYeUHLuu6IoZltUiRM5F02+PuvQIjhx3MP5fzphRrbw/NJ
bgZ0toerNR0aYSYqig767MQBQU+sW1V4rdR8UkhVReNtU6LpvzS65weLdJl7d7ad
lqaeCYJ4F1PmkRJmJRI+XdlbV96ZPOvW7XqH6bPzrhZt6t//SaRCfQkCTa/mkSR3
CneRLS8IslaGi8PumUA4zxWN9wbUL1Pj/ZOZGPJg/XQOaglfF40DHr0ij5fWvWji
cUkioEs/+VJBntqlwWmy147xeLqr7mPqoPi3XxC/un5n+h8ghRWMXmIx7GmQ5U17
dWSo5JIHhXDU0js9ffSWD/Fr82iYWKfFgxjm4o43nHfiPmJt3E5OZc0sz+ikvoUJ
WX2dEGuCQGbeBlItopqh0RLTsNIp+TwW6qtOB5YlRFzeAuQLtsFcLy2FlzX23NDU
V3zpxNjbS47azm26ZXiZO4MS/fcsrAzVrI/dErfkpxFU6LYJ13wiyuMUYLFJKVn9
dHbtRAS1LffeOJm2PmO1PAsCix70RRwMXHL2Ojo1/PTmGZQgS725VpxuHYsKvIfh
TPzfpEi5hlzuZcHy6JyxBWxCWeEpd3e3PfxTixrpj+Cae8kOq8k4pxH3mVOEUHlu
6cBLbJ8epaowq18X2C1cf2WY6vuU4LxPI7gajlmBNsS6enFjAtnye0zL7K++6k+q
qQoG1sH4J0LDLD2VMBlRb0n1rhw3ycfWI2qPOl7+rkh2t7FAEOwNxPFE8JLt/m3f
yuieXI5n0q8wzXnTYQHAKjoG+M3RZJWQwcjHPWU/wqXnTTsdESOSdnFtDYfu8xLX
YkGjSO4UVtoziKIc6FL/G2RXTUX88ccBzqSEmmogRSlZMYUrE1bIGd4aEy2Qrkjz
o/J9CDtkMKfyfXiF5l05jhM+OM4H0Fb1RNlGixpR5jtrtwOfUs/S8IQ99ztb6bAZ
38TYCpK9gOhCD0X2XIR0hz8dGspYbxEzfEC2CWvyP7cfl16q4rEF765+pwJ/2ZVx
fFy6ZhMwf/0NTgpitmOzdePzwuc6JBuNT+UhTNC08Eu76ejpnRUNuPVYyzUSSsUQ
1Lq1h7GPfsTODSKswOWzn0lv2b5pjxYVrFT1vjm0pX51yywN+QOXOVkh4/CCkYWA
m7nDHMUi77UaMiUXrA2oFwwKy4DVML+B/2EYmTWZPkkXOA04eVYc5FECOK/4O2HM
XEumjd7qYEc9tcftK6bgAcy0iOWV5FWO/esVLwCBCX1p3TqVDInb5PR7yN8HK43d
6YegMszP8fOf3BVSGhkTAuVPLD27FzEFHJVLc935RzU3DzNeEyrO1VsZ7agWmJml
rx1MTD36+3hFPtRRWRZ6T4s+AwOVp0ml4N3rAXKt7Ew7vU/CWNrXqgQRgFhPG2lv
mfoOZfo/EbtEWKfEj1uT8yCT7Z+wdXDK3RBMgfFM2DPY4SHNVMYfCYREBoJChVio
BRrHUVWcO2vIa5VlEbZdfcmLXxVqgN9ofMDVZSpHC33KdxcvPS8LRSc4LcUfr1Ce
UHjXd9zrc0H7JgEG9FEbupPbyXDt4pbNUt7K1/xE7RGoQhUWt3s2QDRTp//erSDF
+A2EFrV3zH/3RNc/kBRKmR4H5culzmUZe77n5GI0mz/anqBR5/RtbR1GNOV4y7Oq
8BKfGVaeNS+BtvKM7ZQ1mnqMmcCLUMsa6KpUqMoyuvpbLL7Jn9mKjruLa7az8Y9f
3hPEsM4zB0BJ8sod4gc7uQldYEtP1zfONdjdrFf8LGmTdM5imTOtjdPQGP8gXkDm
oVzAhrdlRmw1haNXHfWSrRAPgp1LK44uH0KO7TI0M97zfynPf8CBkq9mX3Z1Rx7e
ooX7VxwbuDBQpZhL6FSouuJMW1urVl5iMD4//um/zs3jCkwjeFZT0lpTwoq9XFug
s+1qy/A2V3+pIvuD7x4V/88rm5OGQMuDhBkEBPOwSXs3xD4/ppzSt61N4anlnsJg
O2LbslDE5+GYfdaS5C1ICtJ0NmPZMGKu22vZG9OjIMI95G5aXwZGEGuaTbvMFcIH
buRmdb6fwjFdJrPUyupJpMaioazHHIHr3hrrZ5MdacDCve/pRVyQkKndAWJdPGLO
aXwSs9yThXDExTvM+m0Xz27y+a/5Z8q6ZXm2mWzqK7hHL+1Wt4/Y6++sh+FO+yi7
kdueZb4ymsmggNhRrG1cZzXVFvbChtt59+M0qs4vagolZ1yDP8CDVN9WCZU6Ve63
Nu/rDOwBwkhQQNbIg0GfGxHbBoaFmSzr1HGCzGCeaelkOuMgKiTMAXJbL0z6tuY3
BSEmDJ+tlfJCnOVjzhZfiubUtBoX2QR5iwKw9UB+EzhSB0ZJgAV+rvKGUx5CNNQ6
QlGTi4Di2LYP+TRx16vCxxU2XcW9i1+55hZSyfBLL3/VThiYKUclAtphLRGTiWLZ
5SsZcWB+WDGlW0cc36T1fvJfmeK+AWT0oUQ8a44v4D0AktF5Pe6HgoR047e5iKc5
liYqRt3DN/JUkwnpBMT++Jx2APpGSmxv3i6N4dV6Ku5hl/rkJPCfaLKiuoKXyj/y
66R0TXewSGCkXREx1FnF+xS7reUyMG89aqN6Oq82UA3BvER8ZJThSZs78koXoYeb
B6SyPde5i1zvtRgNaOApYPOiOiD+5wQeAGeTFv7R5JJMlxvFxI/vzwCvoM48eZuz
6d7O4iGqGkkY9YDuLjgIBe7GnbVmtgY1B9LV+fHlQLUCRfDmf/bQKB6R8ljgLR5L
bobGUtb3ohJAIE1uOEA1CPDb7GJcnXKkuwyU8t4M1rVRI7Yb9MwZGezBpFcG/PRv
z/bYsWhSelt8O0yRi2VOLt1dLycQ3xC5bJ1Rbv1DHF8PmVs+Q6TSPA9fJLhk2QSw
PQ5usRqW2AFalO8VGkpPltimyS3TFdnS8jOLbQeJgZI0V+CWN+EXazQJfv6V+R5L
RVl0Tv9OqRVx1y6rpKk8JXuuaAZ6lPdsUqWtDgHHhvfhhd54ksr/ZrNY830BgeIx
334F4rhtY2sbawSxtBwMkBO6GRDtFfBPWPfJ3kY3JJUMJ18Y/4AqkptLaONzB6ii
6oqZepfeGZ5CaAyFU2DVnBH9n9E44IYByzWvp27Uq//Ru8YVOtI+w2O0DT58/8Im
V6mB1+/LL0AgLK11A4EQVxsEfumcjGja8soAQdPdKBhCeht9g2mj3g8vlHzDGmUB
YOPZURoawtaS+axQTc8p8yeF53TS0jIrq+6Dq6JUmuBolQqlncdtAj9m14zn7C/o
+SzkgjE9LzQCI+64EaHaITTHnnucxcQEN1GiLe+82YYOYAJN/kObMMHD/A8wSzF+
EQAu85YWheuu6sgfYJSXW1c72txai9bCX8jbeyuo/wpQ0mXmQwfAQc7o3U4GhrQF
chs5WWYROg16Fo7jPemCihhDn5M0iBSOWJOiTp+Acwo54WanGLEKn1kdsKHtsr+F
lAcLzoOayDQ4zuSlsCYjV+nFlsEbGVCCUF63tImg3r0mFjT/sqTy0/yW4whSxdwW
JvqFAbyhW0z7xcvCGk3867xOeVjHKElcwxWjgoPOfymWQw7Fd9QqMD+yDvH7gzsP
SPeBFmDAGpr23FJG+Ae3OH2ERT3elpRQn8kW/k80HX/zIZUUINe+rq5/HOUnk9QR
y4E0YdWfSWvNGrP6mt2J97F7wrW0U678TTSQYdJEbMhBn3J6CO9YN0rv/+Y2dTMy
4at7Sv8gtTJGYdzRTFUSZ9OrIiUec4Q8h0erWeCR/nAFYmvfDVwP/L4WTdrv3uYE
+V+FC5BmIUXHooEvXkukzG7+KHxXB7HGgkDwDTsDGS8zzRX2prYINAFDIe1hS5+k
bbe1O6k/St/0Pw2Y3Pm7+199Y/O3mTWrdc+bad5l4FIcE3HXTNapSl/ZI+FD8/vy
tRv7PJ6WITMeSoETN9Vggqf0Nlq+JyNQ6MPXybjLboh/6K/L61bZaRNk2lJCj7CO
i150fcVYjIMg5QL2ZrCv6Jre9pmgFNFhGUF9Hdsrck9cP6u0kkKV5OgC5ft32efv
lbM3afFYx3JWcmLJw3RsrtiCM8xxVbsLPB307PAT1JnEQC8yOu2nIJlt+IRKZuRy
376C2fOefglZGvrFO7ry3wGcp+3KQv8vXR8/zJVKS6Eb4WvBhb6gG34N9gyneWjx
e5Tw3KzLklxi8VrRyiyO12YbjwMMT0c7zomGmwvWjbZUMaimt5tY33K9mnaqRtXq
5njDDxmd3Ib4ZW0yUAz94KFHjsqO69nhYc55U6uJUnQH+dh2g2BcpSKdSRpWZT8T
M6IBrGh/LoOkH1B5VoZskqsi3hZIN4sLeUlCHPW3irBIvqcUlwFmK4Li/Vt7h/wv
Pbe2GSuD+loMGDCCGIBw2FDnOeniinKxGZJT3gYIuGaLmMe258ima2jnEaVxxEg6
0WkKdfoCJUq4fJ9VAZU+q+jnWp+oHNQTphpF3B7acuko6YCIl0NBlGHNE6YTSi6j
vVBt9iGFbuGInVdl5iNQ/reOPCWFBTqIVNrCniz1Oiua3d+tBm0hUMp/U5jmhrNn
p+/ttxfbsJtjvkaSg7fvq8TG32gPmpAs2uJ+2ZCvzkh47Sa2IgZCp62rxxNzkzkD
yh9fQgF97WpShqPCAHBIB4j750IAOu2IfWci78n6QJ1hHZB+Fy5pyi7zcdcuDnM8
OTcnI3Ijg8E+C5Mx/YKAichSmFF44i5B0YiW2+I+53J4kXq3BBEuSKRPzip+BORc
CwMUxsfpXHFleBtIIJRG3GIBXEwFsFGRvo/SfUlesfn9kLIWnTg13Dj97oSzUPXg
1L5QG+rYpF10KZ6YDG/jbfk/hBOdWX06or0Tkwpag5rYUldSiHsTgm5egH0438nn
n3YCVMPblOj8B+Sws5U9cH4EH3SxuNsP4U5F5OfAfGi8s5itHaBr91hzlgowlsel
e4iJndd0xdYKT7cJIrokv9RXMpQsz4NPpsnSk4gphH5qQCn0A8neuCcqjXHSBJ/F
KCMg/6vX9Rh032MDHIOa6L8rFDfSUkfsbV53zKFnnUlx7JtbQTYgN7FVy2YxqEPn
dyayW/OCfbQm6djKDNHE0qxe2k1tMa5PMsdSVZEjFbYIQDEsfm7dk+nDaUkVZmgq
DT1Y0ruEpLYejmRkoBSC8gd+qinOY22n8niCZ4s9HiBWYaYTewPbdYzSW3aidq3w
UxatadaDhz1+CD9HkTVdGAW5cZGf9snmDMsmax+qlqyO4xKVan5sRwRLpEr2V5Vx
4YnxyyROLBt9lN3/sbWAxwfU4NSUV2sDKNKjCmMhGwzIbMBbfstFn65SrjLBq3Du
Y6VJ7HReHDhohPua6gmUSdMEwebM/apjl2n1mmMI6NYw+UjD63jUxNLaxPvY6I74
HJ2q9VJmHE9ywr5h/HBBrb8YGLfMERPBZzvtfaip8I7uTclczBfnbp+YE5zZDa/K
jSdH3WCHtLu781sx834K3LEe3mLwCZxGSLqOoYboeHc/XEq8MU0VciTy18p9I+qa
efIJJzFKlzQAPPuUJQpQ1nb1MxLwfI2kxTNlvR1k+qz6uCxxcV4HnMTSkE6lpQ8P
DrR5cd4qZM+Jb94mBi2XRCBXEsztXM2y3ggKkjJX/cz8CY0RbPulNDJ9v/uLSU5q
IAt3gmUO3jgb/hxK7KQyWGPPA/re4zk3Ff4N7BhftLCzH1cw+lIQMeLKd3w4sSYt
U7lXxv+2YJex6tQ0YF9lAXUqGlAylLdk6ex+gSHy5Ips43Hh6+1emFm0PJV6kT7W
qJpi3aTDqu+qA2XfR5VjHYCcjq3hRkAQtPIS/zNJzVGjwwz0ZIZkO/IvzDHFoCUe
x6UXBi9fp32LEHj2PwgcCiBj0E4uUt6/ygB24ld+wRtnQs46Kqr2K0GufeV0eE2K
tesdMSV1ic5ADCbDfj/Qbl+7voQnHRVVSXJ9OhT9/gVKYNCJ40XZd3HcINsbkCD0
iY4TjJbnMcL4NxT2WHYAUvBQtBhWwQD84tK7mFqYMZsleoiUBnKvAMjdzmRYLAyA
ZeqdA35jNhL3fGLxn//9rND5CoAMWzTaGBs7Lc32jfKsI2JAupaErW/1VYZOSN2i
Y3+Y4fg7s3UMyYsu99VnzPSvle19NbhxbJFd0lrVKl5udF7nIIgBLoYDxIVqHaiD
9wMR1PYh06NINiEJ5POZ+EiQrfYdB9ygG91r6wO8NSw7lGxf2j9cx8VT2TLVUccq
VSkEwAA49O+Ww4W1T4xmD63+I95O7g0C+IbzQOo6ErRGscFM5mVNDFUPiKolRzWv
i8dzzDybyVEqdroe+gLRwSNsnoPoMSUpI5ivSkDH6Y0z8vq+67AcEPoQlf0eDXbf
KcmRwJZLfAQa6H71KIchGkvCRnhKg6pLz2VOFCgeAQuJbwBxNN6fOJzfcR41Dnr3
gFl90hs2y9jPVXUu59mG4hRUNLXKab/T1l2k3+DwI6gHE5oiSNEvF3kI4qGP+gzb
qkal/BrJ4AKT9EfXoJgpk38MhBkEQpWbslSqDYlXHO/zOYb0i3QTGcSRnPBUJIzi
LQG3yMveXUOjenI8j/ItM5IWPijj0EYqanOYmXObk+HyZ+rONAuZTEkAD1dYpPtj
RfHqnXDTnh6VpUu6B+w1Ujw0YIISHlLNRK4QMOCj7GlTEXC4aDOlYDFjUKMxnWrZ
Y9ov2RaJydBbtkCkJHAZK4CKKc/n73wXm3gEOsjzdtQLG307zOqlu1F/x2x9u9F0
7ZgGtIbb9YqyC+sLA1SUTF3PN95WAb/oBdoJjbMn9mJ6XPARCnEPp7HO99RsxH/A
J3O2/iUMd1ysaRyf0IMBlLfoevdAWr57gNnOcv4Ej3KICX/C4c9iIUJTWa+IAtdr
IHsVttrl611E/jP6MiZFtFXA9ftHxFo8rjIwEy2WY3jP1PDJADbfQQdL11o2SlyB
sbzEfom/hwDgqoAY4NflmbfFuV0g63WW53ITIPP2+QqD6Mrrl6UVKzaRhaYgWp5k
RvrTdAkth2bHz2ZcyX+w2fsDigiMhvUWf0H72CeUnZ+iRMqdLsKQsY4Zv+6vWU7u
yoX7G/FYK87WJf0nZlmbdMsJzb2wDC78ccVUQkXT91hGsONLZ8ckFkUraK/2qxwN
MCok2PZMjzhAZvworXvWXOHpa8+HtOIJxkMnFjeNJNGxu8M+dg9szwgemMFSIdXA
MgV0PTfXVSvpjL6K7JSMWuuEgtWVejgSCOJlVL2WtbAFSnxX0Ey5A/1nmNLZlVom
RS2Q6nofgdgh8yLBbRwhw1qOKoF8IIqyqUrqzUJSp5NYdpDz3kQW8bKbElwr9BbX
8Nwj18MPTc8gw8FPmwg6UPt0/oAKKCLMGlDLEiQDg8dViUbRtXgzjtwEkudgatNQ
UB40PDDNwzYmtPgYmMVHNCzMWywDxeFGRCL71zPqN+QZRf8qzI/4d9B45DE1ppRe
ELqMm09YQ1BqRVQCOIxFrdlY0Zidh+gKuUG8MbOFWxHJJIJx3r6GPJOBPCvWUMMY
FpQQwPrbbJZSCh2OHgdWQB4VzZVj5qkHdwGuqMtb38/PT1mmTmqS117JzFbXCZ/D
5/ZObzvbpTmbP0VbNpfHDD0R8SjFAwmP3xeMoSEYmDD/Sy8Xpn1LedRGe13VV7TL
6YY+suvwJAdVtjGrHIbP38anexQv1HcMf3Rf3SF+djPZuqjuYeTTR/WJ9hitC95+
JtmBixVS/X48cyKXFS4a0FLcWS8C5E23NRMBJlpB6eefaONGli4wOo6nw3LAgQFV
NgTvzdvklPGTzHlQpCOronzQPEPgqdDIPoZY1lhv7nx0MsAElZ21VEHtZRISUY8Q
CwQFaiVS88nmZTugBx41q6aq06N1ilqsMYIHgKHH18WCBTyPESpT0IsCjySfNOhk
ktzir6opXI2aF+7SKcUIlyuh16Za4Zw/KabNdtMvb31d7OlGzg88iZjXZBB05u6r
0C5if43tCgLcUiRxEbIkemWhfbms7T4jOpRCUdALQLfoYpxOnW2N7Z1G/T9+Gnd9
Yzuik1JZiA9QWq9RZHk70M0u24tvAKrXNcBYzIVkdELOatQLDxghdeEalsMRWNqT
jW96s6Wnv4fhUSuNvBCy1OVgbMtqsJiCNdyqxntlclx1p1mawcM1IwP0b62nO5pM
CNWV+Ezg9B6/QeNWrRtuE4vcFIQfeU2DfHLBuz4vfoDePGyfiAoxps5yhuwjwxo0
0WZdoSFQbxHyukxsuFt9QFVXfTmY+jwLTHXhaiYfs+B9IUC3ob4vLQRkBVqCqTRz
DrkzGfIDKDDcZcPYx+whqhn1LPElyBCUE5VTtHYJ222HF0h0axIuv6j6QRWqT5yk
OGa/Ks7kOY3LIXXMIzJ//jorrHzEiYjUncICwAc/YnBj8gAr7bhIkO5rDSj+niwX
//tSHg+sf996uBTFmp+p7iRCoF8skBk68uhZ4LeAAXCGeeW9VlMCGszFYQ9G4wd1
8CPz1i+9SqEzrb/hAyc9NgR2wwmIMJdrSsuzAJiK/F+yyp+jUZJjtQQnhHH+cKcA
KBUHIj8iSCQ+pMaUIogWn5tSNvuE3SU8a0IG8Jz+N8WFX8wDA7fcjXZZahLuxyVH
VuVJMnW9zt9TnyWtWAheJwLgGLliGRgQTVINq9xIYafc6T5YG2tD9xQEB0kG3J+7
8X8D35nMV2LIllhV4QSheT/lFQvlJEAAvla+y/eMitp0wEUeTYRXf0WanzyJ2zQ9
aAWNu8nXPeJTgx7p4IDTj4F6DowkKBqkr5OOssf2VmDLBJKf6GmgAu/4HujYVmIg
Q/E6JAP3WOxMRCxYlA6djEU1UHprNuYl4ukIdmhI91huSTsrok5S6cWoEFqoyUiK
OHO/tqLhW4EfoVrKxO3IWl9AhWJtWsikPOFU/H5RIhLh+WHzr3U7fSicJ2AgWaeR
VUZpFR6vD6LQAJN3xN8tbVBPhcG1glqIFkjta0ko7lkN1H2gsezPuI4/gINKBfG/
90STGh0QVU+b6o0nxzGiKVfG9W2houaVJ1P8YDdkRyFO2dP0S5UDZURAYvRrkE8C
2PwBCjnNYXRgRL99KLJ0H82j88pm0ckZRynXj04eO1VJtmnSvuSV5xa16BbTAMFf
+NF19JeoieteToY25AWeZEAq3W8bPV0CmRYqe9VMMNErRcJgf0JDipq54aWX4R4w
MVuItNNUAp0dId8s8i0UtKlEOARl2DD5+wder7grtO+ShlZ9s1FL02z1miCbozFF
u2OjjgbW1lze/l23tQAsO81ki/450dqf6mC1ZQ2P8H1JiS/CCpMGj6GwiV6BnBfJ
fBVNhxr6dDz2yEPbgIfCBkqF0Q+dFBbHKWWjkjrGU1vsGjd24yU7WCtu6CJs2LtR
U5Hv7e12Zo/xUZVIbi+dwFGkpbze866K8SswbKOu3EEvK4d+hJxk9rGwMItYtyR1
4N0SAdFGUrd8lJGWPhYREBVlbtcgaiYBPCokqo5iYzX4r+gWB5bqwA/MdFEXaHhg
tlD9KN4oic1g02m7Xj8MdukaecK+Lo9WZlz7JYyFMysiV6rLbeohvfolS9SPSAVE
QWJs5DDv+tvrmekUVm/4k/M9q/jsVrt9+H2wVPoJsl4LMIyi6KQM2p1PVlKhaxlA
V7tGLZZ4rrvv1fs+y2U05U9PrM7x0tCcz5hq1teFLvNVcpwk+kvuwNdLqkDScR6W
1kfe9tNLitVqwU4ddMujTgA/KjP0reugwiBq7dnXtWO2Nng4EC22z2L+o1cavWJV
EQj4nMSqoIYx8DKyU3FbLmWzZ/JRFZqNwNP6H1ZiVAIkV0/7M0akIYDHwqVoRQVA
RerztnLgKJpJvU3OeMEQfsZ8+pqjbZdIS0H6DkIcHoFjk/Ij149GTzUGPf82g53F
fsqJZwSfkb+QcSeHCA+Hy6BJsxfBGwx7gD9HrNzUo82SKb+vhqZUM85i9YG0//gS
4q3KKm+vEcwEg0Ik6m8Jd3dIU0pgAWzMFVVg4V8/5C5Dnlj0jhcED/dehZjpW01i
PIJm1G9fEEhXe1lZq9yGtGsBHpvLI9BVKqthvwQsqaddE4y3lLO6pNESBzUj/d+e
CEGFhzlfeBWX7l5K2PE0JE3m/iH53NCQQ4z8ByBM7PokDHe4VXRlh45ZmGAjMACi
XqRVCiJvNGY8OqCnfvwlqpB6F+SRwjHQSBWEPdB/iwo1mMHMYYVv8BwcNPXutt2w
opemiHwmWYBHNCnFHeNP3DrlDJ5yKQLv1+gkWpG4WDpdF+iWEjnMSSTqG76YnuYN
9YaYWwbwCCiO89wE1rHwnk2gNfU5Te7XcMFN8FyV6TtZr+y06g3IQhrk4DxR4kzi
Rr0x/nn+Nn3yKh+kq7a+PaCvPV0ZhVaSUvn8Byhqe5OJ4WJuEIbjkayr00bBwxus
1BlzC2w8V7HGR27NVRlhV8ih9hzA8EvlZdKl+xn5Vr5jM0xR9XSYI0QKvEGdLNVY
lvg6TyLpqUOEyQeJUWNcXqTHtirfka/zVKwmkh09eFF/IKR+CKX5iazQWeH5FjcX
uJ/o7VUPe4P8MuNFuKSziJkANlAYpADk4nSNFA7farLhat3UBrkki7aeUeKDNyA+
WpHvLku4Yr2P5PM465w8WnSij738K+LN40oNwoPGdbU93NqGouiWY/xDkwz0uKLw
SLDD+5U48zO32NuZWiKQENcZeXgNBMOOUIVDLCmP4YeMJxw9Qebg67nSnHhUtt+U
b/vcQNOU6ZAjT2uuz6DUoZ4gB/3LgDYknhGnnvuUnDRmBMYIHx3lwPhJ34470+HL
vwj2E420emjcCqqzwxKXIzvKtYPpYyKvr2FtHOjjzs86ih0UxAb0skWQ/RRayB8O
hH1hzbTxR3g7JTCxCQcVbQ+2C3jPP75v3CKuFtETYA0daUdpGRubkLj0oASTazRw
Ypk5z8MTDjmKDA3kJe2wumtQ1ChZ/LniVtoRuitG5XrcpeBT9QnJJKCOaSVzINbg
Gn6UcfyibIusupI1UHQkVVuSU5qLdR1li9w2mBI+2r/dG4aIK/g3lCgdW7DsOE9k
EozkkYIJapFO9Z+OzqGYQ3g2nkiKv3BHp8YMK3ebhk7mfSr/fasNd/SOFuG+LLtV
MsRGlcmJ/xuj0A8vzK5zuD01scmkZf6PY5IWdHGosIUHmVPlLC/BoU1GM4DjisZ6
y7d+f81GbY0WNJ8dnY+LOUi2qcmxN1OW1wcGN7K5RcvHPrJSjm19PWE4oEKuGKDm
YAlER/mlOXMVZ13chkYqaRGs2XtroQrXgZFx8fnAl54ghlx9nTak8HppNzJ/DMCk
a0W1aE47JPYTUPlw5Jmywx5xdL1Jfzwc5269yl8jcVukLwvRCTvDN1IqAQ3+gvva
ASVfRbhCnpq5oYwvtEMQgGCuOjaZzqCpFluOAsMxnGzwxQue+n3sUBQTYp9GeOrJ
dAJhrbB62zmayn/7yuUpCOprssHd13uvMuywT5Ok5urfV4cSnHiCubQJfkznLn8t
E7rP90YH8rurhCNncETLHHDVMxs2IeGbjRN7Mg+rAOPg3Sc2X14a4LGzF3mUta0N
hPDCZgcyOW87FLLICclD+BA8OUE9jIGY9jJ9QHjQ5X+NCgsdmzpylj4l2nbGn6jW
XefXMbCPNZlB0BsQWBFyUdpWA0nyHc/dP8IGhj8ZWDBmnk27i2Tz95aHgxfzxDCo
uBW2x36oAHdwHGwltbPQVXgXQHEvqfCUAkrDWj/twUtxfXUP4AbjZWD+IIjtxm5n
g+9DJIVVEgBP52zXC7YIZ0WkbqIHhtfCpJo5eoFrvrAYF8ycc42FsCwyBflh8h1F
TnlCfOp8qpA/Qhjck3ijLf4oa5JQDxU2H8n8oyB8Azw1gNbMA3A2A5qsSvsLHr8F
A5h4Nd+32h6OKM6VtoaCqjfwHKQlFRC36QWZF0Iz85aC0SSAJ7nGQ0d7aFJ4tfMt
LwewHKgrR2OYLIhcbfp7XBp1s6amd/PK7H2c5sOoig2DpcjsMP90o7i6NLGZZcWY
kCs1CbCAHg/5isrPfIyMOmRNB0RgPtvacLt41JVm6v99nsEBg2e3K2Qjs7onv9cV
cTucokRDeoWHTKCTPoO+fcf6mzeKLxyttXi9XI1siIPircKlTu3frJrUu15zedob
6tSj9y66phe/7z/ckKcXCROOLOHJ0tYiFdCPDgU7adMIFtzXbpjbXfisWz7btZLU
XG/CuKuD/GLxjrz9PhHv3wmkKo8ooIrEQyFHy0zN/HotnTbn24J1yYUsH24RW6/k
euiMg3dJb8aKF47qP5SPtBny0EuAKTRzaJ3kQ3VftEkWba7IDMsyxcbeoBSvTVnv
23FdichmilIza7pIwwYasVkL7i+Vw5fIiIxYnNGO0Ss73mL6SxaRFlLipA2gj99i
IYGt+SU7uOuNGjRWsDJg2jYUOmb72YgiLa9QJ+ovX8eDmCXzbjYFSl5Uo02e5mzi
5QVCou6Kv7xgdMy9XQk+K8K0B28GnIk2Lni+jUWJOb2S2OSydkFiGSBlr0JWuZlz
03rNQv8TXlCjvU/lmvryZRh9tGuAsoZBtFDXrzpJlmzq3KbpPpJVHgOx0excqBpN
rQqd9JZyr2rXOwBkx9fxx9ciewxvIQNH3U3fKGp4oPF6TUuQ1FPZcUO/+nkL7OW7
PRTViogBbp3yLpTcw+t/3MDMfWVxj3j2vb2ZlZITLS84CiidUcvWLsrM6lMvkr7l
D7xpjldtNrGiwYTG5gqiwghGwnkJ+5RwxHoNq6FNUPDCd7f4DjGlXneewhSRuwTA
OOHRPHMGxSIkm39Pab5cgTwy5OwwYBMrUGanyk2dpFZrRQvrVt0Lw6WvBosZE1M7
/2tLOv/TDiDMnIUNKOhMYRz4Dj3DmMmmyi/m7ruSeXykTA/lXk7IzDUxiYZSj9za
y6+iZpBOCKTcqGqBzySf7CzmNqrk55OvDOC5be79DGzbXHxmvkO2FtfjBi54+kee
w5McaEpC0tznMuPs9YmKqlQ/rE9SRwpiUKmMIFPOFFlNPStOZaR+6JaTZgmID0u3
6GRao1IrIYD6iz1QIA4QCki3a67btNCa1I6gcp5yCm2A8GGaTl2ZLtpS1+WQIpYe
ZF7y4c2BWMfCLjlBvixUDxZEGop+XnrvETV6wJMk7Zv/vbtTXd1oAGIlPHLwhRI0
lC1xhjBRwakJhKYT3oZ7o1T2n8FVVf3GRXPyGGhOiona3ghmCvJyR0EWROGnvQeW
saNFyX3+Nd5Iy7FAS532/9fyb6X10pDiLOxkW3z6NP5tru7pEYb3u8oQHsN8+tII
xxHWj7eKx5PLzd41xSk9VgDDRHQs0GWGISpDEatKUjiBrQ7qVZSfl7CTnvkh6dLd
e88VQ+HTtTGh4fzIC0/D4B9E2onAQ+jI0nTOJ4+4R5i2XS527KD5Y/bsGpT+H1p8
WJIL/ED+WKB45C3hpTFUZbmZ/pArS4DczO1lslK2cKBv4TSjQanp4l56d0cno+/H
RR/N2MSyTtpKchZWBu/UJcQSznAIv6cOxNNfnzCbsOJ79OtD9jIns9Iht8ysMmT6
uPVpYpdXP3B3vEiU7aUiq5vakMAh/sej5RqoukQd/kSRUVPMhglYX8gHGiZqncNi
Al+RR5lxDlb664jQMBJ9zy/aQW9/iOV2OrBKA/L6h5t5VCd6JJp+EpuWtCn7uffQ
907f8VHMrpR3HEjUZo/O5K62+1ETirNGEw5yX1wjW8yi/ie9l70hIyySJkOUTiMs
tDPX2ms/zybhUosMmEWOGH7ijEHH/lsZBZouu9vlE94rbyVD9WJ5tuJsRP1UC0jZ
88lVZ5SUZhEgcafxnINSu3e/55cT/PdY+KmXJzzMJ5Ij/aBnuTe1sqAk8SMeYWuH
t4psyiwwm9+BRZfFTBCRcjA9KjK3Wq5Z1f28524l8Mu5eOIQeS7nN4vRFmIuTzR5
d08hgOzxqZGQou8ZP4maY55XzcnoeGaPH+vzBb+pqU/giNJsJJD42tuLFMAhSqzM
SMn9IhgYMwrziUx1svzeCa+wBftbUuTVdPiPuI4IhLSks2EYUDs0gwlcyX9Aft0x
mbkT5y1OQtXp5l6M5jpfqXDQENp+CYaAG0DSzyNN56AfLTbqVpR4bIk/E/2Cl64r
mH0AmVnoVokQ3F2wHQlgT4QGPCiWcsQz4pvUH/Q/cyNLGOjR5I9jruIfbEEpfzgV
aVJJv/vBNCPoj11hwEmFhsEfZz+WVUZopG5Pbve3+Be7Ke5/AiMC5lKnYGIX+i4D
g2pqQa6W0xNBI8bZzB+jwarkx5o3L5qj0jFWOFv6zPYEf9EsQgfQuhfUcAFo2oka
RAElKqQq98/dyiFu7s16zSSXQkPds/iEWH77QBR8csyNv+Q9BUnCQ+VrQFjsqI5+
h9AeGC/vuW3b25koavymbTVe/kaPSJqD19TLrGRz/1n4MNtZScx+Gw/9nAjZqsNE
3pxtP+tUFpsVzlYdKDkmhdX0KCA9S5tE9JzcQphdKibJ/QXh5zxBpqGrC4vR/Vt7
0KDlBmjTEXcwwBx3ecWp1P9FuJivGSMvSb06z0/qofyscrUA8aPI8hIWM9lJ9k5q
ZT3Nh4KdHTr/kEeWjkIL8CViCDYWRZqhEu6Xv5+G44Pui3zTXudGrrReSAF3yo1s
7LuwThcXVWNkIiP7WPGxMAWi2TmcIm1zZ4I10syu7RkAQeSodnIuuoL5LwGzDsQ3
qbQ2/om8CRbTXpgl/BWt2QQnTXIAaX0X9mhaPvjxozpBi/2vqkXsEPviTXqaQ7q9
fRJwyxkyGirv383ubgP6LxfsV+vWYhS5d0ogQcbe7U6bsbcOH0w0p/1YcGF13bJd
m9of5Riz3TPr/8oNdY2WZgNLVaL3gac8NN5QUdUUQdlF4rIFo4D0numF2WnRMbIe
So4QuSzZhK/lBPtF6jhpq07ASAvsAmJhh5tkyBRQmV+VmLkVjwJKEXzXoJ40G9be
6SXV8qFsBLp4tLONGEh9pHOn3tMBkwOZVu7/KQ56T/MWT8gndZn6/DxgPOPOEzBa
U4MJYxLtf20ndlidqkVCx7of+GKpPz3vMWTNsXCJ07+nmGf3x0OZBveNMEHNQUwA
3Yz+SzwF60//MMZYitJ8Hw2D2mUo28orhxYoQhcb7PwLXDAb6uEJXntxYBAhWj0i
avLw7arqF2k2lXwzhFUppWYGF20PE5k2+EECeWGlTHWpAVZlJ9u9w8/1f3AmdbYi
ju/3I5fmwCrYqPS2XNtq0NV0JzgJ8RUXY0ibyvAVpfvA1DgtuhqyYZxmZvI0kKRC
PO/9AqK+TgnwBTS+cNssOaxAdfh6Z1PqQL41o2wREJLC5/9NuA5UppQlTNOybLWj
79WmwDd931fo6arUhJzV3lRjwCDc4e3gi6rGkiytO3sEXPg/libjzY7YMp9RIAYF
dxbjo0EC0BvuJjtFXENyBlOPfUJlutAdWKdmUvncI0oD36t83+eHe8LOcmzTHNKW
D1rNcEujqDElwP6T6oEsTS1ByLQyiWKmAjj2I7R5HyYv1V4gPEujBdrCRitxsxRx
fQDy8IrIrMpAaQQ4F9oCGsh23xg1Dd4MekFRZqHAxS6H07PE/a218Ukl75LA1xqR
+wlxtG3AwC769Ul9Ji05h+fQZKyKlbwNWaNRzGG7GtKfm6k1ylFNGtb9rApyAc0p
j2SdAJ+IKuWbmvyVkCyhnhGBlzk46nsf8i1DwJVT61cXEKsgBMP6qWBT29gIRKPx
1+MPCSXv+W9Ishfz/ZCFOVPCZskjYcgm70r2nX9BA8AukSiTIyjFgmTel6tlfQP1
sX7RsBwD8fUOilwO+1izMXNwjPs64WualojcRuzTBRQyoqbIDqqXD80e1skStwIH
QO2wfHIFEPy2C4EKy+1yz9AzJ8+xGshY5V48+PlQ03eiCjNruGItts1B2uX5Qi45
GSav4EP1k+yrt9kQNLRlQIT+W8lSeh36kDxnZN+lz1Tk+KmNVNlZsxZsOAI8pl4M
Dd67iduyvhrbJbr8rHHdNLYtgBfTjpSF54o5rtdrgJUyqp2JU9Yrb6lJJ2v5PoUe
YbrrkwUoj2DrT+CCoaMMPjhhfZCv8YbD9Qu6/J36okxp9bxkrvFuanF4KuxfF7oH
/1hIW6GgVtEMM2eQcIhljLDdOoLgn3Y0Oj9ETVqYeZqnojpU6AIAxt23S22twNVf
ZutU5Y/sBmBQlSy2Ufz9ShxFA5lH5SMZ6C3uk/GfsaZLCkK0lb14UsSQYoGq31Yi
Tjbxj+UMCIpyQJmbjYis30nmxqKLOC4S7heU/uxYLqLVmV8XBmqhrER0dLa4WFuP
X0LEScJDbDcljzxe7qSrVg4yhcnGj09J3Rnw3Uh4JZ7HEDQ3aafl19y2OSNGJGvj
xtMJBuq5DD8GHZ72Ufj3ue+LChAeJcLg+qSe34MgNYR7awvO4L0dheHmCMjkMu5i
eMaW1i/a7LSny3PlL5YoY89VXRyaRkVVNITUlhdRmd3/QdFzlvIta83hoMFjg8O3
u9EgxbOSfI1SbrRP+MaSpVXTDdy3jqvmBGs7ALbXXsJHCPBwHTUuy6jKC0LHKRgw
82QvtnK/0jsFd0L6qlDd/bjVf6qwmDm3aSTbAnvs7xkPOivEO4SQdk7W0ZETFOUL
HhUlryJVrPf9r1iefihk7N3ExDg9YJA5b1QsDkDgZHUd+j3hjme8SS+0IxBbn3I6
7nqg7wqj9Ih5qig15VeNRxRy9Nc0J9kv+cEh3iVxaV8MVLOCtNtXgDFfL9lvSJMX
P5hOXZSKGUxAsPDHc5G/ZrA6qr0uSjE2CJi3hOMTQ9/AE+LL4yNRD6iFDBDhizb0
U1DRH+Y3qrwkU1gjvrQY/2x9dsV8pysN2dQ3d48sEduMeBhyZO/UZCFeQi86EoLm
f8PqZKcH1zy14WPWAK+dVKjumn4j/jZj0mKLQ3R+k24LTgt3LMNou9KtOQRMmDFO
RyyJCxpYKwUt6QnM2oOxgx+HDTI+j1KTkyEZ6rdgyyMEuVM3UJ9CsuJQB9TnFxLG
GY4eQ0gfcNcALASITbT7tGBjXlZjODMqPHF193Fudp5HiO/LlV3oTE5VZWu8wfKU
C7taS5huew/q6k25IXsR/hRMlPIvXFibr6Bjr4Z5uE+P+Bw+6xZrG66VcZtnHakx
8A0f21zU37g3Yu5a4OCAGR9cYa4ZBWMa+Yj1RtM/8lfMu9TilvpWlfOjIBPUYm/P
2lTthA1rDVNRMeFP8bQ/7+/Vz0fsBwgUi9OnXyLtMVZQ/Na2HKZPLAzJaCkCI3yT
iJp2oBFYuAAaFnIfDnymz9VWWDwEuifeVsujBkRVZqw4RvFSTq/IDakXOaz5pmIe
pWfNeLZUz36lBlkwKmkD8Gb20ZmZcO5lUza+c3Et8Hu+pweXuTYhRwdhhCa+LidC
KyqRhjywekmM9da3A7SDR1z6tqywdhELkxJWMmU/INcIuXocthHul9fDKGz77P0d
ZsGX1iaCnTMLIYhEis9WaOgVgoy3QSG9kbjWJ7QZH6hb3V6M6CbRXHzwkb1IPSRD
ZtqsADYdTyX6k0xudWHLAg4G0tL7lk1tM4GJioZtJT/nui6DO8su371X1/obyYBg
vLe8LFrGbG9Wjn/8nKVqxLrnZFeoQRyJGjeD+GovkI5y66KyStfO5G10ShMXMtc6
jyRjXiaNaLQZEWszxaYvcc1sKbH/3sLGTvQATZ0Kxr3D0/BYGrOx6sNsQ7NWeBEz
FmmuQP2/hkzq8FCUp75xU8N69Nq6QZaxSbF+eftqaTPRau9saOSzyYAWS0Fqm1Pk
ETBuKCuKeKWIcpLgQZ1Sq6gXmEfUzItcThDh5iFnT8z25tARJRLY5tNkCjyzQLvS
1ZNzD5BACukteouALPuK08KwhVdN0vB4o5pSqCTRWR+759VAQEGfxC8EPDwOz6Oq
YY5yjAYhBwtOOcrRgh2lqcGArDOFoig/CjD6e5rwnYxSywS+U9GreJMEFQbNqAEP
ggdezOK1owh2T1+wfaAWBKgH7bCzyE2mBnuyul0aiPqk3RMBm47py36QMl5QZhtd
NrCJju1npx03vzb85OVGMg0m5T6FlCuYlC95rryC8NDFKa2vX2GQ6g9OvzOiTkNW
pGBrKFhMPookDdY5xRTEIkGQXGAwlVdRyir31oihIPDDIGf/WN9LjUwsBypUQI6X
yjRCw7vjBPBoRmKOzxY18BujV4QC5o/BRA4V9/vTUSb7mHYUYD+XXyV6pSkmgJB6
Mj5rLiaoTzPtrJRt+q+iT35g5z7Q1ixDjLnAmco4tRWV4qARZpvEbL8PoZoRDTCD
DJ4LSexsmqlsCAflCHDXq61aecHUV7MfI3JvQLfK+1V67AMcGD2UsxjswEWc6KLO
3saRVtw65Afb4S/UBUpneE/xm8Ro/8mZ7VrcpTi1OChGuXnl52S3nXLHOK/XU2vC
SseNJSxfzWCUAJ1Xq8TP4xaxIMog6eeWBif0qUURWGN7evNkSBidl0JmLoJYQ+G0
3f4N5EXyCdoTTQZF6yw3Fye9wSnT7QzVqSiq+r3lI9m3yqqWftkP3XeThmNQA4W9
N/Ikp9j+GQwxpDFkCgJ4y9f+Xx6eAnPDjDlDbMN4fO2Q8/yXUGffzIFGf2OQ6awN
1ZUNcaVWFNsuR/XavuL2Y6ZJTdc8GbjZYOE9QHEdZ8KOLKFqCKNqRKRGI1Fgl5r6
SzENcR6nGhPZ9DV0G+K975weS9Fvp2wM2XuH+96xec9rJVqHvLQd5ehtojNmV36O
Rf2nIbkT40opwGV58nUPM3HvcRhkpIMTuurO7ahYmvGRkYlcByoH6y1+Ffb6YbML
w3lw9LdEhk9aIE9QJpnjzUJ7KMjz3oenbkNSrRjx2E7X039vMRQUmS7QSGzIDE+X
x4vvy3G2uVvBYhL4OopxiIB4f2QST/iEndDwlmjtrdI65mANBRbJHjcWK8W/vjgs
OH7Gz9NQfCI1XfhxDRAqZlmvD9fgFEpLtZUdepJBuu9r79AZOWw+8ez++glRkdV1
CZjbKXqfYWRCFR0urDEqxH+vmMQE60vBOK13ZELXiN+B+SAngWI6Iki8RzZSE06V
Ffum/8LuZfLINuCmqRmfq9sukGCqoCGD2qaEp5wiRc7x3uOtC2ppnq1T1W6aK6Wf
4EgVsd2mUwGVFHPy75BJyq49tAe7mSUDU1tMxF0Rtq25XaTZwr8H6jYhXTiHhf42
zBGWmsPnm6QLlK+fJqDaN6h/uS2XiDeGzTUGJobCI9QmKtDvXJmdFB7IeexzviXc
1S4eAF2iHRuh+RonEXMVwuinNRKPP7zsXNxUkRNw183NWfBoRKc3mamRxHKDf4rn
2JWsRdAFsRA7siTM/e2cHLwkAq1j5dSzfkXyvQVbteAK29qG1nZ3vtexz90ynFXe
peQ4tfG064HyCdvKqrbuVcJWKquR1TDzTe7mUYLZvQEzHyOsNg2/DjKtWmqqlHKE
QrZB1FQksUP/Q+PWIgEQmtO/xDkgiJK81JR0+cQNxNfF+uRgQ0G8dUKBgDVY9g/Z
zRpZ3X7Ttjm6EGSD0wj3kBZ6SInTQHUtY7XsZBptECoszXpAI7QcBUIqsDyd0Uv7
S1Dwiupk7Rge29nMziIJNCRStuoUQdUDCCJm0V/kA22KtpD4XXfF9sPZd+a0708n
/TAEovr9YbdjQzPaAUQbNZ2SFqo6vxoAOcVGiNtHzjFvgUSM/prb+V5WkgircBN/
ZBfJ8bnSA253hAWtCYM9sYvPyGUBMs75OnbMUR1Yd4Nw7Huiy9Z8IXCdY99m1gAA
1L9HadSg4rW0wSsUtfNtWvAvi9qNz8yB7HEHeaxcVVqQdHacRrJPQFzKbOAUSIFs
coptKPeXeJ+MnXQcXJpmbIwpWFhvBfx+cUNUI6/WJrivsF/2wudpkMYbFAaBG471
iwihJjN9aEuWW1lyoJEaoik8TYOGAzBOqJpSEhKzcgQ9AlE/seiQzQcbteg+CsDx
DMoF5eU8C/jdx8DaQtoD4mLuyredE9FHLIgjnQ8OvMQ9HfR9NjoVz32Pr0Jkkhey
tW0EL3MWleV7rjtuUFHPhaesXssnO3DzUa8V7ICWuRR0CWJHKgTT5lDbSxfWrtbX
g1Fx4cUHLjJRzckias/1cryf93+k5zamhdopvZHKFWHcZrwauzazq3BfF3TrcM9a
1WXzgl01/ZypuH8izXnu5um1yOQMJSvXDC1Pntm+RV4WYOG4a1vl7gFN0M0+8xnT
oiZv0AH6ZULj7ohCX12Z2aJ4irwFwcMEVzfmZtW0Xt5gqncDRdu+bOWW8Hl8t/Zw
hZNUrRZunoq5mENzkFAnWVhIsBAi0jMxoSMRXw1+inPiYIMMyR1wl08U6pEnzrxF
wIsXOpJPBariGQVrnylHmR6AYckHOf6nq2dXqSeTsQre50h72B5MzRm0u9678hvt
fuJhxySdhQAUzHoDmlg6g3Ir+BtyQfqa4Yxn7dD6boXoHhwRDcPDAoqZIIJlVwIy
j8iwXosko9kXCxQ+W9Podd3zYHRS/eO+W2Va5z8N+N+Ismcn3al4Np4UFikXB+Qf
KR6uumujZKUHm9laruZb2TIMQe5MF4V+fLl8C4DAGigZwospXroZmXzVBWNvZOW6
v03e1x2jktlfY3dVOT/6R5YJcWQ5GfzvV/UMe4p0NJhit5WHkwA4267kfPFwq6cF
L+hHdkCRZYz1ZbOneOtbxIOUNtur/0z7zunYPeOPsAeOGiE0J1eaLmdLN3sOiXk8
mbZ+w9LoBbh5LxDbsXuBiOVYwNDtKxiyYzweFB2rTqhM9RkCdLp2aq7tavdfhQmJ
gQMlMRTRohLIzqLCGyuq7SHXh7DXlEfHqXmeuL3SVT3OWJHzMKUtCGNCdxQPiO4m
bopc7hG1VDfXgjd8KNGiPszV3MYB+hib4loSrRPoc/x0ahtoFC98xDDOyGHLZhJm
HjLiceX4yGNbUi3K+PtAjlfngXmoUR6ZEUCXekVdT5aH7n0FVzic88PMEjfJ3wEr
JxUiePNYGmloHgJweBCcJQcYQurjDKFYnnyKimohsoA3CXzxawmPZIYHfaQWNri7
Xhtyjo+KCGadE4i6/jApGS2vZ/Q8lsHZFzPbOUbPFk5fEsgPFOfeF4D8U89rZ+/m
2xyxjrrEl4ZjYD4beSjCEQhVRAe3QvtFno1EE9CTc8qemoNBIpkWm26ModS0LOfw
5qEtSmBAhdIMBuxYgxtp8c8R3oYfQjKPUru6/3cI/61T75TCQZlO4WFgcU7ZefA4
xp545ghTOkGvU1mZfdFsc57OM4uHX8YDv5Fxoxz8TavB4w+JyCgpc8M3HFwmgDK5
uvNqUJveQ+eRSrxe0U45rRXkq1P9VcqWKG9mX8FMKVxEzxlnnjBgEXD+YskyfKKJ
r7osUYQ8SGKzPzgCBi3hfsr0SQxXzBQHVDvkQY7F9ZqK4mvQnqWIz+mmXiB2qea6
dfioWF/COsAW8pIhiwJdI5FbkhXveG3EWOIGgzAUM44KrJVO19LPCtaqwghBES1c
v41jDj2jjLClkfkMmo87XJwGbbG+84VmW+/LJ2Me178uzaBOArmbC112dtTSz8/L
kh2axx7qcMgUvkX9BkX61pANIoGA+mDTEayKL1iSCtXgq4NeKF6X/qbdI4wjan41
r2FnmufgBo4+V9c1lsOFDpLX/1MvE1xB26LKdZm/SQcz9xZildC3eGaymAkfqHOS
hHH0eTXEdgPqKajICznxni1yWB8wt3VaxfpgRffyOoQh/EoRmo2tKyycnhvSEuGb
JhFd0vDrIcpzloBK5cTChZgbcw7K/plFqCMFqCBQ1NpAkQTBvU+e73TXucXZ7ra7
9+LMLxaRHbtuvE7AY17UK0X2vN5v1HxmhlNsHa1jk2V1WLSISyfoNuUKmmei2IpZ
ja+P7MjMdRpzXpu7/IpNtyEgDkOR9hecM71oErDX4DmjKcPH8B8yGoPpGJIcYvq7
kN4MWXOWrzEn8f68vR98clyv9KW9Vtnig4PHv6aZXAfhyPCn6bSygw02bdLTmBea
AQZBQoiKOt8KUtD2FmK3DUplU/0OZgNR5M3C0GGmC4ixhQPr5C+2muE8p5A3Mr5/
hs0LNwIJMEryUkbUxolHpqEn46bDc4K262L9EPGj8cmvtBCn3FXSMmdzY21to88m
KUOSfSafl7q33vir0czCfCRrzjwMu/WvK0DOW4NemI7OElRAlLsfkQWOKJbYZUDA
3DDA6k94jh0NT67pY4mFMdHGuh/CNCgnzqIzVutAdPQHHOlalRDLQl0s4MMgnK40
70GzqJUd3FzDuzyQPeat0AIowoePN2/w8Qd8ic7TSXdYOyeA42tJrgKSqyDdafGw
iYQ4zRIRlDIzybbNBIOUhB1noYQRutotsY63JUQjlEMjJb7cnWWs1MDdod83FrP+
wktYAUClKmfNHPFhejoOTQki+OHZcfzAoJO9rT+ioeoTRk3jGD+AJF5WUqdaGkWA
E/fB54adj1tlyYo2WeeBprRFpC2cVVYwukkwBs5GPX44o0zm2tlDlpdU+DYkhPuL
7Bx9ydoNAX4xI6pR6b5y7zGxnj583SDmYt8Mz48Dr2ZCFk0nMS0+vby1tNNWi2FX
/FNyFYPsNoQgXnwMmii6ECFiJRkK3/y3GA34DDqv6rQMdsV6fzej8ftQDQYQY+6W
hTyFXrugeyA7MCi6+AFO7+uXevivB+SerJA/mXlam6H68YnwaJu1oceuiSNjZb9h
VmUraybCNB/UtOXBiFFpdZxTJVgpT0I4I10OVFNYk5Chw3ooP5o9Fyrajy6fNwF1
G1ipoc74k21EI1LQ24zha+8uqxCzDT3WYgp/M51ZsG8+AKxAoUhIouCZwNL6alo7
jKm0yL1yYE7UZkecgf4dNyzMLAPxRiv2iNP5Dqy7/BU7U3ZAPqpoMwDCQ3jZ39Py
lZpKgE+1eQn7SglaO2O91fyUPqXYqg3gTCfXo4AbJ4neWtfs0A7+axbXiMdZ0jrY
OcSylONXBZvjtdipzMAfZUCWwclHpl821yW0cN/f8moBKTINR0zcm3tSBsuKQeoC
ZNeMzt2v71NOJBePeZTORUXPEAjw2QVLg++tSK2UvBrdpkX4r9ommTkYJGdODVVd
Kfys7HXiEyy7JySJDOxOz073FAKRKmiw1+7rymlzlfoMR6k520MeJI2FDNG61SUg
zXm8RVD2RhDWa4gWoQH5VpBHqz+TQT3XFNIWNHe87sSfuiGjA2XkQPGFg77L6LY5
Pl3ZXaRasu8Dup6dMEwHFSs/SA5SL6GtOWGGgRLBo/tdAeMvDiQmVQ5uK0hrnRYT
ODz4ucurd+RzHfo+nB2tqTn9nc2RhtmgFwDAky44YaaMUg+AFD3s3//dGZ73bXPg
M8360WzevNoQGTkkJXZp5gOmKEDtsDG6vM9l6spq6fX2Gr1X+ufXBW0Hoz0OjCK/
Y4YwfN+rwsVj2vMaYIQxn4mbEj0FE2nyuRM7nCivMyaI6NetjKTiYcbX3mKkTo/R
6d1rcTp4u/vuMxoyTXtadigPTzwGDzVxTRa+TsSUgDJ4tZ+6ToJpXgGO5P2eEVMq
aWygfGxqnlFqF+WHrPKYYv1B9rcSOhmcfQwXlBhGq7IAAuhnLIqGHTD4sri24A0n
oD0/JEiiQSAZ0epwvH4aj34MARTZJ4+5CwufR7ULHBW7nCnSWmo/tbTPlNap0Z9i
yn/5GCO1sKngFctQfw8XN+itJZ1vxv889/w+nNRDWmKuefiI9dlmgzseUOxyBjxF
A8QsBaNslkBt5qodfr9HUYR6FAKKBW+IsEKCwTSua8JA3LbpRGcSVYeQxxTrGH74
3ry+TtZmbfX/VQgVyj+MPbCKtqUe4Y6PSeJfO6orotIriclCQYH+78SEJ8U++JVl
LJCF4eXCvwSXykyWIdQToTO5OOKGoYtCSobkfzxcXCl3u78fsX7BtuDDmE77ss/B
9Jjtz17yVfV7q3Hu+BAcmWHuQ1CDoGWTltK0eKj/bnF1/xYIONsowYnBHdoq4hAA
x3O9H4Ys5hLahfY9XS+qba6TVMVFLBZjn1f/bE0AtEnfoONkVD1lGUzG/us22Mn7
GsGuSw++x8ceN0OlYG62GUwgkF5w0HIABO9mlHnb0bk+BXmgqdK0YPTSEh33SovZ
TYvEUU76iSTMTdv3KPuL1vxeo4S0+KefY/dQVz1QS7AzpAH3XPQv1lutoIZaJmEg
1lqXwzH6cqCB8A9BElw+IFNGcdTYyXyvoNLoyZt5HLtc3u6HNcEHiBXFgqAO+t9N
tA/9iEorTX1GNcGgDRF8S6FdhqaZoIZ3o6mZU0XYp7PVfpjD0trN3nnSwR+bLL+B
xvA/kcbyDCfuF+r3wVmO+WASRErmHLIRpAiVnbabE7ximwP2FDuy63bn+ns/bJrJ
6GNYsF2blNCg1cXtDjZJfof0niPt10LIsb35/4MFCMEeseDsbXcAr2EMfuVVJqrZ
12gH1YAalkxWrDBPjoUmbW89HLiJeGYHqMHPB20AqShVr/6+14jkshnYCyeIyymD
stnTHSosZX0ubrKIbvY+vUeV12w+iESrCOsaby+4SrUErVipfq5IQlhGTQFR/Ymn
OcXdP3HvIBbuHEEK+bVWgV/tDkWf+IjSidmAe9l8cH3XvTcmXOyjZ6mlqExKGjfG
sVjU462sngQHSzvGp+fphYMhGyAPxzaalEmPv0H6XU767tDtHUOs1H/JNrQCyUgo
Mt7cVMgoWOO+hMW/qS2nB8boLeixtdxEvpKb4aNt1lRmI95ynqT62khuSC4sK9P4
t8//+h2qjF22NML00j4k1AGLE4MGbJO8scqMidoABAZJIoRP+o+gnOvzdrRaoYBF
5w0gbx7TkBY+yI50y+P9mU2LgDlRfoj9Dwz89gxe4zRmdb+z45u/vByERrbeb1vy
yS6f0KHX3sfK2mg/HFGxVaaQBSlrc5N+Vc1FYwHzuaxDCQneBIF2jHFWXewyAOh7
eVZzlIl8y5obP4wSnCLuNkc99Jff8W5TcF1ydNCkJpU9h+LHiGGAqSYrlU8ooRWh
JLRHudHEIG8hggn19bOhjxx6Lw6a5pj0i8ZaFFB8YrpZDxt6nLPUpj2X+KyljHpm
+eSSWOx7P4ZyomW2+5dXibhetBZGG/qJNReuRN9l+lOrPkNxP9ZDI0sTNQZIGNaB
ssHZ64rIjBnREEv5CeV+Pi8qqr1JcedPUzl9ie+tFa1/ProqG40NHrKypE3W/aZb
YVba5NYc90ZcjhCybhDdTEjZ2tVt+cT2bl0TgCQ4nt+X/QhsTjGMrX1IU/3X8g2v
ZM/1rFSGWi/BJeYeDVHe4Nylf+Y+7pfOTdMPwXfW2L6bwYygmXntTn5wpJMm33O8
2kc5+wTM41I8lopgaDSlYtjZrjzxKnOUZoEwN4k67pXXBwBIWkipO35ZgYQHIpIF
b1Rgw9ANFzDZNtwScgVSWw384AZM1xj271GidfgQwCSFMAJh2el/jwDEENtBcPBo
+AbWfHUp2AP8zeab5wzMBMvGAXGfBNYGC6GpOh1yrBpIlQLajqyXcyXPw/OiiS1b
IOBNP42wj2+R8WIjGuj9nKBwLRzdrwS4TWiiMJN7q2a4g4XpWl/sqEBjP/7sIegU
bkFolMLr0FYMLC+HFKNXj9X+7sHZ3hAgI/SKBoyPI0WxBSKKw2PdPcobXhvQ0IWM
x4C63wRRI+p9D6ToOiftHRSkxWRvoZyWGNWu1SIC6XrBdoWftiQ/KVNywp95W0SD
HxUX6eEDTFtjQdF10gm74jdM2cVyXoL7dhj5vTbGuYbqbeaC7msRxX2Jj4XsHOog
sA3Mj6oEIIxvF2FC/bKmTJ/x0XuEO4gugAo7tUOV64nZkDmOB0QID6l0O+h0AotS
Oe67I4KrXvv0KOpx84jHFMJW/uPGkizAw0gH7ms1Cgu2wYnONTuu+5U15XXTbnz1
TLnaYe303pZOeW+OC7xWjuZVG1MxB0yDfAJOfVQPATEydp07pdPHkj2JiF5jG16h
Bv2GJ2gWy9HOfU2ht8N5TSz3rpzTYN5C7MwyynQE+d7K4FVvsumwzR5i+LkV57D3
WNFuAkPIRIRPXENJ4DhLsS6ojyDUTjyB5DjaC7cGIQ5J+mBEaGqf8Ht6pA475QjR
d/hc6rC2J2orSopo14asWClXFbeLlrhvEyGqe41806sfWzJITl+DssT3T797XEuS
0/uogc7ZDdsAhbVc9shcbAydJifCmRFfErtui+/HbU4C3V69ll7fxlNaU12CoxKn
P9dCh5FKUXZktHJrjTCDDC0NB1aabg/CAw4cp37SwLfOHPIkJd+XDLrBRitbG9Fc
stqYvA7IhMg2JfngiM3e+0BdZJ7g6Eue6rYCDc5V5L9IshGP2+yggdyRYfhL9x3Z
SsNPtxtMBLCHPgAgddhhBRgZQX2yJ4A+eqG0UEG94NUU5sAVesG4wq9pAkuKOyUS
JI1qi2nhMboDP2vD8Nk+urElcsAKWV0YurBnPbYd3DJp01KeDAmUjKj7P8acnYgu
BKDN4E6xivkZOPm8tpKUeLPluf0yvLo6uPii5dDCe33BiZlppu4qSdZ2iJKFvhc7
pzgVypgXHZTa93zKThJx3XHlbubKQE6GfldRuJVPTEkEJkGZ8gx0bnvVcDAELOQG
AUzZ0G6iGyHYxZIUbLnrAEZ0JiMDXFjzmCGz8hA6IiI5x0rZfAisrl5/fd7hX86n
EfZYvCl/sZGRG1ljSBuI5XlMHoz3LJqKyUjQfb8hiWdS/UjKV7SQ/0d2Ue3aDD1h
/M5yOdl5G7LgZLfMtHaV6/JRdzbM6gB7np5fIoChz/JGZ03+uGq1rSJIa2iCO7u+
hmGNAXGXHOCXAHm4FNClqI/J7P6YcqID4sTBIh2nibje+lCDKnXz7yXf08RF0ThL
DZievSVriaeRVu91WSkAjKlzyf8o0kBlVTmYU9wdhzjBXa0JvY/Py5PPsvZl3sT/
NCotdqMDrQMlFyAIn6bQ78Gi4Ew5m3aETj4Sc5x/mLY2rk0fpL9AL7x5f2m/KGTV
HjGpwYkfDuuW6SEkpdZTb1gnInbRPymvh3QuVFgUv+cJYUbf9yyiU15KkfgNqU1f
R6yBL1OhuEcNvb+9WbtolgNm/aQYrEmC1iT737999NgzBfICZImlcwlAo77ysM6g
CfsP4DkCOEJYhrUvzjmp+1hAEeBB3Xa3MM43HMrtx2mVcOL2Axx/jJN4zGCKpP8n
yIF/Mb6NCM4j0PTfPKfKmmQ/HqWrkbXM/v5FgZMySLmxd/LcZ805Rmh9FID7oxP7
y8mNdN1Hs4JUHPV6uW1sdL8qNr991Oqoi0Z3tybJ1iMSg8I2TLRY1XY/ub3WhqrA
tdxE7iQU2WBTy604LFDsmROyb9DMUZFt8lXyiVqCy1QTX6oVLhITzyl+dFL70nR2
AJMRvzIW3nJ+cKgmNp+lF2OKdP6Mkhyvmlh02UFYy39hjaixXJ++r16NwwhvZYvm
RTjMCXEUziGCE4ZVq1WGoemyzUyCVaHVCJ/2N/6Xylg3yIFQKT3NMn2es0yOtFU2
tCM1XcjnKWFaW/pROebMSIaSoWOIM5StOyurzTkwWesEjmo7AS9aXFEgw9pE/m6U
9RVnkra0liA94/ke/rxn59mRAYnC/kxxvV9EZb/jbvtPDkpKpID5PyY27ObGH1T6
6oKQtdar9czXzXIOhmN51VKorQK6R8etaPB+CdhuuD2iSARPIkWP++xXOmunNZFF
+ln6i3fwbKZirQyl36VALCI/p3c185VHTb4sXdn8C4/I+ZcCCITNeRt31CqV1IfI
/rRnMCzMZwWPrTOu7tIazZPmTlFRbo7rpKjhTZDO9uemMTGoPwsxH4fdyyl92Vws
xF/wPAkaechAieF954Ho1wsWqigqQAdi/MvM9ys6GUfqD0HVnbgFSuJEUnkb5S0x
scYuAEOt8M9GuEwDlynDhYRvCj6jw61YHUEDnenFukXQ+TmpdcXSDtXYkH1AHYjn
NsKn7cmXiNmp96ETXYAvxA43ySFLquusTLqjF5xwldTCxwTYBIV0NfcSe0q2Xu8C
zTjUYhpxLBRvckaTkR7RWthckmIwkFKzWSu5sfRged5WaP6T6w7FTX/hWMVJpbrA
bOFXcDuhItrdrsKQRfXqreOtjGjxxfHU8+MTkm3rtJRtbkJ7/bJxmNbfB6DdwsO9
vM4nru3oVe9TIKTgpZqYQjouBMMFCpWeIXBkDwdNf8tqxfgh/Xt3tNBkuVcaVHwp
hIAj7Nxn4EpXnQyusqgChInBxp4f3HPSYhepoh2GSSLSesSlSlAYwRsXzg3CVWsv
nemvoz4W23tw6/tjZqAWTyVp64s/8lA6DyhScf6x28DioxPL9OqOaoftBYTDrSkk
z0oMw29CXzxwWIJFr6ME0zUeIGbBVA3LPrniyiL3QbN/Yk1o2tJKRhPJMhv2sOvi
U7Gmj/UqBf0mlVdfE5z8VBNEC/u+P6duD1zmGqJ5SczUarFflPt1j3bCqT2uZ2JJ
ZMOqexSJumfrugi1yEQPlzXK/m2wqKhW2eWcOs0ewDcauOFuNZMvenuGlJFI/mmP
psIWJqy6YDvIUnrkPV6rWATzyFIaB2bgdERXYH40UPtPPTRxLzjWYsyu8Wvy6Zpb
qTQEApbGc25opISQPISiQgMDj2oJKDDCQIV8NXvVmRb0uRjxbrygkObH4xOildPj
HP/PxlnycvMJ3nSW0WMaB2/ZtDVryJF2fyvQIndw/skDhBsJUsR1gukip8mSPBRg
4LuR4bU39iz2tSQcMb5DLZNmqwMxxJeERZ8b0adRJIYbO/K1nc0UikT4DvEVZIk/
OF+BJvO7u0Xr6AZie/7Eb6byK9tgsG9/DO7bPP9vrX60OP7/EgoLksf7j9YUKn+l
Vjrq6VGK4SJCm8Gl+Kv0M281F8FPQygdnBRtNFvgj2iKzh18FLgcx1BMHlOHYKeX
GEh2e5t4i4hLS+2bU87l7tqYP7okjIFsHaZOXifvNdw0XakXkpVTHTLSApCendc3
8H88TZHg66vR1c52pI7pzLMcMm3LK6V71v9AhhH3cxD5fJXhPuls67ep6ROjUHxE
sSBcDKTWyaOxNpVENptIcFnYUG+4H+onOQj0zxYFhZOVXkOg1E/gKW2cVG1JN8a/
LaYiC6mdHYvSfDw1p3WNlcN7/TYPOd5I2GuZPsWLsW0EIs9YpXmeSJtSdfXyule2
gxfBFDtDTCH9w83XL85cbPSJ3+vCpGLrspKA0cBCdELoS64httH/wINdoEslWIbc
951LgHYU7jSdZrFGN66ETj+9oh6IDdB/p3/BpHjjehy1/hHy97vOoM5Ca9ImJWRY
hi4TDzoJeh5oeOHEaLn/dbRBu4g7JyyfHxZRhdaEkxEocM48uKYYvGcfaBIllQyi
CyCyIeUcbaNkO6aD44g9AmbdFjkZr+v+/9cPWsjbZk6WDBMHgCUVM/wqWMFupqeE
yVFppTFgWA+DvczMAIYfJ+Yl32MpXyfF3MWkzQjZDyNoQ1R2VWWuFucaNQftH3Da
GXF31JWL2o4Lx9l0VPEdYOFH9kWDftl7QcjnVBztZxmBiRLstwajqHoqvDlmmjKW
rwNFEnMR8zNRXQTS4KtQ/Bevvr5umEVoaWHtCFxP8DdhGGSmUUarcqUwRj60A01i
PWAoZSS02XY+kl0/ztscd9zLa4FTfGk6HTRltqy30tYGgPEeiALbWetth6pNrcyi
p5AGIBIzCdXlL4ohCRyQ4htgNp48UbFD+eWbzgF+vsjBWi2AKQS6ytkyAMMGV+vy
eaPE+BGGJ4u9Bb+ndvm9ye8+AHkXjJZpZxtPgmVWUzk4EpQD4mAv7krNOjDHZRfZ
xpG7cbQiEZTwzQ2K3lQ0x+fhqNr5e6nZAEHid6ZbfcYAEn9UvrJT5S4sgTS3G6kr
nq1XX/5UVoDWhKH2RGmAAcfugXGX38dBWl4lXEixPzKCaxmdIWD1qbnRUXSKOSZw
ZqrK0ja2uQc2mJuInOJOQ5aa1iGigtc04vnLXwYgThO2FLHdOCqr8VfzT5Xrwrgz
zIbPpPaXvh9MIvgC8rmSV7z/T3y1/C8MaeQluG+X2/NTMxUxBZE537ITvinEYW9f
8h4a9gdezeII65ByRZX200AK9MIEYTQ4dpb7jcCPn+fyJwlf+K7RV73aQOzqqjic
R4RPbSdIO0E0BAHhx+SFgaUXAsJKVG6qmngujeuck992Yk27nM+46KPViNkF94zK
apPj29cru7dQ1ciQ3KMzBafXIXmmC4l13vZhkIaK6UQ2Q9BM3/JXhhFn1K5pbi3D
mg522aHOJIpuI6qyWwd1rUrg4K/cmJX/Pwuef9opUDgoq8HMiCR8e27GsVufvBQF
05d2lf59oalkebgOd5vpbICKlag4ardWbfrc3b9CGy5iY4H/OGYWjkA6TzIvyW+f
e7iOpVzZCamKykBrvsK+5gw1ReMXs9LBndZrO+DlgdUvdSdzxGIZXnKe9SnJYR9k
NCXafVRtCfOFE/pG6/k5OyO5UhUU8+esiiFhwgAjExJMq1Xv4ORtrJFpOqxqrzg4
7YJ7CDxE4eBsma2FSmzr4Rz6lQBdWRRLjC3pycIDMup0gQUkg1FRiKi/wuPkoLZe
p8LBq4haCrcpYDV5BkYnSKjMqb91HToRFiVEDxRTb/ofhXCuB1TOJjrrx1m5Xaf6
a993FmblsfU1cj5iKUiOhqimnIOzBY/ozm3jlQR4Q972e0AB6vRk3pA6RuD3k96L
28FiqyHd65ptggKGsUW8uGgf3rO0gatMYToJXex3E/EbQXD0UygFiCbhYWACDjw2
bLykVJEPJO/OZjxjKpe1vGMxiJk6qTh98kjau/pLALsebeLPr+BHAtTtlwL6bMON
B7b1VhSAIjAWz7poo+LoSylnz5DkcrDNieHdSvajsJClGmxxum6pxNgM8sjL6gO3
bxg5n6VstjeMESCIiKlVnEUNSiTH9cjSUBN4yMc8FaJriGVvekHaVjt3ody6tYcA
P+cxzk3rTQKBE0XGUS5UaFiAHVKG1eFZVUeJZx1geuD3tQlOliqrlirXQ6qS7Ijq
Z8QYX8WOAFoHI1ZkdUbbNV+2MJRd5WhjagarXNJClIwKae5aIeN18XKsGJNxmy6e
R37oOsZ3qxRrVyClrM+ImY2oiPTEfyrImDr+XVVYB/ZobhE9vKpndeY9brIUL+MY
mYeSmlXLbuGw8+bGFygvgkHKE9rN2cu78ZTm3N5bORferLJX2QHNDSd8CcWDkWbr
ftS8uNiIeIwTaAXR3Rdz13nidHVgxjwJhHuHSYTrp+GGUWL21kwZEqIJTJDrhoNG
rsrTtCV2kHzAUrWZq0NyTjhSP+fAjqD0J9BHNW5qaVtLnKK7tmEgMZSsfoaJ+CuJ
KOQUpJNLSkYkMZX9Ee/6atSRsM9g6/HeBov2uAn7XWd5OnvHm8e74Y8lnfU3+6Gr
IGdGpmySPIFSnZ9/DjRPSqmfymhdpyK0ms3KZ8RcnxBJWNZ0brdirUYMz1J7RdRA
9+rjerrDa2QB4JOEaKni0fl9dh4ZIf41eb57neZUYpcAhl+n8AmRxEO5e+t9eZgP
IX1fnlUB2CBwYRwxIfZwfMCFnoHrjl0525unnAiGrQI2+6/tmbYgQvAbCFyO68No
TUJX6qO/7qoDseGBcyNw4AlLjYqYtWrgM3rTm65M5IPK5vVOtYNPC30HeDLC9saO
jSxZ0wBxmM7hug+gAsWVgik1QHma119po1q+LwuJuIgCEfmLjbAbiaj+xnBU/STZ
/GI0gmfdo5C1Egptl9cI+sjj/lYLrq4Vkk0ULMpm0XGLQjUJuFKHqqr5KhRXyq0a
bAgFAsv+1PK8wbU5P9/S33hkInTPpmzrUswihqn4zDSpupXHgiH6SQn33v6kI93i
Dd3TCmjRI/BK2VTbCtexIrTruXkwqUyQnbzEnyTltZG9oV15mrKFrHpqFIPw0s8G
Vk7mRijxP5wdwE1z1UP1tou85gkf4eJPHCvY/Fx4VO1XawqvwDTJy2ejr/bwW3rN
hYQL+cVuUPbVHcFG1/UPNLFUAwh3uDreml/XpDcNHQ60DR75nCyI7TQsJi1SxiRt
BMF21LxGIvx1pGzGKEBRNgiFLdi6yJdpu0OE35g9vjSVNPWz8BdN1Vmz3JnPaeF3
qFCjErgOegvm9PODqM6vuFap/evnQdaPGEw04BwlpNUq31TZdtcOx97G4bwCL6aq
nCVUAvtzSK+Fmu/Q332c4Y6sNx+1yRPR36xOS2l3ghfBr3567NLQNEU6t1qxrvKy
Uwhxp56Ew3YUkGxyyHQ+JBaPJ6R2Q15ISRR6lmU75hHH+IzY1AaClHZ4PbPq13Yl
aEyjYmvxrYBc6TGTcFqPlbl38os3FCexy4AqCYZbpmty3bObRrd1XWuxUq5ASH0Y
vjgRN0CGlvXe4QFOL5XslQWDbK5wxMRfFMRoIxKyTANhqTNAIc9nN6OCPE18FU6x
vENJm3GAXMDkAaAG/n2IZhl1RRUrha8/fDXs2XSTx80G2zfUqcLTAYMChlu6A/hN
4mBb+sTbwKnd+TQvJXW+2u8v6undZKoswdjAWMOvSMfO5DwbgkJ4xozQBw0tvweB
bpXHaKsFXYICf7+Jnudgp1PcA1rJV2fHOC+nkO1QZ0Ij3g1qsQeDOMWxHs1pMi/L
bP0g1S3hQVqlhBx4qbOUCM2jSad4A6UBRSqXHhz0ZcMPVchKM4zZzAfmwuy5OJyy
patZS+IvX89mWcVNcz8C8SDJHIzfb+RKmxaxexpr+iGDJh4S6OIblRox20CqunJ/
vnKYoxxEPA0K7B0voKon54A8/qSTFEkY3Iu/IFDMs+4OfI9WJx/Jaf3RVpt+F2h7
82IposQmrSzdPuksj6Fru9//wB7fuDbQsw1k+T22+QItSpWmdPC+zYZBBBJ+vB9B
aUjB9nsCAUcA0f9gUiXM9p8g/dmd2hKG1UEODEE91NousvHcGmQNAQXTs21sDDAc
IOvkG/JjOmfAPszYMCjJ0JVtHtenvHiyIjUgh5yA5BnrqUkWSUvUfIwM9iuW/wwN
xNua5hlu88jWwwXFfdyKToCyqOccUZyD4Lcg0fd/BJb03l50BsFkICy9RMPljrj6
EP0/4r8UF63PuMwf5AuYrrpU0bmw0s/MObopo4dHeUOWFfSdWPPnPog3docAWRHW
8b1E91XmkCVerxluQScsHlGhpFtRVBeoMHzojoG6d0IqpZDBDa8bWa3Y4nWwztTh
e0p4mAWID3FZVXtlVmko6pX/n3aRmfzlqIWXu6DlDq5gUDkvI24wcWWmpZRXZXkp
0yXW8oDWu34b2d4LZ9Oqzj6uBgn4IgqpvLyj0T0g8v0/3nF+ZHknRFIyX3+80UA4
Ky74j8RVyhKJpqF6Kiylp9RDSQ9rnl1SUMDJDxYLPdE9yPuXqSxvXkC2vO4MMz26
o5kLVHl/2OHvkAIbwh3CwcGKMDWtNueA5MkbZFmQS6WRWZRz+xzK6qbye4IhQKN9
X2aacawbrZtxIh7IHPjVpRFcIr98KFpunntUHvKEpuU5+EbSBFacmrY2sIhrwngf
eyvFiARZLoSmzgP4O81JfE+zjSM6QeAa6or759ymGcp73HTvmoYXe/Xu5pCScXTv
cGtzbTQs9NNKAxlpO9sCzY+43Jdsb4Eya6SL7+HRqLqoLoUObe/U7RpQISFjZe2q
oOyyQ79+uAg9/HGOKJSsNWB9L72fEwwvrf5SumU0j+Q4VoY8JolpTuPSTgIuAw0G
CYtM9LyBTxA9zgQyibD3XubeBgXdg0VmhilOLPQki44qaX0SIWLTxji9jsNhfJPh
w21DRW7nLUt7IfiVpV3PzeZzipCsXAH4HiDexUgZTFwsa9um6KBQuge6gIVCDb2e
utcmowFV3pU+FD4zQ4pQR+jiBSQI3euDbowGe/yqLvtnFJCz9q5FipWvm8OEpEv/
lel3xSeatYUEottKNxADWgs5kBQRCaIAeaLYpVTvDi4Rg42oT7QZlZLWs0spAUHO
6x6n70B8wO+PvxgfzFfg+4j7fxAglzw5Igz1ztoEzoF43Cuc6II+RFS6FxM1/cAf
34xUsc8P5ovD+GBogG6mUjI2n1l2bYOTPU301IV86Yb44wb40cA+RKqB1pEPpaM0
BGZc8M2UImYlbsEH3S8ELCDbvXaODC1EKqiGc2mW89cp6byJ1rO6OsCsfXBYcTo2
f3INv2YafNlJn8p0FPnBlH6gZ3TbTtgQAg6neioz9Vi1LhhfNJyOVbdmCPuVxlJm
WVkoYJHN1m51wq4npl+A7XiuzJonqdqeeyf6zZwzxNYn869+yz6HyTzQKZlMgyGf
Lr+gvfoI/YRNv3Z/a9si8hFpa7g5m4WpWqTwWzYKGgoAdV+K0ZQtOtBlBOKKdrAu
dq3cFnK/hMSksLWt/sbzLuESGtzY14mNeB1XZzLeqh9dYIRZwmTZTiwpIADlDtVT
mOmja0y9iI+GvYs0XTgPYYDIbEvuMTz9pRbQ8l+mXQX8lr/efBCdRJSsCqtXpuQL
DBdinZGbie0wHLa/vh+yl8boBlgEmJ+/VeKG7sRTD6sYHlyitj1QIitOeSORdXvh
bj4NS8X2z110R3rCt0QsIa1jwqWoRKRBjd3zVHERTRK+jD8D6A2sP7pOPJKO1iaX
kgF58961KEJzXkJaqS2S2UyTedIYyrfjxLuYEmxhK+6oJX42wpJ7eRV40Q7cUMhK
aj1nnInVN423O6Sj8mPHEgGbu2XxnNZnVbZQyr6if1CklwMRz7AVZ+t2aGBa3hme
b5RpVcsMS+5bQ4xGh+hJ8itS+eq4x6uVFTH2ZCozA480QSbDRAKrm6VdAQF+a5HN
O9WTo39/odk8wcbtRP/4PClr/L7d+KKouNY7YKJ17xiQcJq0z1jE/Z9uaiIubyNh
zE3E6cq9xHPgXbMYl2CTHRfu6RENbLyDUupNW8CBcJwKz2JM+70DccLYmEZ7FImW
+v9P1wwVDJvZP1wvl6Xyb1d2Goz/d1HBPa5t5M1rNtgc0Qh+BPgbPCP4lzCg1XYz
77D2+3L9UHnh4cRLY/u2cvbtRUYxugFRV2wBNUBtIx3M1up/eOK8N0VuUYmlI4Jz
RcLuMAS1ntWue6qpwbeYn/LcQLaDdl6msriSF3t5Jvv0CAUHNBNGt3zeRmAwIV7D
1q9kMIWmpi1yyMXfeLRsehFuYz9nOmKmdF7Js9iruZ2F+DnbbOW+fVvXiScjVEDc
I2xWNDJXqWQw6HwBlvWN8+JumPgdW3qCffPoLrPx+oKo9uUXpc0U4dDIi1TQ0EHs
Y1y35rW9BZhAVz8PXsEIncEuQuOml8VFp25YlU1gCErbiJAKXkGuQMu4NOqSzSM2
Fl5PFZpG228MiVq388iEgVA/1z7Fb70XQtiFnw1nptzK2q7yH+jYYG20nXcbcIq3
cNTRFpzKPrSnd5Nq2NgAAT3/FKFO12NRj40hALDDLVVGioXW4dxdQxwtqtk76REm
giWPvVsDmFmehawXIMkDK6nUdy31EPaBaHSgYntuC4DdDcrQCVSIVPoKLwjeYjO4
/0Rh/++tbMre+hlrLCD/cFvvCQxlY9tyX2DaN9bg0NlG5KZTkq2w6uAwmJ/9mrpf
CUa6QjTFjL0duNLBhZgipOu50/5tm0BBc8GUIpNdAkdpu+vWvkOEgVqbwCnK8NLd
4zPngkJlpj2IYiT6ons2j+8v9EKV23ykmO6VnxzQyp4julqAsEeoLDtGqv02pOdD
Lbb46ys93SokMWSozPtB19ggQcDNIOBcdZnntqFRau5nkMXiig1d/EXc/RXq9ZfH
mOso6iafeY+CZMpDjdwWz5XqBZyC0VfNcwphdV1A9QGsfauJxufxRVRsbI5RVz9d
5aqK/KlbKnB/KapcBSEqBkXHCK6TzuaKo0HS6Q43xhjLF8h38hsB4iTbW1aiL8Y0
EpXp/6QTkQ215Rf8rtg9sVISvlPtui2eaPGtmcbw7YyNfQl32y4jEYEENONbPv9D
kuaqBjsmxAtSxG9aACFstX8UzozXvy78CdXjpQnclZN9HJeiKbMbceUZ8RXAHHC1
b9fKveZG/iqctAHS9cwXdi5pZk1V5n+yFC6U57WKk0ZQwZtFUbPxb9fDtCK8Ssu2
G9+B4ShVnkhSpjP3oHSwe3XhXud18oDuj3ffuXTSpi+6jd1UuaPCD9mrxj8ULLhv
zzzPMiVBUAMlaRFbmFpwG44J7zzZEbI1oquQclvq4xsFoRQGrrI5iP9iVSCShKMp
myiDtNS11UJEy53F1CD+ybq/Kor2HpxW5II1Vz9hM8H5R8NviJbtytEqgDiV0GvG
+vNvYt1xQhPfWx9b3TzjK8LJw+kDDOUicBCUwODwmUGPcxUZMDAC1Z9Ajxq7ot+b
A0gggDQg5+1b/0E7sREy5XsCyUI9MiNkUfkGN9n7QfBGig6SWrBhPLHOzak2+Qbn
8SvG06G9lpyajdspK4jV9+htzU2ACe22dukamWTXz4XU7KZn15rfYUI+MgPVkSqv
O6/xeKxCJG5OgPvi/7C2I5GOdMjsPlIME+II/XAH2VSJqkiKrnrfsgzdN6L+a5Ei
7oM7GJw1wvrI/QMmjY8QcQXsasei4re20jqNfyTzS0kZoyUMsIyCmJ2V/OpVfjLA
UXzHaP9ficvgae0x5W8KjuIp94ajmdbQHmNt5BxsoUMnZjH9OE3avTS960NeZXN4
6R8ecYOZ4fNi2g0OKUD3Fv4VZEOp8ta2ZtTDfFILy5z9ETS3WxN6ckHZPNAd7C9z
+4J/HJO4ok5s5FQLqUbLrKG91f+li+1O6BKPrzRWLILd2pAxxQt7WgwjvjuT7FkV
x+xatXJKde9tgm3WzLvTEtF4voSx8mb1uvqCZUx7REiyZIwez8eAq5lVaydZ3BPN
YAU5AoGzgFHjwxlHSXIB3t5GVg8kG5ZxeIrzoUxDPsLuB+auy+FbsFx+6aJT5k+l
yAw5ZIqxJY+X4CCJWPnVTntZvhlhnlRcjDt6L5rPjcbk6s0OUhEmZO3VsM1gSDFO
LgObYsjkW6meX5UZgaT58XNMRXmndud5Q4YmdiCaW0/AMqOKSdngldaYvwbKqDVv
p/1k75x+x2poe3mVf/x8kZR1SWBG3bKMhZ0Xo82np87y2blaWwZJxUpDYZA6eCT2
YcwneL0YruXQm1LGJC7VmYKm+AMYy1OogS6Uk2wIY0jawiJKn1731o1Vv3xm1Hqo
kWhYobH9ZRDEruMlaTzI8RvUtni4vZ+3ipCLDsNah69HBtm6CdfB9d4IuQ9smf4J
UgIlrcpqvwb31ku4sO2FFC3ZBfBPJO9SbJ8Oh0isyFdBIx+IUzUugUFET8VDCILh
rSnTvzYAtaINOztrY1CkPfrgVe2fHd7SjiPyVobpP80+6+rzE854u/JCNdH2PSxs
SFbm3zxdJfdV4Bs+nO6RXYontov1TWb450Bg/iDYM2vvUnsIGXEjZveNoHTL5HlQ
cuBLfXo4TpdPZbZ8pvpOUpl6ICYvjRzixgAlv6YlIDLdqD83gCP8nvnbfwab5h1n
+VJZTQlzdTph1yLCdPUQCvi+Uo8OwNX5jaP/qQz4gBXELRc0JOdDBZdEnYMDt5Aw
BF92IK4Z4/BBrG5abDAJghjOekLIMYUakNtK2BoVZRzxb3QrnnlxPhSagNKjbZNI
fbAyQ88US86KPH7QEve1fEMFs68N6sL6PdlBmlbITGVqVnJF6p8N1z3PPFuE9Br4
dbatDIIbdbnrjcljomDFflX6MbG/U540AucRR+mqWIn8cpiL2uM2gZ65mCHQnlrg
2z/26PCY9zW5agGUv/Uvl31zvZbCMMfjSAfBiBjVK6B1r/W646gk14kqp11L30BH
iKd2rX/cu8jtsZjnkre6jGi7yvOUsLYuSNxeKQx55J73L7BOE1QW23I7sb5GccBv
zZIgM9mkFkshO8SpB4PewBFCMWfa0of0HojpTlVAFqOUlRMYjGzOnGH2H1i1IcWq
0BDyfeRb8M4C9vN8GmtGq0WdWURhyaxWknvC29p3IApmzJCrDJ0COLwBus1ydQ8e
IYg1IG6xHrnK6+77n7Bs8CVpF4Yq4otbjJeyD9KcoCazSg6FFkwmgjFTXwsFbxVy
mxSSQo4bnIhqX0+WHByPBM3WiQxK75/tsLj5iu8hbTRiNlymE+7Nj8xpCDFJqt+K
ZwhyjDUnAkHjQ2yPBw7c3gY56PUIBoFrD1wEQudb3VL82x7ggQFMbCPKiOnCIjQY
DosX6Vj7KYh8UZaus7DOq27p3cSxIG0W5dz9NKZeXR1l1T9YDOwnspg4eEY/0c4H
PivO8b2Hy0VQ6+IUjQavkAI/C9XBo5Wsk+cwj1oqvc6OAkJEP0jDupCDFJrcupRK
4O5Fxe/iDlXaDO9Bbd2O0p2qJmNhzZTLeAHrofkiJMUJnA58RL2aOiaDggOQiJ2I
9MVSRY4wa81lkmTUdvjSE3Wn1E8/Otyn40hRLUR19TY37bctPOHLe4inpWNtqY4T
9uUIAQR8L8Odnog9p+ZdHXRrj5on3BRkxRaaZ+CVM0HG9uNHtya5+n6OAzTosOgp
txIRKwJeAzL84zt3KlPap30Oj7FzdVFb032a7Ezpgk4YB3ykE6r1Q766u1BnxrRX
jmX/RNyRjGXEvFo5HgyNq5cR8CRyZ/wjwMIxFp3CMAra1guBbSr1NGkRhKvTb5a/
zIvjl9iIsXj+nA1rQ7fY8TQmpdLeJ68edH3z6DH6I8ViufCED60EKtUYyKwNPaN2
+QozPEgMPva2GNTHE2L+FMySqaJuDR/mk1LqBR1RrZIQ6duP6r+QXD++EI9beHOK
CQ6ikZw5fpHtnRK29yDyY8guXqIS+OqyCQJzzSMSY58oxBQY/YqiHCDXfkW5TUPU
8KitGVqWxInCqQKLj9nNvenBs6UHeQYp8DSVrg9jeEXMOgP6sZxgl+k147UHxnJn
iO7uZKsruVkHkvVg5RApXlI0qykXe3R2bcJK6EISAulEn0hfGFL8LtYkvYFSRHO4
rOH/EfpyI3li8wAbiZLBBwH56FLyVQ0spuTffjAXsVuL6ZYwHReN/M5vHVqfMuWM
z1FR/y3PP1tdkrJ2GCcR4WvMe64a2khm4QspA9qel+nOxeAXSnYmkKBUsXsoad22
lw4ijTsrxuMQUVGo3KXiNVqF/dO323CgPl2NWAiaQl5KqcBn2tX552QSldKe2Gdi
G8rLpgNPTPK/Ov3ApjnUa8gU5264nxDRPCXvpPqHM15KUjS9V+33UD5JyN+TwXCS
gTEtPP/9rP5ZJ+rJ+ey+VZl1oZjrBJeW7R2ZwIAViXIIqoLX3z9B7Ffk19ieClrk
BMQYWX/Fp3JlDh1yJCq2EtZrm+7LxnMp/XvaOZOGYD/ZNc0CWbFhQYZ+wbumB3yL
ve6+9dOWsk3yCQyyNItzasbz3ScSM1pBUbzNM6oan2jaflXoFnin3YdzbAQkEEyB
c/L0aN02EvdPv+YfT6KvBUwejgoRdtfbAKDnxWEz32a3kestOk5iqiLDxwSyHoV+
ckRNCrDHsuj7VP66zyZ2Cq9V3iO3Gnv/Kh8H+GefuxBDT8eHRmpN+D9ZxMHlqLb3
KYkJQFPR5dknF8sW89CcZnvIFcp+DhyX6u9ilv7SyG/Z2235+6RS+omRLZgR9swX
wdSY0tSvpo7omlseOr835hWmxEJ1PJCXagAyq7NaE0N27BqPrWSR2GtqwmZ0dqa4
nYQeH+mte/iKp/DjILKQ7fNfe/wsmu80jth0Tp5hobKUaf4YdW8yFJktsyNoA+tH
IUqYupm5pdme8CVAm8DPjAyuqMFYoQZK4dcywYeTUO0FPRAK2P/9ad36wJODJ6g3
2CNkTyL1oc+W0QX7aqnjujk7mDq0N3rl25/kPGkWnwq+eiXcWEfuCkXP59G3F6Kl
Q9HuT+73Qs5JVHLYnx5Kn6L2kToYOh4RiW0Jwl4ZCPVSBrHUdCIFXfhYA5f3Ox15
iSevSMuK1EFoikm2ZaKeVDO4tDqI/yYvcA5tH9pKPl2whuBlCTw0niE+T147e8sq
NK5Vul/D0yuQ4cJc7p60twmIyPmEBjkJpEXKj/+jlpMMJJKskxJLNvjsPr58WEq/
71S6UuIQBdBgNAkXY1QFYz5ijODb59mg26rHyorNVAAXlWWWDWjOZPa9Sk3pQdKy
RRJMldIl+fokBNT2Km2NUvOgA4ZcjBNN7qaplMxmRnkgTS6TV4kkdbmVA0ElgomE
fcIBJIKYZlvZO0Qf5GZ5dNxeMe90qCP/ayu3n3PBDIge1Rihuk9udLLoZTSacZgB
Bki2Qe7HgfG3XkPVi10KJTkeUB52zJUlkR0JUqFouW5pSQNEbbgbe6JbA+1R6HtR
N4FgSILuunc6r6tX6AWCdQCCMVp/92dE5CFJ3mbfFl0/xEfHRPEdiE2wATl8DzgE
KgPc8TjmjZIqmPk7jrMzD91wQsyO8JsLusXW5M5uQj1MFIcKxH/ylFZwnhrlkdiq
hMDIh7cmKg5Z9Ky5mpgfQcuFnZs6GJNwI139x69AqOryEbUgt/hllosK/rQJKivE
FSSGPPmxvMNbYk+IuVRBzuYYyv+Ep8pcP6JD9do9aSYZ4fBG8AHckmCR20DHqyBn
l/KB+LIewRaISGyjbEhhCT95NYePqfxQQp2QE+Kh2u3iRXdAEc/uLWCOVqwnXcc3
zydmFfRrHnQbYC9u3D7wH89GtpfEGe6rtiBzWFtYbaWPJH11ljeJmtV/7+wEDJVz
4x3/ZPy8C+5Vqgk3Y0KPtNpHXl9Cml0nBysAI5qWtTwDaPSBSt84jxYPLP/2Rw/7
HuwklZWw43GoBOFuhSdYNrCKukZfeJmO40H70FV58NuLAR4hF3gPlbPG3u2njOAj
q11sWoDymR2KhghpR7lOYx6KyIr1oR1p2Du2jgIcjBLmpvT1CEQoFNOfeGBVVUWO
yYcmKc/soAmJFfNSJr06q/O/TcM7PonNESfAwGVT5D+udvigA6qzZ7fP3ug5wQGO
+fJKy2KY8i1OolKbgBi9TLgMZErAAKsk2S5EYGWvvxTKkGVNvwnvTOHQpVO1cUMj
F3FosCHC9Ys9HRRk/OhW19rZggu100WRvDv0Xgm0PT7YpvpnjJOH1laJ5yUl5QJP
uUhF9Wg+XS0D6mjaaF8jaPk2+TGDgeAsbXJ18+gOTx82WWhpjW7hMj5qfluDg/OO
XSZnSkLKJeCtmLLmo+1M10Yi2aMiFpy4YfiTBR3bcoHk8Qp/k7WJPxyI8JCJCov1
Zzqd7JRyHhDKzjmWhGguIo2c0IF0BY8dxHzdX+D02IvhvsbgWed8ySrPG+387tdb
jopH8AdjFmNhuonuRKEyLC1Ar0UiXrV3+ohyLwGgRLM9IwfT1qNqGZrUReHef91K
nxHUwL9Z2VOs6mV1kbDVFsLNnih2NgNW5XavivCTwKZlTo26PHBUNTSoaG0eeP1u
H1tY4KVHyi0inuAl8hYuznaMTekkDDuzKTGrW4OnhZjeQ9bn2rLQkxSz7bRAnIGp
EE/ZpxtLuC6u4/8/RG870XHSfunhNDBxSg1ciKCCOAk1+TtRLq7CfTWqspxQ0e7y
1siqcUYJyBCoOFAniDWNAT9waLvyo3dOn7Xwz/xAq3XefEkWzQR8oVreLSv/swZx
3ORD5b5CGVzKdHG8a0T3u4wNEGzO976F/M4eVx16e4m6Jf5sCp8PiBcRYF4rLpgR
/H6ftK5+pr0SSAY8uMrhGBfm9/KihQ8zho0IvdowTo4E/dPvq/3b4W5w3lEZ24Lk
/+wHXxYTov9zHEQ1Ox0ZH9k0Jy2V0/egcwpTizY2SHaRd3ug52epyzmfmx6hkzaQ
Nh6QQPYrfSs9jZbtO5x/k979SgTYpLGXGRdD9cT+8oVrD/HOX4KLXy6Jq6Gjr1vs
MDI2IP4fm/Hd7/LmTFPtEiArJSaaF7dK0Wf0XGaSEWpY/cbGq6SxKp40acve8qWA
ifj/LyK7SWNx8voO/8ryq/fATtwVlkVNFsEMXcRMJmqcShS/LIqO2fZpGMcBaNk7
QO109IlzwkMfbJwKhSFXfRhjdW//cm13hSB+vz/G5daSRSGbAcxmkGGOCnXPO/ST
cUIl4ebfp8WDs8TizeUuoFENVVHQC1Rny4I+hvPsBheA444VEAkYIE+UeP8giJW1
JCaM8xmVd+bQtUg6cpY3Odx4W78eqVxhYpo66QlJtDwNFShI6bJUfIq7Jl+TqImk
wyHj9PY9b16M3Qw1Zilwe7RVDamg7s7xTW4OFnZJAJBez7kqcQkGNTpQ5NgATe3I
vWGcPco4p+ZUTddIr+FfF9NjoJflJNgvrt4CjHOyqp3ZhFn9QYPT2oP/MVJViAF3
/lAolamwZSuAf86/ovlIXoGyPgvCneTjYRXhdt1CuOv+WYloia6QdswCFmAOEhoZ
w69wpgotGeDv56KDdvoXs46VcX3/hrKHS8eP7jLB595oBB5bhqkliBGAonBhKgpO
3kzdSTmmaVU8q/WgrSIVejjAK1frmy2XJJrqEOJXTgkymfQeTBM39kWp3AjB1ddh
thpVoOVQKUTvPix5qRjXNqoeTrvwNeAM+HtmHhYDhmy0/i3YMlN+siQozU4p24j0
f/OcMkz84PrhLmYcLpqTbhngjA4MXEHZ5N0GVus7I+88ye3goR+3DTfEpSYUmp8d
2OWcHyz2UXZcHQuVj/aU+mt+S/qwO5MS5fTGuY17M8Rn7lUiqhR67G2ivzjnGc/s
S5sPdE0OKfi9S4fs/lnYH7063AusMmEyLdMcW7El9nXOYBwsjcd8Tsota8YiJ57G
f4IaT4cLqePRxp6JUD1OLtLXf7Spj6052LbmtmxFW5y1vc7OObYL0NI4mwYDCbXm
gX9kCGql8FjZH0V5LcYdGfZ3rm82tfb6ZMsMTcgUTqq2NPNSjueuCXE4aD5uGE6i
aHDzASCJ1U7HLY6aTsEv7YPTnpsVchg5dU4bJ9gQLPQfrg4dU0LDDzqXInxR79Xo
jgOzeRnas2Cx+dXD+OCAhSQ3LCjgkSvCymwKkmR1Z8X2OpEDW14T8//4YHaeyG3F
rwNURW/TIEaYGBn35CNd1WWT+shwyOUQZspvt/DnfNMIiuG/VviB8IqXCFG2vBjG
5ze7kyej/yFA//VgJWDv05VQPJN1HLrEL1fEEoece3G8/TA6WyS0BlAhkOugW1OH
mU+s/cq7BJSbrb+UsbtB6DDQISBvnUVOvjg4Sz4lSgf+8RvOYtXr5zYRmuHrNaKw
jZbRDYY3D3vgoWfzcs9ThD6ktUpDzdIygzFMBF0xw4wscriSUMcOYFOlcVkWi9PY
r7GkFPeuqzn2t66G/2Vh0undWmpghS9k1RgHvoVju6NhSs5M8L44cmA9FRAhurl4
FQp3uBqe4jeuClbWgwDTRFe36hy7/p2ICdE/7aX/28TKV0E7GHK75e85t9UQ2jKr
xi5Vi50K6LXR+48D8uj2A23LaJ99BHwqztgKntJTcLdctUV4DphhdRxAv8Pu6ixD
hw5umDuma0cmuP7vsnBS9oRDz3EXIkI0+XOvsp0VMw+VVnWXT2UcYpQp9rrpX32V
mYKvOrNOGwKwe4Pj/hGBVZ0WuuawWhLROCWpmgkcJ2PlWQ7zC24dblR6mexpJtYS
HGIM5GkTboyruswmGHIpzVUIV0HAVOt7K43naQV/0Uzg79eg9V1DLd7JXmTxuEPs
oU3FH318vRGgTvYFWGqWt+iSIXkqw5L3QePUCX+XCEZ5bJGlVwFxnCfhz+DckGcl
t94TKrhXE8PGUWWEx4fNzJQHqSv9QCm55zrIPLr2rzFvaKCXRCcyfEQe1U1isZrM
1SxR+rw7R4iK0Z9U8JgI0q1lNb4cN7o2wB1znJ0YQbJ8YBCcfOvE5cD/OZNd9O9V
QB1UEbhYB6aKA5lqoIEUwFnYcdhdx7E13tfn/E+mJno+P/+1ym72lykyfapUwMv1
XvKGurCVjLdmYb23wZ4h1fA9HBNXbVRqFtzg0zTXOkzQwzTf4XgxVeOhgxDfdGdB
VJn3fga2GDw2Zim0ZhGvocZLIfLdcZ2170pZ7DsloCZNrL3me1fgnUoBy0JVq7FH
pCI6Dpe2sohHGzCwzVHunXM/mn3HUzInyogls1GTTxU+MDncFbTqWA/K7yD+Uvox
uabyGsvxnZLUwoB3tWulPkWpmo826RHBJrM0AhDknaTwONBttlD3Na0se1g8u3E3
KGSbZJd5MAKfZPTnX9WYVjcOm+BzlU32pPbmCjwBD7x8dL04ZRB+8Jf4n+b4HQ70
3XjPks4/+zaWSLZ/2oF0p46BW/0HRMvc4wSRUJasIXhOsDRausSI44K6MXqVBBH9
ZqkPA09X1ceDoAVnF2BPg0kdObBFINnSbaWq/f9P+sXFo9yJW14I75mZZ9t+v04p
VPK1NTB1zC0/PVuYPgMWmIMORnpjVwLngqTzdnChOFHbQ3VVswdCvQRj52sXA9y2
wIAdeiWb2VnnU1rcgFqtIXdojwg6Hz9ra/JGEY/9bRg6FtpM8Us8LjgwJohX+/O3
j7MuB84luYiDmVGiYGl80YsR16WLiksf1KUvdUJZCwRRTZMmsr/KtBf/K6qjSyzm
036f4Y/xtglj/2vFTFQ9r9OLPJSjY/s8iEkl7yUjKwIyFPhR9oQHVemlWm2itCd3
EY3FCfVIUIcMu+MWPnGwkTEZqDJF/Isn8cSQS2VhtpQ9cXl4sRbuIgq/uODkt6IA
ofmk3eOUr+3m9y1arx0CxN/q8HDotx9aFUQ9kfg0pgt4DY11y8m8kQHDq4GnYycm
NbFuE0ioPDnV+fBkkwOOA2TJZieRgjpRqPHNKKkeu9dTDbTxscQPYKtx+P5XxG9y
A2x6T9tDk0bzdgVVncBAC960skNaAqxfnrFsUKwkavBbXsU1ZD9OyinOn3so9YYN
Qh11dHm04fhf7DPwDn+dwz+4xcC6kLwrCYXhbg3BzW6/5/1uVhTtPJE02f2PNQTX
BYMtmuooA8upoopMXMO/TygRrxMxa97eP5Ll6AJwMw13KqOjTewWlDCcvBxHbg0e
Grl9oLfxWReUQumEN1+XZcRHka4Z+2gdiGiFY3mDSvg/W7OTwivYnAKknh/e/2lW
LtzQapcpeAb2CpVE+rYZOwS9qUASTqWaf95kia+zMVTo7LuhVGf9wp+1NC8ziufJ
ITVVOxCqTvtpMRtFNV+ab8OaGwKXgAMk6L7s1UZw6VmQ6XqmWqZZuOQdHVZiHvp9
2yIGAj8cSILaTOXBhcxycM80IXpDIUeaQMjdpoMDf3rrttXiN7ABpHPSwQaQmGXZ
qpHuIDDnLmNvHrCf3aJLPYcLeVTSHSmu2IDm6gd0nt9HhkBM5QIIGGO6oWvAEZ5i
JEv9NjapbLcg5z91gWJWnHrBrbp6J7kayXAVOnb8rmZFDd7ofNrbYYQFQgF4EYPT
7IdLaajyKS/xmpHdMV5ilIsFd2lMtGxEU80MHj7TqRdqUdEadjgDIWjm0X0EIVcI
eZFzAc5pvJCeJ7tIHFzvocFQzFUt9kML76H0tCPFAX4Anet+3wmazs1QXHeUlhUN
68J9M+JLvvkbiZyTAQk2GPkBBb8VqUG+QGFJGH+LXfvz+0mEe8eM95kDEMoSCPjO
EtfLm+PJjap6I+7UJm3iepfbTT/vH/TwBi+rjuzJeibt8SqdqCIxHWxjVM21mcuC
Mkfug2BXsVZMrMv01kKw1x5p/BU5U9Vq5xsry+VFtH6+GdBEKjPz5+4R9n3g/tsv
+56G7D23SV0HRR1o85rMPnFcT5wlOkU8NoNOdycPrxad3g4iYWZCZs2XFcxWnvaQ
oakbIuGKARI5DCxWJ90WZcSGfb9gmBzG47AePKRjBathw14ev9Q3tIqsu8wlrkk+
OHeYqcxjWohSaGpSdLyN8WzFEnntTPBGJIddPWH++6surODjaD3tar5YHPfUqpI4
VxeOsL3CdBHygvmALgB/erFPkVLjR4wTSo6vWab5IuS4jhFNi5WSCruCV/mq1cfX
9O7TrqkM9JKm87OMRza2SpJY+TBUukDfNFSH9tLrTy/knKt8wIO49XViN3WU56WD
c1DBGpRMbWlm3cQcskXuY+g6I5u8HcLcTeF+FyUZUxGq2XRHTS3PbVr1hesnSVvk
1HjsLTiokh0X5bJcPAX3Nc57rjo4tybI4uIjrXR8sIJoOeJYS6YHWN+S/9U/X92Y
n3yo4V+i3dB6mI5XIkrlia4YMKiM3h3CTe32VEbkJFV9iOMUu8HsWmLdDPiBM6vm
iOlGL4X0Y01l0Y2t3D/C4syhQfRu7Ab9a3QCCMvi8jxfLzZZqBNwklYbJDPYlMZH
kCQE4vH+xPtrYSm37e0B7uGopEdmJRX9gm4askx6Y457GHy256oCrkqa2jEh9Zw5
nGtk5/vIwOLTMcmmRPBRrei3b1T7Eu4CcRXLp/GcISobWhQ34H2JAzDsBhHXc/IO
pKLTbtMdaTN+jY3VsprZBrjvaBXqF87pZd43iQKh5lIo6kz2JULYgWKsKStjefNL
YQMY4GC199doX887RM7CLL/musjET38K7HXPWilff5UISe6z7JX2ndcUof+sh8Hb
LEQPIs8mCrs6F6GH/k3ZOC3InLpdAyyXecnflJCZUiGQUz2SYsX+yhn/GnqRibJu
5YAT2FOZiBNZEsUfBMSNtyvggDiJBKbSQjur2Cp4Vh/8tPSzzrHJLOZsvIzWWdx9
uT+XecnxKsEPvtxhtBc08NGVxdTpZx9lWU3R2wosSmqqswoHiVSYVIz1wexbH5nX
laMMxA/XS0pLr1bc2n17xSJCzSg7eMGGCVarxiXoKMzfY6I8xX1LHVjVnXddlEQn
dkc1Zzh5BRKmF4F5ZVfOCVuNLytJ+3XJA7EwHwlNNsftMu3ZrZVLx8OrUZTVIdrp
dQ/Be4hFan+jLXCtlbXCFw+C/j332C++eURi7iAm2HFI7CCHYX+0vE6ZBRkzus1v
bs2u7/TO7KzusCj/reQUYmKUmp8s1Z9q785T2PRS/kwrfQfuannIfB2tDOXLQbmu
ICJropcM1aR3Vp+wg1YD5VEfKbGiiX2T/YxO0iHx6zqaKAcQO+a+dTrWVfYRyqN9
m9zav7yDzHkZLk1K+x+vG68qqa6vZbPCASUfQKtlLGO79frKvWuWVC1WGPE+Gm5l
50hZcOIrTSKSuXV5IAN6JB9LrqpYtHHshNRqxkK2otUmw4TRrDKYHLm++YQCmZjB
g/DnY7p88nq+6RjkSK7QyiljqYiNTN5ttubz95KqjWgKZKz/D+NE+3bCbksgu4SA
hJuHU2s00u3cbypFERetMJklj5+U3itZI7QjV0lqZ1CfNNfkecWXv+Aoa+LlOkck
biw1xg7DvQPY0Hfj/62Cs3mh6bdvrsbvoKsqwDgWyQhgScCj/xXZVYL5V0R+wyUG
J2GF5r9ZituSUPj5ikxNqfOzaZ9wZ97C0dgidYKoLgCJcQL9Q3CT1m7ZnzxEgzsA
/0ZB3m24VWhuDfDil6OTh6lyFHTUSVNoMcGwOQgtRkPzlZ3EA7D57CVwXeUa6POi
gB+/yzc5FURZueZ5T7PwotOPID9Yye6jF+0vqB+Rcb4mNUYDzPSVs16y4ck76j4a
Ve5bfs0oxEdkYEvUUfq3L8mMwSy8VNkPAdcLAx4T/lQvZVQFUnY9o6QisCb5bcfT
+J+riADg01TyzN1ko+w9oF3VM1ciPmOv/3RlUBxmPfOPAez8aTbHr7G63q7bc3hS
ztjKWK3jBlAzi0gzkev8Th8cg/sB1rsRjAL0SFFpK/1JQORAsn5cH6RZjXUCLXW5
xF47of05dR7aXqECiQ9uSzTbD+A/GWHcMsSQtyzNeQ6fAVa8fTopdXFoGu+hUSW6
3rs0005PCDqrJ4Ej+0/KO+oQybpgqeE8KsnhL0Jd5cilMITJRzVlwke9LrSULtQR
nc0Pt25seMMXjIrJcuwvySRmpBPsvqu8DWjDwnmT0PNGDAXx9QnNGNgzNVplVKmQ
2erK//SPMiB4x/Ew+0nPoTjIy/xnAsYF3ZvQfEGcx2nYA64ukAvX6UfOzOZ8pDXb
U1ifbw6ekgp1P6uCiKl9gTjFf4IR/aqZinOJbGGN7yrUN9NhC4gl3XaNlSFAr1Bq
wpAwvgNrTjKepN/Jfr8t02KjBUpKbHDkPUoUaLei2yhALswZixEeZiMSh7QIzYHB
ogQXRDVvLsX8a9/nlzH2M3+LRpj/KnM38M6Tu95cym3Yg5izkmVu4UQ5Ge3bbCVC
dymal3iGTkgaSzCAuwzYwVh43EeT4BI7UbIoNlbDLD/pMVuhmgozTwEgOW2ANHiA
MyPDrmo6m1vzZYrOyEzSugYLDX5/UgyzfvR6d9dsbibyG4htOx1q02/EKMuPWCCb
3KtaXXGAKFixafxUanMmc85csVDDKfFGxgCwr4gEWQbLgmDmkVpTYcXXRXSo9Etr
lLw00YSQG29baT3Rk1N2yjU2Xtde1nypEs/GvKFkNrUYW7jCchP3+CBArND+ftKF
w++ADffbqUL58Kaefwt40/pgt0U7o710nwxeNBwg7/waO8qwvw9BoKavcUz1zIBJ
5K216ND6ZHhjS0Wg2YTYCyiB8y24bhmJ+oPl5LaoGLy6W3E67OSQ1QJQ/ni2Fsel
4MDi9wzY+HYP1NeiW9ZYwk4sRJXSAeHCq2sCl7e15TkAMxG65c8e2uri7C+eA8SE
DN4hToTDAVFm94zN1iP+r6B8oK52x+0hWSkiiwzFmMSiDuzl3Hcm+mp7IWRpnCY6
7G0Kje0GCQwwkrYS9LVwJXSvNFM6wrhGtNAnixNHFI6PLwphlmSAb6K2/+r1gSFy
yi8OTiJCUBw1OJ6/03hXPM6hBLRcs8bHNBB+WUYH7cgmOOlZ8e9XRxPr3xvnoHIi
pYu2hYAG0K2h2ru9nzyDkV33ArMejhvKzCanO8ZxapeoYPnPtGUWoY5NX9EVqg79
mTKrepgip0XHQLD2ocgwvp82gkG96OEILLdgO31ZTbmPas+r20h9aWAAjVbxk/fI
CJ2ki8nEYHVyM5PIXI414eNDAE6zTRIiQdAC2QkxMakzmyNkaUarlVMAFccqwMu1
gd3ZlCNdkSDoA0oIbWlpU2N6EGDUvut5OwE5JSs8WWRsHnIyZffgtkWvmkl6GYAh
Pi1oganIToZ8bruK05FJ3xGLHe8nNTQsm3+SvlQnrbnV4aei2B+a54lqbtlkQmGP
nuA8N7FWcWIj+tbFLZDkibq67JhymTI9L97ikRu8j04saGI7blLN4rIYJJMr1ZKL
YziaXcZF0a5oFP4GMKm4BVIUuh7rCJXIYE6ei93+dr3zrp6YsXBWJ4B87cbHlyYy
idMgTRkloLdJcScTtVWvvYlI8L8eWcby/O0Y6LhDtuZhfTGAu444NynhlHwuFHGk
QS7uMYN12A9rTWx0Ai+Mw4Tk9VKAtwXXDXPyD8AOBC12Gl85wm0sZyQ0f+mm+sEJ
O0mvA/c53RcOP6zeStMTeCF7iE3Ktc5W36TZyyWsju2iIgK0yUJLiZCjxtucVZVP
PeRVYIO7vccXpaWENREfrzDNMrBVKJDrwHqymdv5PpaGcog7sVzQ/q1ii1J1UZPF
AZi3uafRHzEZp96aE7r4zEHqQRq0wmpi7bbGVicoBPwqxBt4VMhVjon0SqchCST6
B6NreHdSEKqrURWHikSHlya/uRh4zX4+0lb9Xaw6akBAM7CIa5Oa15Yd9Ua6N2lm
KG2BMX+Xt+wgcS3YXo4rqj4Q4yR1xFVfBUBBgJctmEOPSZMZsuGxhajh/BVb4GEF
ZnMuBMlVn+eIRVYTA5fdjdG4rT6SLv1Pnjfjin01ZHPOqAfLPnqulrjEP9VMjjCx
RFD83U5v1+pa4ZP/vdYI34qtec9fsuAQPMffMDfzdvx+2XUsLzKu1r5zEaJSDtEI
2n+SJFRG0/CN1ZoB32JOMkQUmfjIPyjXVvHF0VIqt98LAmKKaqW3Ng8f1EzyPLeK
82sU7HJascLFa9Y2+aNJ79HH2zS1b3hlBh0DcwS85WM9MzNAkQKDGBcJpagzgpPU
FfdbCRFXB8RCETNPcIxuLvgtoVO+B1fGFfspD4S6q4nKIGQ44L74hVJwCmI4jy7T
f9W0fAvNwNzhKvnl4zlLOXd8ChGT2shYWYzonmUkg7JV24dO0IX0EZPhFPrGtta6
xPQ6wHcOxp540NwVWfN2gwljPP2n68j3uYet3sP/u5c1krxuex6LSfaAGU8dAUWZ
DphfPt7CRKs+Z9Frsf+Zazyip17BPi4oUH6PdIR1gUEguzQQZvNpV7flnSIcNY+I
Wng0Nge/ddDnaarfTKj+nh+oYnkmAzuiwxW4i5oKHJHg1j5TwXqflRRHV7ySGaux
ZAa14MwAXk3Q4u9hQnEaqfpXZI1uaLbZPMI6vIGwpAz0ceqfZuftds+WGrSdBuel
OVQ/1yaWsg4CKmNYihYcLOyLSnW+BuiKupSKwBhsb6S9mpTFER4+Qb0w0hld3Hvq
JFXX7ztmmrb+dn1Nf9MscyfDcYNRKAzHCPPCKyhCx+aK/br3HgHNb6A2H9VkE3Ap
n1C94CYA7QKocM8wECKVLjwJRBGuyqjtId2Hw8M/wH9LZoEPmPjxW/5pgEQVpJnV
PbUid9sK9FnrgzKot2pzBtVfZta8+/JlUTDrBaxDncwYEhZ0e5R9Rj+YHWTludwg
MaOYfRDtF8j0dK3g0owntgqPrW5m54IZ7V9X3A0uigb0Z+q+7g6/Q+e6V15psdlk
XMDNGre8Le1owDJD5Ja+7r7Xw3XrMdNRte2jKaZ3pgCbu5lTctZDsYziU8uyi3bo
rymOCGbGzQON4Rcn1R12QQkWQxCAXUKLDBdaRJMpcE4urZai8noJCM/ke+arDbFA
NJM6gp79faxYrXvG2uV9Klzamqycl0vu0AxfRKKvWl/wsN5Hn+aV7Q6JIsyo3nCj
t13Qg3ilG/5I8zf5hvSI1EuMyjtwA0CRkBsBOkYGCl7gqJBXwkJNpS5Cpz7lbtWp
KvFqEXsOwuNSX9QnI/GTtX4RaAS8fSSBZd2C7L5I8x/SEPseoBEJ2pj8wiY7pW1C
pwJleGbHdRlK8WRIsnqjo8y5tksKgjgC7cyMlix+9eVZaCP1n6aMkWcG2C9ITM6X
DbhG4nF4f/o5eH0k4eie4t6NbvNdNG0WeftXhGjgo68tfG6zDemXTXNXqnhS6s3C
gAcJgWaXDTHcHCQIxrPX6HLMcOI6kj6E4vOO+HVVjSsx9Nk7JQpowJqmtPrcpJ0z
/2xLnEx+5cyLEIsbWopO9lB+1iC4J+yWjkChdivGoqLRnUcFIQLIV+AfvEg35PH3
rff1zKZCbH7LuWfBcjfPeggcqYvVWjyV1JSfy3nMjjhEGPD72cKJWVrbO1r686tt
9S45AUsgIA395uFpC2wYSqmpqxkx1nthxWnhU805W2FhbK9R+L3hP+H0psNmidQL
5HTadFGfPE+moCrX3FlBm8ToQbaJXtXnoluqM0XQ8p0dLx/zB55WvZREGJvavKi4
IKLc+WZ7OHHgp1ZRNGBWsifL5Bynpm5PwWIXgtBmiPfbcc84fVZHqEP5sONiGy5J
XktYMvDh4xTAvvJkC+5k5ar82Ly2FhQIwwEzAW7yXOBnxizN0HzrzQP7O3y+cp9t
2Wl6FNFn+HhwME2FRPIB/ChnwDEZ/fPH7xPZwHhAOnYfxck1apPGIQNQmXXcJUdQ
jnuCTm5beA3rDwzxD7HyB/P4I9GLR1/8+vlauQ+k7tLWtK6376XT8L8E5hHHBVyp
+AxdzZaSksDnWyHNL2FT+qTNWrIVzMbXEcILvluAozV95wj+kpSrI+ctOlnQsHRN
fYzW1IwsTPP8SFp/jf7MoWGpxib6S+FIW19JksciXTgZnxrAPDZMwpzTNauOED2U
cqLiDBfM17fuVPOiJWfnXBVNRRlMGS9Enl3zH2TBkk1oMjndpLuJvF/w8vOBSJlY
xWse+M7mUol1FtTZSsfPlTpi0TDhZDTAPlApDb/Mr+tPycCnGU4Z0i6yr16Im+nl
Md+frUYW47uxgDM3j7kc6VK33dANd7gB3xfAzCBkTa110UP39sw44btP0WsfxLnk
r5ACowvImex0VnkEQKprpKUz65m/jaMf/O52srszHCCwp7tv1vxDV44WubuQ7G+P
bhoF8MRZQ10kb1AEqsxGTVVMyVXPraCkXw1jNBeZeT3DmJIh2bMWrAV1/KU4wy3x
srIxxgcMH67LOvwfEuk+Wcw2CfOZV5L4sku6nxaz2uHxv9AC7q/9niYXLZ1VnURz
C2SeC6eN5k82YXojVEtQDh1pmGHe6JsY7z98AvDdbBCksiSvXTbN+jgdDAh9KJFO
geugFM4WiGtXfRN+RA1IH40Hso6e35uiJHlHglt2hgPGdanjluJ8SCtvV29frEqx
3mwdzcCum4ZhyN0N7vj4dKYxSnSNPTmOh+rVV4E3InUd/KAIzm425WdtE79gGmP2
lq41Li4iYgnJJwu6QilLSIiRKQgLL0JH1V3UKkDxNQLAy4o+9SyEF0Dn6jFaTelP
Wc6BnZZthUZO0OYNrjN02Za1DeAlHhV6lyDSUSrBaugg2beq9A4FJOQbzA1gn3Pj
icJPxy/Vu3BIdn2h34mDm6Yyp0a98sf//SDeMGCVmjqlDX4tAD1IjAN0wAi3s+u2
Tgp2WY65KKqkb1aZkWCsCHBuK8+22V1v8ZHUgGfsBFthc8c/lR8IPZeIuCx9JAUk
muZ6WS5cURrp31VLPYEywQ46+YCUwKTCgUEktPfGMPU4V0siH1SpJ56rM1M/EQjl
HvVIT34lX/At4/YomZ/k5TU2YPBeUON7ai1MMhePaZ4VpiQF/0lcsiuIbMf9qwWZ
nyQUddTwYF6DATx/qQQayN1w8cdcWHGgMkotFGVRUMPFqJCkxwaHYHQCJtL0Yjp0
4n+eMRWDoffOiig0RdcdeYm5Fygdpz9g8tRpzxrjEdY5/ivEkAzmlaq7TQQ32J22
SdFvxg/b0JzDmP1ykw0BkAEhcTSOiNiWBpba64X+MWhSw8gSgRwrkxj2vmSeIcMc
PeknM60XkmQ/59HKwWfGj+BkZtZcFkSnKD4wmnQjspnA2ChqvkKjMlwVhu8Qz1tU
g0iiUaVn/jVdz2CgVZYWH1CfJARQ4jTekUvlf9lAhBVZP4QNS6Q7I43PaGRHbgIs
XFNaKJlU5sB8KMAR817Cc0v+tw+IZGRYRSo+jMg6I7yWRdH8IapGwTqmyuW3Fe6t
3wybvmeX+PSd7+7hL0jxtBA5E9E0U5yE+wpvpp+HkOM+B/qw6wQveUD79AMN9rZV
X/AsCKdruDeJYPbylqMKN27mf2VNumUj8936mwfhwhX23KwbYv9+ogq7bYuTprtX
MbDTzQGGFh2hsmfb3yTOFjUPvkPBQPVnnA1LjOoveA3bMao7F32azfeSQIrcwjTe
4SLBu2QWtR7jblLbabd53dU7RPOC6uMePQjQyog/spelB/un/rYWfuHH1YP6MDUN
9Vc2cQlGbOK99ZwrEYeJ4MmfcedulM7qOyXlmusytZtGR9znrBUdKS/nkrA3i5RN
ic+HtpTyS0HbjrknMT0G5Yx+Nv3oAP2O14N6Vh9LOsGXfdftyuXMqCwGazeClD22
u8E04irW51pDgLBurJEAOcl2yzOfZAHe5WfW0zUOmA8y2ZN3QPw0kCAs7ExtBRxK
P/ss2LS/xNMcJSBTNPkvWLyUxSJ9Euv0SXJ4uW2lIQTEyGy0hEULQ5qxB4BXILSZ
b4TlHsgkGkTd4fwRw6abxoht6TNOB/X4+7V3Dm6Qb9FiCHs7lsKsrEyrbv7LRbcz
9s6ZjnMs1X5ZtsdbsYCTQ2GMsu1ttEarwg/89urUEWqML6tDCUDg+0d5fx3O2bHb
CFdczUoUH5m+3pwiyS06yshaFoyIBtm446ElVp/qb546VMXef+pR3t5h/446FtSw
moir9hnvP88JEmvTqTVMWEuKUBDxjwlmi3h5ahKlqMur6nrbMCP6mpTzKPB9deEI
z5RVO322n0jbdn0KRmEnM4vRcsxEner8zNfypvlRo1NhOm8yVPXOs4zvL5ZErfdE
jzOkpb6S+aa3buVkB4hoJVNbNN71KhwcnpORQFTOm/6BUrjNbely/E2j955lzPnE
uPUbPQLEzyD7KCMhDsmCasxVxWQasf/zZZpdOILKPhC/jEkoeESra5G+4wZYnXbI
SKElhpl6iyD495ecUIxY5/DHocDlNHyDPupxYl0vmolXp8H0ZA3ixQy5gNRakxYO
hcxv9G5WOrHZS9PvLyfJhLhNBXp8MGAfAkctSVW8ETck1ibFz/OklYcmZflpFDVs
vRLvhMh8F/DnkF9fpXwFCOP6K/l4SZ48syoC6tqiCfLyo/ZSHteyFulPnASVVtJu
eCtPWyFHLNHyQYsD5UTDh75uNYWpdtmSMvzm57sTfDlsEM7+nVQgL1yWNzhaLO5K
TqBgDPqeUnNsDEbhGtXKJ+8We4MvMzfMVm15qPVodRCzSInI48fCLZEQaiGCzkhw
O6/o9C/usXRmi+kEv9k0qpHOHn4wZA9VZpIDw3UjzGPJbv8+HguVMIHZKON+4Jyh
61lImw79OfnPFgCNgcygaydK5NnabxAJkYwUIZpTd8j/g7ai4QCV4GkReKUgOasq
K2lP/oMKm3HTcgKxMObznmMEBqyIU6PdUXTxDPJK9Jcz6rjN0eCd+SFhfEGNdBsJ
aHVapsIyMdenW5AlxDUSeFsMSFRH1oC6qc7TJbhXeC1Eo0AJULmwSI9Nylvkigpm
Bu1Af/qIG7SdpOrpjSF7LTXonsizwhvnMINHWqjjvJ6zR2ezJwvXJE41HFCvZXA0
mIJ7YeR4XLEy1v5FHbE7xxrMkGnpM2idUMV1y0uInaf2ozD5Mi/qgvr9wgtANtdd
MF5LtV/J7MUy6r42DdVyRghasYSlCWagtu2/r1X16mtmEAPurQ6+TO3bRhTadKG0
XtrK4ArDX3mMHlkeGMpH5XH6ZzZhukJrDCk5XX2DNUD6Dlm46Uu6uNRD0wwL3GWD
JYH8tnVnNBhk/6J7x/v0DzpKVdNKdnaPtFVToo9NGXm9TvbyK2aL+m88kb160CVM
XGWdv7oX8U7kHEy3AUTe7uAWh5xNhkkjxFwfArMCE1WbC4ob78rrcWp9LX/SMGo8
LrLrJt3EHL5uoQL//5VabkRvAyIEliGCvstQXVSF3qQCQafGpLJn+YNhcXMMKAas
4RrvUdV0PlGBsyur5uIEQqojbXSheFHTysho71omaIRR/KjDBlzDI76DuB2dFoWt
QvmVdNr1Dhnp8Wg6dkA2tLUJyAmBbXh6dYUWOp34tacvb11UrHgaMXRkFPUYzX6V
SyIGwqoS2P6o7aEQtC+evke460rjGc0qUswdqSIA2PoD8O4E8TxcjKxKm1r/FcC7
gReNX0u7ZGq820vY0Kr+222Jb6hmmJxQBHqpTP8Bc6n9ktEmNdliNaSIJtXPF+/B
FPlhIXzbtS63zcvT3qb8baZyOJ7GnKtXR/3c2jLhr2MKXSqeO40YmPCiWWJbdneb
ykvNTGjtqXCPU9mEZ+Eyq4DmWBtW+tQiP10EwVCW5M4nwhf8i7SNKXdJeO7UA++2
xxryu3KGBeXDhoWq67tMbLNsYZ4NCg3Xtr0LI86Hn3EuuhUEBilquOuU/E/QuTdr
wQsT6i7n94dYD+0YbJph5e4FR78iCOOfIQSmNWifJ5jVcqJbcUs3mH1JnenNKcgi
f7ywhQzPRTAWoqk3kQ4MzO/a7F60/FoUbsuyO2wJXvVbVPZrCG2AsLopQvbktuYt
7ETmOoWeQCVqmRfVBXI2IvOyfFqD23/KAmcq3+8UEs7sZxN3piHQpksU8FeddEZm
8Q/jYTut4VUZpg+w5x957NLfXvupC3m71oZQiTl1FrWNH+HR9WFTnSLEyTEtxalo
VOMCYfNqOn/cOwkBMooQMzGRTfUdr06D+aEdo7IhSC5wd9nY1F+dSa4qlHXzhrqC
dzSxp6cTJ1ulYZGEaEDLcn+0rYS+QOVwLq8h6bnyvW4eqjNwIi5V1FeShFy9VJD1
ozybx4z/P7gz5gJrvCP/5+0gy8F7pGPDZehTPZFs4DZLhvdgFle0twqKI4xGjuQ6
fth62mtN0rmtpTpivRwRkYhUISbRm1FlvM0+JYbIUswQivBwP5Su+gc04/esxEUB
h20cVu4ezZHnT6mdHa1EHG7w9tW2ZoiCJM18SfRWqMyWlCdw0bBEiAdFx0P3Us/R
pkIWiajmSq0L6UgegGp1YkyJ8WWLCT8CcRGtFFQ8OHeBLGhlZpnxdutfLIgDc+jt
wxcGMKIz78m3+WsTV2aTuInAoJhln0qSycLyRS3Gj9p4moJJZKtJ+MxsjkGDkEa9
ueGWkxcCFJ7KkipDEj1LfDbahwE2EbEVaOtats9HJAHCvSl+T3/m2PORbACSVd7Y
jtEkqZTKYIrkx51oXnNzqeeR0kZtOYTB0Zx+Um57WPuLao+Lp4rabiXCStk0LB10
3eM70Nj/M6gkwNVQfRBUfG7cq3njTR2bRvo72YtUK9b1W/R8d+k+JAaxxyy8ykxc
UsQnL8zt6Wc/AS1+dl3F8O2VInu4O7heuMj80AcQGr6aV2V1EgFiYCPyhzNUdU1f
9AO+LE5Mln7HI/bvHCCR7hwQDtVP8bK6g50ezFmODcedJmgZ6eGswdkUm1GVZAls
stix/taIQ6NrP/3QXsVOL7Cb93zYjm+FL+UfCIM7w9mBcdq4GM20GlK9UUY/mOHA
kNk0Tn5qTNXgOCea2TGy3w/TOwQq4CXfNmPVMQwv6jfFFSgPf+BBku9v1HRZIMXS
neccr+SJ1kcH+mf4bNGHEu77bGG05Q7APe4Go6c9XQUe67BS9V5+KBFQbIVbkUuN
1iY87kMloJew5Gkq9Z5REX7EUsWHmHyBET4x52xQ0zJNbUG8UrBiVRNT7bZovrdM
5KTl2oq+699PRyFaRJIDnmQfmb9yJJcxhIsgTdaBWMR8dVIVUn4Z0mIRZaMu6RAe
6cFV6f3eWI+i6x62LzxgRWo9hDsGNUEsgk1AfCGmvQ8FQmSxvXkjQkhF73rmqNzZ
/CwZ5LdS7LU5/yRtgmJNIIRgxol0BLeltMY2zgcmWEzB9q7yd3oFSoY70myTfgis
3PHM0sblLWBIh9zPXjLQcJ0znyeX65MWKnbPF7zxMF+MvFYelxqVYgE4727UEUPN
u6xTnXtj81eYve8v6Vq6aEGckV8OxW47TPUcmVWqfVYTOrg46brHVLvc3eSm0HJ0
mn4x78DUthvSGE+pdvMtXhRIeAxBsQ5NaXNmXUGZuIOL/VF5U50117fNcRa5+j6V
B/M26j4WJGI0//7Ri9KlzJQqhjZ3ALIWFdCuVOnEJTARGcMPgj9/T282P59GStNf
OjNoTr/0bFwEjA/kqiqJF8+oDDouIc4VydhUpXG0hAWXn7c6GbM5J3Wmjmit9TTo
eno/ahHifDBNn2/AtmU1ANsZhvTVOjI0ZP+67iQVZLTKuACMlFgXvDMZc9VeJGKW
Mql/Nk+FoPJ2kegPjkL5Omtv7SxDF0/D2zYs4JZaRHKd/rBELksEdHwzxmO0rIC2
YZAfPxI35VuCKQuVFTSR8b87tCvD8woTBr9ZLhHsEkI+2lioEYhYVvOgSMB2wSWf
YWoEBdwUO/Dcl7vXp2zkX0COxcTOGYxCL5WvhER+2TNzj9XH3HuvR25Zp70uED/k
gCIUx11oGX6QqjXdQEJuUQCsVIFrVH9BxzNEVvarnagI7ptA4heDk2zWKVAQdXqX
qF964UL3ImQkW4pXY/dQT9TdWD8wgQAnlQEjz5MXzqa5zCR5KxSxPJ3vnQjYlO1H
qqQzumiM3YhTUjnfURmVflAfBIq8MCdQDyhfsqj/kmt3/1pZkK+JiZT2TvUBUAO5
wggZOpTMIsNoL8xjhnTZiLs4MS6r8IIZRrgj8I0kjPDAZYO5MGyz6sRfvKb8lBuH
uqUZpU/DDVK9iawWcGQLIYNErMiVToTSTGKTGtTdEJ2lgsnM34/bQmFDUE7xNreH
YY/ounPulVV33+p1tT8HpHtfMuocYJD17U1h7tYiLacD5fYiAgvToGvw4o8VYxaS
6ReAB8s9PhMMi88nAT03Hxe57ExxTJym/t1SPGmPaE0BRuPqBl+e9wyfPSJBnYvN
/FWzdB6H1QyWBI8CD3FKXv6nfSdqx3zSQJx1ruc0WYbwYk+E1U6ANWoaIGKtCfSC
m3QjH7C1dsrxvFel2NOoV2ZhJsrv3x39kETx4j1VDJ9SrYtWnFQw/ZyTJ8j1RBMr
GUZf4H6rAZcuGjR8MCZVzDf/0g+GUoxr4+PBpkjUsun6iy+Q5VjN0yPVjXVrLBJ2
f5SnxEWY796TAJLzLkxHAMxjLOycIkFHyXfQsBH6pG9BnJbpW1NPZ04OgeoXoUxU
DDiYR5t+XpEobbag0DO7VzLmt78N1+9A39JSFEtuq9v4980lnNk3FPisyT1deQae
sS0YhKYzXI4QEJ5kBLM3+8ggmUowa0yDkgEAzLLdW1sWchAp0y0cme0D1srUaAU7
bHJzCOPVqm53X28/MtCwa2KY2DQBU4AguGuVl5f6KnOF77V5z8SvxIo5gbM5aCHQ
a4dak3P0ft0HLIMuXVRuAPSrWLfxSdDeeBG7LNgSn0IYYSNdg1NRkG1t1AIHqy8M
oeTk5cwYwAnHCsYYkANkJUIIzn45ZcB8t9v36FK4yOmJ3RUisEemyBfWURf2lIaj
xwb6SbDtou0RwiB+laIf8pWBlGYaxlA47xgXc5UX/Cd1NWzP1qYn37RoouKON/SA
r6HjXLjS+KI2Kd/juDfneoCzIU+9ieewP3OkmcdGSsBES4vaUIGY9n+cKILONXHX
XlYnStiPh7XooyiUQYZvpNMjfi4Poz0fHD2/2gnCfLAyPXobiWf7GEAtd2ORzNqQ
sX2HDgiuGKCb/fbbB1qNIWqQ5CI08LBHdmRGaBs0bgnXxP8YgdDWwCeYoGvPSgKD
aqCy9X4+jVDRpIbTpq9NMKTxL3Zrtah+pp98MtvOEmz3jurAH9zbO95+1wNR+tXH
8PWfDMkZYX55YQDCdQPfwBCCCUAZeheuC7YdO2csUr3Ieq6JzObNthfzWsWrygCM
2YcSSCqBlE8yLZ73V4PQQqSdAWvBMUr0JXBoTGo45LIM1ATS/cWesxnaeTItw15B
hVS9Uv2apqVkhyUiyETsgge7hHje72YHJZoQqqA3/cLwQEk29I6ducb5ll41HiIV
bmmWYwAFHVBcHKBuhlauBSIwHWshI2qs3V9bb056+8FFW3Ejad9700vercMeFQJk
nJkeW6roA7NtWTw4A+jOD2l3biLDKkm308GjFbwJ4L6cKeoBIvB1BdTtYKVrwPsT
Tlg8ZYSrS11YgQfHzeH63kJHO9z5D0/5YhPNZrcUKh+NVMqwz3Jzkmtsd2GIaUUO
uoV4sdq5MMe3J5cB4Y37gfItxElDsG3OX3ofJ9bZ9D1bpZpe6lgUpyWh5i+J/Lby
FT4nNvAJ9DB/KTnuWn4XZXH3Zh75CXyZMAXzuVnrWNWF12Yf/PlT7V9Tb5WdrYbY
TbAa5kbc03QBtWdo/Ux8Hy4AGPFTEKi4AFVbP4ew6x83tFNaFrQPwzu47Bvqsea7
6qR3dxzxMGHnBAue8jK95oYNEioLZNVlxPNFkMYCZH9o8dx2Y0SkOgKFgCWU1EPt
uACgsGnV4D6kpGc1I6xyg5GSHQ5UoSdrwXvAy0KU9ZHlCwQCC2/w1AS99LaUKbLJ
l4wXYqcqpPnuZAWqe07gXG6G3Mbl/4CBnP+bBMB8gaiibxwa0GUliQvoHooJKlPn
keS04C5aQJL8t/3whp9pD6to27LZrkO++0pWmgajKCnHuGJfrRB0r+CWDiLf/Cjo
VdNGsJKrDA2jEaeaDpD7nOxSFfcu7vbhooZQxI2s/SSy2w/aDa8oEluqd34JW/KH
f7PTeNypWMoDBlO7EUDI+GPpmWAwMQ+hdqPz8J3FKdmmL9Y1gJJuYZ7SpMj2JJTU
RDf4U/RdmurU97gsbTXcgiEzJuf9quHnfYgvRIO//XiIBqexsgqF3SWcw6aJFNA4
c7ucrTtNsfqsk3FQsf5BJQRjD+BviFdJrvx0mh1NOxUpRj9SdtU1pUQlhdffasgd
ZCLL6FYogBdmEbXf87OgOuqAVkppURyyCAGMwONKt6DJv/z/bSBzcFs2q9KaUmcM
8HWQINUd8a9f7rlk/f0Sd3p+1G7myGfVf8dGf/Jaz/MEDcxUAoQDT0+r7L7E7zud
nO1wOtKUFsX7xR8vlyxwlGa4lnK2Hnqz59LvS2weZnB5SNZ2sy3U66luP/HDgt2m
mx2DHTFGOF3xiTDJKlihO2GeukEbNeGLHjSjrtoOdA8IFGfe/VUpIcDkZwjWcoBa
0f0JLXrVZdHug5BbQQzBt4kTk6S9pr+jq2AdE+Pwb+kV1pnkYPZfSZwhQCy6KdX9
5sywkHDfYo+vkCOjwvZhWvsZQ/RYmUweYunKmKJqo3xxnf/9HR6uf5j5Vz6kvkrT
fkzVRufyeko6VXnCmRqeh4YnElkfhCs99lr0Akc6+FevhRcwF1WRYJhLM5tq3XPO
Z6FXqJNELbLn0937HK2xAD64N2nCzViVhDvx7EXvknGRgJu6NwWwlaOyTWSgB/DB
tAUeIq+519cpJfBmMwE4Je8zSIdNICOOvm4CykvMue6bzgMPRXC929RG+EnDBWB3
bbHTGWX2QuO54CSEPqJhzwlX6AmyxEA+qDr5jMu20MC6gFDfuMJ+19pn37zd2kQk
K+70lAZ7CqYTGGeQuxaanWGZ9+n3TOb8PIRrvWxsSHy+DrkBf4wkLG3VNQ5D4XGD
+ZD8eb+f8fzwbNfNnfPo3OClXfqq9jAvHvc9fPA41/23OQE7sZYpDuwGvfnwPyQX
SUj2CIUL585HtpjpuQkGM85dZhhcd8auOaqXjM6Y/ifodjc6f8wmx2faNSFy+WYn
z1QyXT4xswC4M8U+KHuYbFOhM8uVtsezT5HWHOmAeyd0n/F7o1mRV5onKlJp8CRo
X8NkqcMeF1/STL42olAP1f+GPNZXM8edJrzXja67GlnO5gozjSi0yoyDmr8Ap2nM
theRnnoluqXQ/tYrYY5F7HOkDe0P7d1RcjN++y+urHo3pGcKCrm5Kx/ygw8xoffj
CQ3B3tc5BspUv3BlYLGQxgQhHeOqG0w9pRnMnKUcGDrK4fYKNwkeYlgjLfuODAd4
wqlMIrVuot5ehvqCzozr9Q3/ZaGy/GQcspE1XObhpNQgpmQvjflSB56F4I2W6nN/
C3gKCxwg9r0nAOhMZLwC1AVnRvcvTOrkx/q7vjXMrNk5UfoMgmVdMNOScG8MA8q1
PkT53LVTRp8vxduXZvyD5kpMW4DdKKqQu2V/4JMewid/GPIIhCPIgV25dU+Hnf9E
MlKHmtrTPC+zedhQBNxVtT814F1UpEGPP7is9+YvSHz3tbhypEkwNVSYQeAjc6oB
ybCj4IQMju6KtexFk1MoE9KvEH/p/S5ooUk/bBfQ9Zhg+Dbf7Tjgte1TIFr8Hr4l
CXONZHUBfJ9+w2lXcc6WqBmZbJdXMgBSrFP5Ad+XFXhRJDv4r4m1TpqirIuKevU6
y16RwhyI8dnIamntSgv50mOYLAYUXiyOd6Pm44J1FxpIFvZQ1ohkqW4GbO7oSsxy
wSJAIjw71Oz6uTTnm6UNwMGU2pXKfXu4jT2uruvXYsEJ2rzHE29nPhdgPTRMHqSt
HLN7GIM8Zg8IwTpn4snivrzYMshq+l2ut4prfAQgAsi+KwMTY569Al2GF9kAXSeA
k3Qam13Xqihml0AdunY1Jjxp42AjKx7KnLrOuVRRgHXCJ6z1trZBzFqIOLJdeq+d
pnLFHAmhppM36lvbHjwfFD7zyWRlles8TBaJmJAXcnzG8Bk+C31nyhKfO6GBsqYq
chQGg7vAA76x0Wrnge3cKi6yZaWmVmLkCcqlYTKqLnl1qid3BNOR5+7Z805gst4x
wGiMGaHYk5QJQKQYktC4HRIvCQ3UPHzf9orh4nJQ9a7x13IHTei/3oqSFGouqul2
hbr4D9eJni7xoP7f7/yqjPR2Diu/ieTEk/0NBrooaBriLkSAkNPItm4rIsclJ3EH
glZFguEeKJPLdKmMCha2ACKzJKlF35/BIF7x8j9HKu2O8qvowda2fBbAd+SnGD4F
zBtOdWc5NuvOGyIUgKWTezqU541O5sS92Vj/maU0g3ET3JIIAeSmP2Y38oMbkzgy
xUIBz+NhlP4XfCyFNgM0RKNnH7Vw8zsAzJ+8+3W1+dwTDf3KsL7OtnEc/egWeiA0
77jJrnR6DvyxvMcyt5R9uHettDH+aqMnZqmCYlwpNRnkhgU35f3dTpnYmFrtbjbP
m7kNhC1vypHJGzWmaKqFw90DzKFxQkoARYZcMCcTM0RYv3nE3B65/gVx608Li77I
BZ8YS15oBzue2YpkK9FmbNpTo2PHg0ZWekqVsjY0rDzKbBxMZz0otB8T0MnWuGQR
yAczG2GMRmqc7pZFcxeEErjcWtergTqYqXm56dZFrV2Z7geiW2hH4BN4nIrNuXNl
pLVrFG9pYmEBq5dTrWRvDa6OdAMxr6dsN/NMvhiN5bp7tbInrU7WSzlZtIif222N
uT4aEoXAV7L2gpzz8b9CquO7YKKA1VsIb4b4GzxKPVXSL0+oHV7eFA3m6xmQtoTu
Nd92nes0XIXBfwzoEeywPxGcOLoPA2N/SfkFhp4nV733hYcVj12odn5OgWzhNKZI
EcTaLWPv6A1TGo6SoPu2G9e7Zs9xvXX7e1ZlbWi7GtEBGeJ1gq1beti+5NgBPXEE
ZbiF6PBo7eu4XYC420nDIJ7QPq0RFtUq2D+hkAv6fiCiSOdn5BgMua54uyIlLtcA
kmUkiwaKULd2aC9tQDGjwTdPU36hC2q6NASoUyhIaLhgrZ2Ha2z84fPnMgEzpnTb
duzANDZdS6ranfw7YdYZJw75lOq4U67ZgGU9MiGPbGJL4Ob985b2O/OH7ZMdT4c0
PJUB4zuTvaPaeCtEsrtewJ4dl5GdKBjvBlzwFq8pXPWnGNkN4BBJRJkT3mzGpjZQ
BeK1OMwvMicaudqus21h04aH4HgR8siCCiMH0DvJ4dzeijj1g6Fj3OrP6XjkMDdg
yaC7+NE0PQlNEdfaiV6SC3ZUTbaX7Ahg2VuSM0vZ6KmciFGcnlar+B3SysLIFuV3
TBw4EAbx/LmgtRR6kDF6y0vZYElHqHxgHJ4GADdGp/3BoaFdTLGCZfX1jClwq4Kw
L/cDwOobqN6fezNbm11cuHQuQ9w0N3muovEVsnio+uhytGFw8+UIZ/5Sm/myrFs7
X4v/bA8nhF8AakvkZFUd7nWDgzY2ApaPB+kDvqgjZGYiKHbRnU4Mw0+0QYoSnsVI
ydXXZ5B8/bakMkaAW0Ti2dKhk4T69hwS3g2dv5EaGeEkBHzIHdmrlxe7lm+rTr3r
l/U/TprdoJ4Rxcd3hRd+kvwfS57bMKEEDJWjfda/1cy8+O8s2A0SXvE6qb5EW0om
fRfPoxT/BiAF5o4nZ/XEAM+MOzd82nvp5PALVCtPKErKQ6acWSgpeb7CsV3eXNSR
mMY0tIZXl/C/zA39h5vkpcGfGsIfSydHRvXRnanoHlqnh8C1eg6Y4daC05bN4zAC
bO7K8OPJ96OEBT0FYMp2EUpEX2U1ce7+r0pjkwMt2tn7oVO79XCJAWMXuawRh+Dv
u3RCqUKsAdKHZbrYx/IhtiIZcJ9o8A+23OaosMsdP+cgIkbl78Jcpj03hDb8e4Tj
fdoxgkZ+TkvNkvF1bhGNxsJ5UfPetDAycYM5/P8w25VshO/IO1VEKbmg7CLENxl3
Z4aqvHxLuN/g3ctTAy6v5tdiYNzSW8vp3LM/Hl1Z9dQVOTCKKcfH84d9aJmXXi7m
ae1ayaOL5R7WRY2aiQ/h9OOSBw5oMTALzUleG21/5NCsSr3k9fmzCFxT1oC55xD4
TysocprY6e982z2CE0YnfMQ3/N+Tz8Y/cvFC+M9nRpBj7LKEL9W3T12eoyqkYiGS
bg2j28LkhE68Yd0oRi6eSrSFYaN1r9JuBvp/ntq+sgLX22DJMf3+2UEVCZjqjUIr
N7TVDfpCJI3aPX760MUZh33T++ezS200WKl8bJipyPQwW0/841UhHU0mF5+EgPoh
2M8BHK4T5ED2Ab3s0Xq0chX9HvdgSiVuovCAKopNKFg6/QRHX0ztNmjlVy/ZQfIG
dNMuYQyUkqHXGLNMRbDEc90IDbxl0bCkvQ0LahmkLuyMkA1wgnK9JPw1Rs++qqVW
6s/V/xlw7gTckFq49L7mt7pvOAAUL6p55kwUF3kZ3AX7pOIhjasDVR6F2cwk8nfS
l/wSohrNyZithB+Z0qqCje+GYU+GmfUTZ0m97jUBh7U7JF47mVGiqBWc+anlO8fu
psXmG3tauvQOgkrn8AqkoFM0axgGNNvdjmLTPsApdrAfQXuXYT6NrvlJWowIbu2X
+adFyuFGi/fCpGkSKQclGUaNV7LNDR2Cwvxt4v5WXk8ltaoHrFhexQrnGxmWuJFB
/taaytzptqpKOfNyqfAl6xHeJR06tvr7y5Tfvrihd5tiCjXEO428ZfBODKYo7q3O
C9C6RMjkXMArUvCHjWf5py22LjY52/PMgpnVk8BK7Rv6fLEC7lWT+p97eT2fCo1F
jRbjNO81Ef31Ys/Prfy1UYs8e+rgZhY4edYr6H1R4iGEKwYuA24mLCmRSGqG+1jK
r/uESFRpm8J+DaiM99+RbNftiwhoN+YDwmfR+8XqI3xsyrikdFK5DOHSgZcy8IXw
ovcj2q4v7T/45Efo5iIRo0/cAcCBOkOKektTeWFtgt9DgC5FZJSF+9Mbf0oo4vSf
ouf+E2yqG39pg82qIqI5fJ+b3rAK1M6krOtKWFfc8CG3GUIyGsWJS8dP4P8Jjwq/
p6kKu37mzP6qhHWkMMcJJatIRU4jLJHBvbSfk4ZqR2Qp/28lkRzqyqWRdutR9Sdz
pCq0JMOFi4Cw8NFz/nGNWdKpdVng5rveolktU1mgjvbCo0WxJmqt3A8nnPsLJXh/
SOsAGuAqnM8PfGwga14iFcVilvfByjjG62f+ryTAQ0WHwQb/fylvJsvDVTwtv5E1
oOlmEb14LVebuMckcVzFCt9EXehTDdO4vk1rq+GgDbC672gdeKktKuze19tx3yhe
1paUPSlXa77KwFZ1mDSayZl1L+gZbiUDNSrDB5axCU/gmB4Rl154CqZvHiK3aNrU
vVaiOG+iJFvhJnCev6BwV3g2oFhBrqxPeo/T1i0EhzRuH9YMft2nivSnI+6cxrzl
9orn1OI8NPYZ+Hy4HpJOth41uJRhfMCoSYNTPtfx0xPlFmIVrfW9PtyW5Ea/GM0S
A6E/pVSU9aG8oPeR7sAwgQLORuW3zmlb2fjvonIt5TYVaO18ZfReVKk0elgtnB4k
NQpftNMU2LXyIyrivyef3lpNbb9QcmrneEKej4m82x3uHI6AhDzW2fxOzmxsQ/Z2
kmSFALRICEKZuhpSCHSnptecZ05ItPrPB42etolYzFa5khXx4ZwdrjuXpl4CL5+9
ipLZ985AdFDZS3w/J3ErlizGVVqYA6Oyzhfu1LCpSZLvlZ5IouwKymORdtI//eu7
t9nm/R19+riwDlFO0ACLv0Jsp4L2Sit33+1n4Rf1JMVJQIfYZa7q2r7+w1476BW7
59pu7yAldRrfnWB61RvhbhWqxlB5GvunLk44G15LTlY9PFe8MndS26zbdt49MDNI
ARIy3SfdBqhJqqGPNUIG/LGAzaWgQgsZNnE0a8+3ig2SH1pjVPWTG/RBSfa2tlwy
G+0G/g7+IzcNNMJL4ScgJkNVFC7BnWxk5H0pKJxoGKBz6Tl+FIQ6vJpEXGZ0sjAM
T0SaOjs5NBo+6UbFKzjXioZ6V+azfYOh9rx+eJUGgX1n9V+d86coe8AU/1PYk7sH
p6euHqsJKqaKJv+D8vrffB+EpwHdjKIOHc0BkNZ2XB+GBFxPCk2ZsZtkf+mqxbR2
vX0WwaloeoBIvDAu0WCWjx8/uJ2rTswthgzdw5vb79creXfGW2vxE3G+FsFVBd8h
z/LbNta09LcGu1Nb84EQUtDwWGJ8SK2aRdb1uiCXzAPTrEUgZ7POGhUwfu7+7p4r
P3MSdXTSihnLSUUER4nvRJ5EI2d7y2egeW0eXin4y5/eZLPX7EGuYsltHp9mKvFE
b8JkRbV5Ef+xTRzuT+ABiHmHD6kq05wXwAjFoh4SAyGqN2luJi5UGpuY+SM2dRSN
tlTj/2m1yUpcp3XBL5fEl+r+gdyG0DLgYEgbLvaTynnZSG2awUyz34UGSI6n80H8
fpQx5MhxKxxvQtAXwKgooyV5cG/73/rbAo1ThlxFgecVnzuLdzHF3FJ+nil1yol7
Zuj55zabnXnPoDJ2LdLoEZzcqx1F7Q/QMc4s6V+cDfwHYCYvtByOoI4QfIVZhmip
O2JD2pJd735+D0nA3ly3L5PvnTyc0+3rn9Y1HMHr6k208AeI64bwfysdHNiJuX4c
l+wB28IW/zLnnL8nKjEQroa6q3azSGZDwDpbDfHeziUnvze2Ei7z5j68JrH4zbrq
Ol5UZ9zgu9EhFkJpAg5h7Of+j2IdUVcxosbcIcS3qdl8x2fGdLd6rMKI111I+kK1
zqy9NVa9pTu8+/0PCYdpW1f/jhfDaqFEC1rF2glNJ3vh3xhWE5BVmGAa0zsjvpYD
R/hlHKuMPXWByr2yom18gJfaBrmQbpGjLVoD0OM/2uJEBBM+AcWATPeMNwtls9+l
tHJ/j9iXuCGtjo4EU2z3oBHfSufopOIYiWb0FvtUo2PYqGdd8BBTlKhr0+gb19lh
wHtHdS8VaRwuiThwQZSCqh9BWOm51PV8HGZGAxsiFNTzk7oaC3Q8BMBQ3B5kYsRR
AbFQKMEiVi2p2FI4M2eE0XgNLoJrjPqD9FlhtFIEI4xbzORTDXNai7wevUyYBr4R
JkrglVpl1tGnVyDmB2bgotE+UUxNXplouO/KQ4MlgdTs2vT4E1FyCQpNWQjSjfEw
QM2fyUvHXNsFvD3ZecV2ZG/jlbNKSNiCYOE8Ab4opD4NNqC+DiDoprHIiSelivzn
OS53M+StgpJtvWldbuHnmX2Nci3tmbDjYIRc6u9xHfl83+uIaztsoV8ABTNmDPtO
Zicl185Rcfl4XPzuBzkz3rVobsmd5n3GY+HaqRjYIm0Eh8zeCSRy41Gn+AtA7nEA
4KZaQiS+FwJFrJdBT3Rau4eTA90BJRN58DqDAn0nPP6FXNWXxPQcMqIRvQrX35kX
9ag3TEotxJyGhwe4Aoxgs1ILLUgvn7l1074HwZ/e3DhbiYr4F9ibIemWc9WCxAi/
mOvLCeUNLZWoprQ+qIoN+CcN7ifri3zSv4yrrUhIYktTtusjBUY+98j5RRNTAtp+
gmVFJjMfX+T8lsv/Obh+5Nijk/rYZDJWY/19sazP2zP8zxb9jOF9VJ971LNssv1t
crEaxoTuYcoRok6LK+PLWWKU4CigqzF1bn21gkldXTGw/7y8hGptizBrRwSewupO
m6ew0QFd6wO4a2JbMsFdNsufoYY9VCNWC3NYmuJTAAYRYRHmla6vq4K6xg/CZBd/
lF9K6XFzM0lPc4zzeQAvd1J9pj8CvNt2EpQNQfVIeNB4F9HmLk6g9zKYUqrGounh
C24jr3c2hb/HjCae090KmQIj1lnQZFuHUUeYcGz4yqkiLPqBTxsxTUV5tBD6zR1M
enDtVcqdPX3fa0PkkiZgwwz6esL5IZiGY5+mrCurSE+IJws/nASW8Z0CC4RcPirW
RYRrwclf9fZzMDQix6HvXjtlGTC3574ErSv6iGwOBQXjbgsHbhDPg/sqPeQMu5MQ
j4s+QWyjntu67LrzjYrigTxKFpIgtMpnKcSB8yqg11XD8RMYgYCB/cBhzYvlde8H
fJi+IQj189/tLTqsTl6bvbyUBJ7r+xiRSpaFLP+eJxq4c1UV1M76p4Z9MVaXsmbj
rIwJ62q+uph6ZeoRpp3Yg4DecTYaEnnJFryV/vZUSz6ostm4cr97GyC/You+8VlJ
tpAZ6oARdyg+W9J2aMfxzvtrVQ6e/t93WwQG3FzgUTHIxk0Aq74rqm0FVK+kr0H1
nOXK8dbj6bt6aZiupervEx36a9Dol9eqvOAReqsKemahiDYFEMm+LiNer+Ub+eJT
wYo2gcUa9MpvIu9W+UnNnxBE5licR2JnBPE2djR8r+Ez/M1Bca6gBQYv5A3QmyiP
DaYLbbzn8IJGeOqaeJcsW9OMXxBQ8KgZUSkvPYmcOs6CAXVm73tAi1xvQYzaJEen
tixDWuiFBlcw+eRo18icuBaLY8R8lGWn//z80tkWG39CCavBzGY6V1muLXYao+sP
SGNVBfmH5kR5owH7PGq7P5UmxsGbCNNxK36bY65SToQtP3GlQ3H6isxMloZkddGN
1vUbKqKErsA96J9XTliaSOm5J76ilnZCiRdz1u4wwuugtc7731RfbxFcxBfiLMgu
odLp9S353Hn9pJbc1WE/e/fN3ptvAzR2QbWa7ln7KAtu8LLc8c+2KKwYee4uB5Cj
XYYkT5pAlvOTsoyvd/KFhFzVpxBcx5kY/2KDfMD9V42FT+h+eSYB59Si3h7/zRD7
1D7rJ5xm+lBHJWKB7bQj1+vqDFMtz8MbOo8bqeDjZIGNBb/CyTMWuR8eStcRcvWe
i39Od3KtJKd3fGu8LTT3Xh3gFixIwTPMN2c5FChNsdHMwbR0UQWYPKSsb9s2i1IP
XnN9Y9BvArPAAqeAF9DfwOmvjMeZPsAzQUe/NyHncBlJd2sal6nyT81ChzMc9BHK
bhr19hk4wu7MPIcg7njvx9yF9tuAhhuzS/0q+kzIi19r53ajHeM4RNsZedgO1f0I
Fbkxpw+GR5WLm4mx24INmJ3n6qS3fgOqiun9oThVNIIDyO72bH6n4UrjFjykf9Y2
53TXSbYMJ2QgB++esmJ+NEwj29808vN+iXTcrIo3+zQU31oSfHbdOgbw/nbnnePa
IUW80ej6WUxdnDcxKU+6ftr9dO5ST786reamNRKVkgvxJ1ceHSKq8cWHNO+iHTHi
48sfO5Begh56JasMpQATmf8YiuwOl7l2ZUbQ+ijR38ScAbl6aAMmvPduIbl/ZDSg
/5c67M/dSah1s3R807lF4SL4bwv/R+SE8vEmbS2hPwuI6P5Shh/h9PBwp7nMe//b
QEwHTzIqOzf5euEwgvajnHbVoaB311FOCHzeQEuOhOjZKmzT8xTsdjM0Z3Tp4WeJ
g8DWL+fhL5F/kK3fBt0PC4DeE6oG4Yh0WTMRUbyJHO4hwJHHbx7M0aRUlDveYn8s
6DFVF0xrICk6Pgw36TZCH7WMTHTYqoIyDHnxqqsIsLEC/oq83NXv6F+wl2qxCB7M
FSxETVe5zFGUGHesZxDrmyAbYH3yIgvjNmdE6RUoBjO8oRZh9e+vzqZStLtBjp/M
AxZnQOCSQ51DZzI507+RpiwEg4+R0iAJfUf53cH+aCCs0+5T4GL1AGBZp2smxz+W
PlsdNXgdv5pdCYOuwUzQDNEtcmJGetocXhH+PsJPZdXorkl3R2XiH03avYyesRu3
Sr5+aI1TbPcM3Lml2Be88BK62v1/cdgvw5vQAaeVsv/e5OQQizYFyfYVU7QNt6v6
Q705LmmlyLF6JIJAst0by0zI5Y1qDBDlBPyNyWZJeHhKwcZ1W//zvM6cQjlR0Sdm
VK4kqNWzwk64qqvWCUpLJr69DtoKXAlMlQ4uRf3UbJbVYXK6fVOiCEBxq8FO/K/K
S3k8zef+bjKBK0r1Sc10g3BmmGf/Nq0aPoRf8NoE/fwgD2FKUqw6JqzhvclvpgTE
kVIqi2esSzzurqnTfOmH7gf9UxTwl4I/jJiWN2xfmD1HYQ0joMfmnXNG/ZlmXom8
BrLFp9ysBZGIFeFo+3qvAApjscuxDO6VxT7BO2j9lCVrRTvBl6a8v2IzHK4rhEXz
8/LkG6oWuBFbuLoqT3kMxVMrBQsg29c1J8mdMge6y4lGVeKsq/g/KvHhFNjoSgWB
w5bE37eUjRGGelILsq6nP9x9dfbbiq8dM6+JAu1n5++qoIM+fEg31lCJFQHs58T3
tjKmlcpFVNDtzSFo8ZzIQeqgALEf/jbrKqdlFpXfjInj4DniDntxrPglQlPgkHqZ
qSHgGEcdD6Y6ok/q1pT3HZzcsiI9USZ65l1SFjhQ+6I6ghDmx8uT0QO4MDVRzCob
fXfkpzjBuXi3E9lJnpjOBZ/MlvqWNvLI5KBsLnDYhKxjNc66f5y6epbTOxJmDmKY
5a2OTKnkkSHf852+lqER53ELoJuI5szIWJ8iThmryTM8HbhMC/rxx9yX+jcIkLEB
8WXzd3xXAkKLs+sZ4Y1+wrRPF+QD13RjJen/ooVtBLqZap/xzMQFkyGqknM4oLmY
QNGEVY54cHvOi+cBdt0/zH1fVjPNgVSV3T/lOm8tzWVj8eqSaM0If7l/pJ82OADj
mIgJyKCrgevDjohwNUQNMBwlxpSSKdrQjX6XPEkUgk3wXDS1CM05HmMxrfHILkez
r00iYkSi8AxRYgYwWBlIqK+G3Mypa2gTTGhnuT0Q5RRlHF2+yAsYgMmX8lFlXm4X
XGPv3L/7bJOJSvQuHTfc5vaHN4xefA3iNlM9eayTYIDrDLUymXWB2iahVjevIAvC
lnTIVTa4oWH4lG53Zdwwa+DG2cDHhxeCx0dpGQQlvTw7BxJrNXeRMy6JT0ZhDqtH
MfYrvfPfuokOneUz4f+da7nglPxkuzpB4M5U/tCU1DkgnQr7tJ0pwG50WxezZsnT
4YKdpO0AeKmjs1f1o+Hq9u8arAYeYhwAU5rY+FEmOcENUjImn8FADoP2FUqVoAYw
AtkPeOctdfW1MA5+vsqOJbK3ZCyx3xl4Jx7Dx3+1Sve6cyE50oIvqH97Z8RF6gqC
a2rtE6tUsK8mFsuVaP6hkdp2HD0kW6IbuTl5OtR9uIPkHpEGCtcnMkeXBUMfi3g/
z4ee/FTkDE2/2+dmQ1XzwzD9ca0+FfCyIUfKegJAkMDQ39Ijzpk0R0Yt0ZYAVimR
lmEYCi6XbMusPvP5wPpcQFHYWVktTkqCx/e1i9IiwYn43ujdyxjrGIIWA6HfZ67+
8xgO8v0UE1OdNmZ1etM4Abaw518zVLab04dExdsOdTlNFv5HSPS4Jxx0nvtvheis
tA2zhftBuBblAZdwPh93Nvxa//byFnaGs7xNMnu1Ll2e8/Vw837T5YIzunbfDDEZ
Bgs46MQ3+o77uDU5Lcbn8P/lB/At6VrKnF4veOmsb+TsI7UuKZUg+8Fj3ARQGKHJ
Q5VSyyR9Gl/40KGKl29k2HjJ2zYPideqQj3b0NVfPHW8J41qqr09Tu0XHnDiuIS8
to5bqYvvIOw7w2IBduPjvGnoNmqKp2WUb/7DmyWyCf5Ngz1bfViWICpv937OEi+9
s0fKEjadlGwXReKxHIPjL3t7o6tXNdGOg+ikyJNlc586NZ9RMKImb523q9rFL1Rp
aVebIXWn62c/YxG5P8V/yyEYTV8BjcaQgV2qWWHkcOIufKJi79IGiQuEne6sHp6O
GG+XUJAQ7TLGoVndt+QKggnUdbALvpWxa66vH3M2TnIMYcJ++Pn6bvqYahNlQYUj
wxBD50mKel5HCMFP8AqtZoMURuqF+ZeHxtY7AAVS6YqnSYFrvC9t4X+NkviCcKzZ
BzqljF0CXmzzyBf9UvIyNpK72XuCM3X8uq6Vsu+4jliltG/X/0yX+YY1RyaF3P6B
OTRkYYvNJqQ5/EX4FkHUxniK77gHdy7c74dzYMIPYNn3Yze/CQsizbGORLTzSkQp
kNdnHbIj3e1iH10DMSrajp7ekgYV0w+cRT+Bqmvq4BmBaaULEcwaVMfNnazqBkel
Z3F/ODRyo39PTz8XVl5rY/0bXkH0lpmDCZusE7SSwPXI5G94pFoRLz1t84Z3I/pB
ta4JQxJ42gJl+/dTIFbcoasTAW/JPlGWKmMcdPjso/fAhCUXsdEschguedvM18V3
Q+PmRw9egv67HM8OLGMrSWQwPQVlvoV+Wrean5to+AO80fTbV1eHZ9evdvHZ6aGB
VnFrUqnHyB0Aim2oh7bzXh5rMOscYU45qbSC+KM0thIHJoViAOLjLWtHjMK1pX+Q
mjruHJWbZXVJTZPyBErgVLpDjKWiPi4IoFg+AI9TVM5q5bavEXNngMfMGD43Z7Td
VL5MMQxYXbTXOQEzKZly4lsQs/8zKE0qVmpazjgrl0EFueG5g8ikTN4h6wZt+yAS
uPSxoZF8EC6FnHMJErdyVHxEdeqJIeexe0dfmifgbNZvBeiTzgMPhq0PD1h2Jqmb
Kg0mi2+bewX4ypUJ6pu//nsQKOzTbWqISQOMG4U6QPcF0YLPXo5opJrZ8WJ7P3rI
8d2LmDEGb0J2r/CBvhyrEyq9hFAR0EdAhaD/lciYUCgo2c3dxdWUQGnI7Pz4R3Go
tI/3wL2TI4vnHHTd0mFjBuvtmrfwtO7UTuOy/zVeCfohVPJ9WiaoF+Yq0UY6S83R
GZo8IeeOXGjtmeEvSckbcmCd9pfCjxvPOxnit2vK6sqPbz5oiYxjtxiBl5yqxhuz
h8r2Et7E0Qx0LDxdYnkkyB0Kfs1nryGK2GlmIgo3XJAERcPdrGhVPdG1XDhMINCl
/NbG6ir/0kPp8KFsnJinXrvUwYa+e8BykchYvIX2hkJPRBNSMHYbaP1BpJwvYIa5
OyjFhsU15fqQNfdq1pBcsEX6Ni2QfNTXXIY0BrWHqlm660GB1cgkGuA/sfkagMjG
a1iQxJZnBNZdTA+l1mq4SgdtGiwpSUHsQg4pBpMPJGw9w42Ig0y8tloshM6WOl8u
5Pr8KsNF6LQlbRXjqlwA6IxYUGzTfFvZGbEJeuBd4ZSnipBSI4h082eS1ASvTRWL
z+0UszhOFGYBO3MVD+FnLJwwTzQkdwLlQhRn0aQ3C47KsZNyEL24uSXb6C6xPTlp
LdTb0xkZu/T7FQpAdHwdVDU8qNO3FEZfhapVaUbQ9+142PR5nybzQsvm2GZpCedY
mzrMDp0yCsrxPhVT2ueO8bDXEIgtgEFrDVOV4N6xfh21Mnfmjwy5buu7LJftjSsk
8oNcTovw1ypn6WkrcKOtq+k1kS7+bMvIU84WCOhaFCDIJZJUE4NF3KSN46xtC1LZ
clv18aP+I9KQPZxNga8OgGdQRKdZeHKd2ncPJSgApLAnvNsT9Ch/NmYRh0GSLJs0
zNuK2yrLCniq5m2Jkeuyz0SMPpX/VXB6ht1BF3DacjUeDEnbI96PDHE03C67tOtD
ucE077PqTQ+7fHlFpJPdGPnFP6cNxRMc+0czSC6YgF/TSvF2z+aTDtin+0T4t5Yk
yIq7RIiIq/o6rNMq5GbpqVIFIyt/nehANHW8Yjecg2b+pujwQtXbVV+hAtEoraL6
KCxR0XiU83Hrmpxoh8MXBHwyDeVVQdek56DC6HQLHA2vwFwKWeAtMLgG7+RFwizz
I60WPSTHE73oeentTcxlDuDt07YKPx29UmyFjNo940QcANY3YqbKDTalB4TTuvTP
Hr4rpSpkM/c8Ns9KxpGEcC8Echyb2at8O02l9JpQVdW/U7E6GlVWwym8fh3hjeuZ
m3LX+OxmJ78CrZIP0vFoXl9myFqlPwMt0yTxmBDIncyjrQvOAIkRKuG2y1udAobJ
11EbKSXOeKYGfhUg0s9lGseAg/BCIvnUyRyRipLp5HM1y5MrvyoIHGEkNYHDziOt
pclPuzYXHU0eN2MjByLUOHWw/DmHuZTwatmyVQ3449YOPVdps3khnAvqBqVjvbCi
DkDLExalXO77peIUQ//LqpYBfFkT8rUqcQKtPT/SP/3P9IFhcauzqXKv/Ubf/+1n
vXHPt15jzocHksAP8ASXUMmUoH7mIkAt/O9CD6hPszD2DtaGM5cuq7J6A1fMPczy
iOyiOlKxvg9GVe4kNgJIsr35/Pp76JgqSprdF0sEy9XUOQUpVguz/cY4+uL2rTmP
NkRzGIl3MUkGTMCKkp7ffgFLTkR3ejPPLaTWe5bytZRjXkW9NrRwTHRvyXGRy9za
XdVpIAUiJMtp6Hb3qesB6JqPIpYB4vhANLEoXuMAAwzUzRBNxFB3yJvYdt5U2LXp
FZVpe0L1+gS/LrHTzyD9+90ORb8Ch4VliMm9HwdiKaSCcCVgKJVeu7GsrFACJcDk
mDimNMtAgzYoRzkadp3VlDO6bjfbyi36w6QFOV124qBzzQcUAYMDI2IXROCq+a2s
nx/BQ4GX1bUZ7q8g9f72rqHTyRCDk2w4RJhSHaqBid8RweFSPtbaewI1S2XQyssl
jOVVfJ8/dSuTWIvG72RwwpEiqmj7klpAG6jnHpXcL6NB2WeSY6/VyNWUA9qBlUSW
vJOQtUGXM/NON3QKRQSkgIoBlYjEOI757loi1LfKRaXs/kC9f8qh+0kPluvU5UAn
5yBkNzWAFmHaE98m0HvYEkl1RB3FO4UejvdYu+C5NJ/WQ+wnMORbcLvbSTTsudxW
lwdo+05Bg5s+ffBX5N/mszo3X5S/gPnPCyMrEyDTsok542KRDKVkfSNay+8TF4As
xPCkJufqvV6/8N+esuAJSdxaXZz8uM/ZP3QwO1Xa7CsbdOb18UwtyLRoW39rorS1
DIbT6MaB/yRxZieKPS8dlmFx9pjCaCkwuajC9QjJsX8fNuf9Uhv9imHZ/Ca7fnjh
KfkIWIgBsJTOtzj/Cb6Q9oxS2uTdcsqHb/L7nCWMEq6elYXQCC3RXdBkUSY7ucsY
GB+eJeM6KszQ23OzckoGd+NumopOhLmtkVFcqtTwXNa2iUmDEKZCAhjgWDt4oMN7
vynocuq9NEj6zN5BxiVV4hwRBJwaW0cWs16JV6ABh0AGJImYQfLTYLrRBY6DWMVk
r5RwrBBuy0Mqkz1AWHoWn51KA6g2htR3HpdJEzJJLw61sVxmuv2z82g6XdAx7w2E
8FczpgwBr5ocU06P7OvaIMbo2w4ukeKGC56KArVKAdcFWSoitBm597OcfmRuedij
wNkKka3jmO/v+tuVTpXGBk8FiMmMAjVM1s+CZHQ7dmoJqMLNXwfjes+BWE2x9H3a
vstvNzQVcOL424L/p/my1MEFK1TyDSN5r5ebpqjlca5/TYKvYB7k0xRUg7OqMY+h
AR/e5YwFyKeMenIy/3AvJWNLWVPLW6ZxL65NImymLEJFlUzTBG6P14uJZrDzsLnv
DTIRSEpTSvexP63dHx8uHgF83186EnPXT/y19okn1vNEuXqlnMowTcI+0vlfHYTv
9/dm4MVm1U031W3rC+qDT92szgAozK/4yudExFirZpSDrbpnLgTnVkjvTOLres5R
C5T6L7+9BjvV6rqjY3xjiDhE0ixLtuq7PhxSQTqLAqrxgS9jDVHnBeMtv+xCGvH0
gtEzNH7KyrgXl/FzClc1VXIgaqK4bHqLQaAO9oAgJkiUyUxtsXDW7V1vRgTi1sUZ
S3rqq3fDpp19B1qliivNAebBn3D6kBDPsRDryuedo1ioWn1VCR4n+zM1L3Eu3SmG
bzCAPO23IUd4XIzWgY4e59Hlk2nQ6NmvciK9s5KfO5TWpRpfQznG/Es/fJcxrnIc
C1MKuMT4YYVFOESSqWrsYOYwcKk7H2Ula5z6N+bXYav31zXJMnTxf4IsJGFvZOLO
SenCc7rQvI8npVlqx6VPaxfgpex31n2hG+OqC6m04ujlK0LzYFfc/+0eG9F3cT5N
FXt4zC0UG57M3ylHfn+sL4zcpvD5NqwQ3/tHtmswppPWOFvzoEe/jjUBwK9i1LI/
CbaALr1uRZ1zNC8ZuEWrfFX3EmYNWyFh4Iu53LrsFrU+/JDwvKWvYABv69UI7HyP
FYOywnkJNL0uoUaKrHC7mgO02+TcWunlnmEPOfomvTtCVyStty8wxm02akXPCygS
Izgi0w6oYxv1G7OSenOj36L6oS4al9VDYfK/XuGrbUC5uXz6qWCRRk1+F7Nmqvxa
0yTIp2u/xiuOYgvRnPGDAn1B0wOmvF9EHEiV0A4XuESHeSud1xxIiaj8FGHuFssy
5kP1Dqaqa+ffSy0RCw7629g2MrssMNB+M3XFIk2HY6T3QsLHK6j5WchlP+lPqwJn
Xvq/++q+ybf+Bkhg4TJyMhqEwEhtYNodlzuzxAYN29nzMMArBeX2Om9b7/3kaIkO
JaFthsoKxX+v0k85hXAQOLtxpgXZhPcqzBufrVsywPHNRnP55uiArDXEqhMQWcab
ZLMvdrt+W4BfhMHakzMBqGa4UTKA7NbPOyTwvEHmHiFiBo+oDL+LO0nHknQTGPWe
sacqeoq7joqoz25epNqaYYvR+NsJUug8yQqCRYmkYIl7Z/J11f+hYmR4b/KC3Ccx
FVO9t/utwVWknsnHckKu3xjSC5QbKZNvXknGJV5SiicuMzRA0o/DNZr9T1k06Zcx
bElbEqSPoeFGUk/LxFzSUpEj+WnEjO8kSSBx66x3kQHlhiAyLeGLzsPV7tk457kW
oKvSxrstHH/bDxnW22wHuZp4QmhfrZtiXPrauJkeDvJ0HfeCa/tIufHZFKO0k9d4
LmlNG7avZ4wWw8HfwnQITnJGgWWUlEJrrFVIRwaWGu/iDAQICkBkvjyjmAevO+tk
DH3ThQEOa0cTdNp6N/nQQOll8OOK/Xp2D3mL3e5Uje/OE2USN8z1ykuekkkSsAEm
KrM4Yi4WGd5Qk+670YpJrIAZ06n2gFpRWi/9raxorCQBuQz5ZsTd7e+uf9YRq0ZK
JlL9m9YwHHuWGFxwwMboUuFg0EU/pVStPXUIJEflkqyF1/Y3UUqGo3lhcLrVIwv/
KSMnBW8uAdxBHtithZHnGhkaQWam5WoqK6hFRpfp7aZllBWXqUjp5o/GY5zaspNc
c4Zl4pKtfZWlOoYDgsyYiqQTsj/nxeBHTx6lPac1lo7GjLjuMx84NcVnmEvUnNr6
AjtrlI8DZdEAN8MgI1nTNhCqbDaDfMgWgDJcRAexsQp4odcUKTelfGH5DBfp4AUW
nas4xKBDC7t4u3Yog7AyLzM3R7bkbC6yRnBV7E8UwSSuKwD6LxcCtAh9KMijYNfU
V2UOlWEyJn2VtM6AcUQSoPIymnFzlTcqgddxVVLyG+479FDQRGuslzrokUSjWd4O
gwW1CFm3e82ITR2VJ67JrhPpyHk1xB7iO8PdujIEIusgo/DYWZKeYGJE6ul9JTl5
1/4mTxN5htTUFqS0BfGfebudHJL8hXS1ez4iOwvdGYvGgPOe/0knbUO80BMmxhEr
BRu0pM33O7FEUt57BJuBRsQh6A3j8le0smuG3G+GKGVoLX3VC377Lt3HCNL7lDzD
Ou34d8mq363b2mAbQmwA9VI183Z2/LwSbYC8vSLEeLpwRdveJyP1fDa7oVkcytq3
9D1Iobkn1SyHwUC1GpgWYyALWvAUm3AiAqLgP9LGclxYifSSMJcMkw33wF1uH45R
I3A8wtq3BDxfcRTR5ilrJRnzVklrPRwKUUbcnpRUGNpSh1sMdQhB4vIvFbwZQZZA
ZRUSScWq52YR24EUr035iuecZQa7hq+/okGzKeRsttdZlWakqohOZsHAAIvM/iWy
3rfu7V/TYKlFY/joFos8WkHd514uMJbU6+V7kzsXQMHNCdwoqGg1+iEqNkFdx6vN
lygWu1YoHkzo7vmpOCxvuEameCIvy4NCh7xbAjoCB/bnNbfkgR/H+Z6aMsLSnz2i
hX6V8TpKrdUon1ZD6KUQYJNusm/BiA1HnG2MeQAOxtmr9QYjnphMy0CYNEccHqlX
LvAHsg97hqfs6rCCQkl0QzH9jvAFWQiaRgVfakz8d1sjF5+YnrPLl2oIQ34pua9l
LtPe8k7+AINQ8+1ekT9HHzEUxUU8LHCQ5pzvG4rNo0mZOBiRNkNp70su6+h5h6M7
8STsWK42sxHd9h6M2mWinH7Pyq/fiGQlcslDf/Aku+CKFZvg+lc8OJUmzUS+2J2y
Ka98Moo7rtaSLoSc5IS7DekHkrKLx05zRaWrEw7BWj667aY1vK8PdQlwAPv0nm9P
ooPk1NH7rfoPEWxsSPcjgBy6sWqixwA318ewsq055l0IFkSXxTIh0xS2q/9ejqCV
Ha+Z2DPuhEFRaRgJ5/Immckpvnzil79VPkenfobcKPQ6wip4vI/4LoXydtHd4sMu
q5och7LP9XzHlRcDYviznj1umJqZ2RHYH74GwS9yn7bvmTT27iN6u7BHwA2ZgUPj
YSO0hlxjIumzVMd2faPulG2R52oMvjmztTJ+yVw4ItyJq2epr/aJntUb5txTRleO
Y7yk+nfZk2hPEa7xtZfTSThjpbMOIszqloXZiny/KEJDCwkuvaGYJ+yytLuIczWQ
iTZG8JIyVXHDS/LU/DlFBexbOqCgeMoIYhXjCAfcnhuIrGiU8HHhAb5wIXaAMayR
8v9/H73uF0eiyST+ZVXbxK5f8Dx6AbSZELGtuFSAJkBIdOsxz+5FSfiIa86NgVJx
6HhoTnUpmfJEoFt4xQ4QyQ5IyGPMdQvEcOZz6nbW0UMSC32lgn9KWfIESPTtuRU7
Bo8/xJkQDyFM2+95SxNDdWSg5oogpOBjXr7GgtlDdxy4/jg9d64rLoxWX+Vc3u/d
oQEcR4XjlHb4b66J6Kynn3y6XyjDHPCz/s33VFMPjJQYJQHN0pEnUdci9AxUHAle
RHM5gVNb18qp5W3cSkTevtzinPQSiswxXgoD1yo+m7LiLQs3S8NbdaZPyL64QblH
7U8JXwSd6/lyq6w3l3Y2UAiJ9kMQMzyLnCJREecxk0dKJRSJlVmKBDXaE31OJrHQ
15Fk/9Kr2F+9HF9sICIYvUAPacko8FERZ+CLa7xXh+Vdov7uzeRfhtuWNGEv3xTW
Hvw+LnhPoF8b5z4SlYZshfLaJX0szcknR3zyGUpPYVZT929uaI2eksCcKGO1E2CL
9KDQgs4ejxiTdrk3nPDiS8d9RpNaAeNdsNa0+7NhROniHpzs17lEx7xthJ80OnMO
F539Aj4Z5VSqqdfOjAkpKYjmLJtNx38oKg4HiHn53avP7RR7QoU59ldUn/2tf82c
va9hmebXgSbGh8o6Ba3iuK37bXae0op/BndMW4f0RsIWdXxbrQ3Lw4BiJR+8Kkwf
yarLEd97dP6PHvTsmK56aXxDBKD90YHB+/Ie8drh4ajnyQ1iQ8RSIcOhhPoZTHsv
C85wXdKludJWqKVGoc2LeN/SEKBL/dPy3eQbsIltLjGI64odekeB4StbetkSQwYs
Oa0TfbHyDFFa0ZW+WDLW6goVBu0anXQh2ZxAFTGcalAeZaXKAstQ+9qNf2upbR00
FTyFY0/nqPKQ/1LPsE/rw3HQnKOIXgKqC8mreVqBenALkgqARY9fV2ogU3OBLRPG
QDt18cOk5lcBnL/4W8MXDqVO2WKb+9vjKNATxZpZHOVKbyyAvGKSDq/l7GseevR5
cfXC4GrO0Id0thTxXQ5d7UwdmeSN5ftxuLP/2xEiQhVmwP/FQzZaM9mX7a14ZzVx
Jemasnq+96vmyWhhQ5LUymbaOX6H06gkoeyxA8vdhJGCotY69JG2NJn+pa6gcv10
fsTfG7LSvvmnZSaTDyxepIpj6g4Uhqj6aC1S9HfeJjQHt3GWBTszkjPLGZZnbCih
uLF6/aRYoOIuo07owaRDTYf/Mlx9kQJFHaO3cEAo0K/YxsT4sbyT4TkHzU/iA2gz
N4AolnMQA5t6ZWHyfJAyIz9DLiAZOjaE1LJW86ApEGF4zfzbZbs5MXpGtyp2LWPw
J9MB/ick55eJpONC/uJ1eoFb1Jnrsia5tSNxqrc4c4XMLM+vT9F4kO3iTXhlnqrC
1YnhNOrcNcmMEYnIk5FzXj31oTVLAtkFcR9yC8PSShDGQ4R2bwxrRgUcPlPdEdOl
u8cBUDRDx3VdD7/RbsYm6Cp0Q0RAnTl5IufrhFK4i4Jh3tAHaMaQAWH1OOTYR1vT
sei+yXBjoWL3z7Z/DKokBkS0HVuL5lkDqlJuWI2v1qcVvW88Rqu43A2AzZeTncwu
BqSOctb0YnsNK1slAkMQwkLNCZ/A6uxxsF4v4qXTH0Vb8Lj3sjtVFuQxPx9OmIXW
Z6A5WgbXYceHY5/SDZmaFTwhm3ROt3EDZcgbgX7xddfXIQoe6YT1gQDB+8xKiWwJ
ARu6W8hFWRKBfsb/si59Zq2IJN/KW38rVkWYEnfNqs8P2hz5YHR1cq4xZc5Si2Qq
aZEa+uIxNele3ioMcllYEI/PbidLUfZerVXgrQVHB4yDxhKDaj9wMfXeEJh3otGo
0AseoQ9d1FZ1IoUtDXWrJH8I/8JSKmVgjVVvLqzTI9qsxR03GtdXGVE4/C/bLlDQ
GOiw2dFVOg9B+dw4L2kO8ZpJ2DWcKGLMWjzRxrCQEi2ke07tiCE7L/hY6Tdh+PDN
G2jhcQ3lQcUB+fvFTEtWJHtVO6w6153UFRjq3ylkASCVVOVVTwwi5ee0Dct6uAte
ltRfwbcbo+oPd3kQe0nWZSvadIUr0VMaaXLo/36T7rHzlhn68pJ7SLXSptX6y5cu
DjBY8hC/HvDS4zRxSACKK+LV1ahr6jw8/RQs/7wuuMKWN6gWyICh64hg0qqTsG3D
GQ/xxuEzi84kL70aGnYRwHRpLYerOtx86CBFSgJsZv3lLxF9X5y6e0VH+LCQNGw1
/zlTJzcvWoqh9ZqCWJ0S3HWS71Abo9fhXZqxXbtrEj4uUHStvbCo+PKprw30j5YD
PU6OB9ICz+iG2eq/ob/XtfMP/G7yGqpfXO+qneNSnEng5MC0aZPicfFbGBqKzHf7
u8V8d09UsNs8LNcidNbF4YjkdsUPHEQ5BJr9dt+gbfzRWmeGPIxVWfkzsCSOFf9L
YnbLQfUcMsCR2hHTEoLHrtzDU7ogAmUFDyIkrB9yflakP35ZBqEEla9i8Laf+U89
HFUOswMoboA0HCwW350F34kqZJlhz0FobXFdd5yd/oYZNRwFr57yqmiZHxGO+m/v
DIU7nGilkl82YDERoudg97c8zoPwaEs9FePYlQvMsu0BPbJsG7gz+4ssw3o4HVBG
QOkHMLs7+QU8K8mtoZSavnBwRiQCKFAGpX+GCkjGvsfTfw0/YoTgoFzk/vjPFEGI
IbStCciOKunNe88bsEclLN79jpJEA2K/ocgAgjtsWL8qhfElKb8CwlWcsqpcakVz
VTJaxqLLRwAnmMN7ovfqDNDivepxdpR/YQeLbWy4Dc2TSpE6JuT3xUD2ry1BehSD
lAxTRwKHV/27Mw7u7OiC9aMKMbi82ySO/oZrSJuET3PL3QnnishMgXWBNGoseYfD
mp0wRv16ultyJ3Ai/RDEvhJ5WP+wwdaHNnRkMe3b+0y1Uh1jpoIfwgZYPQagmQAZ
ElI09oHatIG3k2ZL/273Eoq0KYPmY7hSWf/xEkVZq+1FnlAzzCj+RBaStNGwV5Tx
VFN165U9E7t3nDBl59tveZd7ypT5qUYtRbvoc5Ma0igQyrXxXM63jVM+M9ns2iLc
3mckxsU9tpB0rqmjxKF0Agnycs8QxutvQ4MspLYN15jAhzhle3OzhiexgdfqDo4g
FvD1C86GCFOHUm54SFgfxDGobZdA6kVzcvY38bpvYMDW3aoYxWANAoNV7+tnH7IK
mTNbUhLYCc3jim2FBPTKNEWwzBjogC8lhGI05VvueR9K56ewmtSV+nNQGXB4fBT+
ADZgSrf679VLJPnPjf8nA0tK1nrBd8jmTUkCyjl9so45kdeZ5q/QESHxRcG/Fd+Z
O13HDupQvh9YgiyeEOingyEXvpD1lSeqOHG1kS3NnPvvHE6QmtlpSN6Chzv9zT5G
4jHgluyq5YAjPs5rVNVzxOW/++rYtswUegppIIs0AJEoaC2o4IXugY+t65xFbVqJ
NDs3GFGWwuEuaI4DRKOORyrBCksU3p5MaNVr0wU8N6tWC4zl24RTPiFfF9WGja6i
3u7MHAwSpk3GBNJpQIiX0N6FqxLGP5xA19GlQ0EzSr8zYICJ3AloScr+S4DW3FB9
82mzCFE8p5/nSNrz1KMf53G4rwjG8hFKYbI8thVqYsrKdglHWf2AXWxPjKjsSCtG
fgr/x8IR8053fjhRbTXiD1NTVaJesFQu6YstiHJpD2WiCGAQjSSslv6f/MZ3AhST
dr51IyLHyoVI76oqCx4W4p4mo4sgjc6mDMepj+hjQs80pfvXcm35/egGOqVV0aSp
iyUg+dbw+cd3jxIxLIvMkKzcvxUuQWP+8wGm/6pkT9byD3pmTxkhoNxZgyHus4vM
BfmLTyX8lDmhPKU7zrJoUKB5KNQ8i0c2vISuw+JqbPJNlybg+FSmNvkVZLp4mi9I
5an5o+nfbOF5h8+uf6K4Wh4Vn5JXzvukq3yXjTwYllUAnMiWXhTPw0Yy8VyR4fHT
IrTry/mSAixWWshkpOp+s13FWIRdgGbKzODDkyRG47e0QojKeWPVmvHcvkDoKoxT
wkfKBnkubfUykKnvyZm2o812IXckW9k08BTfIeNuKVJHrSrHaE5uwJmIWgtt5mFE
7TeEXCit740RaBaUJZyimN57McdqQ/yC8oZaDzPpU5A3FxZ7XE2zjHJ8Xv/8c01u
EhcMPfQYTVbQ1VQfNpt3qoXu65dfCkW07Ld9wREkrfHRrfYtHbu/opusmnp0aaHr
JFlTe4GvbNXshypLKods/ltZ9K2yHvITve/uclRP7GrEDUJ4kwxsrCjThvfza/rS
mEDniID4KETYy7B8wDt/q9wp22QZHd3s9xG8gaunij2/bdQSEJW5/hVtWLQ46y4J
4HmKSpx8EiKz/JW0dcd+D+sp+hIFuC7wWmWUs5KWEwihJ4QlPeh9w3x9y9nD7d3E
KhQyUvncr6vC/vNFioYCugCbz5Zi4SPi4s4cNZhWRbn0Gg7Q/HxpXoAnFT2SN1IX
SOPEOphA2iwXeq8ni8XERnWgylMec0w0BGwlPds69r0gloRIkMGBfHNp7/YaJvCK
ANzyHldoV0nYRy0g2Kk9t1DkomuO1w8m1g6EsXonCw8rnfI9MBq0LjjpT3Nsx9LI
J6uPhP3prnCL4WmYO3T1wMbDzXIGA+XgiyA/C4RCkBo5OSvwdwV7H0J8PuT0Xjsc
F/Bq3zl5siR4UmlJIxhG7SThJc4P6miz+VJlaHYlIOwKQPVsIsRAW3ArtWBKVLWL
awEp9mjPOajnJ07GwOiHPqUsSkY1hVO1+oLFOzBLP8iV6sJkPFPUVXMjZZvO1nuZ
tUY02TFStehBj3+01eD6+Emvo7TJ3XTDmzd2n3KKjGapGJDomhVCSwKO4Rp1xGo/
GNbQs4v5Kx49sYjG7xp9fcslSMHs+nUCUt76Wwwt8y0QiV700N+YGik/4TmaJKk1
+edcrptZDdMXt6+hq0LXOpN0SNIeRUCebFJCtc6cOEn2psZZhULYQr0Q9aJBPmwR
txBmBHANQ+j9MA2+nSKll6klRGBAUa5GqZzOpTZxJtsqcg3xh20cDijOiPpTuMrV
PN/je87/++BqQszRyHIa4eg32DWCW6DqUkxCjjKhM/TNrX/leT3sJ3fypMi0BOrk
DG9WUihfdVV0RWamVFXsstKZR3UmZoUD8q1fPprnwNtQXy4umaRfoTzRyW8kP117
Sw/CjdDV0of/wqZT6ORlpjfTmcO0yN5cnE6iacVhKKOlYh3borU90GK282gi3+Bq
10vBX/PhmGFJC5nuxJkn/UdOkofpoiZrXs1ky/H2/fvWftn6EDUdaytv1y0Shx5d
gLK0snxUGuU0QIBQx049UqaWnK6k5256UHbxzn7ExusYAMm9OSxlxSV2zALC/v8Y
32Zsb6HOzDhkNy66aT63TJugz6E8SC8Iva5C1QYo++5c+W2bHWRAz7YUmXSV2pVQ
xs0uZzivzbN4LUxQsf/WtPdRKgwUee/7dB+e+coRSylbo5+JT4ApouCm/9t3vXqX
skuAr4atTgHlWUn0DBXsAr85epJBqtRRKOtaPB5AHxZ+xDYJT+7Rk121h4yPDEM+
kGoK0ITIrRY8HPZFsvov/AFYjx19TQ13TK2lJSYg399HMNkV/vXJL/KkYr0Xj37W
hcOo17HCWeMb4XJLlU1BHx5+h88A4zj9kv6IhUm5O6B6BmwMmOQZBENYJNuTD7xp
fZF8AoqnsujjFQtG0k3OwteaW7R+jlaFcBRiXYL+kjG7FmzudLezWa2rXlMQPwHM
2GOJM8kLj6jesI8rSDGgT68p6wg4KCN6oYslyF0L+5/Ase2iQ+1xtpLpPKsa/EjQ
GVDJ4Jn1617XSCYfdByUwqLBydcyS4uuhl/e32I8jxwRA5vVRvQQGMWubJz1e7UV
cuEm3IraKZNUBB5zPQxxCs1e4rwhM2+DpL7knYvxYaTSuvR/epYvpc/GfpJCFtCg
T1VggKa34zI5tqSoxOzknNJMFmW2gxkApUgAo3OTjbnntbQAaKnddZ3EoJKNmKxq
7uIfEvu4rfF4Ax4qhTqVVhJPA7Bp3HubUfv1m3R7BgtBM5gGtMhBoG3AdRlDjTgo
wkGe8wjI99V6/d5425xVhfJ5LjVMec/j4kVDZrR9ABzjbuLGbZGubiI81Bx8jFWK
QHJEpksx0MPQojhJo9d9reIuSaP5U0uraf1Bs/QTFZlfwj2kQLsAAcfrp5KtNbaO
Lws+8kDrU7XOznkKQgvUj1vDi+/dPiT3/D6U/IDBR5n7YrE4egKbYeRWi2XJ64xi
GPhIvHz2upebI2Z9Cg6eQwdNe/PXqmmA2vcDiQMcDfReMqZMrd8HfnVw77EJkMLM
L3PGQK/liiisgbHE2gcWNGJUj/TjLeyDF+3weReVifexct+V9CP8K9JD0cupxADW
S4r4qEvIzswnY2CXdkCQUg6Wt7rF4LRBum1yleJXvPeOqFgsm+YMtCwqWjnK2d/K
YHJXxcRFwUJWcpAwmIL4qzMO41VZEPfW0qSyPIoZ3FqMvUi+11VDn1QxEaczLTVH
dfLdFMxrUT56jdnQMeLlf1GjjSFvKOQkCPVQaZMWK6QIgPCX8BSHhRlIAKPbh9lX
UGjkOT8nVtAx+OzyGKJlJfTZvDrA2q5+m0+Qf4QrFaTVfKNMruayR7tj5qzwfzTJ
uIEoIIiJpipFZWomlSQ+bggNvaimuC/24/iCCdE/7JPdEuEo60NKtxvYuktcve0i
HRntLy/AQW2rHWmXTe8DarM1qnbwqxLTA7ysyYnKlEYreXkuRmpPr27qaMB8mczo
Z4dj0sYhTFnbELbRmEhoqSPIXwNf0h4Oo7tfTyNKWg6uh9yzMQYWINooInN+deFP
EJZ+3RKZOTCNwTVh3EV2878VjwLBMsnCO7MqqUwq7vK44nuKTZ/KXbZdvxSGi2Yn
32ikACOJ2DaKqJV6T9S2R7wIzfTvbMrjydg3H+Ow4+/K3teAIm1xy8GC/wU6C3hD
p8UQSOEyGOR5XHazcMU7pXc5GIRZtYlxnnj3+7iOxobHVHAsLCuo4WrXdLtbQ2I8
clv9jjc6wopwEBPAtY0A/BM/Wyv6xeuEwIU3lhxNNEXF5Yk/7FsyBLe1rK+Qphuu
rB9hGZIAqEbYGTtxr44oHGkUUz9IPJslGBohfDywRl721YNZSwj+9EqWMZQVTGCF
vOAqM8lKQFxfyF/aL8CcI+q/pFit6HhBO07PBuYDlOHQwP69jhDk/NhM2cHdas5U
pZo64lsz5j9uK2EKynhzdBbVzMOgqh3EEwfBbx3EMAwFtwwTE3LIK/uwc/o6dldp
0EqH98Kmyf1wVCrYSvXCO3W9qzSbU06SVwGujYaSIPGFO/WGVhq34Lr4WaRjHKkI
7j0wddS64xvfGmf/YI2sGSwPpo7A1C6ugh2LC+eOiHdIdtnHxQ3P+y1HR89cPmej
ZgzvUi9xA9kacChQtHTKUlW2gBAXfVuMDxzHnGAO3SSH40zh+rsQLh5fHTnKaH0t
Md11mTknCrkniaRjLzXdUc3vt3t5wOgXtisEl6+uLv2x6sRh9h4RsVOWYpAJQ8Ic
DBRlFKPCID5QjnXUwpXr5hEAIQJ2nKPWBneKtoMKuBsQ8M0N1p/C+/wXI7s6EmGP
xLigXv8QWPxZORIGjlG6bA8Fd5Tl4NvQDlQeGNWA5u3GhxlHin9E8jZ0Oldvm41f
2+BA0YERtvqxyjdA3IYuMXE/i1npCsU3sd9F+FVOKLmrlkwd0Q7wLpMlqxsFVxaA
wIoJOMTbZhw9v/Kr+G3C0BdJJj7edzg6MwGcAfGBB6O5aAfHod38rNimXRR3O4oN
bluvwNep/cbqtILhQ0DLLeLKChMRvK7qp2E01EA+G8M/CnJ6ChYuKggsrGRRmyu6
ocF+Sa1ZoazIQPAQeDPM0pyATzIsgsdXzTi1xj1WYDSz8vsa5hC1BOhknH/9ihdT
r6Mf3GGUHb1Cr9caBzjx7LTurV/1sFwrLSEr8qBZl5Tn7pmFjcVxmFwD73vmOMGn
AUkoYMYXHQq/99mCPypxy/AtViylP/qAtxLAsvh6jLn7vMCchUUn84IDVA1pHIRD
94BYLsEJy4WVRzrmAJYHStd/t7GryQvhO4lRu6L5P4pJfkBwQWLeRI2uxzoiC69o
6YgpF67tzKm0ndGmoJl+DPsgRYy7gvs+hVdwtdl0Z8e7KBw9k5PayD5Dj+qdEDqI
hQj7fJViI4MQ0zQBCXAGmUhUGfOSEJOdiVSMlZEprNmM0U5qHHSMxL6We3JXnbje
XxGr5moDbY+MZorx3EXLw3ArZcgB5dq/dOzoB3Gmrt8/HQsYcO/57wZsTqgIIwun
RgvIfgQ3hNQbqTGLlMc/9UTSM8d0Wp1HoZz+qqpVdsTIseQX/+IyBNQ4/KzhltdD
PytZN/byrRL5LXL7WXP0DBJ6FNecPgP3QLITBW2bt5lO1waf9I8aGxfOLu/kwk3Q
TyG+lEJXYK2xJW6dttBBQWJA7K5pVqx02Geij9HHcYslmenzPn0vTGPlBckNuIav
89qsAmS/rpOrTafC8UNJyQDXHO/kTHyb5vZVfNZPlSSS/U21Kln3URlyQJJmvl8A
voljE/hWJfnJ/zE9GveUuNYNWETLiTKyqBvtqMlOE39unkg4cBHf35Y3rSRqtKv8
IPpPwbnM63BxsN3epQZJ/hisUv/T17nT2Q7sh5PDXy5/nLXWRO++wg712PmZOQm/
caDveruDXY4mVBNPSGiONg+v/2JBEJtPPsF52SWqMoBpSzZYyM6IWqoVySslJ0xi
HlFD7nGkYEIl/svF0KdjDemgAWmRcFlRsKH+ppio1K/jPe4hzwfXxbGygyBDBc/b
rG1g1530+YHEuC00IPJ7Zelx2lgDA522D3Ch4QL4R8EwthABaqtM/cojHXUjNC2N
SzmQhI2kFoXMBun6MuEX5Im+GSWKj7xx8G4x2CQRRQ38v53D8UPhy6TuDyWZvxiK
YgSwK3TU5G/xvg34pkSw+7FytCHbOTwlLRxaUV2VIpelzDSWaoY3SOglH+UM6HrG
4ODW0PdhMAQYUdCh1RpZF5D3fbERdDOdaYobzQ7pl1JALZCW6d9Fd+J71TdU33af
sv7xc+kbRk84OHlK9nDygHfUzzj4a4KOBkh6vZhYsZYnPCVm3g9l2tWA2kQHZ8QM
sOFcmk2G9lqNFfKMWqjn1FhoFOK8RiH+PG8YYqmpni8/SCHUAcQKFRSOqgCCAAYZ
bJKcyK3E2GvRHgPdAI+91oCXNWgBJIXuWaRoN+8LmRFIczApF9ttTy/bJ0fz95l4
fcz8pXD9rG8eMZAqvCr9LS8Dgrgr19l+O1kgzIOEfEg9RM7vc5wy2/OzMUvG+Cn8
x+W8UecLcw2uGp/1/sZZNbL4VzgiNChZaN0/YOk1b4N+T/7p1HXJWDxlXk4YQesP
mgF6TWrKmrx4BMCJHn+L1sT8ARHsoIYI5cPOYE1c2beG7+7j/10sdQaWu8zUY3iA
bSSOnVVmcy04J+SibBxRPj9/HesXDQ5TN08dGGfB52/e12gXhfEPAcSpNzpSP6OR
kZyJmMVm+pL8Qfc3aJx27K0u4SjnxthJSe9O9LkEho85HYDIcWNAw2Ft20EsquQH
sCgqh6i/1fOma/CXYDW9cLQ6MGof1JlNP38vet7DiCGf3E/u4HsJXLZNX4mn3F1D
mC3K5qZ1SB6Sgx8RdUvHe9zgbf5eVPSztbWLjPCgQ/3uPWEStb9N5q7wcAxtTIq9
rC31Cg3Qbt9+dDN/IGTt2M/yfURmOPrU3koDuRALEvm3p9n1Lc38xSeXtYjSaNev
z9c8vqzGc5KYw6Ty8D3fc3TfY9/3UX7WGKheC0ZOt+DJyZoMs4kgfGuKg18s3XZm
qOvy+UZbpZAKrUAIsH67HxYREJOv09PrT7oB437181HyPDf7FtPlwe4GJQgAjpnq
UyHbB0UgEpcSnx5CJ6sczIizJInue5iyQ5kjFRlEKCEH3vrTgSw1UMKvx+583Loi
JAkvvlOKPlq9P/FnAVjtbEQXzZYY4A2vNogXtp/BnP/DMD2B/pltpT9WBGWKcifL
g6QerYybsN9+rp83/l4i2C7F1ZHLk0apNdev2ScJGZp6Tbzhb/xhyJ5UXtUsqgTO
bp5aWN/dq/PiWb6Bmd63X9Zc22BZ59Q9IbXrMesXoNvem/1NTcMC4yuwuvKE5hHh
oFYca2QicE/hZXNeWnEqIsMnoKpCL2bf7aYoCy33pcQmsDjT9Hz+0CBGrNAGa+xd
Ym4MKyU3Gzl+lhKz1sc+TqB27jYP4pbma7B/nVNXShtKw7qq0+ynkcYddJaFu4/k
UxtO2BWYMmNBCxAyiwtb/9wukxt/weURWROxNS67729LmTOUOCcCJsE70KujOAAh
R1B8+AtUEa0Ng+RePCfDBQmk8w2g9qXlvTV94mg0L5U92WB3ZLx5dBZTMgHYGHSa
0+vq18xlqccawUoEzenOnNPlXuiCH4499biXnhofNj8ktBvh7Ci2/tcWo6Eu4ZwK
Q4gd4Do4TV8RkBwg0bGbiMrUOkRj8lz06eHDsbofbdOBHe9gUtXUisFs8pcXEAUi
p+LbHeV6fIXPMi7E/aMOK0Cp0cmfaRg67JrY4knny5eBQTJiv/DlPTLK/Rp/9wzW
Iht4YK88x1V4jzE0dH8ef36+UIhpu3ZF6eBpc0OryW1nrsVm5AMHXkNF4KHdZt7V
RQrrMKe3aWM38yFuOfZsAaxD/+zghWohrwzdj3DUquN56vIaytEXiBCP7wDCVLuV
L91Gk+AAbh1F7jSAnBeO9oMzcDMTbIz+2tMW+mQmdCU6u+nOogBRVABHeJYuLYfp
FICzCWCgrOX9X4kQ/t/rGDKiMKqWQun4us+8rMG3kwGnMqgGdHHGt7M9UCOhp12E
hKc1A3+oJEExpbN0sRLn/CxlrjwWdEbFWs3E/Asb97XCxGerzuHThnuDNQakbsE5
HpnhX0kVgZkdAUM4ySCFCFoxmyRlzHC8LanMIRaUv5XJIx90pegfAYUjmIu1Zmg1
4WB5SWBTKFIQSe3QkYfKcyanNC7VnohBGjiXbzCxc9+Ot8DKlD6k1tAWeXKNp9Tj
v7YIK4JIpzTwhBPDO1IedLA3Yxlw9WzIizv6B+9Ef+2VoDpbRAFU2WjuqXAhdwx7
TGsRSzYD4xzadcUwMcmR+mfozlXfkCvmFp30QtrqAIHkJ2xWf1w0z6B4x/RZDWqL
5RPs8BLp6giR+FnSshI3Knp126qxTmyAdSvao7NcLDVTYOE1iU83E7MMZMy1AjtI
1C9Nmoc1YbZnrFh/B9twkf89NyTie9KXwQIP3wTSA1zB7MbhQgALOv8pAwKOSAeX
61Ng8tCoI/XMVKlJbIxCZ+dnuk6heixqSQa8mvz3CK6jJcPqfhbhVp+C8elHNIRs
Y53g301D7t5BU7eFxJLZy9WR/n00XhaJLC+W2ixWpXdmGEpyXjMBvVeRvb6treKO
DVk7kGecPA8xR3upoN/H8d9mRkjELjT/32uJyf2wOl2iHwEUpRtTI0zHrjPWcupl
cF4EAmr4ircNbXKn9jaKDx9TWzp40FK2OVIucrfp/M6Ck9Ig2oG24zZ8u2GQbS9P
zk16EQvDdJvyyUdIPmSTXVa/03tvXgipGW7aZ1PgakWnpFh3fSmkQQCoLWYbKr1A
13DdxeW6os7zaMk0zENQ5g4eBUm8KiOoxeGc6EfGF9tfClsOlR7aPwVlaNjh2a/j
FlAavDRj/hw5ZgnGb5S86Qh/Ot1EKKXfEg8BGnI5hXv6TlMN9iCCiARe1qZjN3uO
5m6PxKe3wTsSBZkToQCCmrzNWPQ1tt1h+f/WF4PPFcC7yzNn3V5w4pxmp46Sqayo
Twlq084uYHa2INNo7Xru4YIUpE8zbad9pEb2lxjzOJM/nhth5AvQ6iu34mWiMYPy
PBovoqqD44wAhig1TpFggbi3TfzMx8GW6g8NbZDTvYDXtjTX/nKMb8RBScEQV+ff
LircnVsv4+vxDqEgkieB8aEflT8Uhe4aQokMn3jWsGkS9umrPNVxnH3FJsGgyFDk
mmYcWWaPW5wG01knFyicLZ/kRfUZy11wmYumDd13QEl9waD7zTmC053UgOf7+r4+
Okya4or2zjVxRMCprPTrHfOrnYulNzUIdhLZa/teyOEJ3fet2VQhOgvCWt1oIzaw
TyJkGpJw3fkgjfqf8kxihjRQ86GDPpKnS9qn3/hezztgz5Gt/TgBPG3CXNKCuXXx
x0w08IWeD06SA+hHM+tTNgMc1SIH1yXf6OYdSuLgdDmHsV4KTJD8P0ne2H4tHvHM
hYFar0uPl0v6wU4nmwcJnTr7UcZ30XCXuUWCJJaSvSMlymPstKCleELIcB7/pvVJ
mHOQ9+ehKWlPIN3ozmGxv67iRHlf+Y3hOiavgpPyTlkk1FxkBhgibqTRQxuNDKpt
fH2gFTyNyUWpkyMRtgt8oLD1IgdG8QiNOAadvJV591f1ZvtSw4Bfnx+wu2YuqVDe
Sml9U1KQv++TFxBt8cQp2IrR+Jzg+0AmAxc5O9ES/27fBulWNpCuDsCIQbApX6Sf
DL423vfatjx7/paQrzxLCF6KZJrZX4AsqzRokCvIl7SM0Xz8KVnuuiXxU3IzoQyT
se3n9x48QyuM4rub8oT3lZUUkTueG8D9ha3EA6g38D2l2zrRNbU9fkYv1/pHwquA
d/G+QHMedyENWmkSo3lCLPgbqIqOZjrp7PHXxed8kBmZZ3PMoxv4qTDpLvpjoMNV
KXI8WfzlYLaNtpm69b3aLZQnmnWCzvHMo8NGhJ8prFhx8CYqp7KUsriHgi2UzRa+
h1fbRMVYy3uXweib6OWeaWNVF4wHzdIZXUzFUHcnNSn4vYth/boUpp3+MGoGCfX4
kuQxLCBP9jnIAJalC7DPW7ltDIHddLeXhKpitXDbBdZtdwncWlk0boGdmRVCgaB0
L5e4zuzzrozk4qZr8eAaJvZQvWetGeU2QsrmyGtJW5htIkPgOwfWBVD8eIGVO3qE
h+aqA84Bie2CYscumlodFRXg/Hh3raExBuqV2jkTu9S/w1o7GRui3Fsyzq1ZCg0Q
h+18jfe5OpllukB9wcOk3JCbKtNWcIF9gnzrrpQI2BQ/l7T4QZBVeQIy5yEaU9uB
RG7voPsjaalp3gQe9f+8YEJVLoofrBo4VU65QEHM+2ahau6z1URCJ/zJmNp54i3g
7pW6QVMTXlIizz+ljANsbEQ2kUvTSb78ycY2kFyfB+U0outIrIS58Zudp5RlmmLY
xUG5oyI0323a/it1XOCJjZYk9nVTT8lD3bz1fMx94agRuOO+t0gRSyYsIzwamhmf
Frt4Vct7fqHvvkYP2E56g8+Tybf7DvUeTGSz2n3oLfuyui7Ze7o6a+6X+oW4y6Ag
Mw2PQjisvsMfF3KrCL/GsZ9/4t1KvdgXXNwcoH0w8o38Ibm1nlj2xm8dYB4YZeFi
qcHqNNtCM3/RolMmt0hMt/tOB6379v3pBBcWuoyuFG+UnOKZQRFCTkLEtcImULG8
sQywmoJOdUIGn6ybHhiZEFUEBKCg5c1ud1+IGjQS5G7dTJl3RwNcSwT9usbjH7oQ
Y6xT86nxf5NpyZaS1ohfs5Bk7+y+psoiy3CwW8jG7+4xaMe1D6bYQPhhTXzMb6NF
kDAvWrw3X7+w+sWrtO9gmc4AkZbneCYTscPV+IJn9eWwxyG80Ex7xmxonISYKLGf
yCg5XALAD0uV4wIUWzyytO90IFldSHdbMiI36doO/G23YoXaHDgNyIMvwdBRmPoR
L8BYyjscV2BFKG5QvHd7l7Ni2fcR2W/jEI3FnfTE+z3xMF5wv2bXndVP9cpNwKxB
zsdwjZEfGlrV+AyVLJaoHAtTsObxRpqULvTHE2Auztrc61YfF7tiw60kPkub00AI
j+mwovkcL5EMnRcpNxllYP9OKbwtZRIVWoize5loSJrpdvUlgv42IvOThq/mzcR1
z5w9u94g77JSI/q2tmvoS5RFwCnem7rxybM7Ui99XmZLANdMYuIcyX5m2KTu/kh+
3cUYOQzHfu9NvbqIYG2v5jnRoAUffAQasZoKc9ohctJx6TXHjGZyT9lLugbt8IgH
re2s+yiBCgt85kEf+alophesaUPJ4dtCTKFohYapwnT0gEjlq9wjTzharphvhCI7
Fexfz6b6nSJ9XMbfHU4XsGNiMkZlvlyyIbS7PpfoZHquidZQ3MfHiNBtD6w8tD1d
Rcp8+8a5GtuLNlNp0yNhQMIRlDQR47/gOoSybpOZn+CcqlCZtaR3Z8dSmpahj6jp
OIPks/UZRZxRVAyDBoqgSV5dn+sBvxgDLGEd9l+X7UZkh8XD144PUjE+qo3rs1OL
2hlGoUzza6+zHsm4F2E/SEaN0v8fpejGYN9Onsc2/ex77ghMjfHonQb11mfy0Zjv
zWuua3bEC18Ts/J/drbvzNgaGerEyit/W2fszvCOqwBB0HWKPh9NTolhyurG6yqq
+S4wfqeEkHE6dCB1Ds6yQLUuX+q8Ka1uaI9oIlfJhigKP2q4+Z7Z2flZiL/kE2X1
2ZUqvg2FyN1ywYWKbWroUWuCywsDI4OWylSp5giZBbBSLJMknqKPgK+qTeF0rN0T
7wJWb+zhevRTS+Hn9I4ebh/5GUNFAlnIE1mXtJS0gP2QUgBakzKnGkSgxFXSOcXT
/nc4tuVPM/clZSzeiS40l/ZOXRs4fcsYG7FCh30es6jfCLf+RDDvWoWPI3fDaAF4
Qc75tQB/WutDqxwxf4K5QSsCBCy2QlJijrm1VikTQZzpCBZCYPuwyDYtzSnmb+bc
jjQZljLFLrq3yQuiNJgGx7ohgZXJ6SIQKEmBBfwPmZYvU9u6S3zy1W2VMPrxLwUt
j5aJ+dZBzvsF/2F4tkdYbK9BoEd7oIpblJ0+1+MV8UnWRIB5oOcio/NmhYYz6W3S
IyH6Cl2ydI0QvSEbfMewR5QTLLaE4wYuTvtW1ZI2iDSXlArnd+Ty7qGsZNMfSv5F
WvIafPphj8GY6tyfv23yyB2dyNFq6ng3J8fQgfGNLu7TlM4eZxAoIKWGKtdy3Js7
8aFU9JvN3mfanwJ4rPlglfF25GigSSQiuICYKA527V4JZc8yT78sRMDUqFf08sDr
FsS5FDVujjITgaZobWx/q45cergbPefFSOb4hLFU+FMIG1oORlAnmHvVDp6iGViI
PgGx/5uk4C7GfoyBqZm0QKdu1d5jfc62NrfiUwQTCfQKLNs+LdnlJKSSOUu27rFF
xdaj00SRQhHgaZhSD6fv64R5qQSeO4lGZN/Efr6wkhpjpoz6m7hjD5pJlVLOkSx3
Gef3Qmti/qdbEAVOWo+CTSiYFLnV3gnArh9Jsta+0zP4gvL/s1x9L4L+jkqXAWe7
c+dB5biNL6HnAr4YXfpAZBtS52Qv2ZiM26qe0seiMfjRBr9+ZuJ96YxNXH/VXpgb
aee5LcMiM/ufFkzZxUvvU5/wTxo/DP3JBKtCDsFG9mc3M/M5hwCw+IegYs3zLeTF
XBkGMAsVgB61mMBLZeDGTXNvz49oaRfZ2lI398r0nIzmTyqpql5QajEZeAQ+NaKx
0G1WrVTudYoZllDgAxP+rCzfKiT5ecaJade569BK6FmFDpRex3DgQZZpiSLyfIoi
4uEH2DOBdQjriQs+SpluaChAs5zlbfiCKWCVy5gU/JGclKmTPeT/leG5forqEPcl
pyemn9B8iV+DQ7BLTvjjL+rGz+mztX/ug3jz/SGHnMIvGG9xF8CSSSrLuzL01Xiw
BSwKPCdiRMwc4WqAGd5vyb44/m0G1fHO92zphk3HXG8tuw55i5Q+Lr18cqkbnRv0
HBI7W40RB0XZnXOl8LFydX3c9/FGm7F/LCq7riG3tx1BZvOSQnNOjr0TfJtCiUDI
R6ILv12Y3JpPSmZrCMC4p4XeG64/yvbaR1riPvkUd/pDZZTL0pn8ofPTM8y3pcvo
SlfsRkkfhgXy9wXyYGOzZd3YYXGaOsspQCqkBY94yP35rZr/gafXYy74YwAWj433
GKlAaByNUgSZWocyiS4tNUytSbJjTN5WlBW9gXeOcSpbQyxRMJsqgBNOdGrTXv2/
sPd2kvL/+8q5IDP3PoYqJnCCYUbJotocLjxqiSeOHLQzz6fXDWxuL9glHBP+iJ72
+ysdaki8UXenYrDiS49y9S5/z0W4L+Fk8RT/rPrcXLgyNGuXqw3+ImULUf1kHQYl
re6vTGBij/V6Zmm4qduYVFumSeOz1xdBQc50yp4tNskwtLkndL58iGspX4u5c04x
//BmJEg2hIaO4lA3xDpJ3BY4sDiBf7w1UaPD7cJwqVGbyw0PVue7BRmoGdZXo8sd
AGfD6smYjCobDml51gD5IZQxpnScypBApTK/6UEUFS/Po35MUFMxCUU9/jv9614r
WjBdAXDQAWIPfaDOHsMgi1CLOaIbrl/+VqkdASzn5eLJNj6dak332jlmU4NQY1Km
yeJX4mGWUnuF5YqGCh7QyGn3SnHeGTRaPTROgQ8Vk4TXsaWsZGc0RxCOuG9QLZD4
eHWYJKNc9wNnjbtG8IZ+CH7WUc1DcPnOQmRj0NTnsnbHJ8VKBJDG3KXwpws1UiZn
kP75xE/5DPBdU3gWzJw22TU2bUxhlRKZ+TVyvB53D4vJK3KhiUnio1HAfIycsWc/
bBlWp8IfoXnN4Er/3O8oEGaXzK0DiR3WhS8XFd7zAmuO7GsqgXVkOk8fGiDJ6++a
vPmVD6NOhaLaRCk2TN7fmUd3IbAOP4E/kjv6JcCxmEINGZYYeJOy3XYIyJ2pG23x
4h9rXBL3Qm4HqxGpw1o68jwte5ltLn87UHkb4kseLiRb0SLx+Hy81GOY5a2y4pny
yAo0Zi8Jsn0ap4nRB088VvCXVIsj0pUKjVsgz9MUzClMO4hfcT1I6Qy30o5nYaus
aMBd6lFzZhC4oGIGUisHAQmiFMw8n48tsIk/elMLkYwht0PUYQpYjocOqvw5oun5
8cMhFHiFn1KiBMDSXvLWC6i2TJ4VPEI40LOBV4qfn1Z/eNew0kF1ZVh+wguBDkh/
7U4cuBmJEKjFsTR2yxnx3x3HsPY+zNjIVb+pJFIqwjL/2qq5bsWD7v/JqgNzA+V3
4m5tk50cRJiVxewm38poEdxMCH6KcIO83rxxQRvyLlT4ERgo5B1KaOGtCr+QAZ6T
IJXo5XZwerrLwCe/AUbhoSRceBZ/FUVi3SO1e4BR0zghs8wDg+P0ezX7TIN7Jjtr
oN2lWvYeosUrZGfsIFslcVsTDAnIkofxgT+13/3WwTZHXJRFpGk4WwhNn6Uw4WTw
SB/p8M4sA5Z1en/FlOT9JQvEjcNMtzZt9OCGQ9jc7REmOWAiAXQ4mp1mLqCzSHLv
IFAOIV5BeVyMs9QqLO6TemoX4DnGV7Pi4SktJI5Fy30PeVGv5aZp52QrVzBIE0qT
CLXarUyR2SFBtAv1o6DDGsYYsTJKGXJTFBaxZPZfFG41ELlVOQhNxsY2Lwgsymnr
xnXs5TJFRufLWDjSUVo944l/GsM2T0O+uoCabxwXhZCtuooSzUcOWx/INqWUHaAy
wwCnCH0GrbIAbH6gfD43CJjdp8UKxEhkM0s4IL/+mmTBd7QMxsDRrQicUOg5j/z5
ejn/zLmmzqBCGXxiMCG8sqb38+6Ulkn4IPdQkfjBoV8zVgED+f+gezE1YGIUtPMz
bzC3IbA4zRe+EOJTpO75w3mWUl/xJkIjSbZiZ4Jkq2WmJ9fqt0TLL2xvjjcX7bp9
7Kqx8X15c/1Vu3LbNRt96XyPRaOjDKbB3KM5tNfyVJPwvc6SYJ5QE5lTe6kS9AzK
02M/5y2DdLmd4dR2qcIziqoLhRX6FS8Jy6lsWk2Gufx35Ig0Z8kxk+ZIVaUdeAvl
4EYmKhyAAsE/2fi0m+65zGKVm/GsRkiF3s354PPf/zSdW7Ysol5ACMKM4MK7AP2y
8bQ7kBLahy+0tKtEiGOm8h2ItvoOIbdEQ59bkpvEkc4uwtgVNWH/5sMHhbWAKMkv
y7A2uAu0Pm4GTRuTglbz/NXO8KHbarXqEhPRceW+WUjiqMG+1nHbldUpZCKkufU4
oecxKKd+Me4h5/ljR4wwcuvmQCsSD39mFjfMPFc1Fdut/CHCopvsJGeUlhZYsJt7
jLE1ewRhRybwhD6zzmYwYk7pbGVA90sr2WTGyPhsz0iGkHxfMxXCQnwTocwQLtdW
PvU8MT61ZmRXPliQWTO0yHhD2mVpl8aFAXixI+rIcaaY0AGPkVW5RYLqwQTkOhj/
TyTp7QZLqpjv8ZiyqGQBmOsszlsmEpID1Qr78n8I/MjN63Itj1nWjM3sNq/f/LVC
nNE4z8vzT1CBbOItjoEuEoRZdo8JZ0io0e987DS+riQxwamIBX6fN7GHaPw1L6RP
vbpQgbuzEIjqHWBMhMZ3RRU831A1zEh6B620ICgQKUQRy0kQLt0grzRMP+obMDkE
9XIlH2CMaiNA2GH/y7u803gIQJ27DLyWS4AxxEQQsOGBFROESmjhIvKS2yxZ9sBr
UAtacza65TPNUcVsLydsGb5sKIdWpljSzxtPF5t9DVMQRt1J0++BfADKxei4CXMU
EkeGd9LWkv5npPCk9JCD53fd1wjAnZT7Ge09JHhMG7qpbgs+8Pd3OFdKQFSurHsI
NVK5nLRKGsVKi0ja0NwT5csfsnHIU3KcYPSxU3TZOPBgxE6zPKAfKKRlynWGCCLv
Q37Dy6HwpIu7BrrWRIHELs2eoA6xHf41uCxM97Z09nCqDGVZFX6Pioj86XN/i8gY
eb4JKLuBvG2TiVEyz27fOAg9+rVY/8v18sl2Spj+TdeprY0z81WNH/pdBAN/7fLd
IYKX5hjJKoG78MBNtSlIXhd6YGAjF9/6YzYzyD20987u6k7Mh4dFE836cfWUy6Jz
WZ0RA6mpsEygbNuQuEOOO5O03mL7Ip00+xFdzUrfOUNE/kBStEV8UYPWDJjzWvb2
Rmg2zJr4PjB+qGb9b5yWZLtvUEPzlpV68oTKWjcrmb1z2tDpCKEiSS4ZhDr5k6VD
syCVxYED6yF55vxErUyAOccuu043CJK9G7zJT5wnBRSbPMRHm4L7U3xrhmS6B1cm
3o5q/QKLgS1gjutQToABP9hGfrJYL0407wr1bcClcKEz3SdcgS8B4V7wr81TgjSM
gl4TXZn1VfO432l8GiCZOCZANnhT2Zy6Co41Y2NaUjFTht7VlaXboXJI/4qYfINP
lA7/BwKy4QjsjFYMk9LkHGQ9aoCllmW70nfOsz2ddbV9C6rmJ+4rb7Luo68z/LxG
tYRXifpu5rk+Y+tWgxrEDYFxi7ZSR7HDdQ8Chmq+LBRxoKcUfv+eT0Mbd6E1ieUC
A4HHaje0lNdmskx0wzV1XG5xQR5mnVLscZNhwNVyPg2ifTOhU1TwWjZdgjZKxJUH
1GGOFIeqYcWsUWvveOUakppLHRp+ul2P+R92UixO2TGimCwQ1wbT/ZQdO5dSlwUf
6CCdKMZ5/iLb9BCEd90eUp51dJu05y0N1V0n3oWsgJEEgAhTN0roMiNfc2wHtLWD
JikWYF3ni0CFlGfTMu/mKTd4ox33K+Y5KBAk/2YW/qe6jtEzMDHN33W3e36IBmoa
0Bumn5Kg1WV2gHLTkosGLIB0J3KeNKPM1hEcSH+zfJL+5suOIgzcyTDQkCc2kY2R
tVxizizZZF/VSy5TfXhIRMVVPnGVHe5mQuyhV9t62U9jI4lrM0dznPYpx8Ajoi76
ggc8sUPZbXqdpQ/WOB5OZXbr+D6NtC00fVAFevi/XhvCRN8MhN0gTps2VtYPPZ5z
k61wQpcJEt4DRvSsA4dDtmqMt6NL+ACbMJmVzT+9KRFcJK7kO7DCJgt0n1JNltoP
+6sDlikdU5wnFOpk/0OtkSrZugzFfn4am2aklvkrIQI5JBGg0SQuG3BLQDFbDT2P
3GvfjcSReOFWjm8VkZCCuSZjQy+q6hrzMVT/pultzF8yeIVvvyH5HWxhro4rwwk5
UU94Kdwzrs+YQkIyyfRTZCUVhnKsZfy9HWRsO2fSuCP01+AoNkwwgpo8ytAkg+XM
RSu5r1mIUtqtpiYKLdGy1ZUVSUC0DfKUVGCQ1KFKFEAiZuilAyDgbeN6eyw3xzT2
FhqY0ADBV4Dc8sc+cgOE+GvTl1QHU3cJEuefwv9rfDvrIUlKd+iQqwm7VIwNKW7m
T98HMPkWc9IqI6B9rjXhJrxdSiNH3JZPVBjICWdvZSLVMYULBmhYRXKhcgMdRlw5
9loW20eSWaockLCD1ZM+CMsu+C3N78NdUpVC8SR0GO/cXZLKv7tsmTH0Hfv6U7pN
sUPeTL9uuSWMs6zH3bsYwbMvahhoY17nxmBJC/9XRCPC6EgwZPoel7kBGM4CVa91
bBEVUyxL+sTFa2zO/ubuYDuI6nsVLYS4IocUCy/qoUcHmZAYQznST3LKvmmREzDX
VgMpPnnG0YcJtN8wwRnHTtSI/uEyCauwqPYx1G0EQ3VFd5If9a+joIB2jgPWkKef
kSatqVemRYj2R5i9ZLs0Geulw8duJ8razaqttFhz5p6PbYHAoq8mpuoTJdGu7G/H
Z3sXLyMktqYRKwHh8T9078bhDoYwmYStDl5XjlmDDideBPwCdcweVFuF6y/coyRF
d5QysHEhOvc4hRS2302ZX4OemNVVsdsIEbxcFjmW1dW6vbZfK03g7WlaIyGX+Q8l
9pgko4d6dY4P+m07oQbYFjfl6a4cELjYdm1Cqrz99jvdRM/XuXSZJWaW2XtlOoix
Z2K//3K/xzMGiz5gHlx03uUkGZKeNAZuLwJe0Oob2xd9xFtKGJkS1QpQA2oLw3kG
6AjE9drqPTYfVeDAKQblLSndIWb1TlWp85qxzGteFGmDb/9AGWQ/rPREqCrFrfMw
HnXp+i/+TnwWnNhtnyYt/cLz/mJLTw50BdNVVIDZyK0lI6dY6Nv3A7+V5jOYlfM1
cF9Klozca8wtqwRfwTypZenDQfp5WboehSTFKdnSpujOqIcpzX7+7IVfKaIEDNVZ
CxmYCZBmGVjRmVWqMlFIez2cJk/Z6ozo5mpmGyAQeCOKWD7y5k39pPqed+Edy4t2
+WgR1mn+8xw35jb8SZVUOnYO+DBUGU0xr3L9dR5ADvwvxy3NfWD8hruINueeZz9V
HWJzylPP8NsexuCVizapNLzVpytdHhiPQaKWDCGXh/8C7IqDrRjkGWpkcAuYhyuC
qx4Sy2dHggrOh/ZydYwC4LJDCPb9iAVcXXjTAYhhjLJS5tH7GgioEn/rkapBAAUM
hsZVfRFCjx02b54efbP7Jbxl0tRsLEiV8542T8ezHbY6mje9eCUsXusugyxgPeUa
uYqmljvOmtjORebJTNigJ9udTJriY8jh3vlXiPBe8200zYUyYNW9ttIsPOBGCFK2
TzRP8/+IqJySVdmM+2SuWJzgHj76G6NOSIPVV9Xf/zPCwUcTF4Qo9nAm6jGGFE4Q
al1STVrMQByi+MxHhjXqi4Vaq+rSBABW7km/9yR2kxrYh3kqqxtTZddcr65yNPWs
q9VNuOLRmahyS3R4qcD0OM5IYSuKm/ZMf6J4fXQVJSwSUV2ZxQEgYh72F1dkLF3E
mKflf80ySgF24jspaorgT2z6z9GBY0bPlK4GvCGYWBXvsp2236NOCB2+US3YdSQX
7vsu5wH1/5hDcTxk35wCmbWJioZEno7ByERK51vfddbQERivaIn1Mdlou0YsDAA/
bFa0Lc4vgh66s/uiXbgiMyo4cTckiiMcGacDS19Ped7F9jqdj7UBK/Vln5uzduCx
X2ht+dpSDQH00I6MZ1gkZqeoMdHMqq4VJUDi4q/2n2cTU3Y/mTTC4kZEqsghZBc/
HZ1NOnrYjoVkKRS53miarxpg6fIVc7Q47llTrH3xLQSirlFtai8tH+y2/9Bzutle
Wa3exTNettxGBSqoU1TZtgdF6Sk3WtpZUcVGazkfuoAxNgFEDCOZIiIeHCu4tDUe
H8fzmJajWxK/uSNOmV+ww7a35kUiiXyrMibCcggeFAOt+I3eGNBYvBas5gpmOOWU
tfbrr5mOtF4bkAkJT1ABDOg/YY+1LaZCz5wazoEgzls3+xseT/KDivAsFN07Ul8I
gAT7hkh763bGJlh4i0Fq69wCokLbIgCxyRzWTwZKXab5jdXLAAa2fWNCxgLUWyXy
ggmkBNTaWoM4rr30+PCWWe9jjq4S8mTxbz8H8k8jwyldkQ/HAPbSlaSgSvnY7Ake
idwJVq/YcLb9dfbJBybXqFNwfGoyQN3yBZRlsSnTaZ09wyg5H1CZJ/CrGzLaip8Z
rcQ8eRCppo43T9bYssZdxy1taRscuj85gPVav06+dgaXY2UQfYwcmRi7HNIAJTXz
CGptjeTffHCZgNFJaig91kc8pQY+E79uY8yewQfY3BHMefjRJoR+zlKve2Ah/nle
nKmuY8LxBiChuuCzafU+9+QrxpQmZmbRssStxkEMd7C7eaiRhoiL4dPD+WnrcG4S
hnoiOfKDNKyMWf7czzPcM7Y5Q0epJobHY2D2nxMuQFjFsApdBy18FTzh8hzMx+0b
tglFqg0qMPfKxV+oJlZR55FMpfITPpXuMkzZ7IoruAtDfNzCzBeogqiRsIX5V43U
xMRGMphgTeizIA9kT1p0qUX/RO3VLGNEPUh9tiy/5qtN7gXXwhkl5sAYQW/8cbMT
nK0KQcFsd3imnMYaqCuZ3HZugCTRKuPDF0SPEQlfTO3nU9GBq5a3yrjzVCJNM93u
Tv0OnYkWMzedFI1UonE725dTdcjrPEk8pvk4c/OmimKOnCcwXqY/dXTMT+bi2YrE
zAa1lowYUd0xsEI17WdeAzX7VqjR7XRUC3nZ2j9M0DTiNH9Cfdg5TAxvEI6085VY
KBKAPbr9f+9w6KqeeC3k7RJN0ebqDLJt/lLgbH4S2n5ZJO2M/+WqX5sp+4OwA6Q/
W/es815i8eafPC8Li1awiOgC+EQfudyFq/qMqtBodl1jNb62+gXqutpqqpp9ndqI
7MwHLhyodSFhwCF+jiV/H40y9HSVai9+T8V6AYPTuORL8ZN26XYVZq9lDSSK6j7Z
WAt+g3XrJFCMeT8YFCKviFQn73J+rvnir+9UgaOLjIt8GJxNcGsSOx5Fw8cBv7Mo
vcSA6iBL4bXkiJTP6CWdgEl7T/o89VDLvJjX2iuGBH6TpkV9rsOFBA/+uSkwRVbB
AyfklDmKpb/QifC0FljE0nkKuvTLT8beMKREax6GffaW0mCBJoYk7c9DoYZnjXfZ
u1vf4AhqMS67BsN5r1FIw3/xR39xc3ts1rkK5joh6UIBJIrtdW3FToS4TyHXLKHB
7Vak9QhxMhd4zoSHSWaInr/B0PB7fJxZ+8TkkuSsf6YroIfsRxT3kSR0jO0nT2tD
FCYAKi20Cp/iQ47Y0qU5/yzwdutsMT4smVhTIiOD50fCGDpESDsBhHCBd566ytzv
RLH0HZuZGvOr596UL0O/X1CtvI+m5FJbnl217m09srhB0qyz4IGRlDAXvfs2WRix
mhKg0SXBuS8CdmtchgfyGwZo6WF+4L4CYIvHDBuVjM42L3MxRzpcJ4RLgqGfbEoL
EI5dVd+fH23m+1Ttjqk2tbX6KUNMhnprCQkkeQl37uQil4KxC/BUR4nQyVBolUcH
FGx5U7PeJDX+zjKa4azlBIQRhVyYnQWV/klboZXW2Ay9kOaU1d7FAssvQR8sNiEg
DsZYYpILtrqoSzWU0ahGDBtVOC2T3GadO5DWPVrv87KVEnAzeRIK+JBQVueK5ILx
mngAcnLsiwWx2D+pK0v0qXEwoPsxIovQIW8y5GrYyG98aE2aCy8ihFeQ+Xl9XH07
Qm7YmITqZXI74d6ABEFr9L0b/jN6DKIrTLCHNl/x32GBzLIsFdjgoEfJWWEFjpeg
l+tYFPY8ZqRQ9KSm+CbBTbDEKw+h34VjjJDLFphTj7TxDrT+vzw4eaCdYaRII4ke
bLzQEokIAYIWCF0ditVGEoQIUL7Ccwx9jnVnxGqkPCZfUeuxKS456WtQnxATLlmF
S1fXK4GwhGckiN1ztdJmQwDToFNhjB88SB4FGaBTEIM+MW/F6bzRZe+YpMwPKZ0g
JSxkgfkqOM4V33zehxmQjIeHgc0WwRJ+YKKufmRhMBPnBRTmr43bIttjdt0I791E
UKKOmdJFml9mg5DxOEMNYk6MIHk/hrHT5pT8VKynw+q4/vqitJxkPURaCXb/BNR9
SCAs6pN3o+X0yKxmKKG3jwD28AxUCwehUXbAERKKdj2pvVdFZB3ZkiXUmwyM4I1z
qfssAuCDCo5dHbFlD37tTOydH7CjGvCZFkLpYjq/JRKlUG+T1GDDtz1YW+vqEcVJ
oiAxnELci/9+2z/lG/qxzwfq9uvk5z1KQcy5IAuYViFY8xDSv/hokit+YsvZQoZ+
UQO+aw4TfZxc0/T2N/zbsz5B72F8mSIvfgF3pM09wpStpg+4qSH50258/sM+gwsy
xDco4fH0SJWGom0SZ8+BQcBhXWUFiyfy9fi9jpVjGJiatlNQXHxB7hplKEoDaEmh
Up3RsnY7+7L2KIMGK7ecPH9eFlbhTQGOwMRiMIk30JRjn2uVMDyYF4JZc51gx1G9
pNhCTP1lF3YDm0M/LJqVJGHkXQ4+b55nV+2wKv8SZs3jqyJiumaju/2i/+VYbd3l
eSZq19OzAgBPiIxDK7/G0Yp8IXYU23BtuqjrlqhdMBwVadzttdnyt+iClmfhpI7a
WARS03eGg+BP8VOgHY1LRK12oC3xmYMVQnkpBpyEZujRb3ePIpufM3T4cB25osS3
Q2RnEy/m2tBKtdlyq+9UHJwVGw/zm1V/SkvDpQ7m5UQcUk53Ggun5t8n/JXPGDjh
110bxvXYEi0pg3+jabRzvDRT4X+2dQ7/+Ti1tE5IsQDD6TLxVj+inYb8KwkPnhtp
wbNIM63xEH29bcSVPTK0Nswsv2LhvGVu9sg/VGGALBkxsLC+nR8/+kMl0TY7kZOM
9nIzJVV5J7gBTZtIfU/BRR/pQ1MsD86e1pj5DnIRG45oaIz0D++M+/re6+93Mvbj
YDKwnuQjFBVi05e2s6D3YSc3lDW2xvuuJuPqhMF346XO8kdRJjOd0FYhP/ZrRHKc
q0nVzjfdVWBr8+6fDc+BiQxGVsHoO4SpfNyq1o1vZ5oUtBlMs3wFnbLyat//VhqI
xCNydr1yxNSSSxrEUhOVFXbpPNlH/5hbX9d4jMxxpWYYDNZOUyVIkvUcTGOm3m03
8ShhcuqRIPxvZCd2VlSfE4Gtz52EvLnYKCx1ePI0hNKxmZGonpr/X7c6n1B1K2oA
pn1x5Js0OA16mPLlibqLIaK7h2Bmu792HR0h5xSzhp1vpRipg98giwGieiQnCBRL
N0vONa/szj6QZRcRos9ZYTnyfjzi5Tnmej+eIAym5AQzOgmPhh2xvHKmmKHv6zIt
y703mgPngxRXjJ/ks7JoFrJN49ddvEgEU+/3/uHaS5bU4nDQg5X59MiKhwwmKv8v
fZJWVQ+TNHrsK7N5d2SIayvHVFVAftC5nOxjVoXVXnyC3pYbL3qwEFNcorQXowPb
A/Rf/z4wWHra5s3rfU0GCTb83JalBHd8tUu8TrVQKOg7a9kaojCtbAJdaJ01EtQm
oTC641bAwEFQ0G6SUmbo/s5BUjRtGiDsAeFhlst8Wf8U0KfCXN8o+UlrcOlfhpK/
eFl9sxihEIzh8MQL2EQQIL8+GP2QaSeZvkPCi/pPxVyw85p+OLQmueppbyx6+Fb2
AdKy1/H9EQ6qCwOzeHflyWG6OChtaYpzlOb64RWyjYczCxx+1uJuSiyquDClIkdO
Xi+5HaYd8sCr/n1YqNv6MBJzaJK/KPmJB6wWattg0Qfinuis1Kmwf75wZEa8N1Ls
hu9lUz/TPz0ugdvCJq3E27UjbuYHo+O3SIzObaBHrp8kuJXHZbmVC7CI265Ausij
qug/sHwBE6Nv58TKZa0PMGTMEtMzCBlEpVLkzUsf/GjOLaOOugcR0vWAQbH5FdsB
crMPrevkrmNqtGTvO+fHczAceu3fN+zcAvaoJn/CqTJzBqLD17bBvvFuBA0B/skj
3liXw1oAegY1K0vAcARQxSVCqXaA9u+C2CSC5Bzj3pFyblILu3fX6gmUehFdrxR/
ukeZLkjXSuLBmE+U7FksI+jwK/ttEDWWJaqOD+ZWS5O2vUaJxYnelCvf5EA/iSM3
orT3Ezsa7ZiohOSfJxYgP3Pm9sXv/q6o/jImk1AyV48b3SwT9vr9cxHUmfKR6ciQ
h6xeRpdmUehAPWQ/W5AmmO4KGiTVFcAK4y+9E6ROhS79d3ZevaHlE/i49BOpNtV2
Mvd4g2J3UXCVlXzjn0bJOh7oO/c0xNiYA5uWsggtfe6Fys3oHR1iICRfr357OxPA
RlKSE0ltEqiutT+noJECijVckAcITJpGXgMcAaYTpHYLUpbCQ3BwchcgnY+fJfpU
EXiLHg8Xqkk5tnvijL4k5hdnKLKC8TYLl6uOzpFUW7OTDXdJiY8Xa8Q+/97TuqzL
SDjCrPV+fxT8tJAEdNEHyfvZe90FgRTrigGRNwsvVOaOKbY62amVw+z4wO8fVeCa
NQhSyqqHg0PthCwpSzOd62ipxApNAkvBAiWJKcWl6mwODs5Il3U4mpKN+aN4olHc
beYn7RRftvMs2pQV47YDaSEZZ0fp9ALznObgGI0gaOLDzMiwkSGSuih5ZzBnDxDu
s3O8xbsKyn6WbgeQ00yc9SS+yiJAAN+VHE8SSEqhAXZNsYhI9WdMWPgN9oEGNuiK
CJJDHJw6sPeIup5ds4hpPaFJJ3sQkeJKj4tWC01gXWEJl5CbCSJLgskexe0wr42G
3ffMVp8YXOvnCXGZN9/pvod1rYW8vb38CX0BD2Li2h5IEZ+37wZC9idjV+TTR6Rf
C+mFJ6JOOuMob5HdlvlfUBRQWPd0YLv2TQh/TYri111UjqCzUzUB7gKNLms/Du/T
XDn62YRj4b8YjndJU67f2wWJLYAZ8w+kWxdwBcloF3b8rTPoJ7dSUCcyr2cojcIZ
YOTwTaKIw2PardN13T4RniRluhVidgdYsX7KDCD50vKQxrWNBG8gdttVzNxxbzaw
Fa6jhSarVXOk4fgebjakniAIftsN5P6SQ+yCb58E5jPohPp2/dkglWAykbU/949Y
0Sttz/JgtN+bd1Y3EI8dYhV+383jQsA1uEFbyq/P+Ezlosp5FC6sHzcKS7JEE6z1
2jCFIB8X5uMPGYEglVaZfvb61wM1SWyV2wglPyOtwYj04mZBuhggj1WC+e8GdLmL
SW8fHVnbVDEeJgCMkVYhnNPFiP95Y4JiJW/9IezgfHYTTQsQgwQsmKSuE5PxCy8X
91z2cwySPV/KsR4mR4Ehr9nKPL4CVohCTN+LbsrZeUeEjJOP7zYsWjpG1yECajBn
TGBupSKjO3zWI8o2v9JWZjuDBzaq8lqqze4UgbGZbtCWEUCSMp24gH2k5B7Zf5IL
9luvsq3UaO/I0OWtn1eHkadWGiv2c/P/5ZVd0pQHJacKWZrgLVDZtakzXDWfE0Fh
arF7Eq+7ZnyIy/sxr+OX1PUgWoHQ4QrOLxqAlcfBK75WeJIa7gkUq0rRAGFcoDrn
hvnVBa+25yFwiECGyKZjRd4WIFcWj8c/Im5VfqE7S/LSUxHPcVsiYoGgLWyT1NV/
zmb/6FxT9iKObjX8WSO/sXTX2LDzV30eOjeNQynDh14vycbpkJd3j3H9ZcBoTCFv
W4tesrz6tHUMF1iHUS+hhGFREl/TFqV0R5nx2yAPSmzxGel2vM3FRP+hchHSc0BX
kvvcE1hqfry74S2Fzc/a9Nlkj1zg8reFuDJr+VDKYyzkgwkQBaBnrpTRcvAl8WzK
f+fL5cfPrSTRJHsZQeCC+wLtI8dykV80SegiI1U7C7dCfgH2I9EYlsCf6I2h2s8N
0wiQC2z/vToqTCRCVREn8rW/QZD/ZMFrr4g4i3AJtXISp0dVNoYbD1ev+DDViSjc
A10qLUaoDAKUfTWsZvbw1eL1KxTXrjRUQgud8aUmpWCdnt2zJd50X193DqtQBwen
KnQV7f5TVf1iaCjBLonQsctmcEflATktIsVHLZZsXh09guue4oGEb4N34Ha3M7ss
sUIkuaVW5lpjMbTioVRetpP8yDiwXon6uzRE1ESkPkDo1SF0ZS9UmHWM90aPxVSo
tHXfyIpbjs2klAf0xVfqsedNWIJbAVbzo6heFcvIRrwgHndVXOerQJF5kB/fgZLZ
CxWiJ+lSMIIbRV1RYQ9jcx20BjYrEV4Jm7Ix/a94pLvQoTIlyuZbNLJ1zINGn5nK
ZKh1kDhJxorawKCMQp2qGa9J6G2wgREJkWZ2FRAAgNzWv31qA01ojZ3CJUCJN2ob
7mbONc+ZcKvJS+2OzzHe/4elITrQfWSbgeBGJbwh6gQ98Bw9/mNkhk5QwOgG8ppN
S92h/jj8XhvfxJ7w8Ow6b6zmxktbD4SPXEJw1LO8ECG1xz53cAd/Wl4ckiYiT3IN
pQrPl8DP68FfDLotKGz689p7eC+TpBEqhrW66KA99Ey4z/OlsV2zmemBprRjLlDF
f7Muz1BOlHxwdzbCqfXs2Ml7O7t7jtX+q/b7SDIAG7ExJlDweBg/qarYPXg98wS6
gwOOXd2WRyRo+9x12hQfmK6B7GXQP85PoSu4tqxHSp6LANc5za3GhEjHjYTWIvIf
8BhFPxqSZ6OCY6T4V/WpVCiGFhVEmlMozU8Z/yWn+JzUZN5v/TP1qXSTA3B6ELX3
sPAIpw1h5PqNNlsxmUu7zMOFMLzrcpSnaUVr4J8WsF4HyCrWRWIP7JLPG/nR3fHz
sUEc2qbO6kSykvAKb0ZVjnuqjUjdrxlBfPjZ7BUmilUmEpEqi/Wb8jezSomvAUEl
wPDzjQhvIJTCGJDBWJzJIkjB6I+1fUAzfdWruypy3mHVjpu1u+aZg0h20Jj52K+3
jC9o7OfLfh4hQyKpHXAoGV+r9d+QGJ00vRGX0IB+t61W+PLuGKq+MXVs1XC0KAJ6
+9uVwYdzhtjFgsKYFEaGy8rBkY7rVjwyVV4v5kWI+PsabvOwhxdWjhvNVKPo6AXr
TIhgehZlUObbAZ2AA8E8EXfXS581/BGj3TFV5tCcmTtGt8Z+iygBeHkiZtsIg2nb
+v8uLGhf40Bys6wG/i6TFsowe5KBLe7lSVlbwKsAkOjUSvJpWEXF3/GjnXreCBKm
OrGXrlQ4V6W/ugLc00VjVfAYpBZoxdNrjXdYsDJNuMLuNSnLUuyu4HE1yB21/jSs
4hCRDOHI3uS45RDQOyLqlwgoOLj8hk2PDI+0m09X2OgBuDrkNHAZfTOHJPBxa1Cu
qjxUN5ILeivetITEhR8b7sd1I6s4OjIWGr5Dx5Z2y8GysqSdZF6o7bIRllTn54W8
+lCxMj07bl5xCI+CWbTS8XK1ej/8vRrufRMjjrKRZYnz6z62/2zwyQFKGnZkieKL
2rpH3HpqOj+ek29BYjF/iC10qWhG6+DL40DWvFefZWc7XtyZbEOVJz1Ikd05M271
91qU5bFENmHz/cite6bWkz7/rHmKTw0ZrB/5JQx2kF+R6UOJ8ae81WbEtt/VmKLQ
nb9egQuvJ1mPKykHvXQO9Hfa2VT/T3xyfbdNsccG2EZBttjSnDLcCweJBShGJMmy
/I7btS9LtKM4BRCHJaFeziMwVaLAzQ8ZhZM/x2sj7QVwrg4dwNKGjAZH4KJv9wMn
Q3GCOHTiZKp4lwzSDICqZrLh7Wb/3/Me9aDdhbTxGFtFnZdNdkk+zLuthYFoaUKp
JzzKafyl3XUj0zNM0S403HvCUWX/Cyt5K/z/Y8WQ4Epe8Ne5+aVag33zd2DFyvms
c3gVQnZnwvfHd/bqubOgCJ0DwQK6XAzJl5j3BD/OLL2CKTboNdiFoRhB9/vQuGEu
e0kfge8mu0qCmVe9oLcNr5vUOnUcJWcb3rpT8i/9tFsjxIXoFIMawPEplQtl9WHT
bSQSKCTMUf1BidiT3EZOCdBjKriDEZpotLmx0YtH1rEqEalN/f5sy0M+S6vzHwmu
3bZFSKdajjFGy+UVe1pay/Bch0CEud9eS6jd0bqFFkI5UP6wq51MyxUWOWGFW2dT
HpHxl1VRh7vhtpqzh9BAT8rA1LjiqlGfqqqyuOlK8te6IAoQzoAvmIHMqeVfKlVP
VnAitwx6cyXnh2rnk7Q3WVcFOAwmD/qn5F15mfL2777//rnqss4VkejCcgbx5Ysm
gCTnpdZjsqtaXTSeJWb6jMnNttXmXuulo2AV57mG46R+lRz0qhn4Epgz38rY2t2T
92qVwPLZ5CT/7pHi7ppNzSsuK7xAZcCzlmZW1O9WILiDXQXON3tOr5x8UzfFullB
3l3GDUmUMzWjcY+G1mRjvMgfri+Liu7ew+Yqdv5Y6htO9G0Y9Bzt6/gQV1M/kIwm
90eK8PuumCZzgE211e57YgmDD7UxKCgVRC3ecZs88ni5hnetQ67R1GvacI3yizkS
p7N/eW2fEQ0ti3vMyYuy336RxXJJWjIytf1aqQDl2XsLEDIAZtnPClf9XbxUY6Wp
sm6nM/14ojc3u36VoIeoP23umFmnbu+eXBKu8riEqPjXlV21EmYLp+Sb5j6HFBHs
Cs67LxkOouxmEyIu69xV0mhotokLaPY6PgLo0OPrJzHvT1GLUcyAOv8uyzLuzIfm
gJPrYgC8bKItsnbUUSaDlM/gNerlQ3QTYRU8WWsbh1Xin8ZgcDsVZknuqYA8iRa/
6CNlr0nRlBivYsrwbv3mQHCv0eXtY2ijKYEL/166MSx/7Xi2+RrzTbpnXr/ReJub
CHBlnYg7jYOMPMOoN7eaLPK7+CbieI3+/3sy7Z1IJbMMSVCEnMtcxEHVmA4dn7yi
awAlpK5ITM6aZ0zFBhbFJbezoQSkOYVpndOD6GN4Ugtug/Bok42MrUwjMrhBP/DR
C8fQbAbxtSijkS50BIqHTpY/PspBAC99ZV1UWA/kNmjGtUVV7l3Pyx3AD15uX4j/
FaTtwt5+Xz1jBcs8v1s349c4S1zX7Rm7qvLXsLuCFtfbIhtagjPiFz/+iW/sndVw
y9bxoM+ZEwbJrRd7vNEeB6uD9vBwUfkfMiK8He8rbAPDphvBJRicusrscBW1RRbw
YzVV4To3lljk8iCyNaeyyMKMDmAlYN7n8DL9Pd7c9X35jY8bUC2H0fNSUN7+zzXQ
MDGZLgeVbpdipSWLV8HUaoMr0nM5QcdFnohqucaChxdsOHF+c7S1AdkU1wdxWwHE
Muq884+czebka2dvTU3BeorkFl5ABtFlCVXJs6yRKU0/9iudwRKvgEuAH3kMRtYC
47ZtaXcbFqAKBH/16P6LK3VafzgAcTUjfx0ThXnTYx0qSnXOD6Q2mLRdJ1UQsc5q
tC7A2b6dpA7mzyHEqGLuIsgaiB3FODmgeiFD0hmnsUmHRP6o5NB/2P4HkMi0DdrJ
KOuZebFUo1th6JHWqXNND0gpPbV3FX1yG0AC/UuADde0vPoI1jc8/zt2fDlhyLyD
TDrdvep8JqZVPgS7oImLVCetacikFVwrh3N7Prs4/xAgeb2CJnStAgoBWP7zsipS
hFgBVGA900q8z2CL71Yendm6/OjrKe/gVsiqFAviYUSkxJ+zKvGVrpIqS3RrZkw+
jBZY7FKRCzPMdRevfGrinidWCNiSi2F3/nieLOHLaUB0qjUCGwRgaBV0yyCW6xZT
JjnDhF0pztz84OVPOAFDcj6MYIKQrflVxEjBeWy3qVgar54nm933snWrtUKw+USW
zfdE92OsCACnDi1f/+oGtmY4KfvyK3Eed5ZpmsBGSrVznMfxXTDQ6eDVvkaQ6eCZ
B/3BkeL48hJBo8VelpPR3PskO+u3wY/HcG0J2d4jvFv3Zv2OjJcYBQsCxUIxFFbk
zxbLTT36OjnBxN1GijgTwNC1lWBT5eRX4rQ+XQbp4xT6jQcrMNrSBR7JR4RIDQ+M
139fiz83b0YPK5mj7gnI1lGbENnf3h1orM3Nr8euqGJV4gUnzAYEmmo5dpWjLsIT
dxqHnsAulGsdF1YagHMkonlxM+/0vjrHl3POPqyrm+00+pLNLcsmtJYmJgW9VUij
CbIu0BknXGdo0NrLIUTgHE0Og+136xrtpTw57qtdjZeJ92TVcja+vsTt9bIDy/Ay
htIecJTVRHyt+ByIQA/JCHpjzLV1RtpU9wWxmRV8z3UvBgDHIywKlljp2LrepI3k
Vj0uqw413D6c8Wdmsmccfe1O+yH2XQbKMYprj4osZ9Eljvm1jUJ2DiCJwmEFn/u2
6Kwn/AbxFl4FzZEnkJa8FE23jc7rs2abeONS2ssJhS3Gu8vvBTb7rPBGHFWD9GB2
8QREfpDs8wzKysZHapyVYy7CYuz23l9W4rdbVM9bM5K3fJCr3J4ABDAi9Ds9g6Lg
CwEQ5SLNyLb0LtThIJbK5h+YCBh0HCAbPRV1f3xoBSGWDHY39AgYur4Upt5zCknM
yLmoJvifDhZWyTfgRBWWS8w5RPNzsNmG23F/5nKFbqGa72gLaFCf7MHYpfH1nEJW
ZpvPKHjFjQO2rzEKgF4MbSiKW754NRA2cRSsRdFqV6Dk303ukVmy8b8lKegj7uDh
kgr1ULsky79dYtSvedWzZv+D6pUQMe9kjiO5xVhgAay58fRGePj8Q3E+wD2yG7EG
AZsEAtKDM+6PJYylN5rfZjwNOd2GCrQGcpTq1ekGk8x8Eeo1eUu6jIFkWP7rz/YH
ad4uW63QBODovxNT7uu6eUPRoWWmLgZxT7emHuDtLMqCB2mTYno97JJv2SdbCG+3
P0UAJqnfS3AOfIlvOUohfTYwyVGzFRC0tw9aeeMXKJ2bKrZn8ijIuuIWB7mAeELo
RaP3dKveW01arxxZuGvnq7Cpya8VNCmp7BhfWm0NnPA3u4cJeKOuydB71IzoSA77
evBokbSBkkI//VQGrUgSwPn6xe7DT3Z1dwS7gPWfNjHaL+hbFycCZi16+kNPdRnz
YlZBgvJNiYAOnynMePivLMWmUWvrvnKBfWZt6g50bFs3GIH+d60w4Q8dAAhO7r4P
PsVLsU48pp7NLclGtnqOv0YGhTimmIoOBhyLTMi2QJ1RWUvNOuXcCRBC7QVDd52D
RODmUj0yEVQyOF4c3fZNRITXPg/TXCT8whqfks19mvF41gCHDQtDQebde9oPLCGa
URvBAxoK5qmsfqqGLrRImyj2yHfl91rp/b/eUmy1F67Auj0VPEDbFqW+aAnFmw3x
9l5W5Wdvx0hK1QnWqKF2djvLYmtG5nM1BchOaXen2b61sOet+1TIm9ZdPmCbx9dJ
N+cXLrGbs2cNUhZ16zdnmZNqDWScBsL/46XO7pRw3A0ekBAhPUZACyl80QpZnN/m
17l/hg26bqEHtxDA6MdIiqYldZjEneMfwltPI5/hDPji1vjORbrnbO90MYP7KMyI
40o3exxGWk2kkcysf3elwEdfipDa92JrhrNpPz9vw+YU+XZe9KVQpnHNUhcIsa3p
V47azy3t8IoFGwLSDIbzJSHIjjx9uXMQ+U2gbZqDZVyQ7Sn7rjjzTMfcETzgNmuR
tEZrVvBly3FZEkdtMFw4qQEKyePOWRoga5uzXIPUrlh2grcRaX89Vuzf4/stI2zT
kWM2aNlbyIlIJkHKBz0dd4V/xeHSgy8qPagISbpsdbJh7SajA3XagxBU7HoJpApN
WwMRjR16mMI2XmtlvYO7GpIhaFoR+XhOXpwY50nFlhVHeyfRh4r3+L7QakX7ezmk
tDGdSFgDYpRGjiAPXuUm/GwytwwezTjM/4WDXfV84vkDFAMcxvRTS3i39PaPq5UY
lJQnMr92YfTZTAYJWyV3DjGZJc19vCA3Mx/2cjj13oW4HjVual6xiHia0e+goS9K
GBW2ixlY6usrdEqmbEjctDyOFCeHS7oMcZg2XgNZgppck4GCW/PNurB3ezIRptwZ
Q2JwhGHfdOuBNjQvpTokmFX8D+LZ8cMO+z9hiXmm+b/2ZSCzHXXHtNxCv9BCxeio
EOMofCi/I1Pz8DzLkRwUflr86NPzQD0xiJfRoIyn+Cr4O0ZQWgf4xD3TPwyd2rtY
4pdpCaqLa/WaEpvvHHfS7J/jB0+W1DnZcZygXnNYZwYFd3f5yycCjX0H4aJDivYB
Nm9mmG1mQPIxIu2ii/CorcViO5bfRMBEbB6tUV3uA0LQGmV52bpTeCfIY51oRuaK
Y9LuFCedn+wv4sWsSsou6eKgQevBc0ivPvJXBrck7IX6jrWlaJKpWaU33ekxqvyi
IfqAMyFeCgrRt64+V3JP5oaVncA6rumMS9Nz8OB42Waouwj1PIFq1g6kDJbvO6bG
md6Afb0DZEhYXkYxOZX/8klMgmgJVlym2iRzZS8ynujeVLY2kL/PgmSpM9TglHPi
XfMOLNIhjtViSZsjEwsnqpakqE7OEhK3qzBtOkMO4PsnKZ2WbcZ1ocBifslM6nhI
LXw8qXGjRVSCqwBYcxAjKT6h2ftwwYUdro5wGQwrPvFqkcFXJSM+Todxfz0Nu1v8
eDZe6V69B3or21tsusOgq7rT0aq9G3bZETH6lW2sDE39aYr9RZS7PTR2DvSYNZGb
nT0VHTSY8y9zjBu82VabDTDobDtmE0+1U+JpmkJ/2OHJQvtzn2fxUBIsRYMeUf1P
m7KZtL/2I+OJ9YRtbIFbZ54A/BQ0mVKXxrg2LhXJiF1quSm50N65r0i416/KoOIs
TWFCY9IUyDd7y9neNBBxKb8xUzWZiG0L2Xp8zXp4whM10JDFeHY7S1AoP+7tj7uz
W7Niwl6uihZwi+BCeLYzdxxzMkAAr1UT2k8LKpNgJtATpv10+kuhih30PNhu1Utu
oX7XdjcEsc0034F/dStNVYGZjxAjjPITR7YC039eFJxYSGC144cU1nEosfdSXedF
hEABwd8LMSjeZ5DA7Ge3+TudYC33XIz6JfD8g8MT21bcDqpMxAXGhYi0JsqeFgap
rUtX9MJHYhLT087ub3h3S0EeWXJVxVi4gA8fVKsrQNqWuF1hrgg0buVnHYbY5JMQ
2oc60dq18aHF5zJ+vnM6byHpPRJ5gIJGrO0L3jDXVhlqBT6586l6dJtIbMAkXpp9
r+xxdJ74m5PRBjsEgPeuep9Ta0CLYTZWJ3IpKrbDubdOHxLJbEQLPKKP5uiisoml
Hgi1S4ehZG2IYIcfVqct+pmo1gZsFEjxoobpmnC/G5kBl5QqCDJxt3Cji25TXj8P
up5JSjpx3Cr6++lXr24l1qqk1lVW/maNq+8SQPzPE1xfbeCHr5TAi9CO2MSlpc9S
XAhog+mSk3NxmEMj6VNNrRSyt5/mjo+oPa/vc66+VT43qbO679x6ZVcVzBNAsdZ9
pmYMl189PdVBaxQL0pcyv2xJvYtTJ9jDyQlsdOZY1Q3kXPvEdS4xEtNeDB/N1z6G
k+mj0zhUpEu3ky6oW5FniOH9rSHd6PhCQvlDxUGjs6YAZOOATzlti3hxTD2vt92f
D01J3jjKMtVpcPh63ScqhKGw+D7P2Lnm/w+Cy7yfMZTvhsMydc1sv0iQrkg8M7qE
rWS1ykpd0ey2QGxVFcokJPbuqM1Ewjg8o/FCG54MJ9wu/gnv2fcjUNVKEjnl1NiA
iytJu+NuxnfG1PTe9mX8mCrcBufgdwWtsfC9xLW440Dp4djIsnjwVqP1CeP6xuYV
bYqWogY9hJr3DwzWV5+svs8lEJnNnSDgwuJF0X3XInJJMEgl+eX1SNZkW6Bn+DkY
ieowOe7tCBAF2W8EsX/pFq5AoC5Oi7gHVQJakzqw1xD0QFmUccl2GYDPbVif74yT
aU0vaDsh/qlr92I42jPQ7x6eQosd47HVKgPa+XJB1IR6dufR0Ru6hDxi9t7Q12a8
/VOcQpWF/abUqao/ARR2siA515KqLmObX1LMAusM6b7gEPDy3+p4fQHdYkbaBhL7
ipAr49xeyrTLy7lknPsBBMd/aaSV8eMCDJD7f3WGsWhQivVKce/4cVR1/GnkQ13l
nImseBylj8r3M7/VnZXsFIvsaE2lTfGcDtRCtUuhcVGQE5M+0l6xJ/VFkYIxEkBB
MxEIxEpoBJRE1ZqbxU+TMDZ/dQpZrg0zRQPKDPUmICAkrrCgMF0OQljC6sb9reup
kvBRrt9RtNzWK9xYPNq5Wq69Y3Wjtf4K/vgyOI/yQxJDyEwn7/ppoF5U7FMbIeub
OmFC9X3F9gnUz4w8ZlINZQOR9C/LDXqIBdHcWzjw0GU1JDbVnGFuiT7p9yEUeNxO
YsVLVrQrTRpj7l2FNW+6fFh5EjQUrraPS8YYR3kn4oJR8CJTwXFPYeqOVM1W7plU
8rf3l1oteHRQCqtJEiYq+FQl8wG06ax2/Xqe7Xi5Fv7BOLf+/dRCbzHfsdDu4du4
7cm5KkfUd916JOAVrTJJ+fz+1F0GOsoW6q3i/3f8h4veKfXJm1VMdCQ6jnLY8HRp
UpLg5dGxsKd8qSjF8CjByrj0nG9no8aQUDzHfKCw9dA1Vn/Pu+Dc0R3b1av5sjlo
PYMT86SpmP0/04VyzrD6ESOOEe8nH/iiKaGMNdQzRqq8HEjTJ3bE7FDvhgL0Bsa8
N3WxIPpiSmK3Ri+ANZZr0OUUhaNDlHl6xz/iyMmpW+NASc6uZZRRazoYNoNzTZC3
7gPpzldFvkQrnaiXmgOQ7YZDH2KrwiOqb+AuscEWi3LkjLKZXBLUzxTs/t2B6wO9
+XgxdGuBswhJtutMqwqO+NHLw5R2xHkQ1QMeJraVsYVhamS69rGonFvKy3DLBSv3
xFC1En/U7Yw7moIU/vE2NGS1SFfE8XcPoj8jb3mMebS42moR85/RLshUMFQZbz9J
oc7FWIW6xn4zQI0CKn6nPMUk+XWFVePc53Q5ikkg+WQBCON7xvUPvNJnl+MHv8B4
IpK91eEl/fsGs9+aS5Yauyl2lUgF0SlfJwt3C/sdkzelnh9PcyoVCgonSTf9KaqX
+kmhgxAvO56WQe+71WqH01uxRiwbIWBPrlbQxhDckBvTJDlrzFiowXkoAPOddR4v
3PRQpobYSTkn5qcDFKBetjG2GabgpWGJLAdrolWnrLHpuF48ATDy8eWp4DQrxWTe
yn/VZeZhP93k4PYo9k34djXOqANVQU4kftKuOoZe87FqLfLAJw/GQWtjXHysVvpy
XpKkpzImnSNkXNbrqZ75c/v21/X0t8LkVHhHkjmVBaACpQIUtpJ4usCn9ibWEMj2
Au+9ZP0+E4xFnLj45GKK3RDQPwxAdiEfkhPld/apgmHo3c1Fxsg2VEdMOhODpbQy
DCZ41KSjxWX2yi4XDAvNNpX8OMjUrEyzlGBWMXNkhyjo88a+A+xR5famHu6Ajs7k
hXQnXwGGzPzKzostkohM8VuUYF+8ol6PXeQ2iZVo644lX41EkkPhggq80WW3nMcy
BNVNW1x+JqYJ5CMkwvz0kNWKb87uLE/t0MRL3d7wjgSPj+ZxZQhUZCErh7U0uYnd
EV/f0exmylA5m/S4rpOTh3FamLdYUdz5drJCT8Lp6OM8UHa7oei6xaLq8x8Ahdt0
UzF+uM/fUyBqWmw3qBKXncBsd1uh8lvn12HqMq3k+MRRkveUA4y5ktcSyVqlnp9y
MepOQpS9DKs6qGURH6/IBjvaZdmyE+lj8aGSdUws0KhJsGgyQuBtL0PgCOwkwNmO
FEb/iLAXj7GQjKMXIWh9u3lMaEnOtdRFv8kKfiFEzjSHO6zWjn/Bu3C16Rk4U0d7
OKp9ZGZ9tz1krHNBCAuFQmZnnjhVON+ERxZ9svYWjw6c9fhu594t6ROL8Sbn+zrB
RJhkIg55Rh8Mmz9CQ+Q0E9jZKRqYS3JqnPnrTwSUuQGsJM/tS8vyGRwAbGq3SIrg
l9ImqAu7P/RUZJagTwINzt7zwMjuEwSC5RQiZltLFgfpumCq9ldFppEXTx4GPS51
8Rt/x0qTdrfgbJk6PQhIbfJNUPV8pkWewSq7aG3ZTm/DohPpl5Jqlnu0RJtRa+9f
3iVMxqDZDehMYnCwYv9RMchWqEVx54CMQWJaHPfJCAKS/fXUGz61VxAWwzXJakeH
aq2yr+yR+ZGSBo3qR9FeGkEc1YBdkKutMccVLy7whsbOE/x96mRH5dZugdDYM+hL
b5rex6xle/2s6SBiikDub7mVtOiOsQb6Uhovnqgt0ciD/B0FHcY4FneBlLk2ZyrF
B1x+/3L6qlvjd/Pb5WI0IQj2qSjhNGZn/+KPgJMDSBbmPVVNhxLqZW+XrHbXlnEX
iM+VaT67G0MH0pxZH6na9Lx+ApkiFVnArfVaWwZEMQdpO0LpkOKqddlDxHBwarAk
j0mJgc8V9gI66qbcbVBWLUvQrBz55JChv7XAEKNkjI52QRsOVW3S9039aOltXwvd
0TTluXAqYV1i1rLTdzq9WPtJntpf+gR20ui+rkrvQjkjdIAaV3ajMJsvpfngCody
eq7Zu1frkAugFjcq49jnTOtMdsF8IUFUfztWtj0FB+mTsPsoI3/J2Lcwbmg1TDVv
MTBxJtnuNJcIRzgsVO9+ouqVXJmZOhvv//hu1ouGtVu/w5kXxpE8JZR8YSt00dBk
77N4RKPqJlpaEUYGn8ebwCBOsWjOIrFYOabUtnImJpSrxknpN2tOoPa+Y9zhIfh8
95fZr7xbNTed4FRZV3bUAk9ad7E/lkqocQ7rJi4q+VZI+axy4GB5SutouTzy0ifD
BOz2eCba99RTi29vLBAyhMAvzcpf2kF6ODTb53Q38g5r9v5ZqVOVTtKKDCFW59u3
Van/VFkwmkEWpXuXQFDT8uGIwTsfMydYUM0kr+uaCvYnZz9q8U64HpvyFg3xFs8D
TXrWxrUOVZWNLcR0A+ZTIuMl5yjW4+N9E3NDAwHFy0Z5F4mODJR1Rwt1YbZ1TvRJ
PWn4sXVnLFwfAMSDtCQf4ge+I8UHA5Kp68H9prrOLTQnIJfV9BUCC8rD8yLpkQRF
Yh4tSa1kIy6qaYfHcAfbuYW5K+5pNhZDu7E1D+fDhyXYKfOn9DajNudpl+vUuzqn
+Rzo3AsxRZkCzDuGs0aLC5zf68EEn6Da8PN523mYcNnoZPUgLR+qRyp1JtH9Dkkp
YHBXHskgRZOlj8rbdVM0M46t8XWCI+3n9kq7f6b1L7JQTzfgAW2LWlRU487t6Mr6
xgVy9wHD2m0H+Z0taOZEQtQVp1V87OL7d8xok2bCAPEtZpla0HAq7hBYIU0jA0VN
zd6E45p7cy+DQH9trtVx6Yt3A88jY44gYISkVyzxxho4qUohVJECumWwBhT4uVKl
MkYxrzQALDMim41/WntnE5I0il0z32ZK24ZobBYQBPpzEhh1j5sQRnO17lxuMoM3
Lxz8CIGhekUIid8HX1PFjgMlFxMV4J7Xoke++OOP94IehcYlD6XP/wAB9/gMdYqd
bRlyLZ+AZp99A4tXjITW8L0XqveqrZngbjW0gjV5n7nZrIl/QO6uEil55uAAgElo
Pyq4DIsIrecI8Uve90Wr3CmJRDb6Un6efObJYy2I9PhHU2EsW+1a5kARx0zNCOwN
ev/J47h2aHcj8N6/cnZz5J0cFRq0rKR4S3eAzCtao+KnR5E3JUBIQDSCU4JIITgs
qb9MVetO9XGKBjinbpar16PUH5S14zKAPrS4cFybh5bg8O3MNthd5TyPlP0OYtWL
MvVbSnrBotUBok3oC/mlvrskus3MOON9XnKFjzEGkBCkfupiXUg4u3LeEHq59z+D
WPPYQKOtAY9ZlXtkIlGKaIkTyyv1xMk5pOVYMvlQvyUCyASB1yBQ9oO5nZNVVHGa
uawriaFD9xwfwfkhoWJDUpX6UNY5WYO7bbjJ6AepLxz1sKKxHvax23WmFOvkQp0t
E6i04J2zPdg4oRPBsJ1xRVSFggc9RZBSrTJ/bf7daaL+2RVU26jgRqVBbN1kFdUl
SYs9YJ1b2IyocYRCWcsLQZJaexCGI8Cq9hNqxO6NQpxPWBLE9mhrhbWrN/sL6+Gz
HRRvXNjm08V+5R0OHrYBM9QI5W/wgIuJ+emWhMwoHLxHwzOaZwpPPPsGGNkZEbdX
61iIccBVOwgaTmb1fWoZwC0O+c8wew5HZ4eiCSYx/E7Hph7mk1vo0ZOjW73of7yh
uRARUyfpjKTqJSB7c1Q+vWlIpqwVtoxjJKSP9xY8zHItVX+ugcy/fgnfYPok0TIy
0QeaJZyHOn4w95zZX3yI3kYzqCNbQid8TdPFpey0nk8l5+PtLVz+FIg/Fc5QyNqW
hT3HChL2NNL+t/diV73Rb3QbhzfSd6PhyZR+g9XzrOVh6RHMVS3nP4yepKq53ovJ
cM3DFCsGWMaHOz3ZE3UOjNLtvwAaBzxpUWfTtvia16DreRFMvBJAv1Fe47Qthzrc
DjATpn8e66I9bwU2x22v4nc1ED4OKT3NyKpqP3d7Z4oBWGqa2G+5HTmwp3ZB9B6h
3dha1KNnvPXZgQ0yueHPHnWouRe2+Y2XnBB7RwGpnAOVWkwegI9PxAv3lIM9EL24
KDYwwuDHLoB+zLCEA25BPFrsqGownnvqCQdUagmMd3+f/G8ftihko3690ReGR+W5
ZP/D0kHYvUq7lqb6D8jT0hcbfhw94/6KQTfiNrn5oWas7Fz8+EOsaqShVTQkkged
LJGBZT1JaXpZBzFtCyB4y/IqorzrDPJ9XMCAATBkdEEnnYUa4RzygQbYGFd5M5hq
gzFl0Gxl4P/97mR9ZLxjmOKM3ml/VBU4A6f8foul+eyzuahIKEqjceEIimuzW/xP
T/esFU1G6gT0qL27vfbyKidqlfsXHdTpXXf9CXkY9PjanwsziIFtyrlcxsTRCRXw
2/kvUMKxEAm+MJlU8+r8L9ZRaamcj6InmtxbC7DodMG0giKIFBXgFnoFN3VfTGuU
eIEKychXE5wR+1d59zcWamiD6B4gH044AHz0ADXrbY1nJnLF7DOVYezvVFaVSxzQ
HeO6R5Da97Vb9l0/Th1jpe51wkyXOGeYwiuschwpvFwpN0f8hOaKdPvCcRJi+06O
NHRNiwwD9aclXULetDdqHZ0Kj/I0ppzxTJhP+dn3FWYDEroclnDzpKdTanHdRytR
KjejlwuvW1a7VMU5urYxTwgeZ1gv3+V5y8qTCEuPmsV5RLH0QQMv2emlTZoqkfT5
JK2tNUyzRwEfwaPzVDJJOthbUrtMxIsGhvVOsNk223R+9yFPkElCgasZK2MNUuDX
Tsix2xlIlMJm6YeS1k+xSV2G7VyKYSi2fG2C9/sItvsluXGE/+t+DizdVNwWbFmm
H5V0oDiqaLMxBFtPHpQdDS20WIcW4VKyD+i/40rDPgx8pjkN5/Zz52bC6mjg9D1W
0hC0jqcr5td7QSycwL7xrn78O0FbhixpHC/88IVsrbzTrGINXA3BDBIhHxcfJ1Ad
JabFpMsaZQbDI2Yhv6HE5PIeEeXeXIze3UQuwAixyPapnGDXiG3m8iJVxsovx4PX
rCh8jAUHJ4zhgRu69Dvsa+ox8QcnBaaO2YvJfVHqxJEXGisrGXFjYJN8A7bRnz6c
3aaV4BEopL6Zx6ghOTr8PrateTjdIGWLbE0iYocS1PN3bBhjb2Jf5QNaX0Pcipdy
aH3Z4F+N1ZbsHY2gme2btcmSX3a4ZOLn+sRGE7CaQjM5eMOiPFsfJExDkYLOlSgd
Pe9bhF4jIPS/8r+sCQ5D8qTzxDa9S1MnimB1BpCA1MYZVhK2yx5iMJBcLiwDPAvj
LhSKrTwzyDEewo04nBaqZWPu3gos/XkPKVdyYY35OtnOBcVeXHtmACnGoLs/TP/8
iuyf+utGoVLbDk7Fqfk2ducYGUvqJ7Zsp+hNTdVai9GI62hzM4UniQ7JlaKljDcB
/RMu90H75zW5CiNHr1tivIeEM4IjJzDjzS/f1uLe//ldooYQuLbyNRwt6X1nAKxZ
b1r0ema9ck0GVHZmJOI/UBOS2F2f40VrTpjZD9BcQaGtDi/Jqc72k8f51AOGPCv/
xEP0hniXi/2SYd65IlgCJJAJyoBIoK4GtuJqIzAtc+2PWtY9Aj2Hs7uSTOczQ3ff
QJQ7f7h2q9Y8wcH8gS7ty7DM/4bkVkHAe/k8q5HELBPlyHd0k3BaMbPmPAtrc/Q0
g6mzJFp7y7DHK+cg+paiX9yunWPGkKxWy6fpypjp4ZyhrsRR38KZDPJ6WNKsDlAo
qp1+tX+xb+heURqBTMqeVOu++w8u5W2bq0Veu65varomskBuVLuSYDE5Bu6ql/0b
jlY2VQh/1z0KhQc3BhJr2Av91ZWNM6S7Clmc4kkMROHrBqhSWm4wkz21KwWXMWnt
eGJEojXv2p0nJ/2wSQxUYp08az4+JwG9dO8JPbuHyismHdBsor168vpH1Frw4Zpo
5v/HcY0vLlhNZobbPPmwJjZBWtYNK7JW15PfdoR51ZmVXt30wxjO2TciWy0CEFHb
5Akko3/Z4PYZ4cVN1rqdlr9XFQhxV5wucaMnnrHmtzZQUL80YG8GftpHOVVvPdwQ
3Y3UEQDIZs61p8jZBXjGN38kA6hvhJ+phOJ0rNgrslcMR2R+XMpPg/Wt4OzGf9VA
+A0oZJHvYGKBVrEFkYEftKi45W3j+ZIVl4K+UmGidqq6X5zQBcbDUyYPXVmBiZcy
FHTrpbp4XUPhprI13M6XplwurUbPfEkX+rQtnFhZ4/RQXj3or4T+vwAYKmIwemb/
e0dEoNdqE7xMmJiTwlxjT5eTN3mTGc3xf2+kCL+f6T+8u8dGC7Jqipx7XxDngZDw
0xqwDJm0IVV4Q2oGJa5L9pN8TIHcg5wagUX2/UCSWRC9zpyTt5r+ahxY9tDWxfaU
StJ3GXeTPct2ECJ/Lcn4M0HzoOlmWz+rhOt2KE6W/80hqG25/STGDUn5MUcuSy2n
DLAVru/yBu4td36Ehyhg6PPCZgWfT0bK0RwqTp847ppDJrQ1ujZy5zwxU+znenZk
pgk78djTz7Fn2op1fuGSqVMJLoqXydHhNj9DhLYvlbr7OF8EX4Od60xazy7X3ktQ
scSucnzgt1BNoPmb8jG6YV3AfM4N8Y4cuxO0oXCx5SygNWAVvqVwS2BvXCGWTBU1
hwugKKd7v24UZR4/Fv8AE8QMf8XgPgPnmsyG0WIkHhUtrG+sjK2kjuy//H+NPgJJ
BUqYPgywiVaCWM36j0mx1D0QSostCLc4wCrDusvTRDhuZuimznUGglvRv/dIYWId
/lut9Xin0YMYS7EwBCSUnM94Gr/1to6Yy+8JgQ3UQDVLoXNPnFoQ7M/qptlVefzP
iECyNYJkVxK3rtXJB1rdrDkIXsdeOmMyPPq5lEzMCKiH0+j/sqinBOBE5mEdYwhM
RH+glWvl5KUdNx7ckokq91iAKAk6x8/vDy04bWuO20Iln7HGG2+yTOdLaEMBSfAi
47h6RAvQjONJc1zEWriORpgauI7EY2rdHV+3E1+OK3em/4d7EYUqCj0uBKkjOnkA
FgCP0uRMWJvqBJ+er1GzjwXOI2DItsHJmQAHvgAOyiT3bGrfxZY4eONonobk3IyM
mPjl9ZxMjy5/RZqlMablyDBzQWXj+mgte58ZxL07QAZZJrLgPDh5PO0rSp2EYVy3
qc0BeH4vGuVywVb6Jvkibzn6Wmyk7nymhH8HeeRcbQJPev+X9HEiFSH0AE5OaCuX
qEtO/IjGdd6tm+RGP4H2AQbf/goWQAt+GVZ1jvqeDzwZqMZjxme4sZQNP0FO9hNr
nFz/MRBl2L+o1scw2LS38LJqcD1CpA0E666Mo3VlU2V9xHfnRBWv2atcN1PPNNf9
T73wBH31Zzw+h5AjdhIoaWmpie5wSBdy8FwzO1ypHDwU+tYnVAowHGrYcs/hwjtB
UeyB06uEuyyEe+79VhID+rETBa1RAKY0eA4DWh64UikTEdBCoQg9sR7GHbbOPGdy
Sv8swb3Z83IU1LCjB7wGvR0YEI2+nDTlxec9AjSULGsY/3eMjFdKdvSBAjj3KlyM
7oJq29wK7yHSvUK4lHoZjBMqHXPgxz7wtLW3QebpWCuS4zba67wkqqB0SWilvAGT
lGiYPXVC8m2c3sCyNw0ywMprX8z5SdM/J+/EWQAd3rclkibJLlL2lhkkYm1jrYAS
qiivUZ0xhw6vFsHCwjrcFfloDpNaeDEhv9gZ5cuXX4u8AWhSVd33VEiyju6eQ3vF
wi4uM4dtT4lInGvfekEsA2QUJT+OqR34HkdK50o2IYI49/elLKXPRD/XJw4QmtsG
y3b1xcv0StXiIyXyElvydqM2bxR0wxyDU35OtKnmzr4EjVUmz6ANK1wZBHgpxPTv
iNFnAZMGbAlY7czyxpvR80bjU87EX9OiQ2l0dIuUjUwEIKanqsfWgWPsovM51bJY
s/pu51hHXI3LgMUX2ea2EzBekPR3le1UMqp3fEjsn2zl7SIIC8zQURQUJvgqgdE4
Gi9xYVXhHMY/T+gn1uRZKmNjDIYLe4n42T35trQbYVGdW7BjD9S5RMIN6ysOGpiC
waP1/khvvZ8aZD+4FjDDSjH/oOwkzxSs1AWm0a7IgwcUetFewEckWtunu6PCoJbT
au/pbU4nts/ZuKEJW2eE8Qo6bIwOE3pv32ATIBQKpMjB/GYPAaHPNqfwYp5OC+0+
lOEnK9PUKZQp3QTv4Zn3bdgQyZBAl4SDSriYfw/YQMRnmV1eyZkPZZGnmsaOlSb8
BzZGzTW+hTUnDbI+PLarP+fI9aDmfQuH91XP0AXvJVfcubX3xvXpA4WAF3wIaZ+q
gi3qswL3RcASGSwawmvKGXrdT/BtBUan2IFqkz6AVA77NXJI21DPCwIUcFUHRimW
UqQp+IUU0VyLGes4gqG0hfvQ9+wZFHI8Ib4C1w3eR1V7Y9Mxz1aW2Q3e3BJisNN6
VIg9X07/W+h+s5gP9mZ2wTi2RWXRiciTcLpazVW85RNlRGd+ogyT4NsD8Srl245H
RJvl8jcflWYfvyqyDpnl/ESp4wLHyfiL9YIu4ChXdwQUhtM8bYFP5bcsQviRxbgs
6olK0X24QD28K5y9p7wzeY4liCUQiM5qA2PzehHR0938hfacTdC7wa/dcju+g6wO
bUUlRo/YPEakEH42vs+m0nKeinKO2bhTz5gdaZSNcFIVrHyA2flaMXl84Kz1hsX3
MewzLReGEyiViuc8tar3bBSBMmzTQaiX1Uq+CwuFsrQ9OalWE1ZzfrRPftMtmnba
cETJmAOHph+3ifIqBbIJqMUy5Ven4kUcGDCH+f6OFyFwVPRa36uwuwEoBYKZ+9jk
ZIPLV94x9sSnXdoMWzn+wdjBldi4JouU8YHe8md/NZ6o86vvU+gS1mwOaC9Du4IV
A/Kq+Lyru+W1hiupHK8FvlAyc15We2ifuXipgRQjYKQY9XOzd3ipwoQcVyOZRdmn
CmQdv6pncbnYGlgEexPHbEoqGYxEJtnWQr2IPrRKRp9vHZndo7L55pLgkRnf+piY
AzWE25tmf1RczEeKk3jWxXHJtbWkxSQIiW5Vz64CDMexbJT1Nl6mt/I7o+VX2PMo
0wAtv0dMFxFTveqiMsMWHiKDLencXCbiD7bwOc+6aQgRB0uhJDyH9Aw5yTwFET87
6MDimYlqsL53Lv0u4To4Opzk09zCMk4gBgrfYQT/oFxi4p2IkozYRPXtZe8lVGyO
7ocH/iGeJqXGNLLTs80Kbjzyx8wXE9qnimR+JP8J5TzH42EFwrRz7Ki7u80imeu5
c+QQNvhE4tVM4kxH74sZ1h+wm8ULzYmQIlpKf/pngPPKKq72KFnfEpYcT87yjW45
vB8IWX7cYEfEQLyn4CS5fxGmfZJ7UGnuI8UvhLJRdfiJ7+b/lCikZpcHDNDlj8Sn
J6eRpoKYUjWV4qsBw5cftT9JJZVDNtpGlFpHW9H6/aVSSQ9iemmPGLFbYCKP2zvF
ucoHJLtaOTrS10GTz37m3vvR8T+yUwBdEqHrmhN4ZV9WSNs7K7+pOVTKjyjy/JSJ
TW0Q//k94ezacl99UXi2Hx6lXylcOUFAyvWK8gMY2KTVwNGfVygZf2UHZr4dlhIX
Bx8z9p2CMhRpyHxMYg8LQ5p23gCVNVHymA8iaDj0WTpT6sC5t7n3EwEFel3NnKaw
uyffblEZQbscvTExPPWnL1JVzel5+H8Tkl4iKPibeC4LKZZ9n4PO6vKFUZlujJ39
urOAlrWIP9cPZ1f6wd2NoOIesbkOfqn3jL79Z+3HcmM+6XDx9WdLJwLKdXtZ0nT+
zbPvV5g3sNUx8X5TX/wFmKPC2C1KAk7G69rZOccyq5Lwn0xDVqHJd0O6MTfO7eye
FqLduF2cPs3Em77nTv3hO9vlnTsvc7tHnNr9HIkvN+g6KKivRS0yZlvDsMMB+9Nw
xn93SmOmuTHMa8zaKK/kr4eCPjGtVB9CYEc98I+KvU6nZi+wrY8Z6AfsOH7D+kx1
gG1SPsdAcVulLKmxR4fZmFcNbnuVXERd/DRioJtZmQEsJ3MfSYAlZAH+Bq6iBa5+
UicBs1lx7JxnJMrVIO86HFXMWH3/+d3M4Vj2Pgah/5fNaUeg6fJ+Iu9HnjPIIei9
vuR2RYAwPP2qL9b1aOrVGeaH/zHwZQtDuaiV7So/JJ+TR0bjJxof192dfR+D5Yig
4ohpiWN5oxjQDxRNuf5kheZG77sQ9TcZ6dOSdBRltIcEWmI9pJ5cdXg43gEfXYOf
/oLH5+uG0CmMm5nNrwiM2aOCme5Kkes0jzZWgW8uuupeRPHIis66WlzdSKsaagNq
gbkKKWblb/S/yPAM26TslNACU96te+/KyeVWAOyN9TFm36M63LbFUeiVdA4qX9bL
FNhf9TR0jtDbElxPD+PxVI1BnI08XemoPjUMmjGESvroB2uXEJ6mde8Co5fUlYww
j9puQnHE3JTewGTbuh4MXd3u3qkNsgTLH7lahCi8wKH4+yE7xjnks+n4BR9Yq2wb
IHBV7ucOiDXbnRHMpaV6Mtb12gToLXJ7LcXvsThyGHosUhr2Y+NCTlGOQzJJHNrv
tmKrOjTxNDqFfwRwzmoSJ/JNnUGexqS1L+ja9BguZsG64IehiTeTHRVifdI52Egb
CpWP1Q+dkLkBfY4bwzlQY1NiWC6HrgGaQ5WNJdlSuOSJXAruTxmz7XjRvI8Uljqm
Tyzz5h1rvbh9VS5ZYAUPqQUeWAnxES8eYvjV2Pvc0EPFL+VwuRceHKbo4NoOZflr
xkLIgGzFropwXZmmRmUk8hCG0mE41/id9pdJ8qVhmjSekmbHuQlk1eiDgvxO9og5
7CdH++EUOMvHPD/TjvLQJ8RvEHzNTxSuGnWFj1C1z2L+oP0TKuiDDuAXSweTILvf
oMQo7oghJ33aZY9kX9qtiyKbJIBJj2qB6AO3cDIn/tZC8jg+oS6y4jXtl38Pkvq1
/9h3CyM41cNBrlIi7WfqoLSPZBIWoHMIpAXRiovxWDlZNK2Eh4mxb7y4BpI5nZki
NL/GlSE07reiF5UkuLrgvWeyh+WWnCGz9h7mH99H7+lwqh3mwB5fqA+Smk3L98jn
kx+o1oSF1iKXUCFaF84pxgJmx894Z/8L2JFYgFeV4LbC0CQBdvzmWqN9FVPl9wEi
cb8gLfxiKN3ZnXt/tLWzYe3H9JlQWrKU13RaZehvOFlOMiZjJkz+Vo7Ocema6geH
ympNQy27W1Pi1SMnaYjrWCFHLtE3TarfYgql6ww/NAMY4s9iWYQi1BsEnxgsIVTf
o+04bdpwS4E84Xl911Vb/cCb1zqi46q7yBbLQ7L1nu5bDAMBhsfnpd96nK/T/vDj
dHTltFFh7LAnYqYCM+1uP/g4F7cEdgFO8+kSVkyn6UQCO/RHn9Ko/TZE7wSjOB+T
o2TNZL9+d0tAF5oGFk9XwNo1++Fe72Gzde20MfhrYOsvx0U+Tl1fQuQpYBmzAgwk
njvQAMfwt8CrgUdCw/ROFHQJy9HmiEvVA2a8y95UL9L/tnlukl+5Dd2TSohcoqyD
qajllMVwdfbBjTg5aG4AhQtLcDi2NxlbW6nWK4elwbCP8ZxbeQxgVicQUih7vZos
UIbVBiB3mPNjbqqpoPfnVmPwGpOUUozdREIeoJlioI8TIYYW68EPZs3mlFvWy8lZ
hiy+DNi5T45i+oCAb2C0YMPKY63x3vCDgEbAe3sY5QJNN7VEJIRdBcHyhhUOA7nm
tGB7txImyom6wG2gsOr3QTc1QCSyRftLND28/wB2lXXSg4RyXZDwzAKDrIdpnZUE
SKJYypVKiLC1yi6WMAwaf/F3PYdSjJGo9MjpcZfBWnlAD+GPyMHR2xzNGCDTUGd2
NF3SGvR3AAalBc+OD8HRr9z+rCGy7/ftwcHjg7H/odPiur9261SnGiHlgONkYkCP
Tf62W5PsxNIb05GXMZx/zFHhZ4nGQ8NPTcbaAiS1ytuJK8AlkRjgFqShaDqEYh4E
RIcnQBm3HTQWpvsB1d5BEQpf6IiaIC43Dhka0HxvGAypc7fOpUuELYJNlQzK73fS
dGT4pAGNz+eqM5QLRxNLRv959efwU3IzVuGBLR6SbAQyI4aIjRT20mDFpX16BQ4c
aeTuN9v2rAoRRK1+IHGNJOGi2jCgYRQwJ8Gq633oO2+HoeoB3xjorhZyGyz214Tu
8pev/UmJuL3R2YRsHzYryuKas+L4JUEALwmXk2+CFAJNC/gHzVupqJyPhamzb5dH
WPMpB/lK8rUxXj+rrhwK5ermoSPJjzW/CfaBTiTzS84m92ND7VZbKFeP1WoAnVev
E/C/5GO5/XPpvsm5SPDnhCe30l2Tx96T+qUadxjA9YkqkksdU384GpIO1LA7xze8
SGfaTcf3tBL5tPfbWmO42GSiPXOa4MCCCWceCCkSOQgFW9OXAat0ywjn0yzhetj5
nRlMcFldAugKbIqD4KrNlnmSFHsEDu5ykKFy0chTzlxYo597IdWQeBPwjQAGv+u7
ekDxfQ1Zkg2twi2fwrjZZWUGvquttUzooWmsDqBfdw4fSzmTDrCNygZxY2hffWjB
28fBr+UmBr/7BtRq7GotHmNzx47G42GzJ/dQun/Z6ZeVXiJQl28NRZg6Pe/cDsDx
eZHIMmvcHrkqj1xwgxqqz/eJr0yz1sOamWpzW5YzlC6ZrTi8Bi7pz58NzpPCz194
aBAxH4Bycagi3KI609a/hQmj3LnZOfgKx1/y7+LGaxQaaKO+W/PdD9Imy0sDwoxo
Vw4vAzvTkibDkkgzCLd78RRMlAx4vse2za2VkF9K4C0VDCvk2M3EUNg8e6Rkfp2O
N5UST4+nylVsFJzO1h6Wi38MDKF3rH1yNDK2pyygmI9yEmW9SnSrN+XNqNGoilcx
G9d7eVswcFDi9SSuEA66S432VzXGm5395M14y1w9uPwOWOyAxOrWVvKzPQHuTuk2
EjkZdAWNb2tl3qGOaKoev0g3NHMKJbWlKCFUKZN2WteBJRnhELz1B2HqtcqIuuDI
Acj2Jca6paLd3eLCB7y+YDoowmJmXKJf/Gn5DBOv4pg7mSz2xodTOq6j6ZYzvPg2
WOqImnUBHg5EkVDc6HpQoM8FShbbBQdICRkeoPjcjsrdLkY4P5sJqLU2gZzizPHB
I5Uf5eoBnaGkrbMfWMNu7MzBoV6j9JDce+VoK+36VGu0XEO8Etc0XxK5zeNfRn4+
x6owfoBHtFktu/mDE063cmGYBKhcL5dX8MDN2hJ62vBERfttC1W3dvWyE3fUzm5J
4bF2UxPoCEB3c+HYbGqA/0JTiG/wCKlmiNQJI2rwuaR/z9U6tsJ8IsV0UpYXutX8
o37uly5Q4vrr5AdCSqeTPViMnavemvBwy/hUkqOsTfjItrvfnAGzKiCsMc1if/Ha
2ZOLSQ3rJ9HCMmqaunyR/KSvSNbsQg3yL3UTSs4IwWu3m0WLzxa2eX0h8DjeHEyg
5r5ar7gkwAxsPyfFbbhq2haPxWuRJ/QkhWFuVR2/ocbKECtDH1vPGqOtVH26hA0t
zYTjH+M0R99KRSLwpUgjdc4n00GQnYE3hexsf6kc0H1G8iX5xSDofzwhaSHWxAm+
3Qg7sVyDn4gIQNGGKlj5uPH8eiUMM5x1LHvy7axLHL+23aew5339eaeToJVOYMJ8
GCKAVrsHcWdAUcxh7Mh485/eGXbaTSBsRseB9cuIZOiSL7xQAkWBQyLLmCLDWbsH
42t+k0ZOVe8lYlZIGfa1RRJ6a02Yy9mc6Iv0elGKtsByWZ4xAjD/LC6uh0aGdG/m
49OnCHN2fweySdhWj57BcUARWeNyY1mjM76PvZ9XiK+0Bn/kaH3+mV/+8rws2U7g
uq6/vDfsI3BzHWv9ZrG3HlaCRwhTsa2YM/FZd+Lyg1A9u/HLhtxcjbDKSxRIIwOw
tOAc+x5pEsI7d+X2A6zGl+63namXC8eJE6McnQuUFKpETTv6N4lBmy/cOnTIB6xj
u2mOi/IzoFdLGeeYxD/Q2QMQeK2PqUvZsmtEmj2TsUtHnqT3zUI4hC6jTA5IuNUj
g2wDnUTmXuP0Q6uznPteesS44ZneXhHrx7CoK0X0EdDahMFvDmIKD9Es04SUtJsJ
9jRaZ0pUPiimu2wuI/Qw0Qq0XzGigXBdKgC73wM74p0Ui18S+o1Go2Qj7o7BfhMU
80+sXvT9WhUuH09SS/1/6QXdcoc3z3c4eNi7+D+7Br1BrCv1L6LiIjHcC7udhkLl
fHgy+5bv9YNjP9r8JK/7IAyP9Wl4jwbC36RCqoTACj3t2wFL8zsDJPvIdM/HZw7P
dUNKu09FVVMqD/VqGyvLZno0+0jLFJEAaIjHNnWuF9Fstf3UuGydBBRjnyKzIbxm
1G9CIewGplj86VXTUnLlBcX058EUJvv/Ttr7cdGlkTQ2CSTDf95lk977O38eaDSs
vflri2tR0ZXEY7kh/qY/FGniaXe/h3viEodHupo/xbBtHBLgfUU7VC6hBOmMUTiX
A9glJbrD7UaoidRudFtsj5cAc9rfXZIzww7VSxhQEOONu2j0p8F3fsxX36ww6yDu
j5rQZuCTHHtj3CTLR/rBt2tG92TJ/VeWBD5KrPX/zgt3FpENlOdlFBgCjrqQwfH6
RoEqI4MXl3tEcOG9aVI8haxd6tegcEAfzUBOhh2a2zVB+P0b+qAQCQ34n7kyrH9V
eBDH1m63XOdbXAPQZ6J3WOSz5vyJSCm+o0zzvxzeszoX2O6/0SB468OWwiArqf1c
HKagDxmk6L5botXxTRlrl+pA0ruJPqJSQ7rVj/URDuzGk6ATXS2TT4sSydfFca+w
n6Pv+PcOdYzbhdDOByEn/gfbue/G8xADkel4IOwUYouPQQxuK3eRmdQCcLVvgJlC
1dCnNMwOHKt8fm35DZZBPESJJPeEZlQWoBcVJCpO5qsMvRdNYuzsgmckWA6eFHH3
HacOxlXoEzhJvaHv6RUmUfcZwU2N2tYlq3YjKvCMj/pvzHRTjKI0w3+SYeuT1Qvd
JM21kgyN9MxOJFgzzQcglvB5VOOxPK8gDrixdI6ZkV5Bdneyv6OV4YVK/dhoVNc0
WlolQp5KIiPf1XtBe4Rcfp4yK2gZMQLAHHxoYleUjTLn14HflY5HsF6i4TEMRe2D
ff2JJVicUbsGH4/Ci3c691Q15q797QMh69zXjmIxIYZ3nP7589+9Q9V6P+Rj+U2v
aPiJrOxYwaWRBJuAoFAhNKu544Kbyg8y/PGerKvk1ZJOLfWvr4njwVCvJV5SEtVM
V+j6mUMxDLm9PPcDRcw7mMGtCA3P1ctTKi+VevcRcoc4ho3ZF/J02y+cgvR25DFz
rJTjpIx34W9nQ5+H5oRkdAiPoQXojxepkugSYYKLwshVulvyNugQaXOEQcy+UYPy
Qrl1qPx78CaiREsNXG08v5+l+I9L8PaWyJOGwx9QUp65qnP+9b218sei2+/IZaYj
jwCTvph7F3qtJSLyJgJJN5o8eb/xYL3A5erDjZNGextHnoyICfDlvtn2UwZV1w4Y
maYLlXV5SyMlvEHc24HC2aQuqs9/m6p7va1XYNk+HtpOB0O/lePku9265ovfCUEp
5W6OfbJApYIoYB1wKUOEC7iv4eEXpdHQPicrGhfXkpf+3X1gkZwwpwuOOkiN/3AI
dWy/n6CBL8VXfJbI7jmA10GTb0Vdsm6h10gPyJJP7IZQLpblRsY96EPLrgAwv+tu
VTyWd3IJ3s2a/43hHXq7G8Ad1nDD7QZ1Alzg+GeMXIhPamym+gs7qt2liZbK/JUT
ECSZsA2+JbkW8a7JBid+AVH9vl034PBs89B1tY3zdwoXMsNirQvfgR32oDVMX28k
gq66gQ8+IvOp7mP2N3syvLSNrxKN+fkMwNFtR6plq+FhlgWcfRbMuvuLfnzoWl4f
T+jYIscb9FPkhltBVAxwoAtGkx2Pf9nq/PRthTymLf+O0NSf+MxNkipdyzpzkTo0
QXar0EAitgQpE52NmZzVlD1Y+LmWkWoNoq7ocAiO+rh/9Kq6dGgkQNop/b7SacNM
452fvPEI9H1ZYruvwhAOQM7A49x7aucW6kCcGPbazMtuH3ctx1czW1eLLYi5D7cd
ALVPKulx8F7mxTDrLSkYbo3+ZIhpyekGYxu1D5yiz08znQPpn9B2h59XhJaoE4s5
QgDDX59iAXKu6dGl3aROFXC2byPrYMvrhlyemfl5wX0GgtgBIYNM3lFHB03+K45Y
5IMi/SR+hvOxnTYkAT3KcjZa+n6ejA6uqv4nCJT95u9jKl2tWYJA9mfFUp2vqLU9
5gtGNGAfOCG8fdixI2U/a4PhlWxfb4dj+H6KEqh4X8Twy0gfqjpTf0NFzaBPlRPY
MwTGTi3Ag+ZCxfMChRQ9b+bC3qS6/8y6+caxiRHYgaVz3Wv9IIVYa8e5mS9RSUoB
2B4weL7FE/wWVezWzBxQQVF15H9SLZJ/JcbGwOdrDtD5h5I00Q4VcrVLbUfOMN8S
QnkeuxIwWSPf1ltx0HHCOTk0y1+ZT9jc+hEE/yApFV1aNbE/esrTgHCtAS+A0fwq
AMvWu+v8jPEcGItJjcKv4OuPzL+1NqQQefap1GUi515lxfWUYQrc7ql650TgWeWh
MAqcUCt1Ob4Vd0YXPKFumcSOGAN8NNU9kRqfSRfxSam8Zf6d3XK86EzkkB60t/Zr
kEQU54uR50+ZblS0NTEd+FdKVQs6QF1aMlVs9Xj1Wur9Z/ynbngoQ/y1x21029yE
SBIP724KbQBn0AvISf+XwkPFZLPm2B7fVyo0L7j1GWd1HGVNPmE59/moiOYYqa+C
UZIz7n5fR6mzuyw6K5mblYVmSM91Cw5PprEPj/uc54heyIi2yDEHN3MXVav4Xziv
MGqqrSJ5QowFR93X8Aj0xNgKLvbG5ogsSxEx8weCBorSslq4ezEnAhVB/1gOeUE9
Qas4vRyYUGD6ZR7nryDKTIR2UH5mTfDN30QFfBbIkUEHww+EFy5y0ZbM/kxX2Vjs
peQqMO6+5nHjKw5U/tMi2aR73F9DAkxFbqY9XwRDvXMRLOaJ+m4J0dqLQ7tc7Mw6
ckQVVHC0K9V3z1+XCYlMtGVjoSRfiCet1Z/YGFzFZf7cZKmQopm/kdJm2fli+h4B
5ydTD/iOvgmEAoLr2GbLP5lZRP0uBZMcpICNfaaiRzx8BAdI9MmriJdd7J0cxgKz
q35qfj70OgyBX/vQAUR7wrFTaifHzMricQLMrkFtDEVKU097xXH+mKvpxemtzMAB
0Pr/2EaqP71rYrZQAhyYofMXQTizGUSQCDQAwYOAGQPRkz8EbDetlFtI0vrWPXZ9
jVGwiqY6hxJE7xoq8XqT2c/AEmC7ka6dGbNKyWoXgjb4pEeuMIgKCxM/2NqMDFZZ
+TVAHt0xHx37PyNSh12BSTLsHlBH/CiXt15U8yIVh74HqISreH00FsL54uDrYBpT
o3eAqVbBF7G/2fZVPgiyvAZN9xc1oHboMWO8cl1LHef8VbtUPFhaooaRkeSTuPFH
eBLBSXw1TUsKYhmjuEebMg4vjvQq44cv7sdwmOXzGA4L/xGbolinMrgW47Zd5I+T
XDoJgBq6n+WA+wyF4GSDNdj1CTZXasHigb5At0iJ5rtJuh9MqipJ5ECMa/NwZH0s
wLQC9jn6603+jbBICuuX2pTDx3XE+OxXeP+z13wxJWCLs33HfpvM/ZjMXXc5MlRs
IEDytYBPqqUx6YAhHh8RerwyiaR+2co00niWVshD25+m6/wbreoJBH0XmOuLE1G+
ACCieBGG/bd66BNSECKX2gKzWklbp7h8GGgwFHV5twLqH54hNnVY54jQVsHO4k15
6nDuSkVl0AKmiKAZMPyAbRKlwWp/MA12WHBkVxrIA6u+nPuPMpt1yWct8nB9uER9
39SdjWVAQ6J+Xd91i1/aUepiTwwfsml8wUeICyKReYUxVyrRiDUBtIqPVRLdXuad
iiQWKHL9Bxcmh7pBKum0W2J2STnYDvgBFWhmHelbMhRcXynnBDRpZHBwQbX8BUlg
fM+SPhRvIfzHCVleFmICRy4sTaez4F/rWzaHi/kwpEOJdcryzsnQdSrc/xBweH6g
u1Dn9+U7Bs95+LdjbYS+7RPDb5IHSJq2yaNfcXue+OeUJpHrTKIHZ/w+kREB/mFl
UMEryDlaBuZUlSBlfs2wXKK/KhkvdPANyLa5UkaJQ7N/QlPPlw/9vSJv868f0eQ7
uR+tyxyCJy8mlqAhvp9vfVVwP8Z6egsr/uaOD73AP1bXE4DvAFngAi6nCIPHvcEW
P6w1PiSsC5nQIzW4AXJ9bapsNjSTTbinTcyA0rUtltSV3bAOtxhci+eKwJm6bIu+
yRVBa3RzjqkIrHY8vaXFYr6VOebqP/QeOfEbZngRku7lDFgzv+axdd47nZmcL3Fo
G3R7/jNdmXswOIdojvBSy6yqP2WZWMXU0uvw4DwqOkFn0A5bp0peCpNO29KxhmRY
OrH23r4ELW4aSnhu9DixcavgWJCWkmkWhn7XQh4c7t/lqFmKBvHLwmArZawUTl+7
GKg1NhMugM6yNG5H8OMS4vuUSIM62DEXcLz+TqcnTU5FBORuffp6IoWedZmSKiDy
toSw0dIhdVK0CCrk0ZrX/dXHez7bHmVDudatqf8iqBG+AUbdKNGTBAYKrEZHGXTd
6rnnl0gDv4LlgHzWqZfntTy70eEK4HOcFZouIaF+5nYDNMTcSrQ0lPoP5oGmPU1u
ReOyHXSpMAeWHrkHMS6HvxniL95r4shmS8Wgum9HlZp6t8NAhE3YaslrNPPV3eXK
QWeGEuKKQ1VVu8aYba/zrQ+M10hgIARIoqP4kH0SwDo2OOig1MzMs9Ao73Z0JdvL
Jd7bh8t7NBw3JlM0x+4B+KrP+SC+k6G41oo8r6azZNOBRSWey8AoKBl6SeFSYk7C
yAo/YQ5s+BGXtkhCjGOEoKNjDE6eG/5+GiR7srLNs9rVM1unEnir3aIpn/X5X8Fr
pTIrikCwDPXCXtT+flEIQHsE0giCrmZg0A/3izaoxtIPA8226JRuLVl2/DmhCv2B
/G6Q2OJXe84iiOTUAFCN1DS6vKhl1TrYVrX9FZM5ZfwkZeiDXU36B+s+vg2mkgyA
e7XLYFwaL50nzPcPDcmFJ+yxlZk1sM7ZWxmSJJHobd2qxFgbjHjfPOoK8tAArA/+
0pWS+07s7UcmVTflf64+7iaS1bVduqZFFXIapEHoUqDm6LWgcKdYeztBMSHubejA
CfFV+d/UwdAb27LFES5VfyOSsiK1oZlILyAzYeE4FpS/XxcBcnk9fexLruBKJv/F
UQ6pWCrnISBHUaK/4LgVyaraexkPHNwVysRso0QNRpbJUiQ1b4oXPvIGBwGfFMQp
uY8jECwHUqoXD/uGstQs3vYca64uGUJDi9bfaL4On6+PeRH3yCWWjXMpfwXX3JzQ
DbG8R/tDa8mxcDhqDdfSKNNOLjxVprbq5iL8hIgLtPQS7dQf/KW+NxPRc8gNY4gJ
OlpiSM1XpG24DS3bcSHlNqZhmmgMNKiPhs6toj4UrvlaySTDXbYl307xTDUgW4mK
M5DYvRLP2deyiDqxHPLbawELG28WiC/nNnTDnhV9Uk+JznrChA2axEW0l01O+mh0
8n4UD2hwlScdMKd7/ES301fncNpAeGY3mWLCuVam/9/9URHc2ZbgzSVrgI02usvs
Mvc1UlUvIrFR34FFQWCQdQGjrRaKMJ28mOngDTEudBy4Q7B60ZoOm/qiWQhIz/RV
064dqj1TsVy5Il0MKFi5fvcqsfqQMzejKOeczbDgoAVd/2suGeNCjH1sFEeXxUv9
vZ2UNQE3uHLf6WBaysCyQwVCP9PV7W5jhnfon6ce/lfnj3VlRnXSYR9rp6yjGlAZ
jPqsaBw7T+knObfsGw7OBC8u8s9jgdZrkOEBIHi4H/48VLRSDMbu8IRKP2Id8wY4
xrbIf9d1LxtRsAKHIVGhhV6XP9VmmVaXAVRsenqpyztc6DOEGFzD43oHapYeDPhN
FhoTi8LuUI5ffDOHgkjuKksGstZ4Itwb/YaaKNR20SHY/F5+3dG4FMw6i5Avlhts
qpfXrW+BA6S1OB4mKNLE7fnzbVWbyhys9kve9IMUsceDZP+SbN/G/liWMOYpYlfm
BwYmNCWkNLfJamjiktsuFUfJHyEDEQ2G0A67Sm/Lqy5b7U2NRJBAE79opxGRaGzm
VRNhgJ0SDwU6Vq6hfEzUb1emYOtggnJXVtHIdCshDHQJCwrBribKKq4yoyzqmYpf
mig5B/b1Pwbeo0dKTT1GMmZbHgxF6XofLqFooG8ajPi2UmvMNZBHrSD/t6liWZP2
xHjaa7VYAXvfkPWGSsKKFgUfbsDb17x/G8PF2utSx+bitI5mJbNyO5sHZ6fsapLh
b8QdGgYbo7R3lO8mWGFxh6+/8u/XG6Quft/sa6VZbXC0wsXR7V4SYy8Dr+eCTuMy
hZdXQcru9kyDKYR5NUGaaK31r25AjmIRMMvsAN7B/UUVbN88BUz0oy9KflsQdncc
e8cdKjMxwyMPG4lkB/E7jeW+2Ax37+WN8GQNV/fHlNvNlnJEnnsswyq3qbHkQHRP
6iZ55um0lHQIbYmczoryfmJM0FpShl4ORgcroN/263Ov5Mk3IuyYmZRViBTnIJWD
2MjeaAvWpnsMuOhOQGvdAyhNUnZIdG0BH7g+AtlcUy7bR4jCUCbY9fbQYkUDjb6D
LiTJsl/BNX7yROtisn/H3CLC5DibrCsZN6JRD7cHZIBW21m9ozAMrQ/DW5xeUjz9
YdRUFzQoTb2AczyHiX882djlhgnYnU1v8Go1+K0PIY+g/C92Ej+n5BdWsBnutmDl
AZQvV8z0DscUyv1YzbpfQyrfXhtxjPRG2Nxj126QDm68Jzs9Dau+AZ/mWNdz1mQB
2/oi0xUrctbaNWRjtQSszD9XaU1PBSECKuXwUq0L3iOxBzVpQ5XK30oceDTxZRrh
aePGHfK+q+Rp7Y7c4p7NeZpqaBexxyeENDfpDZ7q1cBknoRGF2iW5IuTUzvdGcFS
FdTQUnFGtwYjNmadwzY05jW+5LeDypOaINgYJhKzUkms0y+0hD4V/Ufe7+bjxIG8
IM1JbHeAWj3kQt9QpQC22mW9/M8v8f5SMpTNnGGMiMiXRZVOFQKraa49aFs8jJbv
68CMJNDxpSsh/iiBLsFH+KNoiclN04vkBujnLu2+nMJAoVIOMauf+1+EZV7EDBmA
zbqfo2u3A3SOtLn6EtxOIuzxTJmG/ZfG2qmpE7paSgFIOWw6A0BXGSRaKAaIgeFj
X+4UQ/+lWXmLOl8O/e31ANFR2AMXbIQkQ8FhDWwihGTzq3QCf1F/l58gZnbL7NaP
3tfY9AACXhCCy4iY2ttbnFiEeiDs0PlR1vGylZ0jiRtfsFFYkjChfiQUpGhSLQqT
nzG4K6sjkp7bo/Uyt8YsgIsVbkMhKJ84v4Fl5F56pK26X2JyiJSCgJVlsPSji92i
RdpvCXOkty4gXnc1EtN9bU6FH/AsKGCNGSli2tYxDi+++Y3nti+qY+shg1oj2nuQ
IwBO5eKojtkqMA9ItdRH0ebRMfK6h/S6aaMw/b4wuFCy83smrgUzmJBr5zzIFEtN
9ELLAIZeHojk2A6HqANsVYQDfLdFEx2TVgaBbrQYWjk60Mnsv+gd5946QM2ltB1F
D/eCQvfJadRa4gTDHMQ2br4453mO/hhSIRwjkBQYd0uLYw5aMOqvu1P+nHgmOFDl
h1XNc/Zf+w1bQx/LSfgfrH/3owuJ1VrtiFoOBXaKSQ8MGMqsJA7hGf3lFwa4Ty3J
MAcBlgxIibSS7IHMah0l9LhKKsK9M6A+mpshcrX3h17VkLIN5bPp0RJ6fiIPiOM2
wXVDX98nJKpEak6Mxfi50KleGvifNJ3pcSU8GBaiSGpWyG8B2gU/PAwGXL69uT7X
aCgVLZ+CYWQjRDyS4AOQn3YjPki6dhfSw8ThAjf1iSMne8j49RZ9GO0oO4rS/Hkz
7J8FMK+2NFJlf3wmK2c/98NaBeM2bqVacGKNm5HsJHjAVVpXdOq8zA6t0gHf6sPz
7oK+NFSHjWIZY5Cw9/0qwbOJ0A8hMIyzlcagSmnjttDRKjiMRvT71eXC19Jp6Eqn
Wb9TZqtS6RY+m72g0dPS1YLVHU+4Azw3jYZJF+uXJp0gSgyAFt1hGQHtFS2u0Gwb
woBVVysYNHpg5A3smE1CA8Bgee3zYBl726T47QKTqeP9cQm9Zevx2WXgIqgBkCe9
rmg4AVIvMCcIHFEMNcWvJlZwSgiqUcapVEe4O4rPh97Nj/ensdgw35EE2XtOD/ll
kryOcDJ/Ff96Z6tyomfVXenMiflk1EeIE3CeN4uhv+M0e1+uvc39WOz8346qRno2
xQjtTkCIwKMCVwAlTBp91Nk7e5L0dNXVaSjOqGiRww6LaBGK60lm+ogJG8YPorJK
11r4n9FZZBtKgmcbSsleFDZsOoiXANLQRu/P3w+vyNfmOkbHKNL2xiYqq0saOmRu
pzkcgoLn6VR93GKl/+yjN4k1IDkBjXjljRXb1erBYyD6xX5Pkug3qKkGRNmhRurN
QICAb36J0kKib25brLMeLaopNvQONYvwFwJQxR729jn+e3A9uruWWB6n7fVtU1MZ
EgYgDgk6wpsPsCPc9KzlbOEhgpAm3Gpi1kvx/cT8pXWoP41aIu7L0DElAXQOtRRk
VVPsVJZUUkHh4RpZ51Wy0eGT9DstJmENXd2cGtRf4zHHv4mjpNjbmgMeDawccOey
ppEn0LSa1k9a0X9R3lCr6mekg9xGsTFPy0pSMETeOh0p/ZN+kfyR7x/Lu5X03AvT
S3hTw7y5T/TlAkWREYhC8baOs9mJE3jEUHSMkKtFnJF3lJvUwpQnGpJZisvEHxDx
O9mRfYIN0vwa68AtUh/EZgmRxxUvyfyXWY/8fUA7QszOo5mHCxgDbjNwb9zQ9cIG
t3fPauv8U+WEWKL1cL76HdhPnpn86mZTeIdRdgEUF+hSRMpleJBd+JgaqDQUDwHq
48NIHitgctyjARiLtLWmi2X7I3T5on0QhDL8prjcLzo5kiRygqHtD1bIbfj9kw2F
bIcacmTpFdBQMmG3qmM0NouxCyO/+LMETRDrBGO//8foVdpKLaZe5aHMD1o1nyrQ
hYrT+r+rYC79qfgTp3gbEfa99pZjw8VfntA6saQHRVqCYopA11veQ2AOsaXSfdD7
9khIWObCuUCR7aFmD7FxxlkC9FDJz6jNJmipJjTNMnMNgqBUhlb60G6K4Efcw65I
1osa407wpziG1oYstQgnRF8lTX40vzhGouUkMiTP9cdNoFvujIDUrZEis5jXCY3A
6iKQ4ojaWG+ceJfc9x0pvy0fWJhitfy/aORGvzeySJc8joovWjGmQBhGfssnCC3g
Zq7z5YG/eivqgD33sEdzpX0V5kF2NkZ5krysGzT8ZmJOOtsYaDa1GdQYromasqxw
s+a583ohhCKlzx0aKWXWYOwgMaGWOWEoGXzOZd2rOIGYpV/3nzugI8sVSM1Zvho4
6qKGMo2iFYlNUT8VzPjMqiWRFELzRanRXl5ADrtxjXpx5vZWZw2oyMf4gvnQM444
pSJvYPcCxD7MjoJ/qX/YZWVCyAjqtf4BzEJvrtoTKZviEWJlrkkORDiIpcyeckb4
dnGEpRxPnXSqjcZBE0m6uDsGFwxJ55YsYUkfsIaDfmaT56KAfm9C+DwyABfRYrdV
r5hN4CbCwnUW8xFUECsLIkYVuD2AXJuovSjVFoDBv0+8PUl2CSKMIOmKwibl4CUQ
oEj2dssED7B+UcYsGRyXGKMcj8Wq2V5n6YzCoVZEmhEADnIdMmXrLQzxudz8HEEs
c2k86okNG0RvIf8PWEI0KHsu+L2uktGmUJxE/wMpf30qjU5dRqSc4/gUXoF38mjW
+fPJ/+y22+8LJsc9VrfjO3CJUPJWETgGznuHg1gv1+uFPIQGkhhhcMzrKxLE5Ylp
ZP7MTOPJTTKHgpwwqHFdkDzQl+n0mb65xuHPPRdReXhy5bzzxOebDPf22bafjWTn
/GwGvonbiIj/4zKRDG9Vv/mYc+gS+cuOoiI/K80r3wylfe+UR+J5JwoN/HGED3Wz
PT1wkUgP+vp5hJWAbeS1xBD2gNv9Dit9bvSEidUFGVW/pxfu36nOwsKDHS1yTS29
8n65iQ47pfLutYR3L0Kin7pep6Is1PiMgDlzJWv34ovvs5A8aihre3npBc66t8W4
r8ltWRB6kMfinwD1MLBrkAndlwD9DZW1ybYeaL9/gjYV6rHVsPE7SCUmsWE28MAO
H/Wj4OZ71wLgRApTFu37JHNNv7JPOtRMvzcYKL4neFox+vS2AvniKnh/M0N01TbR
JfzAXhMao+kxLJ22PuzLyG4Lh5kh79pyLsv3AfMl1+u+VMSPQlNENbZNnvAU4CKz
uv7NjrBuYTSNx0cBN7vvLgPqhmqCjPhAhIcBgapqnWxvPNFmPmuWBBZ8UWb9uFTH
VrYt+RnF93vEFx63xoFszRHQVAZmKmedsTF8b2q80VbmkGopFIxGve8SfGnir1Rq
/FIunXj1g2B+sYK6DuD/wNy7lnZ/744PQortajIIYIHblpsJ0XmFFBYOwKZdLsm6
SYurP0v1cNPdOq8O4ABna0ns7AkhWaXtLoWvswr9eW6piwYv3sTKRY6i1nz/imJq
/e0lQFkPbPgCnZ7H5A4L1jYA0KihzqkxjIuwUUyiHn6MUb0uHMXJm7TyZ2Lwom3R
OmFf9lbT4FEj+d73aTrJb/Gjze57WjSx7ZSja2dDhHe3WJajsiTSt6bwTkEhuj9z
BBbE+Qmpz+kHNL/HLcfV2fZA5jjmn1ppIoS1o3DfxuERYWvGDhg1X/hM/Mm2MlQp
d66Qq8wNgrK7zxPifJVOtnzBAywc/4IDrtaHIrGB3s5cFLAjwmj6zlZ60ltHrDJZ
MYUBZiG2UxmjNJ1d3TRjpB4cJ5oJZUh8H3Y5X4s87DYDIkY708Hn6LMDO0nhnZEC
cVGPgawjVw1uH4CclueUb88hMk/7mbZTFck+D1b2qVaC202L/kyaCyul/kuka6T1
FLiXmRL8dcvuIUqnrLjY0uTQanfGmlPB2mMMsJewt5U3r7bXH2QUIFVr5PepFw/V
olEjXcioXz5Ma5zGuURERxZ+FWaDdOaFzJp776VYoLAeFj5e+VKJtU9s2Xv80Jsy
U9vcKZfyZYbykWGefdZiaW9qOFfKftzMYOOdl5m2AJRv+PiTpGb/jge0uRSNwq5c
l/bm8nFgocHm7ntRYDyjmJP/gfLCq1RE9+AK1Xte7hAb8SIMGXPBwEt20cT3s+2z
r+0em9eTSiPoNfCsOSiNFfv83fJgyBiHXUNSm3HhbiJKwtvBwxuhuEUdwFhsixx0
jLKRd+HCKYc2+6rHz0a1Nq2sGfkxNQPMekjqMxonKvduDIE1fbozqEKPCYyesNuG
l8CREVm5xwgq637/POMhl+pSCDm5hqoEiBfTzfJD0jACekVTgbJY7GkW+n4XgUMz
P5PHeJTuS0ygJ5W1tbHfd0Z3fdomSW5VV99ZLOc9I9w588w3U31B8MEZZ/kKX8Xc
FvsbG0PULfLP5DpSetIYuFqpFAzRCzLeKwuN9yoGHDQcN0PnPB4FgJatpyfx6ODP
nPWX49LICEGs/PuqFahcjDCXPb1Sn0zdhXUrBogVFR/Xtr2BQaLM9BMPONkzZ6dS
UqCx8qV+4dU1DQxacVskIcglejEvAS5y82igWJy0KvwZ7MQIQyuFmXFKDOHED2ui
EajXSeCAkJBk2rNzgKpcZGwhj+bpc7E1hTs02cXr/7SBS1FNVG1gRuDVJjEMoJKs
oXu9Mb0Iyo2BVeDy2p1m5dTC4ccHOQRelt0bT8vtEgGwDVgf5EMBpsiPGm8aEltu
oRPNXG+m2boICQUFIs4RP2Cd3R1vSM1E9ffWFyirCE8di2VI+glSXkKQ+M6+GJ+I
Klcr246/6X238KW1z81oe1k88ivmre1eouFZAf4L5bCHZQFrbbBfjzhmDFW2kuDV
NuQB2KlRA2LXmgaLQYqUQhdYn9EDA2jFBLTIjdoHMETAFq2+BYfa3xy4ISJ/cTWr
cka9MBW0ednas7sGwcGjmUacZRwLDOOfGxqlIBbktLpADDbuuEQrq5K+9JHixyTo
J9YwZd5x5kwgkUc/UedyljOsWyVW6aLR2B3ezYfPhHUa4fXiFdeZoaMsHwA7kGjt
qLJRQCXvuN0nEm+tso6A6Sp/WoMVzIP49WKgltzMFJ4KIFq+DDwrcibWPBYcFkzj
Ux/VKugH59dwU4DjA2OuvXL2rz1kL6TtvbxktIKMAZuiUuJsD+MM6+xIxpuFKVaL
FQS26cnVVZyTNdCnTSjZTJ9sL7CNek9zaYMyv8nx1dhkZjZI7w3txGPl1quLIX8a
BmYgr+zV0XKAECh/NurcABvjxftlDNuOq0/w2uyfxAX/ZLqE7aHze84rbZsvQfoU
LasKm663WvrWlqovn89SLPih+3ukYW/A5yCromfWrpxZHOAv7tB2V1dqBfEzjrGK
abk/dGkZRUytH+HmTixxNbrsaBDLE1IRRJjWBuAO4i7JlSZJ2nYY1N/dW3RfiXxa
IzYt8C+spmtEpWmb6mXVqYsU8b9gmDOej+CNzJgEBwnpFvZuDJgNApxT4o46riA8
jytLcgw5Tgkyk6CBU+13JHO/zVsb8+eVlcqNuZiVliNasxUA/4oHX/4oUhpEOJNR
iGWDV81JF6+HULipbuUIGZO9UFZaTXOovcAPoqxUXE3FlmqLf3yA+LiQyybPa0tL
qSdP4j6emd1HNpzMgHLek4R82B52hYA0SQImGwgWmsIWHtIW/BWUMkM11vLGVivb
BcDPV/DrdSqc30fczUV3bNQHYD3pdsq62ATVJX8NOPt0KqLgLK7jpHvWFuv3bLj7
LL1Qgl0ybJLsQNhJRgnPgXhNQskdnl5rn0u8iDQBM1kpX5gFQ1zB7jWgszetNcjR
gjsUUfiz/+HhBek+1q3Se+PepXzpHAP14P+bfDHrJLXTFxLU/vw/tjPep/nWQ5ZV
QsK2D+f+0PbawFfOmBOG/NbiNXcrpCuZnD0IDzcpvq9pasbi02MGh4vIISWNj8lI
oxPKvxL/hCKGE1iRrItlD2n/R6/KTcIXzAFi6X4ad/S7w5H7XczdxwlLO3OraGrh
lzf8rxTnwLv6b2AF4/Za6FRUGlIDNIU3ZgQ4TnIIjMnlNaLcapuAgAF67VlZe2t2
sZDNxLP/ykYD18llgTac6QKq4K1CCXC6AalF4UXP5nFeNTKFYsrbkmiV6tlQ/REc
4dR6L7V14L+il2lgx2G15/Qt8+lHE6X1b5lQFlGpzXQGDtCP3rJvhkIdH1cvK9mA
LtTLmAX2BHVwg89OlK72PIWBsumk9k/Nb+L8ZBZyg7zpyPRZyDOpeHuT5n8K2sHl
b/VjT2B0MqhTKdKvjvwyMdi00sZBN4u8EJb2wgdvtqxPIYY/wF8Tve6bN4x792yz
r1ZBcuxDhM9NPYfo/6QUM5Re6nm1bsptvVd1N7QAxfv1nTaWtZjr/TImKFsGdkrT
uEPTD2kbr/KaLUVksoXeQFDngN1EEhgubaBad1ETMgYzhXMj7iGDONq32Oc7R+zo
RsPSpm6dcGnmc0OHkvlagdTA6At0T44Akr3j+lLgJGO+rg/WcWzv17RkKzEKkWW7
F5iptglgU+baw5f1nkpuxyHBB7xNe47lK3ZwZIQnlcuC3mvAqAneNYtOJZ4L/Ixy
ABpdPeWrk3dPmgW4efB9iFua694AvWcZ68s1Zf77Bb1GO6Y9JpUe1VLgzKcIc3FM
FhQAPUEcB7wfrU88YOVA7S7n6a4fDeU1/WCo/iix9dXBW2fDWXDoBGw3emRpCIjn
cKKhaDSQSnXsNCI2VpGR23TwGcl+NP03ko48WDe/8lEqBmp4JydeVyFYBghEsvfW
+HPiUzN85syI5NkpLv8JVWkWhSl3F/T9BGyuAJi9JjuovhaGmj8EI8leUv2+IajR
DAuXhKKVmn63E1ZfHwn5Dd7IrP9HPdmPlreU4Tk3NtIaf0D130KCMmc05Bip2Khv
jxAw/CzsFK7fLIc/Rq7h06/LcSHOED2fWR9CPa+YoWhKJvlDHmqUVfrTnjC2v/kn
KrHXNotT36E9nfiALFZDaP8UNxak3JedDVxpo9BghWH5nuTiIHfZxdPxwQBq0oXX
GCue5GyZoLMvrmaNbnbKefNDqcZZApg/hMW8dbgqwRWy/Cw1iT2LrpomPKhWG3jS
SxtXpbED/+A+H4LwIYy4/wykib4ZlqFpPDPcu7+k9C79vH3md2iYCw6gFmH/PxoA
A5W/vbxYP019BHHgguyOhHOGjbup0qfrLVznSQZGkqW4G7+0ziO7KulwiHQDhYHm
g/kJ5pZtXHJ8LQr17WsjUEWIMxPMoKc/sm/IDyxEAOslxvOYm2D92QlE33xfgP8O
mViEfmBobGptLkM25xS9ezyrhYH7p/4U0DJqX+ds/8iBfMgzvERTn7iCb6rsLpZT
QebHDotpUOfISFdbX/++sP5cZ6Xui5zp5bNLmW8BTrZDHkbfnZAtR49pBXxfryLf
JoG/uapnZQ4o3USv+V8riX49meC4JvC5zowlxRX96v/02xAeFl2HObL3sE0hgppT
ti+cKz+2JGj5DEsOwHeM1jRw5z4ipc1tiepcwh8IB0+P22nCR0PwF7ydIP5LVhLE
xaRE3cgCfl9v+tY4ZLNS9dCLwIVDHAqIxh+VKX0nA0Z391nzF4LK9btRwaZWu7I/
+2g2UNRENkuyYAEXYnjecWgs0W0qN2IKMbCX7JS9KRxEpNZHzfxBUOFg+TGeM8Tp
Eay0/KuduJN7IaYhfxf+Yd7uzlDiE2Ci3AEv5TpcpsyUOPeHWFVDIWT9CyYILA3i
RI38FSS6NyUmamciL682YK40YVcpXXOURt/jVf+ymQyR02sRX/ISvEP/yv4gTg/0
Se4OoIr+smrKL0Bc6S4wNbKkkJZrPTfIcIdn0nhaEfGAh3GpEMq9ibMvWUXGJHBO
g7uZQWHantw56QkWBWrIHKgQwsc80/39VAg8yjS64GDWONZwJrmRv9N8/mpf3L8E
yJ3OHyZhoFuiHwJXgYznLcvaG8ovIBvnKdzIr7oqUvnedZ9rwxHVLAF2I4KYhAHw
7H5ViBHGVv4dbdb2QSuOFh8ArDqRZucc+60k9RyjjDFcIECxjmZPDxtgQpawspSn
5JUUgGoBSlyanGK5dVBdx4ylZVYN9HYVF/OuB2MjqEbbGq4GsnHQtMiADfLfMaE5
vLAdEd+C7D0aJr3QWtnSLAjZVuiiL9J83IMWGXTUIJDGJp/4YrKPkh1taq7zb1Hn
eSyz3nGYUS34alZY8r0Qge3aM5QIcgh2qrovBXWVgXhcJDh9+G5Y1cngDDVtSAF0
X45uCH2QEj6aKJXR3ts+4srJS79WTpnlDtRLefaTM03QphQVq7o+yAwjewjoI2Vt
gIOesQJapk3+4UNQDNKcjDjgnG++81/MlkbgGuzm6HeM301gKSkygZTTXi2/7qzd
1ZQ05EAZd8bL/mLMLB3otryjxtwc2nxBZWG5TQmbNWtey6+EC4upB2701XGDT20j
YI77881hIjxIEn/EkjnbYyEFFedzBu/4yAMbW2WyUJZU8UBtyhpsvZqPJksib2FD
XJcnQpSI8KxElngXDRfLzisHnDP52rAOdHS3YjQhE1hHHTEoWnvDXU7n847skLPr
71/o9iF+77GDOlOb7/BXLuDroAZRPTB/xNgEp4GtKND6lWXGt3GUwQhix0vcLgnG
vt694x+KMA8GTLDe/l5VaQYLePyBzm65nxUeVZ5Os6L6++KRn1tGroVtiyoQ2F1B
VsNMxZehuM+JG1gayA+rfRLWjCarFoRG2vMkL8V4e7j4wm5K8Cn6aUMGzbR/VjF/
9lj7NR/aaF9HcSVLxhfRPO2BXsK9gpwvIBUbQ51bLQewkTMWTZgwqzKtoaF6z/xl
UPoq4eJOkHuhmXSGLoQ92voZXTMKR76irjJXHHUAEdY4eASDbvESzRCZHryJurQi
3SHJBNg2eIzxZyECCfmSk3I1KcvJ37pQ8SZtjxcVYRLY9lw3c9gImJVm0pGxf3cu
gyqKBAg2BQKaGUOMdPFQUsYv+RHaCZ75yQHyNFKAOJHyWn2GM/IWgABxE6KWvlIP
RhGq0Xiz6rrEO33E2kLhd1OfnV3gp6x92nWirTOg/bqVClgFvNQg4srRALXpSMa6
07Pt3H6IzviBODB3iqqfD8yi/MJC02Ti1Xfd4zBJEMduz21DQYtC6xkrnYeBnR5L
FnxgyOLzlRHJdZbN061h46hezD+IuaPN+28ZImEb/Ep5Vn//Bg5sP15cBOk9sbbj
MS9PPqeOxeJDrXB21DFhqn1JxsuduFwu0RyJeRTJ2TSGR4G+XEMYlyfsYntM9n+L
qEMSPWQFXz+4tX5k9GiLD6Wr6wL0TyQvzUHn/zjR+yK/bglzZNWVXWE52GtP00AR
NH2gyyKvw9MAN37aXf2RNMaDj6+pawpzQpqd6/Ky0gLKuQkgFYyZvFbG3zV1JpIr
+2UUFG2Acx5plvSX+jw/uDc4USpC0Nd2br4f4ZTOT8kPWbSpJ/1lMupHhMWhIxa6
9AtZa2M6DSZJHs+XzmtHYNOB7Ly8ExrItJCZpjxyE+CiklolR/5aKGfM51nVAz8l
5ptR9MV7Pl7gLQOtu56rBSQZTbP4NdBnpj6EoXND6AsdZLF/GtEGODZatnCSCBgY
irPMEZkYJcOOOKaFzs7Kt8l8Z2uZnHUX87Kfmx2OqgHY0r23ZokTAz8t0I0Z/tge
+fmrRe7Dkb6pewWONSyah8gF3ObWyYxSoW1EyjNo2m8f55qnWFrUwPQzrTZLg/GW
yPprqW2t/NtXdAnucI18W3hBjEFekUita6WvbxAcOBJAS9y5JjQnVv3ul0AnASnl
sqURZz/cVylbRNbW43+o5Xe+bIF3h73Zb4zuk5o1YZuyLNxsHpdnWpLUvlRQ8G5I
clwPPI4ZFpQAb5yuoSnc7AnuMzo7FxaApsdU+HgQixkXHfWaAo+oYuuZw/khT7jA
+j02uUKDv1jTpNkp/loEVGJB+Dyv+TAqi8AiRnnK1uN0YltnzVqGxp0l6TfzwdGL
+RP/dc5XHm8+vizLPjcNrIwm99pWjlt6RbMod20YotG6l9VpD34WHG5HQUVR5jV3
OSKOj0aVR/n2pX+Ls2Cbs9USGogyPBDns2rz3jFfHBPwVgE/A6XEhA/0vHmXKicm
B9XdQ98vHVHphPpAUJ2E84HdKBMoW5u6iYRHTTPXZpnjQCzZVRSmeg7ruhfjD4r1
Uf6PHx2ToaL361qHO5ltK8FdEK+gkRbU6qaBDICE8G8IDAKjmrgFIf4kExh5HTwH
jp3pDhzC8MYNILsAJN4pGhb48fV2PUZRCDM7aKXQI41uuLSc6uHMq/2lE9OG4d8l
stiuNorHMVcdPaXC7mrQQ9fz5hR5f1PQSHu5hYv38vfvUA86uCgoZ85ZS1/HcB5f
JTWit3DcgosgKjF6sgY1dv6ssVO0iqBOOlCIGxqGNgjFW6f/wzNlgMVKnaibmaGZ
b1/GpgDiL6DNppWLL2xBqmGaowZyLwVa9dj5Y9BtGh/0NvMXWl+hpCgIkxUuXlqf
eogF+9zQmxBllqQrZ8Afu/i2Ry/BFqVTWB5VCFlsEDhQfmyhLno3OEEZZl1VFoZi
sRThvQO1KTr/9BttCJOU5VgWJ5ieaoZaGpu9Grthzb4YAHT3IjnQU5i93mt4a7Ei
+rj8HFrDXMrZlPUlFTXRNXdQoK8W/2GA1+ceyVcGUr7i715l3p3QsHxfgs5BkAOS
h7Bi3SWOUt9VJcpQzJHT2/Us1x0T/hmChgwHWkyFp7c0BeI1JFMa5e/DMbORCCvA
gaBskaAOMWuwTVk3dQZlrePo3e4xiEO5QGA5XxJPjNmO4ILTkXyKfHRzeJuif4Wi
m/YG/QAvbnTTl0Q7AmOSIWkzeR6GiFIget03oYprZkdf/TOoB91dLBMDvrkVC4mH
+y6Tb+ZhnR6iGtizGgjQ0XHPEy71UJMafBMc2b5O9A26uGLts6lI2XDuA2e2iuww
M2OCP3sjO3DOpOhczxDjkeyeymSEyAgbUVOmaqLZkHX+Dqb9JQcQrw0lqIOgC7p0
x8RPWd9Q/Eldm8rrCLsKQZw/rvnfQII6b7FdwFCVwz11L78YxWmC7ahoK6k4irOS
RQj/5yW9ZN+TQPLfD+3zhuq7z2ibyFZLlsQViLCM+pcN0uqLScmW5xfJQJqILz5Y
lfavks9XBBRFuBtuaoNCMQXEFMCalQw3M7o88hhfdFYG+ePWDRt7+e5WwO3J6fEz
+zDV+VhtVjFl145LhUi45tgWgqLgpTiQta8OvpOhSYYFRZ7nZ+l9WhCI41JqCw15
m3nMLgVSCJu3yP3cwpxt9df+KRa9cQx9MgM57SF7I94b6cy8/DjqajxANJgbELG6
ngXdP6VyYtBLkhoeayLkqG46ZUuXuPnblHPvZxhEZ/UFB1wT87NHISSJ2g/39jPL
3TgFP4MF2GYTEjkD7n24OgNsGc44RyBixPf56wZ19HKZ6046Umlz0A7UMPGbbPqy
i6N8BHlIunT9vEQR8rtNONpJt8LzT+BZmWqyavxf0hs/q1Fr0k654aFZ1Ok3Mc34
1hxDAhQj8cWRgIEUzSYPYI7KZ9w7vQ6Jc8OoHZzjPnZkY1Ynd3fZ+gs/Poyd3tnA
C+YGlV+Xnj6jOK4wbYV9bwvTI2sQpr3mZjqWzNQ3rN6vytjNourhEZ+SInTNrjiu
VKCN2SywcoIio1i7M1siKeih8xz3N/Nf2SBfpXYB9IdDbYCmSLGr8Q+wKLk8wg+4
R5Y+VCiVII36IaAOJRgf/Wj9Z66bbKIsZLX7EyTKOnncZsp/bfmb8HXB4ZIyoHbO
XlSgdUstGIl5taqVq2ukgf31+RhhCD2HKCfGGXEUocRfl/oacYUT0Li545oNXQxz
tIHU0ksW6E/l1kPE52DBpjaPKuvAZLdBRxHyT32l8NQ1Ds7f/yKQnxeWpJ5XQgrL
zHeeb87pQunXDnLNfA9JsTOrUKjifAXXxFl+KO1QfYYMXnxjMrTjSf7pN9Nt6ork
x2XyA9qx9+GCRFld2870KNSaL86Oq7h8CUeXqJYZdZPQBx89M/UmbKGjkcSg0Oa8
KZ28bOZ6mWn136DfLpsdk3xRr3Vs+phktnrs8YsrMXSzSdSW5OlyUgBB6t3+TJg/
OrheE8BsUhLb8eqmPWyAVhwBjJVp3RFRaRFUHSb4f4a4NIPi/EgCnJBOGEiqwwCc
PYrA0SaeqaXSrYWQ79ixx3pguoxdP7qtWmqMF2HBKH8+tZpLX8P5u35u9sxf26fp
STvRJGjvSGDQwO8uyM1ffw01abBV2Nf4s/GhXEiRClxazG5qS07dLA0D8/6N7oYJ
XfZgMNh8xmNvcb+OcgANoW+U6q+m37akAa49x21TcmSvfUyDwQZbeLlQuI1mAv75
e6KBgPFMiE18V3JvA8i6bgdt1kLje8awCj1BaWpU43iq0k/hb4l8iSyhmAPvXUjg
6uR5d0MwTssg585QOZR3tjIzlVG2rd5NK9RWwlEgmRmBgA0jjRC6b9tygZyquuEZ
+nEDvmosY0Lcag/K50a8stIVUrBuqsvEijT2O05CDm6pxuyrfXA2Lwzz3UY/QMZ9
5tlka7C7DYnFCLiNuQv1so4plmvlMQAJrxXxPmsshvbWk/tzG6hPMNsJi7ev7lAd
xxIIFlG5HcB2u+8PG3EKTwaq3hNxwy0bFPmetDGRfVj9NenYgwicsbMF772J/WZj
Bp2PCgUbgtu5qf9c+axQvCKV78WpPUcrbLlysH/PCnrR/ELdyd8j4BqRi8PPtqgs
xkEw0IxpfRn0Cw3s7EeDv7fbM5g0Y1PBVa5ol4cl45tKp9kkUfepQD7pEwgq211K
jFwHbhL7mCJHdnHk8SfcuzHngmlKez8Wx8ho6Gzd9S7+X6KPbr5izRo6iMEVN2yH
7a4ToYCow5eyJbzMdXTJzqG/+7/AvijsDBZEHQ4biMcMcNSuReyr06ZQZTnG4lwK
t8BEpsXJB84LdODUfzDK722nwSvBeh1aApmlhLF2OHSTy1Tkj9aQKse7luVWCYiV
rVuxZtpytpT4BPVjA/OQEM/br1a5e9c1xwrJeeIK7GkTyL7u5hdAofoMhS+9oL6l
X5xmO4D0Wqi4hQvHPdpg+vuhr3DvZfaUvT2t8BIZo6fbIiJep2Z8V1P2Vbz3udHL
3VIYII8zHUbJxnUVzGeMkBT+Q2L7qtatCoDKsAvnQ7i52GFUEiU+NzO75G8HlYzQ
W1RjvkpSZazdRxskb0fwGQGpqEu+ajNaM+B1Sc328ylntu5sg7jDOLSe4Ns/gUkS
pNw6CAxPT3KqWkmYKZ9ayg5Tk0yGZdJc5wwplewkMfEwwGgn57WS47ZU22Rog4wH
ycDMhyLSh5Q83skYjhpxoZWcfO8cdrAr92CYSVb7jdgNtuSJM+ksEmWHP8QuNDVB
DjD6i+Pa7uXZ9Kx5E3rpB2Hvkmeowd5p3talFIPr0on98/VqkAfZL6d6Qxm6aBrV
0Nspqv/zgWBOwzmGrSLewqIp60EZwHC/SLLL1n609yvzFhFAHtweAJVz6iNfs0cC
isNuqlzfbED4udDkMEFiWmv2yS7WdpHSClWR8YZPUF4z32y68Y33fVQDCSAK+mAl
Q4aIaeP/XZzIhtOdMB1U1SXN/EHka/QTLzmH53FWGTAkQ4KFaa/oqDUtxAj9rYGN
ZMJA1+mN34bD6GfSkxLiWeUHDEnarrdF73pg03sTZA+XNvcuU7M+s0Qc+ELYty1Y
hdssM1GVLIirilgUY/xde/WJ4X0S8cmrwdlafvigx/d/zWz+dsL8/NDeG8j+uI04
eoeTNfWahYhkBQl79m6YnXy1VNYYfoKE6IsmeoIQmRva0lGC7acuFheESkDRhYiL
lopjwmMhOWbwke5EsGIFPX47f8WstMsuaHMxVs+fQhS4t3Akf2muAqV0aD8H3e87
RxSxMsTJDCvjDk0wUc0LzRf2oOIF2EfFauH/RW2SuzMFQOwQ+wYwPJHJeT+Uj0LP
uZtB2smrvlo0Gc1huf+hM5H0RKo8IyPwmlBoGTsexKa/F3qAF/uZvNT4/SBIn83S
Xhfdqv+xT5KjY8oNeiR0ljhRnLQQfXX81rc22ax+PGm6AkBwxNWHuPmKHvlvCqQL
ESK9hePnB/Dvmu1OSGH0fZdw6SZyJCJHyvLJbpvdHQgQeU/WHV2Zxqf54DGPAbOq
DPG2sb+shFMvMjIWvm3lK0PU3qSGYtwvKfwqLwP4g6N9FE9wSibP72wPu17s45t8
G8js9zBQva3bMtEfU4iAQLKcvhr59GLagB2L315CRF9KmhpnG2WC4CTabb/pH3cw
I2rs8CW6E2NcqVQ9qbNChJemP61YdiA/RUISTAkjvWb8upsQafBQrCxOO8Bfs2Ek
gO8QVLSmdaP7loZ1BuXC2er+ffZzc2XWq2Cu+JjDh432v/79BkEw1EZx3MbmPMti
9Ew4CWM7gVzY/Vgjol+0OSpw10fXbj+jcQBIp1/CuhyUSShX73/SJ6xu3dj5ujlb
BoRC0uMvBXqFrfAnDG9uLypZYpwn1jj+pBwz8EXdXzrR+BSyXs4zqABgDcd7+ayt
8Bxfs2w8tdkaAL4F8qx9FtD9y7aMR4wUK2LdeSWdzfN5lkW/5C7PzJZVBKVlKxHI
LlzFVnXL923EKHCWLynMVEekALnvIbBocKBMaJFdr8ESN4rm9+3Z0XobXADdM1gO
3RP0I4KNCZF2F3+tCO+aYqcTu01IewIV+YYLHWo7FvMa/rujg5T8LXGl+VU8+I5u
7OaoAoStRcAAL+iFfUZg1Fgg10yHfLDjRSyVnvExYH1QR/4PJU14aQ6EsQ+J9mhb
IxuuYuwCTQpegyNz5A0xG6+zjUyg8mmElcmroWovsC8Xb8yE8PKZhly7cgOy2tiy
iWaOaZVZy3RCa+99hvQBpieHihehEs7xn/Zcebs6mQfJJrDuzUCwEQqXQp3mZdhD
8IulFDTZGZe+/q3UFQ4dRNGDI3cB4JlweqO0rF52gLmuSoDv7dkMXYVT//anDWGd
RqHCIHhF69b2spE0aHH67Xbs+pPiAEZGQ9uQUE1aUfNE1XRePa0wDEJdo/fJ9xvC
UZcbzSBVH13evvFJ2Khx+6CM9d2pkSnr6rGXD8TLUKnn4Vx6n0ganvduCUUdkRRL
zI5jZJxx1iGckdECfBmfgQVMUFhYgZ7i+LKj0fKJiDrxB4YowvalPguhucd/pPT8
P/eA2zQ6uzSOKMYeh93QshfnNuYRDneQ7k7OVkgBUx3fIGlPAohGRsVBylfideuV
mzj0nbxGQlWxQxYoNJFYHlqElHCFlBictK4evXd4qYpdSQq117q1SwOc0atcWh9w
pxLE9XwFk6XaI95ROKMTd01MmDY4xpWS3ULIlvvh6/C1+SuMp9vbwI7YN4pdL2dw
kAwI+3wamCXrS35TD8iJ8GR6sFMyyx088SGTtovFwVapRgv/Jz+eZrfXoAMkcFjQ
CJoAADNrNrHx+wbSu8qmfJSLZ8nLX0sn90vLoCvYP7bY5YohE5nTjUWPFHJjBLwS
k1zWn9QPF/vxNf05OrMWjvEPEakSRKC40N/Gcwmb4gk3kfBgs7uWEv+BZmskia4p
lrcI4vlBdniGciy9Nf+fzxawwh0cXVyxgOzDunRvccHrVCFyNWAYXWJVUH14sezJ
ufg+tu01V8le6ZJV9/i4gexUqR4fyiZMzfiCIfXpWuU67K+e0mGSslx7ClVnjECg
BrvsFzquGYYTdu/D1q9fjFn97lQ+84mIrY3OiK+nNn+J2SRrX4X9Ta2Mvlw+34OK
MbB2SGNNCtRslrCWhExtGeBQcwWlBcY1Zwb0YU1vtA3bj4dDNVu6qdjIuOhO0Knv
RA2W/RLUG9A0q4hJzDbhG28nX8HlUVs0kwhJ7HeuFNnyPDCBbsHiyiB5v54+lM4T
zq7bW2yGsu2X+YtyWVKuqcExlNbBhmSB/Vugxc0nAEaFFHZkIBCSSqcw4ofVpQ7W
JI/AimHaiMR7EGg+/Pcy+oB+4jlmfRVRIjKhI6QQ5pZGX5Wo+Yn0fHezaVOl76gi
G+OfBW3dZEcAPAn1nLTd6QINHPUPwrDmkXsl0vc58bj4zniXGekC5CoTp+WQFEcL
wyzUhPRrqn14VRQdP7atBAigMD5stWOyCdZysH5+a3sWm5BtgMZ91Oqpz8MjvgYZ
wTSxGNaHIH+yJu5x0O/rt9PA8cx/e76tC8BWJQdTiBBje1U1ltXpjJ6QE8nbXoy1
te8C8SjE2sxGY+zc6XbKDg9hJ+vk0CVrMmOVHfhSRWRUBoR14u83sCtxgEa3rH8+
/CLRgIpEGfykyJVG9dSI7LXH6OvHVRCufW7R50FZzS3lkf7ncQPgqMTcwSOGUOBe
hjeFhbvVcysfv5d7a+Uf2jNqTzPNcVYl4l7kJUMDt9yeZI3dTrZjscz8oDH0GXzT
kSkkrpYrxIC1jhAY9xncn1pkuFkg+s888/azNJEJVp+iNnrJ4TrGwTFQZFzSO0V0
qh/JSzp4BTqrwFkT9H49LSWa+Ha7zpSxIKhxSS6uDkkZrgrj2zGjAz9x5FJ2ss88
4KlkA/tEAaC9Pu/htBhcHCdnhXY2WH8TGuMGf4l68A28Mj8fH73BYGmf5THdlF6P
b7daRhv77jgwkhk/wilKDxZkEstjgKntaIQ9l9Jgy2lCx+c4MGQeSTr8pzdMXI4i
1rOxbBOGjxW1s2f5CxUXOA6UV1g3BkaFcRyb2KncEkTMkiSuKACAfLhyX+uC9JyG
FNvhmwz4GebN7ijevzuqr+a0kAk40ICsrLt4RZmIPhrA3Ph/5Sk+kUz+6VLO+0Qz
ySzTeug94+mm6AgtC5G6af/m7GXtBp24FnQuU6anQY8SzwB1b3fxXmt0Y2BVdsi/
H4ncT8SVDTi7OYtdVGqPP6ZsJjMu9l6Eeif3oCW5iXWWsH+qwvS/T9PnV3OEkpRd
eLKIPg0sMrjBRjfAg4t2LWDGf0VjajMwl5aZQWLbzgw5DRslXESbiNmWaKviLgrw
g5jszp1ap02/SfYFber3EA9/wsZtQ6rRKOaJ4SoyM5013BjGQnHBcRfvrqiOTd92
VHoQZr9gmNBRQX6ktydShga5wXvoN/6wGn29mB6nA9pP6XEQ9qFOh1fObSJywZtV
hZzNjUMWYhloJqdJutStk+SljDsHdP80+3rwr+IYe6ryCLSqw4sJD4Jv39UdXc6f
GHsM/2bqGS/c30PBVjfmoCnaQlWK4KHBCAPS4A71Cm2N2iyrGHJWijuRn5kOONtd
ji6LT63AzVKzEYifeq0UgnZlr6ikEJHNw1JueadpDApINVXGalZO02e37dBHhKAT
eW1wk0XGlwPAJU37GXy9Y0HBV8c4jkuuhTo6CsPXjJmuyp3uHBLoyoArfmcLKPOi
y9fTKWWNKRognlGK2zh1qY9bSBmesJIRI+LxPKyXbUrc7cvH19Auh9gbsBh1SAIZ
moddSWrpsR6LL1UyfsIBXi+GwN4BcizXx7fI5ZLPv4nsKV5knFrbmlGBPWpqQAFH
4h5LUYqLWdAF8g4Zj+d+ZrZN0cv1xsCXGn7uafHLoPWFMdS3cn6ahx55Zm7rCr/y
xCCSSD8FCuwyeaiz3A/MR+9suhWn8EyzYfDCdIHFUgOcVM+iBBmEDNlglsT8FsAC
3aNeKj/GZgqUGPBwbrQXDBVriaHbO72kxOi2SoVjDSeT4iWcbh6SAhAZ/47jH6Xi
26TZvDXGeB//1MJT1SZxMC6NGXMd8QH5mTmMVjOO1IkeaRmocEhJTFOIXRJz81ei
VJbwuJZbgN45MnPY3zDDgys/NjxXyrI6RZpcY+8pcATddEswxgo4XJIVPRupzMkZ
AipVLeVcT0X07lJvNO9jyjRfcmDN63CsHxNkP1f3ZvN1APVY2twxQos8nmnuzA6E
WLIgSUnDiXQq/3jpTOmSL+pGtJSZ5wPqjsImyMVul9xt+svRSNA4wZkWEKGf6PGs
0Ge7+Pbzwra52Nr8737NujNueunZwlQSSca4/XbLxehPjNhyy8acisQd6aFocnhE
6xuA4V+vFPT/e4Rw8WUOy7DOBTO57GCUix13SDLTY7w+HXSLQ7QqqzYs1gB2bcDC
XHIKCp3VTv/D72JB9gOOhVgA5y7vNcCNEKBoO+cj7oT65cwF8odoizFco5EROVn7
rc3BcUI6OHXeAUWmmFxi9KzfAljsee4VSYGwAXVPvM9GFDFbYHVhcuq4wsI96vXP
MrC1sVx8nFcm4zXGSpb8DsRg7djYFApq6kyl4dL1Xn0QsCo+g6R1yChopnosK9Os
Ld3cVFQtZ1OZ3KJKL67YQ0fiW8hn7qE6y6PMO2gPGJglknL43aM1WB+HCCy62JKT
V2C5QQfsKzwauRVaD/e3hlPeo5arDc9YgY90pBadWSX6vAMYLvpz7l2Ze/JtmBs/
ybx0ohdQ1WcJkaYEtcItZbWooMJ3cwLz2GYRl7G6El8P3HtRfQUWGqngzWzPF/Xu
6s1tUMs2TmSN3QFNwl2+e3cI4lwHgU4lBI25bSAUdS+UngatrPm48hCszu+SGaSB
Lq757lSE3mOTZNlTlN6jfzLU0PowTXF997QYwlZjWIfHyyOjh0geZWllZtOIUS0I
le4exa8ygqzqeYYuKMKfEUZ3w73NPuhbx9iN+WI/gIJA5W02DLM8ougX71Ns/WiN
H32MZkTkmTCu5CucIBYkRQgYHb+DZC23BCbzC+xmpvNLmg0lF130iQTP9mAQPiPH
KWgMP5CtjCObTvwOlZFbsEoy+878qPmOBrrHN0eCKMkAZO3uE5kvl63C+siwwDiq
TpHHgN0t3tplda0cCiLXk/bWhR44kZfmhR6ljSfu5BEqNTXCcsDSdt0rv0XXr1/c
lJ8FDFNZn6n/H8HqMA/CMFiWth4x1v0afeKcH/EsZQPWerP18+OY5Nf/tV1v86Vj
LCVR/mJg2qGW/hMAzqWFRHtnm2esCtEOareR3vKeCz/95mEqUaNi/TXZx9AKJfSz
AExcI3GFm1Q+9EVmTBdTxMZjNz4u6khMmNni6l63U76vTJKv7FCN0/wL96FT2djB
r72OE4cOrBUQleCdaO38RACY5QzVgR2ExKe8STsiih7sYriRKrS5sJVdaQCKw7KL
Cv3VO4uBx69p62dmvdg8jUlnQeQl+YEsGM0Z0fxnpfGquwfLbt9YXKn+eHlYg+f1
QkLMLKeJukJ51aAeW3ELWWdHMw/j7dl7ry+5Au4nCMv9L1TQRuo3iyokrZdLY7HG
xTk/2H3YcnB1cl4sSYgj7JW0mopAJlQ2XGKHUi5op/uNmCGPooXowvW1I495NrEN
tSZXgJgmC2DXvphhFz6v318ZIG32Bs3XllSA/Ie3tt15KW1DJXpHNDuul0ycRPag
c2TQLBtK+roR8W/nCANyj05OqFzrpkaDhYn5Z7BIOnVy4ltOSBFknRHLowMkNj9c
d6M8J5rSRmcCnQM8KZvdCFq2rwD9ShWAGmmRwgWc52wy8EAtkPjOXsXyrGybl1Co
342GcKxOVTHB0DIZ4oLgzSqFajflxkJbhp/cUeeWitPexUxu0j8ALxijj8mEy7VI
+z1hg7NdaYLjxmq+n5iA3JWJ3ZYJWxpeATgUBHdyBK1rABGnJXBeY3XZ8qj6OtVP
quqs59tFL4izJ7JU1B0MFD4I8s6Vp3euWkjukGpnfyyO6RSpcUR+a1k9c2HSipJC
Io7bzvegiiLl4wvmkFTk/1W3oeLSWi/0wEKuZifc8W2JEmHAarJXRnWy7QCfQ66I
0pYLPTjrNNtJND3kzEcFyYjTzYk2kYouc5lj6gcVRWUg3S6jvmnEPQRZq8VJ8H+d
PbnM0MNZ2+/4g+7R5aV4UttgSO1UiavGtNeWg+fnKPwYJHE8smj1T5vFkioe9MGr
1ph1LF9hTivhWIpNE6a5CBSkI19si0dlAXPoHibtkowKN57cxdI9tR4g4kHlMTmL
imuUpUwv5g9CP8AOvxxGnKGUqACcTU4jHqkZLAoDdEtccgYuvdTyRGeZA+cv3h8K
Jqm+F39IEpd6SprO1fSKXgTRKZ4jx5hJpW1iQ2OmOaHaNsK0ZcV0RKb5Ah3kFs34
kXHFu1mVpqux8tgE6aVECwVdr67RGL2uHlSvd+9TB09rhXm2yV5J+kkKV7tTqw5+
xTuzyTvNbIaJPiF96wulFPvYUhMD0rOdvfbBNBTBSXFrUjzeuVF1NXCti/Y7Yi7o
wQBq/6OhZaAXhDpJax0Qgpvb544NXaISwEM/fg0zawxTyn0axVIReU4X3UKWymbs
Twpu7In8jTT6iw/hn596EEwPjL+qVdAdmwLEElyl66N7SufcZE1v+Xs73WahZ7E1
JlJzOO96THmg3mBA6fwlGVDWSvSR5xbjGvoKkO7O0hLrPgSoEcubR2Gm7TOrnwsO
RxzGWXz/oK6/nTekdI76qu2+eSjTAFPVygDrJXtwCGUbUqHJS1RQCPPKCuQxow73
wSsxhsnHULA3DJUNhTq4iGzl+N+/Sk8gMIG4k3/YaJxgNa8s12jRo4VQNNpiR0AJ
M/mFrrTW+KnzHVE1yvCQj3E8Vfb1t/pb+KLZlRziXt0rFTb3JEUSLUE5PDre9LR6
o/8e6D5d4a/LfNJYCT80IZhi0jWqA2Jfj7bbNgVe2lsiV32IUhDT7Pi+DkqhKBfR
bGV5d8GqmCtfz+28ZKHuNdE9rV24nAXgp3etIwn6X2Sh6s2PfZPFRue/efXQhqEB
LlS4P7bt8OKmNbVQhpV05OB1S2Az1zK593zboI0qkr+f95g0x2444A6wiAom6e5k
xC4NmgUlp6wlOpPVu1BzWpLmkZVGMWdxDpDm84AgFgNFEaN74ihC6iE7wyq3sunC
v3ib2nivv6FydcZwZHYZv72ItFYb1u83EK3wgbvwaUOgWByyqSZzh7arZ2Qno9AO
sTKysR7qLTZrCi7CCqgk8v8j2o1Ag9oT2ETp0F9Cf7e2Cs7EaFAH9tR13ab/1Hdj
bfiQscnelgnqjlRWgTU+k7qQ3nf9CT8LA8G113+xpgFHbF4IDCBlk02HracaNrfK
NnDa4u0H17jQHLFHI+SEfWdP4j5ehQzobEACoL+cl3Jc4uEfRssCMqBx0OmLx4aO
7g85WDc6yhjVXfp8JroURU1V734ZSZuBe0yPkOcVCCCwfBMGvMhw3iyJ/JXIK7PK
8n6HbveEo3OmoTvW6D3qWciNco4N7lffYHkygGC40zS+ObkJsACdX7mqURYwD7+J
WQLkjtGzgbxDqieTyUXPCNI4nDJaxN3mKLa41PqPlJvJWyfzqeVflK8+569qf9vn
VHsxWiz3iYRynC5/++EpEi3aVY4h7gSJdts7p3UtyfO53NKj0thznnaLeW1FXKGF
/ZUlAH06CvHhNXPGoxhs1PdDSNV/7SSU3H0DULhdRjstLKKPQJPotmC9OVkwOSKr
fch0WR/prhOgnAJxjQL23dgyvFCxWf6uKmvL3iJgnVV7bTdidvoW8pb74TRDhNTt
FWt4fvFFTNXI1gct1owuarLj/ug59MtCLPpWslJtJsvq44bu9a7khmj6sJWOOYdx
oHwXbMBfRq+RDxCbm3FOX4uuT071KnCpkGA83RiJjfYHMwRUTt+XYPiwhDMH7eGy
palSvlby98HRZMGxzx9IwnZaJE04NvWtZVseKfnJfYUoYwx7+/vgkcHrrHZbVhfn
woMoOgB7up+Goi0oFNfcsNV7ynf6TiViUhzhzuxezTiqDHGO8pEjusgcIGvILbjB
zwL14rjWY3T8aB8jWxUQAfe2QXRxlpvSMPiI+L1a1XPZFL/rM0bkZ9YL9aJt8Mjy
w9Ke2QH+cWbF5jFxDC9ksAXjkZeFI7I/qA6eQc2KvoVX5GaPA+VjDo4b/KhtG4+0
b7Dhda9FRy9BgxKkPfb5mfy6ejRGMEF9vEn2hh6I4mFuBQ37SRJw0h/GnPPZ23Gl
bLvBNqPjED3pqW+0P423wQgZ0vrZjqdlhOf9xJPu6ckTRk7ntnsk6RQPRXyFl372
7NAnWdEe//2260U7q+vj3lTtbyZL+eSrL3dUidYQ7u3jSi3fX7i6la2cgaGrJQjj
+vn2S5rAFNu1GHT60IvJqG88e2fhvHAeX3NyMbcjAsn8Gl/+LYYfaCt7WPAB4UuU
alZ23m/Khn8P99oj6P/XRKJavQpx7dWtAkxnsHe5QYwnHO59ehVaoS4u+i+lEa/G
y6peq4oGMdofOslUG/4w1TSlahjX9zWMJ6PbgmM2lT5V7qT7+QWcEkOHwAqQ8Dp1
4sA2TPbYf1RYptHLCYq4YdX4uDgpS4x8y15cBu5UCcZ+05FH+LJ6V42GHvqcdSWF
iea+k0eg4uUYy883SxhDrcSSqdTlcP5rbCkNCGtOmsi9IkTtnwE3gul/7/PvQ81n
iqD7hROM2Hs/v2YxEelu7Z+GW/5U56xaQsMktRvAj+FGl8weDNjl4yF1QkhE/bqD
1a9sdu7Iyh2gRPrFPtY2sW87mRuKj9IqAEvMx5t91D+ZFarHvyDRHof9ZgPOA9/a
h+JjzfiLSQOOfMbQaS8dbYqnLLuF0PMQ6E1hoXDWsEhOF4hApR7SwZb5E4lPsGTy
1POVCt/rr77G1tWU46DaWh5k17AhuIZfyec3DuWYepUfAyOjq5wF0W+UXLuyrkY3
E4x7yw0FenzssMQgWKMP0D77YcVC4dgyztzbmLuNMRfoyeLZ9Rqqyg3f62Cdb3tj
x3p4Lqv09/6SBoyJ90fR/XMJvhgeG7BXQvfRszdGevl+YnDcRHKgMdsqtsBuY7Ju
4gnV1LdB5cKK6Aytm33lauK9KrLlkDgv5KZ/ue7XUWWnJV3ofL8Qz/aFdVZta1WV
6WQ7mVIfilhkYxxM7DC3xfK+DyPgOra+kzDrXk44dcM90NM006Q2LFg+eygqcqLJ
mWlVwznh+nlu2fbOMjLW8jUeiLuGpwevc5ROccquI0+/i5hAJDMpHyzd6Wy7xAXC
r6vliXFhBJli5WPxR7RYlsmYW7VET/KBxlJuoYZdYZ+jCBvMB+RJs8BDdR+mi4nt
OHGtBNwSGQLV2RcGs72HqDtzlY0xz9VyaJ1n48za9yUre2hspufm7myp0gtg9oU4
rLOgqxjsAJKPKGuwyOnkw8UOpzs5LWadweLiyEqfuRxqumuIdhkrBgx5f1807XpH
0WtU0EsxEP/cBaFbAN7ejIPQORt58cNq6eAy0xl8Rsf0sEar9TbrMX3Fb2n6RmNV
ccd8Ap5/E+uY1TiPkdGa5VGFkrENExJY1cKJxA3JsVRRpfRPTVvfPZWQUG3lEz+L
YEcIVrNI2mEYjDDFVwXdrdEbQxBwY/klfoYMYQNFHqdgSYpapLgjPBvj/KSIRvUD
6K2b7TuLdDAYVN5iTWm3/Wp04UCIdo28tA/6NbJ+ZaAX5J7o2/ZHq4plWtvdWCwk
duohAY0dkBuTi7dXoxgPEfe4HqGltcpFMUR17feHRjZENl9QHKZDMoV9BNjsU64I
I6iYy/n8UWgialJTOEZ/fps9Pp2iku3aZWJ/D00+Sk4H3aEoNDdiCdEwI+BjVXzU
XYbU84Ije7KT3u3lZwjUgFsr9Z00cKoKEP4Utm20LwS2w9y0aF4Z95plH7bAIGcH
md9LWel+bPuve4ThQWczoo4mmHPLZ3iBqhYR1eUWgztpIzpvDL2P1KPHSoxCOa8o
PSzBVvrg1GFN2JkioaUT+FFSBcnnh/tvQNskeeTluEDw5HEgmkpT31JJjbSbvHZV
ZiMh101Hpc83sbr2cxPHsO4PIhgRVv218fQu9zRMXHP6Sfrwk1FwM9SOk3Z0Qv15
vkIi+jiplgFQF7YdkVq0R1Ylj3VEpHv0Rnx5H017Tx2uDUm5b2LjZbojNeiwMfvD
+Nze3Owd0kyFXqa+YRsrOCryCe93bimNAZfAAsIxYV7IPWn7lE3kyhtLyL8XdgCJ
uv1yTsXXUGVzHuI9JmDOpgx4Nxv/ReHIFagiQkVYx7oIOke8xAzcfmunX9AS46zA
h+Tp/FzV2/OcCwP4g8KwZcX1JsH/jzAeLMK2xyAzUx3CEy0/pqrTYHzgMM7DqELm
aquIEa0UDYN9IKZmRLABPL9n17XElKeg8zKHlDXlMukZUweJlBUrzfsejmW/rfAa
hE5LEXCjCVIisWKXHTL5ww24/J7WDzBQav6k3uFyWBkFgI3KvGqE9h5lHwZBhKf1
HzP1iiu3qra54UeKm+tRXVY/xdsfM11qOknFtthhyhnQ905oH4Z0gTz2r7rer5vo
OCTcVVlbxDi1POpQCAhXmGASPPtFX40YZ1j/YMmadZxUrIQmjNEQEcDZqnZA8YDE
2cbnUOHKu46WPfu1mAn/Zw+4jpj+2WOqRusatpgIiTH2KY8a+fDBPLyf1qIYBYW9
1syGQ1w4XmOZskWwmW25SEQxGSlEYYN6IoRuHD53STB3ZrPIZxfGNYz+XmkA4/Rj
12QLmBT/uHgPTmUpFCtgyaa7aMGuWrPlyEcTXbDPKR1U4tWkzW+aTDrgQ7HZMGFv
wyIAP1TFo70vDcudZ9zIvEkDq9zU8SQH3gPeGABckG6kJYnjLNKmBYns+UzfGk49
9h/FTdem/AgVCq2OuPEdGeXJ9eAk+kU8P7avs6KUKYECiShgZt8TYZ2knZeK13vN
c+I7s3hqxAwG1+eSCvpF51V43IwgEhM7ks2LiRLR4u+Nn3M0/WZ6aSK1DC536inh
YX1lC6ZmtwwT2WpZY+2oWdx3PqW4DKjGmp5btHC6sR+MoN8ARfTBpyGpuiNVC30B
RY/C9G8Ys7myXyVqshB+IcypnGh8JZCN2gJD+rSlk2KSrfBwsIIlO6s5H9jOkNEs
6+PnX2Hx7E2sF9A/oNmcBQR6GTFZXnDPjHnXBjd4y9LOlmi6B4VAt3BBkUpf0lC5
nkQkAxratyLSj0lDw4xspm5pdQ/+l4J/WgvAmSn966ba02ArE7TJv+Mp58Vv3/r6
c5F2EsWXtkk6ItzHzPAWqyIJcdJHdGf6TBdkP1BnAK8RLkzuk353txPEp0rp9nQ2
vFuT2aL8K8OQIGyFZfHg1tPxTlB0MqdbZZYENVq0CXTuV4kXd+jGm8qeXybjMOpO
h96Hz1YRugpfH21HMjxluNBnNL8E6DwqulbiJ5QqaOcFksa8GO+aGILBvb1UNDhr
6XVBQM4Dq3H//kgPas+saROYqUMWLNtVrvJXjob/uDj6Z+2+Uf7+mLdaLBjErUw3
B5UjpV/Gj4hX6lelwzL4tAo4EGnzqNTR6N5e4nbjawsQkktXlT/DFoyNXin/12js
pTG9dS3VRkHBKWWaGCIb6JGYhTEO6GUKK5nXylWolH0yJObXozPAr0pc8UH6CzgF
wKU0aGaPGgDeh3oqpUVYGrDhTAjTHOgsgxrIRIfeDgSOoACR1KR/bhbs/LAjbr2y
JQv1wC7/LDUmFos15oDqqm6ie9nLCjjD6pC+qbQ7BV2opj6MBKHQ/SgbRtKKGmQf
Rj822o08Uwlfj1Nszv993khqglNWDtMpwsDdO79SIFr337x1VJ2bu37LUVW4eFqZ
QKX/QZ/D/LlCAV0Mdrg2kalac1uqmFtbo0/mq93z/FNPXp/FTyXl2T6KXT1i2pvE
4gWKYt+ob9GBlYkyeoUv47s0759647Lbpo2T9+R78Q/6mbEP+D2fWMMZkrWHpoxO
qixy6cMToezHNCvGcIWexMtLUtB+N/geWhVpk7guJLsgE2pfg23Odthzl3C0t3XY
2x0j1FKnVpIR1da4p1LVhXvvMjXIhUnvjyiHe+wJoAK5ezG9Ctik9udkl1AL4PSf
79sfCXYF4H5SvJO2BRRKW5rcEXXc+BL92UjQ1fJiDLEemLZpG3T9q7b4AWcdDLnA
RxdhchpUoAktHaFnLL7trksbqu29QJ3R/Phh+Sy613xZA1uapPqG7ehu2/qE4Oo/
fDg7VRw5sDfvAR93BtcEhBE59iBXRRHyTxoCiVzsC3URQ4H7uy3UDzS1UDPSX8s2
3lcZy8gT55dlRZQs6KEuLyXfb0BAb6scOj1RE9JToEcSsuYNG6dS6FN6NhHf4+0h
NsyejJ52LcTc8yAjs5CnkZVweGKnERe7K0Hkx8a18edKgAstZozP1JsI1j7EOZ8j
yz8ijvJ0G1qSQw5WIznsMzlysGmPSnLjbrESTuVoAILqsFGozvZ2+sBYFWaK79VF
wu1MAnoKymiS3jIVXJ0Wy3c/ES60OJaWkrGxqs2AKgA/gsimFSWVFbAeu1RaKpQs
ZWntVIrm0zbJJ1exRTjNr588RVaB1SxKTArcjPfSGEgytH+xBkNJKatD4hGanmLw
TPBFciPATry/uGuEHfTkzfWuXBNGcrUSTwPQ6XUTGnhhlKErS8ySF4pBWV8oZy63
uMNlz0+YY7N4Pc32e8MHJPwXG9LeyFj4ChOJ/xvcx3R+nXyTNdEp8IBTh08FnJzP
l5y0vlSUq3PbzxX+vAZsdn9gys3gd4q+3sUD+FK0Ff1LJIvfo3KuNq/MSccXYTfK
8v7rfh7X1VjZN/k9rJZtuYS9llmOCn/HQqhtRagJmsdLb4xlGDwXB8jbqdxa+rrP
UUDkukkG8+wG1lXkQXZZekx7OKF46c46gwWANKPVbg8gPEBf98jpqvowZWuCduZ4
50s69zV34vWu/UhkasWVp394hBjwEfnhwKggh2yp575bi3QZQ/S+RNcelm839SPT
7rSYKpqyTXZUv1edP4ulFCwxwYK5H/ZA8SoOhPc5tKk/bFsFxZQt1dl4OS1A/DBj
7x+JF8IgJVMd3ESZNq8GBUQF+FZI0Uxly8k1HjYMKTXmw3NUW4ZH5d3UXYMVFLwx
UAdtFIxfbZvqXxx2bnT62G5LVo8fTGWr3yTuBis1CiNqblYcH2X+IgBda8zvkFSg
teX7v9lifGyRS8SyTXCzsc5GYbVzLvizc4D72U8mmZVXBDJqu4PCv3/NAfRnacjI
tm9iLB0hm3ACRGsTEpAyTUyPyqt0KZ35hPcCffLLzavJOqb7MF6SFDHDhtG3mNgj
vtRLith4BiEnXy5kDTjnP0654/KQftqv/UyRSnU0AMEtBJ+wY8+R/465IQUcgpZr
LVtrcVgQPVf/ItpQ9vH1TyHgx1NaIv2tdz+khvs15SmWVzJDSM/sWPkeRPuPqeZA
w2HRb64MR/Bv+y0bFoQp8Shnu5xHaYj7rcr6pP4vMsrfUB7Qt2p8mC4pykoueo0N
+t8w7NZSBdqTl/44o46R63X54rKfYLRxtR+VGgnjlWASeGRM0uxVUmvYca6+YEad
cBnndoltmNVJ20re1zS3a+HIEcHk/d6B/+Hax5Dy9R3QXiP7w/0vO4rxlDcQhbkp
PSQiYWMmbm9wlwb2Z+uFn4A109BGte2j1zHu2tjOTHXUb8Wlfaw2I6FfYfM5K/pn
LQ2OyRY5YO/2oQVqXqOhRC5e9nPPNeATcQV3PdfPhoN1+50brqWZobnRwgqqegSA
mkD9X6cEn9p4+JEThQGzgGvzzMdGDnXMlO3LJ2jwiekaLKstN5uZCt//TKATV+A2
HzoBBpP4xfSF0W5UB9+TqRbl2MPs9mtlAdk1FFQ1NNQVp/7hnI+c2zNNZKdY54H+
WriZn/i99ZlvMfm6KLTh8ll6twMDNVhJ5vKowp0qTmo87LU9ip1I45Gev8iNSGrC
dP11pf4vl02BBtzWMdChkEq+IiRaARbUSOU7hOI7LH0VvTqTd4sZY1/JOUESPp0Q
YrR3fzlcnoTME2LpTvpJxZ3+JRH4jMka3L6bhCN362p7eA+Tn5DQeseMcvXMZqRV
MSdKFciCVCYmeIJURD11fSKraDvjPGkatDU1D+1ztW0o4slB+Sbp1pgDSAH12Nol
aSV/uipkTUDaE9TBLNJJjk5l/82JTZ6YPlyMv2S9kTUttRoMvdeScsAJZaYiUXZN
LC1HTonmyITd1IB+vmYFNX0+SQHQCEE/UzBGuzsVd1BHb4d5dd2QoILB9YVSY4i1
b9NF+FTHipmbF44V0mn+zJ5EOPanol2XeXgdBXNfirtg6HzMfGDJNBmvxs8yRuN2
fuKD+haR/exN9+NOqien+3WXqtqMmZQ9jMPy+7lh08QLG43mtfjF992wTFVDElAJ
7/X/uY+buXYU+o9ctt1f/Xb8xE5MR/zBuXlZDFSBTmwIoodUtFpjEDCmykg5Pqqq
62xccS/DqDAxHOFyAdTdW8Z/BOx1yIqbgXef6Ex9kWjwIrzVlsN0IeO0UqRHQkLC
WPXbEC7n/+v7fHIpuZS+tCuR134PHoLjECD/ydjcdEJm6u5U5N72bHXL5ImLgs6k
ErIpKg9zGOxlRh2vOWgaYTOpoFupKjL2ROkldbCI/l8nzlA1x4Y0+Tyrf52E7yYV
2DwBSWn6NrFk8C/cXbTmB3tvVYqTrC2HHTd5LSf303p/5cEXWWy9HgVvrKwmbroH
AWgefwL0ebtjJLq638cokoAbUkPyB5c9IzbQpE0OtHD/z/gJgCNm71bsEBEu1QCb
K03djwgvoj0uJ75xqwQu2KHarkXBCOXfJ23EwPenGqRRJCMhciGSPXB5uQg9Y6P0
n0J1TgTXa9eurqFnihHrWXSatVWXXGgAi5jDLfDQVDwrKI6AZ1nrR/W30YxmaIZ3
W9BhHhxldjZyTFp6GVvgzeqhnLIrn/65xw92lFw2XvixxDoOJXOIp4LwHHzhfPdh
KEQzpOmKLFYWIUczzdMozUVRja1YIn3ffc7rrGTsI8d3rYWGeWnciAxfTgNPGNxb
DC8ba1OH185/FireZTmPTZ/l6kjKibXYSuR5Qj/eU2ZV+zhgPGj6wEKQfWS/qyut
blm2fHrnO0CKakwWOlksdjVepv1jlO3txEpGPfnTDVVLEYCDo3J/hyhg6tBiUgAY
U6i0pyXT6e9K01mquxjGvQLlFagIrfWjwdXxq3Rw+HDu3OcE1BNB+j8LtYcLXOgE
tO1yQmcrXhiCvOHqwx1rQMWEUhcWhmo4dqoXuzCUWFJCd1b082niOgYg2/oelH0H
i/QP6WQC9bTPVZNdLzM0f2PaRGjTBhBfpa4bcreybFvbaJ31qFeQszxlKF4BacyM
fDxsgqnok9DRmDJNbz8wbSL5C3yRanzdD78K/cq+Ul851HKN7yHa5OuM6gxT8rea
ARYYL8o7wonP5qVXJ46ic0RgYWf8QDl8gXpmTceG/ybIz8LGQPy/be7uSDRjGJL0
8fWydMcIWwx9GsFRY/5kx3p6G7kyofDXsIgE4FuR6lPGUp0zqpfxXDSm7D+9WQ0u
av4XWBjYteL6Phnc5oRDgZacAMQdXE5dmin8cgHo47cKx7BOb9EAUi+FTXdS0b4X
aEeSHyOAifmNG+2mlyZ7YG3rIx07UCWwxzm7q0dWWD6yeiZ3cGNxfYvgWrNY4bES
Gza1pcKlfRFL9OH//ByCLtIkLUzmnwMKpz7NwI3jYxududZsC2JwKauFeKDARCjM
NLrD5xZhTHhsSI4EfVY65u8BvrI7OClRa9oVKtM7eWGYk6ah9+pUV0Kjs58J2Izv
Hh7f7vOPKUM5GXXKqJG1D6rQ2x8NwaLg2ANZRJxfPKLBVmvmC8iDk2nIyRbt92HB
tGfdKCM16waaddoCd3a19Un1GRYmU8m4778644a5Cb6Ou85rxiNT83tLYAuBCYnO
8Iu4Gsr+zXuV1qUIuy7w8Bs3hyKfWvIIHnnalt8MOMo0m/O5NJ1duYUtrneAJ4ij
ITnfTbzHH54EyTpaG1lOHqpeKj2YouIazco3sQmqnSgXljBLzMuaXRAKj9SI+q5n
b4dVTKjhx08mNVMaJNc1tcuwRHtflrF1FGiL2OLQ18/F6ZN10zX5S6ouBhUFBWIA
V8knXnZ5S5OE6tAUAN46X8qXlnK6ySLTIYHkUYXFnHbVZDm8qdyg3fSSuiwMHtFA
IZ7kK8igHIIpJUAx9Ea7A+P+kxmgYBoi07O3IQbZCp197u5WcoDg/9O/v4J2Uj+C
5AkH2bE5fvLnnjZab9nxdXO4vWB4EWiYwVyFBGB6keVTvAw5tI/jI9AxM0mlk4VW
mg3Mwh1fljIioiu+MsSyBKFUbCIIpngKYh7dL/nbnLEvOVyZaIfq4RpumYjhGbtM
6LM+zD7m6Mt+eKzJav52Ua+jsoOgcTreTqzkUZGRO7Ecvs7nG+ooWl4jvmU0VlnY
1wXPn9UGnYvC7y6LteeQD99GJwSQQOZt4GSD2ZyC1RgfBoEuIg3k0UMLwUFN6Fgx
vXTe72aJm9P0AnmngZSdKI5bvB1hjJPJlPUCe2UpONA7zut0USht9pn8FBYrqFW8
eKNB1zwFgz3x6J1cYzQNPgMcq0HkPRDbpFezsPgxE9TGASV6Hj74Nnhr9sUDAa75
r5ey6vVP3Y2T6zh2lxTuSmJvjCyP8CWbDr+rKbeb3nSOeh5W1BpVKF5cND7zAtx4
aEEQPLuivxheWnaSrr02pQxZcjPt5XQE948MB9lna2JaCKUqrIGECMBgyAzsHpT1
hOdjoOEK39UxQgi1EcQxrGKhG+tb9bE+0QWExxo7CsXmoqiSARIwG/izA//IAZB7
UFWjKXtfkTBSt1v0dGHj+dD6eRY5ueItFzkYmByyAUi8VB215cxJVrV9Fg7jHpGp
5pC5cdHP9bFQGRwfPoBbclSUvjTe/t0xOGRp+NIdZ6zgZm2Ag3uFN9WyWNfqoy3k
5GMZxh6cK/J80eYK7xlsdiS6U9WSVrSI+QmiXYGV7pOGjcfgOcrSZsoIbbf8fZho
aTpcP655LSGLQeaGDk/vbAyqMcz4Vf9TVC+KXMjoO4Bsr1V9d/SHeQAhIb461Vhq
QK8TZstkkFScQWdO/UT1uG2S9TIE5dxvONzT0ogfCdWHpYWRxdR9bucSQ1MlD93H
Z/mOdAH4EMx/RPPQKoKmKbreLjePbdwCB+lyv2C8tNoK0HWrFVzKKEIN20iUJTSY
3m9HrK94C+8tFxqaag5lVd+FJUe0TwIGcdRpTBytVOAIAMxXtfwlOK76CtRDibrb
2CmZElFsh2rpDVgj5dMt3/6K9WMO8jVD7zmIqJQ2WLTmHZzcKglrx7Jp6zLmvstn
ndUyFPtrAeTFDMHPlS62GDut0efwYdc+XNGvRTxpcUt+zBTXSKHEtxLmxJ7k2HTM
R4TWAC8DJnWiC9YFnfgwy3jypGmKFsr5CsbboKx8EejmEmN+7ejIb9M2Qg6q3LGo
FXBtza9JjreOA83lxygJyBTkVoyBCRtXTFyZYSue0F7fcSQJGctYybHhMsCXbrN4
yWK8zeFHsGTZ/DhloFTkMUeyGFLM/VEgy6RcgBNpg59dS7y359dsg4TPBbt3HvFS
4hxOG9v/rShFGPeZsFb0FmIYCcsRfVLXwSmart8iCLdA1m5oZ6O9YJxg9mbWe2Oy
zi1Pv14JWEh6im+Vo/sLF6G0lCInhvFs9U9DgzEMyTh+y9jjfzH3nHPV3P741TSB
GbHqPGk0rwZRScETDasXJR71gkpEwNCRtdpeYoyTywDn2G2IWNMGJFawHOMG0BX6
gOHe+5AFMsIdt4mfh5K4tdvoqwju4V6+taFvxgyDUQF9xgmsoNrgijzTB8wTR1GD
GpdVHNnrXHvJFJ/Whhp6pnzJ85xiuumvF1DoTjkHZjoEtI0eMX+kw3lhBjxdVeJV
pB7AQzEPzfjmRScZDkn044aEJJLszvtIP/EkAgvDiSPoNUUgszu9eXBtnuXvriRl
D92y6zyIgv3cGyXpgGPfF/9EmQ285UUmRWcq52AOHMyeqKFv2luFNqlwR8QRBJBh
B3YJOjli+HDI3CU1eTWlP07vxa9N4Grn3IGApDVbz2NW5VoS68thIPsFVvPdI+Uh
y1n1Fg6kFx9hz4CT4ESi6CoSV2008+PC7xFN5uzWYgqehpeo7s1f3xL+LTjWn5Fk
4c+kdL0Bj3q38R6NVRApQzMvcMFBd37Ig+Adabh9jSpgB/1aFkOl2+7mJRtTA1/U
EgPVIdwPOosqio/+2BQpmChiYPxTsNf7RGiXLTPQhdSgGHi44QyAuFnPLxWFY65E
szeKjqV+kmOvRVcI0mfm4VYDzjqmxN6vFMNcgU9vfAsKlURvod83ThXns4BbNyLw
EgRBKBG8SoOYjfeJYYpGT6nodfgVTYX3QJRDxfuCYwKNtrvV9PAN4KwVZABMXA8i
HGQaXZkxHECnYaISqcfKX/yPvUBTZchSZe1F1TI64OLLZXpvSjpuu2RWLtkXEy/M
l3V/qxcT4kcJ6QRg+8eqpJ7eA0sh7HoxyqOOP8Xr20h6w2hepdAUmrh+mc6zm9wL
YeLh0VUroC9JjOz470Zr/9qeLqdZ/HVWTBflunepqBHWO8F+DKf5ZpBRS6PSpGSk
oFe+KVSeWbNUYVdBQ+3pOUBu/UpVtDOMbq5WSCjB64gDs11mLwBnMvtpQeYt4+k0
d5WegNCo507hQvP1rBvLKiq733xlv15vBVPY5AOlT+MFkejuGmF3Da80pTC43++m
Advnz95nQ1gN8OrcfQhNdKwqTbeshf4+R4Wbkqsu8BEernkLF6xRRyqxMv8uYZZ0
cnIRGcqARTODh65wSLTPIOjYb22Frg6ib7bru8ze2SSAtXLYKfWNADHSugsmt7sC
LuaDjCIIdOAHvlPa7Y4dsBcW5eagLEQSmdj1n0E6QXDYNTjuZmEW+vDT7vZQJHYJ
i8hdnEGIRdrg1Z4vRX7sfLSniGQy49GqA5KCXV5H7EGbjT9rtcqADkC37ecwfp52
GZ8Kh/y4x8UHADRrulFkQ4Vsx9CpXFZqdseB6zUdu6AoazT6wkT4lewKlyUwIZT7
nRTDokjXacZlD0ZzgQ0YRTC+er3HgFNUDEt9jIrj9Ht0Mb+HTohMD2NbnrGbQyQ6
k9t4GvK242FU7bNmj/sxTJXKKNgLD+ajxuch55Gvbp0o7lZs/HEUJWcz6Qyn4c6I
FDeRBN6LipUPFUhHf/zs1q8dydSN1Zd8pLI43g+Y24Od0qjGVppKyr7gJnYumSXF
+fuCzm3Vysgklk2Abgu/iDte8FAFi+0dua4vvMiTi3n0w/qDzl1AQjcz2dcPkaIM
DhqxqHUyuQKUawsm8vR072D3D3kxkvieTmwJGXsYoM/b+61DlQ22OwS08rzjIjVU
T42lm7eQbN5jtfI4kvlYjYvipjE7PQDa4t05sHdkq7H+17fqh5UVrrhH+D5B4VUj
1xTcl091kNyFW6d4ZC99Ydp7B7ZcnVwElQCFrbusPHkXZyeSWBlrTW1LwP7GeF1j
yiwfiJznmgIpeoa7vIucBgRsA9ULC+fPdWi1JEhWNA9Gt7s7LSPkoIvx4ZOcE5Ek
dQi5Xh+cLYu9Ei+WVUIhLNvhfaQl8z8CDLshi/QnX8EgRxEn5qRb9eMQL0RYGUFv
QpE84G8cJebymqJVqYexKYsbf3vi4vb1ggRqnmGIsy83dwyFf+/bLTfgqRIPLVbs
TkmGbn6X6aOTTy+lg2Qay8HHFFxUsUTfnpOCzrTzXAyuzjuTruNZbXnjUHQsUTLO
SN5wF1tdp2QTx8NNVzEvRBe4sA/w6IjYw9zggEbZSdp8P+IP9Wleg5HiCwR93onb
3Q3NVTLnmz3OXSKZViUpTzyj8vOUgwkVtyfH9k7cs2DQ/P19sfcWoSSQQHtilGcg
SEUNqriDtEGzKcdOD4+6CWzKZOdgi5Z9d9OPCsrFva0L0LVAGakYF4o0Xid3DNCD
5amLCYv5Sbn2s2rg9vaKPGdGJ472rQrVI2/Xa7NvC5PmEhmr1jAHRozsdhkTJCOx
gL9vM5OmcFUmvVXMU3nbIt3+nDdJemRS074t4rIA0UkOoi1XN/vhgnj10HSkQV3S
HOacmarCgp8OjBaD1mJ79pULrl2svQCNEEtfYuGe7NkJ4Qt9xP/mSDxlmJfnikXU
4Y77jPjGyU9droeYs5qeLQQsLgjVCJ7KuB0EKdZUxpHhWJ1mmnHS2aLXpj+89FRc
Ze3KmwaqtDuKODMDihlkJ4hbyCAtmjdfuBHjNCd2Zq0S8VzhvMxWjoBDpsICbjQ7
XYqh9+exWOxM+trQezLPURJa+YE1xWiPWHdlujw1xEA0Pw/NdkhQYWifvU9zjbPP
qKI3CTzv5F5odWlirDXnBoGozi4vP8+LPwjMpaNbwB7rdtVfwQP8fUYWJ8+XVPEN
NYZCJ+FXzUMHEgpk9aLgHCJRUg3lvc/dX2tMXjehokBkBQTtWvW9sbv90i2aYk93
b/voNuZlVlpgutTGAUrzm93f83ioOi1+r7Io+G3IVd0nWX/pQBnEyl2WEFxEPxmC
R7MXOa+PcqmNCT98s13tHVB72vwDDsymtShPSjfUNqrAn5yhCr6jET3AJDwC/KLy
/T0ORkDluK5k45ZCzzhF3/lUSMqHEcGgW9pUYPs13gGlIGUGHo452nVIeObYQUit
yihjnTV4EJ0foZ7HOCOh5+t8R8WeUXWz27lnz6k2wCsHSkAu6kqJXPgGbTMzc4kY
NJnAWiR1xxwGi+74sxC3CeOsrpjdYmMhQzg91k1aq+RjWSZgYHlkMkDXFgr9e77H
DU56uAHnCuJ3cl4GCw5Io2Sj2irDQNrqonhztJ3v24b1EJZXiCc4//cvP12Nr/tp
4ESI4L/qEfTKfRuVloNcoutcyEgms+cXFg/U7KlMIfG3IlG7+5KUkz/GvOEk4OJk
h9d99Hag9pC4zM2zifaVk7b9onx6UgxFYdv2Ozw7isc70ovGjvKxP5gt3/vt/LwD
6zayLWImnTpg2k1YWbDzHfESElphAGBJ9sDINjKDw/KnoSh6xZ92pypJHauNpXKb
NQ8xSQjAPz4CzFB/7nZ7Pdc0esEVJt6g4SxB3EVVZCypxTr6dHSIY3NUeTUcZ0+b
3LynSgT8LX04ZdKvG2VsQakdksCXWd5AwyaLEY3lKJ86EI5xEYuW8lws/QI28KMD
k2Q78g+FTFtWx9xLvyBr8V378QzVI40Gpg9T3+6rqFx9Mk8DPPgNQ/VAAm6BLhe4
P+HaKhURdG4TV4vfywgSepE3j/g5cYSW+lyM8GFEnGJaghhXUAm6ueVASSCCWGdZ
LCQxn7mIzEVyYbPOGtfegCFP2XrD27rnnTZcCUcjhp8jLEBzwvw3w6/oE6TSSZnR
9HAXaSzfLdbLhlEJ5JtEcS/ZxEyz9zKff9kxJHAzdGa8Lq3SM31+jnhyX5Fa77bL
VmFL4swRgHQL8jkRW3OQYjvF8bWahnweBqjvf4nr2cMzf1jrZaR3U/QETgKVF1D3
i07LBdZkbc8aJmxd0DxlIFpG8tlvuUDa8ufxIF+Ld7Z1JCxwWtgZAVveYPcwwcR8
IPiV/X5xBO4+kElUMNwUGycE2snbdHL6c8oRkCujMeCfGoA61sZLF3VJrsDwCSfC
30A0qGxhD/4Ptsu0wgdsTOHkxj+QQO1EyXJ7r4HIioYu9BXwhcB8YP53V4WJ7lSR
OOjBY+T95JcIp554wcXAY7aqZhu8GbLauYvB+hIfPGzcGgOrIuSaTvIhISYPH9rV
DYbs76aaEMVpm0JQzliI/VRoi+lnWa6cClirUoc9a0m/BDh7YtjsgBzcw3XeslbK
scqrxkG5l03LaeLTwACDU6Y5EezBh6Kvh/rPwbJ5TigKyvxApfftJaXpNIfdb3Ce
B2zD5OFKREU/uaimPPRknkTfMzMkoandEtnqWatCK0L8cpSo1jU3sgf/CWsM5zZF
E5pbwca+KNzIRbAzyBdeRd+pzTY/n143G3EybEC3NLZyaSiCD1k4fX93inMBXQ0q
zq3sLkLtUgy8p93FkQXg1OBxczZeji1dg0w5SqLhZxPFfIqYAc1Erjzb5qnUG3Bc
qQH6QH5HSlcagHgcEpurRu4aaie7DCjWZLdrN3Y9KVGm94RHfWEiiJGf9uoJw8N0
G5mxWYrhuRpxnYchVTupSnDSybTnb1rt0zpBUCosrTj3UJD3U6pGR2CluwSjb7ZY
gvNmtIwGYLdqYVEOevyzuzC1in7LNR8YlpICFmrNK2iaOHJo9muhcyw6G3KRVnjW
Z5IfKiJbr8bGxuk8jpV0fiQwdLfTOu7vqs/jKr3hrTfVES8sg+1RFdMvuzp12+53
E+fnqrJAspvSN4xyXIYBfi2Zo38AC0S0hBYMTF7qB2M0Sm65o462g1ogY2+b5ELU
9145K+jEYiv3JHScGZDlAa3x/k3utmevB8jbTJB8O1Soq3ZdkIGlPENB/lw5Dgz9
7JXz79JlKwVM1CyiiX8i9G27Jy8ykh+y8PZgElcaHwo2PxTBjlWtniZ5cIM/tgDP
QorIY1RDGJp1zQGQhLY5NGzs9DjGq2K1GWF7QbHKAAho9g0ogaGic2gHUW7evJST
9ETZ3Gpqe+Ae2o0XCXM2WLnZeZzJ/vKd0q4Mc7AA1zJiBrHnUxjeXbc4Q7BxJMQe
KwaaS5BmkpsJgTyIw9IkGwDpmQTc37xB6CYfH2gUFcLhPhpDikXxQOxCIlauRrPW
OWvoPikSl8suPhrDqcYFsRftQEmX5BSRveV8UocYV7Bm2/JPMc2e88BYmQQTHYHk
/VEaSEmGdL/EC96S/qFEs2jxGU1KKTypprLKm9/1EYiE1g0f+3pFEFySRIy5tn42
N7SRvuIZsXoIw8piu7ZaIXSeQzKzvDrOUpO57pm0r1suZ4n0e4857wVo7tG5vJ5N
C7asJjeFCvHlZupzqYCpRaWDyEbUCH1XpL+vN2xfNUwII9WlLHwJbAayKj4QRPde
luJatwYzmCMUqBIx4nUSk0uA0LeiT9KvpBDpKU+jUCFTB7XezzMPKiPEnToT0XFB
6L4mmGUKE9DtLtpt2bGwoFWfMOt5huap/92+a/WsYWuq7kqJ6TfGLl8w6C+Xf9gQ
WwTA92J2bWmnr38pYJJOcLmmJLEbZ+x9wGoKaB/R4PC0dc+RSQmSaHsNcFHBVOVe
xVEj5IKdvjBQkbzzdZhkjf68sat5IVf3omse7lrkBRhfpjdU2PSGMH+n5z+wAkvC
CyXPMq40lPVVpejrYYxzvekFE5T/So/VDi0+UZ4b6bVfA0QG0nlUs795Htwhw2Km
ggfwNYzqcPw/AhoKy7l3kmMHibN3MT8Fl0uGwq+Y/Alo2mV0cFSS8+YZLUnHu6S7
JT6gjmAdFTyvCffatR/CO5so3jHKce5uiQvDE22LFfbGKqa1f3ZEtCOAcqgnU36E
5zpipjndm4ZIWKq27SAAnfkIbjMhhQ32Z57nMsMZ6+qB23e3r0Nxu97zVeKBKHED
DFN9v93JWNE1FKfV3grrYH2x+uyki7iE5GDp/E+F5teRH288GfuaOdtQayD3IzKN
49nTUZXlHp1oQ9VFrgHd+ko0trjYbf7Sn5w61W6XNMiLqIfdyQGPGLRC7cbkdFTA
uWT1CSuM+wkWp90f88sdEVCNt3pr98hhTfDieoGMf6n8VPItyynlS1N3sMoiTC+h
JLl08X+Aa9In3lhyEKt3UQssW3/ubxWsJawSx25VIg4fQzvctORvbDIryHs2iBv2
zLuvcuhO1xBzpIy3p9qDMMEoIbKxL/YQbfRp3wV+Uj0J4pYbtqOFmIVNdca5zp2L
V7FocP+hZgFBHgZDwJUdFzPTvvJwbCe434elFzkMEdQA0MuL5AVjNw8AxeKYhd5n
3cfQP65VqOmmNx0QJt/e1zIyaphgu916vpCfJbWmDj9i2LrcNitliDcgUf+3PiAR
GPbkqIz/JInRilkk3V/ktDmg/5wxE/Gd0eiPNpP40uLBd6x9W+H9Uwy9d3B2oumg
MqwiC97zZSaSybOLYysICE/Q1/lRxYkLtHqHkoFaFv8YTYNnlPeXPXJGRUcfk+SK
9Ds+37fe8KnQolxP362yum3ACmXFSYof2RGE5KKV+HGzE8x2xIIO1v836uZJL8As
LjTpDQ0U+REswpiSOX+l+CGKwSh9OcOpdeFPqUJpeWaCY7Bg2R/G4+PSF/1WtcVQ
aSZkkQweua2NBfAVxLwHKCWx5WrOlJUCnlGUyKKQwrNsLvZpemgN6do9EaIJfLmB
sZfGMtnARW3vvU7yZmfWihJzB4GUPBfsxzXMc7WXQ7VzqthO9rUwN8IZ6uY9vHZT
e3VqLpPtV6DF/8c1seazXHMo+Xp4jY871SkzP3SDAfws+rtflsCHvLGseLlbdZj7
8YREpr5iBvVkhDs5O8OYnuPNQw2lQCmAZUVCL+uJ6qBdeujpDryBDUSSeuake9ub
zluKk6L+dO2+ARdkAIZjGwKHnGS1qAeNPRw3EQDkqKXCd5R440izHSSSnZLDZ03b
vVDzI8Y4N25/qjh0GqR8LfdWG0vkxfsK29CwLsMO5UmNXCEriZ4uePWCqRMECk0/
sKvxctb6c+d+RwLGIpXLnyzSUTwBQF+f6ObnwGEo4Zmk4OlaL6pZ4yHQYZ+SG+5a
wUREuYPIPRtHxBsVKlmZUZXARrml8s5Hk6LKv7GR1NWtUwIgZDDi5wx0wQM4sum4
46TvlebSNEEBy1k98zY4ICkrABvpxKprsFdBTLCcdkrLnwZdZoLO9n08cMbfEOjH
/l462/k9xlbUiJjYFVIorKIVtFuHURaAHfWDmZQ3sjNGibk0FKjohb3gTXZLS0fU
dPfhHgnJXGOXWNdJBhb9G6EbZBiiBGz48pzZfHEH6R2mkDPpkxkratdUyY+9+GMS
1Zcn/gg84Beigj+dz9kvBr423mHeYUeM4GlGulJk3TLwCH1uM2T2vbEW3gzXB284
H+xZAgzFFVkGTI4W/ku8eOZcV+N2LPSQnNnRA7ry2j/sfHNCFMzDLx+gBaT+4BKR
XNSv3MaCfRWzg2mH1auipozDEUxBgFsWZQwX/0UuAGuFXPC1RGgBOhIuwR1CWlsK
RjPRwBhEbpEwvsGXVaNKkOASAM6eGaFatKEwxdBraZd0x1dGzAXe2M/4FRSWgqy/
C4p1pwq8GTWijIax7PvXDV84nowa3AjJpjJkAv9sx5Z1qso+8zw0UG7wov0wmFgk
x8ItzNsY9hr5P+5IQEZ/5XYAID3+RSVPxsiyvCVCbzQvY2UjIm6181rHbm/V3ppx
Ls2iT3p3rAyIqR/3+ZnFW3ITSH7DmUrx0pRNLYGrkbBGB2g16bI792bU8nXob9du
WM2eFRcPq/Gl8Lpq3L/uxq6Lzh7dn0DhlKoWwOt1yKk8xEsVLSLbk4Tz2BqVxsF/
/KKxnb2FH3vcSUfxZdLjUoWyw0qzfO4z8G4SX1/RGVo8AVPw3tbN8xPtuTkAbZWo
WFuQBHi5bmSK3mLXsxornUxSZIIbvtn7+PKW/+fcJdq1qzDg0cB4lv1gk+hFvCU2
d/i4iBPY7kSnk39n1bWrYajA8GRwBQv8g+1IagfwIyY9oMVtub2zO+v4KxuuTCar
fuei3KF+JVB2nk2qXKKZpYeJ5TbvWwkbXzk93HB2Xck30QsHsjUnoxGGjb/t0Mhc
pHCu3LTwWygvLVKrswbMBZsPk1uyomS0Z1Z4n7ffRPz+JqMWHEjrUHCCOZZCsz3H
rKf851gtgqg3zdfJexCkuEmAB/CaSGtwPRddep/4swkxjtLX63U7aT39zUMAPsdU
kD+JQX7BoZ9KJ4VS+d8XMJhK9LZAlZOTBl4YeF1z/QGs/xsqJxBZtG6ePqrnua6O
dn1m0tVhEvJH4JjWyCPP06ZwgrqfocvUa79SzlbmjYbDGAgfOYC3NxZMrXsiqH8M
y2Zv9A10OzoX2WSbgry4/b3SEMWaip5GCzcnjptNMuBA2pil7kSaO08xEY6BQbvm
LdHH/k1Bwo9FsoI2OMNV1ESA9LBwV4Z0qxjfDfdF/oTtVvGk/OMcrZ/H/u9KwgC7
ZNfQwu6xaUNE7nh7dPFuNWhuGzOnX6sgpUkt36CvsVcxaMS6jf7ESR0kGMLhGHkK
C0xNztBMSiuYuCXeUbcg7KpWO5aHMo4aDJ1zfaBP10ZF+6PvToKhCDhysVXkHDoS
wtrHOz6cR7U0MQ/z7K2/krDnuYjRFzXXai/eXKfZar47IPi7NOs8n25PpTseoobq
v08sMoJytOSrG2A4/6igY8pyYpNpoo/ftrq4H3o9EEXJG3ys0hN2/4dR4pN2PL9P
uN8/CbT2fqbAmb5wwlaIrViXIXC3Dr6z+pEG/4gH2zjq2lHwhzUtKtmCuhmVb5lA
LcFvZuyLbfL9lqRzCzK7KCHLP/N7I6RWHmxFb9n+xpm9LXddVX08OzdltMNFNGIe
G5+sFn1xbXbEyZi0i+y4wfYO3uELK1oxZko0iOMoTXu+1a7TLOQIDbpQF6D8R/xk
e7hT+SYNBA3ByrC7v5nWLW2X2vBfeqf7/HDOdSxfhtY3zd8L9izHty1T1msuqUN2
h8d7c7aLr9cqXhQ+vS7xp+M2+F1j4jexXKMvjZzltXsFmKUovETDrUVHCkL+z+ZH
XyZpeMETdb4aCYmPQXOO5l6dtKZ0C+J1Z5P7+CZ12euZYSMwx1bbqmFh98cLeiBI
+cSpiygK7D7BVO8MsEnVOKLPmdBoutxifHuuVdLHW7Yff0izVh0c95rPglgZyKei
xCyblFFqtDGfygI/7VOMWWGknMwBBwG5iefgesg6lAKcO9trDTD4wZa9ALiqOYW+
Rei74dvwqFfguvi+OrlyEDOm7kYcUp1lV6oNMKZRJmcebxFt7yHn4nGUcPOX1Za/
nvnTgEfx9ECBCpVQsyX9yGiTSjWilfNplqh2Ktl/RqQcpcYsUo+BHJkFyueqHPAM
OtRv/KJxQ1Y10nyGG9TlGvkE/Zj5JqLCfDzYh57UjsP5hdT7fUhzx0ZJ9yo/t+W3
qIHTeERmBUZ+sgBvSSrqUpSecjnSdIUra0i/+IpRu8WM+2jDtPqpzr+5GoPqh9lZ
m2LfUfw9VTKrrlQVJdl/HzCDUbUnZdMMpvk2gW0l0LYJb4rBFA/zwp3wgB1zSuo6
CTbCJBboenWjB3N6brP4SJOuz00SyZj+TnAPUqOKSjnArjqg++iHQYigH2uRoOCh
OF8GW+lQ9FrqDZisFZ7VP1CstpnIAYA5s0TqAKceJEHocu/uubxPjr+R6qVl6Tcc
3MKCuGHWvzxyAojumNUTjSusQ96vuRllGerT6K5Edo1DtJKL+qRzugsDX6R5nfUA
fTMLmilgJjxN7hyjcuiCM3TvRmA6wAIlvfIJHrHgarQWI64aVt+1HXckH8dx2shg
vHVGSwgfeYsYSksrXK0Fb7fHPjaSlYC85H0uGoaQqt6aKTaAaVeCRvGydRTorEYv
85SU/cDh8dRqTo+q5FtnVVtwcgo3JiU2h/4go28l3/1n6C6S5NHrMWSpFThQ54mS
MRBYT5+2SvyRciXbiNb0DaawJIbAdboFDNcN0V05QA8cIwAM5KfAyLaTSAoNxuxD
5PVCPH9cd1Z2NHLd7f9cQgTqSZIKBOJKpWw+5pMqXafR3jOk7LA1fiLwDZIeaZvj
PiFtSvTFB4w5jtQRmGZT16dWG7HkEIZAgQmT/RfKIVltIr4eHz9/qByXXXC2rM97
PkkB/MGYHf8ohWM/7TolgKj8llYaq20/wk0sfrDhkNeFxXBdXpKuCeTVU+GLPP8d
NfjTTx2s62r5vCxDX3CwnOZuSVNXBKQYul9zbqQrYPWyynugNuJcwnoawuyv1SL6
93RyrKMEgsqTY8xP1XUcq/yhg6whrZS/Fwq2XMB0CWA5FvAoPGzDOfUUFFnBs4er
UOAfWQ8RdkDzzUfZJh0ocmcs5NEmYDwvwOqC0KaR+taw6ozKGdR0MeYjQtThnLME
wexVU7UeLFjQJFTZX9MOCKvxFoFKH/8dsyRkZqBDI+ga1vZWR0fJJN5F39RtQN0e
A5kn9j9ADHCa9E+/x1JAVYyViob5pp6EUS1LavDstP4V+U6x7Ik+8ed2gr3rL3Ju
8O1z/Jwp4ty2eFaUJm73159vzuMQi2HmFNqvDJebxl1A9+ksJtkXnxe7m1/k6Sg4
HZgff2biRPFjtshVNnjs6pCFHE/DnM+/bGqF67S2zu/R66uD55CRAWZIzyKq+l8N
t12jfS+f6HcJ6n8zEOROyPCsUMH8WIthDFxybcUFMUAwNLXiGVDyGyYDh3Ob+R2D
fFCYhqUCQM3XaQ21fGL03eKHYVs95KWwc606o6LBS9a3oIqkH/2E3LMRj24P9pTC
Iu6lPfRdmDmLrwoFcaTiGw3LaA+zmbiwHFR3zep+ugWaj6rFi67CgnbvswJr9yO4
bSJHM07Zt8jRh26SDx6zJ2J7pyH71tHN++mQsvyHPOL4Ti1qMX9G68CICETIj1dV
1qjWeNEAkU2h5XOhaTuBmuuH610oIZWcL6nsYV6fv7icYXFHOBWRYQglpHl+J7PK
RnihGP6CiM43Wp6vpGV8jQMpdodj985RPNG5R5Lrx4nUVv5HYzd/NOzz29vUvGqV
akDB9L+CaO3mnYqstxGPZtuNpOhp/WtlBMEi7rxYqKGuKmajTRXghdfhbCBKLlDk
N0WvIjqi3rUnfPO3r+C6Az5bz4hZoR/iFLDCrC1yKRiict1bDaufOjsVQjg1niNV
R8evCiaZpcPjdVq+rXRxLl+SjaoRPTJQGZqcR5ejSG575ogUI9y56q61XB9x/DYA
7pIUmHfqEILbLPDDCJ11j/AX3YLEQ7LbtET3rtOedp/FEv2q369cQAT2OZVb6LBo
P1wjnHvH95GqlI4qd20xhX2bwffKqssG00iwG+G/0BLBqdrYEE2UmW6FyxYZGo8e
fhvNDaEDyt004ahcysPG0Ka0uzOa80mtLB7UJ5XT94Kvc1n57/8vUfsIJevGPBzp
K2svkoE8kM/bm0l0s7m6/VWrqzjilgsXwtwzKqffORsyiD6r7la9+0r2Zv/8++Ap
XmwZjdJjZHult2u7RVoBfbo8BzBZjnTQx6qcjJQSyPi/+YGJiG9Ox7/w33QhaI3Q
y+RNRvvFIuCzRSiyGPQtWcyCDXuhS2VmkY12ZcsH9OaXnkD/3vt+B5s6IsD5/aF6
7j5u+xCNG3160g3P4wTtNYPqJabfsLmFWTM47zIAAtVgoGeBsWgD/OYDzO9etEE9
uZr27FSTfzfcghOrmp51wWRr9QSKFyz8ZmC7NiGhHo1V28EoscVQO7fva3hozotn
muLcWm2Z2vofjP1cKDrJ0HxkXEGcTHrGkZupauCkkVGr8CweFpAHjkJpZgB++pjh
tEDufLrEjzbewRPFAA6jrhfQd5FAnQRkp8nm8m1iMZCDqCMiaHxsucVXAkqBSf0n
w63MA08qizotA53AjBsZAcAMjxR1b0/23nf9r8gb0eF0M7esut8etLsMI6MVV+nD
LVAz8iqvAYL4hnsPjwveYlJpBnBjFOZj3lhjRZ4Wmv3zSTDiKn5ZAo+XlsSEfqaZ
R225fzdHrbCQ967/DOYXcOFrMbNWBNhu6UGwSps8VC+cXaHy1FvcqEPu7rjjXXsL
LiSHO+VMMU+ediPMQD+XL6frcWbqCd2uxtPjRZo2+ieIIc6uL4wHjzXIdCciiOVa
rDbuMoO0ScHJTL3/3c1A1U44e9Ks/kdslw3J1lUboOjXjJztdQ3s3rgqq5f0DERl
2H8C6pIrjKmZBLrNdy8sQ8Y0CjrH5w942nlAdv5oEPBoo5MJ4/x52SO/4YrQ+qM/
wmYcAmUThWaJxJcbMpnjyQMQKoQrx5YDf4MIGnQHSpclM8jls6sB3str85x7cMhf
vZgHyzYTMzwkr4s7NTek0oyCArOKx3cRbXePUETXcQ0cY+lxduX+rG+YNdmqIeTa
1oybRupcmz77pL90czJTqJC0dnh+fwqKNKdc68JuUqFLsiIvBWPegXbBGmiIiCKO
wLxLsPiwWYegileYI0xQumQO+RF+lNTtlVoHyqp7A0lor4yxILaKlQk76jrEJe3h
EmxWN4Meir6lRzh29Orw1k8hhR0cy+XgS56rSeMcrHK+XgyRouYoyaVRjKa2fFhX
KxLmuX9d2cbSEGgJ0RiGYmXefhDgb8sb/3o5ESTxrKRP1OjUlV2OBlPwYoESDIi6
BzSJSY6NZNoSg1J5add2IBR58/kFRsV1P90uJhcAZeLeNPXNoNccLIJkl6P297Zq
JPLh3MWtsbribW5Mor9BxNNPVIsde7t9f+rNCtClbVHxt1MqeusT/YYYZfovqpqP
B3rr1+toPcZGXAnKD001AZ8tCIO9YAloKK5/bTqFG478ZZczPzElwGyN7m3F/lej
RNCyElrQh5q2hTN4Zid3vulYctaIInt+56AvYyxgFvnax1Fm+fOcHjDBgqtgg8TD
peWYLhrqN+OXU1woGpw8SnD3mgc2+8aWQGirQyv6rC5H8VtZcY/1tRX0zrtKhBsc
mfpBBSVKP2F3bHYQ762sgOTt9d40R6O6P/uxLu5CuHQEAdVJZmOdHqN1XFgDE9Gs
HZfggJt4uKyPWkRLOKWEGh4iocCPeXnWGcvow9wDGRHfIXDPUnVaaJSyv/ujF1Uo
dz4Os3EOeM54xn2o+6f1+NUV6nBFYbQm2Bv31+LdNmW3Qp/gQiTa4toGaZD3fnbi
KZzFdJ43G4leuXF6TxWryA5g2/znaA8beK93A71jPblOEO045czOMpngBl3llf21
06RgxoDvUaY5lnTSjb47PdYC7ltkhnszBKIjpkHd8iNAtb9YfwVSL9Vx4uNJS8uQ
YVyrySB8fXmmeBrayU5y+/NjpP2D+50VcNO60dGRcyWsbAwBfT/+yYSjG0xMMLxQ
/Y4nxWw0k1BhKs38SG6HzSmZCNNQDSCrdpGrz7GV4lAeEdKNqcLRpuItODfCDDWr
j3iy8v56W+njbkNowBkkvL/BbdzxsuS4QQybEsNZ+NqWnx04kpLBWcfyB7kcgVtz
LfCZ9HlTGSSPU4mTkdmsYs64FOoPwzXXGQC/iZ0Id+SH/+NKPf2kGwonTFkvsbsW
9wLuWJ0DMvTj48wI+o1OZGRCbn6NGIwGv6bNY9wCgq3hsrkoe9NNw5xByR2vo648
SFWWFB9oKquweTlPbRJlsT5jeK07hY6sOJT54p4b8mXJN3uwvDeQvyDinfrjGN0/
nrZJ5hC5Dk4qVYab6/AP4ZDY3YpulLe5QJwlFarqzr+Ryks7QeWr0Flc0yl4rHnn
soM1votXvJ0gWBvUo4TqU4oPcPB7tc6P9Ot4fYsD+fz+Cy3oHzHHpFkhjAlqKJni
IxN6PfBHXdU+sPvqOIafxLU8aB3b7awBE/LSOUMfbANhy/B6WW/cH4Eg3P4QqyVy
VjfEY/bOSD1xBLu43rSCfoS0FpMcwMXk7UHKlcfNzCqq2c5gS5a9cW38IWqJ9fxB
74V6mnVAe7muMgg6JfquKKHbLcsm/IBa1cXBR3q6DNOgSo3ctsD6mXOgAWck9WwG
uU9FAPQPp1zujlipMwiZyojzBERN1RM/FU76CmNocMTH+twufETmQBsm474o9Ga4
S2xX93lEnpOrH9jmHb8/Wkzmwy/fgAMuYx+m1jMYZq7AaSROTXBMvOH9QjfWYA49
iioHFIDVBpH1aDpkZaPZmyBdadCHjKUYKntNVEQtZ0UE2fpVorrACrEk14LZXQ9Z
c9O+oGx6w4fYKb1yH+rJ3Fl9g85nL5hd1TXxw9IYREqIHEJB6cxwwB5O5VSXYOih
Nj/m8FFl0GmF20b/OgGQviqRpncXKzqjrbtogVN/j7Ym9TS19hams68ub+2bOxKn
FFutTUph2vvhD9+EvZex3MbgqwtnEV/Gm3yZCZ4AZwJmMEpJWTKQ8fxk3OMY5P0i
dVZQqZeKxi4MixcQAu+djz5Y8+sui7ZhdIRaV1FryDDWCZVSD6kdbdpUhXoqKvkr
+AUck35LMmIyddn8iiQcK8J4wO8M8N1W4n6i7tW5l1MfYQghaRpMfQZfifYn8q/6
I6wGvjkJvL/WZwQLoXgdBO+KieLbdn44AjYlop0cSbRTvX9UAYdLZAaFmO9QzxFd
SAB0wQkIabPoxD1LgzgKJ5m7Q97IBrBdslM8TS0HWLF/WaDDWU9WN0TYxqIUauxi
hIox+mY4gByMnKY18UlzxVSQ0CCeL7/ghE3yEZQ/3ScUpCczJTbUKtGH40N4qAXx
pEHPi+I11q5yECkdBRJ9K7Rf33Xg6TDwclY87D83VQ1sfW/NkAUfr7B552mJU8Fo
kjSAT/M1txLfYbULHoz7bi3ic+fQcvEIjEuMHQ2rQ/bL7mfy1pvF2CxOyB7tZA7h
SW9GC7DVM18O5KkDtCRDsz0B6Ut91/ftnJB4pqyVCf+DkPVqP+IQdmqpbNSlyeI9
cdbEkYyEkyspLI+xn7puQFWirFin6gMIoLH7CIprrbwLiUZjwfu9I8LuzYjbLmuq
j//MmEI/x1uvNji6mSsIWf0l0ZjPH6YZNyvF2cb9Ye8/FP4WRry9S6KN2rfM6BVu
fbT7/x1X/Q7OYD+hCmf8LHjzJcQI32oIzpPmduMjaGtXeZSAsL9mi/SMVTCjrJrk
II++6Fc+GZPDf09dA2at/LTz/x1hMQMCHEX7FB0WM4COXvaxVkRDGRaCz3JzbPvq
oywTx7Aewfd6pQ5sZkbgImXIkzeMQi7De4qvariEfznWwg1apU7/n5KbduJ82ejl
AWhGd2iq4ChcJ006qxXlIbpsU6W6J93cao2OACPPa/tfQeqsL7Xp6S+7mC5S3J5h
KwAj0qgIkC8ZFuZYoFor7qxa5tx/3eJVj9eEcjr1SuGikTDmtkMTAJLv/9bRfVAA
XbEDim1hoM8MAThZxwIXqKN/vYk847sTss/PA0abh66lAJskEe4DoUio4N16S3OE
S5bpOwcjF/PcxG9i4ObmEHYRqlcarfp6wn/0voHAo0IcIlAivzOSAo0Ft5Tuy6Qr
eTEOE5B4v1r8gghVsE++kEGipvDmkumpdCpginA1nhn6E921UnW8QXvfL/CKC5Fn
onZZuX+SuIBCLPYauXLg1JMhGfBksrIECQZiaJgExkmRF+bdxe6zPFQAZpHOuvzj
7bKUcIhRK/fZMmZev64c3hAOsn2oB5SE2+WSD6/EBA7uk17Dk6yhd0kaZlWUEGJB
6Q9ER+iIt4NysjqF4X4oKiPSaNcl4tGQhd4MT2Q39RIXJYN+0qeulM9ehXuuqNHg
fYNGUzHk2QeefeaXR2jSpyWNiS1qWyTq3jBVhTFq4ebAiF4Z72B9BkQ3PlKPcaHA
QQDe3W9wDoq7RJ4p978B5hrkNU4E4TaE7f/Dv2QX2rIrnvjshDra8L6nPvNFVRdI
GjHGEHgrF6pCIr+G2/dJHJrd3aWoel3LuHOBFOXGFRtdMpI8LgezoFPks4YVG1ml
DMV7pXqRg94/qPj9W5CUBuZDIipEshiTIB5UGMOdeXCov2B96/pS5H+aPAF+Wr/5
Rres9Vaylw0BeQxd0Ow9UWsKitZwePxJqoID4O6eSbIeNdxkqXKfQhvhqpa631bX
3ipaU175JySATJna85Od+9bM56JzqTClTb4JyHQ32Ib14ia5hGJ8yeb5MXZZv7WI
93AlpUCSLy9fux+xSQmAcnqvAqZkqpDIXuR2Hz24uczU4OqNppCDgkEOmnnkcYgq
kDN7Remv95UoeGm/PyySgfEK9uKXEWVwo5hyio2/JBOJLmFM+/055Kvk+kvqOM4Q
j0QP4gBrHt3B71ruOG7/2rQJEYQ1lW5Cd8sa8hOP4sRR6QUHMSDELckR+uQwTxG/
kyounllWR+wmVAqHxgBWn3wfY3zd3BtsZRjzRI90iiz6Qiv/DR656Ga5oFJUPCXE
SwRV8Xr4E68FdWBz2i/4lbb5qOkdkuz2h28O7RkfWn+RAdbdEdHzFTgltlojOYss
N3lf+1kalI9tiOx9DBnd6NcFl1FkLSnVhqxQcTBOjWDLx91Et2SWA9OArPT0xTED
x9Y1REdsGVKfzcds/vLm0DJLBAnzckudy0R+AMYkOUo+AaODBYBry5xFkKZD0DPz
/f/0YGiLIXOHoO8aedGzh9Vssk0SNyEahehnzbIwbVqqztsIRNb8JdCcjDCKZ4l6
V7e6EZ/HpPXmiuTa8Yiy5Qvq7tVHR2olXroqeEtkx5t6k5DCoOOF7gq6BL4jjoA+
tfy+kioFVAzUgqeOSP+hsFT1DkFWZ0lX0L2DToyAl9pZB3758gDbZkH5SM9eeK/c
XHAtEHtj/TFkceSLRWjGVd0LM5VDxflqvB9rFvMI0GbgqHOMBXa4XQg2cJLvp12A
371tNAI7nvrrcg9eTraJ3/v+Mlcm7n3am2ogVr5f+yJNkDZTQx+o3o9wPph8FWU4
oUdVEQL8+5TbNsjXUn3lAVX37nSSFU6asAcIommFyA297wHf9DEM6J8XhKqq4TSP
m0lqBnkjB3508Rn1VGn/dqBcGrXrGC8FYwll9KeQEk+4UNH2CRKVZ1YTVNdavN8o
kMLNjO9PNfeWOdiD348dOiAunEo0dYB6mz6ZOTww3SUJBKXn4tJgTcQh3+g6MGwm
BS5QL1ZT5vc6xrZmyN/qJkDnGXizg5g037qtpwycz8ZTJ9wGBO4e94HIswkqGiSc
3Ze4EgezhVSzcs5/sb08P4MOz4p5Yyx1+mEaj4QFgdIVW71Y3C6yqLsLlAInmAyK
pkIDIVxBCQb9KJyB9QQOWemF1FkQD/E65KQjtlsDynUhiuHQxVOe3B2s+y+grX4q
s2qRrVjIzxjydgMRInKmt/CRz/i6nlcmuSZnO67liYk5sfXgTWbAyDwlV+NZXP7b
WjiGyU8klnYP3zgKNFsU1GIsbZXQyOohBeIs3n/6scZ1UcUv8WSg2+OPcWTYRQDb
hOAmFEi4hp2AVW4U2PtS/i9keuROjnTLGSUU8Iz/Ciu1XQP2emPv6GKCMsbubmV5
DtbeG5FW8a/82WbOhin/1KllL/aIXyyBCWLHIBKewfnpbziHfCtyWkuaQnwIs8Ha
epXoFfCdqSKvb36j54B1VbCMgPCrpiKmhghpPJfRdlN+YyMKhVXXhInS/IQTMKYO
TNpgIO/MzN8VAFYrJqCm+ewvkkCzeCc5vsyyE12MCo8PGt6hwDFlL/i1KuS1pqV/
7soIPkMVz4aIUO+NlItwtEK4lEDKlBvOdV4cKBkNyrM1LWqQmej2we5nhYJeISos
y5+o5+FZinI46zL8drh+++iPfCbppFtgvjqXAUsWngiY82bxqx7vv04gz7sEc3TK
xHTUs99E0XS+84femS+URtkou8i4+eXkf6HCBYvqd42LAuy72bqClIWMl2fM97Eu
bzQQEvLKcGa+hZRjuKwRdbMa8IhKUUkzhhu7QYVl5k6NcMTN8xKsGe3E7od+mDE7
rHj4nPhz8AQLJbmCR26e02ju5GsXVWju31vrLQfdv6dC3g7UF339r40e3WYQIl7Y
LEdVvZ8V0SiitVZJbtR8kUERHRKC3RWZaPvSTUb3rhBNPUXvDkUYY+cIb2NKCAfw
AhBEXR7nIKzhcJMNBsw8XyMN4mSLNybGy3c8a5bl1YT43c8GliC4pwf3753bvMhQ
3GRXbxV09i7uW2wNwRCJjUrhCJ4zxqu4cfQIsm6Orhs4euomb1Jq2Z2As5QI4sMH
G6xQLdbcsKyabE8KJoJme3Gke3cNQyiCBDIx1NbAawKPsyZyyXcKlpWkZzzQj3LP
t2DxCHAyGoa24RUZLtF5W6kNdfoiGdHaLnxN6f74YGyt9zWYiiYdGzflT5nWckMU
1/tfRq9snUju6rQlsp/HJUUB46JOIZo0hkTRMsoK2df8fLLaEDdK8aeGhYIZkQmd
jEmW8TuzrIJ8mFN78xXF352O/mOXFtGIXVDZ9HG0YLGl+8JxEFUWHGvOjmFOdqDR
wIw7ZQK1RNVjDrhlt7P9A06r79hXREKaZLK1y++BrVv//JAESMRZRdsbicZdsgYG
LFuK+Bg+3YdYEA6u254s/DFjv1mImuAWZL5dzKQSBfVU2hi9Er1qemJHhCnALWW9
2WLGp5b9iHKFJzu/ZoWlse2yCvUCpDAxMQQvAOKtjFjytO4i9Yv0yNddN+erQmc2
l+lsh5MCTcd/Ztp9olaFy+X+qTQKhnFp8CbR8IEEus6amv3qeRo7woob6kkR199N
jCpT+aDyiXfjWdw+i1jiH6HZdDqiQ+5/2nvT+PYUzuSkHi1Dl/ggF3qxOZOUaH8u
PHQ0p6S+fWX+oACCbW5mtA4vLjgH+F1OsAc639/sJtYUStRRjKtZuS7ryYORrw/7
ZCaQosR3F7B3hA0ZeKKh0+fQM8rVIcAFgxI8caqVJtbMqn+BAv6qM1p8Np5GXQXO
vQ5paW7y2Q4v4o5KlavM3Yr5qMRzIAeSjpoPOhYLWrykBcniY1Sxse5HEeMckJJz
NSkaki6mj9zEXRxojL71Gl0gnreMffHh66Fv3nYmLDz2ZuXlqgX9/rriPlvSQPw+
w/coYWSnnZCO5UUzK0wv9yoHyLfCr50sctZuad4yVzT7M5Tkrx7w5/FYYAvss2oR
8hTmEkaTs0VDSzE7ipD+Mjdir8iIvjxgLY9qPWLycloB8QZ7hkIzI/FhV/ulvzOA
7tVke+WfgTSeU4T6l6C+/+8OMoZ18y8zfx1bhnJUVW8r9oyLl9bcFT7yXFKQvfBz
D/dLr4Cpdqyiin4OKCfncaQ6J9Ex+wH/alqbgESlU4ZSGvQWhNhaadKkdLponvB2
4KhJLwCiyS37jTfSfTraJWeaSSS0/LKuGJlStnnuPpFquC9/DFvodNm4m5X8m5LH
FFYh/YmrOZJc+inUWmb/DdXaPlEAGu+9QX4mJdmc1FfODpz6+Q3y/XXRlC55fGOS
NeToqL31kW+vyC8UNTfZRf5IZz0bsFrlBGTbJxH+G4HLHcEtG8NN5JAT+Jcm+pgo
2+0GaoCvmDQZqps1kDcyxn5rfVdLCNs4S/Bzxju77lVyiKjBeK06TjkW7b3oHG7e
xTHnZoFUMxVsqX9Ow9ohrghbfL64VFJEZmh4Q5eJuJhMVW6crYQzWVImwfRYmXVC
wUQLBSjQwZEkoymHAP6Lp3LqbePDiIKVF10pSACbV0qNhZLUKgKF7c+O8yLW9htQ
Z3qadG8c+nJVSOLWaJ+epi9u0CJoRH6FG/25mNFopBFc6Ex0UfA0XB9rMDmE0ZuP
cGkbux2T0QyYxeIr6pgWZGCDYdrp8XD30p3o4SbWV3ODMrQtcTklXFjutayOBO5p
aKjZ/M1JqXnut0eo9RGm1WEPy/mBbuu/lql/vmZBcK3ozrpIE2AUMXCucR58WILl
Vpw0FwUK/VbC9EdruWCno/NqtmWq5Z5PQs2Xq/uvly10n4jfFg03Sk1iH5GVsc/+
PY/RwQCV23HT5YP/5BYcMNGWcHiTc4dryNVwS31koC/YJbKf9TMAKB275iivKPmg
cEkQy6EOm2u2ovl2+9o6xE6afe4mHb13vte5GaE6ScWti8nfKgTHvuyjCmz1RwrH
gxnzEmt0ePpRD3BpeELNss4P3rIo/R6dXuLjTaZqgK/lZdKM97ntbriRmY3yLfgM
aheGlq108UP1Th0K2IIhkSzVOyutSgG9Vf0IIHBSLCBiWTEGCL3Ge5SRvWPq6I1q
WX0tjP6D4jMo40oeXlsIEPN84NuTstU3W4N0LtO1qZs03LGVAZ0RW8l3bglQb3Mc
xsPrl4di0i6u0jWhZ/yHPlCeasO7g5iWU3iDtnXX0HXEvqizArobOyyMXfxI9zlM
daQULhxqPBqfFQnFoaWPKVg6OGDV76QYPvvbx/FpqVMaMnSE0sQkEA0kamCXe42Q
LVlkdqNx1tQp2+RPEtPOGZ7M4JoCfJk5ph+9eMrzendzJ2/t/YQnTcVcw/lI0iKQ
FFYnD03N2xtTG0D+tsUsVpz6MjnFCsMeWDEF34sQ/Vg5KDBcX48Ryo0GbJmSbYn1
IedQCvGpjfWk+zwEicCRagG4I+L+YGm4KG2U0SvlrDlOV1r56gcwYzR8pCXHuqkq
V+YaX4M9wjn/Ogn1a7YcKx1Uji/RJ5VLOMaq1tKBm2WpmiqYNigTxntSnIqZduMA
4+EkxY8cb088FEIaUvwT6e13sZzeRwnfiSfDKjYVWFxP8thR2+5VfR38Lvn+agDh
hkkkcG6MuLFwq7Uig4zQmi43gUrJ/jMUE+UUKtcuTIUD1D5WGeYTRfOnVvPT7y4R
cNzfXyyd8wrhaWvblMJOAsuwLeK6RnFjc61LX73BfbrWVgceucqxy0Czqlkuly1Y
OZuW6fbCvf9rfFfSeB3yQVksKJL2FdNx5vaix+6NdoEsFqYsGCUqhvAGjiNfNP1c
F4F8M60MUDOpiQ5iDJVDJ/sPRffj3ulzsKpc+u19AO8KcBQv7YcgEyikeFFM/9VE
cf+xzgci7Td5Di2Tv0ntvYbpFPjl9ZAkuha/QjHqdPXGEaw8y2vhnD7RDuS88DVu
i8HccK1TddKalL3oJkbNwiqZNrLTpZbkSRvCa1uXJdhkYsEs6DaZX3vOHxWKRspb
vTEPnC/XffQ2+B1HQ1iufaGvZ+K+sXXy4TBw8e3vE3XC8FugTAKg44ibfi9vrcBy
V5joWx9+M2yfOBvE69bJW2IbXjNDNbehzzH74kDxnAteUcjQqJ/3Oy+JN5PpnaWV
RuAlkLXPVtLvfK89SV3Ul4DXyqjWIyRNhklCKI9ICfFLsU+1whjNWab9mAMRA1g3
8mgBcmf0aVEockzzyjwPr6w5pVQKlxsrqOs0Lghvnaat10IvGJAHzaXabJcy4kLR
BjJQK9FEiks9zJaaSGCSExmHThEx3sObp98U7Fqddb5VCIrNwpeuipZNtbpfhEKD
k1lENMW99LgsBMM4XfNHik9BIQ9o8tv/BVOR/hGavrRXVTit750QyaULoR7CwL+X
MhQ5n21Kz5o2ss5Tn70R21YrDePGXeYZbPe9oUeeoFjfmfYdAqt9tsd87anlFrZg
6+UX+ZFt9RR5OKRXwtaZF8uNxsKK8jJiWEiUsqb3TM7cn+rIFvUkpGek8fBYeIhK
FyioPfUH131K1TTJX4iIGme1Q+DpKMCy5pjDgN0WZhHTmtQkbeSaOIEm5AJe+eZK
77AmBzCgNm09nwg5rfAj5wVa7w4i4EhcOER1eJ7G8RrVbNs+W9wRS0rNYjINFFHY
byxdnQ9CX+Kbj1kmwwlBU+80KYqvtUtNnV9eKKhUFXe2XH5/A+kJHVV0xOhd7xGk
DYSGWjlhYZaqVZ/rDocGfuBMaLQLyfFEqUZqX3Qhj9toaz4ntAkZJTcSwLm0U56Z
Ze3sH75pm9OLMuoUzrtpj44sKKJxrDEo9ABfOROSywsv6a+0/RCyAPFDs5CN/lC3
N8iq9YpVXyQpKIJSJnkdr+B6YwzQkuaFm03e2JfWYQqNgZ8FXHCsNKKYDPwFaEuF
NU+Rcld4HXQwj6P17b0I3hgLN/cJ4TzbH06jSwBzUIG7umvXnLHzpytYJ1MZx41/
pZpjpRriVWEWUVJkbtmmNTq7G4Km8kVG3aO9tjzzGOITH8vzALPj60VhsqVlB5Ev
GVj0EZjLwXtf77ar+WpUz1066+8sFKuaNVa5KRUQBKKZ1s/7Oy7FHfXvmVE9NvIf
v/piOQzdsAcbwBIQXbXnSzsfuK7QvMb5F3b5ydr0mUlS/zI8nOfA8deI1v/mtfpy
wWq1YzjbaUZ0B9cL3nhNFkvVTYSi9cL+PZmXj7teber4dWlkCS4fkrdKBgVu6v9B
UToAh7hXaT8JsnP2TK+uuqaLMhh0StjakZi9RCqfv292jaZJgHa0SEHNDTKYK9tj
F7MnlVPrhpTimdGHVKwTdIB008H2Us1+Qzb+5bhbjcDu+Z678phRpZLUGuxFo1iQ
Z5nSvT+TVVBXAJ1AS8FbUyuFRmmwqguI/81ngjZDUrekNr0EMxe/hHT71FPKv3Ac
JMf65XfhN4XoTPZPEQooDZRtj8ynMzi4zkCtXYZvxOKv7OfgtruKe9gxEe3D5dCM
igBtZ9Km5oI/QlN0P9cnuPA89hjwQvPYIxxzP0y2C5+OoCjeI8rpsxH/+YKrVJW0
Rz/bC7ZijkqTuXr1Ken8Bwc+7fwdRfPdxXjZ6LiTDQo8lhxD4c3Gejy9Pi9OhchO
VKQTyL/op1ONjHc5N20lo3gvMyIfKBxrQtLTf7YspjiK1/Jsic2fqFgog//wMGcQ
eOTkkoqqE2cJxExVkpPxMQTpNeHCgq0WYJPMVWeMKStjo8HWhyGrfEFXbsIXdPeT
zKPZSqqqqbyVuXmcJUAbfWec4fXYK16ldlADDyoVarZIcR5SdA4NlgFjL7G6OpzL
39pqH9qMVwBjvubMj3Usb4yhN2LpuOU1OqBY7Hkpx4bzqtPr6qZBdh/TJd3fnFL/
iz2GQCdseWmQlN8jNdQPhU6bPiLcAZcSdPqctYbpHJxGU4KzbMgvmucp4Ar0yIbP
+6vuEBfwNqFGbrwW5yQrZy42nuwBbJbth8HvDBtey7yUkVxbvQjKlfrS6TqW8cyK
WxrRVhVniewiEG6Ev76zJ5GahQzH7HDPzf6hI0RpD4AsTWCUJ9ygw5nPnZppM7/K
ZOiP257XTKTWMDrYZdHbRix+zthrAUc0IQwN/Q5c2eMcQgTwWAiL1WXECc9M9aKQ
9fmngNlveVlpVpWMLm4rIzzQtG7Q3FoOPNlYZoijt6/TXglAgYrPB0eIjV/Zu357
5bvE9FunsZMpgysoxgrxGV0sAB2PpDgOo2RWXyrz+HMuPkKY6w8sd3IRGWKgsJ++
x1UUh/pf7kmNHEAlhDZ25RTrTwxBc9uvXSwZwxtjAxRxPIsXIaYnVe0Xc6BJ6GRb
7qVVNyY2xEeGmGYkCHI6qLF6Hw1tODAHJ4wEmuGHMeKPUMFptRs0iwmFUxR3aE0d
a7ei7Q2zf2aecRbLRknoOqmodUxd4ajtI5zQXquvAtsF06Ij9wbiohljMeoSDmQQ
BQ0Xw5AOslLxBxcui4LBXSMlaeexlEf/RE2PHI313Xy7tREwkNnxSRc8ZWsdAHo7
nXs+yU4Z4phEXOR+OpnoDGaxSkDxT8Mu2Ef3mx3p19BCn8f0NnlmkjrVrgFKTnIm
YEx8/cF+P91SJi4amJi0/BNQYBHq788eqi1inBs5ZgrJvxHkW3Wy5PK/JwuocdWk
p3A0Sn5bt9BQX1er+jaMn1oAqaryF4uxN2sSVghxzU9925/sKdyOF5Hpd25zxY9E
h8RFZ6UZtqouvtpKX5n0lMWbZbDyZZjoX29dHcI+6cnURiUXLdSvx68E2y/ZcIKO
spV7Ve/Hl6ZHfj1nvJyX4De2iwHDoZAXCXdVXs6kb99WFgoBXBeAEe3YMvQ8QO4g
Pqg10Tg9zmLu8bXUnJASTYKDIetafke87DRuH1QFQulsMMQDzWQUVmrYdBBYFCC9
6DNWhAw60oQs2cAWG4GsLasE/5Rm/y7scEIZMQ4jLKIY7qca1mEaS5HhxpWzOzbu
OfZ7TvCluaW4KrmDWJ6Oyxz6WHA/7nsAeg1o+TD0t/kxD0AD6DREBPrESRx7AoSx
5W/FG9TZugl0OdW4EEfla2Ju2rnPEguIFo2Pr7jD08l4h7FRxvZhKij+YmYgncw/
xtWOmFjJrzmZKnttGg0QsLksNKvSpAKiZEdrtbKC/MBrcFj1OzVuACLIFTGB6rG7
CoycVVzLRU7nBfEGcoyrdHjzeZ9nZmsS78noadpiQy0U3DFSzvSM1n7zgFQp4qx2
h49t4zruwMrzSPF8NdPYKW8/or0qtG42yyim+FamfyG/E9WnMMzidPPx/jnIeMbR
0lR3oYNP7EP6iAPxmhqzztAsTrDV9qcn8vC1HtG7gEH4mOP3UHpyaYgab7096DjY
naxt2ilj75Ul6UiC7PLgPp9LH1f9K1hW4/ttctlt4dLxIBCo2yoBOxdj/li+yDha
SLlpPg+NZL/purkQ7e1ncE6gKWwwwxiKpDKBzbJ8Z36Cw8MrjkJis8m1J147hLze
3bVmJxiGONtyIHI09WWwkvJ2ri/KBDiLN+psoKokU+DyZQg+218bwB5rmJ10GQDW
kK+sIhV51kptoGg6WizDJjiQyZDS8pXiNHmXtoMr6SpJ4MIM8vJSqdUaDGuQDIU9
Utg9URfX/RMjAOKRFgwQmH9h0kd9KtWmMM/Anu2RA6Tv/HAleiJAeKS/UkJnvqBj
Pe3/9TlV47eVkC1V6UQMf8xV4mZJ+9knCTURFDMQXPhphISyKLTRO06MZdn0R4qb
Tm82RjloKZrRWNXHP8kopp8ms6w+zGHLCTBkGlbk8O0gI4GFdjWDJFwmgP7BbjIC
RxFPbSy+2flZ2C+XRB9246OInbCe2xkZn30eWW3MQpzAqVxstyMDRIFa2aAqrRox
I4zsYnOAkbiPhh1GWML7wXgHj2cqbiIPqTaSiK4T2ksHGMPhNiod3fqQvwfPvZGx
rGEYBhEgj6oz5sqfSn/f2Yx4YZUBshOkjDQPQn7wQXBJc8yYlbVz0O4oLlJxAtV7
mD7w58YLpEzrBggy0YWNXV8Cr3rtiIaIpjD0t0L7qe4JbeYTjcUSyKXdfQrg56Dr
n6n4tpq8pubnLm8cMnFRmOT5dOFFpFjksAmovUOF44DaJwPtR9Ez0CH2cd7weNDG
mtd4G4YGv4B27REHfgux3IcDX3cckrHhdKHenrTn3UjBkpK7p1RG98Y6FuNaSI4I
PSv+khj+EdDv/RiUiTwUqCGXBxNLWfWCZ9ZzgvpgNOFGQKFIUvw6OZzbEpefmyKH
Q3EOL81StyYjEeA8PrvZyYfSzpHVqNZGydLRToZ9vrvR/HE4bKPl/ZyMFdhKK+eN
NlbzCOZYBgTGl+LXyw7+pc0HNVCqc7qDXn9fAXZGhcO0/c28X6Ew5VmeOmBW7RMi
WUDUSO8ZwvQ5xmwGt48QRYL8rdnNFUEQvUppp12sgDhOofsZjT2oGUL9WItseJ6s
M63uNeYac0nXOtk2ytdb8RbX9iQInu4IG/01AFtff9V+MV8Wc/IKrwW9bSRwHULq
gTVNaSmqhNCAh0XGpUy98tbYAPUcLXagbO0b5Rr4rigkJuI1pz40TNA7UeZx6/g0
nZODOzeFJEvJ4e9DQC9evy1Ulr3vic1LsfYxY7D3AxBd6IR7KiEDqNO4U43XwSpq
QHUAfOCYYySHCAK5qw8w3yU7rcyi1mGTEkl6J4Gcvc7Yib9A4b1YBDuniFlkJcZQ
7hcawz9uCD3EZhlogMNDFELXsfazYLD11sSr8WICQlA8AKCkFzeei47TLQ9G1T56
hJoMcoX3Mi4YlaBKgkw1Yj7+mScLPBgGiploWD2OLfh/0aQVdxEU/TaaNJ1KYoX2
a5BKO+SsdD9gYAkd5oQlrVcmuWhiCRdjZrqlArBAKY2qghCHp2iOmc3HouwDg/pw
hnxPiP9wCehKiA+yJKdv5OQe1fusHs6BGveeEr1BsIK6sp8VFKvwGX8/Ghzanmcx
BTVWvUNcnpy9w6Ny+t/EeA4xj9aUK2+cP42ii0TDUX4VOBqeo5XTd+VmUbuoRsf8
h/i5WZEXFqV16gMjwYSfGeNPRnuIdoFRmy2QhpYurF9kVQto1eO92uI5rbVyIw6X
0gIRIFIdTo+uioDjaX9hTU81vtnr3oUZj3EQZ3r8Z91iMpyF7Bv5ob1+m8h69/T8
p1U4KFSZffrUDxroGupL0RJGSEkcjrhJZECdVTz0awN9JEujMkSnl0EAyxBA4NMs
WLWypEzd3FyqBIHuPNMpVxVlVhm6aGmo8ci3k+HEPrFvxAqKpJo/RJ05MlpYh+aO
j8Gshpfph/hSNjxPspBm1bqxLZn3+JohBGaOb4Fo7QJun4oEtHxhC8PyIK8iZLCX
QZ2VcWelvYpw1+4EZ1qzLB6HcHPkBAh1UsUXRWaKn3Pa0gH3KZgo+OzZAk00jd7e
1lTaDSCAaDAjGnj1rtY70P21oj3kKYHp7FIfRpMSY6KvRE1wiAV0LAXk289DU5NZ
b+gisGD8qd7h5nFnJMyS47424GFiUMhfURDau07xt27OtiqfeF4E2oY7ZCUgpKL6
iadznK6qJfId7NlW+1Eg7dvhgaxNjKj19in+P6bjzYTGOnT71GKLR4cInZMZb+3F
bnnBlPZrn/T9HxqkrDdCqa134x5ajrK90T3LVcYJCbj/HfZ4xM6cqxQ6Z8YG0Q8O
d4CHt7vuI0HhUW53lSxvUTatwpMPNe1wI9EJWFtigHBZPIp4gchFBtOvHv2QGbrd
JMbR6ij4JlpGL1FPlMzfkCHceOetB5v2xd0T41HHJibz9C5HaZg/uWoTnWS1Ygwd
5g2hyyIpSXguHwmpjVc/kIUJ4w0iV+tE1H3QsFdGDcC7UpCc2WQMuFeSPTo+YSxT
N9WCDiohxXTwOT+QvpOcYrf6sJ0o4yfv3TKKiJgFKselO3MsA79LJWedNS5gU8+C
L/bsfNKBHZwtbWy2dC9/bO2MLSes1e1gUQq+dZLq+1EFCsYQztP/zMC6SI5bdjcd
Fh/v8T3n+uG9eQxbBnccu0BPNr0ahnsefjtmTytmuMUiZRsY/LlFw18rstwm7T8K
rnnXoXF2mGHAHGDpajhG+ydbUbo5fDrZ1d9Uca67LYQv/MqI7xms239vjpwUfAXW
0h68ObNGayTwYNh10SFiCEVCv3B5mvWl2BcxgXGWt+rKZKV1g2GDVZBrV0NAdVFH
qa/EFTZ8OpiaVgH1Xfo2ypQH7P5KylOHkp7/8n24Mj+HwC5x6ij24lj8ItSonBaS
9wa/QGpLIvKwsVLVyCAsSJsAR1bINqCZWuu0El+WrerSbF9KjAorh+hZnuLbh2bl
+Q6CRW940zF0Gl3wwEyqkE4sOjs6cI1FFcPDzT1YpEQbcw8ECm1vUJ3Awzf2oFK2
7YLlGZoAwlPohCbvt/mBwVRwUnKIheqjtV0ZA306YjQkNpBM4GxhKl305jpaHEYu
ABEthzykVObJBzwy2P6vx9ztp5ERZ02AW8yDSj6X/TlDVXnPufYt+e491v6HA0bs
BBxhLCu0AxkMCuAM12FojMCiLvaNLgwQ8OZxG4nqkB8aFyoNnltAHt7otWyZTV/9
hKtEWXvYcFjDCr5jthlUL8YCszL5/AZNoDvXxQ3DD4PuwYTDeQqYYYBFh4RdbFKW
nAEJTM5RcSwe/9bumCww/S9+zJYDbps1x8gf72bzWpidDK6ln+2WHccc5H3/EH2N
4PssisrXhybw9OzZyRWMx3sMQ3ncMslHYEtH51DCgDk2Qg0OpoU+NkYVU6spq/Rv
0y0euul7Q7Hm5jBoXH4pb/kFq5046rK0aOALKaoAxT4c8QPdL/8NkVWxUu09KRQn
2lwmRRgPPq0fqw5ofLay65nq3nFJkm5/Ims4f5Wb/teKnNIdvvvc7Z/26ofoJxUa
EbVeR774zxs0ry3KzJMmfiLkzuPld1ChlioaDANimY/47cHacQC1OCYwGsY656nY
RAnH1acJ+50grt0fF9DmXJwQDzCzk40or65j8K4orx5C4Swh5NWYJQGS2ugqLRwc
rzsKzvEH67xV1+p5XQGwIAqKyGsBQQwOIAYsOd0E25QQoH3mJgCA/crO6/+4XQBD
022VmMuUkrSE/M65iWdhQf8hGA8HMqZsEe7tRq5vJjojNz+fueUAwkz6ShRCV5L5
Y8Mi9a6r2ir0rpUpyWcMwjg0JBMAbwk+o98tHopmHGkTkUXzj9VOywsimKgl0iWM
Im7cP2AZfbRnBhxb/Msb01fNsglArEoMBlE0oe7gdVXgrDuJzpqBmHG3gTJu3MYN
U0YRjgdPlI25VYUht/DA6WUDBcW0klMMXXDj+rrisorgosjoP2bc1sYwHSdyziHY
1at3+wzS/afKiqB6gLR6QeJF8i0JTd0vcChl0jMG6Y/Fk5xT1pkZYIdsAYdDHNKN
Aj5fOTTQL1hepH1YwjXM0O3MK37dC7mO8SxD1F/cVj0zUr0IU5X1ewCtxaptzi8S
TNlQrgW7CUfo+eCixtSj/rTL5U657c9FEQyIDDXRSSGGHT0KnOCrrZktES7c3QuX
BrDjpRP2Xh9K8DB6mxqUdpivhk9fuOfO03jMW64MVAyrRZuBgtSp8pHRXr2RU36e
nP5prxwKS5NHWqKKjGuMT7MXYSAKQG1/q/KErmx7URAXyJIfY8QnXi7yYg4Jukov
WOEG/LpPIRKcQEmaKBs8DSLIBMSd3CE2rqRcEj+v/Jmlb6W/QMXTQJHCVbJ3v6Pt
12RHfjfeJcGqAI7kUbc4NTcZK3S8ezk2gPUkUc0VWBEmzEaKuFdCsfWBaIv098Vn
gjlbI3p36VKWyBF7zmg41WbQw6JKQid3Zuxn7q0yMJAnscGRoDchh6EPr+oll1ek
1ZT16ahH+R6uGltFDGnvztbmxBvLFvFk16R/xy4NIG3IeMKjREl+M0qTqv0rnAy9
hODbffF395b97LrYnlhItcGU3A+48a59KUUuCF9NT141Tg2+h1WqS4HyH17rUDmg
pS+VRelfSmKwlBHWfehKYMPAgXvPnHsRJ4H6bUb/P+i102aCJ4IugCAL1Z6EX+S4
37mk3nEXaryXpjwuGRWQ4S5RwekSvH1twBN8a/IxNpv+1160ZSt1JQ2ZaUt7C9e4
fJWsGuVNqAbE3Uj/696DIb0LCubjb3z89CulQ9XprmIlP8Davlj9YTcuQlFB9e0z
CbR+OBaE1q8+ZCqHoITTLxGBxgWwPuh5YcWUueOrc++YcizNn86DU4LXHbj5nlrs
KCDGm9qg3QF2hhuon6F1QsQveQjxj8vrSPwhOkURGgz9sPKEsp9yq1fAdJRXej+C
Xo6+64RCquiS7gXrC3Ym+WeYH7uOzqcbBnIcnKWhwE4L3236mcMPNwz5+yu9N5eN
oxv1E5N9eIqszgKg59aIC3iRK2xDvUT7CuTHGtpz7xmj1ElNrC73lOGBdjdyssoS
Z9wFiTSKtu5F07NAB8mLMxkWdOUctRu0+Jt4j2RUi28r52Wo4u8AC6+nsPetYNJm
7wH+oYXTV32mGPe+zYn8eVXmyokDoabuDPOE53ihBCKX2lQ2KGqHwY4L299eIUJ8
I8+6bQIy80G/IGXhBKhkmPiWAQOXoDmsPXG3MRUn9FibwBGj9IPlNM9BQyUSN6F8
FUjhfdP0mzRvUzXQMGfDu5bWfgWTsP1jQbaGteAtiWbHryoAQNY1Yn64SY2W6O/m
I3iojuyTGG/Wpj3OnH/0YtJ5Nay6CGoxNx1RXoPjIte2GsuT4kCT07z5ef120LWr
lXWuKl1LQR/Fg8Np6f1wgFrsRRTWNeymyMxIMj2Cl75i+gBgbrR2mVqMVuDh2UOS
Jqs3C6NVwergupkSSmtYJHRQGdpYphG3+BXIC1a/FZaVqu/+igcl8Bu90ekvafDz
BEA+/UDAxH6aPhLpHDxw+3BrwF9/H3VsYL4cHruvNBa1CaD9LsHauc0ZzniEIRgl
kOo20CrYfaEMPlMnhyokCibag7Ne3oR1d9lJuqmYdef9ShofrChHrm9YV4e1PR/s
kMft3LExVt8zcpu4tDFS5ZVf3jEsElmrvHA1hQKfX5Q0oQ5lRpy0aOlgjywjv6lL
Y1anjM7uQGTu0M6GK3Zq3nT+MnsiGN4shCcizTvMIenq2JevFZG1dhadqipillxz
/qn1s0ClZMcT3MdsC76HQy4+h/I5oIkUfEN37Fktg1K6CvkcoafPRE8W8QurPAiZ
/177xSWpMMLJerzMhugyR3SJkOrTffFW6sakaIhqwfnwuS+/D/36N4mf1jLLxhIe
9OjfZED1ZPDo2/hKfLO38iR5Yy/Fc8KEnRIHXCdO/8iLj9Sy3kkaPDT8hV4cmopL
2+Z29cJX96ACOMP0OK6iYDltH16qe3bJjJAZMWGVhIc18KPNwi2cZQK3YE5XwzMv
MnWCc+R0kSLvd8uyjEj+Fra+8Lyr1HwVuj8SxSSK7pPMcuUPPBFN9EWi+DzWhvyW
Eu7oRjQpZvm3Qc+7KFeVrEd5PfwhCsJjVL4ps/dIWVmOMGVorsMqo1giDeA6dEx7
1vXqVJ//HxPv6dgd6aIEPLLnr4wwHowQ805tdg9rN3852IiUMw9SrEYK54ZvMm3p
Lc29dZuwkG//Ry5fQt0l21XaMIE8hlDaj7GBmvQW5CEqIjuVvw654tNm6L+aD8zz
D3dxXL0UUFDVSefIl4rLdEdEaaxP2xrM9ds23w8KSSX7OOd0Xjv4FMvUybwc2I7T
GdwLh5N6FmmzEYx4n96JlutWRbImBdfp0G4F+nuPcIFLlRO5nwzEaHw1+y/PVfVb
VRZatgllSG0V98fa4dU+AWsmPszC5Z642V5V7Z9/y3SrFgZAONXW2k/PiPrtUA6O
pbriRrOeTP/8FyHxiblEhRG5u0rLnpUcISTo1QZytSN6gPnxYKJ7lS2zDaLEnD7m
Ppe3L79TIZDSsBqWEm8Rg5TrXqUztRlTUZHzqYt/WF9EYS7P/7nYSQrr5rXItw61
QH/2jAngscyyc9TCyeDVbNiQsE7gW2o3Sb5659CBzS5OlsNq75RdDbrCRLtFzfJD
HEXgjf3VBwuffGHgShNDTAYiEL7asGhwYP9cg9gaBCM0dnjTfIF8JxWwiz9bsCQv
78v2OfZDw1Aauz3e3JsuqUT+MhD5xCbwdrR+4SdRkcX4UThUup8xciKe0akRbgYC
T+MgqhjuM+GnRqo0onbM1EE/Puf1GiX4SneFl94225aHLRITgx5mkoS1e7wHfUSq
gOTCF0/3JUw1EpJnFjLy43lyWgbg8PFc9ZCWRRz3be4DSOCKDqdGNVnDhXZwY3TA
F9yywgieQwxauym72IHsGOR/r1EiTba86RIU/PQ2LLoH/4nw4h1ilTBQH/nqt6vZ
8PGFQ6vqDf5UX97oCdoVo+zSeIiF/ou70c6xFbxxqfrrka3MB6mFji4PHRCMXZ/a
tqFhYdVq6FHCi5nuKjC0kYN5Os8khA7llseqQmF3ERpctw6GFK83S7FZmSSMkR3G
DjPl3XlMlUlzzXOwXm3WzaNY92Hv6UmzglnEcZb5YrIgkCzNfIm22G/6PGFfxaXe
9OANCQdtW+rgzYB2OOLF1VGTfBWQ2dhp0jJYeNZUmOcyfKD0MCTaNNf2nabfRDuF
xBjdrQeUAK9bOs4HAyRvYZ3JQUb8Ocb2mVk/IvFrBOPs46KnJwOxpd3WMFw/SgTJ
tbsNwY5pWeRXK/yBGTGsgM1wX16oH4nQkmG1RWzaZFScWo3su+Z1gnvUzLVKVSJN
Bdiwqw3J1lAT5vazH3EaACbmDQAP85lNBxNawj7AqtddnnqnSIYSXVO8KZUtL+Lr
bIkklP6PM/TUx6GL0Do4iteOQU0fD+oHmipe7bcjxuPzlw05DqJksX/WXQpBqSdU
atK+yXHrEiZjrS+y1+fMmhpK8s4Ze2Y7pnsaGxbpVVTGeAsCxnvJNz17cgrgdQQU
68FZjgee0+aiXTs7oUGb89M4NfECNIEKP1/GpKe/VtXPa/4DoJUjCTUcGDu+JMq/
8iZ/GPYX3GfSzZgYArOaZtP3PI5aVYbJ3y93mCUGbxuloZ4baYMIzAZNU3gD3VVC
1azwfV2NHRoap2IhRXCpaZXcjznvzzBUB97uuUbriuhgNDRTGBEkRMTWJjBO0L6y
8e+A1SMKY/v8jS5/IYDs/AbdVlXwOyIcQIwHYb8WjMKQzbzfnO7aaK8ENJMboWxV
67Fk+63Ej7L/GrdwXmiKYzFVuWGfoGmm2r9Xbei6dugMGBSxQGJCu2av/xEak3qR
/jix8ZNa/e67dImZU8cU0g75OTiHySByf+4Mvb19ky4qucCmSJz8srm7L6ChY4yA
KCW1MnvLf6qFQk6h6dKgFObEzOA1kxB6VCOQFLfzEUrWJJOYJIxJ5N1jEFKxUiBC
z0wppHlg3zQt5YVPotifDIoAPNLhTx/yrTSET+DOHHb8JUWksN0KqhVWuW3dEgDS
aD9tWrGIbm8u4sl+XxfomJ58bw/ueQXSO8Y0bGrc4KVZQrIGxIxPXl+35dxfN5xD
haRVPveKYORk7nCOwkc4xutXNnb2opGd+T/KcgKjK2fciby+ifWhKEWkCnzIkI5y
XfpdZ148jMqPw2GoBkrYeCFdOEznob1JEGSVHhOj2mkusiagAvveiELj0XOmCe+j
vPYL5wOOVypwTIUI74kb8Tl/z2Q61Y9Ffh/AQv/pkFSau785KV6Xe5ybEz5uc5x1
ZcQ20/jlpu0+Yr+axbBbZCl6FcYxZYXlY1ha6eiuA2RO9uzPTaj8lY+WN5fTp2SU
sl1t4O24QMO1jWZ3X1Lzx1axduIo6ewN+ZzE3GDR5Akz5wD41sQCsGI85aE1wKwx
/EmHX2tZkjcvbxZtGwNAoVhzawFQuLsKkH/sYiLQf3B9j+HZjnn4S316sg5VMRjA
zguU8QALFLjbw/Yelh3wh/IlIkhkfuyYL8FYdgkrELj+J1bWtrE5bDFcB7WrJFB0
SiiLOhsCc/PR25g+R/uHqvJPuSRtwKBLN2pcz9rX4ikfzTgvO2sVaj7ydZVDB82r
sLiYwmgC5y9+ZvCeDmC4unmGW6xiopbA2YUr0FkFQHD13EPyImBq5C4D7TQqQuSc
JmzZV5Pj7Ls5ealW5H8+OT4qVN5TRr/t5/1eerxadXaOalV/82zhRagYbGEApuc7
LwTQNe/y9ZO23X9d2I26LQ6f3BLQ0cqvfxkOMPgQAkxmQufBtn/MsZ/98XGx3K0y
z1oG2NdgVShFwnpBBe8Q/eoVYbfBn0Hp4MspL84CceMh/D1zFM9L4rJq2nuhtUq1
gNexA3s3Ud/4zGUoyflQ9r/sT8llUbflMqeoNmMIFxwr/sip7TDlM2CLf67Hf7Vi
/bxEuV4DlDQ37Utp69CEewotzV+bxzDueif0IKvYhRlh8st7wzVTG70k9qr2BewS
lihu/1pzztW9NNaLVNocB8e1Ybulj2mk3NhLjrdypPL3HmAxJSSWE+6E8XvzzhoX
EwuYsDj6WG7KTLYjmvIdsTKPak85wcjrsaGMxmF+BgEBTyEW/gmTC6RQX60WEdC/
3viWDbN6R5/YJq7HtQXtlzHBa+RRgibLJSYSiowDHp7Kwv60AsxDJJOLGA0/ZxtH
nBzKFQUqBc2CYLfkhY2CeFmVMG+nOsX2+gH0Bc80VY3EU7/FyndRQDcjncSQoffK
GqIBrqlJoOkxbGFQ1vl9r9jciSJD8yz+KTfBb24rTYgTQSjnmD3EPxX/HmESQBYx
ixA9pvmIlxyMyjPQ6oSyqVFW6Gy1WRLW9q6zx+OKAwqTLJhaJkN2XCzspe6sZ5SA
su7gRsiZNw2mvUTA8DPDgo/klhxp2P8wTBwO7sDQhGAu3yyBdIp3ResymTG1rSIR
cnqZbnWIrYLWb0Fg7nRhU7OS9G6du+i0Nzxq1vFH/J9po3ur9pbInbgW0Q4tJy/V
/FO4yiLTojZI1U8zCAsApA66yXoNVtpKMCOMfRRKgegZx5huKNfF2X5bFb0G+NSA
2WyzyR3fAEwZGBjBi3RR/ybsIWeKG6x8SH13TLX+t9x2O2XPTrJwwZlsGQAC85rE
nGI8WZhvZWBcgbtlASWbXg9jfQ8xnsGiXAgO5kz13DMItaLywTmfKrMs+liODJei
5oDr5f3a9svAXAvbW4S2r39vJA3s0Xb/gc+yPjvjAkA/FahSfsH7UAfVHx/fuklP
5iftyyPZ/HCX/xnxZSQqzVHX8g4z+GXAuCh5SRlo23EhP/MEOLi2l+aS5AUdf9r2
UQQxPwiR6W3+ZIUSLyKpPK+9bGL1CZv5BIBlu8WHwUTQcCeryTTCWqh0IqKaiiWD
dvjTqb/4gkzWmFmLh1XlyWjuTdgGCGAMFh9GHXN5F8LfHVAR4Ey4JKgm94hj+Tgv
c6TqjwN1OkjxYQyB6EU3kW0BILnyUZ++7C2i9EZL7BMdqZ9WkvZXKLcmhjjcX8LB
2cZ9Yoh3rNh/7JoyGqWX/6P4+ZxBwW7Ga2KMSLp2D3yASH/pSPuHiIODbhotYJQ5
WH+tBKZdWVjJ7Tx4VVuMhs+3TpXcab6mtNO7O9YujyfmcOfd51aVYuQhQc9+F3di
aMoOnglghSDJ+Z4vUXFQuYRObkC5cTv10s+cr9CtGwAfxf0hJC/0lR4HRpmfv5V1
YtoL58yHbAYmjIDWOPexou+0i1ECkd6eDCZ1A9Z/uCr05sYH9NcvfK7WiwdwduDk
2DZXro4BfyTHEUQiU9VtUFwfHls9vqa7AdYou1zNbQOhuVDX2ZEl5XuQ2U90O9r9
2iCkXGrC+Ql8vK3mIHuj0BbEJhn3Jqb1ZkJZvVbAvJESO1jnkquMT4b0F/yxMBOC
E2uf76H9W5k+NlxDwaJdQm74lsWoPDnssQ60z67pYX9Vn3iJJqVl9daB9Imt4mbv
qx/i3dIVIDUh+Df1IyjA0dlAtn3TMLXYs36O+ONGsDwh9t6LVGFQS1nYQM8cWsAf
BEg+3TBhQzciJy0Hl1knFUnCwiRYDpqhvP2+KwxUds+FSR0zVU9XjoJSHYLJdjIv
gYGNtmsjZz8XskHGFPqmbOcmzQjEpIQP46nvAITt5Mtf9vgXFPsDJCWnOdO3s/Pd
bi1HPOuBTemqigrw4dVuh3fjK5mEA2zll0ydyRR242SLIcZ2hPzMwuHW/Sd5GgKb
6sQYpwlBkW2h+aZN2178X3JkE6LTCzkxZ/ZomwR11+hJz+0Ql0Vr78p/nfDgku1B
2saRC1hRV6xloP+9rjzAXtlcWSpgIJW3AzS0x5DoJJ3MlU220ywVoYUu03IshXFT
KEnY3eftyauWsmRIl2TAuWxtyUGgPGz3zKa7agFI9HLPPl/VV81NqZdF6umYA1Av
BakwTwCn533jSDjqERwH/EO/JI0OeGN7rRWEG8HwZ6ZwwAbsuV67JlhqV5886Lgm
80peZ2zy7HuFTuLsuhWhY7inVQ302LOwg/JbwfhORIJpFRbRdXn0pmzU9C0mfoHC
pRFturG03XNSz3wGiLKWBcuuCKAOJmKQMKkYHNaxfF9Xdeu7j4kwr2fv0MdxCm5y
qghqSmHYSsscUQgHwVVLjZPNWn0ak5ubhdPBnJLxOgMEor2Rv+QZV73VUZ2KaCl1
PGA7tzDCH+3ElYF3UKLCtQ3aDLUoHc/JeKN0rsUZhsSQH5G2fDlcndLgpTyL0qPv
Rdqj9LYsiZTypSij9r+ZA+X4/5o5musiXSpMKJclp472+fB8yaVsC2e0giHOFwUw
z5aMnVRo0FEJUbbnZbPeCG1cYztbC6fPy2s6H6Ve/hLVzgFfeE56EM0mycdpMx31
aJ5b7Y1f1XurNe+Bq8+nDHMX5RN+6aptxBNA/4GiV+gBhv4Nc3MDJ4XFdZ1vfGRt
svwJTH6IWPwXyUAY10q7iVexh3+uYKOopQjYzYcV2OLjtMO3/h8jRM6orzo7rQIc
sSmBIMAk1dmar4SGcVtHOFCjcYcWHNcrNpR9EPe/+gSbgS3agM1+UlXg4UGZJBK5
uc1Fd2TAD81kkAKUlQyQavHL7ESb0X/zpomohilg/mDtzLD6nJ8fzFr1NNOgC3Yn
zr92rQ5qrG7JYProvi9wh3+AnhQsHLnZF//QSIEMYbXIfbe4Mhdr/XnUc9BrWURq
RTfdF62vGA0ZnmH7kUze8HtiwBBQ989SVl+RXVNk1DZwiEvfN0FtgNqExmoKfY90
DOrN+aADJTpLhDn8FLQstMxhkHs++zLYl7rNrMmDBlt4GGLUPesQ3oBHIXkO8YSy
CpIeSMxzopzvAOsqD34RGykCobiTLZ+Qd54Z4v6FPgfA/Y7OkY8Zuh+fZUrXYQM/
yAPo3q9/iokStsqrt1Yjwv0mT1zqwz5dDQ6jPATNM5mfNMOXDqDKpbLzDhG5ycZ8
JICGMf0SHDOnadLzQ0Q++jlt+uJgdhii5Dto4IGiXWoa2bGvxpOCJaN9X3Exu8Bb
d8+PcGP5JzGRSROcRjXBF2je9hLeVuUx+woQpuPVXGSBXw3kPmiSP+N+XYCFXgV3
zxCUhdjijttP7hoItTmG+uX6pqpK6jl/xF7rViRu5eeTtMbgMzi9q47p+PthGIrm
9jmyfp2VvZIm9IgexOqgOX6CmY0tZegESB17w5j6PQA/zBph1gVhWi8fa72tzCP9
H/hsQ1QYGESsSIYwWz+Q1FjDaZlueJlMwvmNKLqAS7zQ4Y6T3f5nQtKryLHBPQjt
A4aY3UWCyGbKCDR2sgVk3ZXVWJR1qkIlZ3afCHgkaoeiyj75SPQ1xaIdYvGB09zn
VhbdRSm48/rsB/Ie6Cu3c014pu+OUrdUbjHhh9mhwibK7TGL/3d1h6s3s55Lf8zt
19z1Oi6xsb5hfXkk3xOgpjgM73h8vHRE4DoEOMdYd0hkOAzColOQ+3eNeKg2ymfj
zVt5yA7VPDhN2syJexO43EBxZakibreJqWqR3GRn2SFzbxdVzRx1HF+gvwKvuPNw
odFAHRimx7e5NT2dvJp+9p+SHto4uwcnL2PRpg0AktW3zeqNaqKkiTt30J9t5K/W
KFmunw+4CjXFtRsTWLkN5XW2GQKCqWxB6FHFWQZx1hf4RmZSiQIa9qKmVyeznc2N
bXm7vVpO/aDqSeW+amnZRe6040WM1Y75NYcHsHGXvX2VZFGSXHX3k1pailMZ5mNi
mZgf/g97NbBN0XaWxdG313GXOIpnJRpzdOqNkWoDa3jU2I409ThsKzKth4p63QYS
7jdjpb9gf1UoedMACjy2zF56RTJLHG2mRAi8c8w2LbOS7I1rNOuEWUnJa9szHU/h
KHdS96Ht1eHW8/p1TGsb6z7sp5WvzMWSB9oj/BelvmCwxmHvdZ1+7+QBTa07JgtW
6CNEpcR8Jan+9jsWknJz09lEGKQtipAxXqLKpv2NRlu92+CO6UabjkCaXxurTQEj
QnBAoWC7O/3ZeTiebNLRgqdLDJFin1W0bw5bN9yC8e7WnlZafhO2CYXivbWvYaZw
PF7ez04DvEkkYkrOP+m1yFLZ99WcIUMHHnmLKvGKG3RADmnyLLTfHMFV4OW4c9Tf
RQ/+nPMGyKV04ZJRGpiUqzw8mZ1yVaOcqRoXmEQRYyoHqsnUrLY8iz55OWCMAa3Y
B/kaCjI4md4a6kJ9VgpbvOV3QfZdzqbdF4wd5aea6n5WUSO06VG7MWrK6NwXzkK8
pQeVPOQv/YxfKWv65UhuApwCtrbpU+79m8CznU6rR2DsZoFPkuIEQpDmZNOjU6IS
RuJnQ7LHnKWC2/rp2vFVuin4ymkS/+mQGYhW+8DpkTwHxtD+g76K2VuIktu8iedK
3CQTSIsCyRxpZEn6OMgpFIUHKcit/k5hynnQ5oe/0SAgsnpzSMuegiQKW23id7KB
RAZ1xRbCnBes4CwJdAyk30aMzOqtPTQmo3gSfUiqYm5rhdCjEoAlNb4b64yGwC5V
6R8xGdngtYNp/Hfw0kStx54iroAKH7hgODvuRZUlMv65UFCUsC6LnQu+izLGdj24
MazhXh1aWzaTFVvaK2pHQ1hU0UXnTwPMVJgdIGAObwc7TAqr4SO7FfbRoCnhSUsQ
QPV5QywsJ5nP8nopBY0NNYhFy2yNLet3XcMP/ioTZxwqvAnlOAFUp0NeixJVTSey
yW7t+mBMGTqd785jC1rXXnkZAV6W8vCcGuwXJee6ZBRI+U60yAt3f/UZvU98CUCY
lgsDRqz8fMpo7dmsplKtQQbpagsdgrOp+LjKZETfcjt4greV2C+PVG/DH6dt3JMU
/oG+YSwzc0Dd0PHWye2tDivhi1e1MKEiJqzoWvT1gmOh/cYxe2lcQAyBb51o87+A
CO4VR/hAn+JoEAcx1JLy0/CL0b71eRCKfzNWssPtyeNdVyHl5WoFMbdYSX4/lh1D
bZ1heHBVvTxi+GCRI9nzUpYsN92uDqr+RCTNdA+zJtOqCvl9mJ2M8vKqxKF/da9v
sAmDB3K9m9KAcwYHwh6NtVDR1C6TpFI9SGlsQM40RLjLtWA0iig8TNEWvg9pIKAb
uheDy5fQzVDc1Ob1DlheV1RWsaGKpCrb60jpdfQZDk3RxWlVZ0ye51MHhmpivVGm
eRbvHu+NkGg3BIFst9Ifvk22pLegp/WjadZ1LaNZJh4rSjMwdXRhIXJ1/PDbg+zt
Zjjd+2WGamQRGQal+5IRUwwjkTed1K6MJwMQkk8q6ydTKkUGoDtLN/0pKwPFq1mg
uKcixVwZCpotXJqRshzXov9GdxvwXq4Tock40iIET7408EZU4hVlH1lfqI4f4A0n
E0YyhaWW0t8dvycy9psXZjUYwzrQRelvXOM00f6zlL/hUT3x0vYSbMIltfWiYuJH
DcDnXS7pU3QaxuhxUMtlvLF9ftWq5sGQjR35BGpdn3lsL/xI/lLNxaqz4+ngJzmR
bT6REmoG1GD+dkyc5Ckoj/ZvNGcpGvum5p4yOADO3pHbZ9aVehbDCtIbpy54JBRm
N0v2fBOatx80zkYibAvNUWm+e9NBqC+LHmXLl4SNh7hTqjC88aHRnzAR6rmQcZ8O
9xvC9fA59xdaNyiphVh+Dnoy5T4HdB+2nhKU+dMvSKHiVozDZ6krhqShTdk0bxmf
Epx2wtg3DWpM2xtTUd6jwtCUpcK6A4/CvlRHWaeMmUY4SEixe3vEjFt+G8TLQKkw
TXLa8iXHGwZBGE+CnaMY2cdxWhkouZBrDr86WDp26VaaTKP1AxNR6m3m4uCdPajd
tmZfJtpUx7Qh54vlCJ7h3Nxg6H54Q+UKvlwPpt/LLVjIgLQiIh/c4SmtAGmMMazj
RwqNXj5N+xc7+5ibDnrfkqesKCUsNK4OdWJXbXkLL4xL7Y1Oi+N0BMGddiOS672m
PGmdF5it6ACRkEBeV5iPvUVrV/VmQBwpOm2DLJo+ZYsk1WZDKv8KzYKX22sp3Jj3
62B60lgQ81JWEZ76aAe8jqOY/4xcMxkP4SC1sKzvldYzKmEGabAnYEEjMfC1hwnG
lefxMyjXbSHKQZ84fWMvE7NcpkQxC3tYIcQra466osCF+qVntcVskBjrL2yEfB65
DuJ1NieVxTl2N0ZhfA6yRh/vg9b+oQAx46nTcedw1DFrLvwBwIxHd+y7NwaPG5Ko
emV83SsLv3P8D7yWrtVZRXKaVRsh24Q9QqswRAyAAkaD2kbFDYQ0WFVM8Bhi3+IN
j5l2Y6ZXA/aVczENSischbA0RbYXFDcNy6fCCXJzKHWNUqDcrNeM3wtv0PLrsSIf
Osm52Mt2+Tlym2TG/ne6IcrMUcWHfyfd0i3aX9v6y5xKcs17Jf2idtRtfRtYErzy
qBhqtonxf2Sog8zIt9d5Yh1bs1pF0tESmQXmLkvunbWwcmNj4BYCCmVdZAzWDUYL
bdS45Z0CiNFom/aamjtHcrKhal9T04LxUGd1tnGshpJoYF3lWCzO38NcMkRXay2H
NDu/uqsEzn921V3bq+eDzo0904nNCYWa9vFhqq6FttwmE6CBYSYszZLZ+zFfm5mO
uOB8EXad8GBw1R5+21zgZa3/1IzFKlAVMikYog8nE6Od5r3d22DtSwPqbUNBGkQ0
AzOwGXtQh8blV+KK8eBtcTfnXU/NSg5P6EShqT5laD77d42WgloZU6e30cKi7WBh
ZSn4MH0tOSgFRbjBuM+EN2O7JQCVl460nl3Tym248SPCDRpgy9TTzfFT8X62cRok
HQcvMtYxju+7JnroVuW10XxnXNSsH+mkX4fP3gMhbjM+fqOTFr3zdhdvkgIgtNyq
V3jwKhlUb2kYrclUjdjL5rTSUXAc3+z5rWyzIUEHixv9z8CJxzQB5PP3fxAf/3Ee
63bCpyHRFD442l9rAXSfBsbflnqKZHcTkbiJ0RddB2LCuMFylhZGP2idANTV/8AY
NdoQX67TStfdHhUC+PcxNiYwUZ4VPf1yFmf6JoJ/fsxPZ0OyRFNx2+xFp5jtKEWI
WfO+zNQjuwDW0StnOOOk+tucotBbU29bkhyWYAXo4LY4N9p4iWVn552edIWhict8
ZLYxX2/mlhrHUuOcFkrSbNhpkH7HlpkkN4W5Tk2sqgzzaTenDR1bB8BBnpkKjf9u
YTgURAE1E91dnbaZKrNnbQjVg3cur+2pszbuPYN6QYUkjhMPp1Kpz+6W/rfvM/Bz
wSL9aMtV2rHHwk80/3sRWXhYGE6NXYIqrSYKwaXVLVBbzdv4SEtJbXkUh7+hxKe6
8hg/fMSKU7CKFj2d0Q8OOe0sZ81rWjmSulpHGJ0xw3HVvO33F8g8fuRoHfh8s5G5
VLI4hR6RXZOJXShhppO4l9mBo8bbYu4t7UHo+kL7g6QgYeVFPz6jUdx+gW3R/Lf/
4+Vv1cJMnuMNsD98NBl6CxHsZfRl0qtrz5pA/WoPnhbsRk8PCe8oBTeeewjGdDlA
/Vam5uwEKdBRMQAsiyhu88duU1oSl4hfTM/xNulj6Wg7PTT3Tqoo0liLAPRv60Eh
+D/BkOShZCwmo8KrLF7e5lv87/VB6UInM8c7aeDqvsgq2XB89dtz3901aT1n0Q1H
tj7PPMWn+2SwD0WSfrGhFO1t81kxNB09CxTsxVi9ykAjRMwPbYBKGQwEprnxQx6A
EKb1zYUhS2mqggjJTD4wvxrC/zgMxmr+P8jxDUMxfgHSb5na7urMreKIDcqCPIJY
yC7LeGqsChcFFbUZ2ETNhAJ/jibLgmLnzpY0wjMJy6O4QHN0vgojp0bH94W4CQX+
eIjv1Ozc5iyGOOBroBc4P2DYxE3WpbDt7wA2FovAwStn7MPl93EYDfPrmH2Jg4Cc
M5K9en9fnBfo5nZqx3Le5+5OnAxa4h3nk6czbuHWB1ZpuZIoEhdbVjmEwaDSKG7E
Wazq9n2NIiXZblzUEsUJz9vUj0S/JmZy6jIvsBxnoD4YkkHa076nLweIwdrV8Stg
zMCb7b65kH4tvWAeNuUvt6i51jc0VJxDBgWNrkYR7F8KWOdezIQEyWHfnYxgyAC6
D8zuInDUGavOjrjkYclA6rTVfHd+jEALlW3Icz2Uw2eE6gmxdZNSGDBUDXiRfZid
2GiMIVdzHfVwo85h2wk6cq61X20k+UqdoQ1XYS7qK9lZaiOlxqRADT7bYsPm5xvw
feQ8zM4aGctdF3/GcyZDvzw1oEQx+zSIiZ4l9tdlqZNmF7JQnSjr1rE1SqbQ4CUf
K22LZK4telTxCG3vMnqWm9H5q/bH8YXKisiRxQMCxzXqhyZlQ67wloVyp0p1qrjN
eIrM4v9Sx4khK3vS5Al69R15aoE5gOqkzC69A+p3YfjgpILJThQ7JjHrXM/35frb
QNSfiwD3OHNSa75JGTJDmg/8gUfsNIcIyW2RMsWVTBDLgUKzNRKPP4fLRdqAR+yZ
M55ZvOescBsPLR29a9p/XP92ijb6U0BJt/GVVpwkAqsfrTNd4vvG5BtNwCCOQkxt
tebn/O/geRbvlCT03HqjGH0ZCb6zWk6baVQ8wIu/XG8oWe8kzqotTHYIf6b75HAc
Wrx5pehpF3EF5FMQlLHkSyr3WrAViXZWGuyOCA2XcIlv/y78i9M8+sfJNnN429op
m9qml/rqjiCJO427+XRtjaxPO712h+yct+6rVzovvMtsCo9L4cvBwPzI/QZEeasz
S0yYSbtlFn0OLB3yshl9z1Bf1uETdiGXFMgwURAPkFDh3lZrY9rUhodCkWX76Bpa
f9g139nQPmFC3xJJ8F/uZ1RxgtfVw2cC0Lfdji/K9xBFVYkWmE5rPb7GBSfDXYXk
XuVszfouuv8UrJZtEfXEl1Ydf9LbRE5wDhFvhIyPlwus/bFGTcZSbfX+nlMBxd4m
VOHKAB99dm15Wfi9AiXyt5tzMn9J+f52O45YmLfLKBUDw/aEN4Qh/QzIDsXyLaSd
kZlRh8OVqvp3HN2+EmddSdCjKGJniIEcOv93Mtr2MrRmlEDjz16KovEOqgvANJ3z
zBlqS07TDa1BLINiLlk/2bEC0GhP1Wkvb9ZtTJ1Uxh4mkt3s7E1vdJFwvHrd4xEY
Ce02Xow7dE119Cnkc0pyZYyE8KoJw4VZtx11P7FaEiESxXjQrHbzi+DmuoB/FW6X
Syg3Se8dBLsKVDg2TB27PbbWgTki4vGyusp9U7yzFxyNJubfzVPMatwoqMmdD4W6
EASBQ9xMm2XXr9tGfE3ielC/cXJX4V5v0fWzGJEvRg+hM58bQoErnivFXC0qhZTt
fy0VOC7hgmcO3MpwNpInZxYNNIDDxhi5O4ofRQV9eoavvdDh17W7HJ1JkywVa6lr
DaiO8j3wadfkuPIg44thC0VMi2agpBPDlp9pZV3GTJjEbAtMOMrFPH1dTOElWV/7
aMlowu+eIdfNp2SxpdrbOSwyd4ylWScWjP2qpzdFLzYWWqJ6mAVdv0Sz63csLMaH
wb6Q/OCZpbHcpZW8HXjZMoEsT3/fDMGaD/9pQ4f1gSh4bUOpSH2lhjDQVW7x7T5T
U0Ib+vvffaScsJlqxXoHKeToVtlwr+OMlYVGUAQhfgh6aGldC+kNoKw7XYnLJebe
3jamrkP5UTD/k53RGxVlnm7BeajfOI4SmEFhv5kFAs1z8P7Zn4pVPQwP04I+/OQj
7y1h03VyJVMT8Hqr0D5J4GKYKyrwGzUcazQpKac2cAFr457FHuBjPiuoc2df3RcY
2vIzrMApe/XXMMFAnqoablNTKX18Z0RyV6LV2uP8TRRchbvxxpK8TeEuOGCog4Zm
huBhTh7PBvdGIntwnXEWB3S+yUty6/agTlFrRUt/rZco5Ze4vat6Jo9l3Z2ZGu4S
JTadwpMi4BVUyjpeQst2fTcHbwOBqLAVE0dmx+we6Q8gqv4wUyO3sT4CkI7NyysE
euk3y0OQWfelRjTXUXFI0miA98cbXP8v0GB64qc/LhuZwrbHlKmesHO2Xi6bs1yz
YV246Ui+KcKtU6IuAsjMGa3pGRBsElsRDdbsYNmYafZsOXfX06UV2tmivKd8yrcX
aFJYGiCXDysUoPDYkJ1/bCqcLAwZZ66HartlupOhmH/308S6IDPW/YE8MXm+n7a4
QO/HC8IJZW9nabx/tTLyJ2G4423lPbgl+/urqMwRYmQZY3x+P/+H+Xc5pgDGwk5N
OSjG3G+u9stJ08PiaFVrJw9o2Nb0+FoqGVFBrWrcJ1qrgdjMtvCOH/UAiWqShegn
22IupxMPJPpAMGcH168bxAtmTg4x8QL1jb4Ib8ItF7wMs2pUPoh4PoI9OJqig7mS
RyAnd7cZceJD3sPHPp4KbaazHY/uklAfkLBw8BxDGsJ4FswBI66PdsHydwLIpbfR
uZCVyicPdsNlJQR7086SqkkYGWmKAx74PStU/nbzxlFz8BhH8LPajsm3x1lgF3qp
iIfOmL4YBRTwmTURM1fcVMNi5EV+QiA0wsmx8H4dsG/FOO/du/h2jOwzPjTs01K6
pi9OIc5gNsc6EetN+YaQJOqVfKp+BoIODYgiooyvrDoLPaeprn1Bf96vRCFCxY2Z
6E8AgIzMV/EVAhJ/I+RZi0YrKe5gqMEX7qFbJL31bCmTIenPqCeiCWdK85YVoYlh
cSRDl8A2MJLF22EBLbyNLQxHbHPdgS+t5mOTg/Quu8TxxltmBgg9fyNRBJZIvuds
ku9ThA+sTJc9AhD0x7Bl352xFxd/SOwazaYdFR4CuoB5cB9ywd5UZI3pDL4spphi
EBe4bddjI5rCbMjYXOU2q2gjeHPpsRD4PYSRI+eVZ1mImvkJzWq332IG6d9uWDl6
BFhdEIsrrEaATHFSdF+att8DD2JX8fJtHPmmnLlymBWsucc4EKEJkHi15lesrEoQ
uhHzkl0e+MiDGfBvZuQXUDQnGwQ0Ac0jPfEXAxtfavBIzIs/dKUfBp50idnL69Q6
uYAG3ihXMbZHFQWxVondmvyTTso1emGzAZhSHG01R23MIIx4dKzP+OU9+BWQqzxg
TXhFWEijA3xPhwlozVPgSzs9yGBoc0zatrBswyALRBEYBap2/P5T+QPv8i5tknF7
/++jgda4bhQOazruHhIw2UVHjAs/zZQ1D2hPx/eLdjJ0DRn8icIJ16lHkpiYeiM5
E109CeTop+543aY2jZHDQDJpTx7VW41ZasEEFkmxZ90K6dEzwRaSVZbz1l8ZJVC4
ezraLrWpU034bpJMVY6I9pNk39FQzxRO9hGI/W2vh0jzMGPBTHWt2tOaTjL22XCG
8EkK7rSBB6cH07lO+RMPcDHYD50Ay/EauiTnA9CkJGnZJs5WVXj3rZ24LSxeZ0UQ
eEh0gLkL8wHXCYWGHnb/HqFey/q1x1fhV6iLpGJzTTi49DmOSfwGE7kGFsrD9VJ6
bMj+40eHoZ8RdrHA8CiYgAHZRHKDBXvc2uEET3ZxbeJCYHiNYOFywNjWQsG/+etg
Iapk/l99iuXcU15yi+CwitgULKRVRHoddtciCNCv5hcBIn2Yoq+hoyh70I05ka9Z
6iWsUlXfA7KTxG5hLUBR8tRK9kPyDfdUJEbHr7pNAIto6HwwUjxUrpRppN6V6Asq
MUfwYeWp+A6lolvstX04VWbI7dy+Q9TfKCpp8+zR7uJdLtI+ZcrRYihOwS4WyMnp
3qjTcSgNmuq7sbZudcthrwGmbs72mxHakkvuBRjqIFGxafVhsPPI2VLLr6FHggtJ
71Meo3/0IfqfmvXEjY41dBKBuRX4nKJV7bo45rRMRvLHj4xDgbfSbKwM9DjFY5K6
KSlXzHeYzj/CxRcnrG95EOATXJL/EWxmyr+VeaE4lm/YQhMrZBWqAeIMZvdjtO3p
24gDPTvgHt6vH+2FTpoEfq3b8N+xLRoSyrXcrHBqvrM1UfWVHLLMzIN8ZQlNt05j
tWHHQYpxZNyssI61OCW1/kdHGxmhOLJ6DKcT+RM9cpmN9dsCz3Ur319fW3pJMwn1
ormbHT4EFoLoHeeG3L86D2xbj9vlq/6vlRdKyhRxi+pje6Jn2GjktaKXqrSuWHdN
Tp2sbRjpShmdn1sJznrHaucykngCXhsLyLjY+tb3jvEsbKCyVLowW6dGx+eQ6pES
4SG1YMkoVLCq+7bk/VrJVb283amtpUBIhl7xLIUwI/uB05fFUwm8jyVJtpyynCjw
whZY+tR8ZTdTWgxvKHn30/T8cBbvIWAQYVPinSlfADVNgx1PdUVUMWm4jL1Bo8f4
DFR59ez3K8ZAUSfU1kzZXv0LflR03S1jSyE0PibQeiyelvHaI4gwQelWV0fP0RqA
P0AWkM+CdvLZBBA9n+39CWc4uuDg3qlJ1cwFamgGxeIMRC2wEX8OTJWtN0gNiRG1
FDuTLIuHy/y4/Utmqt2ArtBQMyPZUeB7EUHetidPkwtGA3fqfWZEeIvGuArhlU1G
o1ZKhAwKEFT9lBa6K7NrT1+XVg36awLeAtYfAeScf/S9NkM+ZRMCtoZFQe0nB4Aq
btOvBmGl43TJTNhdh8cvLlmnDWQYnhpE25wj28d837wYgze2ajAi3gFVcCpDgdNG
SPbLrSi9Hgr12Ev1zGUIItTTP7oiFx2/QB7HX8ORFnm0vNhQdgCWnl6M22XOirdn
uQkUJQ9On0JxyLVgrEieqW/FL53g4eLylEQcsleeKcrL7WA+VWLI5m4hZRiJrKTP
+80rs3a0dH2FIFcow1ViE5fRyqipzAWp+Aoai8GH5WjsmUR1Ux3YFJiyV0cSGIM2
nUvZt1esK8XFQJsJeQXDKRQjd+ntSDmcL/9vygUaJm1EXQiztIpHz+GlcAQmB9EC
WOFpkOuS9K1SUyyTo9ACL72gDJp/XAZSMiCBjzEMEkTutRUT2v0LksBEI6zdPOpW
09xt2xF2rnK9WY+cjs6zGoqejwh2jMcOveSU4/AmRwZUiEO2lUSC9uZNKOcQuTd9
ErwhhiBtvWCzHY+CcPe1Q2NtlT2EAFG/Yqmqcq/NybAUuo5cN7hsvFtqIUao3Ss+
k8i1XadcQseZ+Kt6uxm+d1rOOaYTuenC7WDYvIvlmsOwiG4EpBSW0nrfrhgQRmVo
1AvDrsW000td8N7PZ6j3ovDxlTBKu6ona8IY6Uq1HC4cLKOva4GQOU6T1wECtHKM
iNICpF5yAYQ+oQCqXfpzTbb/3P33SX3cUwvRNbHMIN9bT8gM4ZgA+etBrQUkkBO0
bZQXBGRUxVp/sP+SnXz8Q2R9cztmCmvrUdRM3DKJXJRc2liTVjfqtWENmox7AlE9
4GfsuprOvY1/4Rz8Ep5lMoc5qT0X5+pM2gVwqpXKhG8SlEDERAUAiKWRELhk7Ggs
gUiEpR7KDeEkUd1BrOfowrsvfe+IS9o81hPVAcxCWq89Hqd74xofuA3RZTtQklZJ
3xyVYUwIBdDUjjg5uHxo4MeGvrhEdJ0s5blD7VWcrGwoCbQ4kDEnokdrOUJbXqDI
LJFoYzTZ83ZM/RWXP4NYnH9GHVTwVbGWt0ac50C5gRzv9PfZZl9r71aNw5sIYE9x
cth/zhoX58CMOQAU2BLFqnWP5DomYDhScDOvAtS+bvW3jq8QYxwkDHa5FuFAunlW
HqaSwmMPGrvnveSLrAXR4Q1w4Mif+VpBqbBm+z4zt1mPyaF+R28LV4PJPXN/qoi0
qprTcQEZzRi75HMa3rUKGX6XXB5nELuIYggHYveft4KSui2Ie6U2j+kEfPE53d7A
qCz7SUHmtPeWBwD3wdauJ5z2EbfxuwpKOCjTERpoMI7CPWfi+h/HPuvDPxGBGAS1
XRuUa+Umdhmn78gqC1OQJxSXcAs4mh3OGHOVCkVZLpwItGgr4ACM95hCvl/X6pYV
r81y38xmwqBQB5V2xmJXJ0H4xmbTeTcylEnDzrlIaKDTUbmORScYnNZh7RQjcSSS
6g9FqC5aKGb5uOI5BC5rCddEOxDFw5ZBiKIRLlpu0g5bqkEwsnqGeD1Ul6iP71fc
vYwjWUkWi6IyQf0FKIHmXiDA+Al5ckH6oZWbSKPYFnk8SdPKPz4tjoPEm5ciVw2X
ZhoW0Ij8bjzmnU8ESVPNe73dnAP1MuzU4nRk2i0Ph76OkmaEXRvXMrzoZMUlsBJ2
IPjYEYOOiza+NG3wSmdu/S0YV7TrMOIxuZqxhA4yW+r9tJSNrFaAKCplp7gMqizn
C5GhRz93j6IFb+tqvtbet1CPoKd84TOoGCFcop8+TQPrnLx66KI7uKkCr1MIO9pi
7QJ5z9JpFiFdg1yJqcrZua9638JHy4tpALjbdG+7+Uju/CBFbsS2TC5tO6fXp90A
u22dnOg6rsyKGKTB6K8ym1fRBLFYEsZ1OpQJQz0B0UZxQRUtmCz7xtzUWr1StbRy
wHL5pA2GXAO6YmMb2e1tp11GjmGI9Akm+ouUqp310N+qdaLmA2eqdA3F40tTUiLE
eFNcC5R+dmy4fulxS9U6kJRYIF+tX61Pe1x35pPtX55eQf5rlcjwhLyfqs+QPJ0s
1Fwi7q4UMwXjeWMkr1yGa9+BAwaPGKDWlHhikvHrrMMRyEpik5vv3v+yTZDHnYh5
Ej9dhBqlRJQNiqQpLOgc6YKxSXDy96H3LhUeciy+1pgyyEYkW0ci14urChz5zR00
cHFd5vhQqdZwQu+bBeLwgf4fUyHpLJW7e7r4F/683H54AGnfg1eL3WmVHNL5MqfS
6yVFc3z2GmuKXRbTXgWUL8GpLOMkC0xplg9VLZLbO1x8xzQMjmybTMeFyArFGyQM
frJrSalzOX2RThnpuceryPK6isonmWtD6iIaabgMXw4SfKIuyic+8GXLhAcqdTKJ
aE9vqGxHY3k+SIPoWHC18FE9kwYCVdnmWydvuFMwhOEQFS9cDNFdXmZRQlmzhD5a
mI8pdX7uf8Z70gX88fXspDbSXA+O7Wwjj9MTGFBC9fZPpKpfqXdj9ph8BkKhaeH+
/4HxF1A1BiaJepxpum71MsdH9XrfdFs04ZGS0i07cnCDBPAszpNRIY4jq7Y2CA8C
lpOk0yAZTuCO7BPUrKdLW2huQOS5g/veosQIlWFksfgFU5mnF9eD2E9vgskZhSV3
AjR9rzf2hPA8DwRUw+zFmlpamyFHObmOBoJchZt3P4Pnmx1pXjBJ9Xp4eT+x63Wr
HT5tUzMwRadKptCcYvqc6DEgWbd+PrAr4mQFlsCrQDNIaaC/Vlbla7Bv594b3M8t
J3uBPJr2RY8IBXYHRCfigjaxvPpl5AbbBntXLqmDNqwA0Cz91pikiMu5/vIfl+kf
JmyP2K9f2ZZV1oKWkLCR1RP6urQGEgvxKa4CZ0LsqyS/EKbYqIzwGAyy0yK/E2sA
1oX3H2oGTmaeuSjA1uRkTASpsBtNSmLo3j8XThm5D8yKazWSdWy9bA1Qx4eFsAdq
4jAJpSpMZ7/hYg4aXNdF+ejYJI534YiA5Ep/l2S740cMQIcM0MIxS3w3qAebcOIv
b8uKfi+pryIVdzBO/nBzTdBAnYSPgaXskBjv5QWMYhQuomPamos4mBC4tuU2Rv2g
iep9FC++0SxpC/XoE12RzvoDyrwUG1K9M7OISou4Wah0Rm1dGtDZfK/vHh+j0ydQ
aSi+cfmaeSOFcmWZTOuFSQdoV8ZJukpyahb8wmpkSio29+Kg61RKaasJk+7ZFMOz
/pye5CSoVgJVy34he/A+G2UWp19/7TaGzVASnMg9S3+0FkyKfVeuzAbYRrIuhaMG
qG4KrlkE/i9LX0zIQo/V0/yTGDYW5BXwLeDchD/tkG2Wp5l6mPRr1P1Us64+rizp
c3DMhZSNWNf3BPRXqlK9+TgpfHdXtLLctoqYuUKKO7V/vx2LHu282VEoUedocWzx
3l5w2ReeJBP4CS8T4UWf6YUE+M4jwNQL7ZD2NXO5kqvl9dCXRvqiEySCpCNvh9tW
Jnno0UnfzJ+wZOQ4eTbrw92FZ4Uot5zQTZNK5jBcN+ebxbsR/vRTD5Mic7wZ1B1Y
ajx0PhyQPApvNzH5jbfDhigzCqvdjcQmC0AAXvwpwlbp422tGkL4ZTsBiuardQqN
8HdIRAicIGjPiWu+sh65Qlj8D/EnBUkijmyMR+50o+CAENipTkld0Ut0jyQ8cq9C
fi7tSPEpVGq2RmtI8sjpiz4mvdS41VkYzEAVa21bVLcHMAj1XmI+ZYI+M+hqNiO2
57Cha8xCW4fkXMTbc7sCPuSL7m/NzeDOZwxoS/JH//5GArperiUsEhgENUQ6x9np
NmkOHOUdv3C+8sc9w5BaayZGZsD+YiVAX+iobi46+masTkpmCItWfTvFiEUYZMl0
Zwr3dJCZ+q6NoVC/gq8TlHPC3An88iR/Rt7GMoenx20Y47PWqpyj486rKf0ekN2O
ofTek8ia0rAP/IngozNkA5qkqFcYrSKfdzl3D1cvwxauI2aNu3OGucjQq81mViBb
WTP3t1sFi7OeUpSu6lXL+VWnvZOpiLG1Sb8kVdrFcLq+u/zn6+xprbkvHef4NueS
mw31k56HMHOI87dq6u1SWPiNOOrnV/OTdIkT3ukZ5EmLuc1bHfTHxcfkg9VOkmqf
KKEwrmvWkxQ8el7ChUrLDrYta5tZ10veTQtmC95/dRuCCFcXXnsOko+g4GHFR2MW
SCRyOC7raS3D/T1pz7R2l1ceCdcFERdyZAPL7UIDC8r94DNBOECxlEI+o34C2xDE
lq4cNI3x1L7qIpTX0FW0Ptu9S2aCwwUnco8gw6qCUuqPKvYe0rka4pP2s8l3PzPC
TtojK3tUnFG/vovgA6cXxoHL7VF+TD6DzbEl5LQZarGX18LHg8SDtKboMVdvfUQ5
ADe7ugXSoHQ2zunLLU1KexhzweiEVkXiBfYfEj6rSKSVK7j0aXkhEryFpemyuy/4
6YTwFAVlyubDhRqrHtl5GGeV+U1Xgdgx4bIZvDemokMlg6TOh48ZhFdxuWsYewe4
S/lzjvmri5i06dG5SYJSM6qTHQbwdRERA278/zRy3UkrNxnqeMlFwrd4WmHrv2Xp
Kd9R5yuzVvkfYkoaXru2S1FUOl/ZwnbdvSVq+mQOgyJYI/rqV14xNeL0zft+VL+e
R+h0AnqX2T1T5OKzxVHV15pOnnjGpOwUxc9gj1GRDdb1D8LOGlcATUgD7yHokpJJ
mJc2EElDFbvjLz/i6y+jsyQ2xgZG4w+l/IDpTlysI8+Gs0U6pK53i34MYVT7EhIO
5CxDNH8Gg34ugZDaeIxgPEtQvCo+R8OVj1fzHO1qtmxlzNHGe5L8530keYJk7bHG
GDqcNPxzCvAwTdMcQVi5eJ1ZYDmQWPZ6D8PFq6cgRirYHJKJaO73oSeepnJ8+MZx
qyibFGqmT7h4BweLio7DxmdAg3cV5/j+DVK+MRcipdclhlxtUFP7oloiGcxfUjj/
qtE/UbJPkO0vNp6j5ErUmxaHIyeUR9wVmg1TCpacX5Uk24Uayy2APk870hQ0I1gJ
J5eaHZNYE5oYdRJIvDcyyoVeeA4L1QG8Q+HuFq8RReq3qIn4UDFD+bbEkw/7UXac
Xh42f1Ydg1ipREQanb471kBAKh9yU9i/3IWjpfc+D/C6Lla4jhELbfQLyxtggx1D
WW1hrLlOMB8fGOkez/i60ewSdOt7Ywm7r9FVvopWf0NNRXDSkedpj+Pv8fAp+3zH
s3ukjVaBBFTAZMaX7Z0lQdkTqUWe01HefzkUW1N2nPQ31QhQ3+vpdb6ovOgP6Lo1
4QioQ+wAILxkP2VsYuchPFnXMevLNHmdrvmiOpWNYTC33kNYwVmLnYPDbMKOs5Ai
xF9rEiR8NXHtd9XcKHBV3b6gpHtApNGuzPz0xTXOBNVPLlN81TnNOOgseyEHA0t/
aGSEDwCavpi8rDb+Q0q7bnJbWLfTEQGHXIG6K71w6Itv8TiR5OG/Q9cXcQWw0df5
QBhsHEW5iplF2LTTmdzxPY0EdubOc8FWu5kisj52XppTgRGOT5OZXfd1EpxrF6ub
FDPD/zVcZoroH2HQCYhb5CYZ77ZF4QIExYcxDwODTahf+LlN3pgGGn9BODmn60GJ
ILyRElu0lqME8NBuIjVUqR2QVjUuK7WuxfZaD5Xp50U99FyKKbHyypPIM33KaTyZ
5KM74znezpHLCA6sm2BSVkFRqePf+/3tBag8w6PA2/NM+6xz6eGflT2jCeM488jD
9SYFOBPR3UtiX/cuyv5Ultr9q+M7vtchCVzs30oPtJJDI18s1cuhnZPm6Cq3z9NI
Q74BuIdthHVCjZ6pVXO2YPRGeJG+JziI7qIkalazmgpsnqGqVw6X8K2qWVTHUDON
AVCt/8utnJZ8oHix/sN6FvQJQyDeABG5tcaEQp8Zgn8b27ZMLk7DWsoPrBbOft5G
kYroN7LoZJUSWneUNerw6usdRYPiiPrF+mRJoR4WJMC9C36K9lEeIg/5OyUD8M00
w0mn7AwyhzWZMqkCPYuXl/wCVXlavy3FitTS4N8zdm0D0TDmPdpfhvwC0wlFj42g
fiuxy1V6Ar4aNafoYjhj0q/2YaJEA3LxMzGhfl36sEM6ickvBaMKFlWAghohzLLM
JLOBCPxqf2v/FDYroF0xnScMb//LW2n2DlCcUbQAJ1yzal34QepIibO//z2Et9MX
a/eZ8Q07WdzCvjQ0WHl54GjYJAgTWhVKzjtPYFOJGvupNv9WcOrd9Mw8D0tCwIU5
Cjn+7p6VqRiTM68NSFqiDLJkNVRmyg034QlpeKp4M2PKg+26AcfFWEd5pAYuRPes
x/DjSqdPEL6dF/cyy0JPp8UqBwjFUMShXOnMU/AQdYhjCtri8eXMci/ww8uR/oQk
oo3waiYEQFqKCjgVlscrLx9sGlkK3Wtd8PugRohvHLOnELEolDe8kxXgzJrwTQ2U
y/Fy5Uv1vT0EbRu/uM2WLVbdN2/r27cCaWu4mjuU0NeUcYNO0S8i411B1TI0RCL2
3DMAPFfsOH4q7S5C7HncnaZ1Lyfrc/PFtcqfKLAKJhaCk7r3joCejIQjxDepHx0k
Nnbkw774BrSrJr4JZeJG5ZIY7bwsp5ELJSYcgRTqpAdsjCO8BPGKFX/ux2oTdScr
nM7yjmd3LjLL6ZishOFNECtAqwB/fogCT1t11NwK+l8Xd9QYSUyqZI9gd/OWBWMn
f+cxyehdpp3Uz34KpVO/iltl+KoeDERXRjLhpJwF+dH0Qve4UmZuEnaDCyBsmWbd
rB33XYVmdFrxHG+xQs9DAZa6Xk7up20N2sa24pzuAIdzenHZtC0lxH32uP8ZzlYH
qpmeeHK22Yku42tceYrZYqWxsoNNadMubZ7q1LBE5CxqIazHohREMQJA3hOR2bbQ
oGHB78wLi6+YlEAOWWDpddqMU23dyQ3w4lzroLoef91xqTkO6pW22Q7GikQYu6ts
u9FxC6svvDROGVB81JLUqXbOoOAUA34ipHAYYgwq4XrtN3pLr7Tq12wRRxZHVZfF
EjKzOgp5ZCgDYvfbevT0+5kxEZEYyX9Wqi8mTLM3oHwwNRVZq9oSqYka51AU1nxD
gEtEeynUw9MulsAQogfWau+53pf06Vu+ap1CDrzsQDK5LNoGYfNnSCMiqn6VGJvk
TKoIJiZGCxyQnAXp/Q9YHyuZR3YDxgLOZeGocjo9zrYOUHlXWqX8qd7vV2jis+SZ
YU3sCfuRwagJKp/gpx+gwnmB4A0ua3g6ODJboMGjojeL/URjpsr4GopyVRLjEdrJ
c4uv3R2QM8PXzTyJoFAtwYWGNjT7AV/BPJiBYEAmuvYq3u9WAf6UeMwjTrCY0VUg
pb28s6ZCkuhTt6i3y/DvgjyjtMuP2K7tZmhoViUaf1yfoNbTcAHcgskazdUwjEbP
757nExR4uKGexnsHywMIjAIM+GZL+/hiusAi6yMT5qUZhAxZRkSjLwhnxi/DGzCJ
PY8Im5qSYL2Ix/gk1jgt9YU4gD9HSvNKveTDZbFHe4c5Kcu+57VAMlPjSNaSiKZi
SMQqaLmq4LYv+ffIVqXSsey5pfV8IYfUTVlIK/Y2l1UQhdcQKD+Y+5v0LR8pVjdt
TFQMqw83Msyvzan1ZSu3GZYMkI9h/4PqIoKkjsH/oYmNbba/rbSbWAsF66X+yD5X
CkgXCECgQQw9THp8kehz6xe2o1++K7Fh1QcpPQxFHSpmc52OOd3g7uxTTMIY31oF
D4pAwIwWLHZF8beu1XBH5PonkbVzByZFzImXkIIBu+l1ak1iGCceYucyOztrmR2S
Oeq7ZoUXBuJhYuET2d4nyziGLZGeWINLEyYCZtzFIP63ad/pBOjV8tyGo69Ce5gj
RIEQWsfW8E7gM5eGMYA3lYD2sJhxIMFC5RZcwTL/GW/y8hVas+7i/x0xcYYW/ncD
iXBUiM0+bqmnlVSGnfmHgls+LdecXn0mADsb69CyDxIjo088zSqG087ARmDtBb34
t4qZzFk2aNjX/Fp5eSZEDGqRO5xo5eokkNup8GUsynkHPQ70OB7llnAwslpPCzCP
olTydgCk3SQdfNXWOHSK33V5npTrv1PzcxHYvCCE7vuwC4f2gzu6MVbFEadEEDmI
OKMwNNmJsk1ZdBoDDxW6zGx1a03uQy2GywfwmbEauRFsxxhYhNpqMoE/cvcf/YM6
D3Q1Lkg+xVlF8vT2uJvQnqQ2XaZxYqrtr3VLJVBefOjC+6VFLTDvqBzvengvCBjE
sE1cNCHtRI6Md855oA0vZKSfZzNJA0IxWcYhm6zw0GdN4nzyanj1NNqxm5Vl3OKp
YMBgBsa9akFzX+2CB1ndT7z41Esx3aPygMXUG6rduNaeftNdRFY2IIOjV783w0sY
g2w0kzHLYbT/ESGrkAn1GcNpEIcHLQpqA2XXnPPvCIivwSCFEyknaJ9b1ODHB2Yb
s6ESFd8oB6iSJL+Wgtko6KoxzDiJ99cyT8HPCWTtqc4m1Ce91m46NuhbEErTdohp
TDeoV2/8gGuZdvdNqPPEMwdx2FI+31Ja1gyhOgUBF52tzrP13X9Lh7UAl59rNurS
ziu2RL4SnBcjNsz7YqUPqfXypdbVWAZxzbNAdzG+VrMjiV1q6ACsVwPqkjmaJIXT
NTZjeQFSLgsAvbNgdTbaPLOAGMkoUHDptLuPP+bAazA+hc3vvv4x0JnrE9mdZNBN
eSLOEbdH1nKKOhbN1JoA90K985XVFwdf83kMt8xKC/3VkdhiLMBUkLeAqdFDIRMI
utEQVWKaHE08gotATc0sTL/TRQQg6/KsRIY0MDKqDmHXxoVOhSZvlIsQO2H2M7e6
883xKOueP9MPsxNBZWsq7/a2367rpC7kTthjEoHgSzJ2LAgLsZnu9+RENSaL6UOq
NiHeyAgpjg7dMJLe1s/b8uJ/O8nfly/Inif39qeD+8BFWIpQexTkc3KA3YL/NW4E
RzpaEi5YbcoZuuH8Zyq+Jo/CH2akjHmRkrlbFaHb7rLv2VCZucVcZA9ciMI10ZJS
2IHpGQLFoLe0ootuy7c2ljeJGIskS0sYqiDv+T1QOnpxpiPoETsKLhZjCIKjU0wF
gIIk4qIqTBDx8H9D6C6FK8XIEc1psgZ4o26SgyRG9gPiyBDu1yz8eRtgcv3wro86
i5vRLM7Jby8TFIMq7SVCCSaP6xQM4xO0CyuhFzCZKJcm/RZCXEaDrO+Ok3JHE0wj
YZQMPqHwOa3bi6Jq7CxV9N1GBouwFR94lnPwFO/XJ9UKMvUMnj7dmkL5+QiIaSid
xccSyJ7c1OwG2+udAWJtWKk5I5i/5/6EHP0iBqUOsubfKc6YTA1t6OADKCBPVIYD
UYryze7tiCOQp+uxazv9SJa7dKG25IiwCCiL1giE9vNUnrI4Vi1YZvz17Nwd1Xbe
IzJf2mCcNq71WsZUPYnn19jFbQhUEQ5VWXDF6nTyRFDIYEyq269/4gATAzEMJiju
6WLssRKR1HjhnAgujf5H2BxgBkRbTQ2ReVCwvrNbnriwtr0lnqcUXBfhau9rhBZW
hQwoWmMXTbm0OZXYHcDe4CLgvg0HAv47tuPRrhmJkPsycuV/Dn8bMTUKHhBouMxQ
J1WdJvwAFOGyjlXc9hdx34fHVimx+bYVOrFn9YHEWl+9A4B8C5GyixYtqRHCmDmm
CY+Q3NpXffC2TL/qG562gwAnujL0Bibyve0zdGvBgh/j1gvhZ4j0jdfWQs4uHQMJ
eMDR3zlcPBsIVTpf7ppA+xAe4QctoPXBC+com2jRVad9uf1FKGebg0827fS2NrW8
/IKrRCxh27T1r3BLQITjKoU0PoZrYvs++/YA8p9lb0krQxXRV1uDNxg7iGkC+wKL
nMUY0uWSL+aPOqIZ+n+wfdd2qQ3ImNvZeNIV4Xwu7u9AT9AtR0u8SE/Q8gkl1UjB
pTfyEltpO2kW+LOYmJUKV2AD38VffMR7xK0jjBuZ1hqCg/84M/RLeJKj/rpFmGdX
yWrwJT9sgiQX97iJNjNVt5PTS+U2eWu5XANDBqEVOsScodHJjX2BowhTUgSRRqr+
pIJSQVJFNa8DaTWhbcbyMJ3ZvNDTUC2KQrVo3MFNcFW+2Jh+AdQljN5EpNyhHQhe
BQxqjcLO6SPXswtgl2CvkrYcdmVNOyusnc50SqBrhH8eNI8z173oDCdZxmDCPQmv
jWjsUiDssmcMAJN2ssj9P2MwZTpV1gyeO0QKd/8cBVSwpgpnBj+MobO7dEE99Ab7
ODsA32UmRRWTlIDRGBNi03c67lwiA67/3cDiHfP/QVExr6wODdLKgh4/FmmIiYDM
8mcRLmZfjP9ZThAXkzzE5bNvwnpXT7L9dImlnAfghTTliHt2+WAq7xTIP/UVVWdq
LmxN2h4TIFK5DDmN+Du/SDiVC51KdZT8Y+q+N7InIELmLzTRf+SzIbRTLgAyS0Yd
BnEX6kqtQ3YV2GWQ0Kt0p90bjVtbhza7CdDIsaudy8CFwMALP9TOo5qSSdmaz4Ii
g7v1rp095W57juv/QKfdc69JaI8/wxkJlKidS5HHULa6ygvU2x+1iGYC0DL17Es/
T6y1IdLUKYwNB98Log/xwQTTmc+TzF5rvrfgc0QVkKG5Osv0IC4tmDsrTHvw+Y4P
omwV8XqQda47S+k78ECo2ecHeOfZK27a8Ahx1x/9ofDsV3EL3ENbqF7WcCAKXDar
r2OE089jZiJbaP9pXlOP13tch78GYf+yUmTUWdT2TaLSggE00jaBqpjX04tcUkKC
LRuIp4ngdBs9MNRPs9wotPK+tAovcBbdsdjam1zWXmFAB2Xe2AmD+ui/NvdO22/f
OVGL0YosaOSEhH+uossXgx/Uu2j/kGGJGOdCHD2ctnOdPNg3Ah1qenDjtmTYNwHl
UsZJtrK0y60Wd9Q5yhkGHmV9dsd0WyFX0agQuXIgQgo+oaqLQKmxcpYyViJB7SIY
0jIczjBQWGiZWxbysAeCWgcB3AH2WrMG8bGIUHRT4gx3hC/qyDJW41MpGYMU8cIt
mDxsM0MU05xhiLcTwe9h6laHI29ofkN6YSFfa+d5jBc0sNElhWM7qkmF78nXBM00
pyKR187bHaxpqBkAcUyrXXmMS+yJ5pbh0a501Udq86GwhPq5zFqfik3fYQBTWZaW
s3pNLEGmYsOU7vRtrC1/LPpaekS4IKire/46kvuD7SsDt3VuTd5NKtN8Z7b5dnmM
OO8XRwQINeD9B31WfxmChOmucqrbq6c/U2r4J+aIQKFwLlCccDcsZuXj+VIPcWZF
u0n821oPCQ5pNJLPXBaa0loRHQ3p/x86sYDLBdwiTB6lt/3iiOAyGx/uvd6Y5yd3
9dI5NHtd/1maITLMuIApX/vsvenokJtJjQ7HXzOOydKfCjzopKdUl7k1gt86HU+4
tizegW4/tTzWJQBNyVLMUqcZ7Xk2ZdFO1Pja+3qWTFIkQQQUkGZOhkSkVp2pqbhw
NpvB9junajKW0nFBHPLiYln0Arcgx4SUeI/wJJSBMrV52Ube5ztqUAJO28zURERd
Jr3aOF3bxmfLnuwoRHta2qDHBVU074bWQ8S1PJXnE1pHkD3mCmVdKqz347AWHiQI
em0ftkzzBFv/dsFWlNiqo8PD6KMcCfLveCNNTAzk/s6r8hOF44hUrN7DTxMkVC9w
9XLwJDsMlPqd2eexXIT7A1KhtwLY2SPXgA6lOyGlNTvsCTXV9s72T1tE6UPgqeUZ
QhhFstEI413Qtq+PpuPYlSCROp5KKlRd9Qa2xf+0ERqY2xZ5EbakzzlMMmQZnW9X
orvtW2YUHqJj0/LjbWtr12oFR/pg6OYAdcD4uXweaz7RfTliWtSB/0LwBBzEEao8
WcwjAwV7Kc+iWg5RxA4+1DYpFcuqZU9Ss638YmbqiBcTo63LhLPVLbHfJYpablhg
G+hd2pnHPsHW9fiGRJNYM3TKvfltiH7aTUXOClcc5lRiatl0Q/tle12DMoh5/E7U
ga0PGSwYr92T1pe5q66nl8NNbJvgbM0iXxqKzobGUQJx4TUhvHypzV511iY09PnV
ZGXZomua3vloVwbwNlS4DIMS0+KMm560uux9MjSXodi5G5QhZyIR4D1nQBsVUFRi
ecrt+oK77kKn0+eNpLA/jCwkQan0Ytczb1TXVNxsP28CI3mDm0+i7egfzSP7pKYC
kiTxLUOTjzDgM6zM84ykujR1lHcqloduGuEmyF8axktAfX38848Np7rEBcpwv1qo
rBxy2V6G/EckcPJIcHq/eBMWVwfQSyqkzbgI64w+SuTPVxQCAGQ9EG9cWhA+ZNmU
6NO3CugcR7Wn8lydLjmmyVxEpno6zJoLUJA0Xd7xbgUP8AM/mpZf6X8doDqCMoY4
Uf+dAR96nzP/kKVkPT7PfR3BIsi00YofDDRmzuLgA2eOOA49H/EwTEVzuS86C0WS
RIDVzQMKk83FUihCVNEkjhv+PnqSevFT3Xkb39qaDclW6VAOb+mBO8wdwAOFyxr8
KdM5Wcl2cy4wqfc5girFL78xK0NzEmzfspp84eQoRGPQbNQhuPZNxtLg2PE1vJag
BChoj/i1peVebIJfGHBc8bZKWGcHO0ZpAX78VU2rI/jLvOIiPqY3qTV58q3p78sF
UUrs+GaJnBIDp0PbR0odfUZ4M+yNFz/AjlZ7bg5UhVbvMX5zryqeIyzjCyg6tj8U
NJgaHiXAS/ZOeeD/R1gTAwUz27j/kW/0CNpQLqMtk3+UD1Rdh5oMxnLY/YfMRsQ+
TmPw9ZilwOB0xPihDE0VY5ZFk1QrZTT5FxFN4KKVzDUQvlqN0YM6/DF1PGI/IPb5
5JA1wW3e78XCfN7ELtsz8qmw5W9xkr1fI/ohOmIna1tNnPrOhGnZx2zXJwbPURWn
5H+sU2Um8/2hmZCAtG6GWvF+XWNBWBTarTGszOm8aTdFT2rmCKOltfe8AtsuQ8Bz
PNnPPSX6tpsS/fxnWJItFDJmSm8xu3nUQw+tkJwI8Xs4pJ1lQ7j1fsE9zjzzmO4C
OGAio8tqXho8cKzquOgRRMVeY4w0oXP5NUpuca/mG4CibRIPv9q2KhCa2qDXjwdJ
P2sT3VdI/rUTuYqYx6zyYiu8rP0SvG2p+qmUWM7QS9MLP98CFsxGdva4bc8qA+yc
MOrOqoJMx5DZ+UJe70isZiQeF9pV1WTuQd6sUlTAPUXc94CALX3PrcK3U9mDWkwy
dYVzhMUL3LZkfTqNG/4tWIy0iTZXj26UN9cPDV3ORyhb1Frp/Po3ul2pZsBjbHDf
lc0PreMnzvzr0HsdPoVXpWUkE5iLkTvhwqgLZVv1VVYBv2Qa3X/gj4dnasiu/Q7t
hexy1twi346BmehmoswC9+9mNl57ZWJdYCqepWMTCDY378U65LKKYmuJjN5bMf4L
i/NaU5BBVn3VwjhbtavYGNNpXscuTwK4pUmlILjYr+6Cpc5jztIpgDiq1ZuiIKPo
vzVY1SLm3ERshtEeCk5VFwRFFjhgYue/X0eptBmzX4ghYuSa0dw+EFcIiFab6WR/
N5+fqp0lMbdGFu5o/ae22iVWb7c9l/WziKWKaqzYPf7/pg82iK9iEjf9/3l7TZQO
jtduxSpz67CzHrsk245/j9WxeFi0sKBh34Oz3Qkws8W+d9cMWwMS1mGBBH54Ydgu
0HtFL/yN6hWbx/ai1NNsgT8vO+wBjuAj3p9JyU75WftVv/Co29svT/B3Pmc0i+y2
/df/k2znxwfEvq6AGtiHgqmQPGQbutPBOEgOaws0ywEhIFo9/ePTvDnvRcRz8XaW
4g2zZRWBuCwd7NYaq866ziGgRGWqYodavoeEW7ZCxwWYfKAGNMs714S+bw88AJ/p
mDB8mGP5buc08GGujADujX6P43LEz76gr8N3XeNkIXMiz75WKihP5MXp7kD+tv3D
WGz9A8OQS++XUxXkddwE40DUxWNMz5uwUNHwyeLyw3dcqviJXnSKsLowZKW9ySnn
5krcI2K8fOVLA4dOi+Yo8UerPUt28jCrmpXSq9d9F3bzBfEu/QK1x3dB3cFxqlaS
3o6E5Eb+00w1xnrdb0Tvmx/47Fu+bsuBBOJ135sWtuj3uHc3J1CIsV+qenrT10yP
LTY0SiXjVKep3au4NtygOZEOfd4NWhisSs6RpYN0z8a5t8xjE6jJjWQ7YHCgx/zC
w0lHbA5jNmT88lvwlS2ZRa7GiturU9vHqs59euAgIlObP4bZClM+fr4XVqjHL6MY
Xe3mKo/g1cYE0RknKZS9KZhhZjP8BlerOYJ5yX6cgIksuQC25H9hj3Kbh4fIx6tB
fIbMyHphROSH82aUFjYR7C+WTO65965PvqbqKfdfsX756SZd6KRTPLxja/439DdX
IL2dcXMmu0jbtdrcz1E5ZbEyA9T6GJbP0fcZcSErL/mueHK9LcWVLUfIHOBg0frQ
vZiW5EO6Vgz2fG3a5ieUmBwNxdHkwPqbFINapWc2+rK4f8Md5ulmqxvwhV9W37uT
D57QmEDJKbsuUF5S8kGlJlehKB9yacQ2NoWvMfxi9mxSro3UzmmLq85rfHuzSsKn
goQhmq1cmxsMXJhOTSh9dC6vuo2XKHs42ODGfbQHiV0b37SHTt/QeaNQxyhTL6mA
oEJoKWzo9tJdoUDxiaAnHDwj0wBa1zwLVafZDxu2MBBRoKFz9rol0CKnWc1lD0ZZ
D3apktj7EZ0soSfXH6BqWwu5QLtD5KSxTQ+pssL06zUzR3ZQdwY1RhA3IaUpRZf9
gCpA0RlkK3BXntgv0XNQFlZz7300kyQ5xrDjpQapGhdBHVxH43G2YI2Q6EjphpEZ
YPE/KhHGzyEQkrAmHTA8I5nyB7cliC0d+fx88YUGypy5CtMeAKDD0ycRzsFg3IaW
nkl+dwzYdJ0GqU42TiCjpLCE2s3FHVbZBQXYKq7kQ+iRDM+aHA3oJ9vn69roIEPi
rFAm6+JXxRMqIGkOmctcugsBc7ZUbtfHVcJPiT/e2tujWmtFod+qwnTyG5XnJB78
cBV7NrnOAA3YSzP6zdU0XkTlUBHpuF3jlnzzkzbhVKAK92Q4tCV+46QBLNvStBKg
e/Fr0X8JH3HgOz7QRtE1aaz8JI7FiirwIwLeyUZM7hk6016x0xmgLdc6RSSQNuOY
3BebT8hPX6K4jjSGNAkot1NiIve2RylXgjTenXBNWDFnzU6Z3XU4YMAa8XxQTeyx
cL4vPVloevhvlS+H++9A5YxtfCa5TAp8Oi9uq23aRJnKLR2t+VZcyRDwl8vT+i93
k99nEdMJgh4xDYWzidz2z/eN3YJok2OtGhHTTD0lFxgD5r0bBszoaWHzydwbPe/Z
8vmmJVKUpxrJlLEdc3+XsGU84XEzMWip47cMLtWHR3aBM1WyuY5vkZQNl2T8TLYq
Gby1fdJlPNccvdJCFEIixvJ2gE54uIDdG8ubWYjwY6HlYVQ1ZFpzOzBCHYnLQJtN
d3F9+K52YYTLa/KMfEsJbkENfy3F3JHpIUB8zOGweKw15e9TCkk3tgP4SftuoMrC
q9aS6O9nDUDLRUYSI2Vu8upF2g7NXv85F1Imgju5mQ46prCl+K1F+mcrnnJliRAX
xplcurRSsaoORopZIxIguRwcZpg1XD5BJBl61kFwc4L5BvGRW5qIIaNGENzZ6I/F
jMRzaf268p46v9PHhuAMoweos3it/fRgD8luHdY77l+wCBlTgUFgXt0W2xQJKTjA
0IYAZVfgUgEDJnTWh/bKHp73f9WVSelkM6riMZQtQd6ZutBp+x1tP2p5LMSVfrAV
BOtdWea1J+NsE7doS/Y1trmLWZWS4N9kJokR/jBthDKfx35YvnxIG3K6Ry6qYmwG
42CWVGDv8a1RQA35bQomQE8HLCx89lyb6yxwvJBfmQVq05k2raMJSLb2PO61oIjC
AgkMl09+a0CIaXDP91R7AYsli4CsQIlMl9w8mvIPc2grgZH6loS46UeqcWzQs2ZA
qNH/1g4w8ZCQoBQuWYyTSw+s+LAAfGb84bHpOa4MXsrY8ke3/ms8NPUsSdpMRO9q
2mRTcqolOLQJ34lxtDVbDMuLmV3LBUGDyfkd68/MeITscDi0G8wyWSXq5bUJD8b5
GbVJwsa8d3BUDtJrJ0rbRpxjhhZDlOYzWmXRNl06vL5877CmEnWPbBjUHah3tuRm
I1N+0bqnGbnBZLceO0PMoayAVnWQWDOm1c0KAehU3XHtvxE2yTdAsiq+loZSXnOV
cvpkiwgLCCKOgQtbO7RNsArD6ivwKCfOPrKkJTIC4k3MeCNvvtj9DxvrIMkUmlaS
C+xNc6hQsXs9innOU2ACl9l3Wuma9wm8BizCiSxIPt+Dnp56yA9xaWephVWJaSBI
Eh2c6ZHBcm85lxdVB9iAuzeetSW1vYgKDO9Ck/GxlPkZo6v/nDgzWmLthTq6PI48
e0bE5NJNckuQ4fj+g8UQd1kDzOfTbPTnZNdwgvB/gwz1R4GEEwmFCd5rWuGSSlFm
J7XcLYBt2ZrCQxO7TCnjNZwQ+uBZtX17cAZBQAjBZBZCDCQJ8RL2mM8muj8ROGIY
W6bSsub1jo1T5wsMTlREz7CCqoXfw5QPF6QUBhHFmVsoaboz/wDmjGpQsO+anHrj
eVGnZJv+wcDTyzyCwz9/2gQDZNPWYaW0nBlNpRdR4xsImV8+uppskkL/NAZi9rDy
Eatv2nTR8yocOXINqy3mwZqjTiTxpgnfRg2Ob1ziOWLODyV+keqEyai5mbdC/5sC
FOGGMOZ3dSDvFM92Zu670aHwkz9j5/kcS2ePGjg+Fxp+bup5TtS6T/z98SZAy3NK
b0ajVjKdVwoj5hEpPXttzfFv/77BKdugq8k6NzqGySydkFDJNKVO5BYj6uxln+Ej
+xvd2NWZPhygyK43e7OkQrA6D75MXnKERiOqLs1wXttRYAEwD+2XEWatT/Rnkr5K
rQDKswWFMH8gqmLDzy28u0fkSwAuXNcV8avo33lOfXWxrkCOOMABXDLMDo9DbMEC
dZT5c8sixvDpq08Xlp6R2niSiDHYIFubLxYwAdPZ3LFmfN8t1V15g1jha3eTmxye
haTSLe+9dVnrKQ4Kuy12cvRYTJGyfCdVoWMVEPHEM0i6pTqElVMTtuKyyYBnDihW
6vN/gq72UWo37vWFuGdWO7ljuCl7qWmsCXP2/lJsSAmZ9moqQ1r5UeIr85mkviKs
iL7Hjg/ylLs00oV+CzGZb76wFFE9a5uqqZ8+wyx7dDimn4UoGXukyC5rXm0i89xO
jYU4MYYDTRS+bnsMyayRhv1Tr0aSjff+P5xmlCqEPJ61M860zLiaYy3M0VupXGtp
Rf0GYI5RHBp4myMeX9nuJTqegq14XVnpOuWsVYVqx4GaTXUihrOqRnCLFSw1y8yW
NT6ouc7OPNEotMQJDv/RjgXwQJ6LHcYvn3jc+RPjT3asofias4VipkFNOkqpmP/1
9O5XDptnA6umxZUz16G7Z/FFajb8cy2CRAPa7mIEC582QXadRcO9fA7yjQdQwFVY
5IVOLkEnCNTTZ98MMQ/DbY+XZSwNIhvIYIzRgNuhM1s+5lGp35B70/oMAZwDHBSN
PRF2bzUAOHtXJWGCSkFxGkDeiF5vQqFcYPJauiHbHEf3u0MoroXE/6njSjrlXhNX
ok8DKjsdbfrFZbsVtd8zNHPGrDdIdIlF+Xt8U2Rw4OrQ1/rBaDcrKR4mzGC+MaNi
TxqoZxBnU7L9cczXMJOSxVxAmFFFY/dqvSpeMc7KRfGEOJmWakhSp15tENPueo4D
rqgnx+B1YDIMSOuj06ncGA8XVPziNHZLWiyGJc0xHd3/qk/XF5wLAaXHseG6hZAP
iCcWyMBmPAynbl0rzYfKrraq9ry+Q5BMjjYzD5k2W0Yf9beOTK9h+ruDNgAvkaHd
8Xaq0RT3/lLjQTl4haLoJIkIPsfg1Uk5g/jVFBvBat17woNYA069wIVcvmxGv65k
ZwmL3+3bLhgxwU367hgWtet1QcWjaxMuSBLvVEQkl9FSxRHmD7/w8lipyL90Y4yP
KOFZX6LOYXS1iORQPW1EEsnM34PbPwWqZOutxJs13fkJjyTcMYON9cYnlpdXGksG
DkvOnf5HZEznpDvkjb24dLKjdre8/M5G+3SiVsNgi4geh8xvlNB0BwlGOmqmhvtN
hfBJSebMc5rdrN0BqfYVa9YGD6AmSTLK50YoPk4TEBdrlLD1Ur2u+Y/tpd0q7lCs
GMWjE1eld+Ze2AggTxso6hh+GefxV33EWfY8Om/BR2qUdzHk6YYblJSe1GhQQ8G6
sw5X8hW/wnRzcgeLxn8XIgrh/IriBvoMuzmNSSooQ5WlhCfNPrjwEm/36dyD7N7w
C0so68pBqa1VZdBFKjp0rRbEbCjiWuMUwd1CTiYCGFsX15JSJbuOi3wwFChl5nEt
l84o1uttdj1dc3HYkj3bjGvx3TxtXd3VGiJDJCXXQqUbHj/yitB8/jQTdaFpC6nm
9nANz3zZmETpUY9Yrpa7ME5YMJ6sOz1xRes3uV4QyLfgUWQK16bBtSXHDQ0+aMHf
8jg54agL4lMiV1zbASYrW7lIEOMCb3YHWoEdwaF+Xb2pX9qLaHmcjXFNvvofsSs/
PuDMeYxf6ZURk23Sf3hYb7ZzXjySkbkvI4GGxYyEJ4T2yyOW2CYjMRnKb3x3HZXP
hYPl8txNpe/4n9e3yJhau5DzBat7SHhVbI1PBpnuDPtyAsvZM2TXQtdFt74TmurB
B2h7uzPXmNc64RLf7Pe5HDRElMeHxK4rLWzL3JiO00QGnYjuVAizzwJz2OukfNRF
2nr403c4E1XANxFeFtD3RLXZkKZ0k58amzGz2UqPO16mxgjWiTutCqEvX1djzc21
DTfiWuGzocIOwKtg6O9upaku6ABn/20MBHryeCVPJyfYmsiab0mhyFqsO28ZG7Xy
DmCcUOPQt9W9Wy7XG4IDWQHQm9hCcdHtAda3PhGsgocUMl5T7PqMsVFcwLS/tG1J
oE5i1Fk3xR78SXlaI2QQKVollvIS5w8qmdXK/cIh/rGk5sCyER1d319pmAYAXsit
n5g+fmxoeNuMBsvJIb0eCK1u8SHwPhpi/fn9fhwXcYpMk0P3aDPO/Tr/GsmtySvJ
d3c77HSc7kYq2QVr/vUI/noXSekd/9AEjhP3qNaMsI76Kh7eMTHoOVkLjqUrLXmR
6fcEj8LUAQnKBbN52kYsKGEFm+6fRgwfoGgr4pR7KfHVFSlu9gUMjAItIVF4V88X
QnRUh3d5bXff3HDRMSm0OZZNV+wJvBVYCaBuBr8bzhTg92lx6T9B8eB5RHsy3V+e
oFhFEXr2k04OGkTH8DchT0QqFiGPN2bWUgaxO13fMFNN6BkjeemSu4Byr6PPQG6R
8ksbiRftLpradICLJFF5YOLjnHCQ5aQ5lyZTpt3Ah+bTkkK4LYtI6Bvp0ppG1xJK
7g6RfTIRlrEozDf/xn6KLnvCF2y799xuHTUn7xITOAUj5d8zWJMOrA0Yh5R1HyUY
vaDNpZebvIhpo2NUjCqWky01CXo4A87TO39GsW0QMy0YEgN526LU/GsTAArsPmq0
oE+APhvSEMVvL3Po6+4DdSvSOtqlbRPlyTkcSgbd3UEpgaR+614VuBsFJaRG9bGM
aCazOKQCk78Y4JXZi/z1/ESxifW90gK5//NdKtaYKB/3n6pk4I4TS03mlRPg2Jc3
AH8BCvjxLhHuS66djyteBNpjjJI03GQhU+1gXsVEYUa4KmiHu7pcpYR54Oyb6KV5
1dVIYIUn7Ab23ZqQ3IcVdRVLNIZ4DVCoATQaxOzL91MEPt/JaTnxuYVlnwiBVwWu
6Qmaps6u518Cr8w42wFlvJMV8KGNRLDtPpx7We68aOZgOwxV+11DsKMV32Mpp16+
EI2l9Gv5G0qIQWpFeeMNH9OuuyFpLR0gE98KQfRfOKR7AB91J17esjYieand58Db
yDn7ZF2U06lUQm/wj9snLv30TJ5HSsL55Lfxxw2frgqHs+uPF37y6QoV9a72zKtH
IkJyyYxvf5ouXTma/Vda3jLTSsNSGdjJF0cGHn/TTJEH6QDxbmDEjKnRVPCFtEwK
jU66Pyt0Ix3NPxVhGdOAD+q+TngsoQtyA8ZLfQZWDyc/D8n6gyrlu8elrvfmM2aZ
f5e61U7I/17jnoKyOtFZz+0p5+jxeVqepcYE5oxgua1I+okdKm/bkwVzzxG6sMIu
DqIFN9wEGhOg+qWNl7Qfrl7v98qMTi1bWRB0MyNcecglz+FnkGDnuL12qju4o6q4
CMLnIL7Qt6/SUYtysWRN03tAh9YC7PifPsA8sIw1QgVzMUkkouU658eC/hcTqu07
sRTNy2dOuRUhyWk9pc0BsTNrcnhhwL5L7tmyCRAOh/nu0W01BDOYyh+poRS7gEi9
kSd1H25g+DCldVkgEXaLQkRq5wMX9DIGE+DYY4wmRaK/HrMpW1AslKniMIBFlxGP
KzPNqZTurJzk20jzaHHyBByhyuKF6VIK/n2rDLY1Z5H8emt/YNVMcL8KtKfRBMIf
6TxllVEhhJiwXvFdhLcYjQ/LACET5+mK3Y30bgMIGv8efVvRv8mXUS/Fb6QCkKrw
cjEmWllX7qWUsh8NQRiacehISauoJAckqBCQGygBbI8gWjdTF5WuF8vJY1toRa9P
L9IRWc/v81eVlxDVYOU1lN6zf8kBsHq63y5eyUlaVjDAmXA45Zivrlu4QYAnFnGo
6lylk4REOBMP7Ej6kowWcwe8CnyMKQcTWM1wXwLAqgTPpHjmn7pQb9fff8m7xM2P
US+HMmkASJRV3IDIXT08Z0OsdmglRiEql+35jlRrTRGfT5WIAxQcNtoUbfwHyU/U
GKF04se5qOK0Xl257S+n0y5p1ains5t45rresTe798rpraDaGslKMcP3o21T6g32
91KGrAAKQ9AzYdMbSqeBfLWaJmGgcXanAdSK++Q28rVZov9oO+YLpRP2dNh8wdKR
IKXra3fhyCim0m1l6W/K3mZl/FMFnmtKz4CGx+z1lUhbjvY+Kr6IJSXU0PSBgR//
SzT3SZxbLlFFB6yVO+f4rYg2K7/W+XVWNra/szYrIYcrCf9NGFVYR73I21dhBhkW
airrSRXCivMd+L4s4tmmQcHE70p4Ni6AyXuyEbint0qeEk29FPE4h1N1ZnjucgJn
A6rSGt6Bfb4xSa6StJ37Fxd26De5NieL3JtsbXPBkG2oJ9PB/N91KIJKxhXh0ucI
ebjQ4BTk/LXQfIrHJuebiVzSVyozV3jnu4Abt4DAZH0/1aXONh8WTxv277De6siN
Gd/T0VQuMti7Dn/xLjTmslPpaGSEuIMnaD0LZIwipRaSA2QcxqlN9zzE3LEqwASH
VQNUgFGJ3AgLAhhhAvg6gKKWbwruV+EwUJcG3je0Ua+wIhmIh3/YvMFr0HKQgUuV
RKRW7k6ps4tyOCp4+/1TUJD0g3Eoi0VgWMVUruv0EWOQW3OrEJZzjkujZcZ64I+K
NMzcdAjXnVX2cFeEU2zGjaVm0ktO+NSusx1sX0yHazRoSxq/GWbZg3mevNXzb4oL
+cTWyxd0fzSWsruU+iT8CnzmYP4TnSLxC8t6vXRtc6YOZnyn5U0s3aHkt1tu2dh9
HjPpKnQKfC6jdW9NZePGi+B0agrJG2GllBpNY+zmykyc/c0c9Si7wFhggBikXZ9y
qemEUaqEwX8FZQ0z6tUhCcs39E98Nmrofs/vzxYyi5QzWA+brg5Te0a7KqnX9EPr
Mcntfdoz40VAuHQXVQ8bdsFu5LxCdSVoEuboS/GQkfJc9St+amlv60WgYij1FKKT
5t92qDWLqOryO9S83NzbvTpl4BKCn31UEYevcJDcoxTSL88n5ns/k62RwbBMH3lC
Qz5R20h9jTzics10tCxGJWa5M/WhyYJQnZ/PIhIEUo7ohWFjbz3z8lnZlQ97gc+e
xyrl/VYGfbHA/0TSng39ocdWz7uL2wtkowAEsfRRVmHV3GFvFoagWlzJ2nc0QlSN
I5/pFr8JWPm6+o2cqg72kFunw7h9/xDigzmVNv+hyEP+uaTC9JOADrjdWF6lS7G1
VdVwnFQqX08dJ2AscxdKfVNlxHdEyEPvPV7InH1BT4iL36fMJP4JAV444+BdAcLL
JHD1I2zQXrWZC4AH6YSf9wbkFMcgJEOB5n89plHsEn+qtVv+51ZM8vbWIzLSI++z
JSDrvYzoRpsrlKCEoloqKnsaDj1enJMdGHVhu3ddeEE2xOTGUuzjs6sk/tZbM1Sn
8bqMpyApi4wLL++lebziXa8Iw7sZ0YJMaS5VNh8IbYST7GmpgQBn1YPGnFZs2FuX
qw1LedR8EIJaNGySAhtfMRzj4i6Ju7vuoO6ebAtncnt1HcU/dusJmAf1uFpOTp/d
30jgbWCdvPqrpfpkDTLVu1AbATLHveAM7W2XyLUNWluZraIWfc/6fSAP90pgeC3c
RzJkRdDm+xcY7r3oPgG15TSBrJ4OcX2wOrR4oQQqCQIsvrI3G/bYQaIjmKxG+ifx
I3enXSV9Urajk8idPsp0sj6asLCuYnCxyn89xTyPkeJVZUMdRNjxiK6ZdRkNPMyC
v0pDW/xwQTBfE1puvoF+bFo/kM2K1jy2jXN83PQ1Mh/WBLg0+THJUGVlE/Cw8jRx
5h11gv2Nw1GshyIZjgTsbKC4ixR/zGxj2I2MmZNuBYDxffywlmQ7s2+KvzbpO9vI
UnTKXoQKS0K6vRdHFWDcBMXFT0LRRPG+kZEdEwLWYkdfbETYnUV/Dn6SxMIKcquT
RuuVmru5SXOPqiQLu8vC+IR57ZheTv0hrn7fsy5BugvuYAJ2hfxUiFXI3X9TCBGc
OdsBxVkiSsQEmeUqHggQIcprDL+MsqpAyYshWAozb3UUtCEnCl/QmhKMUmluZafx
BhhIL0nuC7IsVtICf0Ok0ekVZUZPJyds269v7N8w1AXKo0QWQf5j9b5kxKoR/Cvb
e6m3gd4uwHOFJ9C7kSWBZIehAaP7Mek32PLrgzQfTRp3hIeTMaLDACKvcFwp+HXp
pqD+FlmSwCuo/jAcdmJGYVYQNEjJVIVgfMxzVO6vdqMN4dPcQFF+JUcggIIbMsiT
/J1NWO4XSj/nWzBo26DuTzIlpArqbW8BYx1WQY8YII8F2o0RORVy9V2KKnT/EQqx
zHrWsAY2ERL+RkGUgBEaWj1Onv+YSKVLZUtHLCxT0xxg5HZAFqK190qWBQEn7MqS
d43G6FJoMnEGEezmj07a55e2ZjxZwrTH2Wvspgg8pRdb+QYm5651osNW1QRYm+G+
g/Bf6pigAL+a00JQX+Rmi/e/XQuuLS0cCLwSKopPyOnFb5FX1McA3cp9gzrM0Fd5
JJ8PodWxbFuHsNxeo1aHzc0/1BBW/a2x8mLaBUFem2aEMqFo3dk+nk/uuPY9OhJC
tsgdReL3LI63E/EnBw60/Il2kZWahdLGSUlCOUjDSlKUQeciiuEAlPX/LF/ao9qa
dWyx9BpVsNEY1ntYJYYC1UkHG3FSTC/diyLX5QWCaA6WhP1WWIYajIlFeXVg8cO9
UEPct8Kn2k1+C07s0o6bhORjX6HQiZOQUb/3lfBrbmN5wrVTOP4XUAFBVl8reHXa
1cPh3hQJl7uruCFOiaCwAAujtUFxYwhE/m+Nv7laX6eB3VQ0sjW9CCxM0XwsRXu0
G3//7IGOGUQTXdHYaEYklgSYfLGuwy1Z/T/05qeMG/S8bYmzTGjJtpuZ7/jKuHm5
KQ0QjPUwKedBKsiPV3xo7Ck9AzSPVzmH2jKytWO7kvXgEYm9lWuhlrQdU1EgDBBk
z9sO6TT5/a8R0M348dMHEzQy8Frx7u9HhHzDMrotKfD83Zq1ZwOD02UJUlQTKyu4
Pb92d+dxj+uYIRdzO3Bk5l/+eO3WxmfcqY4wyXc3ajLP/pFEr+AaBW4p1a+WaCr8
F9wrPzY589JEupz27gv5WjfZW7a/uaq2qo59mTgENUxALoKPEd44RiENbvaxcE6C
C3JxI4VSraaji9hog751oKDNFUVTub2gHOY7rSZ60ZW0MCrPuROybYa2WnRdougY
5DnbXNhR9yEUj8dfTPn1vipk4h/H9f90sFvtLYSm0qLwxtNqvkd4ct33j74CERtO
EOZB+aCIjkqP4D5+Y1VvUVtvLPTjdui/zn/56VvVtiUB9CfCT4ALpG5DNSNLA227
tEHCt0W/JKtp9gvt1zzG6DbZe32l/bX6vmz8g+2YsGmhaWinB3zavy12BSZ5g0q7
8ezfkxC2qQqog7uLypgKivuE/NG+4MjwhXU5xmCPUiQUKxHabGw7dw14VURrI9yz
CT2/jY1AxU6oAzGn0isvaLxyOiNtrtrjHWmwsf/loNd252cU8/Dd6dR0SUBmz9ia
/95gidO2xZsVRFkPSB6HnhxFPP/DTfxgNDP5Fvl75kC3Pl9f27U1rZCf4PI6wEgQ
J5Wge7QqJWkhXmzBVykphzs3nvZqnL/PzstNgOstyp+474yGJ3Gxanvnkd+MGjRl
6L+3Mze54vsCXcTXFMrmYMXwoM8Xc4USxJEQI1N9DPXpyDsrxzweMA1u+4x5V6l0
O0m7lS2HqGtcUC/HECUTZWvX6hhG9bpEh2HuRV69aObAPFejwQWS50IRqVObJWFo
MXi/CY2s9e+qmC7OQFIThl5qTPK2cXpRGMVVpaBNZKtXMfciX8gBbLO6Kp7Eb48z
l3cvRET0cwTmdfk4vQDbnetCGz7OTG6MBb8WD1mlykxhC9HCISZfNdk43RiBQEmz
tqLS2rsRfCSDcWE/FtUcusNdJWt6AD5u5Kemn/+2StIxR+uBTS/7fTbxG3+4Z/Em
OgiNX84eKMkxDtyROtuLLfA9F2PbmryoPJNEHGVWw3YQ2PKxbjRhAhE0BkK9bjKl
tq917BL45N3uWhuapkqSpL3sg0fL7Vnl169ZygW9YTNgmh5+Db9aEvS2yQ9Ew6sM
xpilkRg+18oq7H/wqC414uwc+qADps9Sernw9xCRJlbAEblSTnPK/CJQw/3yyWXV
NFmS0a+PQqJ9yL/p96Cr/q4dGgWPXm8Mn+7YO/z9lhvYtNFE0lYifCIy80Vlcpin
P4SaNOFpQ0bKb8PxCW7Ek4sx9BmeP+AeEHVFbVEEKcqGfbhFcVkX6NUanpuV4qfT
hVFH/Lk2+Zk0LRtP9iVMtiJI6832br5SHGEqQ5OdBfGtuOOa86HCYYasQH58Oljy
ey+1ZVxGHMi909YmiaV1IDyvVm1lFl6YQggw6FqlXSQXUvMln6GH6dKIFC+GVOCn
ytQ61UU92YZ+zQFpCgpt09DcMykZtSa6C0udvPAY/GyRb6lnK8YDy/gur2xJ2xX4
jfEv/hVxE3le8lNhxYJOpl/s9fEyDzhUIF8PsEmNjVybHV1pqV+IjbtINPi6yOZC
N5BH1SAaijpHCWKzlASqhjXaAMYCHTN28mzh74lkuiSgJ4L5U4/TrZnHh6HPTm/L
cRulxC1ImDhtlvAUPhB9z+GAIjmIhIWEOmq+ebv8skRrEhXhpyV5l0F+Fb1YYAW8
iacapGf4wuxDe8xpXVxR0qDZE6XcPEsZ/OyZgO832EEhCod8DVeU3etyeGxYq/I9
2SqRiSON1YJHRfLNJoDjguGUkxQkPZxWZMxRidGvLt9WmjdRDqsZPYE0of4uWV7+
0Ezl3dtAGzMqZiqn3FiUsim3cWFoBkGXnpbfEFwhF7c81Ihgwrq6xRTtnFaW5/UE
vt+Hq41mGh1/C1QxpjrqF2+7QGuJ3/8Nk1BQBPGPmxBNHga6UP+2cT/BOlGl9DwS
X5ezJ06uDeJRw+mjyaDS2jDIPMaaZmAKkJLKgDijtiek1Q6eR78fN/1QESzhbW9j
Y02uFEgEq+IrthoFZaz8FzN2nzv/xL4YJL8lbBA3wXxDOoTx9ANVdWdkKStFpT4o
GG01VhMLg+RzW1V/ctVCKpdGoFS77wiSw0OPDelk+xGaj7mwxqJDOSUT9ORt/yKM
5u7bGC2dy2z8aNrqFhwueVEtyOvZuFowQcJAbo6TSrhI1fxA4/xKVR9fPp47ymHg
RzOr2yZV0Vhicdn7iCfs3EvRaTajQ4GPnBtxHzDLprXoGVtFu4QIl2xGw4djHScw
Bo0DIHtCHBPcbjKUUDTfz4K1/SNxVENuFdv5pGELJsBKSMdGdV8xbmigA/yqjD1t
pbjyjPS0OAzq310WTBpTyHpnzRgz0Woxl1sWl/y9JrLQrBOxFkDrcBlpgv6BL80n
IJAQBZWfxLq103YZoLSqLi75umolhFgAJwBS30OkPCcKAeLerKYhZRKiVx5SkNnC
ekNTFzYA7Rtg3NBdIm+3UL9yEcZlocnahGbMRCDrXJvopPXp5cfee0+sI9eWYC8Z
o9bATd98p1rV6FXhSUMDYwO3HcIE9CHymch7hNq8qrY9d5jd+sa8uTP3tsspmjWp
hFwanso5GZLbaOVqXtJvP4SzjriAO0tpDoz3IWhS4xrmV407LBq0JumbitlwxRMW
fEBqawvHASmX10fG+5iVoDH8pPiEkAWq0OC1gsJwRL7AzZObfMY+dFco2qG9ddDN
t5xWBy2Gn5A3HSkICtnWyWjGmuwPFXotSwNvX0SCHBIvWDOlDJZTLnZnt6O0jxPS
O7sF5d9/kR9mJ1kbaIJ6Xa3dwLCGAFwmj4EtEQ0pHbMbR9jg9Siw8oL6EvkLJyho
JBdT7wv0P9YIEVl7wEv7H3E6xrnQuSzWEHMhWAeWU58lh6IQ1f+mR6Oicu51mVrV
BdYf5C1C2+VKNLAmwxMklZLZ6YbWMLLxWYAMA49cL78egVRxtri0brp/c1Ei2df+
HCWl+AOUa3WfrG9vZICmAuYrTmhnKh82OJs4hyupf2aCHqG0N/0aNsOa0nJuUpql
94SZyjO+WqVl/N4YP5dVAAT2UvL81CsT1EFn4wE8kVtJSRXwpugJ/iBRey0VC0Mg
s6ddLfuqhdWYYlUknJvN4Q3Glf6YpQ809Bgox9r5MFRV5pedOEsIp8x67AlzeH7D
3TYiDi78JM32rBr7aAr3q6uLkpXhdt2hYMBb1dpy+h8a12ZTnfTyxPAIEZkyMIR9
qI2OIgfEFmnskIx13xdDQRTrnM5uF3Q1xlYw2aShW8NlMXiS2+Rcq2dpaqq5Zt8h
g/OdcSvR02i7zSlUbPY0h5e9uxAPOjZmy6rN5iMmoSwN4bgtdUdAjqzgzMaHvgih
H5Vhrc1n45QUTEqSbUMqKDASxTm+wbGe3I2IpdW5urOAVd0Ammp0Br2W7IBQaUCX
n7FyzkmoycrpTkDFmH8brgP09SW9ieFRqmVA2gRyBx9jx1zGOZsYYn6Y7W/cT0K8
ZFHl1z6ptPargjIAkeIRzZTfCZgJiRPz3NVjh84SCp75kecG2oat27H2I2SudPq/
gUWSglwxf3k0I9owVAnvg1RP5qlKZdpfCW+NfRMQJY9OA7q4n+OFeUe8Mcn2bBtU
FfDgdayWjEaZDULvmAjl6WYHLVAcTuczKG6tV9yjPrbiVw/U+eeFyKUQCCeOU5iX
8m3SpBagMLgAOgbInlwqZV5DOuPCmHV/KxSSe28WbHNNg2sieg0B9T7kcg7uBRd6
6V8DGbAZeSt/3x+HV5kod1Kdwo/aiBXY5wGlb3IKfA/VOvgE/L/Y97JGL43l9Uwb
wpPirf+rdv26I3Y7kqdOvikexfLlpmt3pNc52zsiSRXgMKM4Irm4FHb5stbbU60D
PCA2Xmh8R8ZfuQREpuh+XoXANaSP925nxD+Sgt2BYL5E612RpaMa6dsfOPUjkFs3
vkl6XsMLJOlmc93FpbpoKxYD+kGRF6UrF7e5ysTETyDkboFMtuxEXHSvk60AZC0f
rbwih3TE1aeKM2SCFBY0D0cLfZoIJu6sMef5oZFxwR7bCjdT2UVTGWewjLabu3Fc
UtOClg0iZ0L/lwncEE/Q2zZFAEzsjax5l7CqzHh6iAZFL9Ey801w306ix1rQodgV
waS4fbjIsIhiIKFYQsGyZ7t0gzjua87KaK12Rfpmxynd7kP2SnwpKpEscTMQ/oj8
Vdrvt3dNvk1/RHmw4sGMU+f31HPmt0N4eMuC5x/BjdiaZ7t8ibQHoOFyr0OAYC4f
c4VaCTSGrZ20Ak8FvBTlpZ9mBZl/bzOYUMpsGHt7sEQuQ6OaLdKfLMxRMhjJYnYL
NiIXuvnWU4wGAiHJJ2AIldarMlxvNPg71FD1Q4TcYSCz7VdY4M5qvjHljm015RcF
Vq7+DdanuMKZjghHCAz0ncan3+GcnpBRk53U4NcsZR0lVAX/6ffy+5iyDbQMGmh7
CbkKOEqk1OFmNfdpoclXvnPv7kfyQ4AzZYNauVNLo3482krDuJMemipogMxXg+o0
kNUFGeQoZdMPbzRvN4T47W91Xr1liwl7Rj5b4jztD3rL6Ta1ngYfHFlFMV40JRZQ
vY3WeuXrJz7UpZ3j3SIAUVD4kkcAlN8LdYXqF031ZnG/wNJn38Q44TG5A8xcoWcR
dTSQF5YeRpl7gGsezzrX6nvWScWAfR2CvwBmq+e7jDrDLTJD3+c3z3vgkQQmRAbd
2ZiTSiYqKPXn/rQyXTE8b7ObMI2vZCtUitN/tdArJfu1TXGlDn+guhMLW5aNjk/p
tRWcGKQeYxrNu05uRYgz6W08hj7yKPyEQEUCpxyOZCIoqiVK1CG1tCc8Ypy2MeRM
cnJl6EH+gyUZdmF2b8xtYH8A0voI2F+/bXPdBgRl8MKPGC/AL5JlPp0WzXy3yuUf
c5LNDRcR63Coka9tbFdgOfVGxVqcXsAMhEMMxxw9Y1xpMQ3LLL1A2BOh6TWDPMDw
kgaa30665N5brGo3b3C5QkGTwV2zr2QMjiTWDnoMvvUx5yR14DZX2z9Va/ZuCJbl
TqEE2RYl1I5y+rSgvfyBZVmutNGH1Kju4CZdeuNBgX8gd7llN+E8IYnEmX650Wge
GahU9MoC1bxffg/pvxt7Dk6p7MudhRyxbWpPbV5KUU6QbLbptdbE9mn0jEHHP0OT
rMgjGm0q765wkYaZQsSFSP0gxCX+jU38Jsma2MCwXjNqF0W/B8e0ftoWJBOeS8U0
Aj/cfL/ErfU+BZq7fFHzTZa19zT4ISFp6ZJ9VNaRK1p4tw7KMOKNiEXVpEPSGKAm
9hnbYoaIn5khmfx+qNWlCq8L87qNswdMLk2ftd+NMkTk9mlg0n9i6ahTNKkVVkky
uJEaoNGzkE0utBsLpHx4UzfQXfcqwXNo8XoU1QASnKQJI0OwO4IEtpg96/rwLGy3
AmP4IEgCyF1qhX6wwYTu/7ED7QVZKz53aGbfB9GdErLMDbVIvU27U6kj3zSPKD2R
YHXam1WIP4+T8iycFLdOaUsjtPLZ0Ydbel/G5Lb0MIBQ0dMg68eBIp3h4GAV7lFD
2K+U7CpSXRNRyoGFAK4WfkhVA/zRfv53NmIY+YmGS++AH9AQUIEx5BkhaRqzdj7u
fYfd5qm0J1SRjsv3hXpr+tzQw8GiRrT/cR+OL1URND9ayBiBEw6cMvHx4kknPSdI
n3peqCFl5i6WmuXob5+V4sge+a/APaSmedjLBZUGY5Uk2IgiAY1EV9Z8Uga7R3jV
SwRO5On2kC2Zg1YG31OnXHVUgKf8mdG+n77qbhbzjJgwx0Ix3EbFPi5RRWcbsvzl
5sb8O2lRTWkk+vkvQ4O9VIlTVD79a36ZzgaHZGzUoqSMvRI3fBY6rsRshKpQ9VVj
3DvHSc1Tu1tr+9o3Dd44dZpO3/+Hxd+iCRaqdIZWSsHlwwuPq09FN/HqmGGuzglB
wLfUUBRap4KGXPchruTU17dBE+hMab3qbPxXIzcE5E8sf+tY8bOYoy8fNuep2MIq
Vc7jVFM8JnjLck0ts/Et7k3EGpD0p76Hiru9hC/LXXWOvUyGMCU3bSlkjGlxtUFS
B5Zjrp9vXqCvPG7ituURsnSy/JuXkbiZgsGSCRd3zKAZSRISafMr25bLc83BfbZ3
CsYE7rPG9a1q/6D01oGe+i289wiiqDsodDVVAmz/4l4OMAOFqdwzwiQWlqoVhWoa
KM87S3HjN81etQN2bSCqcsqVNSEa+PulDnc4ZRIss3Mx1qoMCJLG1jrZ97l3/Y48
pADunUCijQurrLI8X6TpLMFhKMT64BUJei5MbDp3az/JCNvn2gqeFTc5B0wbrDgm
kOlGg1E4OBJnUaFZix2T+zopYutBlqZrj15WK4q2NPYuguaqzyKQZmqRdFwPD+y9
dkhYebmAQH7QPX09YeAlZ3wPg+ke2kmh7q8xDlVkau1vZax9s11AFbvLoZi24zLv
qIraG4CC1ykHMKbR9oFXvR3ogYytjtfhWRqe0I8tdvJVuUrW2bzR51qCDkgkuAMW
DBnPs7pogRd/hqf4dgJ/WZCU80Z0NP5y5xJM5JisnnqxUeMJraP4yNFGVZkhwOVw
UWutme1nW9RCsqQG0V4me1tXJb2RJa1SG7UpSye7f4/C5ouwtX9jWB/7P0syePkw
NEy39KSCgZWHPIi7dusYhY1O4yCR6UQVj4tzMSr0aZ73G93KORtJ6BXr+2P/Rppf
JxXsypOHqlSXCoNK0Qs8lesMG7Sld+tLSyigRdpxqBKrfZZdN15KJ24odAM5q3MP
f33B06ZreTC1041Orw7Ra/LjHgOEyj0EMhdSKulBve07HDn9gShz77uYq2Fbig1x
wTHUMKQnJRJmI4WBIZqEE2tfvy/zgB7NPssQB1djqF41pu9h6ay+RnxT0aJTQZFZ
U3XeSBS05Yqltpgj82nyQTDsr7sQOgtE5dzxJMcVfjg1SrrIuZUaQB3m9HeE47Z6
ClxRnkQcSd11rt02kAq0/t8mHo5NWols2QkczmwfjImx1NoCKkl/IIi/ssDjbsdo
V6FlUiIX3v9Ym3KcMAF9gbbYQa0hLEHUnUwakCSA1bS5zHzvLzFcr6vBPKygOyVN
KcP/C8/BEcjs1yjWKxlOZ54NsDSPO66cnsEO5rUlWxmmv+A3tDGsxrND/8xzerjw
5p1VaYfLnud68HCAjkG2QN1noReoiRkwYXhN60E4E+elPDUrWTtGrBi9cglmop5n
6JgedOFxA2Jx1oZEAsqw8ks4lKG1GiAluRUBEdXJkuWFBCyN6kRXEWZ+EONdDsRx
uCb6uQIB2yQLYZwUfVHrJ2oDebsdEMm9224q2FuZcZrYDDGHXnYlaogk3OfhjQJu
W6LTHDOlYORE6hMjtPX4qD8gCxKnhOzvEkd6p6rYiH/fEW0i6uMsJeNVJuBPUdDo
qtjZMTDkOJVWCn3pXpryjjJqW/Vdh1f+wTIHK9WXXE3m/x9w+3/ylGNfM7lIREY2
WEBtzsBuovK9vhfFGc5omSs+PKZZfaAsddrb9Ml9GilJUlqtQoDse32Epj+CwLx8
zCWke5xqGGqLC5bXR1RB0WJCnZWTW60+Uo2wJ6U5Pri7YbBTr3f2RGixv/hEXAbK
TZahYxjKnJotUKeoVGJSrq9xRrRbDrAX7FT8CRwCoXYzT0rUrmSlLjvmFesE65qO
QOuyFZNlgXDhQa1+QBqeCkMkYwCpX9JAjn5+doaGI2lvTQeypilTEoJwn8/ylh2v
0Y5mIhKpfy3DHq1pvdTgU0UGXvw6Vr5vHu+VotxJmG8ho+LGdrig+YYTfqG2dAbo
HqpHRHRCGdUp4PR/v8KvYShq9EclRi1vmjkJeMHUOTkoIr1Jq8BcUH2X5qq7Ojpc
LkqZ68fMtrfNqvDOfGbxeo5hxeOt3uzx3/SK3u4q5+6iEVS7sMISN5vYJmrGR8y4
5V8Etg2W8N8gp+CDGB+fpkvcdPeJ4V1z6Kt+obJBgSG+BSR9F52cA/TEua7NO7YH
qNxJr5RkaVx3/TZdQL9PuW1VlyXQYfT9bosFrn79yXHDK4yop5NQIvEm8HHkpq/u
RViHLQp8cDWXdBN8sPQwuXA/9hxOoo/gBSKROllb/HMQML29Yf1gXqzrKbT25mBc
WY793bs5Neax3VaB/ZLcigjTPlyiZgSWyT7IVY9k++g2O9VH/7veBg92mr8xW534
QMdqmIQV9nT0SxZbihxqjaCei6+/PvKC8pld+t2fzdznN/k/QmSKh3QZGC/dy55g
KilSWVTlCDnEI5cR3GpV91vAPQPrdoIf+N5uybNg2FEGxReEVpj3BF6pWvF1k6Wa
pzkyoS18c2Gaz7fCu/hA2GLPjLeM/Lvx48sNJ125wxmeK47n4JI5TW0GBZSJJ0JU
3RmOP34EU3vCQ98hlLvue0NJuwdmIUhxJi5Efg8pydshIo5lDl/TH+IwWqJnVPuE
nBDkUYxxtlRaj9F53+NCiNnjhxXNB7CG/hHztTlVGi36vpCVpaOsbS8CTgftiKQh
wHOB0jF3eln69/YYam9niiICjsbZEH2fxzL7B/bd/br+lViEyUiW36mCklm9iP17
MUg6XDyh81vBe9FaKDxzxQ+zeit+MpiuVFW0LNPiflMn9tmd5gATixHswKJQ02tO
sR6MXyCRZQINwOoIThNPAB6/sJffJtgTW3CpLelz7CevBNF7NdKnD9hxNkKI9mDM
vGqKec8P0/kI11cavPIC5Eh6sQaQ0HgjeHz6tNDh6S5YSAP83ddxzSy3SO7DXGgP
pUh7jfImN9jillGGXDdEXPzcYKoI/p85uuG2Lj9OCmvETtvgbZA/Qvux5teD0Xgt
C0swKIT+8Up9N0M2GMlKvTDZpZPl1LszA5Tc5U2jJlBdO5pt1pFHf9/nqB+x8asY
n6ujgoPDmtCh9O7yDEZ94DYh6607W7oTgrlcPQX0XNE7n8SV7y5U4AgusXldCpg/
yQtKK5ixMFtt0QUTH1wS7KPwr045a6cMg0++MjKxgSyF16k6M8bPwJxTTU69eYyd
d0+e4BbgITWFGd2ZCSp0bRq/yVF+B6B1QsVmdarSlH2grrzXqD1/kp54WZ3pg5LN
3NDci24+fZDtkQnE+gqLYp2kCtMe8PagTq0FkFC/OTP3s4VerS4qc+ba5ZqTU4eR
24Tno7DlJDQcGN3y6GrVfq0lrx9sQ8HHgjj/GFhuROYbd1J/BfBary4DGEN/su48
jHHFushDEGI/mtHO4FBmwXSS53ktbehebP2Br6OMr3558Z5RUfxcfQchUoaAHtSk
EoUfBLg5DICF7kPH79jPDjJXIZsyHVxORWgmlGQYFEH2xl4ptsWUzvC12hx8VwGT
4cPlVW7m7lCqyApyyCeCtKg//rCwAINygRDRf+Y9vF52jM1ChUGJ2DGjr83Jyghn
KRH/o2VGMt9gcTANVU09UYYWFTdvL7Xn7LY+R/h7zaFelpGDKvnoBEUvIg3Re2ew
gJT+WT8JBUYotSiidjpldK9w/LcjUxFYAtZe7na5uObbcDHXRQ95ct3hyTVclwlH
eMbbm3DyNqWIzywUOb44l+9m4koew97yNCE94zlj2SKmufb218W9/VHMs/FwQio/
FIXA1nDqpb2DVVaHsaUcrk/662TBhWM3AMRqhKkJAxLlCsB4kr6sUcBf8phuD9BU
KNiSv9g11D6UQ7fw8wM7x59zceQlJhdgJMRMlZ1HK352YC1TzBoIwAjPjhmMYMnq
YnVBfoypeW2k+Zoxdy5kW2u9frm/abn8yXKCFGd7tNanHIxvG2x4AOu4upE1vKIK
SesCTSkyzx2GgRWTPPyIZq+v0kbTPWSbCxNdmqPNIhxan0qxHzh2WHQrUo/Dq7MK
9GipO6enn9yb6UWzbaHg7oXMSaEmRtbzg1iUZsvDGGYy4oCZp0YVEbRZqKwpypQj
y2D5GIgWvNeQk54WCsj833WY5c8Ngy2GgYDuPU0xqI6Yk4xlniIOGizScc8FyAAz
jxpfHL5lLG7xKSqpCqYAwBWt7+vVNjQkRAoKMUFwLToRjXqzdoY+tzcru7G7p8SC
8SynIUbIO6dL5FNM3JthzvoleIvbFtdpsFbiTXLZzGEZsTVZiN7OQ/MbsIp5tVu3
Yvh3Pf2GAJ3q1oQnshb0F4wbHebsb4eBYxkdPLpkUWflS4hsB7yyutK91vVNCvVN
CPAd1J1o5sSQ+gagwrWKc15AK77bKUdyNPwGpTiaeIu9JtWP1BI8YXCaPEljJgIh
2ur+sgu5my7dGWYVjA2o4ysgRGcEMFEPz+SZzn9OOOVkyAt1W0vOgdqhXRPmMvsI
5wBr9QCcDKH0eGh4lslqV+dTVtohF9ECerx+m4ii8PYVnx7zojJ21WXw07F2xi+R
LTdfEbfCJCfT74EFnfkAmEQgP9uzWEgcEb3IlrmOQGDYbUQXlW0z7jeqT90vcONe
ExMZc864kJx1zir8GeSbQsT3bKH9h5pfPhhp/dQYgI4kp0HssWFQnFaQTC88jPnT
p5GTkjfVzn63bwFCheKFfd6N8Zb2PVts6j3Mhwj7Mfff3S/82kT+2PxUNXVbpFp0
s4Yw8JlqB5zK2et1Hm91DEBfQ7WDFa8KcJ29MjOBm3szrPQ/jwKiEuBlKbWzosjY
IhilgUmUKVpSs56atEjBUGyKR+DGMERJuCwim5z36p6dUy3cfLOPapePItwxOn5L
wMEhjAA6UJ8Ld54lDST9cD+laOD4bewmMrOPngc5kkLvntW39xpTDNmpHFRr1Qot
7EsFBMJL9JKSNg/GBWhlCk6KHEvlGZ25g2XNybkG39MCcM75DbBmOMs8gcH6KJGh
rraKUpnP8TL5BqXgx70uYIr9DOEHN8ZeYS/4TyDwsyH3Cwq8hRrDLtKF/lRcbMIl
FV0vBbpPT7616QgoBmFL0ure9BbL5xWYQkHv7rF62+UjE+Hwy0o7cJhEVOmdFs4L
Wp1eQAwLcrnKIwi90Pzz92CyFQGmHBlVqACoNLEmEDtc90gBd5tbMo2nSB3YVnFk
bc5CY6jb1NOLaxCMDbewLaWgbOFW2xxFkYr+7biZgJUMIEJwmYv5566SoSqEKUxX
ZcP1sJ2dWg+45sqEe24PhGv/XQ6ZGYhogRRSh82DNqJVv7ZoBqxVwfYmW5I44U0+
HOM7S9WIkE7YWCHQ+LZ8BxS/yM2+gLF9sBvl+CI/j91MQn73rN5o8n4FUxdyAJow
LZeIAlG4aks3dUcF2FQvsRSevm+ly7E0qhzEuB6s4cN7Nj/N4jTXqKuFlhU1pOvM
YNlJqAaqab7fM7/PjmwLDvHcF6TB7dWodnVeYPB5d69ae3VLp7ejpveJ2ZTk7woZ
9x0m0du4E0K9FOc+yRS6KjQo8i/5gP4kmfNlXz/eFyOQKMVNRUqIzGsLDSqrgogm
V3j1T8rNkae4XnImhehRq/fi+xFNOMDxnwgvu67lbVFcceL8K/orgJJodc81VBYQ
3K4/R//eDiA53OzAsOWTZNnvLfFnkw1psJxVWGFe5fF0bzavm+/Wu4CCIZSvQVCf
VlDjl6vi0z8vd2ZPA4QGKd1bHiGWl8IAQZtOtGIShB7aOWX9xvMxQvhGXaChWc2L
sxCAO7kv7R/bdJJ4f6aMJF81IS7665OeDsdBBZPANXWsBcsMV1m7yiagq4C7DB9s
yGkf++QpnO2oA0pl/wQK9Zj1nh96w1TZP1/vtlXJgwFfcdP3xmh+ErwEjnfE4DZ+
zHkt5v72+A1WGUmtvHw3mnc5Tr2U+SggDpkZvDEZVkHtUugh6iNgo4YIVuImpYfE
vA5LmQzqEe3KdxhuApChWgCHJdtKfl1X5aYC1U4mD8m+mOT8j4KAHWRwIN+rKqmq
n8bph0IrNBVdGyAccrXH2DVkEZO8bjCqGR1CQ3sXBXjgHuk+zqBIvk91SGY7NhnW
CLjmP8zmA8Rd5kMOSubzNa9xlzVf/PfbRDwM8LJhZozqWdu4sl6JCA6qRcYKv6Eg
GuRD5N+URyFZ+oNARD7GO95i4fOZxisUc1bDx0FJhVPMwJQSyXlmWWcZws2YzxK3
JthqyTnkkduH0Lgr0k9YzKBQ1FLxGJC76MIhUJjRArOndulc5FirB4JlRppa7w1b
YDhc7fRZ98R/pM+Eaj/mSGmS7PFgXOSrwDPdqnXWetdJLRSkxaWgHjRs92bxw/+o
EA/BddXlUsg5hIxPeBHk/MzgJT7Arr6Qc8cnVl0ulM/RFjo7RAbjr3KY+4yEiO1+
p9dMptrOhsox7lIHGBW6r6AGJ+/Krpjl8fgMQ/KrE8DLi/XHI0yFrxlgYwawv6F8
7GJObeT13eDMkF7L06tBh4d4d2cWzOTDWh37DeULZDwzi3Ro6142yzOJYabO3Cp9
vWOnGWlhuJ3FmtNSSha8Qk2lTscxRy2jG35Cf1yAh7UhTNPkX61o93no6W0xaeTH
XEEXsIFD23WB+3hD3uDFEP5XM2iNFKSszzYfs0fY1t+85B9WNL+EkNhL9bypPsWZ
6w8u13Irvka3Md3CHs8Fbi2mz/ulY5W994h/ooHxSERgaQUSdhluMeDjQtqeIVcC
63XPwYpcaQI6e/mHtTlJav7EXkUgekqkSHEnb02nIc/m1/bqFoeHrtZNqQ1vDXls
C/A/fKhh3hKNZ6p712B8lmqclx9Zwd+EYKcyOoarVcNbdgWdrpO8Tif8aAq1z/GD
xgWRp9WXIxpiga6dt42XfSwkjxw+2cLWEVFXqaz+CDrdCNYM3u18NqTU2/pnB+EA
WUfdWQ7QHnLe7pkPH2tR7QkBtUj59kaiwFV5RKOantzrAR6iMuDBVVOksYqVn5MD
zKbDzNzi6SvFsYMV22sjBp1TFcW4dbZkJ5c7DVSFlmDLbjpzFsQvzb+xiAurQE5k
DIz7A8hHQMCavzJLvrrnyOGw5B9DlSetUHV1Au9goEUdgAUVFzBd2FZ/yuJcF60q
RSct1msd2y4cw8zoNnmGjp86/kRuCOuZTbHT0KMneaOwhv4pgQYHEXVW1WnrD3Ns
9b6liUgyfuQ+924HUnrpgbIXcwj2orRQ+QSqOHqq/gJibQT4Zu04Qq7jf7K+iM1Q
w16cF0lCnM2QXJPLw952Rd+PGMDEl+myIXlnTH6Kw1dHaa6wO/xly15HMeQzOWhU
qApHMOOlCk/tH0b7kngBEovbe5gMKFLrEW2+Q6kr3vA1ZDDdobBpq+tZ0zYztmqn
yiAbDfeGyskVm+2m0x2onL0XeLYWyVCTTZtLGzCL8gUmBNtyNRlNancAfFe5lX1g
CmKL7xCRVzOu9M9wreD3MMIPmSkXmCHQZIU0KCIDBTfjrCZ95tNb4GC7bH1yTI9z
jG7V5a+ZG8P3PvDQJaAQP5jVpYlf5esE+wp4Aw5vluXg2YyXvOo3Ks0Hsh4ZtLJg
CRWiTEzSqOKjunkCDtro26rFZKyDRInbaCCMpljjrKrMO4RP9avfHnJJ84vgnTGG
sNHVigdzvK5RM4CabL3wQE/Noj73XD50/al7NqLggO98VbKxqdfvIB3b4i07u+kv
ndbIuuHtY5vIGEGskamhGBN1JMeC/q1ACRMJoMd4TUjQ29jS6DcIpwlynWjQ3HKI
poVc3bvdn5q9OFhXRto+2jKVrprDSEGipfXIra3D679NA/RkakQTTp0UwicmwQ43
iKVr3fEyzuHod4+BOsNi1UUgck3ZfKUx/TuGO8pHM9x43OEVBysRcfHPt8or8Ao/
d44FhP83EPS6RwDXuWQPvF+P3dFrWoQvOkIAhwinGd1/gqPcaZxGjM/i52sHpOfQ
agkTqtOkGNNt9ITdeTZJh2D5HM7V5NHCPXK38zF2DIPiPU1vAiKnT/l3m3aFqStp
kPXsa+cQUj0d066I4a3NJId2/ZDwZcg9kg8UVZVpcxOaCWwoqK6bQ3RjWdKjIxvt
VJAolmQ5fSKFLhGB2MMXqh1KqOi4lgNjWzMx3mxTVoXFQB9klvL8fu60EoHg5LCc
Wh9p2f4OmCVNhNzlXkM1QlinlzdGV6S9wqphHRC4JhP3S6rng8raxyxo4DkQNvfy
A/2U1U/wI8CQRI48bOhcl9fR4bJCEtWhH71Jvmcjevi7qxsiEhr1rL+l4IBoSDdq
jO5zcE3T7PxUfBlI2/KTbyYXLjxUYrbbz/jo8OwwcBLzcsjN9n6sbXmo9Npv7eeJ
tQNOV5zvmA11SoIqrPPppzUzEK651Q54FhXH4NyX257vciilpGJR7DtVTSf3uEXT
4LIvO41TEXD47dFstt0NERO4O85gbMTNTPvV26QtO4jab/Hbys1TNcf5YCYOnQs/
zb9zVIBCoZLnWrimGnZciTQ4WhqnRoCuH6rvFLBWR1tHWpWYAwH4QsBBLEpKobSD
tuG1bWcU62KhriRATMsgAv0ibfquNvsR/YzIctl+m/BtZroy4XBwiB1K8331q+C5
qEUGb48seWh3wJET9jwN1bXnebkdNiwCE15YZrx8utWDcy43a8KOnUAnA79z142W
w/2/CFi6CTPTfDlR8z66rztWGfnEQx6aznIJHD+bwxSz9U8GA1sA466g+tAAYPyp
IaibCiZx3MdlVmry240Rb0f+FaOXMNcXKiLggYF2jJGJk8z9jllpctgj06Vt5sAK
YrwxxQL5qseKBLP0F+W3OHSquFvY9jZ7MtySAKOyfQK+Mvxe1vT0t9xZxMsg7ov+
fU6Ux5JeEOQKq2+V4LeMHdk3pkH0BmbOy/g6GBs67Yf3Z+scpROWCigmljX1Q9ND
rs0jbOkbbRmsgnWfFLoJnGvO9GP+xDWB6ixzk0xOchAsORp6aTOHMcoX1XpYFjEr
VjtNTRfDH0oXaQS+nRGjgJdcgscyqOeOCYDzwJ1NLvGjTmocarv8yhBeWpP0waJ3
bxnGk7zJ+Ht/UGunk7CwobO6bFR7maCW7DuGxZfD0JCH2qgxGd7mxQsE+Z4rxBRv
BWWI4YEMfByvrHFluhaV3F7BPiXCORUfmcoFEw18vkYgePBbVgDeMmijwA6RR7Qn
19iMSYWfihu7mlwm1LeZhOVGGh+YOcYsynZJlHZZ7jmxCNkIHVbEvOALB0DpHCw+
ASPgF1TyqUo5pw3Cl5NR2pbpwOSJSV6nWsyxeEYazql3Qmno9NCw8Ix4+jxs5ijp
iBjKfFGm1PS6Cs0fP8e0tANaMCuvY6aP523GyfWnyz6k0/hZexVqOj5AYTqiR4n2
aZDUJjbvJc5YnYNKBSAT9qq90UvOO+XVY0JRHijrZidb8QZxBfUdF1YM/7T3ZwNy
BPsS/rYF7YPrQhNGiDSx34Scq3cULsH5KYtwjAzbLEApBfg3zo1SuRNAyg1uxWrH
xT+KwIFxEa1yMvAg0A8sB4VhK7D+qNZKvcmBCoJ58+egl+s2O+y3NzIn2zSpgR45
E3vKIIYzAxp6Fv4C6+IKkklDweOfICr0vOZG7q+r+eUXmo2SrEshy8Andayb+AVj
e23tAgcnz6X0Hx+Ph5GyzXHjpJg5B8+ESu0W5joqYkn85h7UB2Do3nDECw9G45h5
ElkaACybsMcrTl3RfBxEml321xSM0RvijA8kETgIJjKVlpWkabSZnftpEG3rsqay
CFBs4ew6eOyix/dcKhQxVce9NmJKO4EXVIJ0Xm2Q9/8T0elyQ01ZQ0TAinrNnsF0
6Cnobz/zqqc3VeCl0UwgYtLPp1KnyM5cTin+psl6Ouh27lWcNV+Y+jcYa/EJXjJB
g6Q64LK3e5GsIfNUFOqWUAfsNc0eHLz5kxGhknICFr6wYBXDVW7KqQ4Gv9ysah7R
QuKIzdfw9E7q/qK3cuECPVfZIwJ8/DyotkH2ngcU/Ez5prt6sdkQANlNzAMioUMC
SFPtD6Ff3xCkHRyrcXmqFQ/5PF2kAmxtTtRpF/CMAfT6ljZ/YQjcGCnEe51YuFZS
DkEj5vad9ASyPzvWzRFCajx6j8MIbUHPA2EmubVmdFnkyb7d+LAZuQnQh4NvNvlh
Y38qdq+5kmOyrG59C86yVnzDacTsj9ieA7SAvqGSKPXMKWgJ1YxpjHLSuPG+q6l2
4tj/x6WDkc0VFBzL9dJutZdEe65NVDNoSjnjWuM4zoVAoutruk9vVLzaSuki4kER
EJlkH46bazWqeyGixeV0COZsxiiNGjR7r3MtlzN0kiRo7ottaGzo45KWQYus+qTq
zX3wHkC6ED3Bn7xiKHpd1EZ4x6SDO4vnM9EC4la2u7Rwxns4QPMvTvjrPhRiSsWl
eHwKIKfyNFBQX72uSy6CkM1vh3+BCBcn4TQtb2FOgOhaOMWYrmtKXPOOG4oM3+4X
g7HkskwmGq5FVxxF5GdTw50U82kLlH8xSsOTPvfnT0/xfhIfdfo5VYPsg/xNLm8R
Ce2uPrz1eMW81d2u0MX4HiTrhZENNHZ/VxfoWCkHOGMFQ7Iz+KNMn3dh04uConQ8
WCNDGhDisBWQVaeAYiCEGj8ukTYuqlxkP9OL3cw7CetQhAOia+6/VwX7WGqYjnAb
ecA0DZG7fvCzCWyLGSLpltQhN0Fp+RG/LNIZuEn3WOYRH4XPgUhmV0s579gtCSyb
5Hf1jBeziDkyBH/XN8E3ZIMZufbRX7AzPzRW+r5N4IzgCeY5gkAixNRforJVC5MC
/Gchg5ZLP+gqpiOtSbw6ey9v4H7VBsjDLWjr5S6tb8EZaqyWU7a0Ph7NYv7Sfyil
KJj2OFmtWcDV5o4DXt8KcpCbkyE7Jtt7kbsiR67FX3fFMWw1C6HV7OT5e9pBYLxl
EvaBhmGYsT6x8NLihLZwPMslFuVXtWVCK9EONXtSR5Nc6Ep5De9YwOpKHh80et0k
2hWYn3Au9CQBbUKNmgoOxm/vLjXL33IvYyL4WyngPmgU83PLXGi3Gr/gOzyFPri5
qGLSoNYqFcEMaP4shOSwR9ZPaSY6AOnGWBWXnlqFX8TJa2av0PJzR8jji0nIwHXp
WccCuo4XxMExTyEl9Z/3FSRMk5JhgRt5DRc600Bn7HzqH5LJsofl/jNjeIB7yD9T
vXZOPZ6Xdvkjd5THn6tzdm1ltRGMF1MMTbftFQ0nt+tOuREBB04AdCF2STyZGrgx
hKjGrTXT9RsF8JsEJft69iCrCqOnnNhrD36aSsEtDMhSNoOrwcGwUvkwQtHzTZQL
p6itbXzwaHX+ud4r5ZkG8TTPbxk7L8wiv3bgiNioNGqeYg1wkxnOKBLvqdBO4K/C
JDGSR/jE5UAyVdAU68tK0scILz6g5SEZHX2YjqDdllNJdbIxzJNklgFecZxoVbhP
G0pjELLt6LX4S/3igYBs1BcDuqTcSIyDDasT/SXGrrtVtHUaoMDlI6TwxncbdzoX
8Mw6L3b0DE+/0zxYVcwSY6MadSyQqTOUiDsQjgPbuXiMbWovjbw7ed3SjRBs08PQ
3HMkim8Dc2n2Ci3rV09BmAlz5v6tzsD6w4dzLiJxVMRkXjB3gTOSvCctiMh6+pgP
73dvK9Ra+yp6AxHG3EfYZrayOVb81qCeN0uqr/aTX/8BKXJM/0XfKu9UcnApB3QJ
uUxUo64x9/rmw+ArM5hQ/3ZDxr57TIBI2H8+r+9PXaQlPwqMfHZXdtoiMCNSq+rF
P3jeIv6BwR4RYLa4W+FVkidrgjeqTr6G0Y/tnkXI/v/DX3gZ2rhy5IF1wYfYYoDu
RyitmFm+pljCm+WwnAZ5ucLmPmR/vE+9HiYZ8QE1LWpJkkivwXod1IU3lTyhuWyr
X8CLB6Gra8zKR8UizVm1VFd1mM903xbLIBshsA//hI+NQhcA37yVOEoTr/O2C/f2
U0sAQCfophMj1urCzFQCxGApwnU6nX0iuo9bNSItZ+CyRlFM97Dd7Pa8ig1VEQWi
6m+sMxExoL3Rly80VWL7yVHQx6rG7ns7Ya6QeRUKYhRCZhaJlyCnHe0yoteHGrvD
RPLJ989i6yZbtyQzwl0NBwXNopgByKTxs1A8tT3dYE5WD8bgUewW/o+Ybn+xRVPr
529MZXXWwKDpI/eZZUtexxVjfG+GjWqWfJ1Dapwn5ykB+aHpSHsJZ1IUXs7hWzcv
vbcOvpGoJiFfp/D+dmMviYVprYocWwqgT6NltPthr1dloJF7cAbnGrps1EYMQSHz
VRbtWHU0oS1JXMDpVeWE0yakY3No0sfc7I5tXSxYa7Kanf9S/sE2JtVNkfjhSnml
Y21dexvXPdwS1tsWuOOtkN7x4eP4XLcOgyby55BH3KKD2z22q2qTmq1EpQG34QCQ
8QmOXt9hv7VNvpkHHp5aaX3G6pkmq8tPtIJNSAEl0TVzHefjVjiQKMFwpfIow7Fi
gRWMR3bltzljErBB8Gy8MC9r8VPPKQssPg5DH13y8OhJ+K/rUiVuiNtW8wcynXof
4e4Xy9bKw4mcW18i53E0KLNSE48zLHaakAjv5aj3ZSGlAhusUjfPnevTt/r1SxNw
13Ahpk3gwUXxx/L8x3I1FTO5TTMRo26KBSApgDePABHqLQ1BOX3LNeT6ehUPY5xi
r3vLq4R1pxobs8Y2iTLEQyM4KeZCCBuMRR8KqN43QIW6g/azeEyr81LPrRo5gLNC
0QVNVIjmbgqEvjIius9rJlD3dpsLT2GnIsg90IK/PYPGBfq0ynAgIVaJPmvd7Ak4
lvL9SlZZQv6CIKiYCgR4kOIBHRXswXAzXmaCIbkGRmTLTJvApLEzxWs/GmbciDww
uSjmh71QjuzWdldzCtXixJ9Mtb1VuKaKVLcBUxKsuFkN1IX9UnBxPjAwI2INkoK5
jX7oyQ8UP1nNQmo2VaS5O4W/pemnpvf60UnLpHh6vrsmkVw0d9wrt63tBDWB9S1D
2TOgw2x0CTL+EM2aEGLlnYaquqBqO7FcIvl8h/RHbkyjCfVFhEadabSFOqj5yyXY
bsxtpcOqzGu64Gw6BTbsxcz4ysrqGMTcynqxSO+8EFNWDXgT86uETD8XhcW25Mdv
+lYPXIcPdVUxnl6C0r/XplzRsRBgyfodGmBp8X+0R2fboQbzUgtCUEb/DwtbnLCG
qaFSmSD8Zo7pgXuMlwO/ZxOnmpbYjx93D4M4671KnS1uNCVj20NEHibiLwigrAwA
SdykQRK2/jzx6zuzrhg5zmvZTbyJ5c1NDww5B0IY/AeQ4gatI9iLWkfGMKzMIcf3
5JXq5UqqDahAqNhnKbw13xWHp7ej+UygqXptgkQDy+PFmsEF6ovtw9/dxNW7iPf2
mOC3Lcp5bOSQjgKvOuFE4Pk0XfFZW+h1g5xXghqSUK4LRcedR8pU/3xDnhmv/b8w
u9GFWtnDAAj8zn4FzVfuSLDxXQopOe/zV0QwpoNwhYnm4rcwhLowgYhz6nmtSPLX
sdHx7xCxvyqtrgnZ0luoaJ8kGKkR9J2VHoMEJ88JuJiaknpIWK6jwuAB23eUypS+
+H6FqzRZyOtfP5LhiBG7Cq5ru9Griokj/B9Fjat+qDkIeRAjKPB5gWjddPA6gXEA
FNpIiS6W+E4viKO587DNwFTzQh8klagme9Skz7hZGMrjRrzuR3NzBiTvD6df/MTi
D2FmjSfvgeBXUl1osOjoyLCCOyWcW+Vl6P1TUiQdkn6OULhgqOPCn05HMvg50WV4
O9fIeXV/Ow2LX6ZAz0nF8Xybkd1v9kAABnIVIEuDD+4I3bg/2XXn9YV6HU5mbNMR
7Z4yns75/h26GmMDqX6qaEF/QVwSxR0f/Xxzb44vxM4SNQMeJXCak53NEY/sFNrz
DliYoJ80KAd+CxWmWao8gg2KdpQFRKJTs8r9Qpwvr8guSb1tHibbFeEHjNb5BEc5
21fELQjnNdbM3pMX7F94ETKbBK9CvjDMbaspn3sb36XY8Jui6j3U6dB97e0p0joB
vsa7OH0jAqYdgn8RVMrmho4DsDh1AR5k8irSj17wTyY4SQDVu/42wY1DFh9P2ZLE
N+rDuMQb9Plo/b8Uu/QwJndgmvBU3WR4HZAwKvvudX9lzOW0FmLS+u3P0cZPZwCM
BQ0ZN1XbqYusgkwCcMcdJsreOc3aPoNYlswBi6PmB9mjRG1/yNGmSc6k58ivwuOm
jkNMebFY4JOcLn8YqCk66JJ8jLhrfWzMAoPbRxov8rPvRuil0F3JMJ9yS9fKH/27
YHnhJ/+7Dm8+ZxkR8w++nuHiHotTXIy7OmSWK+FkvpRXpO5Uxd+oelTY7oiT9bM6
an+w8uzo6ZZw7eTcTMu250V2A23G4J5CJ1OG9hzNyaBCwsUBOCnMkVCtVEPtl7Sn
iT7rWXwKzuEXbtslorUfZx4j/M4GJWVLWyWfIYNdlsd9jaGgC/fg0GEYAMv8IslL
9dRVst7CTS/Bx4x3C7R6yq3/hBYbswqKgq2w5c+Lck1i46dKSa6wvKr8Sp5Jr6Ad
tS8M0T0gtnnER5MzwPgkr0EyFhm/Yhsgyq5JCPlGXqqJX1eUKgRMXu0cI9Uak2hX
R4ZHabIBqWobrKwZ8oealkUCnVYyoKKy3wU0NfomBWIBNVZnB8l9R5dQpAFeVYdN
wJMKn9YVJpRzQBfLgx6+y/rLz+TXBRzQfqvSibx7WxYr0CGdfZib5Nyby9uXu6b2
lez8DOeMSGe6TnJbvHWLMEu0ZqAe/JfV1awg8ZrY9QBjlMzZovebFrn44fbrgIje
Ok0Tb6ATNn/AGqrEbyMJ5QdiMCIw8JjTU0v4gfHDli8BH82HJuWoiut/Xi9MRkUn
6A+VqLZBtlJriF6XP2UuIplY/emPSQIRa86HBSb9doGnbSQ8Kn/kmxJAQ+ARb5Ag
Owvb1y0Txh+d2rmReXqpfuDildh4TzBNBHd+w1IQYRzuSH+6x9R4IqXnq5xvWVwh
aed5oPl90K6xorWEIgTYJ6i9yYpP0H6YyW5sKUwD12L5xw1lxJ/fpMJpYrp92PMa
ZQ8yTGjZelTavUelnU8sQtcGv0aSgx8/rffjbgdZas11P2mZKhyHtueT5kHu4D9x
yP7Vab3na60hj9WPIVArnL6ZYcftJi3jHHUziTR321+Q5DioA+VPF0hKVKMQAnks
6sWDeWSHDHJSRrNNY/VGGTAvO57iVP4WeWCjGx2SZVWQpCd+SGSczF09wRSwci7z
QLF0FjKLwDjOo6v/ka8qOgsC2oMuogHVy13V/oxU12PxwRagi7XMMSVCQyeItoTn
WmIEu3qi7FAwYW+TuD+7zOXsgkgngN34Q15c5GA2076MoZmhQC8Ambrh5Oc/eGLt
XGLjm+21xYMm5bVWlWamkXYMvx9otJV+NmfLc5YmC9KS4vLyoBf9QHHKa0fY2e4G
HpzPO9ev6uYPoS9HlOmOvxvpzzjANafJI/3scCH85dg+qa3WnBdcNFFlzCM7yRLB
maooHpRcqv5s9hI86HMpq+jsW2lerOY9xC5k3qefj5vtVbsf1ltlScF6iNF3vsLk
d7daLt1utGiu2Qbfz1TCYAil4LamtvtzRuRdrIKA9WCN52+yvmG/+5rPNM93IfUx
Wz3UzhFEc+c5JMrfl7cTKTQxqql95OfMXyK3lEa237t5/qtCHPQ4e41T/wblMYzF
LlmlW64hSQCIp0aujKX3YUGYgoGPRtozY6q2nKVnPe3Hv0cKm33MtPE2sdOjIqEW
hvTRkCpMm84qgAlBje0sYnuvFeCFgHVDPn20yfpQI744hsnM9C6TGakAIWT5T50A
YWfvoJVAv/p00/eYXq/Ul3bu8KD0OZvQWArVXs5xU2VBihUGABb1PMC7Qj3xtur+
+g51VlwFwvh2p4wCjqTrukJ69vOEaD4WfzXucfebPv9IVf89u6vXWr3lqZLUqJ3k
XkhD4S2luO3MM542bcrV93j9YHkVSwWvfB10VtQTj/i12k8M9DX7ag4nz/6ZEMCV
oQ8erxuZy+Ucj82+WnSMo1gPVo1XsfDx+Sjjah+RYlXuzQwXkXpFRmC4m8oBU4hO
EmitC2xbtAgZpJNDVuWLoQsVjD2fIXdp/nymKuebZAhgueU4zmvUzjkjlcBXjuCt
htvHppmaSDvCaL+OQWG3kZhu0jhWQhU1hZq9FjsQa06TiBXjw7MwC5H+0cabnB9o
wjdvW2IJEind/xz/YHWxfbhLA4UprRbWjZ8XKtnIMMjMEp8NWx3qurqrazEvTmZt
CaXcD6vETjbwaQ3h1+JTPbrcUpEQyM0GLaK264xk3cbqn0llxjRKDZ02xe43bENP
SPj4nDpvo+FSB1Ews4O5HIvgVewkT1BVB1/vKVsSqg09M2faRP7YU6ib99/Tif/j
vQmogn8+Q09TUMXJ/pL1TOjFGQgbGDRilMqaRcQkimy9CHnjDUC+3k79Mzl5Pzno
SYpx91XC8ajtuhpKozPCGkqekrNpOjq/swmSrjqHGgkt56n9mONRFDHAXHtE1pJ2
uMK1OB/3hV96xG43dKcc0+VSjU9EEvjiYMOLQ4/qF7AAX/NrZcd/6zlZXJlcMc7h
vlGzz7l65o6Bi4MUFs57mkdm2QE9fNplg+2dD14VH5i8EUAa9iyu996E3ExsuKkS
KUJBBCrqY+E7g3naf2WNgNpKg+eeZnf98hyfxdH+k+FLRCQ685G03TuJGQXL4GVE
yTMvtha3lYm/oMqn6g3xUygVd7m4Oqcf0Q7EqSESQ7zdccmpe3pvJnQlOCfXhTrU
PJJtW+r+0UHdZfcEtkpwfThSaQEIIdSfBEC3B3jzFFgYNRnD/fx737RB649UmcI/
MaG5UGpwttfF3JoEwTh92PVbq/sVR+DBXaBryd/OMb/m8M2K0sfyKWOxjUQZTs79
a4gVCKdaRpB8FopJWH049V9VJDdCa2XYYo5L6xuHOOv+/ewGv7N/ypQ9/wpsrXJD
UcDzep3VhDqV060yYta58F9QaxPGk6Avaa7wkRsPKv5F44KdirNKqjneKT5EM6vF
KTJV2IVwFLid/sHqC4xWiId0rDNL8bc5S/tlyq1HIWj3BuYl7CtanRI4/Y6en5hB
d3/ZIQbpqGRM7stmT26pm+lOaJTx+NxeHS9AEvE8OfLPmlBnyfeW09dyY59tuYTn
9mHLYqhjdCOAb9YoRSlxq4CC1+Q0OwqgoZ4nKCuJH7xD4wW5yMz/mi90fSWTI+y1
8Lq4hljJOrQd5Ywa9Jon6MI5K1wU5nr55y3W/URrkCVoZ+tLcuNRgczo6uWhvARE
13W5hkQ1cI7Mlj19kOkxITrirsMo90Qk77w0TvUlCwMnTSFoDaOkq0sozLxgNPWh
1CcAiNhBgDdxUpTXNLI9vB4S2hSHc+WEKeChp1k2D/quLjYpTJpHh88VefWK0W/9
ocEOEbVUDMMbJlBbT6v9IBSSYksaEoZKu7D2rMHciGcdZnH8d54H5iw4jSXgWDoQ
v4NXmVTMiBP61RHAtUqn0eINnCR1ZylyXX2w5H4FxB+283iZaK+2GHiqieu9PQeX
aZP718TWoHys8B4RDZ4498xda5qCeHISn62tEr8ulUPItkDBrhw/1lzyPzH0AIaE
vBJFGk3oRscWZpiSDDJ2c9C+/ZbpEiSTpE709o0vlrH0gtEGu+XGm4bbnNwmi7pU
uyrqdZebVE1KlKtEU+l7Gvk4c/6B0EQcZVLshjCka4lhJ2epq+8NGEi0JhDBw22B
bk8hyWYdDIp8ZT0TlHlMbHREJeqmGtSFoJigHOZuecXnYdtE41P1F2DhEH5s3df8
a+kWIUs7SaRo6EN/mHC7EiXJ31Cr+dQ4Yy/u3NJpQBSFM9mK61nGqDfPtwvbCdHU
qZsRGNDwYr0RJ0HKLQ0UhYcuACmweVW7uijOcAU0z8m9wsdWY6rf2kJ8L/ao2ch7
Kaez3wcXh20g0G2aNI/oxhynvB+hdkljUZ2k7Uvoh8nWkdP9oAw7u2XnrYFno4I+
peQ2PKwgUfqN4WMUekw5KorIJDSMWxSh2exFDZWXC0URwMs0JToySl8/ZGzZDmcE
vHHWCS1/d5merwgJ5TYW9xG8QFn26bvqqZMgQB+0fp/v+B5Ih/YNZcGS+G4ysBbm
PEfBUqnn70fglxnmkNxIq8TvRKg+qY6FlFkdJFwFrr8Pq2eXEByieYHjggr3/NbB
yVGJ+ujTy62eqe070zUSNm1mkvYs3YMFv77aXRFecqZQWpgf95AmvHFTn3G+aq5i
whpJTFeGRmf7kKiQZ81TEmQjHyZKdmUGr6sIE8A3ZAtUOOXzfVsUhMAQyn92IDzW
xwVg7JiB3ShcuwLvn+h6ns9KzB71WycOBt80AJcHVvS8ZbXVWhIEJxp+LPxgFO4A
nBj/IVEZx57YevPN7oRrA94wlbeVADtIS9KbePXOgyRqsNPbCKkzyLYpSRTf7F2D
4yonfiZW53MB6j/o4yqH1xZI1nOET39Kpqeh7IBkn4UpL8SNG6VftE7aHvVXXvDU
Pq+L4cdXQDygJCvRtWiJl//pu6OBtrm1Vp9Hy+XiPIdfrcm2tAhKmblR44NsYCHK
hi0lNe1aEKmifN0AZpVBY+oygqCqepqObMcHMSpRJTS6zMr5n2CPsvWIwDWLot6o
6B4HK3u/bEJFikNsXhqSNEcX4Che7rjHW/4yowQuSWj1MEmjHVdwiV4hRH94iiUO
JdZG4TERw4yi4bBKn/sRJA6n+5+gN2T2z0L9ePEmykDvKIlbGbm0MQ17R/8wqeDO
/3/pP7rw5yfzTY94bLLIqhQwsD0v6gCEgHlYxOuK8RfwRgqNvCnYytHhn08Ep883
5q2H2MqYWEnLBilcjfMwy6zTn91jbiuJT0qy+0nT34vu7u6bK2xmc7qGGiDOjZ0h
rqjUiP5WUsse9yfGTvUBBXA5cPLVgynqFCthSDLta9PcqTaelwt2iW7yLgZ4/TZi
7xBKQbZw8AEHgAECpN0sJGFpxg7IMTXmTnYn/1cap3P8kuPfU3RyzCgAnlDzf4n5
8v8wKjglbw+YEHxnrjFRRf1TnH9ltW9hl0C10jCax0GiPUkA53HHe0KkbN8x/Z7W
WjmBF130qH6gPXRuid8V2ndaphk5Z94Eigjh4wCl2Fb8BvfaaOHQg/BLD6EpeIYZ
NEmw4gTSpMKFUljhWtNYH6vhRgzL4JHvmGqIUF2dEq5NFIERLKGsxorwLTWIxCuh
mvRsfawX9z3wE+mzh1GA/vd1MJjNUqDGhO2+N0NSsnvI5sICAVjzCagWIX7AEd7N
RUf6kEVYFuKhLgKbg+mUC4sSNssI9ULqV2daNyo6qSHrixKjGIE9ZlOPapjLy0oz
tqe4cOJl1RW9FnUHX3z6XgjVj3dn15fDBxOYwVK2Rm1PcKlBgFpIUOvTJjkJmASj
UNgboZWQiLSA4PdRfHVgwD0wKGmciKbOCRnf4o/dGHCHlQwBd7iNSHnXLlBAUg72
Z1rfUwrlD9WiB5iZae957s/pRig66egK5YS7Z1buy0GaGuxCMDbInW2nLsZcn+IT
W3k9RP6V28rB0V9q0biRueN7jZ7skjryqPTKzSVH1UTp1ZczhP7gmlJ4PmL/tTNE
Fn3NX6Ap9YKoEn2cme6fhWHfV0NdEDnDQmxErcmSsMVANmr8n9fJRrlFKOw8OKs3
0YEH5av5Ql1hiB3FiWNijzhIrG1eTUScIVs2J/HziM4ewVKlFWt5Rkh5UW5RDfhK
erQK7lxO82gZdjoZw2uvEW28GhVvvK5RUhw+BSYt1J4elv6sMT0WIMmPTq7Ud7ai
jd0793/7hYX1KpUPnnIdXuOf4SvjqNiVnFjNP6s3eW+KSozih+meNagplq8i6EPD
FFSyktvJLJj0VnSY5PH0eW4tclMAW9Z3uFY6bCUz3BlVEZ1dXOEaWIP9Ul7N17hl
EzU06Q//e3Qb5UGE9XhAp1fEtJkAAjA0oJmQWOhEXZjg/7zJwWNQFY1ExTpzYcnG
hRalK4srwGFldX4ZWMDXcXh/XDbgjbXd1DcASUIy10A9jjGbrOMXith03d7WA1Rg
itUpdrLNijKZuzoPMXGeOsUHYpNwX/uIEz0vpuEBFdzWAN+Gzj/uTzvGNtfeq36F
7L0J5AWPJeNl+QmgQlTl8WG0iTm9MFBSbdWcthWTmjE1qxmweqPmLYy9+NsP2kRY
jp+CNbaS46LOxpEpawiMzGfvwa1neRjs8ME3320YV7Xcs9/74wUSFllqhe1uQgYC
/gES5K4VgadW8yN0YDFUsqbqYrVx+cOwacWzv+w8HUiumjR8Y860pCpxlhtkdjRj
2X6eV0zW1BH/lcUj+VJjXYz+Ddh+DWaaszoKS6SlZTiUqrp0tqW3QGQU21WKyg6O
zIHXG59XK1CUIMCTMkb70YCqz8uMf77nxqE7ijadbrujBaLWMoeBxkBfNwcD872+
EuWsxqr6KT4Z4YW2xSUmtueCGy6yk3iUHsnrBrXLqmCUFLxeJNN+yPDpXzudj4+Q
FxFZJ904cfm89vmlXdmzFZCmV0/p0IkpsWEntGpyqD/ufhdtWYshOsAkj9HhD4yo
E9DpYSR9JeVUSq1F8RSlKOMgxGA+yyRFSiCcobTYrz661u+fTme+XAFUGRhtlKpj
NlUepQdwZuyGRi8vnJy6x3j2AcUj/yW8f7bCa/eibQg3A8DkI4OKuKdY93dXJWU6
rJRKLzjsnNM+9T+qOoObLZJyyMZ7fGncMTg+vT0inyaj4ENVhrJ7y+pwYGIFbsTT
a6figcx9fUXVBO8qzwgBImlbOPNdksOq2udjQDh/NMBTYPrpAZmk0Njvkeh/uH0D
fivYKGnQxg3/0u7NJaZaE0uAtPpM2hFJkJUqeo53If8JIcpathOEDsMn0bk6tlIL
+tmZyvMDbqHmBRy94x+dz+c9+MMiD/WGqcOm+bj/BJ5XaKzWfVtWWYsS6OQyoyeb
Ko8gvzUYiekegUsUC21zi98wt+LTe0pkY/4JE2sbkVuDVbu0ni0Q2WFtMihgQoSe
/S6bKdDrPMMZlwqOPiLUMZNaEbmItc65de4R51stBlBXdrqHImekjhMt+1x5t55W
HfFaaWrr2w/8IW7VAPyhmWR3TYqtv+ohRl7xOXGsAgkuH3mX8lbI7UEKDeRSJZNh
5mwl76Sy2Qo5XJrBvenN/MmuwVfFDGtr9g0CIKE00skLBxo3WOkqacaWfL5Dapi1
vtv5LdDpOOA19UcZHa6/RG6EuR5JGRQtRt0MVzizyququGpPhpa3JYm+yEZDuJmN
I82nnpBe0C25GlC8Z1cvNAWecLYA9l/FPPJz7r8mK43LT+dUtgnphEyH9aoLfwdM
EU0DWpPbNYrel7Vi78fhuYpobVoShTRszOdNDAXyLMDMRqMMNtRrDYEx/s6FE2yf
Y+WMBjoSxbiPhbF1lh6OvR4ZrWZhubFg2BA9h6U2vj2Z79UhjlWxim/0ZGf4qyQx
A3cE6NiTHh1JuVg+U0eq9x3KR2R3A0WP6EOhogPZ4oYyoALNNBeOiNy13S5wGvH8
eT3Ha99Va0NlLk0G7deKs2OMfeTjQkT4V8kll+XOvqPUuVE1fz/dvd5TsJ9Jf84u
6kFBW3WswOJyk1mcmMTQh0ycNG1OKGd/0O05DssgT/GkQLTc/iHaiuktzGR9o/Wc
AiBeoev82SAykdkIU9lTTJry4PcnRErp2cT3McCgU2RasewfJw4Hmd9wC0ELg5Oi
eRzYG7i+dF4g9UMsxC1THL3yUO9EbfTyLE0LzRkEptv4KPGm2vB4bkKsaP3ZXti/
nLzfbdf/9cmzHCydVR4iGzSYgFsIqhKiTs2sI14NztH7t4xZi4rrHL2t7uI7+xxZ
+d5JpNlbC0MFL7DUtoelQhpGQmvlPEZ41Q4aHQ/aZ/rJXQS2lA56K0H+wQucXdoZ
zR2Cq+xUr+SFpuroWykKFnsvRD7dghEUrSZDbE4S304T4rSmOlmV/stQ6Hwv+V/G
nbxgF3aChm5aJzWpvRZVwlVC4DnqGLMZU5CNJQR3z/3Vqrrs9evF9kxYfNyP/yj3
CLbi5gf4KXlXP8AbwWx70Upvw3cFDAmIiyDCQE4VJVrCTIQqLXUrjmRc/GNrcFwo
7v2FapOOiPdh+f0Dulh8dpxh7uuLkQ0yQs+rTJUsXmhcsXMvD1EbON0nux57a2E5
YZEIrTK+oReBonMCqge6t+sAXN+tWLRCjHGruR5WJV1DCaCplQfuEpM6QuQW+6QI
iOmDsuwanV0XhcEHCatMx9SBarR153S1Mpa9z7BOYzH4vqm27bEj2kfxrFBJ/xni
USfJJONGh0TNWhNsxAZPlc/hJfa/JgFYbCv1FlHoZQ+D65Q3ydmOhOfmuJdU5y0P
bE9xV6nGDAn89WS+71pe3cmIREaffk5IyptNkh7pHCIhWharTLZ/RAtAzN1/XRqX
wefNoTIETiqQdblH0qtRJB7W0qvJEmySGI9gdMUpkbgLtFuQQY+5EzZdn2+RQIFR
N5f1+guPy+TtPKEEJfkgz6HMZIZG2NtqFZhaamtP2TPnwHmoFvjuqe4G8LojEktj
kHwoAuZmT3YyVz5rKzqJpbwAF85ecbGgpeM2PIT/7gD9bi9vrAsbujgC7DWKxw3b
knI1uE3AxKL/y5V+fNGXCfH4uiTmgbiyG5QNMVDN1Ed95clKjROmtC3W9qYAjJmp
319wZ93tYo3xVlGrdPsyATUunXbwuKJY+8p6lz4JLUPeMx5qUfx4ronwucFPh1ny
MFTwlZoTBnNSnhHTTEqI4f53LyEXNzqo5lUENwc8uf7jdzbQ4Gf7ZD3dRJeNQcG6
AQdnRRTQxxIfUeIoUV5SL0NjGpqebDetTS1Qxq97ghko/HIQpvgVMMBUluxO0nv0
XQlxiuo5aGUEjtWoEHqVj4z9Sz6mJzK65PLDYr5yhZjWKEQbB8VWpXIhRZzZQbDg
4rJClS4VmE3KYJTKlp+/3SYvMGCMXqzyaDXdIgJiB9jk0VZUyzqM2JCtDOlZ6rw5
d2AQ28D5iO6VkyF5AAuDg1o2ktRzG9bazj6jhcFOAt5c7ik6N5SFYZ2vDCsB7TGs
i+dcQTuXFP9sYtRgDSAflbyirkuh6TRfompYiMepExDD8vU+d5Wa9Xcdx801vuf5
Bb38r4WMOkpilRB/dkrkJd0m7UaA4lweaM1SRg1L2SPJJh1UpEhiTw+NfSjeCtxo
XR4C9W9U2YJ74H7SOXvcHCxX8tr7lGob6C+l75E3UkWmc/4K67TN0vj2/Lkd8vGl
VZZwnS+nDqPPxFXm0NUN/Ci4ZqieS5xmS1zBPbGicF+KkOLMW7OEQ5tSXJnAn3s4
1jJSq3tQSlRmhp/RM1Hf/ONAoTRz6+jJuhErr1s4l9NsGVzylG9BEfHlj/puZHIN
x7Yb5e9wtvVTitlLmDoCeV7+VkcWi/E6qZSQ9f1CI1hLW4M7To29hQKBp76CB85L
U8Tub7q9Y0tbKdp4DUx8uZhmWQg6sxHA4y9lNKik1ZrgKAt5tVmPWoZxqY1qbool
HOsVZMhIDu6EwqCGQhAnawmTthmv1DY1QH5YSWJZxmG6SWAwLMQ8ScKheFlSxk3M
Dna8rOb0dRHP15g5LpLQAoP5VmJuxfmBV8JukT3qK3ntIG6952OaGHFRA1dLe5Do
JFx8TN33sOve7a7QYtnxcTFr/jM0oe3svLqk0U/IYfcx7qzPS3n36KbrWPqMvJk7
ybtH3x68KmgxF7a6E4HHR4o9m5+puM51ZCqxcuOqGV3ftZ321ofxhogCOTBDi9QL
em3RoddhYS9b6hycpT5NAFiVR5RCDpT6swuN3qDe9BzS5ernYSMmqY+uxz9t9YZ2
347+Tku0E8g6MHcOouJmGA7M1GTxKDRsYmnZHzXLSpx06mhOsiDXGKWpMz5lKfdw
lBxzluVUSHpgSld8ti+VOnP/AtCu/RZkPHQ/T/Jv3Kr2YVAZ327RPC7mmsAHPHT0
/SF8SL25Az6X0VJylm6bjkUJazPV55dB6wgfdCzREsd9p/E/CFpv5LpdCJB8HhPa
x5ojhTY8poi3Jg9naFeEaSLEms01WCLzD0UW0GXZBAVejNDcV3QjVTeHVJsgGNB7
GXL7WcPawvzyV/nRHNfDB4C12a8BsJtCmUOn3k3RANcyVHJZeE4olIjw6oFZS/b8
iB1L46rqAcH7MvLsPNVx56j6XLXajaLxBIx1DygoeYIQd2HSTUCWrUljybuzxepf
tquzvEIxtqlb9mRE9no8hCJrKQPHccD/6sc9KxzY0syq2A4CbCb2nA1PKyEBJROJ
d3naW5Rwhvs2K2uD/9OaZVHlagF8jlXURgoFp7wTrc1JH/NyQF2ShHiU5LenRRfY
fOcovXVR2kUeZfA7bvZFNhNpQgplHFtfh1Oy1AiYbxSuz7sk1uWUTzvo+zxtPE58
28Tk2pEls+W8A+Hl8cf3YeRsWRGT1TbrFAdd84A14xurTcK5kRsk3x9yza0tnf6G
cYB5km/SbamQHwewKfavnt7vyu52fsjMW4n8qRVAB0gN91koNiJVz7UjiuDLk/yO
8hRfWiU/1syTaC3LXwg3nhJ0a8ZBmrZ7FC3K6bkUDvibqJ75C1/dKLD+z7semhjp
aMzS6pnJHeO0gxF3k1iYBjbyGeOpQR0tYwyo9VVcb8LiS8NuoNhPhYb7fBHMCM2H
tv69q/DZs8Ko+hgr2JSWYDPm7x7P/EAg5cd6l9PJ/z1aG2lnPOCPCswuyJXJ8WVU
KYtWQFCMOsKC9aNsVvU295NrI1YQxDcI79qcadNhAQa6lXbmOOwWcJ1AVhR8mp8f
G0Yt09WFKDD+VUOLVIytqtg+L+y1+VXuFfiVZX1XxlsR8Jap1TxLTy8iZ7LHWMSO
z3xMuOYwtg+YSEgICNKTGaxImLhsOHMl6IZoAqjdq5eEvoisr7vHhOjeFZoRqr3V
rVZpYUOl4zUdxZzsOV5Im98nUjMyoO6GhmHLSdtLnYcrzcwM/g8iGfgS8rcWsWjK
lTb/AiMhfl+7B30umt5T6LaNKI/pxPVoN6moxIRU/JPUrREpj7CRwJtLgtNKUzMA
va70jbhQWhUwtp2Wj+8MFqhyp0rRF/gqF4NRlUi056b9WlqvFxS++ASHj1NtZLVk
dUYjyxLvrJlNsXuEMrZb0JBhwueihsyG/ws/bYRB3n79Pu83M+pffNsbWTp0zfMj
o+VSA8o9bvsJI5bh7f5SH1fW1FvCYpa6qFzEEfjiRcF1V5hiOIrLkkHCe2+CSZXo
g9+s6e6bhtWb7c3SZBH1dRlstlenFjvO/4QrRgZIwXkCY7rCdAbTiunS6p8LEOMd
SPQa20D8DOs8cvLjl7hSnWwK83Ix+bbJLqhIw6x+mKFdsH1qU4Xsg4E6CoHhsAgb
xXCjm/CGmx1oX5XkahVNVoDV6666yJweEJC4kM8feEaM8pqNQsZ+h+AuVAJNAClQ
+080C20Q4mi8et+4zD+njmpslqahaO8MKUTG2b8Xcxy+NCXdaFaNLg+HqVkPTGKU
61RqtB4Y6CuNj0lf4cP846rCimYXjj31GxZUoSfOQ2+DGc9XKb3zbpKpnfvIo09y
jNGvNnN7bL8zXiOYARcIEnl+axq6DqnzDrOIsza8jQgS96YTzw+hyCkMgEU6Mchp
Cr6MBzF8SQS1beA/V6ekNVf52fXYt/+QkhZjHU+qUedXe21REWSAVfBAL38TSKi9
3tngV00DLOoVcGhFBu0bmcHWir+yFjK09WP43HBO4j9bLDPpRAL6Yo3VjSKDvira
UiGBPjeFaUfBYGpCRu8k2QGtdQRAiW9T1sS/5hxy3FAnE9XGzY703kFR4PqWbW9n
TQ/2GbXb/ODFVKkFgsjkR4M8MFIF4praFKDFsaUGCoTzINfMr/qFlmOdTvLwOuHq
PGWxASjhaxrdxDQnKHKmybUc36IR6DlRcjBvnQsbvR0DOy4CQa8eQhXY+/9MVSeE
BR9mBE8iLqaqd/UUeoz7wS/20UUuEw/LYrr1Iya1dab1JkhqX7ALcnJeZY+ivlp8
o2DGFae6peM+rUAWsDort+F/Mq9Dc4wL3MKNU7MNrBSj17MUyICm7QHDWKEh4teK
dxAZ2HR0ivATASJ/W6NYeZWVsxrk5T8bGejDNCF8zlWZKC8xhoAJdbEwyoiOzbs5
T0j6bVQFZnHlb/u5YzWgiFS4SNkvlqOIkyJhVYCUmBpgKn6MN8cLnKw3pyvs2Nwx
WcgnTQcat6zgvipqgN1gmFso13V4hY0HlHakJxYH15NrgLE6Gwm7k0krIp0goV4i
YAcnJP7S+BdJxcuQKhQIs/GU/eO4szgACd1rqtAMQLaKvi88oROXPLa/FjHx0yil
bpLO/OVvhTRVn4/d1YmgDjdEoKe3qPqKnmdkOw28DcPXFK7ZwFtnH2YawzY2jBd1
d9precHUstBZezzs6lnugFcYAKhAyppfrkiMJyEyOfmUQWlwGobCJ2b8TD8H7S66
/5LFNQQ4J9ygWde36VCzRBXrWrZFdM/sgq6HgCVjdS+M5Vk+dXbA5/Jl635HT9Er
ACKXmzceREoXhd1pgK1UkqD9GgVaSRIvAAQNQ5EumG7tgX/lpRs7YXMFhpOm4JzX
SNwxl6GqKJotHtkwJENEE1spAEAQFwBSJbMMpAaPjYgiW+4/WE/O8KPaB8uOVX2h
sjKgHm5HxHSBVEvkAmHGniU2ts08sgcUYCpFKZN2OnyfBXZevMHNBlVSUuBppm3U
RI8HPHwdlJmJVvkqOrOqh+XQhyLNB8F9ZuHsow/YFBjzN+/BD3Cq7UwTzuxoFduw
z2mt7YKpy3/jj+STsercVLQ5zWpw22awFyT8yvrjFQEe4dkP9dVl4g2ApRYRj9EI
tFHBd3j7GJh55u8bWr+Xll7nuBFwk1agdWPLdDHoCYSZqiod+M7Tg3KyebQwzuTN
4a3qxPzA5yM3AhAAKFwZztTtvUyoIGzw/QrA4qPDFBMtgd/LPoEnMvb45H7gqLBm
kLIuIyqHohwbyB8sgnfPn89EI7Y2qmImHTzI3KoqH+bYNf8NNXBZlzoY2neAk98U
Pml2NUPYY+kAnJHmk/1xb7KtSas4tMvDic19Zoez0T+XpA9vEDSg2WsI1A4Y1aDx
lCgZZZB2QxL2/3qA5/hWpR+Kj4cLi9bZ4r4zbq+MaEGnYIpfhdt/4RHLPIi1W+ro
JkTPwpkFSusoRnc1ARZLX6SYdG0B/bD5Z8ODFeDuGrwd1ooAv+kV9o36LjChlaDj
cyEHKzTY470MQkB10ViRwpHBZuwoOT1ArSNWNMbf9wS1fWvt55esdYpMStaHxOte
b/mx17/f00/kl3ye+u7FB1qWiTxNwFXSa3ADRA4Grn3s6hTSOObTuIluABvY5sGB
IzeRYTPtd5RcncxmP+lWvLehCDTvcyrVhJcdCKCSy8+qH/3gAmYFRAaje0ooA3qn
E6Sy/yn9e61HuwroP6JXTMO7c3nJyaqy490TxYbI7jKCxN9eC/e7pIXzf2jlBv0e
KY5k8ORqFpeZWyl7g2JIvbhVVvlFU1HYriCquz79vmunHJquYGSqx+OvznbkOeFN
3j+uPMXQenmvlzqft89aEZgIzWktT2Dm4hHhq4TkURVVnN++c60M1pxJjfyHBpti
LWTVJ5wKipFP+U/L0wAi+HT3mgH16nTkanjO4Tev8OVJ+9CJWqQdIjkwygbRZo6K
2uN2yzmKVsL+owU8M70Fj0ZJXoYl9X4OPYJTFJ5h8vVWyZ0G/7PzqitaVZwbChrs
ULJL42O5bhEU7Nw2l8Xi6JB7CMBLOZ1Ax64aITy5b32glH1gNNcDnxqKH8bhQ+KX
ZtJu2H+B8FSx31RhT/srFSdcohRQszMTX7um3Cwr8tLE1ndAaFofyNG0X91LoCpc
kPfeDyGVM/Wm2exkB/s7kITTp9Pa0qlR2NHnvNowpU19hy5LpM3p7cVeTiQ7/eNQ
no4DQM50eQsLmAyEad1PzLZayZidf/ft5H0iKVj2F6N1Izxb5mvmPR4xmbV/inXQ
ZL1t1bMp13c6folP+sSCvc7a5KvrFjhssguBHfvmBhw5Nc8KoogUmEuHFhSXZrsH
5ow5Qxp1lR5zaQ/77FAlWl3kXupDv2FieDfXiAUcdfAMVe93Yot320D8hpcFz61T
MR5D2ri9kxYFq94BxjBwJRvWFFmoaHeeCJ/hKf1KPUX+hEB4cZKO4W9+3ySqiEUz
7mg4Sr7nlM46dBDlQsZxCXYB5kIt9tcc3U5FhwZQTOw6Hks9RA3zwZ8j5k/FrFQd
zBHwt6JYCZ0SALcfvtRcF1l6X8shTrN6vmYkZDgqskH+xCa/57lsFGAEOCO8cSCw
S1SoUfnRydCAxtVTqNhGIFvrjs8jRP+t7EI99MQxs9MPVIl+geO1wOp3ZizbEdkj
vO5enZv96b++VbsXyGfzxsF9cKJBL5m+Xc9ZsOXrSuOM1bI1GNO4T438WjVgrBr7
ZnDuHLW4Vmm7SCtu7Xgi7rP6yNYtntekFMYO6HxhwyvXSeyyqlImxWS9qL6M+zRp
XiJaz56oDxp6B0NTaEqH1cTCB2svg1JCmt7yScZ0ckcY+PdqRBxIAeRWMWGR52hH
gh4hRgZPzYuojyJJPAqYkvXr/MgLiN8swFiNuN4ymck1IJ9ut5BmzjzGW+WFcTWZ
IuvzWoAvkW2KGjTA6h/sNIUp0hqCQksajI10akM75DCwEl3PKfjWh7VL6Uri4wrE
Ad19KGBTvZT6AFc6j/OegUrPPx5FpOX0/RT1VjjPQPBlwmVqfjkn8sB0WPXzwGFY
pTBvaXntNI8r/ldAl8sgxGswZqxLbzeNRmaF1FsMrvay7FraB8fzUV82j/SCg6I6
eNjj+Vykh4SoswyCWWP19+Ziew8r8CqXs9iQaE8vq76/XfQvLuL8wHVTwFF5FzOd
IaMsibO2Jwuzmb2QlPhpaSiK9NGy0YKuQUZwyKKn4aEjv2JNxBxrbzrXtEyTi2e7
/V7+ES1UxkFUl9kQGnTQkxyzzfnuNkoeoEjlh3Dw9l4+tAgAIrgCbo/4EoZbxGq6
4fIPJIO121I09qS26QrsnW9MT+IDHhnA3CGMNTUei/i4QBBvEJtZSYEmcYdvucD5
HQtzl0lAEuFEIcsCkWlqaUXm5QuMrmjWcl2T1hN0/NpCky7Nsp3Ee26REHXh47Kg
wuberNmtiqk73Lfh8nO4oNYyH5YNzeQBAUd8E/Vl7GGsLgeOz71MyFz5K4mhlcT6
zMUvHgD3x7yFP+45OiyibJKrv4X0+m9cGcsBFE8myZhGAjYTtFSfR86MgtIcJFka
qzctT0DtTl8Hlcr2dE/ypA2zglWsmYXTtiUVKjHbGPAqFYP5INI55wW6mweHNqgy
l4akDSRSTJ89nSHV86xCQOTUSCw/UDVyFxko1VENm909e1qBUvIsHWHsxVCi+bKt
k0RrK/hBG7lhLheXqJtXs0AFATz3zF+iCsqUssnCc9o/v5rjk1AQeJBwVZD+DEx6
N1WpoBSakBtb4biv+fHmPV5tuQ6/d0cMuhELbqBQ7f3C5poYRyx8QqL7tIfnQaIi
lclzwjOK1d/6PSO5UsZHUpYIMYRyBgvH32VhFne//hVEZBUW7q+BCK4lMC6QWjuK
SpZ7Q6VQW4jxZWimBv2xjNfzmr82kC0MuGogfKEEtj7D8dT0RPINcqg2mU4ebkm6
4a6MBLtpdsgaAyQZx8FJbz4/iCLm2HhA7Gp3Kh6n4gEfLDptklfk7fwfiJpBonnh
Z72FATDUl1PXXhStS7zU4zrtgxfOTIWn4K5qM5WY9wqFUwtUcc7iNss0339oTybX
9uQFms6EDP4uvxQ/BUJVbMjBghfDEdFfZnpTC8LU4SH7DQcMIXutrlSdMlxHWahN
aB3pCFn48ntbQSjq2NaKRrzggT3UBDDHjitI9BYWhN5/mSai9YLJIz5q7VkvrEuA
tvSwZs4oPpRUpnMMX+xE5cP6+Q9Skd6n+spIZWtX5DuKxI52a+DyBD+Po1EZz+p5
XN7tApdd2wft5aHEVgMdATHe1KvqPYDqxI0vyTU8R5rl3DciYFlhrLVAghN3Fedy
5PLIuD0IY+yL3bU6+LpBUaYF4OcWztfgrGkdBp6ksGhesCvTtglYM4+KKuM8lEPO
FB0/WuDV7d82SqT6oKqG+lC7hC6xrTs+vmmrNDnHvqiWogRLBRfJshgb0IwGbh0K
45YVMMlbkGZV4LmSdEyW1DJCN2CrIJTg+8sVjze66glCpcUwN8UqNU69ZOcnH4k5
daH8SnY6fwBlGqg0c7xKt7KBB9NvOjuZ9ToWsUFnp2hiq6aJGu5gYFu398BR+KKj
AoUihykPg0+PBcw57udPoBAA7H7J9eQFXRJhcDL4B4ANBGHMcth9LZVs0Fsouigh
CeI5If6RAdPodXAkVRfZk0fo8T8c5FgwMSQ/UD4SyE3hGgRsXNXimnjwS/h/V/yb
8ueu0z1JXebK1uNC1O/4oysDyoxWgj/rXJhbWAgfQh1XKREsyOzGx79yDAnePseq
QS17jH4TlacDcsIgvPWcf804Dms2hRnshwcsKoV1kmucB7rMGAdb+kjM/gJ5QHNd
WhtB4IPFzjzuDb5BNacWXJRSb8qvyIRMKtY3Swy7wpCmJ7zuFrqLSsCn2r+slZ/K
keqpTy5lIe9aqW/JyjLk3xtEdirxRxyk5eSv5H9qR/2J1GbhB7Xo/wga4GucgdRJ
Qfci8AYcWEhHUyOy05swuHxsiRZ3dcEO9kshZw4i6QtSaVH20iUvQiAsuH7dpRnI
2R7HRnEomDnOReuq46d5ARHVauhTxiiZMDAs0g8KoaV/1J+iO7XQW03IjFMAfpE3
WCOZIVHcPFrT95ELw8ZRBTE0AEl/eBmQpghbprqtIknV0V12JnrIi+/syU53xaMf
ZeskXbwBevVr7ExA0Xhh/NfaD4OI0xdAGoDcnCjCtKrMp2saUSpSHXiMAU4gzsgF
zy4nTjjLKusdCH3Wex4Rrd1p3khFQnKZJ/S3/3ebDrqRQFkcsBknPcdUxLuGXFgL
6BfVFc18GmTiF+CcLOY2MjL2k2A2wgO3jZR/POdhuy7VIEZYYj4s2ahMSalOAORF
A7EKoWqagvMxsd5Zj2rw8gwkcWSyp54sih1DLsaQXg7BxmUqa7OYekpfNMI6d825
R98EFyRDljAuqsHFlaRN9rTqayA50yBW6/wzfxyEHuiGSr/zaYtkdTjkEKXxCm95
lq80sZ0lNvpPh5feByvRsshhRqlQy1Iujk4g8AfUXlUBLYd02ta0ujv/P5cnLtHs
ctomvO/pIcjJQqkOSGxzqEZXADdnq6GGwjvF7sQ6UKK56zuZi8eeTuYNE4JZkmI3
xkFyTwIXeMs6RziXGEezav5HYX4syiSsNgQlQGAKIW1/lCLGwzIHflBFCmWG4rXC
Q++UWEkCqZwGqvJFhyCkpCbucl2wMh4orrBB5Hlo+MMgeyWQcisu7LPpj6Avq8LS
ypWyqFAzT2zSSaFBIP1aSVWljEjhaFtQyH/PEOEXUbV7ndnlJrvRNijvtewvoOpd
63Bq0amEn9kmlwrv5bbA60t+rkIuAHqUp/BK/Y8TtNuLKveT5KN2h6tRlv5X2Wc9
Qbo9vyiU+JIzRBMYKbEsDtea8QKHakXTiUn6apIKNnOGRWuGudHQYrWpPq0zKrNd
Eh+eB4O/vGmHl/HTXWY2vRBKVFq6pkRszt3b/Jevju44h+giShKSyLMJi+KRnDzz
39eMECJkvV7LLih1Q2HWg5w8xO4O8T1ATuX9gRwU8RznhWNZ3ArVbM5RHcZ3WWAX
UIkr9/1Gd7Tkx0QFRC3p8ZUAQB4Fn6VowSzZIBHUklJbO6Pq+91kLXN+iFQTrR2h
BctHPq10+bIKDbVKJjsUfymb33Q6jdNeJVkJiGmcM+edZ9RBX5/mQz4vVdhxaoLF
53wBSFsJWSCF42Au8ThoQsL+ZxeDU/YkMuDQ6jIrO6vTRabFqJgdKg0OFUZfFR8d
68QdjbHPbn3X5Vhgz0KLKEvra8YEAovx3GgUp78pDurTjEFWxA2EiZJbzHJ5mYCx
DspJYoDW0YHhBbTL4Uypp3W+B41giEe7Pf2AhpCI8SK0waN+kGhQJyIdzq8u/kt/
tVPZANzRMSRw1k+zSul66DD4pTq6Z/6+LOrGckRRo1CRBM7mfIVyw5koYzFNK3Fi
8r+olq2kNAWeYG+NSGY/0W7L4YTtT3039YfFg/RwlFzhVzKc0Bg4eMqW20WKL176
vDN1++AtiJA+rH7tEAjoV81FpHQeZUGUDce6TggOCSjWEQU7bXQpZy1dGwXYTIxB
ol/HC0IqA8ggGscagODgOix8z5NUToyAH6rUgbM4YfQGj999hFT3BW4bnOPRuZSx
QXY06UXNXVXo7dSDBtix9933YqQ/WWJD7Nl37K/ovXwBhMpNfaOZK4x941u7Us/K
rk+W86aG6HCBPETDFIR7RLuP//LUlGqCjqAavJHPTCpOV6bt/kRqcZokXqneC5L9
vVq72J8srS8xG4jd7qTC6WPeFHpeetnmTZQenJfU2l0+aZ3Dq0nw6TT08Pdzp4oF
svK38axK2ETU4x96/2qQAxYXOwdVIaLGIsaVLz/x0TQZCKliDdTC1v9az7NP92Kf
UEVvDO18fgt1jtTZ5o/9SY05GespK7cfqLzj7VE4o4GSAo1g/E5vlnXq6zTNqP+O
1nQkuZvE41wwfuuDsEThXOncKSYNy/WyHAN7MFYolw3eFcYPz9eNr/1EaM3ZkRsg
cpQ/xgkURQP89a8994YW+Lov/fMai9BH+YeDTsUVjeB6ccidK9T995nm9dBo9aEn
mSVS/RQKGXDpuHo5ubswFQHM3oEPsBRPtk2vyeMWdIc4BVEIsbN+Afxjg7I3Oigb
X6VdYggDQ0sM9lTmi3I3C7XgtFLeImhDy6DbHpB5iNC56qvNCIlCUUgOcNDrbI6C
2qa2aZefxMtMSWgcUTZCeuEHTBFbkTN1JCXJB3oRhiyL3ym49iyqoTs+ayzZtDY2
nEEhBOVat/p3tubM9sh2y1Ea90TJXbScS/R3aK4eFxYeodf29f1caFUKF9MtxNzb
gkmWLKS+1NfumPdQhRzf+SDKfE2lKfE2MhpOx/hge5FLStb7/Qc/pFwHnm3/5uly
ueUVKSi9HAFJTQdB41QpXZQrSEsZfEwpi2PucfV417pww+XttHKk/KsHLSjmsQa9
X/7AFlLpmkYhMijeV1XMr00dmdQxfzjCPmOmeF+zaZIIfFHYuDmsESLI1bj/ErV9
38ZiEROB8E94wGLOeAOtisCPNc7lewVDKzLuc3oFuAHqb44U0MOxpO4X7gyeWv2o
jS2PGp65EUDUAQKT67h2VQjImiUQ5XEgpC4VrP4RB8W7oTSdcnWQY6xbuBOC6lFA
Ko5Bns49V4UBk/TT4cQZUk1oMMlvJpTyD3Qxs0Jm7xBQBX7cz4NU7HBZzW89wsXG
hXDb322YQPrFA6VmzQBh/CpKde8x4k1X5LpQ6NzaoN4AmM5KtYw8eVH1ZGcAGwz2
TjPa+Up7Jf4ar7vGaclMk8/+3iBiIb/DbFVj0U5x7CfikeQ0bcTwzyOK31XLBdNb
AbSUUUccQZx3gkv12fn5RSdLKG+q7EJYWzVwVN9tLVUXQ3DbAis0aX3eHcaoV1n5
x6TncZWe2pkR/6E4mc37A7oNWI+HOl6l2Pex+KQ1hq4QZLQCgprZYq2lV4ZFWXoO
P5BmPwLz6OjfuoFgdyMvcE3IqmdmJisLD9zUrnRbLWKiTf3A0DDUJ7ozG2UALgyt
qm++A2vzZJDX8LFQANCqFJy1A94drmANCN2V4yCsOB9+qLBlh3P8AoYCMgSJVra0
JsfTpyNAQFyiQI2n1mFTT6lII6+tMfpbSC/RjAO4Sv3EUklWxq1sD9IdIHm96T9h
HIU0iRoTYzhMSxHZonzMzyrlGgB1492gHMW5/yHuacQUe3DxdzE6BQUsvTO6oRvA
MMmwUXcLQhllpOP8sporBq+sUl8YrdrNooJthzdwaBxwQk4SwYLguKEHPvmpt9iX
YbqzrbnckVR65mEJh2NSZx76m814tSJEnQniS1tLU6FnKRsUXK9Er0nrgUvKeuKk
aR9nTLUiXN7lj6y+/4ExWhJK4XR/u+STnVqL2q4paP7Mg+ngxaeY8gs2uoCIBh6r
D6VpFSgvM9wAsxWMIamXEGn3jVS7GHcmJ8Ad5asbVCdXy/dpvLG3k2UalLiq8crR
820rSSKKIc7pjFji82bW2KPyYq0a03xYIgevjTB/W3so+/zv7w3M5uMhV2O4JOpU
DhjZQY/x+0YrMtIveyik8leIH4hrLr6SeME3neaixmC6U/T+Su+Dm5hiDc55Qw2L
WZuWa9mDu06JRjQJxrQftLKV7lC5F0FQ+DEOSSI1rBfo/VJGb4f/pJ9xk8J+dhEf
8VfHXNfcItRUShj1FCG4/KE2dWDqGHSYgFQNWBrVCwandpDFQn9VGEtl9kydRQ8u
ef+3KBeX9OuedvnWAKrW8hHLuem9+5nD7SkF/n7OAxtJuDvAJ9/zjiM7rCCKByqw
6Qu3OFa38zSkKFf+ZGAn/gDKD5mvpgoPIwt1RCl7A+scuGn0ChenqdViMsobnGXP
Qx4Xh6xODSGjZ1WWn27jmmKm12hg9zfyHghjtA9hLCo7bL9pfv2Xcfw7quLPphHb
hRPzL8tLVsce9gWs0qXhPLEUVW3cdDsAQZTc9bUDZFbkKAKQJRER8n4yc3qwTrZQ
kbst+TVpbmYwzfrM32MxegCsoffUt1q1/ayzlCMwEXuw7qjysJmr3XrpnvTpzq+z
XwNUSPYJjTM8VvcQ0hRm8nBm3l4yOABFnpfWCehqsOLHeLeBYEqbKvSFpQTmJjJ1
SV+9TaqRL7QX41qqGC6IR0xF18xK6rlJlIXxzzuivBCifCEedNoZFBM4iZgAjCTL
xqittsybSKA/bZKlx61mKreVhELZOdCZogc2c2tiQ0upafEQUPtkKTeOlHQGVVtq
7EiHPBI9qb0LG9nxwyLzViKx2oozscMHkDSi8eYRbS9O3S63UzoWUZvMsnTkpYCF
xX/+ybkc0of1ZR6KUGNlbr8zcvaXO6GrT4KsrPa1TYgmQjZRO2zrONBGUbqZ9zQt
ZFwUbWYhcr572lznZYmMnChNokwYEK45Wm3iQa0wIQ1dbNjU1dCLFqVmFE9gi/U4
J2jqkmdJJeRwkVVtQy8IMA4uNeZOAIp/Q+Rxf+yENtO76oBeI9vYsGkbzButBe8P
6tMxe1T28W1ZOnm+OTvRLFKNlYI8lv9TLCbZDc9GU7a2pRtn7je+xObhBTmqVEb9
we+pFH+/1dnciV77pzis5TBw05jky/DdBhgk+LQhRNfmjKkX5RM3+0GjTE/+iSAY
PR4ht5i8XAURoG/uvV62KIXg3OcShK1U7vKwbpl8/mFujCvVmyHUFho6PvgrE9z7
efeGQKj6YKGv7ztEcOJX6GCCcWKjwv5SdYSyR1RhpcLT3e2AfNtuZ78jmD1fT4OM
JgYngkcGUYBbmEuFhxhzf5Sz2BkcmuWY4mufRts1RItxA5x46Csg7fqkN/ZqjjWG
3VDvmyXR9vwDJv76SlJ1Gz2fuAQx+qpTle4aCtZ5nGB5u0wsAzw51yVwl55b/1n0
hNQ4SEGaXuheR5XLRiHzFRdzhrK1u9zxk/lqT51eKduyAMvhjT5Zsesu6OZLG+MY
QTIZgyWacRmcdiSh9Ym1+rB3Jzoq1RC4fAqgCf+zyQzp/+aczKCMWeI/RQg9gzve
ne6KeSsQtE/EuKbpAeFKy2mRrT72bHd9vdHq+x2T06+hK0SuZCz4Ayu/ylv/1D9X
Fmz/Rf1aZNFlNThZqRBRgGBipYM/XwWTAuw1lLFR0If4S0n2xuKyRT2x/C542XGD
dr++UNmnyxmnwcNHDp9Eq/QYBzsavRqK82NxLK+rzQ2PhG6s1svdI7Ecg2ld2/wU
Zmevd2nQlvpHZOiJqDAbWkYOJ4IhpfdgzLGYGeC1vCmbk/DMbAQVC02PItewO6qy
BnSHIEhU9/xst0psGVO8YRjoZpdUG89Okyc9TmWX4YEOA/XNsBeKNIBxyb8jglmY
iSLeXI0LKMdHUTF/AtOghMv1hUHQWl+Y0jbjB0mVhw8YmHd/F2yW6X7YWmBa4GXl
MDKDxB2BSa9vezdZpKsExJpuMk+SeoW4jprGnzLhFomAbHL64/zcfMAbDII1fg1r
xrZQKjyNQT2J5f974PcT+vaK4Q8acaO08sWfVOIGsp3NySBMw2oWrS4dRZZ8+X4V
ydKythebtEXKeDU5YkbVolbERTSV9+9fitEWrRFlVd3LXVx18jnNpwliBCLrZfF9
fUFO97UPHaFGdl76Fk2wEG9d6XXk7sOTLy3IrlvWVGjjgP+HpiYg1N6vPs+9ZlIS
5p8uZ4bTLenDXOy5N1Q5iN+BP+KYEg0OJH73x1whgNnPI++GynMwD/zVWeEkaNwf
YFExp/w56C05r2bNb8429+DURl36/m0Vw75cNWJat+2RwjIMSM25lE7yqL4w/Xes
PEbbew7lyxngPRkgrzx0LWtCKtM8wjWPNSp5NiXkiD4sujL9FDJN/bu0jdIm+ms7
1lWk1p1gyr81nQgP157JJCKXmJHjRZ07CG0aAYnxLrzGU/4w+B7VJzTxIlZgVEPD
PPtyHI0HpF+0DpxCDh70CT2AkLSRErkGBoO3g2EOROw0PL9gNI5o2TaenT92ayqd
rvnmJb9iQsEhNMqBWoDKoIHcs+DbASvFZNn1l4yg/aPNzb2WqSqzWjgka9BzS/7f
NyOECYn9AC4Dh7CL+P16ELPcvfs7gX4BEFJOGN3Kf6WF61tppkpHyjUcGPczCptT
j0LKH6E9+hzo12OVAu9F4eluT+BLIU90wRpLdhxvROzJnYD0tBTmOpoxtANi+D4r
XsOgLS6QAZlFFEhDejPYJ+dM9YU848cQg9KCsFEthaHvZivdNBG7rwK2d6IHUXJt
8ekZTg/38EaIEX6/cT2oLdCePaAfuEYDDWYJtYft2/SZp+KX+015USMI7LOTuueK
lcGl30kWL3i5xv+s8riDeL8wDu22bQJkAeU6uti0psovem7q+Rf60bVRPakuNDLg
IersFkz839gilIxSiKM6o3/fU0RZFipeDWdLCuVnhMSiDVF9a7dbRjblTGXF5eQs
68ywK3AQhDoAvYj+ObZxKFvmXQemPhuuy/FrORm/B1Gik1+W2MAMsRYuCdMQEV6w
HARRUXzNEuw/yJbRZviAwpacSRR5xjS5cX+1cl2KGtPw9hAVBFRQ9Jf9KUId/nR+
LP55FXB7cFz6Dslb4qPUcETuywFf8rJVm335/t/W7D9BXQYjfN4JUhpzVWQlsbzs
rj9PlJkWEyqE1BgnzfWnZVyWOpHO6tsmqgTwFBsUF5FAg+RGSIm+x4yOZ3iXibF0
JuPwqrnO2aprHYoYnPsSRTi22leEhfiPjdzsGOOluZv5V2TBD8HLb19BYkSQuu27
1VpLb0BMI2m977WrNIDvD7Jg366Iiiwi/A++gx4Duu/RuJANFVI0xMx80rstgKKD
xYLHa4zjiHYtP+j28dKdbywQZL1vZJ4k1x6wBbZjHrSI6TW/oEbONUoWVAXNLpD1
ldPob1De27ds5cabGcvdo9GA2jlTY4UY9Ib6dnegJD+vwv9/FLWAfg8GDg5wROc1
7Y80e7CVrRsBySEOPKZ4zGpRPeZ1/INc2R7YPeU3cJsoYJ+4CSVzCBYxp0O2C2US
1TI5cX6l+5r8Nhv85a+ZjSHogM1ktRPQu+thA187eLZLdOwYa6gZ761+SFzooaLr
yPU4kcW/HBpeTSJYUoJJ1qU6p5Bj++F8ydwmdLEU5HQNsvyXRnl5mmrfzKa7edLR
gAgg31rhEhkbRItaGGVPBqvzJsJ2FUCY1RZP19IWxnek4w5AovlxzZHoaaYAietz
L9y/CoF69VlJKM+bp9raRxYdIWJ9qBhE9RwcRWYp7j28sfddxBfVSoSwDE7rCrwV
NwxNbFKE38LfoEc8W9Nq6Dg8OQ6w918FuOAo+RO+wiIyLgakYnw+H2w7YnA7ar4u
txfy22z5TdjwvuHV315HEQlldsVaxL/gXYjKC6nxD+aQX7xJkvB+Yhl071EnXZOp
x1r1T+6hoan7EzJ2u86EZfqsUCeZZ3rYwaySd1E8rMHEvnfxQq0eGJJwvqwI7zOh
J7kSskj+JEGlGU7evdhjcni3pspianf4r/4zTamynJbXKN7r6NkIzqRx8yVTSnZo
Fqr6EsTDgyd/Wl0hMiF1jwnlqKaEvTBDSggYhZHPe5f1LdZ2ndNqpr3VjmP3t8et
Eemgz6FGSMLYClK0P5TT2Lo0yQt7wBqL5TXg89x0kEvf+4h7dll8QBKXfVmk7uKP
kmXNjZ9vXhiG5+y55J/YMedoOGQA0dJR2q7WSFBHiose7wMZ7frhItRf8PqmBJSD
aWbVmZSRXRawkCOPLwh4dVtzYoZOpb2ySDrHTlisCDOTi4QFxqu7yR9jk55LKafL
790mAU/o41UuHZmSnqaZ3MWqRjjeUrikkMtC7t/HKiIq29l5ZKizlOlIyykG+xkV
pwOe7cUPGiSVfkvF8O6d/K56rWVOZ6zF9jIEEXi4jSDSEJfkFaSTeDOFwxZ4Ix1A
3KlUU9dHe/IAkueBzqPFERgw4AALvUgH8aEYrLVdzkPsKn4qCFLKFDqQ9c/v61HD
d/2aHhepzDlCyoxPbxr1SV89Lu4rl99qfUzZhebTzOK26hUtxcuWy6ui9lJ69U97
psHA+YwHETOQ2pGKk+K3DiI8rvhAbIREhDZP54EWlBpF1NLfFRYgEimVVuVdQjnB
Lk0w89BaDUrHKExgwCHOdgxIm0ztQm6Ev5QVUVTueuVazm2fnOq8TVHC01IyIUfo
a1Mzgb0bY0ujtynN+xM71wAsbYSmcMeQdRlN4Uw3jrCmZZMhB8wYOvWmssQqeyLy
kfAxpLZSkfc6qwJN+AnGxRtMHXmDNofBY48pprmEtZ4U05n8c1cJJ6DPYuswhw3O
WX6cx8f57+gJnH+XbFAnsmCYGBi+mKUxj0SMwsB5LPuouvQntcg4+EWn7vydR01/
bkEnGY8+EnmadBxG0rwjrqp9GtQC2gLtbUdDsg43dIBGWNTMkjQ97bO8okJlK2gx
g287+eS9yj0xdLKzjp+T1uirP0bpJ5lSnCtenD2N+VKfdCHD+RzhNn4f5t32Ssso
0wk8t9CmZupbLc9lvfopgpEnsgnO4RSYKHaiQ+7d2S7ZNwyB6qKFvu7T2Ale0qIn
prHsmsueGpmi/9fdCDy5AjZGApPwoavbC+vB5hNU+WcKwOiV31M9DzAoF2BP+Wwm
fWxeLABUuoU1EXD3OWS3T0vCGQqYT7mJ0ifbRrYxZWlZ7HRN4/5BlmU8bWhCIICC
YnmVbjbQ56GT7tz442+QdmpdDO1gGCK/T0bvd9JKXtE4gYWtc0LItmteCAbp9meO
vWp7HXwW2d1bVNzj+G9Rei6NB+FtztFDDL01bulT3I4k0lDV+F4Q/+IdGbTKk5WR
8ov8oPkDiLIpHr+EuN3kIyZ4RTva/QEOJc+irC7rv+KDNpIuvoE4gqah8JT8TpAj
hyV8QBPgZekBQpJ7im3dAMRqwt0ymg0hkXbAa/nyoebgaeoebTnhM/Ousc+Gce40
RLZeh3EfDU1V7MLPhddvCe7ayaDE7T/SaeLY+8mF6z/QNgERGfB1/aNyZ4VbtdW9
sa+0EkUIfNOHeAOL75l1hPn3x0IgrMCZaaVocokEIhQgewuG0GRf4FkwrwpPj5v8
zx0wle9ZnQtHHqWagv/Y8VJlY7wZeEFjUbmAkKsvOiO0aZVRcopkMQe35YaKxVbW
x0NGt3WmxRGtRwoi19KTfQDprLqiPQy9dJd9WIH4Mehs3axsNK8fTNwA4+DN0xeT
ImgHcmFMrVvC7778XzmIM1osxUd2yp80xkdiH7VQ1mpm43IRsO4sOGdWZWMMZgHp
N8Kgjn7/KgABK8F7oZRLkxDiM+mt69xZDRtMaHKYf6epPsXk1RIFcPnQz1Bx0LTL
nBq4NvMN5j2RLLfd1kQjJdvwauWoPyM0AVY8Ex/1NKKAvZeS6fE3TAfPU5Cir0S0
f4oNWTKu+MZSTXLaZAOuz5bxLc5E0+kHzD9ZhNvHQhyn3Tliygj5W1xOXD6xRxe1
q99vLnibk/ZZm7Jegm+gJdTaut1lJ51hQ7U3o+OogsPEMmNVibgUHiAwT/n1QNg/
CoLP+pDg77FF37hHiQahvagjMyjes3TjfM6W7rSQNIXJ9CvEEZS9GOkvQNRdk2wy
gBw9Qn0uNY3KQlyib8997692RSH9MaAr+iwdSNzGYAKMpmTKqdGQtQ43HY6scM7B
GE2dGXgvXk1q2+s17ttifQk7WE1n/Q1tY/dNiE92f8b4wi0ucb93wzQGiAVGuo8s
fXq2WrP+XIb5Phbr5CVRKLLSrrlKKo/nSddRTtXaver2vYUUhNeGWkaNy7Cb2Wno
mpSh5ThGNNkMXCRN8Lh3VABon7gCpGLInMj6If8tXEizuXgoU83sYJQCxF5xUBAX
8PmvdKXiRs9Yd7AG88Aey/a5wca1M+xJbuOY7OA042jp5+wuXitJRp2Oc75tDVcB
9tFJ6mUktGuEEjm7/zF5Bd15UTk0dZBjuGu/TKfMO4P3RkW5qvi9LcDAuw+9aJTd
PhIl2Z0PpH6INvwsakbg6kEC45XX7Kq0WRuJGU6SiA/2K904kqimEl2x2oSfORQO
VmykpFRYjOsJGd7eTgpuz1ilML9SXZqN+Cc5S2TJ37kWMAI/wxtIBaYvsZOCT1is
s0qqDhSKWSwHjp0k4PqPLDkaPWe4Nry+YAdDM5JW/XGjDuS7nEpt0Gp8bVmztOsy
/w6N46ZMeI/M2Oe/cTEsPYAiLo5Utxxiso64F86FmkG7j8kF8ReXvjwIWPNeApH/
xyaGjkq78NExYx0ekkULJcYW3odexbhxyCOZnWuiq2vRooRH0w9A0mJvE2t6xgyr
5DrD64onJfBc5ho8sMEcUoT/iFaXe6zgwpJ+A5ZvYDpLfRWrqZLISl1cke29YEEb
eBaC6deD+Hw+nzNSM6b7uBZeSDX6nn6fw8YsS8/ODLC2NE3tBfRff23Z3Ki2TMXx
bvtLVGIaKfY4Xj6Vcp5FvpySKHcMbI6ok2CAdSTb1kViPLZXEbYXxepVi7wFlH99
9o0A0l8socHU3SxC7vL37pWjozb3pa9ubC8VJCFRxHFXnfgnAHVUY3Z/zFYJjELi
tN2eXde5O7ptqaR5IUq3U2k/U8VZ1BBPG3EOwR3a1Ew5NzjSUMO+qr0h0OvSeGud
qPEBG+QamYytuKeYAddhgLPFk1yrB+R7saSTFL6Tyd0gP6REH0zQCXVfMe/ni0d1
fOZlmPQZo2pcX+r97FwKpLqOjY/GbCYRMGFLgx/wjD3OsTo6lfWQrk/57AVVhFsi
TUeq30ywTetVd1TennoTZmyaSjuNedENgjU4INvK+XDfK7x1NwpI/25ml40S7JeJ
mh4yR4psqi46gaF8ldnFz4MtRUbY0MQyY7k0IxdUa8p9pTMllQeG+pzF0R0NElWh
Bt2rP9hyyIC0oi3qDyXFM/G70CgFGSnfk2/89DUEf700nu1V/QN1x4HmoiAkMG3E
IPkHj+XEL+OEkfU+jgqzxHN1NzfJ7e1xn2TxffK3A8QX9OpwgedaUyJqKERq1kpg
eK6aWqp80qffSWJ1w4bORs9krCikmu5tEtOfEvNE8ddrgdWSIlCPgzfnjZxKcdyO
LpE/b8e0AwouwQ4qvVxzFpakmRGuAMx8hW1FPisn56HFi+eJRcdRWMHQoDJXGbOc
YqGCEmdyFJAolYXFqkz9BwzswaGOjR5p4SOuQgILY8SnyhXv3o6PD8H9XgIxhx9e
ay6/9FomtE/+y51LFl5u/9CanaS9FDdszjYhj5xzR0Nou5Jb3H2qDK0XwlsDg/Y4
PUhxy2vIs6H9pBrEweiIGJiPdeva3mvUecN9p5bkQCWA5eAK4jZt+JCtEGU19D37
O9hOo/TokG44lAcSzoj6NGuL3k2+5PFj384VvC9NEzgKM9Uu2RHVwEvouz3ZrRx4
nw0nvItZpGZXcP/jiROyN2QEZcGOrxu3IkTC/wsBh7qULiYr1wxXWGYul6oxwacp
X0gfXN8w9OxXtkoSrOg6NS6HEv0igZlSnDO7R3H5Mweu0yLrOn9G6MVBfBw6cFnS
pmi9lAh8fcmkzeBM5CUuYeL6uH56BUwxS0N0Biv8vy/7h1gPk8zZw7OFT9YLAR77
+RkQEUabrg3QWwph+imVC4EEhJt78du4IR15WFccRVbX/7RIsRot+6wj3mFQC0al
d2REMLrIk5zsc6SznsgjuDbwipOqKFrYoZTRuD2UBrLZIpeWTfYutGsN1u554y8o
4iRC7/t6upyED+vgferRNB56TALFnSJzn7dg+2wQ9GvWaU1guSQO+WEP8Y5CNSLY
pd4eneLYizox6HAHwf/pfHu5Zya8N8GVc3eZmCx7x3AVdMMZVSbliSZEPM3A/nDc
1UzyHTol0VsT1cOXc7Rj789Sd2vRGd693lvzWdcWS9sSZRhSMrgjTlJTLIUVFigE
mlWD247q7z5epCvh4R14xeStZ2s9HxjiTTn2uFUbFe4bts0QUJnUv1uo2chWugoi
cczm9DfSSO5WvPlzVpscQsLNG1ujelzb6EomB7fkmDw8ES/7GQ45xQv0X7aWxqln
U+U+zZu+cuKhAfYg3bHK9ug6x96asjfrSQvXfFGdWxTdlKk6InIagHZIx/SEB2uZ
I3l8/XSxgfOErB0RMm4VyFCFseM/0uAc/EweJI+63BxbolLkjr9rjyFBgx9nQOIW
FzhYDPhP/CPsyxkZQ8jRPpnsUH+jiAlJH8HJmqY9P7qz5lAwpJyMPy8oaJWDa2Nf
Z4Nk59zY01uwALmWDkJIfUj+EDxAHbOqWjf3COziWIsLxSKMpA6fZ1YoLlVcfAWU
icljVZ5vDojEB94O8Y03Po5ICORg9W8pHJ+/WbktKKfMgyJV+yY2ZrgkKq2f7C+w
ojjMCv5KTGdfyBVN2rKMo5RX3nkFpE7gSj55E9YcaeL9Fl/KraXkvqDGhXfBuQls
lUSnQvg38Ur7lNZzjdSnzySZOUuVUz92btkBA8n4ikbdfPOEFPuFs5OxmWcAEV0P
8xHSUpGz/JPjV6pXCmtZZVCYnrwKytBPa+l9qQGYgN8pHdNwCi3FLULXXrADeBzY
DLrFd7+ad2P08Lw7rK25bqIjOgvLbG1CzD55+VRnRV/pc9jwBfhGHbWcKmAitSxU
ed83kTdgnSU8+YygnhyUkvH5H8Bu0KatW8K75oM9MS22avtLDUKpQKmq4GMFKcal
1VwZ1luVTtPFcK+JErnGpHesyNCsWNIFYVztoZHMEbIQQjAvSDQx2KTxu/mnGq9I
UtU0CONU9QwF+HZyZUX6pQINCw02FWxBUbcJmsRIYl+666hCYR/v/cgKZWUXec9J
KTHt58haJl6BKHHoncDNLaZdt/SQ2BlmT6qpnD29Z0gejuIz8Yw/pEDUzk8TMyQn
mJYHcbb6ILk0WtXIFfgzeAFzEBlRSqYnqtKrOFMND800Qkah/Gl0t88ZmFOveh8R
xbWY2t3OpYQGrrl49RByAbD75qvTQYHlB+oADMGkm76huWj4rsMz9/baiI2G1w5Q
UB7dmtX1zq00gPRN06O/K11X6KbiTz+cPFY7zaXtldAdrh9L/TJOXcMHtBuNkWYT
BaknIPbyPxC7bkuVXjBck8pMQB8Pv/xUJWEIYqwjVq8GahuW26kEnB0XuK37xknL
SmnBLMk9l/TasylpRhzGhBHX4eHZqsWPjnolhRbWbO23nvJ276JkfmVC5WgxvzTH
fsd7bezfwx/vZAumqLeIGIAESur0kBqUm17M5Lt+AoU3Kc/92nIHpN9kfZ641ZL5
Ja3IuLY3/U1pCYoQqwMl+JbkgiolAjqprigWcarX/TzzotXfGPN0TvBqydUXSFqS
lsSuo8sjzgdqPfXjh4EVFnTwrCKFOIkbfWGNJj5UxHsezvzbSOaayPPDQxuN/1VE
fMw8+uF8pLFAowAnAifmduZazODeYf6RfmbHhhOekUJTeRFVi7EXY4bFyLgsnBIj
FOBs9q1Zji/YE+uMEKVd5akoOEoAKubdtywUVHwIt2Uhk5wy3TCQNenOs2133Uve
Vrhv5yUAF1Ny5im8E1hn1+Ycc06+XoQRentxj8Un0pCZv9H2NoNpfMzHyUKPerBU
AvUciAJQwSHJ93juT5nGdtUQWVc03SBmyvJVc2fGvvTo4zyTpY1dWcDYwP6LauLF
rWatJGUFfovGxa8WCkc1AZ5kxruG3ZSHduL7fs3q9tXDfkCxeKWBO7ikzuh5nPWQ
fYoEmU5U6fIyxz34h6p/41X3jeTDlIUnMt3QW57ZZd0bAi0N7L9Frx7/FLxpIVOH
etHnkKN3/Z9qUUYWLg3f6CeicB9v/ZB55qYkL+D7B4TF7b+PPfJ+dZoXHo90tHVh
ykUHm9Su4/zIxjiFrYhVhEF+7XAOxYpVkPHRJDS4h+Aw34RG/30LCHvbMF56KkM0
S1Hzu2mvSSBcAS9TpulrlafXkQ1jRJheNmQFnkkmuUWe3B0YVKGly1jBlm3PJNgM
ncyCj0vMMfctVIPAEr8J/aalIaZ4YrrZMVt72UH03M3v6OqMbrzpDlhFJ3ZXWYVF
XyVSK0cz4mO59sFfa/YTQc0cjAYzjAmz4Ny89YXEpX3lLPZbVu97or3/bsVMyemx
/FBVDWKiPoSnb3859ww1G+UL7Elfp5PUY8EQx0Ybsd6GSWlETN9wDLLXr+Hpp4S4
jPv6/VQzQSD0QKV2YulLsPPDQo8VexTILqdDXyrjqz8oQ7zby7WwgdbGuZSJ3NrI
LVYILPNgzCSYTPdMLo/Msk5KdpjD2+XRHbfgPSWrS4OQtvSZBtWg6u3HPZqzSndg
kyskOjplo0IR72CU/rycVUMjdLQQfeAtfg+Biq+uVm6yuyiot+sTBVRyD2T5HF2f
QpI/yqMcOYJV1rTHYxLCkpfRrq6Mws9w8mcEeLEG915BbYnviZ9jaBJtFeoMfSXE
4Gcwq1aock2Ne6hAW4FdjMr8rBlI65HbkYIjR1jNBtAp3obj6LqtHU6BCD1VLip3
EvXB9eM/S74LuKB1eqzq/kv1+z8NX37JIKO9U3u0oPSGZFvPHuHWWXIfKt74S0pl
rvw5xcwwkYWWWmspVLbsoi51pdBFzG82KoYF4osqejNwEsRMlWD8kapK3RpdNCcz
TeqJdSUKSBtcJheYbL44j8H1UYDn4ZeRi3PGQxqvdILHYJ18K8XwMiUCKnL2B/+u
S/jBy6UO4U3g5wMPoYvFhj2izFG3g0VsE3YHldloTFe9YhiOU1qXBptXxPFpt7nl
e/FkC7cKLulA1vtyZaAHSV3gMm/tRoNrw/HjKAsG8WRazGZjVhMX+ys99xEnucs+
y0qFCPlmiHjJmOFnMPy8MA9Ky2YwhCpMUGsJqxuD4xH0RT4RvSCYxf7mPPPyNIXM
dvDjjUrwXA6cxQ3UWadw2nA688cS7NqRC1PEMqoegJqRu5pIbje0S+4PxgB//0Rh
gdHxzi4CrSQ+r8GL2fOg6g4WoEW1gANbWZqKACXC4eehDniFCF01loo+yImxx6rf
7mUo++c5ytjjdvGnHC1ciY8YdC4hJ/0eJLHrlrWuSrH7WK2WXHwPavBSGyrrj0Wy
LqyqlJzjLKND3LJflg+ZQH2eiI2XotcTD619MwLGkeZLy35qa95bo9UUWBCL1w61
QrDM5XV+WVJOw4jf6vdd5/m91leZNU+6Cl8JsQY3mT7Aio6xCpT4NJWKUheGARwA
IQm9faGDfkN/OjjZAzc7AQWLBnr0mGO+QEHXSWOBHm2tjg//T5jydoa1pW6mB++L
Tt0CzTuS8JY+HBDwG2P5Mg0mmtCl78KwrXhSNEvpngprIgmhn9fkY8bkMmaAltCl
6he/f5dXy06DJeLONGoqHfeIRqa/rsp1IBpHNDLrdU3NAGm9RYNX46X1gPZZIJRM
aNx6MiZyUXiWGtoSrmXo8FvVu6ZqUOeWv7GuMUCqpnqf/4ruke/jFign2jYNAy4D
dCgIzTtb7tGahaq3mg9FQo3GUDkF6EehjszNKynr6Y1Ejoo9Yq0H62tj1U+OBWJy
FvPphgsCnVYn2GmY0xIVrirEHCGPuli5gn6TqakIBKGalz8ZSCuXnDilKOgg7HJE
exqrQRmvopJ7Fo3NMWoTBthtK0jel+x+Uwgct2of0cELHRrEJOqZVbuKoDh3S4n6
TjjPlEyzeGA+TVHxFnrAjCbex2fN6WpQOVF+zmPSUbQ7gscvmimumdNZHFP+P5q2
iu41wbI9gn4nmtPIHXehOtKM9DTE9KukmB/PDfF86Q1W4ADC++HEWhAuZ48ZciNY
5WxpsXkOxUdHVFlFGzzmMqsFSGaRJd3tHIpLFsIFHVMDpFwMdsrdli5nhXbK9ayC
xWs35fFeAJgf5VWedgu66aTA75brdpehWLFhENaWxGfCOrctc/spD5e86qw07q1i
viQ2IezJYIGDacbmXyY3G5Z8DVv1WDRltNbG2bXFDYsRXO+Tv/ekQ/EH6hwyuY2p
MBNdaa1KzYAn8aO/5MlW0yUYPrUHRX7dOjOCppWBfz8kkmO0dyCCrlbT1zLIRmeJ
SFpNljNYYpdPVtzgvIaRVmUJLDcTgM9IDLCRE9hmKPq7KXeMFZ0RDWA6vIw+x4KB
QTghU//2vHOuaETbL3YT/a+GpRanytWXUrOZLPLiW4FmOpgOAZedLefytAxOIiAv
e55E9XWio3133Fhx4T9/RYHypu+TR6NyQXwgP+xdjzpE1vJA1/rsg9byRWahYJPL
Z2Zp0DXAsde3J/17kioKyrGot+v/R0GXSFq/6fWultKF+3axlG//OGLvl5OWSnCR
ofk0OIPwXJlaSFc13dnzIh6HknRONqOGtCeEDqPetSTkJyLUz61rVtrDPSxwn/qa
WMxQm/XPsqqLtjICtlv1Gux3AxWI+YsW4q+TYvDmXjlqekrSG5kpXaOnxGMWkeYW
mUu8TOaAsXrc4CQvnq85YHPF5uzSnU++M8TKh/+m1/VzoLzUvHriQX5gOqJ0N+i9
bfRXwumHmkLJaG+vvXLxrrDNRCUpGw+g1GW3xVS23MhKQzePNS72a/eR1NmRbCoo
Z99UaMuP2XKn//FHqK9dZ1ybu6vPFrFlxxbeqxVRCb2KQ38IQ6q9deezQ1wg7/vg
DWrpq9VRD98nWolpH5A4lficLFTbGnDiQxSS5iqIVld8SCdZcgPS8wZIAxTe5wU4
SY+/Do/5p9M2dr6hj8cPzkcSgLvdlmlc4SdchXdg2qxwq9zWnwvnHjKCXVRT0H36
bxSH2I1V06+kjKzUwjyOeB2sKNNvp2JTRfDOCdMp6rHgPnxxibKzEWSE2wPOqxoj
Yrh3axragox773N69LS0RHYewhFTEc3MC3+vD9Re/8SWMwOWWXy7Hmp1T4t3dEC+
LPWOp7i2QJZ9dzb4hR0F/FaNYi42Fh2aaHjoIWHHQHCGwWo2d5gC991y5+RQg375
FBV8K2ojhShm6cQbH62ek/dAFipVObhEBfcti3N63iCc3PvvgF3P+9qTF0PWecFq
gaqdY9CSR0LGx/lF9T2bF4XiMCS2nPZflaNDMik8lRRABD/VJb+tLOjas9EQ2ul1
6Cwy0JrNaMaWCG4JKHIvnR9Tyet6Mj+szS4MvPPYjGORYKlGhYKgKFoJg5oA9vdH
Y7tC3CaLPkWIoUGznjeJGe6i8FRR/VCt/R64/wezfNAGyNMWTg6VFAbiQ89A+b76
YG5SNGpIwKTNoN+FzKlwr7QdcXv34oFQ+yKf98cILgsNNP9l9ewPj0ILJ7GVj4kz
ktmnSg3CQ7auVfLLvEyxwfnQpFiT1gTMEcJzDTmfepO55uLSvqpV0BbnLsgAVUa/
aEqYdBcSMbCX/UEzjQ7MWHIfpKFTVqdqgOaD02nrv3WQ7xEKTJSqoDqfG0fwyPgj
jbcyYOk8LHyWbnzLfyGTNb6akVOVja7awzT68e9LAQ/4HVncoSbjM/hvrIO2IxAp
6vXjvfYkBjSCndAw5M02ZiyihojD151KfRlKb901ew+Gt6Aiwtsoj+SqN+tZ5I/a
KHWciskywAZZWZc7Nk4cVk1Y7q33zXDjuhQ2Ecdy5I5SzT1XHb+eoHmNHj9gUsvm
/AUoB3t304H8cm0FdeAuL6aHuPBSVl48l/wLX34Em9fDLeIyrYLhzVxoplUrZ5m0
/0oiyxp5APbyVq11qQJcU6PjGuWK45GRsk//OwrYDV7wTEt06kNx1+OHDyWjeyZq
ly6TscpQkdTqPknMZu/ONm5yDxaLQCFoElmAK9iFLMvFvy5Za4iYUE1COEdpz+Aq
AbqryIjIxavuSsab9w0mhumlhQPxqZE12k+QqxypdllpJSsgjjCx1hvF6bFyTUOL
cuoDeHk+6fi9CqmfHMDL36by/yBilE0N7CFxOeURed7ic9O3rgwEjhXIGV8EA4CI
x3GKyqCrKC1Y4PdHDD4fdgk0UMMv0cz6ONiJHb74ptISYDYxRj7MBgIAsKhmcJQw
cQAM4FTASgIArI4dc3L4JQsZN8PHuEarrCgq+kz/Xz6T6zwQt6D5SaG98xv+HvpD
0EfiSL3qpUwCzQa0+LaPPUod1PWsW1wiBjT7k3PFloOfNMJnIig0pVQn+p/LRfEl
ax1GJnFJnHQC5z9HT9QacpYWd3FJI/2z46fomL6/ZgWkUh5JMGURDEhYZbI5Swha
bKRa/8J3zFzxRkSUtTkC51Ns+TLrRvIyUY570V1VSJtvWUY2jrBa8ljIlTceRzpn
g56lf+djumX/uUjqlnfQ+TOmjyhgkavSp8NEmLELTzkVr3Oro2gVYDqKYva/Ci8s
avRyNizk62LPLm/CFywUZIeZe2XOTSJdLc0S8OsH8qIuSEq05KWKe3ghtolhbb78
codMXPkBOOQ8SpDD2RXpMaDnwhrgFJcVg4XkenTHgEnwjJbeTDWSy9pbxHe/Awu+
3FOLDYAk3VOsXPBpvLukEEChGAFMH1iKLjLPDM1n5nmiBgsXDz4/ve3mptCyiYPA
Gl2SeHHyiEeepy0f4UgPEAGWfgd8aYuY61THRrLrlAESTCHTjdL74k3Pvtf7GGY/
sl5oXVF1w5b9Tw+sKyhR0azJhoCXfeKxO3LW8LcK54UIm/0BHv14iape4y+WgSlW
1Et+KVl70K8hVslh4k1CAIZ/TbX4Q0nVphhFYVYVPQvlGaTU2sg8pRTyWSprBPeP
7nXSkW6l4uolcJtgEUjnQvMWLOZdDbjyvXNKJZh0SbC1PNvEhzApNxxFgNK0r0jM
Txh18dr9eHlWsk7BH+LRqe4+E7ActmqNM2iFXv6uX0uDPNdGkwNq0P5OWlHKisat
eclyA+EAxpv8r1ygIyUIrK7ATnGi9Ze8aoVaxnsDwVulSw/TkK8TxwGjUvafkgms
y0De2FM5cVKGFx02KGlr/ETtVAVYtqXmeE2VVEuXNVBYz+E3vhd2OazsqG3pskyV
vD3FkAVytOpItcy0WqFpxOYjxTIJdW9eddMuQ2+ZNicvS844ubbG0AlakVGof1sB
3zF2fzrJ4xFa5B3/0E1KIFLDQ0vQix1YorWxJTK3HTt0gxjeGMomuwG+41GLefFx
8QghwjT2mUGq1w/Lupc7L+gsXf0jBlmVheB3adoWnMYfeNwhSERfMBFo1YyjzDBU
BK19ayfJzyasWm13s/OypmtGLm/u0dDRlR0DbadAxRdv37JFOh9yBEyN72/HZW1m
Og1QLay3/8EqHCTcF0Rwgmjrym/hga3sTWWc8xZprsYD7Mive+w9uF8zNhq3lRln
CbeNbJ/7pLkJph4igheKmyk7/DwmkjCIGuWUWSky1ifc1WLF4jVr2Saaivk72/EK
IixOm/lPNE65TsQjsxU0GfEf4/bnXktYeQbGExzCL2sR0t/nktqptEMnGLst6TuI
2JPobXfbNSJUV7oUO3MyucqR/vxSSRTa5d22JqIXlVPPJ2VXebZMvIiwcA0OXp0Y
Z3WaC8Veu6ipIupy+qbwwQdyaeGFIMB1ZIlFriPF7L6Y7ZrENdGLDoT3uiBeE6Dh
3Xy6GpaV/B+mHyfqtvcI2PBxyC08uMKIvTnk2+LawrzI+mLyoRtwnleSNmrxi/Zn
UB3z27NFVhLywbxXgxi29ZfPy6pbWbeiMvWatfNIux9liVcRUyQtUVaU3R6DUxiy
SnvB6nC8j6CYdfX2Bb/1Xslx84q9EC2iUoajtr3JJmm41pllLzH4cOMtIJhjSp6P
357QkL8DNlMRGph1TbyTTwMCZuqZaG4YTAGvIjWn19/UhuUpzvgcruqWEskaiS+q
e1VB+7GUpo17tJZVKzv5ojxsZKGanidhCZkjQarc53vqgMaWaJtqQXUWtkEsvFeP
ZN4botmvKQ5C6SkBmpOMN2tQBESsXIWPDpGAbQrbqPLzow7+S/ZFINAB4LIZbbvH
y95yN41CLLYfKZcUadXahyYOzRwrQVqfLHc526y7bhVhGalPd6PBx1LEd6vRAJN+
BRYpX7hwi1WE1cX4VDaFoRQmADL9tkjfg7yQ2bkvREFGvL+V0CDH1ATUNir4krad
7sOlzgCJK4e6le4AvKTOC1dtDJaQ3ht/3SxtWJYBIkSHhaRXxV/zPcYwZPvJKais
E6/2fD3ywNSsApLs5znxwzEUZ/CsyC26WG45jjQ7IhzegmaVbSyxE5+IBvn1eKvm
hJB4ZsQunHOe3KMuQCa43vut1rdupdHSIOQfxRXjFF5ZPpS5+dQlPEs49hvoLJIw
qYI5WKZ2YxyXf5Th2/LaRBurFo2ViqRXF2jVCXAQ33fA7GsSfUj+5SysvhzwGGbK
1ay2FoPoydvqG8fdp/JZNYEWTWfm0N6fpBy7DG8I3KAmG0hKozLsrHN7RW5xpHck
x7t1q2T6MlMgQug+0bDnCKc5sfByj3xtOjOz8ewkBGK2RJQDSNYd8L9jzOSrD7Mj
FZib1hyTbGMShLZ0Dw8XqohUY1oTwUyIiu96im9VqHu1kh6JX7/EiOloqWjBw5x4
TzkF+PUYqOjuVstW903blUVMmUX+LwDC4tel+Q41Ge8PD6HfAP4avrwOTPDCK0UM
2oUVu6vmoPFJEkkMWKukqD9drappEGM8pTf3q9CRo75t27m4lOpTVkPS4rYTptLM
hXyvKh5bPo8Z9s0WzIsq771qHwm4W6EcQjqG9tOASI3mRYajK2zW/ZeYuZySHXSk
fS1KUmTOSnyb7USheSD0N6m5zYPnGdLHm+6rtknvBfzoUIss9cxOu//S05HTsNXV
iKdfDMFefLyZAwlY33sR/5/S6J/tAfRDuvwU1h+znDTXF6EcBgvDx/K2vZYJNjoW
6LcQWwnMDLqxDMaB/KNe6cHuC7SjGXFOxDI6tYj+ySXzdRuIa6EMyDgvFFicPy7L
ESYIJpgH254Hws6vm4fKHXbZtt34GD8QZJsT1MDNR1mFOoZVHXS94scH655hDP1y
W5axNocxuP3W3G1H0AcEAQgUWzwO3gZLi/FUzZ+KbvlOgwhZ2O56FB9toKnxlOkW
p5DM+Lz9V/kxOr7txxT3vEQVL+MKn1qvObQcvMlo/0g8ldvcmDEoLht41BXC9x77
f4Wk1VwBcOHhkxNaFZq2K9rDNr7fLgHRnZVAz/817+z3vudqpm6R1/hpQ8s9ozxb
Laf09rTJKwUWayxGy+wnuSxIgfKYJXbaTVh8R+MmGoYZUhlKiuX1NEXydmg8NOXx
bI+nHTIENlUgOQZF2aV2gvDEPUyh/RPoaE4YoL9+FUYLRc3iCscCeGFtm6JoN6w6
LJGZb75aFX4AKd1xLuXyJQatZRXGemrR0PSWq6vyjEJaScZsEwbT4Y6LKmH3fpsZ
AVdUc5twtOyHoignZq4LZ3sP8Ui56Opu18YpJLN0xNV/5LeiOUCLqDqDtzX9pR51
Lco57gumu5ZbQcM1MIRhR1bGw8b1CEojtJQ0eDfI6L+B3cWBxo3EI50JzxDJJKy6
Kbp1JR/KZXAnOsNKDzq1825L5BZmD+a8QvnrKhRTWLAF3enwlCxgZfynD8eOPdHJ
xVFoKJHvIf8IAOa0zK1/zVQOZDV8JSNNB4P33g0kI4O2ttFk5KisDFucmoF5wyLa
CMAygdzgRJx4EXoQC8vQ+qbEbHVrdYMoQyHogVqoPAlj1Q4PBB8CFM/jERHRctRv
ZFfT/CoZoi+znbLa7PvYQMLKoLdItVQ3MFHH7pvzLpxTOfb39TEMqwC7wCwIyM6r
FryeeuGEUcVXpMcXphGU3bMMtYMCXIGz7B1WMsYEUj4qIbAjxUTR6b6VIATaCyCL
J8qARdM9OyM16FQM5+VOA56M3OlirQcqn3FyCFCto0QktAqKKGe5wLufZ0Hb6PBP
uc2txlRHM1mYDj0YbatQ1xTaNsybsNybd7LXVccTIJwUU4AX/v3pf35IXy40ra8i
JGfvC+DDWB6ycYb6Yi//qWU6h0y98sjoi824+nEC0fr1Nz6z0+OpfP9Lp5hGRfdo
s5sIniMy1jR77TPJHdpjCm9xVn44Gs7ct/OJw/zq8OtDRZ5mCjZaKbnFYQuT6IkF
NEepuY9dhIg/wXy6xa0MXbpH41riQ2DwGS7KF8NAN/wVN52sj6ZXR+NmVTiEa9iU
e/GIP9kap34Jdnq2QxF4zXBCl6T4KiwfsgNDpGbFtZHTSndn7RrVHF3vQfZxWRph
vwkZTguJBzdcE/8XM1+VztF7eInneXJ3PVEZzVzW7gREvF3U8YsvLzyw8hKaQ27t
+GnnQwZ0YiKa1u1qcCwBZRSqp35UrqSvHMeTGynImJ2C56WCZIiufjePaMdtx6lW
OIrsrmDD3HsgqmZ7aHRT60OCLPJFAQBTKyI4Smq2wVoJcrRP7JnAGGlgE+vl2uMJ
SzOBUgtKsFUp/8029jMf3aD13GGTC/e5CrFVDM7MdLqeEFB3XZmAAhCnyuvkfe1Z
iRV1Yn154gLTGzi9AGZO8K8WBogmDt3F217PXdjr9whDwglBrZ66L7Y+pojhnpWj
u02e8aYrZOSv1Wm1os6LyzBYsmFC2L48xCI9p3BfDz0WDV8UKfRe9aMZys3UGms+
fir6Ewn2cXwQzRrYvmgILauk+Q6wmfw0uCAHV0oVqQSYKqwcRjhnRgnT+uCAJZ2O
OXvpJWfl8TQqmyXry9Gbk8vHDsCQ2qvgNwzFtLbBsYCMcn+o6TRSXmg1LyCtWeSI
jPDqrkAt2dyYzq5XVhFA4Y8T3aDc99nFxsRQDQNaUe8TQRbD05m2pcQWe801e/nu
XYyUL/k9vHO6QeT64ephuIMrTZxtw/26C/GXS8kuEeXAE4zLsg+ksnvRbzK4OlrM
JQFcGNexJS2sttcJfv+wtx8ryNX6nk/cIB4NefvtZUVPHDhwS6woUXNvhnj4cPPE
aCUb94WumVOTHNa7gN3cVy5c/rGqmEsPo+0MN1+31N0wPOrXVGIpYYiYGGbhpwTa
FBSWunzFli+4VoGz5gS4ybdt6I3svubQ5dVrcx9g9+dNSZ7+sjxKWuQwuWdVTMYR
WqbWlkEb8PZmU2cEKZ83ASUfmc1PYtHsVT+TFbhRNWBQ1tfnJzaJYS1RBO7CPGIP
wxBLV3WeOsIclI9BPj0Pe48SvM2SCjuBgtGjEgfyKUj36gcqLkNAQkw5MpD7BM/p
DLLLBX6N3eNY/HVk//sbnlgmL6gFriZ7TN37AcfWBRhXWGt9NIYpSDIVo+0FS08j
MXk1PP+BI7ktGUTA5ey676FrAbzWIZIepC0YNoh2dNcHrDMdDJCD9didLMBpBDZr
MdQy3adIlC5J/icRiVdrowNu/jsN+KXv9AGCvTV5wWTakHeNz13WupHzmVQ+lQhH
RCZEfIiMsk7ZxiYy6rs2eblKhHkk5vBA5aFEnC44oOzybHDIUXf6IhVCQyERxpYG
tUHbo7kHYTs2btcHf0kvIM6gcEr7IStC50+0lG9S+dAv0lHsN7zUcgdMJxRIu+cT
/jP1EpSUwIgTQjalhL7ujzfPBltONxheEtJXARdNTKsoY1CZUXL4ZFVdrTgKeBJv
ZEuRfrmyWNWwBp2BHPbK6gTz1sdDXGLpvvoawvPZrnigsEwok67vGXVEwGLbjun6
UOeFvrlp4W6w6+pLBSNo/bY0tNlJ8IRruS2E/SmWHrisxPiu1GkjLQAqD3eXO5LW
7X+SRR4Qec9ZvGFg8aZqH/YxL0hikxL2CAaHSNt8E1EiJmlQ0UfMSAjJkVZCFe/W
GEGiH4hJZuvK2xOgDs1tTsmFfS5eYzpnYI71OVyBdx6lkVH65aaNprLdObYI97Id
lSNiG6wCKAHCriQyqiRPuKCZuqcOIWLQmCTOoDAXQU1512RouIsGCBYHmOEyzznw
vxh2dPrjh4tYORLj/6JCIEnC5tRPKaPVaeG/by4MIIcP7jfMCMzmwt5b33axBOz0
AfR2FIjdyQzeUECaDKFVQkgjAGjBaJkja0hgMMgHM65QeI94/PD/qMHbTgY5hIR5
1UmqeKY/+4/Aiuubk3nH2BLRATn2g03Zdaw4EeNQ2n8meB2eSgOlRr5SUck62veH
NO96cjNnKcxSnR2N3jMc2BXsBdlgXawdYnkEHRsKmG+oygPppolHqq4S3am/zL1U
TCHSRqtgrvWymdQ9YETJpI74P0sc3J8AY/CiIqg8XoLtVd6om4EmnC392jEpwwqh
u1knuEZeVqqIhyd3wtPOJdRA3SrgvBAUunEk8M65d5sR+rKMIubJHQbqc7m/HuBx
HCZxRdKgS3AvSweClwW+KMxsH9W/h/Q3ciMEWIUBFpq9ZIUFa26XdeAsy3uyHNFw
wBmhJDi3XDqElb0gKM1JcnCzITpTMtdoTaJYOaHmtjwopZ/T8JCi4nEzl0Z6jkVP
KTTfP0qJpYfDdMhtmdjx/WkSdb7D1h9u/VWmMCmHPpacLf0Lwqi2x10KSx43SQPf
sphKHolfMEfp+FaHPyVQPM+F+I3DpfNqb1XR161vmU/QrSwQ4ejVCwy6ulDj+w/P
icWdEXfINcUCPU65QgBtmYy3vRrqx08PTZ4xb/LINQ1SVwOLTb11JIWc0Z3x4Wy4
SDncb+Ja5DH4ZhgcZVx8uYMaad5lnOeNjM2Cb/O4FPFgBk4qNJkhld4/cRXL19aS
jvMM/DBdPGbd0nYggwJAMaZ3ZfKHkpyAxNAGN/71koaYUdkNFgrNpJORPUYA64In
EFYvzuwk5lAA/ty0u+k3BgV3HlZUFjin3D/MW4dxixaQixh/5dzBgmkhBqSXeh8L
Xn/NxH6xqfVo/j3v/AtCftkyDSnbZqB/Nv5N9sLqa11d4uLsZjTwVEDDLThSwu9O
NkvnjN7hHL0s4yslCvTBTpmKhORzXUFe27abDBval02jtfCO1fCeXxumYBJHXBiE
b/vriwSrXWX+jzMdbjhSLgVdwOJErx6wTgWMCZt++3BHXNRed5sAcu2jiulm6p2U
POH+NgV5AP5q5pIx2ELZNo0oJsUrIT+pN4BIRPoGwucayA8Jg9glkyhboJLyu6GZ
gIsC3B2lW42E6H4ly2w46oMXuftRTvZsXCyrFdGt0Z2JOUwB3tea/sTZD0/rpZIP
yIOql3J3Cl8FECnB7dn6sFU/JxyZS/wMaTREBBhdIWFpjrO2PML4J6UzDjm+3uoW
YpT818LHQevW3GBee1k4qeMyXCxhCXBmpIdTaJu1hOSs+6OAp7nBtHMh9GXwyNjO
EP42V0hI03N0dEmvq8+FKPVXroSllXmdtp1YqAQuEvu7UtO3k+jKHuna3XLhDsib
kgmucuVDMNdkKKlJZ0Fb9NgMr0yZqvOqb1mXuEmrb3xSZPLS+TuRK1YwFofMWDTk
XsAB4OcY0w3O8O/OVEW2aNs95QvaIt5Yahw2z1V25qeVUDDkwTurSOBiwE2Zor9c
j+bK0EcRUD/8amYyvpH6ahmPpY/M0HOlgz6lgonZR/tpkZt7F92IL9XR00eYVgji
oyplcZBSJ673gVy82Ckg89GW7w9+96yqI9A5bhZtkAhWPwbqFaZGrHXzdKoyiuVX
Mv7QXRuLJMwCGsR2kMoKhcymC1NLbIx4AbDZQVk/NG8hu/tKx7DJGTxTp8AeowoH
HqmJH8sbvXcA+LSp8arXLjcp+7K27i2/PAByK2VhbZo8U2Ks82QcHw8obymaRnUB
kuUBmq1OCabxfRgd5NPhO9XqUAg6MGv7mbZpw5XUQ04XpJKXjnDUqTlT1YEgLwsn
yIjGoaHNAUWoOH91cCX+SVwM071QM4Bo5RL1cWXwSwlBCW5LUNIypwbL8yaGwdbv
wj9gwnEj7nkqNn222uUaDEKS4DmblFXLAPPo36Nv12Qe8e60rl9jGqLYM2zfZNh2
ZfAqSxoM2QG2v2x6UB3IWeNg+TgXKiLXwkUHGHBUkYyMQal6V6owCoLv7AWG0B5b
6mTXdiirRkIIvsLh2IsnXLFrrzZj7d7H+WIOvcUKXNfYSnxU0MiW0OQCljdpTHCe
oi+xgWyuWJr7JrtgH5GemQq4oSV+ZutgZNgA5gtdLRzKJrGcmzK2/YoezLD7JLzb
4IH9htRIRvMTzupfNKit3AporqZ+L8iIRM/sDuLdwhFuFOldvmPBffZLRZQ94vWf
NkjYwiBlDMMB3jUgdamAvVKaAQjzZfwZQInf1sHGHQhGDnrbiCz2/V5k+rc5yOHr
AAFN/o3JJlbZR7vaI3w/5+zbZaEkOO399efoq9FFp17SlVEV+zroSWh33pTNXPEb
peV3WR5HogqfV4cMhololmak2hrotUTEWN8KC+J265p+pZ/uq1eeilNrnTdl8uMC
jLv2RKi2o9AfGhraBXW1MggAOJXqA3bX8abIA0+vaQnAWH24FyMEhih7ffXq5mP/
M42P4OaX1CGhC/VgOfCUJ860xRExfpF5qjLByA5skKq9qeF2s15/f1GEsUxHCOE0
rKBx0ywsBvnrs5MuNRZibpb7HGi71IaXhzOTYo6Q6svfxXMdtMcFHA2JoiC6w2h1
VDNxdCNYMXi2OhMgqNVEvMmwFfwQh4rGZva/4kFtxJFgCI5R+DFx5l04LzogjKKG
Hr6vwFNtTrsRZmnJw1DOythze/1BYNnNhHy6NZo8BGIyOlWtGZvlbDCOK2lPLj5B
kT/dIZKZg7YgJoo6DCP7Xv/+3wKNrltxal8ZM/4OEFlIEfRGCHtZBLPxpfq6hm61
ZGe58K1qT+qFmzN74yM1YYOM2cOK2IenGX1Bg67GasZvJGic0JS1ZWrLSSx6oTMz
22V7V8nxm8PBkZRIjoD+tgy4VvD7RoCITRGcmd8vthcNM844L1AWeZ4d+5pOKe9M
v1V9P9xG41xA3jmg2kH7DUg389mcQ8Nd/KaW7SR6Bipkzgo2kzgznxheRO1Ym1KH
EKUleLde87eiA8FYouKzu9kuSkW65jxOHU3kRo12emhnch9R32YQIXjPF4q9YyWo
+AikhncepeUP1XIy4EmOQEZYWZ/x8rT+DLxT9/y6S5N6v+gosr65+N5Q5uHp5J2e
t31v4gCJOZsZkdc1bDowBj4KqVaEEir1xzlXLUw/Px7U6OZm//P47vvotw+KPP3q
5rwkf+dauNrA5ydZeY9DLIGmu6PPuUoWznR+iy6Nlg+SWtLvAdvFPN/fb9qqjqfT
AXH1vjoDMf4S5f9zXaxia0PqqN3h7k5WIhpVyFsH6vgusmxWIyqfTEr7EJpCnYMS
wErqim/4tfnb4UC7KaHv5QOnuzsyf08IsWdCsNLqMPXFwdOs3Hz68i5qfW5hKNdn
H3FBuXHoBwhTWl+DGIaUmnFbspPo4tFKeWkNRnNqJ6dOJXljCbUd2g3bjXJpC9QN
qVhm/EkuggDcEaggxjKKA2E3zpnYIoZGZRNUlxDh8j3oFNxHHjh6qEtCBhtdli0s
dHhCUPqowIREK5RcuZ/BCbCToy2FFfo4uzak415SZv16Y5XeKpgrVIJIFmuru/5p
q/GBZjuttErlVtZsgXISLtjtjObaVsqbEOaRarJazXyJrZs6/lpImZUMbB7ZAShf
px/rQVAG/lCJzCXRvStYdTDEIvzaCp+J56OLEAOF5ynT9EaZGxvPR7udrlMSs2pK
u077BT80+Tp6tMlW0nbE1mcoE/iaB0/JO2Y+9jXkF8AUjdcTDOhyVQi2Tnv+IdYw
P+L22xRKTL1ZzU4HyKG0VyaxNokTZ2gANs8PeJmRfCDcI4FbrPtwckndNbj0wjT3
a0xRZlNzBJOHchllqNr7w0JBOzPFsBO5Uyg33EJ9hmgTpl4sd+Aar6nc2yZOpG0/
O5s0xFXw/CPhKY/ns9LvyiwP4P72fFvm+fu+XsNp6kOG7Mt0PAIfmeOfhsrvu2zh
l5nkRPsC6MaQeVpRHbWyuQbup72lxoguWFrj+PAX25cMde7tsjRK8F3kfTxL4Hmh
tCO0MXtsH8Gxy+Kvlr1kAbsG4zSWm5CQlLsrHL8iPMD8THQVW149qM8qY2MpxHv6
5q61qeN+Jiw+5zono0O4XZj49fQJMVJK4Hau7oKeBBEk07+IZcgsKENhxL1xPV+S
hEKtTmznvxunp1Qku1GzZVCbbGTbILDahOppJW/wje/zdCF6oJ3Fcbzuchckc1/L
23wmsfQQjQLvJcQWGAksPC2TJB64g/R5BAS9xV5ffbV7vuWayb5xDyhmFTax+Uyk
+Ej4p19CNJ1Zwa3PcDD8iAOXVEsxvsQPvCNPS+nIHXXbHzIcLzzArbXrA4CXcuCT
LQfTqZJSvYEMGUuVW/gjVgFjr97nAMufl3aQPLKoc7CwkzR0Wu18vbXoA6vFZ653
HGKyXEq4+d9+Yy4q2MUTikVC9kbH0Gbu94hk5ZQgAoDPvtfGoTf7lvYJ3WL7O/P5
QWZsBD5ZgsgtnEOLj4S0G6ixCBwT6U9EqKkzvTOB6B7MDEgVtek4sgjwJf85tS1R
JBI4U8fGi9Y0LmKsFMPeu4zu1JOvWhm5xn/lRS8lKb7W53Y4D7vU8UW+5gk0XRsP
J7ErSr3ihDgxtiMIGUGexGDz3wJaYqhCOs/5xT3JGoxD+cd2oX4HjVvF6iu5Wab2
t0F52Y7d886c8lCWU0c+9fZGHclMIHYRNcsrZrKT7rZfwgB+VAC2G7A8pW/ySXSf
M1LIo7pYyixvvBX3LsReBw233OmX5JaRfwFoFXIHi93jpBE7olf2ixYz1d+eZj3S
sTJyjsD2bnC17tWjRzqo7vrkINsBel0BeOROOFKCyWL5l2CbN7/Y6QYZ0M+j+lgU
5L4LIc2rJ1lnfsLfAD/Jt0xnmsL+kgx0jLgVxZNk9R79mh9k9jcDmMEkGwkDawaN
Iot7ZcC3hOjxWStwJhePaF5GzaB+N0paCNEr59Zf2poXqzF5aqqZ20YBBZkFGHNp
LsEsSNd2lLC8kYUputBj/7BhRfFizlti3ahGp/iExlW6z+Yxyz7mhsNCA9c0FWJy
gnTAdzqYSzdOlyKtRz4EJI/pnxH4L5KjNy/vbchR4U5UxRpOP7i0Ulx+gGmVpwTW
Qy77/pmzjSJ+xm4jcnTiC/fTNXrwyrqCnfkx4kzo1I/TM7Y57dua2+ZhS715I2qo
m/YiXbgYJJ+ksNPrweCaPi6WeFpsVp4UyuTuSaT8pSzhZVrIDrJgYM4wUvXP5Cwz
MenfSSSdDIZS/K70BPWMIooy0rfPTpw6bIANLYv2Ds2UdSvkCN3Ff3oE12BHtuj3
ekfXHFFQV27YIzBunAeKGKSSvFysstu8eDoaij492Mjs/G7vqkQUlgO+60cgjBlr
6is3vKe+SZjk2PG/GmatculVL/B/HlcqWokCd0W8u77Fw+0cyP8M4uWZZj230vjm
IGS02T8HkaCRbf0jPubtLP4q2PvmkGclPfyXf1LmrRfS98/gDczp5QwJNQygq5rZ
+d65PT+/7bORY73NWW4tTZVmBqUHUl4fyys3JBarhe4cgnf2UPbi+3HsxNezNNRc
d5oCLMtFiQogCFQs56o2EeZfjrCmOZujUSbfLTn1Cu/L7X1You18umnZRKbvRXq0
8JqOUbOVrrbik1usxvVM90JHDtOgeFS4W9pZ4KkzUe3TcMRIhSpDl1wuLYDxc1fH
d+dT7MRnx89pIDkhfAVltchC+eodITzUyytxZ2vWFLex1qww8/p+ShmECLzIz6Ar
NMuB07tybH8+Ka8RnpbsaJyshMLvqkB6vkmSjTDsaDJ/JdmqR3Wnmjy+4pC8LSoH
hPvIHgx+Pc9A0AKcY1nGMZ8ZHJ/Whm5Fo8viJP/z3150VPbzmHbQq0JNIT25Idh8
d9EblK7fXXIOjMAWce/kGkaKlt99TxADfIyRAl/NLUz3OXev90vidVvYS81qp3qv
k136dqtqt/0UDNyQpDyvjIUHVPDkt12GocfiAME5PXxxM2vmR8mfd2vfF/jaFCcQ
QT97abYounm1n41nPqzMReAAyEKamdgRgOiHBRvpu6I39BxwMQCZtJy/Vv0g15oV
9NHlO2Yo/Tc7KgtPPrdw3WFK/0MhsKpRkkBqmGO+VX3CZLesqN6VkyU+yY/yeJb1
tV1B9Cl9Zvi6ViO+DqHy+sI8TgUdmLWnUgXPWETJ2ubAvyIl127yOGhLVOD/XRhT
WAhkG5cgkHRslLfhlPRjg8tFPj37islR8hA1urYnadIvQ2020QsFuzJeVZJU6Cph
/Zit9REkOol2QXaBMSvDLP2313qcvp9O61bE/zW5YBTBuM6mp79+uTiMoHLTX3GT
Crr13ple6wDwsrQT0jj+yrn3fAL/IeCPoHDgUTVCQGZofAQlGZ1cFCcB1OtCJ2VB
GRC3D3NDTa0u4pwnyOy4HhPjFwUCAONe+Cio6VOEWINr9d+WQ92er/+KEo6Y+Vc3
G5E8FxpADcwfxsch8XDY2R4mMKhe32i4IbYm+Om6ETWGP8ZK8V1N8gnHQ/Ft9b0k
X2PNLeNZicq+JIL44DkxM7CBLXrlkWStszY3VH2ftAWkPzeys6F9HmjrDPnKQvqX
JwDAeOR2MoKKpMerPga7G7ITvr+BdY8FHQ5O63rKR0+08mvJn4PyMe9BIsS+vgGj
A6V+L4alZF3UCwtozp/5VzM4sYFAICR7xYaZI39rynhuYo7MH4CDSKlbaZQs2BUD
8BdlOfwinOHML45AGRNvl2emkxVXEja/xNBNPTqOaFDIei26rvl0D0iYMy4kEu5n
N7VdnR9SX98uvMtWx6d5qdaayUPlbWZq/L3nkyQoLa55P9cwCg+xQ7ZDSOkFGkZM
OjY+N7FT31i53imh8p3qK6W8WQBVTFKkFn5sygKqzDaza8Yh4kxzEPKueuOq0hJy
bD59j6WvNglysUXApcyI4Ru8qFBRk+Bi+LxK/vGguLOFNHz7AF9YHrRSnnkrsWYF
iCvefl3va6Ld6ntgcc6FjrpP61/7bZJrEg76SL85WSplL5you+wI6Qe9mCFpWAzN
kFH0go+rMREkLkrmDS3GQK6qb9PA9kjZmvw9i8L9I5jSE4faMnIvy2HLEXW6h3sW
mkwkazR0fZxhrEoBW+VgXo2f7eyqLD3E+XX8XAR4BHMo5JXlfQ8E1QBW/7iUiZbv
lsYUKjUThT3oe0W8KwCEG0h3T/YtoQRumemiVHfakMMOUWmq87IgS21PWCK02d6K
7E/pLZSdNhTGLnsww3vMqANuXBxAf74SntgfaNFmaXAoa5Bmf33jp3BYnACtgT56
DIasFua6TdMpGev9eddUZsvXEhScxaZedCFOR98isGNQkp6MuQ5nmmjGmAaON1nv
UCAW5aeEAH1UE3twfTHgGpHum+9SHA4hJ448zi+3HP8iHKsPgHRpjRYNaKoPzKb/
3yV9QBVLhE1kxkecKoDH406rXSFcHMHd+0HXZ7oJA4u4EwViM2EOeI61+u0uBIyZ
nrcYh0zLm7ui3/HoD1zIQ7qHWUmrTMEC4nsIS0FaiIK1RKwsXr9PprckEhPjLc+B
7zdopoH7YNu5nzch4Vd4DXI4YpwJDXldwgJaZhvPCmJiDZjzAsEWXKL7lbIZ5wG5
afjk+S2VJ8ZsAJ4AgSWSEnIUv+Q76DzLM0l7V8mFhjFJRcb3zbM2Vj/VCffqg0ZR
RfBjUl51badZYbzPj1B7/hK+2p5TUgn9xgwTwKiiPr6l095SX5QAT7l71WrAlA8S
qUYTG2IYT1uK3TvZ3GxNKdLmz2xF6GCqrXGkaEPEf3RXnc5gMgthMO2+xFtML1Q3
8y6P47/0fm0phmQReGiioOGRvGPruIJ75Eo98MFgKBnEIpA0h6ZZW7AbIrm4UjvH
18Lk0EdMW/crD7UVr7pI0OksOkntKYMIt1ySYUUohK3iAT5TTjF4uhviMUf/+jr2
cD03VCOZlUnU6p0kslG9xlmu6sJVOsJggg0sgGgxt9suSz3avhOXRQGujaDLTCEh
4v5vZY3s7ZhDzmfZTDi9Kiw8otZjZxtBGjg/7OrTXQQ2sD4ZesQSQjnapJl6SYJy
As1pCKk0HlrV0VAsSKauotqfvyxHE+Ie+blpc53iJSoBtWbkEkqPKlt6W9NcxxtB
Ez29jBOmvd7CxE1DHHys3h2LJixsG/7cfSl25udjGbL5B9k+BboWVRGIEbsP7bKI
Cb0r32g5I6LCXZ3e1sHb8r2B/y95sykdm3W/2boWRV1lBcHDWE/fPm5Fy5hv0r2U
QhWdP6BmpZ3TEZH4gc59SsFZGo/o/Nqixoq3lvbp8F9qnsWJHWgcmAQm7mRS8R9T
uD3voUaokDD+ZI3nxHtOnFSxobeIohqTXctf2giyhrAjNy6mFOC/JjuQh1Ih969Y
hZcGcF4DIyZmbT8Xx9z0zFfOpyyotvALvjUD8MmIrSPP8Fed7e3BYoQkWaqJYayD
FZTJLPyv0BDqbQ80mFaR+duFQlt2IgBNziIhKsbhz5PEW8MCeaLYVUO0KSecRQQL
3RhSLF57KAhiiOiHrBNyNzLEeOS5/QRjjKYvtTY4Sp/Jl3BmrE5i/xCZNTRqJBHo
LthRGXebJsB6HKLMJs7EqaBclMllav5N9lWovtjrsWFrGct4mEk62BpqFEyq+m33
7DzCfH9VKLCAUR7oSJO0KUp++9cOlFO+rLZ3R2vE2xgDrYniHmzOQSlBYVeJ8Mr5
HhNXDsUpOT8OOamIq6P8Q9FY0UOmGYM7MdUpZujPkbwTa02H7Fqu4XVTkuc1NSkK
zvo8HwG9/ftboTVlNzugRg0ydGcGMVx6i8j0qNgQ/nIXZozO1IhX+kZELVhUy5MI
M9glwHuEc7qXtat2F05W8LXyAp9Yi7EX1BKekLteM/mX36xJGve0gNB8fUbIQImL
nMzyLbUwFl/6/xEyk+wWLnRBYdzwVJWzo500phKiEzT351n2dpNRTexLJxAsYF4D
qhyn1XkIJiQOMv1TzwM19VTHyuBsn9RMnwj3v1b0tfZP+yKoZBppbXYEuYSzfHI8
FuDNOYwWr4hSz7Kq9yX8Alu9Qk89YntzJNj2dj0hIPawEv51QSNchRINMlhqV2EW
QhH7oRmIQOmpBaSnHIMNuDGLxaUB/RTcIYGDMZ/puoKAYC58ELaYQPwfqZ7d3tbd
ZjxxacIPJkpEujKJVZfkQnOwS5omHpi/UM/ZxvPBvujnjxMuo5VOh1Dqw66sW9+q
U9T0LHBL6hXUwHKJyP+4WjlwPsl3UVKlgYz/eTTriq6VWMzlp02Zp3edOmojUyjn
ijlKe1ZGcQ34fV9BgUQ/zENu8uBK9vvVLNvQdy4tYioVu1A9vBGrtGG7HGCX5XYr
HeZe7aoswVdM6wJxJAdgkm8Rzo/sdrAfVYyQAuhK9glMzj06wZ4XWm2MOoKtVDyq
8ofZcc9t9NgL1diyBMw3jRqUbU7y/o3yTiJbuRDv5sjWpNFBZYG1WAwKddmvqGOL
prb0+5mvikMk505YR2m20aRQcnFFnBlOp/4auSsxkSIGkfefNbsyQEsOJyceHqMj
xxc8lSkAOxrGi432LmJt6Q+ZQ4G389hiKkXbip91SdzJrRPcNzFT4r4X9ido2sph
SYFQzQL0iaG9XB+pYNCM6ZtU0IIp7/6dQc6zl+j706saw5dCPTjRxeyi8CdryT/1
OuwyQccX/TVZCYXWZ8fGVdCKJP40kzywD6gB3Z1WKy2w18deuxfPCZXXkW//dI8n
0qsKdOXA0h7pNPNGQhekSHeA7OWZsk9JAObMJfXWkwUlRrbasIsusF2VAoKvMBt0
bAIJv0n73dUIlYu1NXvMdR/rjb6Onj4gE4rfOG4YUvyuzbV5E0QKYa46qas7YQLv
WTINr2DhBcc2d4WS3/tBO0Q2UFYimDydcg+NA//8qt3h63X1OpZakoo+fZOdLIkg
5UMWvF4//Xe4oTdjkQ+BxWlYMZc7M3JzapSqlXj2V2X9otdW0hQtn4LjAwTqdtep
yRdY/INSfwbsABqRy3Rojy2JslUrFZhTxXHcVucpdL1qbKVPgaFnp8xn++HnW3QH
apIscrcwKu67k4U8OdKD5w6aJqPAvfNwLrmDlrBkapBxJLaKvGsR9lVy5U7pORSz
rEap5eD8w7BP5BAElFGKAUNtJ669FK8RxqT52OS2PLemcCzM5mvnlO9+viIY08xU
puTtp26pNbMwCzsMRKLFpOfM5d1QM77bqy4oEoXraY4GnFvwqU24emNCO3uYN5Ue
kLKWOZuj7jdoQMokZhk5tpP8hl2Ex8o0USJTN93WtxMsiJSIciYPv6QM4I8qFbJR
HyBn/iuR9g7G+erg9/TVR4ZMFjd5viwgfiGXV5Vb4IN216lucQtEMl6FlQVw6LPf
xGBhxIPebB3SQumNEKCnvMbIW1R/BNB32tIm3y+xDL/xbrKEAPhYXp8k1LfNCZEH
R425NVd9lXRw60CidFrw5ob9oAjpPlHT3b2pD7ydk4u2z8qnATTMB8YqXZXj0eRi
mF7k8bZybA/vKdKnyY2y6VdWzbcf3owr0UpkP2F+szgrPbCO6wgeg5hLKDa4tyEL
XtznRDIHey4Rez3PhQwP8y8TOeO0zznFKbE8MaYf5ZN5HPFodj9oJPKyRLcN9Viw
P7dLP8LaavR2PYXmUok817DyzLk1e/U46OERyqAqoPGl8nxwIorADN5giHro7T32
r/EAeLXTxdUasgP+2P8PGROq0dVMKCkZAc4nIDBHl9dBDHxs5/G4q0LAlsJztQ/M
u4SNshpzDbWp6XD7F7fG6zRQRBv06uvYRP3o7/MLLHdz6T6txkXN9NJAAxniRcsa
FS3iFKcWakJv8ZjbK76u2GVLoHQ2r6kqGKXmtjuGknXSXj7kO5O8ZksG6UAeW2BT
9dtQ1GaQ6qIlToBSUoBrNGG+Xtbk6bOTP72chCv6BuN2bZS2KjwYEBPFCXr074Z8
s9EvXEt24v3kRu7F56E97MKzGoaJjiL6y9sgZAny+DjCtMnF8miJ5b64jGGueESd
r0y71Nb3IEkl62YdYvfY8ELBaZOPBG8rj7rKKh7lLDOiA/mAkGTEs5TlY3U/Bxe+
OKnm8nVxk2zF6eHHYX8D7nRQRqmCCbJ7FVYMpd+GGg1XZ810cRMnIc1fVVDw4TiS
DFBFH8GxBxHFHEHRLZuqdnWyxy0o0htbqYw8pBuiuhhApv4+HPihWBJ1Nq6sEcKP
5eC/OhtAfmz7iAQf/MVICw3ENtLpSjRt9JLmKfZtcP+WOoetUDlb+2QLSgjJcBKB
GQ2u4pHqs2MZQr8nUhSAi2p4xQ1elPUn/LvO9e2b2tiT32LdPd/mPsMsndKcFGfs
IIRqQOgmgt0yKDEqn/O+sCF8T3U5S1pIJh6Pn4OdMYzBD8OirubVEAzvADoEZXfI
/UYHuLqSZ52wLVyfrKjaGPEQd3SwiucQl4OcFK4IAUQh5AqUzf+Ip8KT/w6vggMZ
LbdJVYXA8XMtcR4xWaBb2dAy0yCbgRGspasgMZBYz3ctgHgBFttOsDXHswYRbw4r
ZtT41CPQiSw8wayXTDHyixRwEMkzGm51XeSp2M6TolGkEgoVfv9VrZwy4bAIe72e
0H2hxKZiDKbTBDNhRUzFgrOhIBNifm7mD4Dup2I9gF6ZhX3Rj2AYwDoq6eM2X8Ui
iq+uK+HX9VSBkshplYYgaZpqPvdDB8EJaOLKrd0I4P3D6OEtayKT4J0bgS2o+lh3
JP69Kl/jIZx5582bxCZdqyEjZ7bWm+fwx9EV2g+HZpVfbSWo71Goo0TP4KHvwtyS
cc+WIwGOQjsb/VM2O3MoE68Q88MM2Haqh6UaIYiOAkyeMz7YSuJmGKdxcB37zFg8
yvjME+kZGrNZCnghd1AxOaUC8NgRYTHcqfJj7nxeyzpu9m+TCgEZmAcrDlR4Id4G
WIeHxJ2sDhg9YNIxYnrOeRsnpfI3qp2H2NBTN8gQ+RFQ2YOTMCx4TIfY8ocxo7FV
0F7bbY14bua0tps6aHoeHXxQSkmyGQpCLsBQ+4xqsluYZdWZpyF1JKH8IL03x6pz
ulPM2yhl7XPLyRRsvrPkEO05EbKZ8M5gW8G65/q96jlcJqX+0Bkwvt8vgdVNBL4M
t4ReABVa0g2IZh9BIokinBOuGcPc/T1GHkjzAXh/nYZ3qG58lteVqojkr7fOdVQM
ObVOQ5ayXmq38z0h+zcOyrgns3mLlpVtzjsAtwqymC40QVhr0PQKo+lFumfgS+Bl
5oI4Q4Q3wQSmByGrkLL9AMjHdDJNJzE7gTaR/RjgY3PDMHItEX6a+vwO3UDjwkNt
WayLsYGF0VJE2MP1doUgbp5T+vcDfWDB8KROwG/3wWD+MMkTGGWlp5KZRPnzS15I
2uR1b++FTc157iIRR1vaUg4GiCF53YO6OybTrRFuT3JBvlRoa8gEnQ8L6seM1uC4
N3G7vWqOPHgMBpDaeesUf4G2s3XLqFvt1UE11NoNxiK926XTx2l4qfSV6TpOxR3a
Cb21BZDCn+V8Xg3Zc/+2faEWHDqiYZi7rbY+3V9/DW9rQM6d0/R2Noj/eREptxrn
9sBWGzLJjgGtR8bKFW7I3vBhNxhsScCPDJ9OyKjfSsOzY8RcxedGidwtir87+MRe
IQyX7tOmPwgfFhLuGXrlz+CG1FwXa6vAwvsJXjp+K4UgS9GYPCBMYVj4bCQj7MWV
iLXXyOq/n8YbtAGcOxVZbNws8iLYSbm1iGib3yPFsaYyzxhWqn+khstngfKAjTdA
MvNcHJdEz2ujtZpGYZ7/F3w5U+gTxvHK8wvwMVreDPHQKm84R36hzt/PIAGfvPVD
F0YkrLrzEKB1gqy7uWvLGAIIaciTtdwqzDaNqmhx+ZocDfCGlZ/XcZb7d8qcXCma
zCZYU/oep6ARQTrla+bM7kv7BHcx/wuwMMAYYygQqalSFzZLZvppOHJJFT6vzxOb
2pxFeh2AcKL02EFIZONgKRrJCtWOEssSQQvqeHk6RGJfdLmPM9opfGiBHS4D/Hp2
17f3X5t/YQUutMGe24EzA1it5EvzCU7mrXi9bfFAxHYkKRkghV8SszGeTVw9bDzD
O0E3YFcRmKuLiZNTxdawIOkh68DWVwm0vc1y7Dml9d8l9DnjDBa+3B82FRgLvCUD
iMDbIsnFEn5cTtjj9VNl4eH8JCI/6NDgBnORoSaDOU1amxs32vwWx/dMmNYLhF/8
77ruz91vG/YH9rbst6WRu0T67FIK29NNMSGu1FfOidaNzrMitUpgQZMnme1/L6Jc
wmdXzRY89UuzF6b+nrWcWI3xl/EcdfsVm0as9a0CUTiqvroQobW6AMmCP3OAqOaT
2dEtgln9K893bSCOnDXXKlsXhcpeD7U/APE4ZZmcVquRwEAM4PuUGv6g/hfdv1j8
9Ebg/wuTu8pnb3Dfjg3FKWASAf4B3fhNazIeMxukg8pzUuA5WkEJMv2qjSgqU9xz
0zqVzevBBV/MBidSk6y/9OPFhVJP5pXgqKueKOTXN+HaZ3CbuteqBhRQkixucb3r
7Xff9AjEKvp0+RCH3Sz+fVCvkyP1Pl7BkHDWDcLy6YcfwYxmSdODJXcyzXR+MIav
CpwuDeLeGxSPipfGamHWNYLIMXCCG/x/roqBdYHQoBW6oLkljFTYKXvqlcfL0ONF
cEcqLyL7grEYqQDCtoEmPytCR/hTJ0aQjLdH4LyrqzUDOdlLu0Fbx6qaDF2tpyAA
5pZ+uIQTRHhYvqi1TjmMZs5ohH6plDxpOkyPGxrTvSU1T/IQ9hYRK0jBbjSNZa/s
EkMBA7bcBZU+MD+QYb1xyf+FPwoHOIVwjb348UpP5vohRz9rAdsO+30oqwI+nO9k
ttVH2pVQCnK0UNEHPstPO1DYHZWy88V/v8GxnGnU8fzNV6oM01fK/L2Tax18jtUD
a0k4glqvShhbuc3qsd7VZO2VdNHD0MxhJR86AnJDlX3mdCF3Yd/sD9TF6h/h9Gzj
2jhBn09cMBtkYIBQ6udsXNP1z8RxtLYNM0SIb8fskykGaPl1K1IO4xQ5T+JjKYRW
qwu73zSiVR2x3JAmcu/ASo9Snns6lO6iDJ8k+/fPuUPiL6GXPVrqfHUYqXcuj+Vj
Hq9MuE/2ddj2b3bm9Ro1USoc/IcJAOq+yaOxmKCRPRLNJsnn3WRqc96TSPqZcOtS
gtKRXI9yu9kHwmECO6Wbaje4dotwSpxaAn1Bt2igbC4ALbCTF/wrBFRQBWVo6XCH
pQ8yFj8oy6bAGhWTsRJR4lA7GApS6y5cXa4rwZdx/11x4I0FDmt89IjGVX0d/+oa
4bHnE/DN2LaR3JcY9c4ZWSm2Md3tpGv6KtprnngHdEfN9B48SqGW1gy3p9fvJMBO
HJcEOtwP6U/KCAFzLm8iytUzlflCqNXGExwYatSdaF73EAN8PC0IxuyP9S7Txruv
eJjoR9dfpZ62nQY/w1SW+mM6LaU3qnPW7sqnsRQtl1ziJ+QAa+Enrty8qW9mtx0n
jJW4ZireAE0odPviMrp0Da72O2rqwnQ9NH1YyHO2EmZxOVWnqudaFj5Vr4fGiiad
mMGC/kvKm72VEk3RxCJkX2NLZ/muAFfmTZEuxHj96D5gHasL52n6Fju8WCUmT4jj
9AhetPp0Vk0Ud59e+zDNjlJmG3p/hd/qqN8CmtrypP0v4JrhmZ227DowA1mLAAQ4
E2C2Y/4fgYQ0FNv0OL5slhhJROMhYUqW/oFYVuKy1FxGAv+Ql24qTQxuG9c4q/00
bf+gA4+jsc/1B2gjPBzZ28kdgUjHUotY//BQm/h0erq/vcdhD4h95B/GZdb8u46B
YXQeatexTQl9xeGgTf9b4NBenZMswHO1AdsEwvN8sP7gIKHB2jHwIjcIC3bOIX/M
LKnTthewj9jv0ZwOo/fFbJiPhB3hksLwqkODmjnce1IbLXoOei5CXNJQd0udpZWB
aSA0NtMqaYCddynLFKwLbg02GFARivYzbVTR5vlfDTHcZv0k8mHxYHDBrPee2lY9
VmawUbZuOXT4Wpfj7kCTVrtI7yqSho7IroobiQFk6dwAldecG9z4TcccuXMtmD0D
gjYqc/Uc0XGwj1/qQprThkZCVd+p7KUt71lGdIvcF+XuCtVteDk09T7zXMTyFM0p
83MGBESWwxc3tE73ZCvAQEIy35Ycwc6hXehzqbh5yvhvfXT3HCTVCZpY6oAFVDTn
NzIdgkzUFseEAJdwgg1o+5pjRqAQVwBEZ/PJmM0wxCI1VXFD+sFsFFwByfKWV0uK
N0QnE0WGpffudYpisewxjb/2FqB0bx9/tlev8ely67Rfam7IGD3tFY/yKMrjQw6d
0p5j2blQb9azLa8iKebf1YiUr6EJs3qc6oryDR0O0HioWHKw8RV6QDa8G+W3rveO
Cr96C7Ha4Lh0K7uEIH4ZiETvacMs17BgA3SvQdUPYOFd+FVMUJYRtWHqikPZostR
FnrBUbEsathXzWR8QwcY8oObq6V9mqg/8AwT2CKL0kJ1OTJF5iR6fuQV31aVGg4O
iAble/5YxeEoXjvXbqSOlkZU4R91PLHG/33f6AhFJWDEMzOodXvAh2hkOx9b6fay
+TgyBuyznpeQ+kZ54bgaEaAGirXJFeYzjGZ6uxbhh+6GC9xO+fjyrff47YoED3Mk
2Bud7TF/vOfSe6fMoK/rmAAQtWkXFgeF9TswhWvzgmGnnDCeiktbqXrb7cau6WfK
7vbCpJav1/1AnyGPVrF57XRKj527wKNAYeaCH/UFw7fX4p9ZXw4DJpIJN66EORto
Cu1yPJwcAm989ooesPf4YP0nPn67R4QCHDDInFIsPpU3DbOvKeY4We9IFMKfu8EW
/JipPLrIdpEVsZNLigNgEO+4B5tJLJWOQEF3kKSYbhlWul7rCCaFojHYxXGfah0E
kQ35m7GKUmy1DdVFjw1pUzpFOtchRZ43hHByeG8RYePwET0sBA++18IfNkbrrZhp
PXP6WlkD7SHyZM3a0qABaf6z8UywECet6vP+d/cW0y0ndrAhYAlgc/DV5Uv7QKLz
OCFVL+M+phC5KT51g5/CQuIwV4DEewZ9p8Wh2QwUv2h/sYjpMqPNJ+8l4gWUoYNy
92VtL3KBcl6929C0ag+cGOnNeQoJ7LHPeootN0kZIEhwdvMcISZ5GQxjry8ib3db
VyDp0I7OEkFE6M/GGEyOTzmVG6w/YyEYKg267Oxc93m3ZZ04JPPocf6vRYsa8O8M
EtJwCw5PCaCJChvKVVVVYRXfeLnjXhV2CwKYFCYYOVDQVf3KXzBbNxgt+LYifkZK
mVWYShrzChtSgB/I3Ht/+s+3wFM49w9iFmC+vyvA8s+momvjSjVRIBzmSfFkMnS4
Oxh9jL8Ln07zwMlWotssUjvJhTQSNgHXhNJHhNEATC3I3TR+cuDXASbK6M57h5wx
fgkvoOUMBjf/1+RGemWXOLdTowLjO/zp3z5k7M3NF45UDu9FQ/l2viAb4UMQ7g7e
irOy7EiZce+iqyU+8XNiO3YNjonVY4Yxs7rGxUG6XwYlPVVnRhFuYP4MR6OK4wMl
vdVfwrY1OBFyW1F0TNsOQf1DJZmnBzRHkeNORj1ZZIrTn7jJaeCAPlEoqRA+itts
WzXeO8vLy0KjOsyKPOvJhOgTNDK7N94t+RaDIsz1qcSgDblIGilpOk+gMTwIyBXo
aEfyU43AiwcTd9H5Mx1F9mwR3o6ZeBhRE+zVE/nm6u972RJub9tKHGkxzZz/50JB
Pd6FgosuuPZ3VAOwa/gTkdOu0PkwIclUDCdxUOkmNLIdNKokn4/NdWZCMDj00TXX
hMnv5jzKxxl28ZomOo/EmPOYHpGFm1bsoVkvKy2/rNORg38YnwOtJdkA0gDHewkK
hwFK/cefAtOesNeRhjMt3xZgGojE9jvgoGylHR4lJ6GF40CmdpGuZcYbOdV+ly7X
HBJE606El89fRCIOXTkwUwr3FJSb3zO50OE94vB7539menAO4PsNyz0St7qkzLNu
qrvGBWEu4DG3PKvzXE9gERNKZ/K1/lsvtY1TBwl8ioHuNTBmsziPzGReWUSFJXfw
jQaU48biKeqsvO+7J5Jrgec3m4UCIiCjyGttjB4knpzTtpFKaDIm2P/f9z1ZQQWr
0N7bZAzyxT0UbWDiiHJEbDrLcGC9fgSblqc6PVjjIoJwdcaSQiGUGDrqJO/V+IaW
AjyHyQ6vAQ4wWJ8xJ2TTHc9ZPa19rvk2SHluWUd/9hOjiIQ8t6e1cG9K9MU8M6Zq
8CA/QBdItPQ7UunCN+CZdYFXo6jAlU4BBL4ipVp1+xc832XHjC9B6px4r8TdVxPu
371WUQyUv/AHGRV7UqJaHWduPmxUyVBxrWxWb+n+V4131E7qM3AKKelEoT4pgkv/
EVo6yQ2qGlQUd5qPpt8ymg+/WRO/lFY+U1PiN99fA1zNclclG05sAU1DwwNNPP7Z
X11ai4CLsdCnCdm5X0dEtPEJz1KSs2e59bMe7R3bJ0N5/byeCQ5AYESofUd8D8sM
VqawztsDPJrBJV2DpZ+nfibrSv9G5PsFGdW+M5QB6uTxhm5X0K+bgPTS68QtrUUl
EOETmgtmFAKs+bBDUqU6VJ4PPc3RUxbhZ2/C9vzTEGIimsNA0ACl4f44RqndoRbS
eTyM6gCjgNKzOrXzPEWCMCyK1oOu2QxBRUV+3VKLm+Wo+/j9MjWatm27h0j+srKG
hD32Wlb1aNDM+3MYmcsDaPfKYMK3/Ax2ROe1wb3NzMx2RLFxdwVE24tFvmtwjmyt
3r3rRgqBknVzJwNsc3heoqPtixL5hPdZRuY8T3O+k/HCM3rSDHD7Ur7h4YwDTtBG
SbTnYrRAGwzQL7CVQZizv3o22ET9GVw23KV67Mw5EL0QfHgJ57BVXxaS7HlmZd0I
56gnQB0bKGpjTEaZgtq12xhoG+1599FIozmd/l1emc2Hg/G+xorjj9xI/KP4iTt5
N4govz/YblDiJki7dvyVD5kQYaaOyONnpw8UMvkKhZZeSLXNGFXDbJx3wYZMdSaA
78KIx2mC16jPyaP1fxYF0MC1EmQFUJlj5wiaruKIEL2KKRUK1m2QmkqKuKssQ27K
fjhAVaIv5WEl24Ks3aTWqJikDGgtcJBdjpVKXur0xsus+fCC+z9X2H/9FezVNZVs
c8j0iK+27h6QEQE71q4j6PyUBKgdpuuleVgkozer5zS4iBlfu+OlBUbM77qiyQd7
uH7PHLgw9KkgJZsbOE4rivkvYgqZ5CUQ7Kbvn3qPkl4Mdg4a5LDR0sSS6JXPcRpz
S8bZ+lzM8t68jkFw1b60pJVkx0mwb6YXEWVahFzdf6EJxmnimVvdT/YL4ideOi97
FRGhCD2p8BzvX1hOgVFh4aXg1wLfLsqXloocjWBh1ty1i6ozGbLeujFHoe82msHA
kMBsZUnxAGkjTP/3gXgasC6O39VexemBV5sDYUA3NRvw858WX98fQYyGPTm+0Uj5
ns2lo5E7LBLzpRK5WKBdEUAZ0uwAc4fhSPJWWIkSefWQfmDI/qSL3h23MVuocPWc
xGPVpWRL5wwjNTtehbAprLC35VNw4yL/IXvg1TxxGS8DFiM3+JDq24Q28VR0wEnY
wCy9cCYXNuz8RD0Y/+mv29UUsAIvYmMN7rWLz+/hYAfPeOJ1ZXfGPIpmFzwXSvds
50azvvzo+B3iXFJuG63tu8fLLGxz3CyKlwG6kXNqQ/7dGeonYBi3n1ctHP03sxOD
T8mogq2gDYmgBBm6064MOIMdd04W0CZn6nwjKWsI3GLzff/nzawW67zj+ML50VJ2
tW2wMRzPhB5wzdHI+F45xFW+52KzU1MPwIa0jReYZPKU6Leugi/a96xwjIXB8mUo
5jmBbKM9b+f222SbDocvP8fdAS2LQZCyZDFvXQoWotzwNHTVRTk8PvB+1ZAH8QWt
SBJgiYKgiaoF1qWux36KrJs+63a+0Cc+4TDrzhRPaf4Wmr6vliHeBX6PncSzhCOz
96sRdGbh4PQVSHi8ZjPojW1lxzypqr3H3+XlH7g9uOAE3CxZ8SvdKV9SOB+UxJPr
6cUlhtgVX2Ei6dNdUFSYv6tRkiHIDDcZNNXwEIXe2fdn8iqjidliFgBp6Lm8voqD
ru43LPY67hH/iW9oRGb5gQyMgbHRy48X2kmmKkp+nkXpVMpjPCIY5EtmjxBm07p1
XPfo7YKSgggmH6KixjfsHoRm9eaqD7jPj5ylOSTq3iXfESItMgPKa8YZW2XfaufI
/Vl6TVgnfdkZf7TOeMqVIuKFzk6km8cwqX8Jxv16APi6P0Blc8ToTa7uv/9ifZbb
9eL7rGFAkuzgnY1xBIm8VWz6P60fuar2jg9yKGTCKun/ZBoUfb33nHvEXrMkl9Mu
fWqyf9dSAqoJafVxMuI0Snr8tVu+eNXIImcb0BgYpXH1N0glIJo0TBG+cT6S4KcJ
yIXW9YFwJRRDdwjTbi4zGb8zudjf9n3r3oEbt915FTtvxzuTIBgGuY1mdyrA3dK4
+BMkCnEMqPFJaYBnaFKquLnxgUKssYwDf80OqYKMURV4U/oybZkqxU/HB5X1Jh0b
vBj/z1AoJaQdeMEGkHrzP6RFCjdYzigbAKq4Af8yI8Z8xcFTsswq36tnuBekboaX
p7+rACmK3avAW10hYqW1rxZolSCJzOIUM+7Ro8+e8FDqGNPkw5Qai/nW0Yaee/W3
q+ukdAm+nZhXoOUs0uM7tpbD9GUStI+TYHF/PHLoc1wnnnb64lNIy0W5Akwc5z8P
nYUaekPbIHkDCUhyq2OhkPrL8EkIF1GYlWweOIf7yvAQvF/WO4sB1Bfs1VMy210r
5WZRKo+33yoZtZCRSEL7QWuxNxTBy4hJiTVlBvKpgZ5I08nXtJHcYEh/HiwR4J6r
/oj62mPtaJhIO9jXOkLwClbh+As844oO6N2C3NslvPBX0eOGAo2trlTTIb5WK7uE
l+BxyZuTT7sqF+xTxsu4jl2dEZYvOjSX7mjA43aNbAdMOFzg6dcFKerGWtupyU8Q
wiX+FrIjF83qr1yVlm9WghXaDRkwE8BiVnTKX+DWbXXTOfR0VUwwhLVRcDrR3pkX
ADiH0ZUuWNCkZcyow3CJGAHqIyuY1qoOl4+8hDjmP7lzNBC8rh0H81LW/lCD7Ceq
RhIqYr724cO+RjqkefbWUM0txOo9hiEa82xA2e/digbJd4pZixsYn5cn5wbjXoI4
AmysXQTcAWQrPiVBmEx5JSv0mEXgNzug9XwYXSdB0AhGqREl2VTH5m+8wET+dhiC
Wb2N/OtFpS58zpw/e06K2FKim/vFrf8UyABoMC+f+44FgHVciu7SpNa8i7MWwv32
C0F6IhH983KlxNixAIJN3D8Gh2z9hgwGjYtRUPYz9QIGIq/iR1LgqD9DbmdLLueY
ULRGV9W2y3I8V9eN5Uquu8AHrPyW5kp4DfRYlxeL1UE4INhzABEevYJWPqC4tbk+
mtS7eugifYx+elF94HVPZNGK+NLwOvSH0Alu6hBCwruRvujwzPKxZ03r367xN3yV
LWz/5AULXckTxp51p80REaCd/7ddPUuJTUhcwQg6RDXjBfbcmAApMnqbypXFvyuK
eBRggPLScAPC5kpQLFFhliDR9uGF5suZaxcnsURIdJh3WFU7kxqdJdS74C6Yp5uL
xL+RKq/fSsc9/HrdCZOEYEIsi7v5m58KmfdBB0d08f/U/6YtgcOTnlDuHsEQjebJ
BdLQnt7sg59CiWJ9zGkY8XxYQJUgalcyMCQS6DWM/J5DzPbmwXwN3dYfCKi6r16Q
Kup7lULF4Ifvfpy4JYfgV6bUBs95xi9zBaxirE9fdmmsp8ySaCDrfr0LD/JNkI+q
PzBBBwi8MWhnfqCniKfg3x+UT54UaCsGowpw9cMvJU6h1Sgq48VHVgodLvyos47h
GP973oWsSzNNF5xIyTz7yiEXYv+6w08bY0ERfb1GXqmfIsD/9X6sFiUEiEo/u2DN
kKa9gT519hUKuXffcjdJ4/8s4QYoDGEMDNnK8LgBD7OKNGCNiKD7E9qgy/NJn7vc
+eqIFATCwpDZjfATJfuNh4giEl6zbTs9CRv1+saypvviJMLCTfD62EtLG741Ng1R
JfnKZ+zMP/uMYm4kZ4NX5iI22s/igv5cxcbCKM5mh+Hf8EXWYCuCtdjrpqdXYgCr
cTSp51tt3AblciaU126jcjIeGRJnmrj/48149PtAccAYTOpw3NGqMHxtW4AkTqZw
d3gHTs0706yrKAXKt45izs+ZT9xEdrI5bV4vm5tMU5qWvYklPViWSbEnZ8MlXAi3
R6bbrRkFd1nfL+k1avvTymxGciHWKGUwv28MYInrakindSvyzRGumEkrZmqrL293
83irIGTk835u0z25WS+wOzzX5gQpqWGkMBACF/e8dRJ4uzFx1B5vb2MZiRWNcLtK
rfRYXUUjvfsA2QNhEtZw6bQcDHvAxK5PaHp1PqC0m6kl3qsMFQBSgX5nvPFvYZwY
aZCiXGMgytPT5gjfFVTu9ibDKpaoEZLA/F/1Q1rFsmauK0bFt0CLy+BlQTPff5Na
rdBR7ejD3QJNU22VjBS0AS+u+IGeHx3FEi+BSL8s4xQKpn3b0FlhDmQWWodrvMmQ
e0hKtbDKnnG0DrRmQd1qnPcBkOfscmNkEvrobXjcPu3Gd7o5bQg89K2oFLIbn2Ft
fZwqYzYU1Odr2127vLM66XhjM15WfV5/MiwXTpdPigWkiFzdYrHmnZ3zdwVT0VyZ
/PnLtj5d/zSCH/xD1mjWzGhnvX+fW3qEEA3eZ0UG0lwYc8orJIebW6bVOaCNtdW6
vNDbeJSRNkBNFVa/qVpWJUdxG8oGgauN8Oqc1e0yMvM3zRpHjiBVkv0RqYCEU8sZ
SS7TOmTJflFDeUC60hhZMd0eHIh0+myvdSdogd8ivvtU1ckyFXPYhfpv3qM0f3hQ
f2HNiSm43zbKTL46ckTLUfW7Lv5K2+hdgGTCQdJmdxQJTQPzat7xVgFy81WeHvyL
oTzFjNNSj9rrnBV1iUTaxF4KQ5AercSV+9Aqa/2vxjcwRW0OmN/WL8l4QcZv3WWf
if2yqpx2kAQDWUWptZXifcOumqTCRK2JE5ZBaUVvx1UobWChcZnJiNauxWUCQwL7
yYdU7dZHN/duQUCNjuknbJ95wvAdripP6vIKvtdlzlCwuKGos8A3tYLgozw1uDzJ
wgDohneMny/hJGDRJHsAyjtdx7F+Ue4RxH7xIFwWawhJMd+68PLHTshvujPVqp+K
afMbFt+CF9LfzSxtoWmSwwWYVAVSdg6GwvvlEf9ID0dgZfn+f49Plku+4v7XNNDW
iMVNuAiGMc6xNcFje9P0z39+q80CRPbf/4oOQiaTGblXGkAv2PDgX0czU8Pu92u0
1y8sITbkIWUEQSZ1MXkk3YDScAluLzulD2mLDgZw5sqrXNb2YBY5bqrMlbnoHO1u
mbTH6+U4G5c1lRI+8qyHYOCndj9Qq9+UrV3J6rSQvr/mXj+8or8b2YYGsahmxivp
5pNUjUO0F3M7EsOdd+lleNzRvPxn80A2wyxHwMix95BnP8wgvwiVOLD+KAnFstQD
Bg4xGbR2o5mQUjknBjKuFUyuKhbR9eb6fExWhE3MqjRXH+e+Xi245aYO6343aIFG
479djX01iJaCcjXJb53CndqtVJKfB6Q6HDgay++8OJl7pdmTkyZqjE/YPIuECJQD
RyDkLHWYE1Fdwzq7R+QAPmm2eQUDQKHzeZFfdgSss19yYw7DMOgg43M8kW4tyTZS
caUNsWFkgT2PJhbbhYmkHdsfdcmSxlwGpA9LIZSwnTB0JAxYGQ0RxzVIDuu7/8jN
yQ3RKimI/M41t0kWH6NoGeWMmprE+p+F+H1nsKgKwBi4HKMfnN0T2B/+h0FAVYbq
xAl1txnasvjOPrY5mSsY1AZcJ496U6Fr2BC0XfrOfnZgQbugPC9PjK1I8jCI7aWr
cy72uG3EbgC2e6TZakRR5rI1CAOOgUcgO3VTaCcfiypoNa5RzcKL7TQGDDGHSteI
+bWCY+Oj7M2YabGiqxNeNehZnVY6d7QQsiotFpqMFVFTNfGZ98hFcD/ECoovF6oO
AppE3sBn1CGdBZPuOjoAw2cinHHGc1nZtsty8DBuuTWkx3UIkqnl4EstT0irg/sm
jUCjBdP3yVpi8j/pCVNwke262Mgw+nPFj6diGPfI6emoI792U0+rKkFRbV7IelwI
tzj0C5ZZh/7COtTgwbX7hPKCMQPTEp6FDzN+h7jQkxj27G50r1ZBG8pFewpg73Lx
PaGTdjbx+erkruaNt9wU5zTUeyQh84JU+xezFa5IaDE8YaoLeso0dLYuXTmLi7dj
X01c3JUBFtVPJx+qyGzvwYjF4q+FDlJe29cl/obZv2uPwEeXSTUtRe9pyg2nuyMJ
MKIZ/hYgq1C4c+0UogO1yfhD41/OI+g835wgANhmMkH8uVqcH7DPV+fTaiKXKwAD
4cCkziQnmNtudsan8kNWYGJGf666wgxGsghwwpvjsS0ku/FXcNk89U6EcQiHXLnL
/JxhAIvwZR5GbQB06qw4hgmjuyV5Gp6nMCHdHBfwH4jsEl9M0PESp1xTCyRwnwWM
bdnSNzU1eGA/0HeseXaY+acU9D2UKk6DHp4IdnlMCBN0GT2/+mswzm0PLAqgR0Iw
oKh0Ryma+zHYpt+bfkHBTEHWJqy0G49QxPkxL57wOorIEV0gZAB7gCUUprds1bHI
84+90ITCMFOj/bD0/Ell/77k1n37a4UvClUZSQTUdMsJsAEg/NjXyDo6URko5Zf3
pzpwzx/goA2vpdH2IDnX9RuZmQXEtBbrOj4jhaVt2qZSfy7z92azpZEKzzcfli/n
TbeZse1uS6kbDWAsMuXeLp9qlI8kJ7ewEc+YrX2+2hURSHsLrDTU1+IIYVJLnZV/
bILi2EF8NM4MiQ4sLHQkUf6jUpGJNvNM0VcIIltASmg5EwX34TJGTRtxAmj5kuaq
53ipeK8cK1HQl9F07uDDm9Z/78t/AkVsnCdJhwNVsMURpzGaVgCOTneWvA2bCDZK
2hdBmeMLaEcTej6+3iw+7yNwhCD/TYMIq+0ivIWTEDMpRC3ZYC+OKyrZ521MICqt
AHviF5wvMPGQhsChG6Z+PMDT5ksW6WQkKIMbXjJ/BrRlfQmJI9n7xpFAQUkfCLv1
pouFC2/WRm3rgRJG4KfkZR9XXIbde7TWhjTBK0RbOu/qT4kfGKhtjDVQcD/SL/oN
VjqGT6YsTxyH7hNtqsDvR7kcv/ntJG7G9975jTg9Ufrm+JWZko58EIr8UV1YH51u
+YNq46NZGBk5bw9VbuH62RppwVgWv2SQw964dVZ5P37xFaRboDssDzp2OWd39Lft
VMuybk/VVJyeSn91kXAj2OIJPDld8/8DS0k9VTl4MO3Yq+pongJJ/BJi3LU07IQg
TleVE/sjndkiAXlVAR58n3tKxLJVsZJxj7/ahvDJv1iWqW10UujdiV99iPNtTtnS
RtUPFEAwL2ThWUfv1GRpSSvfTwgj+JlZDJT/vkvbQwx8Nqq9KzwOSihODOSRKxWf
5aLH0fEtHn8YsAt8Wv39aTJenGdE0L+5PY57O8a9/faV3nVz+S0PvEMbOOC63VWm
lSG0p84XAQMstgiHaEBion03d8AcJoTsamyP9IQEDUcU/EM1L7l6IkxMvl/RFSi9
LKmdWoeuJONRw5kfe6UT4B+qpfb+YK3tqbkWWXvezOhpFEV4Kqj6bShNdEXR17zS
xVs8w/mUpTWhFq7O7gCn10bsz6HyQaY8oQImSuVJR8bDx0wm3Q9t0sW16gyRMYMP
CBfXbCZ/siYgvuuHasDQwSELAL5A1VxwAPPwm1CHqKmpYj8Ay7NjG4/YPbOWea9u
ISjXnhl49VutvTSJltKteA7JmE8T4g4SJCCWhuSCeZK1Ad9Q3z1f2Rq/pjoYEVs5
qDNNj0MIyRMJPPPTfJj27QIUXQ780TmsIxkBWMSxfvC5qX4Mhpk96ZmMjD5seeY8
R/rJvej0gclg5of97bd8L2gdWjB5GQsiA+ewlCTN3qXPhog5xTAjJCZVxmWvK4UU
SjZJ/E07BYvHx/jgZVL2u8dwNcts0unGMQaH4C2cbHUETBqo/TXFtUbHRR32q7ww
Wmx3vI8dI48SvakXmLwOyMfIHuc640BEs16FLjMF9keNBs8KjSb8dWLs2d6y/VJ4
xQKDrudlwXN0dE4+SHm68Onk9AIwSp2yBqhoh75D0e+CzTFhCaZB4e9Nsu/dUi1s
cQnOun8DXZTYymaJaIEnp9rloBF2uIB6UCOiA1Lb9CxTOjqYW45neBKUtewPoOhL
H0/uHTAnV5MiE21A+bbBPr2djBPlgbWg2ughd3FPMTzZwXlIKgjISz6EAmEbpvA2
YptWK1Ar6OxwGyDiIIDDn9o5l5gR+8NIycoZWdUsG9jT6oGz1CRY7PA6iRumshz2
olR8Y8voo+F2huWw3tJFMgrSt8SuTaJ35sfwshkJrUY9ZZvRWgKhqazqO3mPu/df
IAheWQ7HiBHJSxBAbDAPsDoczWdmJGOL68tNMq9nQWVmcBRdnRVEGPJXuzEfnzoK
kPUKL8WGj2ocA+h112rd1UiA8bfxPmP2NV70r432pQYXHAArV1Z/u5rS3D3tZ46r
TOVIKprIf3KYml9s2T/LbukJgqwHb6m5QE2r4MECbkNiClU9tVHeLtJCvNGEBfUs
58D82HA8VI65EhaDaHX6Bf7iUWZa+3zQunAs92sptFrkCT9fFYP1Ol5/oHnjZMQe
Zu/5Y2OCg9+5ahBKlgmPUYlE9YKuBT6ncwhucsShP8vWWlBCVWVQpfeE9k5KycRq
/wQ/gPfXCdLiBRRRo33PVCYEYRQe+igPHfdVBbprDOeiy/lnZTTwYDtYgtO1xANV
8DzezTLFvg8Qzyk3pxm7fFnZGz2WbAvfV+BKWt284KByeKSVi2BesLZ8PylZHTwU
QDCdOKl4tgwXDvy5LIBwY63uwjSwsCvb5syL5oFockvmp5OATU1YMqTRjl1pSgwl
1jQnxF3vLuzfmY+qTngwG9LWE8vrTvPWenc4orowcP29H8yQd0fTKp0Zsf/dnAIv
O/EQBS8om3GiKidcYiBbXPSr9lx78Ew11o0+0YT4LhPA+sUa3gH3DIUySCBz1c/D
4U6YuvCLcVn7DJMbLUx/OrcR4Pl+ZbkN9+sa4u0lQ1pLIDtMLysDsu04AV1EROAx
Ca/q0Dycxl2eTe16ovUa46dp++RKzS6KIeTH6jMA2t8gRwT0DsHzwTUyElhiKnZq
ZLWYSg/r0SAXqMAKUu6Jjtr2a82MltG6am2+n+SGYGy+JT+X/bPhmUMaPgrKBaev
q+F3IBZmn+6wIITRPK8VVs3NpuI34Nt9tfdHivHKmY/62KgLnfTm3tAzF7xilhAA
m4thKTK0MdMFjYW9pTUjnzbOOscMndPA8dbmz5j7X7oxfH8d6OKVJtRH77zmBJkL
fpk8duZhBOgKSUBrKAVfX+AxR7cI96goms+tDL6pRQ/r1NMt1/hk0WRZMWv8B9A7
axKLeZnW7GlaTT5AeyDEs5Ad8NFYGdKPpdV7BI0mm6jKYryppgGz72pyqrcFaNbK
h97KWdBubeOLbVJkg3SCqc/582HyFDWIWWTnO/cCis+EvaJwaBrTVfg6BDPr3r/W
ECp2PwqU2TqriDdL2rMC8bmt0lal8CGpGwCeFwDq0x6PzqPxRj9JAmtjwQ8En6Le
r19Isi4IFrl63JyvNSvgrtD/96Pcf8fmOXb4lwX9EkbSZJMSaCcNhF0YyQQNyYNJ
HHO/wcdFlqcaG/y8f2RNi8C1t+uLkCEXYu06JYrIsWw6jw+emc3Mph+PAI2P1Cbz
SP7vD1xJnZRe9QshTajmpwAKj+XE1qqTzrcfHYJxoH5KXU/S1Stob4NqVLskqXVG
Dskj33QCq5rvAaNnOk3DBZr+Nqwnt52sZyhdKGR/p0u8i8iRD5QNoTbrIU5dFKEn
yQ0Fv2+o7l8SQAv37C1yGOCBvaKy9msmzVB81H2fiuH3bQoH6gJnLb+K8fZX5MiC
Hp2TPHJcAyvsRh6rESQFHcdsh5k6hNPXJg1fXQTFSDjiZV9EqTvlcZp92oJ76vv3
vy8q3oqkH04vaxO8R9zZRUI82d31+a/9ZzlaGmzCdt5qe+D0bmhBxxvkLS7fbhtr
3ehEm86xH91jLIfBQdI+7AbO9r+/HtQ+7Bz1LDt2827hq06VFTe3e6qWVaYpQ5ol
ERvBjlxTMVeeCaAo0Nb1HUOblC6luL5YdqPhhk5tE/Wr4oiu5YENfZaeEJ9WwVn4
/YISfVRJzO9T8meiB5scR4aP/3SgDGKrOFboedgQqEMzpKeGrKxPKsnxxpcDCPuu
qB271f0KwqaJ+ZwtRrqXXBatY5x4YbahZ02D67IYF/lsoilUeUFcSnpwuzKaheDU
dU7Fj4tTCzcH6S5LIJw4v96j5oW5UfDSEctCSYM7zPJbkWNwfEDpvTq7T6GhNPH4
k8zXH/Zl8FZZb8p60vdA+n9T6xRPnwYaet/wIZAYLyTLzV+9XQNnyPDPiyiOVawy
QtzJg5A3cldh9XxGG3Jgsgd6gCGeTWGJjwUszJ5+pRYhTMxs5atowJOKYFX+vl3+
+4IVNmmrFIOV6T5zwx/D16kTK7uelymyRwF0gwvgMSWwqMgkRNPO40XDvq3inXYo
OKgXXlhP6zymwRndb+osJZ3RaBKqrtTDQglVOrBgwyNq34Xbu8gUoFZVdyZ+GT5C
7nEICILFvwtciQEUfJM1/CSfOuckImfRxYkaa/okMU980WuOqUjwApWECmIdLJAS
AaiuUDx7+3Ur+mBWmYk6QUMpAZI+Xx8nuR5JLjvOTVxGDNV3ndiTPJOTp/zf5/Iv
3KFyYPJ5Td8EcwQ4lePnFlYDajMxg0zXjDLMIhi/woeubhfFaKY3MAiraZqFRWIh
SoawZNZBJ/ZHAFmlwuiXrbA5cO78uXxpGi9YNo8enM97S65hZUa5DVRekW8SY4hO
NtjoKmhx2rdaXhF4HR+WzElQJd8DS5WH9KenEqM8s5Wdw5FvnlIzkMrd4sCOo07P
MBeP8lmHT6wHaIWYwzhNMpGERWSDXll8Ep0rrQk27qscKdlCmKxBs1ACJ3/Nu1vu
hGS2LxfFeA0VqguR2zsoW3Z47FS05luj3X0gUwIQWqio7CkEt/VTIp0fxpwYVoD9
b16hzoMTFjfMA7WAyp2mUsf/nP8fRwmc5WFditftPKbhJm4rpRrBwM8A4H8SULj8
Pmh2t6S0/yEjqxmh2RvnbjRKtDnvC0AIHNzJcNNZ00ObdKx00/N4kxwK5xbBvZMv
1Ec7ZlrXj8JRI7GrQH7l4J1pA0I8A7gUIsL+jtJNHaz38wApQRw8FDMf6CCsGnSa
sGX6ezozrNHOg7YwGVxn5lbx6qLuTgQOAZvc9NlZj+4bCEUdz62mCgDwtw9MOgiz
KnhW5Tyh6mrCLUMppKGWDgRr79QnTK5r7pkILtBAyj0v30tGsvExr4TpXXAu5lqq
+jpGESlV0fJlRblJdQ2QsGFHzyAwBzeviQb97SQov0pBaiksJNfS/kszwWOLHjCR
19oV8waAH7c21sSSp1gu2Y4wX3PKoNlRcedkT+rUhv1SbolgKHPsMfE3S7Y2hDnO
eqxYdFW7I+eLWXvYg1+/Dsa/3mnHWXy7aCECCi8TWzBvNI7oWFkWBgF3cjDjWPqY
T75neB+9Gxn/MaCMoqLFnppDut+uOVXeDl2Z4Dee+VTcj840Uv+a8RHlu36W7qqR
UBmNEd+KYmfA2H+7YG7g8KmEPr428qbbUBiCTf7F+OHkcKdyKDH45qgmB7djcUom
r5IYfhZ7wcCyciY565IfVKCRAkbLUkDgtd6+QOHS4+/8MlVhD+LAZ+2JFpTUIqIQ
mLoc4K5xd9aMjd1gIxr+OxwN03fFuIh3X0B3ShtovI1cGyjR7obKP8mUJVTolLOw
zrutF+13ns043EhOJ6ke3/Gxe52K8cs7Z4jNJFgygp5hBEcSj6kpkXOs9H3vcGlj
8xScdhGG8OfVp6KVgJXeWYDtPv/qBfunCBg1mMz8mYVrBYAUbsiOcYSvA8NnM2WJ
zFPF1Q/yUqxpmMDNSXAKJrvCt0idKs7zgz4xFLn8rDfDfqaGbS6TvGcVvymak/IO
syauTZ90hABR+rb53+Rb/WBi2MKsGqj9W69FhVGGaST2LURd0Q7pNgCjp/sZVRok
y2i5M8eDlqGN8F9+3iRubkCkN2WLsqIcw23ayTE0cU8EeGfsisfTQSplc39JwHuT
goMZkpaoRvs0BaBrZQdB6qwboJyc9mpijbAuWwT5Dy+sqnAA/Jm6PhGxMj2U8Xox
R1BrsPETuROOO6XyNHt7xBVSGushn1jqG2tuMOJund7Yu+VYcEcUUBnpwP69Tx3h
t8W1TXy08iJjoM3nje776ondAgrGj6EaWps2SVgFX2zHZpsxh/5YKnMjUqubvRG0
d+RpFS8EWcFHSQ04rFGSxWUvH6zjRSbHpmP/xJ+/HubF8igalRfv3Di5capHhJbI
M2ULbJ7RJg0USsm4AdNjfLJiMU464OYOefz/BgArIqYgRCSez2/bW6T4cyujpfrl
6SqPXQrXr+PNnh0UUl5CU9bMSS2CjEyq5Z2DKnE2YF3No8os228eTz+CCaMb6VY7
o3OiMaHgcETZKgQFe0gQj8ilpuvjdSwwXWPN392ZdVvIBRD3t0N51IDA+wrVSiwm
yFYQC1EnY7DY6Rqp+MipziRtfU5y2NgREc9PuAhDbeAjZDrKeon3/2nuX4XIiqDd
0kNwWt27pbSSvJxUgnSsKqStBSdmjpa/dRzUgi51AKBLQkgDGVIvrchXKdXrFrxQ
mex0AB9hgczx2AARuA2ky94qeOxGqBcmAH9Sw19o/z1QUoUAIMeCizPvhL/K6xDS
IEi3mT591EvdR3IcxseHM9zgDRyWDaJ77bzNmzXugJRjd1ey0y0cXqvmXwgHHcZX
DVDbGDqFvd7avSMeNPrjA1IXKcSpWf/ibhbPyQe3fDutslj4TUD6iRolLdtKep1v
EG14BgolI9w4DDGvX4lOSi+fqS+Rzx/AGZpO5OjKQtJsXtEaLyRcDoWi57pkjQSX
A4BHhcnd1ejt6Mzfn4a8O9v0/lMWSuwIazbyMfKCPuVHkrYefZLbYebBbPqg7zjn
J5MHQcBguoGbz3/5eK4xP/vibDyrslwSv+NVXm06/rcswnhLa8whIxM67bMxmlzW
iSSAvQDNWAWmbBvYMYNncG+2swiffL6JM9C7XYI1PDiiDOsR6qQe/KFRBCzqQWub
GXRWp0J/KfJ0NxIi1O5iTBNKMsE6ZKgL54pIE1Jlek2tBhVm2MEJmqVTkNBjBqO5
iJuQkMrXeFgpJ7kjg1Ff2EIyePl4TScXxRm1koF7USBG/gLdCxdBfBcbIZ41fj+J
w1kb9PP7UZEiQeklpCjRCEfzmGwcmaKRzuthcFYdxHXWiXdErAu98l1G2+/8caXB
Js+T6Hltffw99A8iAZWc/SM+6LfLHNk/el56z2gZD5CXJFIWLa4CSMTY9/UdFyR0
Sgw4pe8hrXRJoL8xWEQslxNRL+4vgjE64/CUwVWqUknjHAjZtLwVz0BhcmzlMxRb
q9RiscSoFrEX+WVTI4HzqQUWRt4jjfAtbp90kqWE/V6ratXAZV4X6Tt0gL4qf7Ua
x607H1bJ4ddrfoBDftaEBhgPTM5q3aTiVtBYhhA9FbjOsFtqtWMPwlz1ra7olURl
EOiHSE5zGC02zglVNepsrBmbnJjR701Q85IGHA/yP+7iqviWDwNC2sc9Mw4fc1Wu
TNOWkFa4uumtcJnhS9mVEMjKtTanQbfsB1f1Mrq0ghITxsvikbwztLiEtiJGsIl3
ris/vEljtDkqjcA9DKSGvq0oGJd1jBfxsJuKBHZKaNGTLb2HG9c5el3gu+NQEYhU
5HqXWyWdWPHtmPKJOyiCdURvgVHl9lSzoCc9TCCU9oh19RU55YBsEKhEiNQyEW+V
NTuM+MIeDftmb0GOqRBamKGiUUHaaiAUwPpOKacDwC/+1IVJSoZekSWmqYiu+amG
gBXCjeqlvK4QWQKwCbin2ibIV9N3FW6KZr2pXOjUiSYjMJfC1YPBIxnN1+jNhXm4
McCyCUcyW7iiB6zfSSEQKzQkcaf4GqyUDVKXMiymuDTf0yeL6HWqnY4555+Bmw3M
2WFRhV9D4rMTSlJ90/N0qZsQwY47rgy7rsRLvKyL6PShXTs/7rWerNJUEdJVWZyx
JXgRYAflnUYU2e33vGo1tHeQZLLllJhtrFYzNK89mK4XBgPqmXFu0UNEVDCwkCHz
n/ua8R7ijpr3YhueAB4y7D7zGQOjAi/OS2YoXfS24M7MbTDNDznYuDMGNlazdEBu
faQySLoDoH/o2khtbOdnihagiH7C5PWZL8+vqiJJqCyTo4Na+OtTBQ0waRJTKzKZ
bskl3DZX5ohtDdXGgSPjFo3KzyxahW1hXbBxhsoOH6UJoAVcXCcWGySEkAbAco/f
0mZsGa9cRy4QnIYJSRngWXPCpOfdHfGzo3ImnwIxcv+eGn4nTq0pTpeRlQkvg4DT
SrtvoYz7RWx5gLAjIx3O48hLITDLKFUuqW1CKfODr6KI8KmKa1mxNSALDXhlwNS4
iUxCyrF+VoqN0eqYcRGxPsr6BYkUBcBX7AisvnELSZzI5lgnqCJczXBSJAqE0zoH
HB9jz2Czqg5D4+iu4hvS+9aye94O87H3Qy8u/spTdnn+My7UybfMaOcsuFzft49m
o1TOuL76/UA6gHpJRSwbPyN9VaDms3DGf8hjaxEhckWrj+IV8VnyMsHsgNosKtvK
RwNvUamhK53jjEd0XZuOwcDNWUPlvcoKKaW8IbWseNgU3C6rQmGJKltE6K+eppP4
diI3/Xs0hdAwWi1h5kvfnw3MHEywFOp0lQBzj1iPnyLj+D7gfpdu89WMPQIKSb09
WKJN5cXxtCSGP+R5pZYZ57mJWC54Nh9k4Mgup1MVbyjR+YUx6YSDXjnC66+qWOki
1hBn7P+tZcUs6oxUPvd5FrjUvCQgsgk5X34rH8XiXzMLkRcD87B98R/gYuzymhTZ
KIL1+TMlDLlIKEuMD5OopJ9Li6a+2QOstO4kfWnGkJ2jF3fJsSMC44rv1hCEE1L4
dl8b6P/f8FRKp5LkYfnRlaAWjt/PpWjdBrOU7wBqYssGU7DS2N0xbPW+d6U8vu0j
dP+7TphS617eFz2V+Qfyi4LYLm+1GXBkajsmj8Pum94qDHGYXwE8r+MQ7WIt0mDh
xXdvPL63GgAPWMGbUQafN3jybUiI/gL1r29Rqkvy1/yiLTPOTgTd7Is5N3KYO83U
svpX6eZ8Rsdbz3Hs5KO0xfzpJ39A2UpnggnSdvwxCwkEj+WufZjYHwu9Mgu74h1c
tYKKeD1/WECgLXuw7T1dDYE4M+8kWQbR/XO2QCziX8rGK9ALU3maVbxrXPxmvbOL
OlmiXi5nVVNPvFDU11Zr0GVncZfzYf16kft0Jalqw8SXjhIVAvWhzuCT9upDQGVT
zi6LueyPo2+h0eKk/9aVLRMGjYzd4Oih12HT2emFgC4/r4H+EAkBoNLSpl8LDgsI
g3yQLw8/rg52osgqM4TxcryMuwdZdqp9kyp9XIrcgM+TWcux236jRluObmRej1Mc
LFp3aFSI8mcQMvzX81xUMF5y/FndvdjdYYtHU3/ZP7GSppZ0T4guTiTbhC1vpu4G
jELYHm1kfF4PYJTBKewwqJRLYoCKtDCO7GRivZaq1GOyp5DNkB+kfO9xo2/6WV4L
gQxvJEW2gz7adQyRPSka3uiQSuXx4Rt4Yl7iTlbh1eyTEydLKhh28FxVJhIOroWs
DGLQYxlD5HC/7seg7lEqxIpTB8DXVKkib5JASTTid9Mfa7TDL1a7No/5+instn/G
TyordhuhOP+Zv1LjS3YQdxE3NkmUR2DtDJDY+sPeM1NUJZN7mxOF5KmnDw0hzxwK
MOg5qhls8qxQzQ8RCtDJue+Z6GEIIwtgZzhxAAZBZXRIEjzvQEeotNVJ/nhkSTja
gavG0EBGPeNjk8lhFYywVyPPysC8MYt22eQOHaNDZ0ri3Op7lQ/I57zLmZXv/c/R
4KwDQLsx3vItpczTU6ppkTxSL82YQEhbLSmMC02mA4zD3BoX/vapdJT7ExlnPcsO
L6TKUzPfSy17mwib+DJk2FXVOWrAp4Et54Ick3KDl6VCBfU4q8p1nouNsDG4lCH+
s5++1+t8BT5ZPzBDGnJK5HiZgXyDhsXaeee7vByE+DrZTka6qR61Ts/7jmRXDgHG
/igykRfKzhefV7ck+pI/fiuVvqv/q1mCVIIhKerxQGvIuEtwCH9xKW/qP13dUgnm
N6TxUjHy9MOBg1pqqyDb5y68WAnfhCYMjRd75B7umSp/qz5DO5zlnbEEaRPBgQsc
rXIXx2mxVfdc3RUUbhm7LRqIghHo3kqzu4GeBqW1nd4dYJpq9b9uEkw8NlZCMohk
jDoQyUX03r3UEWfvyScj+HDG8sNn1Z6yWmjOMXbrqKgFgdj1lkaMdaA/CzgB4VWw
SQHUIv9JMm31p0YifAB6iNFGNgora4HwmEdi3ZCVWz+sEZlxLmqfRVE9QGxhNgef
Z6g60ZUZt7oLXfH5KI9UQFLZlLw3Qe7lmaYX9wXAIhScFfdvaR3uplUMUW2G/f1j
5HEimOkzq4g4BOMeFZXuT7ZdH8OJVyMKiWQEEStJOCchn/I8KBwrb4oBGetUYluy
Y1Ztu3lin7IsaPGEEUpoVqGra4Yz3NSwTetLisXzj2Ts+1WOqbuoSugKSCu7ovzP
lXCK5drU2Zg/AKG2INw2xdOxlcfPIOr322Ed1KqePrI7Gxfgfsep8v+xYhuEvGj/
09/mtFqV/0I+qclW0fanfDw1x4IaOTw1DjBSgwzeflHjc0mAFxTZJqfYaIeeyEaT
n9EyEeYYOqKni6NKnjOZnKTP+FZ2vUsY07i2XlqTzbAzyZPlKYEqFsaqMuJU34Af
muagKvWs5FTiMGQ76R6gu6M7PMheh10AUV1kiXvm3YLJWQCDOpL54Y4kk4mUA+ko
DA21eO9Hf2170aIK5BsmDnS4u+H8+exybfVEP5Cwy+jZgZHouWfzPFwE0zNBCnms
SpemVwICWnebjwXg4emVxdzXL9q/EuBTMOOt+CgFrEKm5d8sFpH7LJCTYzYWbdSj
RZk2YoM1EEl8UqbDrusxsDdF5yaJAwzmRHBkvIOd6nEOE7hZf4jA6f4mV9FQ1Ov6
aNtJ5wYSuqGcgV3F30I6leYAOiiM3PF4LIQDZ9mog2uhsU7yvpP9huvRqBu4kg8Z
en6mEOF14uWyDODgFurbw7cBMwHUBprqwiu2Om7Boh/1ZBUY82/MhjkrZQ7lR9xh
xTGUJZnb04L+28NXI5hJoxFySBfMMyw+eYYgbbDUPdZNXcOmUrrYCwugkUQK0nhU
o8C6RDSwLvJ4S1q6rTohfsQ7mUWYNImwTErp9WzDyuyg9RkvBq33/abzncHsRfZr
zoH053rqCIJe1UL7Ffo7zzSMspFNsGHaHlzq8foP2u6CMqsQ7kEAjD44a8lnLIAt
sXq3bE2K5cSKJUoIWXr2jrd5pSjdSnOinUGABrCDWRp0Yg7dpx7mMptsCQ0cjLil
7nKKHSNWgDzH38jBpaa7oc5kXMPOufLeCLyDIuxarXIZCuVCbkWTIj+1zpFwC2us
oBn12jhKyxdcAz3fYQQ0RhSBQcFAbJH/xWD5cCEMijUzQq8u70AI3hPGcporkrF9
v2OCLl7cErgHOfWZJJ8XhMSm7XikGLsSdMV3zDSE3MYSbjDoy0AF4fPPY8fsNk9V
zuqN0cqP6IYghOazWiX8XvCc6w36ey/Yp/NMdG1UOjA1VZ2UXs2Texmx3eir5YVq
m8zVmfKz1kxUFaYYGkyaKFTzL5pgHftzqjLBOurgnIhoZYCQXkrYjsqFFPRBQxaN
ykDTu2GIFEK2nc1UZW1YXlqnnoOSDlIrNUdHH94gvVYeB2y4C57M0hRkJZWcshvv
b78WcGHVYn9/s7Jn5NfFsL/hcPq4kAF4yTB5hxLAcDsXffn/6WHIZuYNSwCrCy6j
U3BoP8oOXUmrmyuO6kyUmutrpAC5Ed/wUxPtcLZxjSL7NJobhcx2QIn/BLzgq4Zd
EnQItT/O23THN0e4wq79m7w8lo5TIDSBVuJvTLhWyCdoyeZ9Gy9zAB4UnlnEvdSJ
2QokNqcm5PVOUpugDdlBj8YPoJoXagfBD+S9FtcnaPfcQp7GB7R3/lHfxXH9Ms1+
BADNLiUwvNfSrBZ5yPbgKcwOgCFct//yN1qKNPKIfjYfe2NXN2YcPt1zba144AUv
O3JdRFSjT6zsCmUtN5KgWPvKHqCaF1oNMWkSb1qVUJ7LQ8ZXkaaAPRoj/eOQPIvt
htiN+/4+jwkO+dvPYIdbyDtoZyets+g35Nw8P9eYuY0YyN/oQzhLcsIc2ruyEauH
FKdFPpmLIC2EZ9oJgcDoc7u+mc2Y4/qzdpQDiK5Ecj9lyBGRoHMMQGG2LKXYaGFk
iHfV6Zm3Yhfo6NaKJ9qxuPs70qhyj+e5XRzJtrVd5t0EIvwox/m3YkRWQbI9Odik
XzqPxUQpfUTowAag/VECfb3eQ0sds1jCy6MXSbg+Dhr1ZS7dcYi3jVEVmrSUwN/z
AMbQZZ42EB7V28OTdNGqk2qlTSDBTVigWKH/oHUdfUaJ9ILMnHSJPPrt9rLqiudk
H9Nq82RWiAIt7vUvzRXDVlW5B3t+itC3X0snNv8LInbdDWhkxW+MsZ9vWSU1h3J5
9qm9aAKl6AaZMnwTD5GSdgbkrYh2yIvIBNBYUtTUS86Xfy01u5xAT+76m80wYpMp
c/eSRe9BukaflfS4qZSTvSYIZTATki0YOg1GulhWrAMWiNrhYSjW8I5fMGGPs62e
QY2ntpqZFsT1XP5PoCY+8UuRbI32gMb97JQ++DssYBNRWskJTgvxzoguC3iNcRbo
RM6+OsWPvfMaKOuIM0qX5f/0/4htBAOP4S/310tja/xCM70yrN9V25VKrE7Vj0yz
D6c1S4DJJ9AhFyeco4r92lFhG/BGHspSySBWq7+eTZYUU8w8PM0/aLaL2aq5uLf5
C2qCOO7fCBTHaGkRLYNp1Seq59EcH+Q0BCuWajau1apZQgLNLH7aQwb4JTrizDPA
kMNpN3RFEXS70ALEIFcEDA2NNoisV9k6PgQPwzBNaTTHoaOe/FSiNKfkOeOpJs7e
G4n23iod0P8wPpLDU+fqDGmrwftz00txgIXE4fFc9KkT/Dc8V5zZ/fBumEKW1Bzx
V36+Ac0Y9T0AeuYX+5VTbJ8GQfRCsi+S1gIVs0W3/ncgAQIr37CbEZQ+eWMTOz+V
gmnRxnCXew1fCUBw0OnQ0MBYjZSNtlkSJZgYUTqR9o4nvTPzgx2Skf3wLYgfRxiP
elkuzgU4yEQD9aDmuhgiy9RQurpQi9vguLR/+TAoMlIg4/x0HVSJDPRQouCsCqrI
+IiHn8VhlDvNW0sJxRUOixBcNUz9RZ74n8pk6iUt6wZNWY1JbTLn2sNW+um7LMx8
E1ROunr6uXI58FrKFrXU271WGid1jMZ8JrVmYQXbocIrCwRINHptZlfNiIb+ztgu
dSSQZY/uf9wO7Tem/kPx7lM8n3bGzC5iW2aYutC0tVW5VPdhHSmJRM1K7BwIjL2J
OhFOlBUytRHirchKX7RMyDlPdd8Km69DdH857CxnhHPfKFVsTQxsUW4b+QzX+seY
8Tol+4/yfslbO2QsPy1jU4+TGvR4rpdlvmb41zKtvXdC4iaaF2iAF21V4Rhjep7m
ay2yxOYO7QNVcU89PxqiRqSbNahqTTFDq8XzU1sIZXV9jwyqQn8FXqubS6XPVS5b
bd2GkY8UXigH9ejCXcsJYVtK/garDq1A9ln5C3KCXMjoX4vz0nrHlOWpSnoYDtDI
+Al4U/pdOlybt1qQ3rm/av5Nnu+X2KMxm07c4wC/N2306FpeQit9xjQckK6PP4df
e5KNSc5TwbTMnX52R0oIFL5ij4TvDBuBe7perh0lYAgo9ipILskp210nEMtGWxTa
PKC3nbDmtyFquYwz2i1n0xHEAOOTEoSmp6hDvmOc2I2mZSaeak2tbnamU0K4y0zi
iQSRhzGdkk0pd7r7wwn9smxLts0dpFRQ5HM7xStK809AhLl4KGYOG27Fq6+6rpdW
NlMBKwkTK5h6m3UE1zuM1Kmh2rmF9cci2V3ew6wGhouEi2CJ9QdSWX9i9+X6Nomt
22OI8i3zt86eqcXkFq6fNTpzhciBUEmqZQC3yfExJGLVGhbx4Wzzl28tpR+yi1U6
5fMToBLASxWMKwbVEoe03GsbrxagpzURKHNP+r6X62UbHF9bzF/Js0qfbu4UlPWg
wH4NrZIzeqVQXEn4/VabNUrSeNszk2htx9+V0tus3ZNbNxgTyB1a/qDHQjdyxbzi
xczk7fOdrRCMtifR773hbSuheujwkT4ywCoqHk576wyr3dXTqGZinRn8EvEjGqD1
JkBs3oblrRh+vHV7qRjAgXFs4GkXIs5QlDfHqpxhaq/GkXptRK7JUY1DP1p5HfGP
iWxwDQUNaMb54Pg3J+OljWZCgioH0S3AAVXQZ6SfBnG+XFjmBMwF9QKju2C94ok7
ZensJwCbYxNOV1jQJIEwJT41vWrvjUX5A5WNpmlX0/aAsM1o3eoxc6bweqAsbaRG
kEuE5WLS/hP+4RalY8waf6vJ7p4g6SkyJmibNFlo7zc9ulI72PbAsExSmWu/JtIb
gAr7SfNIAneMxIFOR0CqNu2HXjvwdd0LqM4v5Onb63SeWhOjdxS7dB7/nbnKWXmD
L0codwWXxCSCDZreuJD81rDQoCJHKI5mpu0KuWMoB5S3rv+XUmVf1GuZPHoaWekf
I2+NV12aw98QZo1aHaDUhCEnczhgQpnAMB/zw1WOUFCGTyAjQilvUP42cH9kVKfs
r9PUBAF3TCvWVtBqPYb0iKvaD7aetQ/C8f1YkfGTVRdIdxgeaMkeFtKBwoQbaO+5
V1c6nIsFmvAmkOCV3up/xS08dZ1ieR1+RHz1LWBh2msxUKOmeM0dLC3b01QgPGCb
E0id1wIvWrBjWy3qpFiiwFNWEY+kPP3XGHYxsrl+x9iykfI4rmzNPxbfx++/L1Y0
QTslqfCMhlDLnhUcbcOad/oDhKofdk2mv9i+zgMDlWi2/1l87EFEWNUrbQDcLFyc
7HZFk9TFwCNd1HtNUFSlpJOs2of1OEoAkrc1S3kXBxqNlXyQPx62w+UimIAT9/em
g1bqhHZiC1eqp46BOOATAHP07PRQReLKV/JBnsoqfr6leIMxITMEKfvoTHxV/tf1
1wBd1on3iZg7k/z9zNRrbxEmb73fFqsGu3w4XT2AruXP7lgaNK2bQJSCIJNOuQrZ
FLKkW3kWJz+KrskfDxXbGz/0f4/y2xTIFqSjrS+otmGEEP5AeDojF72osm/TwanC
foGQk1eiwgAxfP4hhhSWWGne9QGSKVsc+7VM2ANym3KGSqeg+n5dLFp+0mYzvacT
We+FeRyU0+OvHGaJ+irloaYXvH/+ypcZgPKRHkp+ICjrzz5kKgWtVVkCFQRrz/5i
DkKXseEdLpH1I6MrTPkPQNboJ3A+P20AcJvvQOqXdqrUgAR9x86emrLdFCx7wxMZ
WTQ6rPa1mSpvY5W7svaEEZs5RESue5+fRrhnuyH090ibH6VCrT2wBiBoqROVsDTq
0OODuUZFPUQ8BHnPtcMeBIjpvzBokNJVmEaE4dhUmvYpgMZxUbwdIyMh1XvxZPvy
QOkFwZciitKr3etWGt2vkCMPSzN+32/vStUIo6ZErLZcp4NstA04IcEhieiBkjaB
VlfuEAwB9eTVuh1txIbwGb9OAaMk173vCOxXqrTc4VYMAcczP/Nbs0DaD76hLIic
gnT1bI0+0DlEWg8ZrXjtBBdN96acSKS1QPGtx4AgsuVa759T/ngeXRQgVOEFKh9k
CEFGb2yYIN9Drw0E2wFwPG0DqGzkTFMdjU7Xuc/pRow2cggBAa2NY/yllp5GNX7+
LLiZCd9N/3Zifp8J2CrJ3f+vBguqsHInysDR/ih9xByxT2+L9RibLizNQj3P83LX
XMkwJIZI2hr/SNBDay85hIiPPFKwK1xJvC7erPByk47ktZ+aWXHbSgU65OtRTUOC
PHAyRDUsa1XoiZpV8WAB1YIz516mpg18Bns2wEXaZfbbJ8Yum4QV/6efhGmiWjwc
Ol2XHzSKBVJbu+9I17SJzEt06wifByyViQjE/02FabT6S/yx0beZrJT9bDYW5JmX
96NrKjtChgDNlCu5nLhzMdgVJi+pNwkYOZUHK7Ek9+ZOhk1liAXrVk2PZbGUuALH
YyDIG5mjM2KnYUKt0nFjaVRQGlECak6yXg1yx28fc8FOh4IuCKWYtHceoN9g0Z3a
wrF0k1Wa+QIaOEIz5omL3RCrwegge9vjUf8kD6jjAoaNyYr7kUe2xSX5UhvWrsuZ
BJQdnEYCvLii3gI6Tz6q5LM9F7oa6PApHBOvRodJAwYFAQVT2aFF065kfh9J5nlg
0PAtaQDgdsyOKuT15tDeCqYTzhPbQjxTWDe9/lgB9NE7f7lp0eqExjhjAmICTgt5
LaOw9C37EMvuaEMAWjYG8uneM+FNg2o6OISnwpEjVnsCylL86HGkoHp8dxX26j/P
CCXD/tfFdOYDeo0l1xhI6LgRDGCzD00NNJAtS4zIL7wk9AFP52symxoLxlw/nXO0
axvZfeKaDVkGDFe54KKpVVKnyTP+TqdQVfrbVwgLbVd1zBLpe8bTjpMzcuTOf3IJ
H9nBcI3Wx69zfrhyz90r/n550561lCsWEJLkhchMqe0HnKIE7CFVhVInzkB0WjU1
qdfBYQKFSWcCjx7wO1PI/HbzBXdWCPdgLRb3qC46tmB613hoKYYpdRoVVpbKDuxR
KNSSW0h5ice4KWEJFycVKLauScbENhMmi/qtryUivHtKXz1Onqp0HJTbUPNOU71G
kTjakw5uUREWanjhERQPD3arJIPkCoFswj14o6ALpPVXJezwMU4zkjhPuxtdrheM
EerKbpIkEd0n2hezJIv+wPVa+o406s4E5ifomECCjIqUWXjmlbVSZuqVQ9ZEcAUP
jnDPZeyfZWYsMswr2C3b0T/e/D3mDV6ie6kL77rJb02spAY6lwV3LILLiWlIgXdk
ZPuAxPvrVSX9vMsruHRQptq+V8VA5yTEJLzN+SDuY1xSca34HY0lBXELCzv/skHj
qjNIVjPnMyHS/5OPZ0lld3KG5y+qSLkNhzFscRtzq2tohn+duGf1gZU0OO8vdDMM
q7z5YvoyOsI7LnEmgPGrYX7eXziPHZ0CVqd3xcYeqaVFmuB3JPK/cboAheZvCulk
b7MXR8jGoBzWZxuUcUF+GC975NZ9UqdaZpd/cqSJTHgf/sjlAwWg+1GDou3Iy2Tg
IL7C8ArNmTxSNJ7bU2F1fGvMzRRd8Zom+ogjKMSoLiix3f2wQ0KavGmoSZG8r+kV
pLb++UWSfMLYoXm36vv+R+KaAidTEWnYrA9+UgFl32zy3ulKr5b8YAQ07de1KnEn
av119S4ONjNgjtjBpKuxd8xnpiCYBFRkLBsl6J2ZfZaCyFh5zyAN+/LZLTUchsw2
Ix6e0SmUIUcg0wAlzyBmXbowMVOsXu7ddyTG+/fTTQfi3otigdyo0FGgcG2QjLju
TRRQPeh3D8GjNH+n8PyWbW88icp8QgAZHIoRTm2Ln6Y/In3796XlC13sOXssOiek
zEfsVD1HS5OkmkQbTpP+JuHS5itT+ghygaFoU3HMXPLtlrHmDFx+391utl2Gzrcw
FP1YSNvi2C3aDwv+kiM6f3em7kPtuBqxRgSOfYtHZ2QVQyeDYONLep/De6HSTIY6
GuZrz4x9ku6rSeJWiBydsOGGmwVNy2pSxgYzjgI6JR5hYl822iZRhTCHt57Hyyjb
fgYgnaPhZO7ZNEFqglU1F2HxE2f6w7OSFQFozlbWRYZXSabdVLtqjxhFp2qgVb9b
oVvRRvGkdZsEUjfGrfTJThF5rsiPMGxlRQDLOKDpJzy6Wm/1hxuqoiBegFT8MYrB
TH/LJI+2QE9F99Z50p/o4GXHIa2RKnuNnQ9qCJ+EH0zORBxcNwhbKAEoaCx24Thw
3z6xH0ONcsrGHBt+K340Opnkxu/cffEq/Cke9zWWtPI/T+j8un1ztp3rRydQJbEK
SWkiW7npWJqUbG5tgvfOqqHMDHzbWSY36UA+XRlDWy7jt03A5E5O04jclZwTSqKy
T1W1p+z3Go6dP0vS5fwfrXz0fK2hRxazqbJPjAX1bCzQWdiL1+oMV3lcK3uwzPB4
KQtwIwozQTczZXDFgCqAeuqnXAehpBeT39AFE2s88+5QXsS01Qzmz3zE1BEpINXL
kguZvzBdGbKMpqn2iTCse4dpxS8Y7pj7R8kkcl4kZCfmrqoyAJ84SG4b+vn53+jD
7ZbMfqUooutTXH0ImSWnd5NTbM6gc0Ak8S7YEvb5q01tpclKSMXU1MeLHmlaISlj
1X8tewJDGyWyigmZWIe4f6SsNJ7h0EGoNXsAdgsrJkM4l60yY7aJmaIJIisHmLWo
hRejTG7eeWwBk/Bsjk9R8fGhYe87ALE5AQljLSnRnOwdrHhRBRR8vSxJ5v03cBKO
ENZgNO2KqoYl4pJfhzZ5+YMKTM1PQZKJnVtfSqJcO3EQv0lM177oMgd3bJ5/b0mK
yTGb90w43n/f+FuT9/YfgWTTu0O9vAikOn7SwvvM+9MyxqXopI++O+pFERgLJxlL
veYzCDTo0weUrtyfTacxke1poePAqEVb/u76jygt9Yg3OjRbSvTjwnsXK5sF9Hvy
Rz9K+RRBu8SEB5h5ccTBbUZHUQNSIxVrPWY5nj4JyVDFTsPnI9ZAbK7Rc/iBwFas
CKn2efm79tMTcd4LdL9SZMzTsGuCEIpaqN9QkiyoBvuK7i7BPkixF1B1gkDNCmV8
u2tBtOkB6/kFeS4AKR9YGYUCty1RQJ8CbByCcmGtbEHCePNd65eF7o2nP6vZx1UF
a1EkxIIzeDr3RkoMVBhmOlwYj0SqzsAv3uIjRzTtRnY3KlrPilstDnyn1mvFzlpi
JhD41M2fb2LeRItiWEBY84gNXIwz0PVWScBiQv6NDVtAXfj+nhKYuS0vdcz2XGQm
0wXzaQbgwVXmf6Lz1raB+6z/HjHp7AAj6kzEtr4zPTwp5EEUvQqYZMdd2kj9MmG0
pKz4j8FEAxpMgH8kV5bRu+ldkg01TjK/Rnma7qMQSuzh1ir+1xFhNaUadXUMskTP
dLiA7yfGJeUnlrjZH6iUu8vaXQmdcewjeA9TBvW9kBD6j1Y/UDDb7YvE/Um5jCP3
1HifUWn+1/+YLmYdWFDFHtfMZ06R+nOVUJ/b5ltKJuj+AdRRooZFSkeWkgdq0WjU
+E+CD4CD6UAIKe7g+ZNgZB3328bTQHtk28MRv73aVlFLdT75jQWhFCc+0WZyakRZ
/xdnSsVIT+fut7wHHVQCeBoy81vZf51eQPFfj8m1M/GVodwK5yM8JdmfbUSTOrk+
uynVMjNZqeOmvKwOoZIE+ivHQy6tlaDakrh3WPtRtreXVMb5DMfftAxsqvtwjrYg
8+0kghSjOvDUaMrmw1d7Iwwpp7GUIl0XueKTfR6Koor1Mr/rbLX1Ad/A3PFIBYHM
EgtqnYc9X0tXn2/+t3XF5dJ8nncMvKW81ZuAYjdj5d/B95m+ylZN6EcaYJPKHcEL
/4dZiBDNedKuwhijhDwC5Tuq5OpuDd6qruW6B9dipHlXYtDYLik7YBSR3pGjsoLH
WGoxctrki5Y0hVtAydnapVxdoDVPTaZ9S9ttJeWHEnnZLGw2l/nQULbp9nANwyPj
WX2ZJxFMPczWiGD7bBCPmHbG2T5uNeB2mqNxPIM7PhYrU1+rvCq4RVBgbzvCY1Ha
vbgDcByR/lH1WriWv5LkBuhwINwVOuGGah6c31e0ugDmx7zS+39rvWRQ4EkysJNL
KK6wtqIBoZp0gtPp9DvyRuEJ7X0BigN05Z5pFAt2BNrvWZ/mH9ck02fMl6klzwOW
D14FoeoV18/sAIkT/KiXFF/D/tEQEZYor3R4z2ZKMvEKuorTOP2rQXnao/nMT9vE
T/SXjYMdWIK//P98Re88Tt6i4+yRzRuhhrVK2jCKdzWEKv8X8mRHZxJGF5s9zRi2
ivr1hCeWA7hbsU8XowkKSH3KFh4XLFx5M32eESEbsMUG1IYmtLhwowFbOOW+SaLm
4i7ek+a1rrZEf6vquZq3vyvXsYtyHExi/SfWjOm/Nek+DApggv6qrOdu9QhUOCKK
rz9TDwZ3uMMVWGNtAK28iKUeRVpgfCTsXYIJg4bKjkaM7CdgwChAFq4zsWH+36m1
Z0luoc1AYjg27P3uGsRC/b07sCR6z0Wt1YFwVlo/ufSJKRzIBM/jeimpBJ6ny6F2
RIabSx5Ewa37saCllZJ9punNT9Vb/50g5OUdZIvpTFQhB4kvlqCrfu2YF0P4HMcO
ufnPBxmFNJj9bcb8qz3XGH99hI4B1EkhH4TTSJlQNZVuprngtXCsMPj8GxCUuyR6
lA778MtynaQRLawxobEvp6Rf8zWJyy6ytgw71+kQhafNNjvpcTUT3mmnTBk2yqCu
tJZtqDd7p8BKsIWg6Sh6ztDJcyKSB/oi9PBgPSVjm1A03ufz4gRlCmHT0hdCQiAv
iO+noEBAnXAIZfSR/n98kK1cI6FQwMa0BC4Jb0d39ZL8AoK2PkECEZAkwxmP0uTV
ixgUDXpV26fFTu35QUQYK5SyW+AqktDw32tdl8J1r/1midXO/L5a2LiuFm/a3+b8
6SCjmAEjpKSfWqDP1UU13gIKRf9FTvk52951VtbBeh/7UkuqmVOaeunY7MY5fREb
xaYx7HwbvsHBq3MH17Am4n3xp0/uexDs+WNqt+2i+WrXxh3K29RKIrgTTGty+2wd
dkawCOuqPUZ/LS7MO/zK3Me8tjYvDoJy3Ye1HKB9SYn4a++0Pc8xCRXP8TZ9V1dJ
wAZVh9amP6DGX34JYHU7lJ1JBQTCGb1nfaF8cL4bAh2V6OLhcmivyzcv2oAxORKN
7I+99+tgy0tbM8W1MrRHjbrxzoyCmd5Sc+qdA8nbXbMN9aZ/wtxhsOxg1T8KEN6K
qlzm67wuWTFRCe4X+riPOhhSwjncyOca+bICrGeRAkVAExpWL8Uy3w5kBb4ilwd+
UHFED76vOv5sLmVTSSSt8x1dYx6X+7ABPLDKoKnXyYVelO2RNf05auryFnEF6wna
7MUhufn/FyfIU1CxN+d2zic2oLjclVYAJudGaVuq7wtOxIawaoGZW49xwVNPTN2x
MQszJQgthANT3hUkSlqb1yuf9l5mqevHhJDcVskvJBm3IwgY90D8Q8YrNaLpgDye
v2NBJqvJTxA3JBovvjFJICDyf1kAu4OMlsq+FxqMa6BzYd3ZCHxV5jtWxug2CA5K
q8XVuYUcFfTfkg5GmZdf9Gy/vVy9sqDYeVPWTOddw3VU1ClXJCmG9NU+21/CaQB7
szKe/Ao4GB7hySk7wRaT1dweqQ3Flwc7cHZ5Kvg1sgOjHT0gKJFdhe0ICn0MYtTW
HRpkf0Gx7mDjO1iJkJYf6KXFvIr/OxvPVbCKfpCgBv27PFurKcbm1DmPNc0xn0Zo
huPDZC8dgIwA5YWmJdqeoyoiCv1M6lHjLqYWTce+MW8Nwexy/vMvqytEA95Dyo15
mEKFFj1rP7gNWwO/VuRDps3CK4oB8CBri5mbs8Y8qCP/Kj2QIkr9BUQlUmC1SUxT
1XlBIaqXl7FGJVCTUnIWtkKLFDwyYjrHvW+vUnOtOEbg4OPV30NHAG1GR2tAkg+s
CkxxPGro81gUdce0Q8fllirUFbo2RZ7kltTDgsu3IXJrGAA6+vJQrgHGa22J8dA8
PXKJElc6RZzc6iaRV4/v0ubNSi5XnyzhUlZsXKCjLgnqxd/ucsiV3MLf3SgBzEoq
rKJdSdnK7nAHZE16hKHEHg5dtj7Q7I96FnRL3EGxOeYIw95EsWDvUAYSK1AIm4Dv
9Vyxar3gqB1/Yp4oJU/QN8s0MCZuhMWH+KBivn4trgbPgIXxim0qDWf/TN/cfSVa
p/xqxSKwpw0vCho2eqQMbFL8tqiCm+pDsHkco3IYr0xAKSDmNtQ4aJUo6qzvSNTE
v2NFniE2eO/po+cDnTQ2tjYxO463ifkWgtGUdqj7vOPb0Z/fA/ebTZMywS/wGv/X
9pO+yN1r8T/7HURVWP4LVoQpvBKuOQGdIxGDbicquvGiJFnIZj8lkbmDf/NyKntM
HnRqT/twoxjDyshFSMdEM/ozYeishu4myWrrkgKqEpOL+ap4Ll37usINS2gGp6KN
wB7eW6HavzZAG3M43LFGV7K5fPJseBAePfhpvNsGqFtRpSzRIP0vlZqvPEHPcohV
uvonks6cuwwJ8PqgGoPvGkWJlTe6UhYTrD+fpjBFC0C7LnCnK9qCHD3JNyCVZT91
BLcAQg0NU5I7TZDB5vVqLV6E7+Gp3Vm6QPfPT0xnTnpdSj401rJMkDbLF+lG0iVy
XqKBraA/hf3CStA2fLu5PpGlJ0pTNYVo8Cg9B9aMnqEI4f01IIRiJvkhaZamLxXQ
CH+atSTQpQA5Fznxd6GZ5Wf0/jFw1LMmwwCrGzq+G/auInxYiiAjP4XK5stdov5u
4SUT39sPDlyybTtzsdXsgwEbFn0T8Jln7LfH4bCcHI7NUbO+uG9cXRPQJMlBm0l0
xYm5ROoeetLGSZs0FpHN2S2/g9mLlSF7j8PinBBalhXW0ApEOae75ivLZD87HqMR
/fnvyCEJUIGyFGjtKmPiCkEo0pq93CrYDLFEYOleZTbTQw6ozSWcSwsC/9s2tQ0G
qrkjTvFCg9FxFlk81yaX/sQbemeXX3rHPzVVJTrHsoc8q6ICQT7lS2XEwHL/z9k5
OJmpK/LAwPkh4IfccPSAAxzsgIKtUlZxH50shXYoIEBTcEPP2+pMPLj1MKgVnxlA
jFuxxNqi0wiLPZrXgHANS+khipx9j53PV7gjs9RiqD3RionSX1TAxJyGyOM3Pgjf
jEpNmMLSQNRI+qOXEthGttDXMDtfzv8IMet3PYc+mP5pFEyRPogAEcJSxEK+YDa/
kM3Ca25fPRDtFvZ9gJzMWOTvUTUt7391oBjGvAauwcbrBnbFmFhLA9oOqtCJrPpM
rrKOJIZCb4+R89+/TOpUPYbDWVRN5UI7WF+0H0ZzlFIq9J9qKT/U67ENTfATEvTx
EKK7SL+rFeI/vjDqIzILp5RDbdlqWqIpKd3vBbmWJgTABqdiy1rjXQji3OFDhXw5
/PiL99jKf3Te3r4IZIMw1TpPNTz0iDTYpccKcG8Sy+EcXJD84dIlDXwYqphugrVC
cjvAoI8fBtpat5OBIwmc2ivfRXRD0kS4IvYlCdKgPZmamyZ9A89SuRHZPzUImWqT
kz9o3Qtl99kYKFdEwCWG1RYzichfY/UkmZ0N24noxIrnBisjSua/Vp3KVaI/+T8E
0+uogKtDy3lA5NM1acMaLy+9hZxxOGq+PwipN/zQbeTXoP+YVYmEscVUmf/Q9Bq8
llWIXfvYcLZV1v5fGsbY9kUPVDi6RYmTFbhTRdrN6FD5rpwCHeOJrDscIQt5QIro
AHVGGtiRRYzwcK4qR/jvU1z6w01xQrNqNTa2RDtRjIV6y22e+xhsasUOn+fdqOxq
3re1pYqxbK3QswSzRHizKxI+Ze55d7OfYbeBC/81y/njruX/+0WONxap7f+SSUIP
rc8LJoBRTmR9TY1THubIAoFHtxQ27vVhZoD0IW3W6zk3icB7xo6KywuI2afEpp+d
OCoP2a8sL9kXuIIcNji4UFFgcGckPw+Myy0PA0SlmBt5f0T/TemHGRaR/XO1LCkD
XeP+1spqZRfEF4bOWho5+vdaD91z2mMAm5fNm33s16AAA7j9k1mgmTCoi5+mT35E
iex0ZsMG62k5V0mgg1sLgDNc6tSbTDoTgAkkM8HVPMGQJTXRQTQbS7U9sMXol6Dh
41QtP746NX/FmHAsceHxyUC+ENDXIi8ig/BUwv9wE4vd+u9uPytA4W0EHmQZIPau
Xns2P1t0s8YHxnkewDMzCMPk8QdDp7D1u3g5b1EudCbZU5mQrw9o95nMBm5Rm4l1
IySExftOMQ5+gMER+OowuSozpfa/kWBGLHwx5jOdsr5HVP4WVRaBDaqYKp0haU2y
I2/aqSlVS5S2iWLh5F8RUrZEd+IYXpLQSOi7lpHWOLqRw4Ws8hdVpMSHkl5GSsCT
g6Wrdj1mV6vPdDEE2AxRxtBSjYJZ9QmlmhT7JS+E7JPA8MP6IjBybgYBbSElJfIk
+3o01+1VrAEO70xGOhUcm3uezNMuHTLqba4+X/K9BxGjcNxJ+NHo15qr/qVD2VYA
d9vXjbSWppz+LDiS36MkjPbQDTrGnxFun1Ud2lCzQ4gkbPHguwfPv+oyEFXostES
bTZzPoOThVMyFSPoHnPFc0XFmsqr0H+VIo1uLslpuudcF9UH3BG2qAkk0ujqfNDA
5h2qwxzWmn3CZu567bHHtqD+cq2ZblJvUniCirssOnBaF87t5xfYq0Kqy6CWyEAu
mg6x3Cbeth9H2MDEICJ/tFakfc3lPhStZR5Hre+mtG6pc9bzLPU8nSBvfv2n5TAs
Uu2wlKhqJ18C4CFryh0gYWBcil33qe/zUSWjMjJZY5FUgUXAcueAHGiiDFEGrOOY
jq0W0h0wkspiBCbtJiGDi07tgxG39ASazKzzP72t+v3ojg1FxkB8QV92W/z8EmZP
l8s+hIqYVGz9IQZiGGLuNjBiEn0B4Cx7xZHi5GUj5kXnH5Sg/bNza3LrdKHHKpTl
hMuczW7ogynj2kFhyZt5Jw0WrBe/7+eZfg81E7hArs/djuqSPiag9sqxTuyVujxY
p00ve82R0mcWzAwzf+sqkpwJ+p2tA4UXymQwO8HPMaRoMoptscaUVTZIYV69oJ3B
+TeZBXW0EWiec9ax2VWdw0l12UoCfHt3LuBQGzpGtfC9Fe6pctx+r0Y1l4zeiBeh
sq9AMOqrOHYntpj2zMuHIdnhNRUQqlIev1dHXd5kR9HIAh+8zPTbDnJjnT2SYHVc
mSm+byJxfmWHnmdZGxscO+onNH5UQgcZTRFOP+Zs2CzFq0GVRURiL6Xgfk1hMEJD
5sQXQU1QGODYr7+r6+3SUTWRWZ9cgsNaf2GJ8tz0B8Gi05LMCzUrqnXgGnEjwRnd
uGtZStSqajCjvzBd3K8G6CVm2LEGt5K/7e9+yzSPMmhwx7VgaAIznn4ErPL+oiFo
gQigf2Vr6RbW/5dO5EPcO50selnavpbGvk/IEBeC41Bjd9AgI81Q2kRXvEATk30C
2HUNlQh6kGh2EcGLmM5XypSsytbNCE2T26CzUq4+rRKeyJFE8net1DWDh5Lg6jyf
2s7ZxLm9PWxBDddJLQBqu1qqpPQK3ihiDhUuYmW/d3St5cPgAghOkecESp66WEh4
y3D6D/VqRgG3e351+1Vf9TXmLxWgMuzz5tSdZafLtO4bJYqox+nxqFa6dN644R/k
0cPP7WICoweGRWAn2sUiyolWveFNr4Q5WtZFnxJi6p52vLoZmv11tZ2w60mdYRWT
hdq8xeCCrWGBO0nq/CL7yzRWBBnA7pfY9vemN6D4G9FH59np378SEABMQoKF5L74
KSo/UL8j1SRSSZKOT+9cDW76aeFBknUUVUaPVsNBZDCcTPVeCDqwSfUQ8Ue79YZl
zb6mmLrdSM5vvrJGlodF9cTjMzhbRND2l70+rCd2Rh0t2jKsqdBhObUzl732mPfz
u9/aoMkoOt1Q4GRJ/nTaxwGJHRJrdrA84TLcSUmu7IvRS25qZnPFYenBhyZNpv8V
D6S00V5VYBBzpnPbFYmjzejAZt6y0eCx+o4WRJk2rRtwbk18rIMpe3dneyz7Kruv
NZDD/F0QZmV1D4F2GUYM2Z9NNU4XIHiLeBMskQSE/m3KucwvpT3ape9wFawVpp62
LxslcZZWnUQL5AnAIo4/rgJYLqHF9G4q9GHS2ByKnSmjigycz/nx2JSFO9yaGofF
VPdhPNQ1CVQW/w5AleUCt677I7OFYeTlWEuLz2bfUCPu5WjGh/IAGVsEU5tBaEN+
IiFygtdrZNAo1zKU7qijGsPqAriukwTypti4LlouXsAef98S9w8wpimDNA6Qjlks
hsItY96IUFTogAnICyGca+ts1bsTPxjoppOvNbF8B9yGpiikoGuSzGRWXPxGR7Hy
2o1tEN924tS/SZP645s6LS+ZZVVi/ZcKcjRQXF/FmDPW19IsNV6m7P6QD1TVh5cm
IerZLZ6APzPoEt9ERYUc8aZ8b0bYm2xhsZYLoahzH9RtmjhupZM0rvcLbH+igJh3
JXq7OKOwdKa4+/rLwF5oFPXg/nhjdziDHBe/cXWjxkYtA671zfaJ2hQdceFNH+8X
L/CpLHYPs1hwC+oyyKc7wQYKj7v5nxVUY1jiqTwhUXGxaKhlrxebn5vy2XgXbRor
kcE5ZP33ShXtiJEMNfncAFBxYGKSqdqnCAve3Kj33K32ccu228zj+vp6sI0uGwT/
oUOxdlM9gybydSsosQDOhDhdM2O6ACfOigMwFt+OJUdpov9p0BIIXQSa1As0nbkV
s/X2JWIqGG37JdyV+9eBfQq6dRgneU+jCJT+uEyInteQnW4i3RpKTHMDVPivZW4m
1KCoStNlvKKQ5S+/rtk7Tid3cJRKTWAyRLQvqFp64hDuB+13sSkRLWKPtz0kPcyd
Ii2a9q7DPHNXjzR1KSVjT8V6Z1DT6L0+T6SKM93QA4t9l9z8Job8KC7Fj3jLeazv
qvbAJnCxQ9VNpB7ucoEuDwJocU107afh6irB3y0wJ3Q2do1BS4zmEuEVzbtO5+Y+
bbPuEatxon8F+XxECz5ipp6FEFcR2xOwKAasRYdRiBEi03NgCNL3oamVIT4mnzQC
WEwrPwj2H07W+haXBddPt7I+vOVnzFhjHdhLOogf+vPN8HQy1hzQiyzMp+d+7vZI
33zbhWCZ/ZhE23iUFVgyUKZ1SNiXc39dRPGUQAvDhWuE///O5LfXly5vUFDQCpdg
GC2r+Oot+/pSx170sjQqg5YWT86CK1dwHENo6w/XCh9BPGj8FDf6PqeP/nwpJpq8
mSedJc/9nyoa/axY3vZcAdvN2B8wSMw47/NQUb8/cgKsxo185c5UPEjy5mnGG/KL
x1Hj5O1JZc7kcLt9jo1Uf5ta1TO0C0LA0OuPtiWig+/h5WNMZn2KWdDzYzSETwZy
v/bhgyYaRFZRpDuGxIjD4VtyzEf6DDyXIWRkGO7Y0y8JkJY9SuLpEs0HidiKtEgb
ZYwX5M4H76stDlC5Xvur26sQA8OgkeK7GusINThr/TZpwBGWCrW6FMBOyYaf/5MD
elwj1TptHkLYOwa1RnPyMeyP7eSGNFGBwCg/qyOBgjapWSk5Sv2RYSnslydTNKL0
2b/eZwJIdo06DsJSJlhuWLqZ/CCx7qpkJ72GLvSIcAtqc7FWGrY33ZZ24wFGR2Gv
gdujwb5QdKvFnm1VcHl4WnlR44VDqgxT7kXEKbuKgDNwnJ0xdc+gKTeo6RfeVFZa
hM6/+KXyJsJ3k5+l0P0Pjs53hK0iuwLGb2t6Buyj16YnlSvpxjgFMyDQO9uHbhi4
ce3LMGrdCTrbst1R/poDVLMZhCLI5LyDhzH503BCM34/wQY0QHZ7Q8sxWT6Otot1
Ok4i8bpqGGY2vGbXhdFwT/sctED3961MUmiRgeRuxF6BvR0m/XijhfpfbA7c3GxZ
e0SGLyE2LXw9/ML2Zlfr1SNrJfQ62wDdxKFNryhtqy8AeheLoCxzjra7J1XELOhH
LPeqZJF++QdZBB22LFkF1MhGPJ6zL3UHShsWalxezTVP/otbYuGmQ+V5ibgNuisw
sW53iYgGgivMVLBU2nV94+Ac12WfCflVXm2H6Blk4pVZ7kLc9TeiJuB0Zog+UUY5
ncjPO4P0Bhnj1xbbcEd4erkFe7ACNopGKaMDLBlU1wOUCiEWGS1wcY5dy1q4LqJ4
9LpEJw99MAlh2Kp4jd7fi/Z22CyPgAXV3alnWOv1p0Cop54XWA+4n8ZWeV2cXeDY
hrg6wy282+ggvM9GBE31dytPCo84upwiJul3bgfnjXBHzIP0l2KK/S7ZhcJgRxN3
GHWZ33jtGPEX5Txko1blCcabaUsA8gMRsawIBg3J4LukWvZlzXrAOBPqY/SektOj
3I8TkSLEgAeWmpxaXFWntf+dHLms6LgmA4hQi5VgvldE3j1cpE4w3PfWP5GlZ5t7
TeDeAn8vREiRi63T+e5GJHNYfeKq9irsLpGAXMq0tGDVh54ARbe+6h/t6I7n59aJ
eIOVVtDZEp87mN2kNH/mJWrgESm8MBuevOjDsSgiw0h/hk7QMlB0qSL7q4J4MsPN
vbufDacfXyX+Zx+yfhc6kzR+zlfBNRtBdIn/R9bUJd8dlDMt2zlSkDzcH/6WVJ1y
pbaNG7Y707qcwaK4ncB5gp+YyeR2OVAwXWi8ME+vcotUJwzICd+PiTYHIfxwPWuD
SUYdBhK8tECetiOY8YtvYsBft+yuNDxfwo0cqCsjp8izssgEX73UIm+t/MVrDfyB
gpC0WSJoHIA7HL38Tz4hAIyf0Y+MYRhX386WORJAEvxe+YefvGvV62a2n1XwfjTj
m1blpXKFo6rtaZC9+AJn6g3RVgy9dbv4O/jlzhPKZAPPzLKaQqHWLJCaouWc+GKI
S6g+6FTaz7eHK/GO9eUabljjfNlZ1RmPAk0LXsBIYwwmYwpq+w0d+xLcB3SfRrtU
HC60h480MeNFeQLLaHLKFKluoC+GL6+gL70tzZt1oHd+/7POBk2QhN41s5J28nLl
nlOqvkEWB+Psb6p3M6mHkhWT9HthS3fx9t9bkbncKGSF1NgKZUZIKzH6rACmbVOG
zIVZAdlTwLldVNjQGZqN1lEbs7+hNhb2T3oL6XipOjqHsfIB/+cEU3spdhIfrZVi
A4LBEjN32EKWF1cUUv8doM+L7BzP20ow4er5n9z+PQGgTlsWwBnSE0RlTVDy9Dgj
a2lmoYRAZ64QpjIbbfJe/8a/cyExMgN9j1d2mFKSPujvhOifNTTWy3u4DyrGlsVf
51umjtCZYZEqKVbYFV5D2uUOUz2dhkZowrpGlr8XFc0j4lWYRAX/r3T2gJBNvKSb
sn4d7PWwBEt6z/szCR5uhxGNY7W5kY7hpcdUMkhqUBuAY0afuqGb6BC5FDZz9Q8Z
1z7xMDIBMQa6rYXKAdV8qxr4HkFkuGNbnPJfrgX4NGouEGYI4Ywhjdi4DHG2Te11
KracV5La48ge32OiOebJ/vWJc+p5cZp4k78VL4M8gJUOmUbCQ4MPjT8fJS+hLfki
VUIBCaLB3MFQDAT8NmdINZiAetoqOucW/yxg97GiuaQI4+gMU+FzM0AMJUagM1AP
MxQMU+uhwM+CzxCk9CzfC+NVmPXqipLDFYZkSKUX+bahkRu4nCIkpTC4xhMxs6os
wQJykWTm1Y54m7ED4zyLhAAFcydwPH23P4LdHvOuQkrQ7gfN1t/0yEqxNjX0Pnsf
125qdedOL1C9WZDWM4sdW6MAFPMtquun1debxKE7MgjPWkBR9U7cmlqlBOHNhwDy
Q0YJkXXfz+n265JMEDE5E3/aN0iwIiHmG60A3Wz7aEG6/TVw00/5Ib+0BIP6zhes
V0852CX4cQf4rmba1vZ4flfg0tv1zMx09797fom1/JJzGhispU6MkUpJVCgsuoy6
FPOJkWhVW10Sxte7I19VY8WswtlNY0+cXNz2vesP/DS75Rb66cNqYMBGCB5/fjGx
0ZO27fdQzI5QqidQhuboy7/Lw7NngjEb0czca+iH9lNe7IVm/a5Zi+XLG7S9BZOU
ZW4Kkd6soHtYWjtrwbw1HGNkb3OpLkCH1Mw2VyJXJUjmSrc2CQ0/cBGpaSm63XlR
8M7NOY270/SswZtNzGaok6iAJfMa4rV3ldpAUohIceyHBeOfvylsnq6Wmk2cEhxI
7WXEJ5ueraZ7lo7ld1PyN+xFVrM+74Sryqpg4UyPJT6cJ/yFzdYhD7J9w8Avd6We
RTqeYzeaOVvldyxj9kS3gT7J6xJt28pRxZI0hhMpvBJOWx9bih3LCsDZUzdNq/6S
NrZ9/cW+pro6sp0G+jErM6R3/246Yqk+Z9f78W8glcDrPlIA1sAxqtbeIk8c4yOT
p8qabmTcgpgXcQxSvSi+jiHnLRQ2HIuSur8Vrd1RtcsKcv1capR8s7BnPtKddZyP
orst5SYjG7lvSLvFkKvE9Ma5Wdhx85JnynYpyFEs0t/9SCHxsHbZbBAI5PT7HDE7
u1cbPh8mYtfYgaDGLjFp+9tUGae3X4tj8t0u2TNXcC2pZHV87ttH7vyXMHKMCqqY
Z4yJVnTTmqK+VEUbx1Ir3doj8L50JJC+8jn0qol2u8YngzObYLVulcTY/Acqwkw7
ViSHrTeCgWXhF5Z9IqybvnNTKTnrcKl5cFyocLVK6Xqb9OCI14cUdww8SYEtrLVB
9cASAUwuQAkW/HxOMgDcSldGevn3Ol0G2qC1ouVCiFVloDlxbKXUoA6AVyVsdy/9
LoTyNdUpV0pksWVy5WiecKo6QEoQDslwMPrtjtmSob/PYN0WTPc4pARPKh+SU8yu
Mu9rAxS+Cr408vxeiuyd5j6jzsJ3RyfgqEYYzMVfmKa2NpnxloE4sbJY1bZ6cp74
/GEYZaIxiGdKl/mk8SWkH/exAyyQqoG7JmqACMywn4ZkUqDsiOAx3T/fnJ8n3aOy
iWt3UxYLbCvOV9rVk9RENxm/zWpHdvTGpYzlTBK7Nfg9XqcB60YwFlLDvWIefHfg
4DtVQUFsCOJ7qZlwFbhhaRecLGAcEqb2KCgIhWmuV/G4Vb7+/Fy1b26idXBbSenU
KQhz2xs6AyF0rhWfwAbWwB+FnrW6NNJoBTaW3gnczLWZZj6UrRKRrHTEF7Py6Alw
9IF+DMrfsvhiT3bobjTXs4C4V+WHNAZCypCvBhUNtmwl7hcIzvnox6ZFFFtr2ign
Z8KqG2CPyNKMKODPbcjlSYM6gBsihT9DTkv793kJky3wYyC34lP4PbwrMBpOfx2s
k/JX3noIR5PUdYJtVaa0Iggf0o+2xJxxKddkKJ/VJZRzrvoUAvvw+UIi8Gp3LBck
pylNkLwDvXGbWUjYQNv1MekG1BtLqVypYhQ4L8FotYDmS5aBmJ59+BRu869iNLZW
mLHv8kQNnWtM7fjqunLBo62CBOns0qMAjXHk3OW+zSWpNmofRJZgDRCdEnMIHqY7
S/sKP32B9kByPaqzpR2vzYRvRe65oPcpKt7r0hiTMiUmNehb0FNPq2aZFuwV7x0+
cla5Pj/Ym9of58dGFay7w0ypgvE/t1ZVztCDmUszSZDAJbiyL5fBV+WRI1RBBJwS
Gx9g4mVo4LVyJONxgvHPEibiOR5ClcfnEe5k1KcNdRFTPTZ5R94HEEm5SRT69TYr
/e4BkPgjAnbX1NMJYIcGvKBf9kwO7d3/buUFeGv86UxK70RFOsUNvJcU/CW6/C1v
PGAblRVzIt0BhCmUAB3jr25UfT8cdq/+dHrvYQJl7MAbji6Al+wheumrpymHAlhB
VouWAA2M1ZOytRzfIzKiARR5hOKj3MAr8Wdx2FfHc6QzBUfUMPJ9hT4RfclL3ZYa
EPOIjnB+b/DMUDLNuBFBm1kHB2yYo/A3Rsh3QX1oaCeC0paEXmhzHgGT2uy7NzWG
43WDuQz9a9+8mniBOg71TmtatP1JaUlLA3kB/S7Fz24PFWosZdlBuJO+HisBAn89
7Foy9RINDVgLW1oTkhlK4V8qoHckxYKRXm0dkshWyBzlodZzu3XNTKxxDFZjVY62
MgplxprKpkXteDHMETEXjcJhlcLhp6e0yBaHmg7De2AwKRiZ1XG5iqxK/e81EyGb
tsAgo491DkGXciadJD264W7wR9Na5eeRyjbj//8j77+NaFkD9MF18wMRT0s8AHzd
O5NWFgEzVe41QgDj1r+VKMNwB56T2qY/1gJKeBC0mOmn9uK2MxfVa7hZT5RstDhw
YIDZi3pPXSRZltLfEbIIjcvjcV98NAiBuAXh5OLBnAdwwxOTVHJqf9dUPT1o3qAm
WltF0U/5VTMENlju85dkCzLB0QWYdrXRFlcGO05BqYK9hUy2KIXAoOXBIhJZN8G/
B0rBMchUyCuR0ShH5hw7MwZNamp/m9cAr3CN07DjE9nu9gUbUY0xOQ+3yE7HhgMG
7UI5ulSIj22fnh12jZ4cH7OJSpR5id1Ht4Nz/g7AD4qsWX/JHkdUmFbOb53OoVyS
WDaUXU5brjz6CN5nmdDxZHcTtA8Q4FlB0ECLSmjUwCpLcEVneNNxiZJXjB0AfVR5
Pme6P7M4s8xhwv6AOD5xkK97zuKU+tu/CHkS40HKXx29kU+jQXCsyg0v/5r5vllu
0PADkroCCbkmHNU7b+9kwp8Mg6kCJT+0MFmT7WqgphMLxHi7aARTuPgPrgnd+VfQ
zu/gKhfEOU3rhOKQgbdjfQsDycTFQweTeVAk3XJ30dpZxmxUno9Q/sb5HjcVCuID
3mwvsHz2Aatv5gThDjr3juBVcWOgNskTDzaWlsboQO2wo2dDStNdQSnpcCWVUSCj
XdsEY+YL8FvBQgRLscESiRRi+/qM5vidP1V2W7TGhhHKQv7Dj0JG7VntlE1CHwH1
9+NJeQfT9WlXm+G7huuJ+vtKXFgypC4zI+TI2mZk/SQfW+lOP5GjYI9HW3TfcJe+
5eQMY8PVNGlhXUZbfs+7uMKsnMrJ+bEI6M/iddCl/P9X3l5vOv6yXcaFKKzNYP8O
NqN6cXq/85M/AiIi6MoclmR9XaNnTPyqniULXTs8hYiYd84trOBAqhHxoiPrYB30
+tLsK4F/PtqYcAJyP/PRcF1YErtxlg14U9bTAdkKRARGyJTnh76xTFQAnKPU35k5
hiBTvXZBepEi1Q1SRbWiisz0vgnXqOlIqELclTA9rlHs34JfoCXduIXiEKRQ+fo5
fEKAtaCBr12KAMTFTe/HxzcCb35fvAIqY1+uwZ/u1dmqWECe9SslMQVJb+35WVzi
7hcRsoyEwyLMJ+M0Sa67aBCnHlP5N2nijVRt4FrxIY53Rh7FR/OWzCWzlnPR6bl9
RMsZPVWZqVW+BSZoFViLR7dCyLQOGe1bqqV7ni/O5J79nZAvfLJq9TbYkLozCne/
yqS1oYP+CmCazHPReVsB3daeuaW7oGh+gVIOSm/B8WOI6YZ0OV5oLXfuClv/T3wM
RCL+wZKxm6sWsOrtkbjf0PX4481t/6gbwPTdpnrCtLEez+zzeFHGCBHh3U7o+ylk
EsNpa/IoprBPZts5zrXCUCp/GJFOUEJkLcMJQCL2XmRyf0P1VPRoI0GEv6VMjXlW
5TCBGNZWkYp/paIaOLaggNGvTjQURNzlY6vyeoY9FdSL9rBdtEFScOfBT0q4j2/3
U4Vs4LJdZPHYn0iN3X5P7MlpHa9iMwfrtazclu7IZokcz3naDwrNroataZoJqzPa
quRM9CIAE9ZdE4IBuEAxt4m17zQoiK4jumSSZhRYqUxbJHrSlfmg9vPjMToLWEwP
YHakmiJIQrl6HGk6GW4phluo4FnaocrDVMZxhHiT9e2RftJY0OCQPnlgZbhq+ynC
Tj+WlZ8sH4782ttjx2X3pLAThxM1UVw6wW4GBIJjY1p9RxkAYJwuwQaGe36BnPwW
rsnsz+eopUYzV9VY4a6l9f6au/klQmKlSd2ntLYJmvR9U6ke008M3/6jI4fIhnNO
o2e90djNIw3KXwFOmDZ+mm36FQwhVSuHH4foHhvPrJDghyO9FB3IAdx5CT5k0Hri
bSUe9Zfx3B8q6IQIDo6TpsbQOl1XQuN7Kq9YU/IaVbyd5vs0HJ4eobul8C12owej
rk8a/LzHcDZ7tSuPK5ICbfrG3jhiYaGMLhGMt5lHSw1yf9VjMJ+eaW4QwRfRmCFH
nyHDcCKhJiRrz6h9W5TFe/wdnXFalLAD73a7xP68rogfMiEQXya8Lx8L2iH3PjZk
SyLTnJ74ddQkNnVZvoZpoGhtL4pPw48NpQZGQ+xJVUj9oIL2PFXBKtSd3UurQ7IW
RZDkgxrwVKL0c23jUWsMwQ03eim1xfWiz/SMI2q/7Bp3w3dV1DuQ4+e76xHNzoeU
0A6SbzVzVEd9z/VlbtL8Ju0BVnidlVsX6NXrjD6gqbXTxA8/SiuChgNWQuZ9DSEX
rh+iV8H/IIaFl7p7HsARCRFKePXeYZJCjhCYpaEFOkR+NA6odlQ4TF+zLAiRUnsN
C1uWCgA+QqwkAXGmb4HSSbYl4Ll1r1wTylq7ookqY4AYD4ZOt+SOjkAAQ6KeGcm+
WhS1C8rRgfIGcAfW3xVRYPPiSNmc3/HJH1o38UDtcbShiD0RgIeEoNcPKtMCCEPa
PbDk8CDhttKxjkLU9+on5Xplf0/oQ5Ut4Xd2sFlFGIb4gGZsJIqmdC2wLiUERhY7
6MTNM7R6IIINRgDfwJ/0jUxMxBKTV/9hErXLEsSERcp1jKXpmTG2pcM4MX7vEPza
pPUPIa2ydLC716my4Zfy7+rS85ZUWjVDb1F8tRw3LMNwLkFmhS7InZBdUSs1rdo3
Qtxba6N+z91XehyqJBqNp/Ifvg0J4V6+B5dJt/Q3MwBHVJwsSp9yv87AtBZIrAAr
42OXhKRZjFu1r0qiQt+vZWngwqYwuJvInea10ujxR+53z7FpZ31k489EOm3Mdcbw
MSh3LrExRjETJI5q9NwTq1izXzuVuncdFsAfMheCacwAS8+Qchlt0Se6ZgOOXFXp
uKdSQGFc92DIioy7m01XQ1m3D19EQOc4ha+2zlDMCicE7bfQuDLT7mwOvj4C4g7Y
LNut4OzJoBp+aXnAr7Nvm34ZMFwv9271B0U08EWisT8KEBWxr/bH3M1pfe9p9BGM
988a2fWFad1SmiblcczMvzt0TbWZmgUPkoP21x4dq5D/KIHDpw7BkS3cp7hjAu2y
S2shDBLnzRgk4ic+5j6zYM+7olpBb6hvNE7mQe2+HLGprbKaDZVDdGcaaUtSGw78
KLPHnDfYMyKjHA4cbNyRUjnLeE23oqPrAf5cZC6gbXeTqgia3GRj6PjsIeAxLMQy
E+0dCZ+SaIGEpOw1OXZayZnfVvalraYnksSAr6Z4p0hdyl4UuQ9Gc85qTAoignRT
CfyAJ7nRcwz/sTC3mar/mtMp3PzOW9QLFHaDpSL+zbH87ywz2pbHvQb1NHt75mM9
UObwobQznCg2cus9IIerO999gFQloh5XK5uNU249kIMVhriEgN3WVeF/BksrDPYd
CMzLLwxH+zAT0G5icRHS1yiGH3oFucbz6mlff7EzzdkX/78Gg89nms2qM1miQlua
MiZxffiV/aC7WeDSHezIeTxLBXr3xnn0v9oqtesyptMDcs+gVJOqx92/HtL0+VUc
7MYRDCzGV3NNvGRfRSMMpW4GfXgchVDUV8SU5dXHXi9Fv4uvHZ8YX4WGOwEfF9lt
2bko/epxNpfAGiSWUm14xP9Zocjyb+nl8lxOMGG6kaN7yd8cBOuTA+t5dUxgwLen
hZHjkFhy5R/X1NaePlPyJB6uRj2jS0oCoakTO/8JJTDnvazUNXSBtwWnOvxSgDU5
Ve38HG8zXHb8Iv1YrnyW6J7Q8B4bCChOuNO3KIvRcMZCf/CPuAw1fN7lGuHvAgG0
pz/ZHyShHvLHA8W0hSCmSfc78HqX7GVdbdhW+iNOSQ5XCdOx0eY50NyN0rB2woSW
dtU0NAaolLx8B2ud1ztXhJ/wS6FZ982Ry1+yuinejtbA3NAc6NCqDKW+XEuVzm8e
2UNnMnKVhQ9nBiTnqJjIO7MJdNvFXIUxu2XyRzcVdKdAQAbTbVwpt/IbXpdhYnTz
Dw2RUnQL4147D6edasUkaknAaY5wyRSELDHyj0oCylkfOwRx06U+sMKwU6GMdh9U
HAbY1JrHKkyZ7h/QZTNb0luhpr+43ygyTH1ay85bbQh5rD5iL9/t1CTc9LjQYCj3
E1g1+NtsJWqQJL9CWhAo5CF+jjAIRYvs9f6UUTpw+TOJecoem1Vviamiq/Ycj5FG
e4w7CV5tXOJHOLNQSsi6VcZmqZ7MHvZCDhmrJARhPkEdjO71DSTE6lG9rBFTQVVr
ewAq4UKXSm5qWsEYvy8wBoKTLQzJBVlZ7wNI9uiIxuPitRIHfnE3Czju2kQH35sA
OQBdFb6cbrm0QczHTnh55qMDbzeDgJJ8a1Fez86Tv2wY0CVPLeGgfxWnAG+H5mhD
0jduia70/BibfVZ0uFEe1i40Qj8K5wb0t7JgmDrikjGYvCWlpMA6vPuFs9bm99Bt
yVOzZ2mUYnJ2PJ+CbvW64QUwjB8DFNpBWE98mFlyt7AYB8hW3uMspwrKxNrQUTug
KtITpRy5bgsh546ZUEBejTWgdKk5xBIqDA9UCuRv/p+ABv9up+7kcnOQek1RNUaO
lccVYwbjesSG4sVRmPZWexsKRjemfYareOJ4hS66UO7V08nmV3QqdklAH07144r7
QfO2JJOsEoV7DibDXHlq85bAGfjeQOHLYng6n46ac1WE+QvlH1noKC4LMRWZAebp
UupPC5a1t1pOW+sD83HcV0tcDmbQ8n9y1UNMa7yvnFhko9AxG/WbxqY8tgWSC6qn
/hKbklNbN7CylemhMIYmZrCtX1LwZ0dcb4qLKF/pr2bR5VgEzY2SCG5Y/I4nWUbx
ceEcwznA7dVhUc0r7pIrn/hwQpOsxRKHte1++9YhuhI4fvbBTsZpG8EMqI7/xDLB
OQKqWLMczCmvonmpCDgxwzvUrXgYlV3ItkTDiVEXPFUltovmiZ0QZoiMd7xwCv/D
T7fdDP2K6a1jFrzkGEjrTcxBD5q3Z6iwBkNn+uDVb4D87WeuAlwO/dSar27e1uIO
/iM/M5Edb4yXmsJui3Jrdp4lO6LWdTQ9CMKdILe85Woddp7+LAm5cOKHahrUyayn
SLoraqRsK81AjOAcoFTOhw/p2J3lOsJGpCht5FLjZCVYrHoIvr55I6hvBgd05WNM
IPANUbSUfsGbgkarpGmgkVP2otXG1vNd4//CsAYL8iJY9zNH53TcAqgdhnLTbt2p
0egARg6Fmtryk+rg42kjJ9Bf6CvT2cdh+Rh7SHSGAu/f6ZSDpkxw3M127UnG9kAS
2TnDUqAmM4sY9aN5vOhmbztqR7HYyBJmNDndjGr8TcLxRCQ/y1iZfFdoNuc3gqna
ZSqL8ZT7livT32bSSLLW1zzWndYSFgDQ4L5RSPF/dsEKwKA5uvZguGtWR1OAifGQ
Kc+b/5tHfAOiHefadu5F+2hS/fA22+tSn+GvUA1StP1lGW/UBpIlr9hvPk13JsEq
O66OcXv8zX1RmBqcPO9bMDA/zyRfh+eGUHJFtMBUqhgsUZFWwXyc4L1qPAWKIEh1
/fywi0k60GZfExdtLlS7qEqI0ihWM0aM88EfPMh8/otsnGTw88Aw1K/EM0ekB+TQ
OFhNwLq/72+HfVBThssszRZf4ELqpTRCCD7WZKLP4Kbx8y9RUW2YXOUt2rR79bIx
72oMHkgN5uazY4DP5Wek2t3mvOWDAkAbxVfoRnFMtpRC21OIE/Ab1uq6CVk1rtcy
RUx7hDy5paHR8iaUfJ2HMlG3sqsSYAm2COG/1f2Am/wluw9p5Jifa5H2r5u2TQhF
ys31OJARAnM/uKrngWRq2X9Am8olvk6dxhmQeX/AQRtgpK7UNnIrRzxNTntlwwZQ
bn5OLRYdcygO1y5+8EN4D3n7pLyyuLlQaR4zbgnJabX9Qw1EWM2NuCRkhMCVYDy8
0wNm/URsiSEkTEKTmCyPnoQUsejYuc1PMcEb6s9I8C63lq+NXYUbfRX7VuBb+c4w
U3JS0KyhfkrsGcQcmenqVOW71nytdPHuKwzl5E3q3goyYGNdgbHXRwGlMcjfxtbH
FsI/CDqX1/Ln8kwD4MZ9gkk+WrFuFLrDSvuwgISqo+ooibtgu32dEEPtsCGXOn+F
VcFECwfIFRy6nAtsglwyEMqPSAxuCaHhjm8TeTA4R7lmLWc1CiYIwjJGnTzYpFdI
3/9TXYoT/sn7cgnoG0gYueBmcAEwIgFsgM3VEAlaB1UFMOtbxk/PF0m0k6GMAAa5
Z8e2FO74PCMhaqgt+rDtnW0BVV+H2TUWvZXOjYoIL2tA0PKLi/3vFHhs29SFuprT
8H6wgWyQjQIVvmPoWIEbNnUx3R41uxaHizsK32lQJbeQ0jAlXUOVuWwjF1miH9fL
0jb0IAG9KNr5skARESDlFnX2xhDPLMdHTXauB3gXlVnHOLORrYg6o4IaNvhe64IJ
T6HXEKbKJyskdhK7zrIv+LNnm3IKe4K8/DjPPjLN25Myy52Fjd95svSh30EZqWDy
VKjAMiQfTKp97MkpaTfafdJIMOL6qRKWE5rSJc8UjX38vBVIONAbYevoANKX4nbE
WkhmZTMjIk8Zuv6dY2YITzf5/JH/bs494E0rvU17rW3h8xRakovD6RBDsZWV2NdO
HXGiacK0d7QeK96hwcco/v3Dtq9HEUg7KaDkE4Tth+j/Y9jPTTfr+Fd75qTJJ0IK
egCkQUqlSDlL/Gw3DZrM6r05pyRFJPCcL8npX1qZBa9jhPHDvdkg+aJKzct6UuBS
6Qmrt0NwHlGZjIptZX5skaGaefRNxJJ1HiaYYdnCr6RMn/7ewljviWJL9eSYjNbY
dJONN0eMogB3u7JuFOT+tlM1rMWxfHnFG5plRU5a8Jl5KMsDItt3vXWVBDY34kVp
kCxDLG/ql0Dli+tqX/SrZ7XknVa+FlS4DV5kxRvszjWhjexZtvLPJ4F1OxWwgY1o
VQwM9jXnwi97k1MoZZ9NnO1mwXJWhXzx4NGC/QMMTOgKOmU1obvg8mOA9gaLUxrG
oXKsPogzG903F4Se96dG2mhof7ObVXuq2heRzlJbyCAuafGL8G3TJxDQRfvBe9gy
0yBrUOvlWqYWUea2R2ppgdBV8nPC1OfOWCFSUfO5mehZGSpJepaQOP2LhkzlMhFD
xSMkOw49f2eEC+siOmgi6xpN89uDW9D6Fihz8kxyJ073fLCn9ZpdxQH6QcTSnPMp
eHpt00ISL02mExdRtTbZpFYJHeLvcCjt/X6DKRDLRXB38SUXza/pBgxGOqqtpM+L
mJi+Devo4TEu1OutDLqm55YwJ5Mt6IvON2sQiA3I2cxjocNC9Sw8EXMRMuRrAzMW
j+u7n2PD4Wgtrkzl3AKbtnE3Ko8OSqcgj2crSqnyK42K69CWAZN67N1mT1wv48wY
dadDodrepa9FP1PVJR7QytdQsbQakk509B0lBZlHAWiT/LxGclP5h5XqS2P4GYgs
TAfsAJ7ulNNhFXUBw45sRl/IvcKYOWn76abeaf63VVmkYyYc4kNg8SsAIs4iYrZo
m1luYaKJc0r81Yc+iEdTW13J7u4UnhXMq+huBVtNIiPnlK0wgxJF6cbnEoN8qfT1
vOG9q7Ry8upyFG9+8DnsV7vfpE/RZZLCUAW1ULIkEfmZLnv1NHxt6ehx9cYqsUv0
jFtxvMu01q6s9ecl6no+n1tTItVlx+/MqjTAYAN1u1B1ExNC4g1G+BuX1ZHvU62G
/03sWG5zZ4/eIbLTPL46dBmkfb8EGRsIdBWKgwj3bszMF9Q80JBfCVEjGDdC7Mnj
vPWmGX0ZUWTqTp09DmofCoc1EIXnwHZ5xbsdRXEIHraXWwRRIE1nHvQ7UTnqD5xx
AH+Iz6Plz/0ApcV2WFTrSQKLHYIAnL1uyXO9ZtYrbC+vhWS7vuWUGncC4bWgX+J7
fF4fkBiNJFypfO1nZR3Oh1UXOuZlLdQmAa6qVGjuQ6q5utoQq84RboTIsFUwqb4n
W6tF5dyaclvg/9yjT9UdtLVj+EJd1sFAu+c7aw8+FLg1xXmDlt79dIE/PKo/IxlN
35aWXNAZXYbuQ0ZWN9RYWa+SH7Zajbz3vIE2zmTpHbFimc1g+sMdGN5B51RFQEPo
hgaloQkzSu3qRD5E3XPycNIh2bQrQuT8H8F5AkQmbZer8nPa/voSFIqo20+mfpG0
+cSpPwBDjPh6Ozo4/olRbb9hEiUJrOH81F4RhVn7G/a3GV6BBVQwbPpaFLcazF7q
qO5UUcFP18eOJMNP+3c6CfgHW+FgiJGAO/ohzPMF2Htfn/p1aOKpwV9PPEJWNogb
pQDwhnwRKo1eu7yCrg5qj13Ik8wsH+DIJTIRd3jd9uPnDxAG608VeKY09S+O/97S
4k92VlB1UCJMZVS35OF/sHnxSAwxvW3c06sXoNCWP5vIn9C7zCT43AiOgnz412Wp
m2DtahDpto7INO2vCfEc7ACjQ7v4ECZOVdssd/t7LoVfgZUi7/e9mXDCD2dQMawq
MT10sAs+WKIZoVdJCFk/eBrMVw0o7vFIjftLV/ajhDr/H9SfeOC95KF+yaUTCitW
BwH7WYvm7935eTA0oEJ9T5ea5VIqdyy3fkgP1TXf8N7ITL673u73LA1fMqwuPVyW
1ZA+O0PVVdsM4FQkSNEyK9dch/yi5jPpyqd3YT9mNEqAvba+WTHk1TF6rVcSBXyx
FL5qAsqOLsQG0No50hEypKZcvBjB/FZxl2YQAmKAW+51P5C02S5f20HRqHyyJTZx
W03sO7z12I8+G9DhApe00D/UCafzFLqcNFpPlO74tkcJrHhdM7MKCWOmxhzUfSjX
vRY38fQpVp4inhG9VZhZQBVtqp2RYI+9oZc5OmvotsIZ2jvKOPvT9OVzVSZwKhaH
hZrcPY6XJ6M7W5k4B7GSX2lmCnG1C74m4BiqfYPOGGu3Xx7SaFuFQx0xPnvKLc7X
Bn4g81N0rhDv5Eso4HdfJKYcOoNOxsNccfQHdX1wCfH4q39ToWdLf5xNtWI3Vffa
XjGEAWl4vA4+oKHFB7MJSAQ+50EcRSnS3FHp4DIYHvNGJnmNzZGM4zEYzs4InO4/
7c9H0Zr/SXrX0TYaHa+wQ8pydmkL+5lMlUfbgvEA5ksMy7HyhpckEqbfbYKE8yDV
pmmnzv1K5mp19SBwY/lddO8MZIVW07uLw8oea44VxQWOF9A34SuCRfnJPonhCCtn
Qn2muNIkfceBleR3C8cCWdnh+cMAII+F/9vUvwoL+rDx2ZLk9kuVj739pJCjoG9B
f51qCbn8DDZp2APWfNRt4Nr2MQwwuuCSny2T8To3SpR4cH7DpdXuGiQMh82zDsIJ
7Tjvgm1+MTDMYxET1+5Fa1ZBP88DyL5ld5DKpWLggesNm+LIrSO8iNhLFyxS0vol
+nS4IdMTB6nFM7Pgv0tQm32zW4F6G6A40IPmkFWq/Bj56yEYsaNLj9XK8Xroziy4
nzPdwU/A4aUwG1Sa9hrmEgNKSmIo+Vy+2Pjj75/o3I4pfW5JqMAGV8JvhP6YLYmD
YpQVOwmlzgTwGYElgp7VF2qfF5f1zhoMZK/0YD5Wo/M+1qvHJIVO/zB2Vmn4q6zU
9xSs5uqDkqqGzI2Sf4fDp7Xrf5euPifR/R51eVvOLoF7VNr6veT3B2qzt8K2Xxmc
uhRaLTrLYQg8TPKn3zrSgeF9O6AIF0jOH1i/mE3cYJktE2k+js1RfMGV2LfKMUN4
gWm/mpJDPpnNuDQkK/S2GB4M12kJexMIcsdXMOZ4dszZmyF6OQ6fwrbSoSLD2/ib
hAzwXdNVZ7IMdZ7PxkZIeO3kB/Rvg8plNZ89hnAFIX9iSo3jbaQd7l2WDzI5kfB6
HJueRojhMKElD36rrs06e+wF690F75xGL90LYcVBi5Wqmkq0LAfw0xB4N0phHb4B
Hm/hY2NYL/EdVh9ZQhx9Vn6ci2gHRV6PfqwJFCP4Ui6kAoFxTlnWtI4eAl26Bq25
pCsM+8192t/zlUWdgRcXRRfdn4DXQ9oqDUquHxjQ5T+onSF44JtH5sznf/iNQTYB
EPyJul97ONdp53gSnck0CryovwiqqpPS/Cp+LSWznnGlAFUZ8S3/kiVRYi9r6fOQ
OiUTTq9k1f03wQflFnYLK05CXzP00Y3xjMBGfAYNZhFLkUrjzGDeVGECnMyb1T3O
8mR9hOAT0aMQ+BIYZo+5xbIxBFkZdUVCLWqzpgNCcl8xbGEeHbglGOQ1X7CGrs/C
gkvu3a8AQt7GH0cRfto61NMZroC8YaGKjvoPehoc0Mp/Lh1rMq8hzpuoPBPmwhb+
0OWNR5xFpajvFchd0YaF4B5ItKN6hlYfQ1/RM8puMKVbs31CnkdRzfB9wP6U+Qlh
xk10LEnuk+ApQfpruqarZ9tM9Y8UsVcVBmfHFXcOOaCbPgFZDCfVj/BcWPJ81zcu
3Y7gV+Eb1648Zrs4PBhZMRxZ5C8gPjij6IBTx5F/oyqKYyClNQp6+d740F41JfSz
uEm7oQYzHoQ2ImopJBY622Na8jcQs2QfCdsMeGwb+a8b1Qb88SIe7tgwlEv9Bq1h
ZzSK8+iAk8FB976S2RWGxyLByfoshKprqYF9vnrjLnaoccyPkX42jyPy6BmlexCp
VqfQYWHTX+XecLlx9X47CKWrlHz9PwRvVstijkrpJ8Ha0G1Emd6oECnU/LCYXd8g
2dG9bn11X+XM6FaxJd+L8grY3oFca2kYjUbdaixS+Ur+0QFZq1NCE4DjdJAE+OZi
jclkpaIrEQOFNIDJXxEgkQento78nUhYEFj8zTmK+BuCYSYAI6PV2vUa0tdAjw93
8854GFhv0g7MFG0z4c7TbfQgEtSGxJKuAowhQYLI7+k4LX/e/zePPcbneZ5R1Fqv
/Polhtp7WfMaKpXlTZIRa+/soJc6EynP4JS+BWZBYM4/wd2Ryi0Iio7aHDwNvrbP
i72oyfs+2EQamKpu8KpNVAj7AuScz4j9akmxtL0WVOaYGeaj2ui+HkdveXqPEp/s
qZaxJN8BI8TEHJVxmdGAIsTsAbbR0CBFOk57+pW7At//f+EI4P/AHmDqez0l3XBr
GqETrOGdXtLvWx0EOExdCeOY2/id9WAj2p6UUwOqyVvO7o/jW9aNwvBtsymIq+o3
gIkDp1M0xZNwaebE39r1DtSyTso8HO27K9x8F/Lb7PtOQUdofx9yGj38b0Haiugw
pOazzZ+QhE1514WM6SKYlR2bzUVtrpIe/UC/LEqICWjR9RTLQ0K0a2I1Pcg5u5as
AsDnWm/M8j/4KMN9btMndH2GcbI+C3IpZm63Kb/sVHPU+xZsfgMYwz+LHEmRUoiY
zMsRkdJ0GeeAC/28ohAPI3JIk98pojim+SJKZ/8dgp3PmmXe6d8foH3pxdvEl82y
t8knpqlv02F6vO+27adIOsI3ZF5FAFx5ts//9APxl+8C54Uf0oBHTolvck9PJeDa
/7jk50LoumZg/shq0XolnxS7yELeewRgozdoSSschung+3apaUeDeLBoxCFuOasK
zPtouPc0aCX13YHBqDv7TaYqpyFtuS+IAUnclToULIfqLw/PgnG9uX0qQH4/dyf3
wzFboschwY0LdMpX0Zi4R1CNhvXfQprc8OEh4JiRbhayrJPR9Id2T3iOuSpNX2Wk
5rty97oIhOEyPcFvAQ/SlEM94/7LfeWV/zMVxn/ht3BAvc/E2LOHQPwH2sSFHZba
xFAo/pRflTV9fyj5smTr07vkvW8bZJsfXKbKBXpVlDQNGD2DCxqWj86tnGqQU3Xw
PxwJq6t44eNfWN7iaDMhW0ax6aucdQb6o30zgBhzVw7bPHytNHQma6tZb6JhxayH
Jv5tiZPYZi+PVWKsCPmk7uSpwaUKPSg8e5dM2BIj+HXK9+MceZXVkwgcnvhdicXR
6RO7N/E7QU/avmxhvpXM+u4OEwSIMxaLXCNM37qnt99WQVd2Jm4rV0pOMO97yQSE
PXRmJy3V2RnyeDznIWtLPYf/QfTfZNvy5O5A+/PTaO0hkeOevEu2s+EnkKFIM1Zl
Pu8JtFyFB7NuQVpJ0H90dewXw6WBmgPFRD/m8laHkNjq3+Nuas78jd3Mgb3r26GW
3KQH+qiFdzHbSzuqerCk9N9MsKtUiYwhDdbG8El3soXDbfmHxFv6T0zF6fJox861
zvT9vfxLFstgHZ1/VMaM5fnxHbKV34RAZ3JdS7HbHCphERZHyTolx+pZMj1YcdoF
9tZQWKtMgVM6LImoOTTcCb9pnHzGu77d66+vaDCkhOxhS9DYJnv0kIarWdrqtKFE
UPoEOBf1DfvVRy8UDmWc6Gvcdn0ZP9vcWKrUxNitBF5ioBPPlk0qIxSPejC8LTV6
sGNH6L1v6aeWTSM5lCxIRuuKr1m+gINQyBQ0XLc+brd0ewW4ahpuAHxd1gtMT0by
hsY7Uy15PnKxRZb1KdrowrjA0C3LdsBYxN2TjTYpD1zgVPYFP+ecZhPI/OwlnfcJ
Z7gGHYPfQRqNendiUsbLTk3tCvHSU1yuHa3lS0Z61Y7O9unWCkrgrPXgm0SbGS79
3KJJZeywp2BaUy23/GIrmMIGGRdNDPOEcQJg/SpBPQ+FnxsFUIiKQ9xAeY6nNqy7
6ZudiUfOBFJX11AN1HUTGMrMTl9n4WuLvNimba1jvqPuqL1bMHIo1mEo+x9GYtwK
7ROWLHQDQRydtEAi4W3whPn8isOs5M4vvWlk3Ddj/0WYUhJavaDUKTUOJNaZDf8N
PbivUKWeFR2CRQXxDygDXG2LzxjMyGlHZ7GGqN7gLn+7kYwgVfWk/L93XjDYv4pA
3WQR/4FTohaYMb14RSXt6aaO9uN4k+e/R2flKXPJLu9uGTB2hDxd3VibMwjHavFA
LvQkq7LmTZGdXjNYla6c38z0VESRh7oYR/KNoNNAYbnz3DgtzMzfQKhOxnQbNUHx
STZHY8RMIngL5HtAz3kWC/nUUBwz1eLrnoNiJK6qnR0H0kSXhZYRna1TSi63LIAb
vAQAzQblcdJ5UtzwwxPihHSd53HQAmPmsMDPyx1ZLluMmmiqRSArKS2YRlApCYpj
VcUYcYEEIExXd+cfLpHvdaF3SNCNpr11/O2lPvzpOhyGIFgVHOfi3sum59SatSOe
pzvLzFqqi0moSl0aQ7u1KktFRKko76bjBifAA2F5s8xaUubGCELjDITz4d+ud/gz
JRFjyh+RwSczQYEF4jZQ5eH0HQXPgTBW5AIFdDDaTMLHSXWjEdlOOIpke8rzy5WZ
Q7yoOBqfv9jhYGkipgrk4tIi95+b9X7e2Y6lxyiKhXWfW+SqTpFmTEUFpHQbdVkE
tQtNT1fZYJAiwuKevNfhztn0AXCJAmGyLSo1mqylbB0lAgQZNcLHqCerod59iyas
HB27Pn9HQywQeDWbCKmzuZVTru/poORpmuSEcN8M18nQ1DgVAsXAKvfgNeBU1/oy
orGfJ3Ft1iRIw0v/3JfD2O63+XbnS8RS5nRCVNhks9C4C8seBWDN1a64Ijxn6p6e
KIwpUmZiEi4nlpLkXt1YDiSmYq8AxS102+5Id0mtH1i4K7x/nuQPzgj34PCZkZAQ
l0JKiwR7b7PZDzwSi4t2Ny3bw8b7B+1aNbHZywmFL8+A6u0P3rIk+3qYVqLabEUo
+eaWgSQqNb2xn1nWmfNER/jlomu6SniLcFBHBS6pkNjL8fzKQjT0em60eS36HjLW
51Llc50I9Ww74IM1FuTktO1xdeBLPIu0PM+Qhx7x6f4k4x/LrfMQ867SSNzlTA4q
1OyU1redpWO8N3CFBYLZzqAiYwuF79Ru9hb80F8uOQ0CBetxGfubX/UIfETThATT
QUK1jY1hInO9LWPRytfI1vt3PbhC3TYfaIPAWovyOdzcIqPCAbDXbVl7Ie00WcuS
VxNwIkaUuB6VOAi7CSe7K66Fd1n3413H8Lj0fQ9NbH0hw7Ih9YP2mBLXm7ofiQk9
h77ejfYd0ZRAGhvSi9TpRowh2XZm4c/DeRSrHgU+7+ext3Ms/7lOODpVSG3DYCS+
oZ2mhDkpKkhshKuwi7/4chK7TvxBlg53SU6C6ABZ21WLH2/gABT4GCOXUzIKmBRE
OQls+BHChLBdGbx3lQFvqXpQAe2D6G5ShTqfjwR1S4FNiZzHgr4lVAKXswZOa/Z+
sMQKGdNzuw9YUPMtLLJl1bT2XI/6IAeJp1QfucDHhYKESAx9ZfJxE1JHulzlpTSJ
hTceajfe21mMxp6EPWHW6cfIOJwzJzcMwETsdEOBVACR/njPDdDw+KNNIWg6ExXl
2ob9Ylbd2DlzcwiQHi9EEF5RXUaYQ/stTjIgDx8hMZO4KYkSMVEo12GBQXDllasp
UyhWYmROFvN5OOY35A+3MiOPF44lXabXPEFaR4MJAw0JYfqCjBaNzZ7v/9xYWOPg
dUXJqO1rTrf8EsMWNZUwzLU8nakNXkgK7khr1gT/HLTK1IQnJbbeJHGp0R5ijki1
TbOOlMaRn2DDFYZhb9y02SSaycMalH78gSOoEInRafi2gVH3BV6qM/oCiW8mfza0
JyUs3EzvSVRXL2pMStbFTQEWOxvqCkiOvD9BII3YOciPbR1gaT1WZ3KRsNqYniVo
9Sea41JYqXLyKfRekPYbNXQqc6cGmhENKreaCdN8Qfpaw5bLgkRPukctXob4DnYx
xorMBH+Yz8orwNDrMZlaQSWxmrjm/JZD+w1WqolRASnyJjowdXhmGrxEHgRsNH3c
vzNd38UlXSocSTV5fiXO7taROjsDRJU9xY+rmeVziqf8mHpgAI2rlFzgtATvFNGc
KgLnALCDWo+wvF2x8PVJpZfX5a/kIengli8UixR39KKPnE6nFiC6U1htvHNM/Jw6
kMcyRWjQY5fXFwGaXsk0KQT3ZTx+OaX3HLHlr6l7NU/D86QUXFMSJkBeoZginmMr
fVadRnt3xjjIGkmLHpO/elTl778Dm0ONf0Biakg/yUnTgLuvEFGiK7T7/Ppv5WSW
2K4gCccHw3TB+WyIqFrIe1nwFX2063OtMjWusbyR233s7hCUfq7cFH0QfQLO6Cik
SRBbQiiKjlBLeFlQk4AN6WfF5lKWlmtZ2sGMQaeT3RTHTxwfj/gzKz09mF97Qifv
NAeVUOJyooztbBCqudd944zwfnHXg1JDkUsaJKRTokxSOl5h7yNSLT6EmnGCPZty
HLbWEh4Tx0E+XBhCFPZ5vwMjwqoGw21iyYkgj7Li3rSevfEVmtjpT14/K59VEBNF
7u3FajT1yldyB0abIu6oJdKq3ChEZZWAFLTGQqo5WG1FIsjQ0Y3XcQqP7jn6xXnl
dCnDVDQF8gafow38qrvgbguAhCH5TUDnqXMD6gENYGRfN4RXDbQq0p/k31upr6rB
QajkjXBa1QAASkIfVhDSd4738L7/xErX2SX5U6JUnV/THE35Jo0em6y10TLgj6Fh
0C5ROpyRMNBZW69zSG5CVa4DvXLJi9X7rv5pIUBmeMI+zV9Mq0SlsJCN+eboQikX
42S/yi51iRxrxk3UUZfTA/aQPck/os59nbqUBoaxUbpjbfMvPdXrSQ/kcUGGlXvt
75X3L6SSFXTdNEIEYmU5A3A7iqktjo4vywdgFgP0IHs95Sk/Er6/3ZFTAPGda8tb
nI7/7d+zW532vHsbJP3XEM8E/lcYOAlfe/qSlA0opXKw3vXGxZYaMoopOTqcvoMG
niklNOaXhqrj5M9Uhv9vSJuOeDeecC4S2+/vy6PlFt2OZFf+P1963mIZgm5rY1hA
CHfCnOMtva9N6wi889aSmsBRLRoQAUlj2CKXaiD5DYvgWvsDmG7Th/AldelMJmDk
kI7vX5OC0yb0ulMZoY2QSmo3Zrr+WLZvnfYH9XO2AXq6+EqYSmeKJpzOi3v6TPHc
WfxoSDrFwFnA+IJvSLvjl/DQeRcWm4RMKLVreLDpEWmydYt6NZDD0+ibldohHcHb
doLXb/ClgPNDUJRNaNrlDmysvGLBUmneVE/7zjUpjQFBlwx7YfAireDUfs67FQtz
ji57kRSVWhvQ9seUbQIlC0vs0eajO0RecrOXbfVAHKKjdXirkaP/53iijeYHhWNQ
GzM30jnKt8GaoMpMvxbrqhFq+C7iUrQGNlazqSST0eqySnsHj79dk6HoxqH94aSn
xLCNbdjhwIzl/1a8TaGLWTRpxGmCQ66WzYolHEsF31JTuXmvKuaasx/l0oVAQCUo
taIxbKwzHVLSumXkB1b/3Otbv5vgR2r5vyc44QP7vsz84e6RChLge9nU54g10wqe
GYnDh68N/9BVdzO86hQDSV+bI4CVfbLaG5kNxF7O/zEa3nunauw5pw864jXEStwz
HthkcZ3NmpOQydg4hOTSOsQxYXt6mGRCwB4D10KvjNyXOcqpBlxaOVXChR7lCi9i
mGwM0Ck9aiVzqbX3M/YmKFTr/ZtBvHwVQC89fsVVtwU+I+kQsZb+m+nyP2c/vRos
ThxK9gGaO7BqdJTNXM7AKl53wSvNoLiPPTO8EjjlLTrVIqUW9lajvq0Pvfe45NQs
rletDyTjx2Gl5cyObzpRetTbWdUhoUo8fMBkjc3O38ezw3XTkxg9SrGmF7lkuASb
VBRYC4jzH0QkdwW1DLLXYPQvFJ83QhYoaGodCwyX3wePjS+yzLv6GuphkdscrwSp
IF+VcYkdB9Xh0tmSrbiiNs37XPaIJREbM92aeA0eh1dfcPLp4GUzLq+JpkweYghf
x8nk9+vzKk66m5TN7bkxBSwrCHDcjzpRP1H7POUzt3mSceQHOAIUZVL0ejQ5FDXF
KQgqp6B3+/aZYlEiNbr6cunts8X5fLuImiSvGxiRg+8/+OwDQnAssdieOC0CIkuH
YDkXIHpyngqdFa/PFhHTaqKHZYX+wgkBG5EzRuiUCqu3Jm91nrc+bjvFxdMTWMdt
2ORFmTztcCpTsxzF8AlDot4Mt+jvAIZ3nt+5f3GGBicoGlV164kexcCF0qNanHHU
3XLNEUeK51LLY7oh5i1ovuGeammpv9yqLhxxmPtLWKguJ+Zkgr1GPqeP2gF/h4iR
H9TSyrb+WKYRPBJiwpClvQKdt2fj8EVYCngPcwBGEo81KC45KHi4lCItN9eQB22l
xFOk4iPHk2tO+U5GnA//5skyftjZAXdhR+H9j4dqx7sI2BTTQkIOo3P/RXKnvZqU
h9jrc+LZhWE0w2R6D6gVouLKL/QxeZpOx4841vAPwrK1aIQokgR+XaN62D3FeCBO
0JP+oFQS2dfaTrmik+p6s7Mtz0Isf5rndL/2Dsk/OK90g8imlCoXWwg+Er0tkT/3
ujwT9bULMkimwjaHFLFJGGwblpL9sO1Bf1LNrLFnzoLAPWzShgyvge/cw9YOu2h0
h2TbpsgwrFoZNNZbnphIs7FgODJ6HT6yOPi66jL1F7o9HT0EQNBWWcuux8vU32nD
Ll7ZF63O1+ywDhEpjVPrNebc/57HATB6/GR/RMY3rxegMqPXuR+dqaL/lWCBHWz2
Kl1ECz4uLepawvJr9xU5eT3Wgwvwof2Kjdv9IKOm9YoE5YpARg/GxpY5JYeuQAAV
6G3vBFnZC7x+EBKYSv0Q4UQbGidjDypsawP+1hTQ75jnlXyat/A89ynbrjJ2gbKp
/PotkgGkJN5sijX8t06p0vz6SiOtV5YwPwNq1ot0Tp986naBgxCvLe9CodfJCdGJ
NAPZni8KGd5cbQy6Gdapeqww3xyTpvp7JC+cRZzRT+sNx34s6KpjEwz7OSmh/y43
Am4WOlznCppn5ji5QXkbZClu6j1TnZYTfzMmwXyNTc3HuCJEmYNRyOfS1EyooO6x
aiJe9wmZ9THrfpgkVpuAHSpHMWDPnvUKvQGn/9wfTiRKa8N66lG3RfQokylbhL/F
VO6kadgmPjfq9gae+u8qX4gL6weH0zr/RcJ7sBsg60U0rCiQPI5pa+oxPBqejw6h
srAGmM8Lt7CbBOOLto8w7/mEYi1jNCI+pa8Zn6hVgkvqgnknaWz8q5dTxte5PfvI
OVjGlxqyz3RD2kKUZFKkYnvD6nxdu+9Z6viYF7Lv7Oxy3UiMKKY3j+wnyxAg5Qk6
o/VDDs64cO/kOW/KglA06LSYBmKr3nDReUofkv72sq0Iveb2+hTEmhp0pEiC94y6
YuPurR7rBaR1ZZtgXd6m/KvsKV+Hr8v0UJcusw7Sdyix7CYdwd8g6y+GlP5RvCMZ
ELWcGFsG8tydwxZQuSLq2yJ7BLGh7g2j4mf9M9DA0l8BgZZba5gcQWNOfR/wZg6K
YK1qt6uwQkyhY3uG0vZ8wDpuMPt5qIY43rvGpeTcS5JMUvDiCGFAITUA9UkN8UtD
WMhu/nJRufSyzX7QKoOUAavStA0cqrOOnvQ+ZRKZ9PMTaLK3k/23zThKJgeW3r5x
2SanrBCGmsqEP9HfyLQ/zyviqtHqGl0pDq5T1n6ISrqVQz8i8U39UJcHNvq/fKcM
mzynE3359VI/Rf3bKpSnxJNVdKhlNjX74rRLJ2bUw2rG9LHEFBJhZFnFzurj9Ypj
WlQS3VqkQrvHPNniSaZnC+IzC2W65e9ikip2TAtgm9M66tNzOLK7y1+GtUCVx7qP
415oy9kKQKNVKwwqfdWL67cbynfhPdjI+qSJHpr1wPmVVba92Od+XihQdzNLBzsT
opCsD3doweV2aSOe6cAZDjY5vI/3XKkVeNdzIO6p958qK09PfA8gKwc2yoJDuT1L
UUwNNoyX8vZX4Ltmr5xFukp/E1zL3/PjeUWThktFaOmmWY9Bhu5qBR0z7/eDnpVV
78mCNBy4iB3USLm+XbJtMSwGrpAgCxgWIEoDUpMbGHZzECDdGB0LCvFJG/KJy00U
v+I3k8ZMAlsyj7eq03HUopwy1Bugc+C2j+HXJVxeCaQGr83bxSP3vzTiq6UH+/9h
RSmQwBF36SSaq4uHNDmcnWlak6+2gP7Ma+/K4iAJfEcn9Pw3G4cueHDigKuNSBaD
7685Ee5KmzoDrUzDQlRJ6/opEyaQYFRc6YH2MBUuHeyquc6XIvnv+QyAWbBSf4Ek
Choe9SNu23cTuwhaPD30QZzEnCAf4vYYPPlXCSkdFHUnK/hu3RIE3+aWXVlbkYH4
/gLbf68DVH2B2gbOhfxPQ0YVROvMq88GaRz7GVSocf8PBxW3TkMvvj6d3kmlXQQ3
TddTcs+7EQFgHNEfP3K4LbyVtIFR3HSd3rmrMw/UrvQkvAZk/C8n2rmZg6wKmfdp
qX/R6NBwtzR8p+lEixPdGjioAPfHZiASSYi/RJlg1z2iOWh4KqFjRzQAU30DRMZV
omxfTmbHcv/LJkUjRimVbJe2DpzkQE87753tZ0vOrgG6bonGJ4WYJdMWyP8DPsGV
JHuV4LK7t4KKFiJjCVccLhlkAzILIyVzU0lrDv3uB3NPF2E2VqQcq+8JS19+pvSV
rncIO4ls3jFVCHO7YPOjevkfMXECOGJhwKnGja+qrBfODERI5dALRJ8R1dlAqbwk
LTcW0BLv7US27mkxd3j7NqJsEI0WV+AWR7ESrQuCBkL7S6ES5y+U6zCOy/asVuhL
Oy6icAFf3uiA4Kh707lkE9uK2tKssMqpX2lhPlYAdhupd8N79bD2tPv1lTVGmJTX
kqobHf6DXpz1S3hhO4M1jwYVy6YoVF0vvWXfWEvZ+/20ZTPESlgP2kYe/Kvmhdwb
2ApW9CTOuI+IktS5c44IBgymrkeP0N4sYs4Wt2oEq7Lw6Fvb+ie5Amv9PEHwAV9s
4P+SEbiUmx6SaGCrPB6jC0iDGWfMbdTvB0tzpHCWqjUJq2yNhzFOMSh3BNSYq/V1
s+SRwJ2Vd7C1UW9QojHGN6Qfa6VWMy6EuQ7zo82+esg/TRtJz3cPCUKID5wnccuQ
ogG6hOndgdOpwn6OWPaZ/bZYBcxD9Wsw2DPWH27xy9/IxHSvQRhGQJm97rKn7LpX
8p86RE0ELrqlloPzu0LVH/GlyEkecqxoLptYGQZbk2m68JNm757uJkt//p0CR8sG
8EqTFvT/mJTILCtm46rrSmowfrMB7pvpOBqT2tYW7h/f+Ijkwe9OkVXn8EBZYjNk
p1Pd7okOngEfyHDsYLyLedCQQcrwJs02V+hphJUVIyHHmnWs1qcQBxyfdf6DyRsN
Vub+72lxEokqPebwjvNSjGTt5NKeyZHMg4rFm0u+kdJUEUZ9x84bYOE3y9RVhP1L
dGYqru/API+frOaW06VK/CsJUDsOSfri4czBx7gjKLapP+vWbct6LQylyIiuwVWn
/r8r4XHtGwlSgyfb8mdAXY4o66/U10mm4d8ku424xziPNDYZLLmz7P38mwylu4ei
s8ZphBuxK9aCwa0WItbEhm2gBv4JX+YkVMSwdfN+zfjx+7Jpd+je7IjoFVf+Xbcz
Loc3MlNZn4zrcTjHb89w+A9b0R69PFsBoGcFxU9k7pSLDLEzWMnNGxg9aGtGOvtw
4aFxD0FTkNzOPJF1VlfN4NpST7AKk9kREG+eRUtG2qhNzH4O9AkLNuw+gLB70trt
K4npmD76UtYZGVugm0r6OnLImDKmtYLJrDM9IDAt+FJLvr03neKprDODXuM0v0P2
IuThU4pCb+dPTET/Y9AH9DKeP8gBhKDdBX8B3mkScMhZN9cg9zr32wYLXjjoJC2T
WelyXnGf/2eARA11LdEjQeq18fLbsH8jyFAsLZxDmo2XSmpWN8u4N1AyADhC39kl
NDoo1hrLaVHzic+kIOhH5jGoSMP6jEFS96HlKj//fsuY2uHsXMabjtOGH7S4Rkmr
fxSJ9qIm5EMF46ZME2afl+39IMpdXT5ZurH1XGHqyhjygs0ZZCMS10suymX44/uc
N1q/+LxNwm/4YhysJsgt89YPpwchVepRw8UpE7yTRyo/9fGZma40UHXUlAaHx4a5
ZKa9R1lSJM2gpSu2r03NhB/M+ztX5x6EAUzhloP1qN8NdNCI8witqiGTrG9PBtiq
sBc2LOSAAAWuR+8lK9aYAinWoRw5bvi53RSVjlp3aQiXhOI9S3BI+890/8gEQg4y
667KL8Nbk4s33DrlrgOjODpQXQWbyjohfQcH+Ltv7AAZS5Bz9Jfw7vW02kQtAxfZ
ll7il/K+350YPwvJfCtr4El4qAs6HtTCKRMltR2s5I+0Dwc/Y3Ap/UnzmZLwTDcd
eAMSFjTmxw1FgrxXGyi7IRIhmsda+jqquYdS+NWgaU5ww3MBM1Gc+CPZzZJs5o0H
sQK4e22QKKtJ/vBOxvKAEusqSP4H5K9tyrTzJfQfGhjzAiSg4LJPIAQkbPMPqR2C
26OJ5cb+Boh8pQGq1OrTbE1l/Nr+3+7/RnIaOB+37TWti+nQov76QRAu3L4wAd3b
JBdm5aOHug4dabwOXzmK4d9XAMXBAOr0Nttwl8htEIZmQUAPjWG6wGIW0lxue/j7
gl99RxN4TQX/Y/D3cDEXmFB6iX4WM+bS63tcFnAGgcIvEvOiVboN9lXS/1/myMsw
JOrlY5ffa42RrSsju88G1EJ2b69L2z4mWdIQ9inJgpGvN/WRE6HY1F7BYRh0XtmM
hXDj3LYOEtq4OvQZnBOwcS90eABDgwfgWpBY/gd4D+o+0SfTxm+kz3jzmQ08xDCr
wLPm2K1mn3Y44Ug4D6ZW7mnzJqOTT0RQ8AUn3W0YDZanv6grvTinBawysRiLTYVe
0mVwPUFqwpibD1T/st0bgMAsL9aALxocN1wuVshP0SfQbQFL88bZhh0LI4cqXxoZ
wk4phjSLWHM5p/YxztpYWrtSDiUI3yQ9MB4J5OSbkFlXccB/RPyZcesc4MYfn+sO
IWBHXQrfdM4rhyneEJTzaxaIqoqqfxEfEuMDVYkUPN7ZS0mPoN4olbIs4VUyhicX
a3Dfgyke8zz+m9abKbBrAgjmRyssuiyKhw/EJdkG1WrYiEZGPIWKZipsmnTY4CAn
dJCaAxeIcK4YOf/4ixYxzO3aTRwTn5gkLcfI0A9V2F9ckxhr66wzkOmodtajknuz
is2LyFUI+JquIWw3KL+xDYiCiQ2v0vf3oGG6HDgsZE7l4fSPt9cUZmc3KtXNPxlH
ajWzarBS7k8dxNy+j+1mgpvkzGtj7QY9PuAu8Chm91+f1Wc74+AC5AUQOxk5ilQq
91nlglvQ/o1m9PUoayqIR5HujEiyeWRQ61mrmPZgJ78Dk8jYcextC/NZw/CC1AhH
tyWcuEPpHSduQJqlRDJEHY7IKko/8k060TGhso9xCHGa3L9qQi359rE2p6MhGw2R
X72dMA1FiB374d6LOEHInI0jhowiQ09RGdjagLvtLwG2oWQXuW4beIQxMUL4cBZy
xwhxHCk/Bfak8kNcSnq54no7P3uiX1WYFCRO/yK3jVTVySshCcu4moqiIObf/+Ue
47xXEmhc8VMCDMgrX53aMSHu+zub+klWJt81MGzcL+n+MR/YIuOaRjpEDMnfH24T
uDYvxVWnC76lUXmxiVqzaMOcG2uVYvQZ0Ywd42wLMtEwiOZ14tHPAv5OHNKo6v3q
LOWOx6uZ0uD+L42waV2AM8Qu2yx/A5XcMaZKm5ARKK9NF6MvRXtMcZya4dE+T+f6
48jqp77U/JvvQJAxW8jpATZgzdxlPYWRx+b595BuVMzXHlV/bOa0nXWmLf299CTB
r7O2isXV7Wo2iLwF6XeJ/GjnH6DT3h4Yle1hQCPp0ijaIknIgo22vrC0yncLvQHI
D3F8XfRGGgTWdua/EI8oGJ7IzA7epCL7DiY/m1BHY0ri8pPMDlocRJDX0t+AlD2L
RWKV4vPlIji87GC3/m+dniWgxZariOIqVOsXNv6qHTTtSRbCtgHjNY/sDOOshK5q
GWJ64fZz4snQ+TzHWq7h9TicO/sQRCHon8rxAleqUQC4EMZXUT2cUlYtEltbtBiQ
NBnwgNhJvt0AJqOVfpPp17DWcoxJ1tOnWmARmKqnaRLZPRp09e2PLHYA57NGPlmi
aW/NnnwrGFqHk9h6vp4q0GAxB/tky32bgXflYzkqUFq2B8YuPTDl9zNZyJ6GlBEp
O51zc2GUBVTss9bPM0rBXwCxF5hDGNQgGBTN4OrRmB5+Ma2aHZbFfh8tzjAGHB0/
WWLxmdEMZCq8qhdu0GsSukUnwzcvooe1hjraACVctlg1ji4KBFyJCxDNUEG7/74s
SmbFnGLylOwo46rN/CM5a/WYEI0T08U//z14sQk5KpSTXZq9qkqTHuQS2BzdC9zq
SXzYfDeWUu5szPpu082wd6a2wJ7nchkFy/Y5rzhUNulSc9KHjj1rsRNm+dSvRvw8
oBMjhY5w+onicR1d0DZy2H76rfqQ8NBGItVY2QpOBtOfKFoobga2JxXWlyHApyCr
R1qrq3GhWjGbR8bIiYzkQVHo15xM3RnEvUP2yzdiy0/4cklIzJHIYeZD1DmOPvYl
eZitaRePEL0gfvTurDDV3rmULZ+uL/FxWB0AByiqyAVftdhekAMAjosDXkplIld3
6VWrkSy3aLmw+AA+edgw5/7qcfH0jMLpw6JTbcX8LYISKFOAMzIdHWT/9IZs3RcJ
UF5t/C1rd0oy5o8EkvgX1R4RE4SjXZKCWg5qEbToGoMA9uKq7xzaW4CojojnxMlK
HfC+5WNcFAEK+G3RsDzeU+2D+E0cvIyR4zBzceo+itSKZSBWkgPKwC0/kIm789o/
DPjtaQcVrdOhIgeJNV0YPNMLQGD8/OnUAUp+DGNlBdpMOs1lnxln/OllNmMzEIev
tWp+TWhA+cLhzW9qdizMuqAqHLaC6QXJP5k81KTUj5QfJQ8d1CyS6qqg3AVV4dUy
1OO+s7Ve2JCXl/EjPNOtJW/nFmWfe1MPA9vJsV1Yb/dL2BLIbxZDEIjtjEFPAYHp
vPgRoiYMVcUyxsHDWT35TYu0XM951eCi32OyRXkJDTgbS+PBz59x+3dW/c4Bs1bD
lq/1W67fDKORI1f2V9PKepLOuPriviMKoXNiz1UlGPazZgqjNrioJ8w8QhIAhm0c
+KTYlC+ollP1KyNhRSxHXREtC6+SgWAckizZLhReH/2N1eFGZZL1z3M8fzAuLa0Z
JIOf/PNLnmQarwlfJdJNj/XbWf7qTVH+HykpeRWrvmIqEB0Xa8oxsJsYc9VjGle0
kcOGqqPK45UzubxkwKyTsw+iGMJAwfo7twwVS05trMIBTtxNR7l9sDESni/hMyWW
91q/e/RHDe4+6n4hx+GkUnU6lZCpw048bYtxb60w2QDxv8tBDb4nJc/shNVt1tlV
0iJDYFDko6m4I+jCUzB7BXQX07rZy4rfBGyWCcNtF5mjGPYfxeQ9C9lOyEoNtC8j
2AZFMPnTr1dDAJFXy6jlZsgyXAJWNYbiYjzHi+uDwQtFFSGeBEILaqGPKHced4rN
6lFsvhez1LsC7fxNhv5JQ5hNm2087VPGTtuGkWlZpmbofGL4nrDxnswr3eTx/Ljk
FXpVIz+5DTtO6R3/+j6c4xuTf6LJod0sDFRsJR/CgMekdiUwu/kdgioVmnbNKLpF
RoBz+zhfbjB6woQpKYIWz4IutoNmkHXC1x7Uo9rO8jwfjBnSz9xPw53pVBO8pz7p
XGKYd6I5qdEPWT4cY8t8atFCoc9jKRAcnA83Aa3jn39cafh4bJwF8YByxHGwgGzC
68C5QFtU9MVynaM78B1q+lV5xfKgxHm8gN3EkLFiT67418cQBck8Z44rn9I/MtvD
MVxnN1SV9ozSByBqhdzyFQ32xwYVT21XrGg4oC9LdQrIV5AqDr3lvmKahIk7Hxrm
cVN5Z24lu9BCDcDEJGTjumalHzvDZ+Sg/UkstvClmxUL5pt08rgxF1aL8D8JHLqJ
tofvpSM7adt3r+HKJXHaXBrnkxk1CSVUfKT9xcP0wduyyN5f3tDqL/MfJ9+SFmjf
0aUwHpgdScKYHUGtvGDBxUQbCvwqDc2Lv6KiYjOR8EvHnS/kzNMn3IYSvMTli6VK
SXZoan861yrhdEisPL7a5D9LHxto3OPw5UHuv57YhVAXcsQxlKvjK+UyZ/gA+jPi
G2rjF5zi2ibc5QPYl7Lq5UBfZnCOfpnC6bq/AwDFTPnRPxeCQ5CQAZboq9uIVTDf
/ydIwoNYtzSOX6ZRt57ljHwXUTxHqyWxzCPlYuSZLhL8UXxrXqr7od72Gsu2cn1U
xPuMGJ6/vOGxCv/JhUUrtFjcbX75AAafjkpqyPIuDE7+Bb8msQprrDqJ4mpsSwBq
mRKouh+gs8sKMoUNzP6VNELrmvL9N775a3NepByo+JL+tVpCZJcSegULkoijv//3
lO/wbDA2uq5gWkqPMaPIc10kx0DGn/frEx1l4Qcrn48HSnKdTB4hszYegwPCl0g2
9Q670L34FYbdnbDR0L470ccej5WBtVoyFbQgHEPMk+DttBTgBIQT7jRlgr2C23Yi
Phqo4Jitz+m5XLYGdc2KanEl2iwy8CWv6wk4ff5f8acdKX61UJEDpGkAAbIthAlG
qgTnkCli3t7+hs19Q2UYGrVQXaoTyCOiLns+EQ4rVcX7UU+FsyVmIYFZ0/przcT4
eI8oVVZkpO7z+zGoq/2/FoD/OO9CTYwsPFz8JarX/XuFaI90ErO/KLj0SydNlHYo
8KaupKlY9gTBAPDPtJdFj40Ulsoj1tIV0kYSjApJpJeulwiJ0/4haJ3Gv9XerZif
AbX13BQ7jGEYZ7WROd5cKM5RQ4jMRgRhV48mCTsvVq/N3M5He0pCU94xX2RUs8ZO
jFSkLfXHINQZl3v2O0WqudWQrzyk2XlPuSM+PsWaEverBSJSNF8/HTdBTdS+ynxK
LssIXgFAmgm4bKgrN4HTiyPM1UNxyxI1tYB4zYcX+ib3whT+/PKuoifw07VV9bh4
rXRE9D+G5+FFwi5V7x0g1JQepYaGpyfmB9Q/4W3NbDfoW0Dmzt8k97YZJaDXBkus
tAu3jRvIXBNpTubt7NXMhXm3JNoOV8+qq2TwjvZMGXX3/9ke9NAJnD0k/1tnqKzH
O+vONUIqVzl14r3mneUJgUkCdO9kj/L41wOIobFnLMpOmwn6mNrXPV77duwKboAl
R9vmApWSTtO18nGInwW0jH832wl0PC4ninmmXFB7FNmh68y/R1qZpk7fXVrjnFTX
S8D4l7dz+ObN+57WZ6mtQjj9fr2H/XFed6GpOAsbSbQci6lWKG/DbJPoISek4ftY
tVrlNlyvlV9+WXJcXx+rjO4W/W1jfM5wW2Zjzz8FHDzjMddslW4PzFo/0ffPPdVz
RYNNSGINafartMhuZJY7XSKOLT9dURvQldvBjKEXApaK1M9z4uv/fm0QsBs79g5B
ZFkA99bw+JFUxiIyk8Vhlr9k2S5YTU2mmUIgfYQnal0v4//XkccL9Z8wzpt29Ea9
eG4eAtNgnyUodhBnxo1QPsYFP+NKno5wD2iWZsbfaMpvfFvtUhngt9LvHI+akKEj
3D9KGKS+s/YP1En1WT17yl/Cif6X4YUmICIlzBVOy6Gmxljy/UL/0vaPQjpzmW68
J9Pxq6qizPwXDnfxPyNjd3Wuz4ZGUV3w0vmPvfBJ5COvl5bTSJyqsjW5ciWIir/z
87xeYoG0cv83/KO2T2zR4J5C50bVXBOPhzWCvFCsuEgTIVAiYZ4RdDVoKJT41JZm
z9m9EqEe0t443LZlLwtt3II4Jjg7+2RJam2eHfJBkacHC8YgaR1dyy6nlXfBmmDd
DoCEX6dCTELVsqizoZ/HSMRJq8sin4yZQcu6NpeoJOX0Fx4Ts/s24dOc8spoyjZb
92Q9HlgoptRgLHLbUhdEHQtmdwbjzmU/0uNysx46bKfo9HzOHTKB4GwiA/552idF
8Q+NMIKaU4B/1e0ocGPSOsW+CHduAH8JVIm4oYNr3zh3jErQxnJyTAcXCr/1L5DM
0GQzfuHeZ966HlZ/p2odUMxEv/uGiWSxN0KsqugnJbD3ezuobCFxDSc2S4sWNwk6
5OrhG0oeKVD/rOXQ7/6Gx7elN9oRjTf7BE2xBWXetd+VehOPNm2mAg4pxV0umv8Z
epvPqTJBkL+VA1eLx8QLnteo9tN1itrRmmS31C+JQyZm/a4MwOAt6i1r5RvGvA1i
/B0f0ei2mhEpZ0vddcLpUihICQNy3P7l84rhLU2WmC+ItAYAJnUWkjf/mmifK9f1
e+gTcU2t7tJo43cBDqdpspupCZw3jGJJSQqT+IOiiC+RnUioHRPDx4aJrF+SDcHI
iji94tgqRp968Hrkrpt5vNTqkJEp8vFyC7jh9LJq7kG0baFLd4WEAYwwugrcBiJ+
4efLRDDzFzK6dRlkLsp9XVnCAkGifaFyjGb59/ALOZtx3/FUQCJEalc0JdWA0yn+
x8+MSsUM00tTzMn3HX/n/cXnv80FDok0+q54IwqEteo0j46tgzngrtR36AdumzdZ
gtHKHZcTz5Y/xQzsyUmnhFMrZzRQynJNlZ+kg0yOgcDfXn8IVOKqOC3s1Vf3qrXh
tAp5sfdn3nL19yjk8+VxZuFORUvPRsg8jaEDaSzGlDZCkMFrIr8P+Wbe7Ur6NjXF
3OCTlHr1T8kmOxcl1/EVczPoDW2TkrWgUvOTebUWMeE8GtEM0zgn2krIfAxJG1Vj
tsFiTTKdkQTvy1SwE+5SKL8yciRZeWA5CQx8cQvyaGx5IAWoeFaNRBHMeGAUK8y8
aTicZFHjLY2C+ntoHo8BXugzNhU+HmfFYFF1PiiOICtGzf5mCTM69bJehwlBrKwm
t7PIbSrFLeDS/HC1zfK18LDM21YM4JiaGGoIv5y3s2uPOw/ruiLpnDaF3dOR2Ayv
YHCAMorrtSAXcMq1pWkAZ5ZW82g9AjfRYEaA+XSgUGM+zkgCrWuFE8IPL1u8nwOO
NYVU0W5RUi8xMyQ7HBLv2EWKhOHfU9bQ6zWAUOrHsG1XCBvRJlha9IKTLKpL5Ae7
yVGtoFB38zrnGEkA00QU0+heoY613t/IOfds6ssaHjxigSQJdXtjc94zGypqc7QN
ZJExagZdZ5IZEthyZYcl3xpv0yh8sRBKLizKL829nMcL88QOFGl2G6GznGN19tZT
eOOvSfrn+ZM/LZpt/refMPBtQOrxY2P4rO+1ykM3kpbwbRm2ejIvyXHoG+iT82VU
aKLAjJyUpMmjMucbM4ZgroE/a8gYTqtzUqqhsdKQp54ZCthJE/tTyzPMu3Br/4LP
MschBUM10W6PFCc3irgpxKe0NL/alYIq4Kk2PtnO8sVuoWkjQuFRPGdnysrdCQ1q
SNG4vVqLyDv37+8l9ohc4PPM5Y4Y/0FSaJgOc/2PYxRsQ4ujkPjk0z9s/u74OKW5
3rs6bW5nrOEnBGRG1p3q8Lwyqr2wvAXETY9bTcqD+A3qEFvcVXamt6Sqi9go/S9C
haHZILA/2dGga8O2boigl5Nk5v4eULK/ItPfE3ZWa1BZgeeXQ+VQTtXkaa3iJbtZ
Vjl5Gmjm+f7hOr9Ppbsr18+YZLZcJcIPvXb8nh3aJ9NSXLVmVNOHRqgIRFyroJE8
fM10fVT2zdws1RTtUI7AfzHDbKp9gts3IcmFMWqiVrfDCF88CDGHaIv7MrDmYiZ3
pvVFJVLDiBCkcpLYqhAsReffRPIXY17/N76GCAYgFhBwK5zk9RhO82RyxWXayruM
URKo/YhGe7oecGSTvZTWSglhhya1sQD4IExGZRHmCKlKk8QOtdscSHKtsSGImi09
/BKExxuvN80jboZ59ZHqGMQJSI5NKo86T/bANTm5gGFgeFCmmrXwRu6nzbwsYKWE
oYrScYEDx2TM6gRen6phgHYGnc7ZV87sxzKhFnndEyWQZ32GFfz0AuE2wCeMV2Zg
g9MwGtKje73cJBROrUjvlay/dBUiik8TROlckbx6uVIog0TyZJk5abSDgxt833C4
qMB50hAK5LaoRmeKgsp92Iku7UDjF3gaYTNmyDkbn+Wn8QxEeNJHnu+549ovdj9l
b54p+kNPEHiafCvCWEX2YVsM7T/gGUG7Glfh/34KhQKrroXnieSlLAVD4SNJM2m8
UptYhhbwE/Ae0d2oggqTbG7UdY3tMV5xeYR44JStSe/wLdOA8znB0yxgUCzxxYho
ZFrQusg7WlqvKF/nfapsPiNnS1KxLan14EvWe7hnh9HRucTnR7hPww1pxNUwzf4j
w2K21OLemTcn+S33UeZj4b2yidxTXoRKp33ZMOmgq9vIhw/LRpjS7TPfk3UMgryg
UXpbat4L2CWr06JZAaKZVHKoTE+koUvwLkoaImV7Ry7lSOPMkCKw72xWW1drX43n
Xj03wivKYLwx3lUlHI/2QPVeMP8ZTTmq4wFmAkll3SQTdrGWOYa/zOr+FJFYPj2Q
EOWsvmRpsPVkKbk2sT7KmZsq7+TNzwU/tAZNTqEjDN3eyg6atyWA36EIufQ4hNtT
56XUsei4D5AnGvOjmVXooWoAQG1qs5j/azrBhcxjOygGpEZIkG4db8+eWRfb5Bm/
4pT5t6cLJNfnr9vlEixsNyFfDUajtMPSEypDi7AWU4KkZUXoRqycj5C4iBU9ylE/
Ryh8SEnFyP8IxQkmuBJOufnUyGkTRkyvl3BK5r96LVATOhXaD1MpYkLfsUWNYdpL
sNI75VCFaSgtbDC8ouYgv2TH+/oj1JlSgjMIdCTu9BW9sETqkEDAfRPEfEatxVQy
6AxXE7rArbeUjZxQofP6roz0IeIx1zELWcPbu0nZo5/a34YOc5d+wvepqPMb7Mf3
qapKUzQeeQNdvra398QaMNATY8BCo+0fCKPfegFB35FkyvxiZSyxDYBAXsENWbvg
zw87UNW1pmSXXDwZR8FrM0LFwbZmMXuwN+8V0OtFff9fQwO6tdkoIwIuA/aDw9/n
ce8F3WLIEHoKdb5oy0WPLjkkJodxB7twgKgiY/TMTHjA9X7zMX24QjdEGUFdr1y3
XX8cPY/KAxnK/ENLUpV3nncgMwJ66If9tEo8I52uy0ZjKkbCwQdVbcWqoMM2CivW
8NZcxTusaba/UNlDIw+LDG50A/ZVXlQ468eBUvD5C1u0FulfTbuE1n8GPVK2Gp40
KflO15+2ZZYe6TowNe44tjUhj52pkt4lYP7RIqQFV5eFw7K49W9Mz23yRNuxMby8
/fLf0sAldSlzUX6tsR3iuqRLri6OUymPzG80Wzq7XFECFQ6hBv/DJgsY/L4vmBRM
6TZm5oK/47YGzASrb3LEuPpjkfL+f9kUX9SBgskvV9uCkTsjtAnHZRmAqLwzWJKG
0NcHD9vTTnOIiI5eJkHJRGUKI++kavtqjHzUQ5teAQuWuJftZ/GvE8XWMzL1723F
OBByBQvYCp2kRaE5C/IIg3ASGiqfUnfcnAO9kR/tL03lTtDuKxLV3PWq11Ik3faP
GWTBlsWqve2SOmkQAY/4IUp7/Ct1IpvvQIT5gqmAilE2As1S9pjaNzyH+pkj+qdP
UNnfWsvYN/yvnnndL/bh1MOqYK5CBZghGur2jvBxbCnZ+5mFKGmGg/O3RTbwu0BU
LGOaQWH9rNLHj0PdqBbCSKHiZ+/eY+vvbd9IiJXytJRtnyOuDblzDVckC3njdzc7
IUruG8YScqt+GzwqiqDMR9P+wDS1SnCoaBMfHR9Ulqa3X82f3r6qETS9rEQSRC1r
pDqk3ApMBn1OxEU15XAg2mKT9WWdL1ZGISKNwDG5sKvQpwdhM1GLQNutRrHJAMIQ
Obe0QcYyg3YSsLMJFpTgkQt29Cj9nOjtmBllYKDwbLhOPElEmTCsNmLLjc3hDwnF
PwFN5czncEBWIMzwMVwjv+tPx1XewROdNLQyaxDqWx4SBGObEbSIWhG21JX1BFCb
0+zrcMnkE4ZWD8AkQ0wyXy07LXgNGxqFc8juAYvbu68p9sVKCsybbT18QlBj/0yN
BdxSsDUge6pV1QhYkU0vmBqOFYixWBlC3ZxyVx+FwOaqtH88EjyIRGErUnTaFuqE
3Ed6lReexzFlugzPIK3FZQ8K1HGCbgPe7S2ecL0OWR2jrhJ8isc+eDqQxxUS2z5w
KLl4uWLnVlEWrMCtRqlRPwvFK9DXyZDgVfrvnD2BwWpQ6+nrdIYqU6ZakT30t/iY
1S1NkA2P/LPNkpl4yIW/pjWKtpzxOLnNjOQBrcvpEMP1Aj9hmqBbGEbPrjGigRW6
uPwk11+3SXwcPTuuv/xR8Bkbh0MtSYqTeNwFhlVcFIGlcUjpQnR9zHu5afUM+IwF
fYJh3Lqzvt3bjlGCA52pJYEaBqjwvgVmpwE5aolNIeAXrvLWqCeMQXWvsKOlGScG
acxGPsWFiSYVDXEtGQOxc/0uAZ6Sj8x2jfXY+TNe7aW9bk8ShuZx1X2XpNzE/r+C
HrblB6OTDCAbLCfCzEl0D8J5W1JnTeHp4Op0A8qF3SIAX3beRVT+Bqlweab57A28
dIxa+467OFqEX/qy9wMs5M/6bI0lvh61S5pHUeYzxIkiHplAZJKLIaH6y6xVtm51
PSinRoh1EpSS9a7Wctfwgw9y5hqmsrOmhKLe7F7lS6zWo8m4gNbNfMk5rdvGFGyk
8sr+BeuOxaijzPKwnjW3c0sr/vhj7Sv6GdAHW+COkYs0f+cGKGyqJA2zq8/DyVnc
WxrLFs/T9wlyZBtfLdZJ7gyJ+WPMA+qYVsGI13vy7Y6iFG6/ew74LUqtZflm6KwR
7UgdV/fIU2P9NuC6ClqkvHqfBc0vpOwtaAgIZufV/L7affjvB15RBUmDnRp3YKP5
D+YBHXHJUrXoucv4RQdqH8F/0SiJ0VGC0j1f7fRmR3Lok2eaiuXTqm+2n1ba6RwE
blAUmNNy0toHsPiFHhWe5N204G+gGhD6K3AFJYP/Ehf55kpraiuaGzKAuo3Gpj29
SOlbIL3VN3epictzlDBgFJDh9LyKwswuMceVVYpTBKCE4IHLjuY5DnLHXUaf3vCF
7JWbxu8gtbDhTarAsb5tbsoRycX06a+nkDiSMUwbpV9R/U4PoqfSW8HIzgc3Qj3c
6efAHyMnNtuEIdTzX3zJDRVaU1oYy3CfWOof549Wwzcfw/CdtFnue+JafN+fCpwK
W0XCoJ0Cf7+1KZOTCPGgVz/mloOKdQVjp+VxXikrW4KGbmRNecR1YxFvDdncNoQQ
vsW2vgBB/gpj7BRwEVQhQi6t1Oc4/eBsEc2t2tVIr4YR7qALq/JBAFGgHrEspCw0
q4JaFawHSiuE/Ziii4F4WC6ySmA3emPYebytdlv5x3ox0I+XkvuV/wIhAQQx7dV7
ELhxLfiopsvKBkt6XqeLqhcAbm+pEihIxyaOy2dudAUxb7cFlOqwteIJcMdjSOJ6
OtOddoH9KxLMqBrRaGhYPuGxfpptl4y7B8Lh6rvFuYzAJXX4HuA1LmjoQqfB7mUt
VXza7fPtNDPsTxtySsY9Korbd8GyCHHQBUf8r9HPaFQj5PJISfWJQId/bLxaIlvp
GFp6NFXuNt7JZY5y+wynRwYOnmY0RdsmxV6BFrbW8caPiAYpFy4A+o3mqI5LgwVn
+5UVoKzfOBHfDOYmzNUGsTJEAXg3+6ZM+mtTYjqhNLqlEUkgBjJlRZz1aGmwqZ6j
Aj7qTRFCyCx7jtRmoeJw20ItR+L9RK7TisRf0r93U6iLcPGSmucczoon+t4TvvUF
LHjlHI2uahpLfWB+fJ2Xpn67DETwx1Fc3PvrDPHycodLAORZdb4sxquC10+KqDJ5
pZpdGJqzTkhtBSw5QjvlNjcv4wY384u7EXaDA87Zlw81EVdZRnIQ+/kJdsiqIdnn
bDKSPEVMRvKSX5rDQjidTyET+jhQDrmfZ2RWNg1KkyI940v+zKq4KwGJ6j5GhtG7
0F08ykzZMCmsrcWHO6N3Q8CPRZM6jU4rnS1bHpAzGIP0BkNIrSqaGomDXw6kNAgq
oRRpH5TKbbz6/GmCM8r3yfaDs/1vLWYuDgfDpHvLUgrMPq6mB7LdKS1UKGCsL7yD
ozZNbUzj4iG4keQg9NPccfTNEF6kM06c+7TcEaRaHAbvY4/ku4m73DQVQVAVCHky
nmaLG/jcs5A/nZSHuJkkAbIngQ6BTzFS29J9QjhqimW/4XPCul2K62Y4oc14i7cz
05U1UIhYuIC5I/QHjHTJQCob6LCYWnHlEvqBdJlcZ2IPlxMFAJkAQd8hcRpHuHMa
uDLQxfh7fEjeQmkrphl/VzEIvVXLze2NP5eGCF817bV2cmdnyQf/rspORnXDkhOX
Xza/iL6s5dx2gg+izxin2UqmH74eUJKb3Uz2o/ZcMLcQ0rAQrP3PxzaECTKB7KTd
wk2FlZ6IQZSIg4cI/CQg1FQ9EFxd/yiqlsUnCClmUBoJChTySwu60mj5fthwWmgQ
3ymddKm2VHFCdUiQjKwgGwRXJeHw5t6XYVXhbp3xn3v8IJw1zvoeNaqxAURhYe1P
jaRqVGUmQ3b7Mt1toUOwYe7+1kOC38hZZeIk6qIuvuJuWVYSkIKzHDe7f6xqyRaQ
l3RGSkPNlpGlFM0H6GIxZ2z6xHkbT7aQ+vHSUnY1+Ko0Bh2BePbFF4OpqrBryjht
qRKVhaN1m81X7bwRZqfvxqPD0RNoRiN//w0Cjx6ioq80AMO4Ko8qpdvc2Y/G/8iL
UXecPj27kAC29ugU7AqpnhgrBWiWPaWQozyTP3UznSOMYrkALcZqsfOKBwjxnxRC
aPBFwRM2+/I/RFQjRq1Np9uIliUCjN1cp6Zpq5X+UnW/yewLxhXBs2Ru6bvcst+e
jzHlMsFyB5Jzn5IIxlG1VjYdteJ8ZaLHHTMNRgA7uuoyqrzeSLZAMjNnNbKQ24wp
S2goFxnZ+laLIJ4/bCL6+Xlxe7JIDrE+sDXHXVsto50eX4FqQyG10zwqf9mt2DBi
DUdJycaml4kqWzySgqpLrGU8jeR26W01p0AFhlJ+Zw5IVCPF/uXceihzghuZubqH
fQzw7f5RSW4O2rkPnGeS0YHx6ZMvGlKhB3gb+NMEZPesiuVTheAs+n2KZ9GHuvdI
Z6xgrU+AHFvngSNh9NtBTfZPgUGa4xYpn48jfkrBtBY3hJMOr2wrzcjNVNSplSnE
dNiYKjY10pMeMiIVeuzP+hk8cLNIPd9IIwhVeZC64BZYJ2cDO8aBRoZfOdCiKm+5
bPRlUhaF6QmupfT5UFDGm481t9Op3FjM1x5KABRi9sZDtlWX40X1VBA7yCKaxF0X
84EzJBiCnENGvzcLt+r+FFAAKvZlZV9PoQRNAijwGi0/IJ9LlDAkwZFhOkJORddT
ld2add354UTxA9hUGWxXrwL/2bwM4zMLwKBrJYNOHSIIpx0cqYbjpABQga0uR/yl
Ccqhm2hYvvvaR6MKjimdMiE344X5IlcSG1moo9syt85Czje+i65WPlbN6xY29md7
CFzIgQ+PfLTt9z19RxgkdQVlonH+2g/t2/usg4PONsB8a8sMuu2if4+FQCcmbf/d
mtCoK/FLUXulbeOfMSQUIxukQutN5FeO1vO9iOkSCj+P19q9adF1Wf95bTbcTdgj
cRpbKtqRz0/0+glXwSAd1lzm0p6/sslDd0vO784Wo5V523uItutaNiIsn0H3DiQk
KRJo8CqedCn93n61w8N8I6LeVcHahn4vkqja6x+ZnyJgTqvE3uIBCw5bWswAXL1H
B3raaZttTzjmWLdAP7i9v5wlrhldamXTrr/RHU8nw9q/Lhmf00bxyyBlenkYAyBz
GeSybLG5Votup7kHPQC+QPt4Va9uMUMzKIr4WUMkewA9lw6hxuKJhh694TXPTyiF
76O95xHWu1bCZbaCIbmOjKEVJjUBF45QTvzzMUJ73ppeDerTHveOwhhLTnINSvFv
O56LV0+79W1/A9kgjVJBuPbCnMcV6Emg46TIWaO30BaVAj2mbRzQExwhkS/3P42W
AG9Gu/XMFwI6sV1qoAHXtTD0zVkdRkTaHEhiqG8nPPl91mImmF7iT3PnoaIEw0+9
7jlmaAB5xPhbaSDFMwMCYSarKNLHRW5SsqAayXvC6fCv6vO4qfwMsMEHFKRqVTXV
3ZEnG8ri6Q1ZS32l4ExrcQii97hNmo39AZFKdWpUT23ejhCcfB+X904q1oZdVYCB
GEsLZF2PCfQOkp2gDN27kMlCm/x1MCHV7cnfhUpccZ9snZ08R1AaurCgmGkDj2Qz
4Bbpgrn/iOCZgrO28dMeSmw5RM31lFBLs10I+8XfsH3M7ouPbs2Gf1IjMrNmJq9G
6xRqEZx4SoMuPEoa2bwDhQXaG4S6eGsMbULw+fRN+UKKwArR04AjxFOC5ge4T892
eXpRhCHN4r+MNkBb2xAg/IrMdqcFdLv4Y8Bs/78lDKcJ8QoaH6voJbdvmM1mhm6Z
Qh1r/MlP7BXZyWpOWimjWdeLIEL6GoC/3H+2rMcJsgJzMQXBmKvwCdsQjnIVZ1TI
odrj/KoEOaiws37ADOy169XaVGLGbql/KUUl48ei+h4KUpQtzHMCA6i75njfKtIS
G6QxzSXKCGo5xCrUl5zVC2DOMKaxN6ejU9ucWAN+rjKAz6isT/nOcc34xyhuxKiQ
H/mffHfcbaPSUfoj8/JbF5xQf9QsUJVvtMiBnl1ha34qzG/3n4LRBeDTonH540BB
Y7lADlwoJDnMKKo9cSLYE+mOo0xZqXr24MY2NG3eRcXYHSzWVsau8N2Jxa0zwV8/
VgHN6uKiPVYVujMY653ijxlEkEafy7lyTaf0hWnon4UUJFm2eyfqYo3miCl6m8jm
MXwD07tfOhdh7u5QdGpPlnzbBrRsXB2i61rJkcNOuOOZNgAnckeG4O1lPsoS7JO1
3+LjZaea8q48eUTX+sO12ZgMUPNkeYCmQc844IP1Da1CtiBtenl5p7ZAer2gbs2u
kB4w3Z2PhK2v85sSguUIdLIs0X/PrcxxMzPkYYsRK6h3tlfUAi0UlmPt184RYGDN
3X1FiHJ8UqvyFWCGO5Eobg5YJfKdLCdUgakR97XlKJ7lNN4XW7L+sKyrcy71l/Rg
lnRVNw97AIIlVAXV6iTvMcln6tuHXRpmzl/IgjefeQyoztHFaB2xR27WdPq9eYFm
AHzxWSh9kg2x5x7tKQHhNKXDH/nD66astxms8/vFpk2z4YeUDpDVm7NZDncPR1NP
qBJFyokdmci2wEaTb2ZTBMf6hBzWfiFsbhXgGPfaowmPgZ6rT/V8h3YmbkwR/v1I
/Bw2TZqnSOARxXnLy0HY2JtlOJIbretzlGoCu/nfzm/dEqwZ7B6xqXK3cUc3MmIW
XLdUnojuTLJq6lahnyqgwM4zURGdHkVuRFxSRykRo5tXFw7V5A7Qrm3Vuj6+ffwT
33fw1zWkcEM/gO9UzFC+lHFnn47weFa1Z+6VJmPzOKD8dfRLgmEfcY/OboFipC5V
awL3WQgmLdcohognSNxq7B7VD7z48BfLC88a1W8yVG61m4sa1D5CQmlgZLUMZqCk
xym1+Q3nrZIigBFfWb4KvkKVfsAVbQh2GVlI3v5b7zdCqW+ddCjIeBTPf0F8/u1v
Bgt1o53z4GVoO03Af8x0VhbcQx7lXjldnKlh1rSvYKyngONuRs2KnK4xddNe3rnL
NwqlxVhvJSRq6l8Y0tBH7fLI+lDm2sJusd9i+XH6yiJMruNtfGHB7LEkHPAZbQ7Z
4RCvPyoxq3Ri6/rc0+WpxwYkoZmpRMc2PrDxfgtx2V3e8KZ6A7rnVafHVDc3BxK6
4nk0OhxQgJ+GvSFagXpmdORdvWkkgVzjJSeEfqq2Jxq3DSB7IQXpH8ELyTHk2N2p
TiwVvl5gHD9H0H8kleE+cqWxpxH1UPTXqnB8GAVd9+tpdIkraYRWHD8PYrtfiOQX
FLGyBnWMyL2GZHnhXSfuyfdoFfuVIEnvnwDB3c/V/Ywyz164eTYxCud14lGe45nX
PAndWqCz1hqYh+8BT6BaTZr41dxdkRasMjdVdeoGDiNLd9osaCC8YcyW15+7E/gf
Uaz0htuufUBPkn/7z0UA0MnpiJc4E9IENcMv0Nfs47Q+R5/4HHCCSFWn5WDbDJ2t
jPCOGEBzSixrq6q2vNXcpoUItiC4sMX4GWmAogoXUTTfG8d9gEuZiuS+qAPAkp9H
WqDQFkCqV5NUYX4FBCUh8Td6gDHKPfCoqLIGrQu3/9V3IVb851rTE8LQ2EyGjdDf
Izo+RnGnwFyrt2zGJ93GrNLJl51Kv2T97uZq8cc/wYPnMsHKXKWM31HE5cVxlAyn
3Fd9MDapv/7R3dDj/oT1OTkI1abRQkMAnt13JBOVwJ9rMA9P4hyLUbW9zETTW1FD
gv9rTQ7i0JGwimhY7pT4hkZA35uT4d2ShqHonbdz6LADk1mcNNLwtXYgVHh4wY7m
zGCty7Kk/I5XPr1KRXaCp4x8zRtN96kx9bo38IP3JZ9etKjrzQ26tTHhDjQM/umH
7BJhBg6DrzJ9OPxnBJJ1wdinaZAMePfbQJmMMG6pIgpLYD1QsCPl7SckIH23Llv2
p+Rdj2P4Txk6szdA8HZ6tdpke+Jhdq0iiFt4FmV9MbTrYIDY4VFscIZLaSZVJbpV
+7IhU4KJpNsq9Lit88Ou7eY7wJYIFw/FSRSh9So5vQm2stx6hSfVt7qHttWKg8hR
+J9SjaukAU5Qo70i/O18NVmqRtYT34/o16Yi5vD7Jv7bBAik7TO2TJUlA1VxZsnn
g+cnK3vgi5i1zxARB7C5d+yuwdlsgZ8yDCJIBKpjEcPnUNWBEbnm6YVNQduudEaB
Qw94LYg6hpG1+nsDyYnjXeN1xVQMfBhcKtmEr4gr7VTeSHiQWCenmt6tG8aDwzmC
RScZFYCw5D1GRvSLOB/8eWxhZ/nrjkyklOSVOSShirwZ3qkK0Rth/hOC0LGOotUA
KSdS0XmNbKQFC7C5TabrTt8+C4oeMdREIyYG0pF5TraMdNwn/Z6vCcPgy5oqXfQo
SbKUSBnHtAOMwGOaLNGWoeA6K0UptlqB5Ur4Mqi9SrQPn7zxqaCFQh287CVFzQiG
YgK65GYgHaMXRtf5Dkc9paDZbM2pj/rYB1JhLvFyggfoRuubaVU9PT0NXReJJ+NO
4qt7xfeWjfSzjSwFCjEAUxkhzwyi/puGOpAzigITWHIf50WIbsp5WYbuaNDjnER3
qMFTZQ5v4pSqcE0z011oP5ztBY56CJxTcn6dZXk+EM5d7MMfPCCXdogSEVHIAqCm
IDfM57Gmia4zTun3G/AxmwkTJBWUN56bqH3x/icXUSv80Ia7NOV/wva/KERfoQ51
QkChS+Vew0Y7CuLPMWSKEqODuO00prc+r3hRKzfAFn4IsOqgv7+oiTw2OqgTtd3v
MH5qKDm+UbOML2impfUtDx5ljuAE8DbryRx4akWZa7a1gVu54W9HSITkzAbnIyXN
v57cDb8OKoOvF6/EXVC4IB9nr11q+wHXya0VDpmz/uWvtEvfbxjFOMKLym8Ly6+F
zWMpQmbxTaY3ZtEhJhzlS481amoKJk1Xy99HL/6JqU38I+cLceBYfTftXw1BPqr8
6riKPQTCbxXeY/vkzkcL16KWgtjqYxS07O7lllPQSca0N+yGFEO5n9Jmmx/7+V5X
h0ej/SRAoXBJ38jzJrvaRKR8OKKaIyqN9gHlVTo5bC+Gqy2tGyOppyUk71+WdcnE
vrVyU1CynGR++BgFLPsZFLhGkmdB5UzVkQ1TmJRYP/QG7UDfO8GBxaEe5eY81Bmi
hUvtQrbFXBAsoGQ3jdY0XWmkPhsMw7wzAmBrq46Zzl1+ZcecAohU4d+XxVhFHJOg
Byfr5y+nrRUuwVIZOwgkQfBBrAOLVUWeN0pS2UdBVluJXTdS/iKXaXQikpBw76dS
UQ3woTEQVugLYcp1iki7wbPHzSRFsAh/i+giT/R74cSxf9dgm50FzEb5edR5zLdH
KhFpcd6YaugYLW1z7w0u96nwtFZbxe9uwWEMqoZFPzYpvmbydxMnN9LtfeOPmjao
6EReVPmpo66lnkSLqXtzB/odAr5HXXRJkAsBvXMdnkaAhMb/S5tzaJoyzcDJGU/V
ZBKWH/DhCnyFZDOJSI7c6AD/P4gBctorUrulhaThrLIij0wR/PeuuA7t6Hzby2H0
8OLmM03hNBZwEWJrz6cxkpD9HU0HkO2TRD2C6iSueKIE1prBPXc5IC8PMjHXS/W3
ntTPJ9rGhR9LK60A0iXkFyOz0TndT9hcAOX5sBdtlQUZyOClPYCxZqUC/Id+Srtl
dqURPF53H9SuIaWl3MRTYs9SvW6VUDX4nSe9QSUGcy3sCPZkNooSBlATcK3vGSuv
qM46irwFuTjLBy9MN2+yy+pZg/y6ECAFabubA6q9DndRpB/0Baeta7IWlyoAkUyr
Cld1ETuks3dv/2t3Lg2MHhg6qMOSKw1U5cDvOvLUfgVEg66NX69ljpkUJLrTfvW4
k7tu8ZHoPNVpBQtH6hkKWNziGco1UMdVICe4tZRHWl+iT2YqVQ8ob/Jg1DYIYIYl
/yw6MMNEhI9S5VBlWEo//C6+mslDyvlqo3Z4qx8pdew4C6HsJKAIQ9rEWvjasTG1
mOx6rONA3pgGfyjATmyrRHqSj4vPQz/wsZP8+195t4LL25uR/yifNoa5uap1cnv3
q3PJKf2jIPxnO89LHIQXNZk/Aho1TcLHagDtQf4uNJagX/Hw967xCnVO+TyNdVCU
H5UjXXLdifEi1YhrgdiqaYSNXxrpsGvP1GHcztRVSuEu88H6/zYMzKuxFqUVOLkc
fjtCd8R9Hzmfj6i37pGuOJ6uXHGXXh3w6lU0c+4ZszQEp+KFG9o3J0kkt6henu9l
4QgYNOrh8N5oQdxcTsdqIw5UFdl34s/VIUYaxPZlriqJH/ujSJixD7A5iIhHXEUb
3zpccz5B8WucgHffjB1rprJIaObl+9wjBfJWDYQ4lb9YdN8eEuV7tEorqnlYIZI5
plov/WqWD2D3NimGNYJx2GNPnDxsvczj64qbawA0lOR2SvdzhDx58HUjeoWL8doo
QhKtCckNDQb8R2FamMr7aYOEHoSSkJU82zPtpC6wapnrA7UkrmWZMS1uTx13Pbfg
X7hRIqng7sUJvzxBw2Um+uq+8x518tDKuIi7op3a8n8B1gATkHrq+Mr5G59RXr//
vhO2vXhDTHedYvG/VEwjsCo6HsTn6zn4m/8zdNBpAngzF+NT+gGBTlmaV3AXpP/m
VS4MsbTgs4YOpKLTMNLYtxSc6pW/OUI2AgqrfozNyUKPUgNnXWUIZRYe8yw3y09n
D7eD4Ok1yZDMzNtIwnkrYTlizr1BK4u3NZAaubAoS5nM6Xrj9tAeF1zDrjWzS39I
nb9sKebEyp2FSGJsHcOZzwUrhj1lbv/PFa5Un84cEiaAkhA4WlOunbMSeBpyZt/r
DpUe/FGYSjAJWliDzHyt1afx16ziROWmIkUpRq4MwAVTze2p8VVzWm/qVOLcH7tg
eXQxravrSqx24Uv/IHKl5AvuWFOMdaOhM6c3+++j6cL3G/ab0HqGM70BSxFX9vG+
sRI/ShtsyS3QsnI+zyF0IiJ9JNKXTiH4AqsaRqa4wZh/UWc/pVv583uBnQdadgGw
3OdAweBxPq+Amq4oSDWXs1ScPMbVUk9taqJFyPXsBxeitwvhfi0ZVQc1Iwq2D5IB
oOsC+9M2hi+20KDP6l37/kRllvx/JUqFLcgk3g9M0MYi8XUNLXrGc7KVz8R7n/E/
bUgo6Cmar0KLsfPVdbELJEMbXzIN6TOZ1rq76wKM8EcEI2O0SJeG/p+FB65V04yb
ovT8p4K5Fo1sWLVMo5IBvpFPrcGEZ4y+L3nlvi29/BCbkC5lZnhzbbZ5omgEex6V
FECZ/v83UC1CwTm9OdWRH+/NR7CIcG/0jj6CUPWjZWbMDxCZcay/DCaLWLZdlw+/
HzhKOabzIvqjdEIltg9gdxf0M3tXR5hbHH66iRooU4271coLW+86ao/s3YOToEJ0
BgviB1uV6nkD6evLznlHdZVFWXJ5I+liUWHzRh9YBKrXm6Ky/1MNODm3YkHrUowL
1gqd22ff1b+M0S0cONnRPVvSN9Bzoem4FX4vuB5AkwhyDDoGNsyvbQwKk3H6Zivp
dM87aM5JPJyzRfk8iwFjQjL7sBdi7bGN1KGvPzvAkZU8xJ3qk/cE4exSm/1sBL4t
GFFNbEhicK+BYqwmKKtcbzKld5fiO3Mpa9NmEuW6YEaUA039eHn42RZgHo67+5eZ
VcFJRIBJRM0CSBvTo3kjt0ZamARmcj8e4cwQFLM4LqfJth747GRF4419Wazr95js
LM8AsH70WOFAukuy4hy/N6W6imnuhMtfMguPJdRaMLK4dI+mNEF8TkuPbAalkxOz
KQiAFRwgSUhtoqHn/Y2DqhFDFspvdiVtMg+HMEnHtorQO8IMbgAYFb6EW7A2Yueu
PQEhujYlU8FsfK0QC/h69wFg4uNa4hgUIRutoGBjo/xNBDfDUKJBejLAuUFAl95G
piPT11P1mNZJJQ+wa1CmumOi1IRfXqGzs6U8zjeDDIxmdJ7Ad2oFtzcKTk410g9R
gTUxPrDWM1vW4S2X+UKbAmqwW8ZXmrQtqhJbbLx+fZ1rOH4Vo1Qow6DOTT6dG880
GZNepMtDphk0eR++gxCGAfaxzUfYQz9talib1oOO+dUznTZQPzgCRUxTW5RMVl0g
JqL9WNhuQL3C1wWrCzijQpkbx/pXwLYIpTRB94K5mIjslg9q3LgnzYWwD9UR5jvZ
/nulZmffzTL9UULeLgX7TL3V05Fy8ZMpD9eQEug2Srl/50r+keh3ypx+2A3FJd3l
PlTyjiW3XJp8pMNQXrKm2Bsy9U9rkh/M1A5TGHXdPpqCTtOasF/zFcrNeCSIwnwe
kj8Oufa6DOwIbO6hf4JyfCkQugJMR8w+y5cQopTJH/nygakIMyZD0ZHieTPBvJGv
S31l2RxE7+mKWAND418rDysM/fMYp4nVSwv2Fn+zeKWpgvGUC87KwSm/s2FuBS1c
ZCwReSkeKR2SLfm+in/Nm0SBXyW3uBkZznOAv+SoIx0jERLx+fV3o3M0lJxoOK8M
D6g4FIY2z+BXz/91TsNpBcfma++xWYsA/VPhhe7HUexat6WxVW/14WYbadT663Oy
NVdEn5tsModPN+ki4IPeAxYnQ6UsVm8H4di4EIjZYtiWRO050gc5bbTGYccK02kr
GrMiAvWy9T155c+S2V48tXxgRxepGhjIhP39o4o4CxiALEHcZSaA6EhrokHB+0Z+
tRkSq6YyetOCiqYFoJtX5y5HfF0STd1X7ZJABVQPLupbiGVQcbNZ5Jv08yulLhMC
t79NABfvV5jfNQbJxD3cym1WkrbtA5rXDZPYt66ULwoCHn1d9xzuvf3D88uSFu1d
f8lPYrm2+G4MwHQrqpElr+F8JGLaJdCnpCxBnR2LkY/xX6V4QkcXckkBpzfGtYNY
Ek6lkRpNNKqw5YFlYB3oNhCcXd1Er6X6rq3lcx2iiqq3Xm8ngoqB5CgCnGJZe7Fz
4savaSJigLleb3iNi8w0CJhBFhXRsY7YVABGbZ63PzpfV9jNro0b6JKxWxkAn54r
1lC4PLVesBquM5+B6xoMNTv35MbZjqbYpRHpOG07hAwd+wuVSXiEm1tSYpU0V9Wz
G3qDHAuggG/HIcLoto3P+3iVkpbZnK2K0wHIp0ZmCzNYBg5hrOZ4Ww1Raffe4YyJ
9m/bPDBb/IvJt+pkZXnod7ueo9kEus39H4J27IK2qR2O97U3VBmjZemyvYBlzZNK
IscN6FdRIOLilIXFvkvnLDpdTe7iEW8VPzYLFw+hGwSYjI/hLX6JqkLqjiCgbCr4
XOCNkO+UWvy9yC2K0BAd4q63TOBKxFIxBcsZ3VmbA0uPKyc+4uAB18AjaAZE7609
LyYpQSaVQWA+9WN9UhQSnN5b+ddNAZ84o1jjHZXsmgzkVsOq883DdoPpyBhVL4z6
+lLdPnUoCbPdp/T5qdw++oZHAlsyLRj0QrGu6ZsLidvRKUiRco0KfktaI1ycSZnV
CwNG5cu2BfajnMfyqaleer9g3ofMgAKs1Rb/iy0FKC7TzqqygkzXwKjS6e2Jlpf9
1GQVIHsijv/wN7BhHMqX1MhEHpZYeL8wGKTiYxbZp1j2qYKsGOvXdCwy8doH3cfz
C/ETQ13iXz2H5m5Ox5pQoKnB6A/ltOropWUlPBD6Ip0hzKvHH4UfCKqwg+lgMJmt
t/FOKxlu3Bi72TLThyHx5+Kpv+ek1CYMHEMm82KGfnrfpkOBHqiTtg3Ju/+jYnBE
Nr+QT30a2ehNKlI2p2JdyIf3/Ym0+tZRWulVVHplEVG1eN+gUpN6BFqSgKtQT78I
jSVyGBxNAw99eUf2dQ8uAJJqCrap2QjO3OWBJf81Vn77ZDtN5J8tFPg8+HZaJ1fM
7FK8HrRPW+AePgrOof+E6vSnxdX9Rq9XtVPOHbmEbN15PQe1usBZLbtL482/IYeP
a9CcLpIoJQntaU60uXcXKB1bwY9PW6Hbkr5IbNXwtJxo8aYDs/amRI0t6VTNs/6X
uGbVZtIqqIAVolYa4ppeD5VFokppxzgawMZsi5XjedmGALQ4dVZV8JneRxtlzMlE
DkaGaIjg0Q/rrMFJXzLD8wHT+Dna8qIfS4rb8zfLwpaj0fMlHug5zl32Pkm67dn3
cQlnd/ujGHQkPzxEUcOqDItaWO+IVFC1rRhBo3J5vxShOrW8jzisPEGLKXR4gAOr
FEzkwhAZbdbA64VhBosrO5TJh8gv3RiZV45qhiaRZ7mikMw/hlLXqaBbWydodfnE
IxEhCOVfoizKOZcUdYoss0DxHKfLDzqOsl+sfJHZfYkyFPzv2iq8oy6E14wbS5yi
2rbdn1o0BkYTbmXdc50+7Yvt8ChGSBaosGg40B6gFB35bTDXEshCOk3Oh8Hzi7bP
swNXoE+lYEDR+utYd/+1JG4i9aIbjPq2UIgHbmbXwoYPKIHEHqMiPXSsmif5ateZ
UI54bUeALsEbrK4p9a0oNF5KIsDuvMi2khypgVVUxrwH0UkIwoZL73dgN4+K7udH
wHeGuSwYN3VVOGVFjlnPFrMzLBr0A25SypkVvAYQmmdvlsWvCeaoFDCJ/nmb0Fj6
KU1SP/pOS6V/2fgPoRB0Wf5jJjv4iTYWZr+CLJKSPbse3uvChTRXjNEBmqXwY3mH
ZFBg3/hbUK0CKCe3tI6iRMWSkOSFn3lklMxHCK/vKUEk2DkAV0ZsBOT1FUaHbmWv
RQLePn0xbLbLUkFekkTePHNyTmuJw58w3qLK5hn95Lh+ui2j+k6SvfVR7hxfSvB5
yIITCM1wMiSIvZL9as5SU1eDVVO5kIrCjwGz1eQd/UsyGpMqvRIRQU6qqZZCeGSa
QXVamWzEBJheJgq/7vr2HezKpIOBkOgYi+0LH2gIplHVJNa8HKwHBAQFKUyOO6kF
mptUa1RRrHIePyOx73kwXZoU9EAynoEP+1NSMlFMHvj4MS8a2mSA+ht2CR8NZRsQ
evqckTUY2vuX5N5gabdd5XzmGjjaUnU3XTWNQEfq9zgVYZIF5jR9b0XzA/B9Ec8R
PUre2zHguvxRPXcg8iL9HGeKfzWSirxn5FwHIDTyVmmwGR6Us9guTT6cH+8kVHJN
0VBgtWjzR7IVTvDkPf3DMZKVjCUYLko1l+ZJdAUmIXoHEEhEUwiJsglkGlhm5rsZ
d0W3HBQUuXn+8ND+GcFC1IgQ/htyN2q7V6QDBSSJiPj8wZFTA/FrR40JlAxUio9F
C0vbVgTdTZ5KRNwS6qy7H9ve08QcdEviy38/nNeeRrQb6IlElXOopiHKLJbDpKal
j8xZBgJ42E0mMf5SAjs+8FfrKA7pu/Unf1GF0Isr9SH7V5AzD3KmA1PP3pf1SPkP
sS3cVRs1cNi5S9OLVbEriZ08TvW0LTegu5jJewUGXiZNIQjdC9OWiRo0ZVh0CHEJ
xKFenYiyO5IvlwX6YZ5G+qsNCddrK5acomGOhngjs0YDTDUDXvyMJGrAdMirWkZF
vlF9jze9VM+U+FHg3PL5xyvT5q+yJWQt4qRC15DCTr/wI4S7bxvwHMLdvZqYArqN
qfoQXmGv4ytGZ1mZMPNU5f27optbJHgAzr2FBu8bl9YAuL9af3W/G6LxQyXCEtcs
Ep9pj7T2NpkzijL8pmgmmdghe9kDWygsjXU25a358+HVF3OO5AttUu1cDdl5qccs
fqXatnqyTiT4DUREwxrRtMGUYj/bOmu2Y3bwfjZEKd28oWGcbaaAILhjTv0TdMva
9ZE1H/3c8IBje19ii+Cy2tFB9btfw6In44jWKviYZRstXacnlM+fEPQZ1IgqhGR0
/+3XGo7koyetNAbfGdtkdTKDEox3U+Pn/wjsZTSJ1vtilvu6P4q68RqgZhMwL2bb
b8zH7mawIY+1n81aNSRkvZIR4jTWkBGavvv+oZbO3bPrQw4dYxxSjRV8AoJYZDjW
Djzjkc5qrjHYLJeQ5whjOCREufetA+TB3had+SxD+GUYo6+S8C9aMwZy30FEph7q
wP+Zz5g6nrx/gwbqG9FezSyz7v2KnRkll5C3kk9D7MPxj14p8yB2imJvtx6DI+PX
x7RGZt1Bcc/+4EWcZlaNTXLUiXaTMBbEBexNkj9uKci6qSlKrTp8yZZaVGKWuguw
CLOYyP0ipiIgJxZbiEltX1AZPimiTG1FOicQkjRwZOmMdvAogxUejczEMWDuUMPV
RDguP0iix0MyxrvnVWlS8yYyAgqyXXCxcmKFHxkxlZMDdV6pALWn6kSYc1sTzU30
AUqRjoZZAqATAXreEYBNIRKkvcbumIUYzveqOjD40DvZxgjbS57vlXMQESiBuFgu
vl8u2PyQOGcFD0fOJp5wlnTVyQYG0MCtBC09z0zgNTTS0ITHVCKvHngY0sLTQ7/q
Cdcr4qOEWH4AcwP31gtI9ezZMTFzaG2EN5SGrYdArf+PIGyDWMIRJEkO5IRmnUsE
F1gVIGpiAJPwweti+gf8t4cbhNe2l3px57LTBd/9iqSuagl++Fs5gPt5jYgIjF/o
hZ33guYeiwkby38oSp6GVnB7cqXBnO0Pa3zZRYYBH8GRXmWiVV51VMXcyebhJ46I
05/9brMKN+uTY48bt+l3UarjH4h3QfQM8HIBk+OAUog5KkGgVUKYJ0O/APPe8XyD
iuwAMIPEVntcaW8sY2rU/MxRiiI+Yn86o9hhtjp0KYrU87/gQaF3dqvnal2QxzbS
kVGvd1bz1mSkOHiXcvSNC4b2rKW4rJGIzZX9bYvr5iPTn/2pCu1Ltm+xuzJhO/ij
2J+7hoQNjuiwyVStIPUB0up3pb6ZMb9I4Am3xsufykqp/X3Lg3Mg0UMIKGcJ/P7E
+BTalBE1bcK2gffT7gJVubUlhPE4JZoFi8FlT2G1wXMyfvkUHyIcW2UoJByuCpSc
l3YNYCR5MLE1Zrxu2dalus30welY7gev/NmAw5AIosgwbAK5UG7TPrv64mbWd3KP
ESpum0fvsYvGNwTcfxAKnec45QS41fPYXwEVefTkzgBXCWWQaVbZ0mhPtRu2g2cg
Q1awBB5iV2idP9PwFGSH2434Bb/X1FbUum8j/cl8CG2hKpw/hyN3OAJOjE1OuLaZ
7YzcbjF2o0QWoyAe81Twyw32vdcGMSvJracl41hK8JbUycRCjZ8/omAgxr48K6M+
vy7hoh6TaRsPJF0G7ULO30adaKP6SdIkpxUImBD6IiW1ZSR/LB7S4XZEOreV34ut
2mchJSESHLGGF1iCBljuvsl+Luu4Eea/BxlfnvnqjVvUR9VVWP9zyVDUkOeh0R3l
7VMz1NDDAcdnwzqewPRDL+Kq73x856Hgz5H2w94Qub/a36UFVkkMPS0z9MlvujmQ
G8G/sSK3nJUBrAjX0kY6biOvFU7zmEBGt3RWEUpSNbIFePbQCYw/Fi1EizNCRdJs
42WmciMeh/2Pi9qKnjS0ohcImIuQIl9q2AjKh+CWB4HoFFkEyTfhOIPCerv4tWM+
UWKclkmuTxar/0t8uE634MzH67Ykia11Z+EggtBcjaYxKGDf2+9h4Ih0E59HtbhA
V8hCoYk0fQ2RTUeUWusBg67s/l7qRZ8eW5s5OgdGVSQ3k8mrlgpTG7je8d82SKaj
6rjDtsYcYeRCH+KFqtlu+FK13sC6j/s+4rW7JjNKcOXYjz1uLU8COfAzyE6sEn9Q
YXCt5ko3SRot1oqiM9qMKnj81beiRoDfCjwLjcjnigS0uoV5c8EgELSL82Ch+pYx
TkcnrwstlL/O7D7u2+k0cWkvV1rOOfaHMFTX7F12fL9P3Cu5qlKeDZ4qWEGRimk3
M20eIAwEO8kW6TaTEUYbOJPxNFq1v9VTCHp5ZY3YgrzCurR8rLbdvYPY1xUI5SRg
heZdvWffCJ8KRrx5pxuit32wbtpb/zC4OHfuOQPEVaG8mxBp0qJEuuZd3tJfdsHg
SbDHgM7kocuSD8vbl/IhCilljMgY/63+6NLi9J96AZwoELR5G/lae9/S+H7gj998
loH1rMD6TbTssy0o3hGKc0At/Fp6S59GKtNWYdeMWG3uTn36MPr9k4soKFcK6gNB
tXM56LTUKEJR5NbI/4E4ZyyiWdF3VJIJlFHONHYlb2+y3GMsSRdkZxNVTiOvgFCl
56Qgws0KqbmwxdmF1VQzucIVhiQDpoRiV08el9eZXx0JgcG8imKJiO6qaMpYC+wH
wDvctDFOgx/exPGy2mKBqi4k1/Vkz5Xg/wOxKeKMK8fonozMyYGzz4qA708eV0xz
AhLchSA2DAJRgKhbjwpkn5lb0dt4wGCU93OMAQSBjY3u2Gek9uL0+kSZqCiERqua
AN8IbzfkUgpyTwb9idxfkTOnZnOzkSBPX4JFpmOwoka3RhZnxd+a13aa7BcHY600
tM3vhbn1I7m85Q6BxOo9qQ4LCF6tEJgB6xynFctkLMOwa/KV5/UmOsrkAOoI4RTY
eqV9mQdy70g1TGH90XNAfFi21kY5L9eUOSfmMLA5Ba5caLdBGLILTnE8Th18OyqE
pI5i+K8Kv/kXLZCKqL4EHcAXLlyI9oa6BFTM+FSOkT8N5IXxs2JZPrwNk+XDHP80
sN9QZIBsJr6QDFAL6uy0cJnTQeQVQPrn0Qu3MYaS5Hl7Ia/NtEoBxT9Q+++D2YK0
0cMU6y3LStX+n4dchoY/KPJIpUQHH98dFysRZLD7Bjy2VyWEhpknASSEEZ5cetE+
nEI1TrQjJ5jKGi73zQ18BTrHOu0SiyIuDJyT9y033YaWHkwQIuttjC9S4/frjgYe
p3BmcAoLhaCfhSI4ysGlpZm5NzOp/fjgiNwlJ2o3oSq6SctzRVzNuc1L6U8qEYrm
oFImEXMLAwxJfIkXY/Hez++gVlpz08qiVkYycl8wzV8u4EQrR3eyEtH4Hx7VTrmL
EOeKCfwr1HpNcLTWA08A27EeXt/3Wiw1+rX5Vc8mXTk85MTthB5LEVUHgb7vaOHv
g/GbQ1ZJ3e7R+thMTFsw4KQYOAjilYdexFTURq4yrCn41Gs7CuRDQjyMN+ZRDyiq
R35qD65AKS6JTRZ/o/fr52T5EFFgLmrR1N1GQlJyBanS7a8xPqR8tJ1vmbyByrTn
qvmV1Mn8q9c4mqyMEYG+vCDlo2Hdu3X1qBHC4WlWuz/f4wd3eCjnzu61YWtCLvId
bKvoMwR18FZzbpEju6KHWrplP6HBDyeXXYSVyYD3cvT4kuIqD0+CaueKgf2ajMWB
z7q/rNlS1LKM7nU16wti9kEK3VELV4ltpsDGDnvyr61xeyCPHPb+spv8W8cO2TYF
2Jz6rbGkTDftIgm+h/CoyvZkDFOq5G9quQllb18JrDoIe5lp8dkvSm7CwD9a69PL
mCZkXkH2/8pmUiPiIIHh+mB7xvYo9GPVUXyrWdJdLViAgRc7Hbemcai6Cobm7pPW
YAx/F8JXq+FtsnDOF9VgNpmr8eBuEhGTNtAcNa800+Ata4Og0BOEzYZdVamwB1dS
MagKDPJw58nFJSTz7hhFNKP12X60K0T5kPPKD4V/mlJeJZpbEwx3D7ZZ3NPJxkGe
gMq2LU9V/8AEM5CBJQug0I9QIqhP2ogmSR/G32SB1C8j35JkdUDy4eqC1UOcPQcm
Y2C5tAXQSEZ2sYAXmEQ0bsT0QgFZUaD0LWfPkFeJdTIZ6sD2/woTwtJVu4AlxViK
FanDUF+3orJl9lDV8Qh/jprRxiRROOwZkHhOYNBSKFVbGc7XayxoH9aLsmx0Vg+C
400WmHCKLeoWLFgHDUzBgf8wDSG6vkkusqeKHSf1cz59/gwoxixMxsvtMJjLBTLm
Rv8Ih36a1+k+5VWPjhcsQyrN8MSl5SHY7H8YxqbX2NH8XaewB4FYF5txPVVIHL1c
hSv5MABHgW0cN1kNh0I83KDZQYoBSBYDvEs2dEDTU8Fjz2NGNG+60Y62NAigtTnB
Tzy0yT2+FtoTWEZ4htfMiOnWbEVob6xDxEEUpXpWawcEfCaTze+LaSUEHppreS/B
Jx/11gjlLKOOHjXsnAZy3VQJpCsc9lU420xOjY+JUxsxQBvHjIRl8DC7MjKzTxFW
Tp48HnVO3GkkT47ETaa8Csji2AHKp4EhvukUmjC8mdrVZiAMwDvAljNkAnNJPGcc
JefUyZtlNFlDzKUf2sYr8Q+QEWArHKEj/1Q1EM0D7epwakH3zUEf1zH0Qodar1NO
nKdGHMfOQ24OoyNOo+rbsHIFqeDxRtSTZV6vZrq8zpCOU525Kuvz/8jjZqJuRYsJ
4k0wBI5RpP41GTDIZvO5r+w4KhUPIQ0G2Rbp1cpkZ2J5hqMmLu4sp21GychvRzwb
zZxPyjfRIEw+lF/MEzA9FNibvGLKZgXgsOKjSNUtwBWCmADxVWGT6BnOk3htsmtw
E9jsfi41NufLbvbhfGwsRN0HF4n6stuwHAD+fjBYGuNYgJgAS3GgBKTW/Nm8X0D/
iasM2rMTwiSF2Enr+OsQyiRiVFwa9vsUINj2A5rDmsayc8IYqMzXct0pO0ZHkrKx
m/S/5V328aGb9p+DNZMYdTzAE01PHUcbU26onuUW4BDteqdlMWKcbq5B7lXYqdd/
QgzppFc2YBirexHvy2hABzf4TRT0pYSqFkLpcJSPv/SCtnv/Q3kX0K4aOULoXrEu
/0LB4dm2z0nh55sqH+1agpVRNpJ3x5zZTICJO2+aDo7HfGXxxBTn802YSr2JkUtr
mfIMmojP8V9gvgA+rqWw74/nWZC+bMSyKTCFagyNh4yJzoAYeY3fdyAZvczuJPND
ePxR2g1GcKd3ZumJRe439RkbIm7f4SC3xW7n7aiV6BjQ0cq5XZ1PQGmvFDEBTPpg
0287HFOOOIASTICe9IaWbjgwatGAd0HLwwX5/NNl9mYCjqB1RclGp32wghq5k9n8
9S49d7ctkrRK1TKH49BscfhoB8XpEidDZBkPa/WZojt4Zf6g5LqvKfC4MN/xPyhv
+hKPAcVhUpczZOoGaVmJwrptMxBBTbrZq5Hr9bX9vFD+aQkqCx+V6OZ9kb8Ocw4P
Ht/aMDTCaUw18bHRFggYtPgq9V1/dj6Kp6FnY4B04QsE7EzYt8oKSgMULgTARFUg
TqlxSGBuxcHOPBxS/ffrbPUA/Lg4GpbBErybVmWM/dNgRaS6XG53N8V3ZCDcmQ0/
Z/T+JjI4JkNJFbkKWSuxcXWQ/XdiM5Jap67G+Qy3kM6bzfSqLC1/RwjKJxwICkAu
+cg1drdnXyogamQ9HmoEluOHzn2Cd6bPMK35gTOB2buD5qk+q1d4vFafmvt6oWey
QICZSW0uQBboZVXElAf8dbjT1Ng36w6HVZqLz+KEwkNszR6xVdxFO2L+QgNvlzQs
RwVjHzduq/8fs5hspSZNzeGirOlsKitkRSYlMhV/IsdjPggnKuHJqv8m85kaR86K
SADT3EbOMWfsnN89qwOukYL5Q3F9ppey/Vx+8jhVVUiHFZqiZfGsWd9OObg0sTp3
bdPv8BUZbxff6JDdbwwcweguBgJ2SsKcERietF+sN3NWLa2YvKgwG5PtW9WZHYuK
Vah3Omdxp1t/WiPqPmLe1FpzjJK+LSYSv6XuE9ynCE2RIDRO8VNzWnLVh1bcU/Py
XYIr7YNwMCn7/n0FR2cJZpu5PXQdfK6EjQ/T86CIPhqm/YPi1PXEcO66qYVSgF5o
J/lbqcm+7W0kn7eLhEzBk8CuDkVB24yDk9mtalC+rGq8TqUG/PAaYT+MYU1OlEoW
kvTBNEXxMnmAxkRj6kv2iePSdZBL9lNbnhr+OA4iGcPihjT7rT7UvlJ3f3bJ1nTP
c3nYfcqzckxUDspcXZ32AwNfViBZ9XE+72K1eExVwwpRytudg1owhagYC0KA16z/
RN+tmDcN7f9TIK7O4cIG0etvkhbTzegJGwJeC58MM7UbE1U3TYYezFaT1yQP3wn2
F4VxhZmMuLYMExLRxTo46PlSGNDiFLLOXCOVSxvFkRWTunLBadeCiFr83SKtjUij
nCVy5V0aXsXpdI0eIFHx7BV33DvUCRqx0ZaZf9utLVECJimUb7Or7K7aiUUeZPCC
biXkk7LQkKW0VQgYvb+9mweZMYlwZEJNTQwrb/sS9rH+kvhBowu2ewAdPYUdbp+B
iMGSDsaE/GtvhO9jFQ9EH81o4wA4p7xDQ4BJNqcMMHBtggaazqWAtN9cG9drAK2L
Kb14hTTqCS2H9Zy8+KgvcbY/zaZDL3gFyGZj14MqWyNJayxkO3I5y7CoNX/GJ7Nt
yA1P0A8DJC6H6kw9zJ2Cd3/nV7xs0Xp410gKaGuhoDAvE85rVygJ2BaxOafO7+Ip
5xivks/wpq8Uk2kTpL05yPtKKIrNfTkU9D0b47B66Fa/2waPWRpLxAdeEDLkD0ba
6iq1ysL+e9XIyZQsoeYUlut2x7sseAnFpe1+Xc8CgH+odIPXdSlHVZFpn4pPXlC7
M12RWtqREDwS5vXx4k/vTDNgveuEyRCLYYa/TLlcz+ax9nMbVKq/DbAPF0uMWUNz
0u25Lw4ehrvggqMJ6CopUkPU3WX5Z/wYL+SJLShFKpQuvjCY8yjjSYMZdiqM0bHX
UWtT61TsY02nY/HdZc/yOo4SFZ6QinS9XZtccSWZuKgFwFg0gxPFYqIR5VowpdHC
IaxxYKz7YcaqlRTwO9zLX8JmJufrooQSEw9qsFQbSNa/YmYtcFUKcGKjKNtoESH1
pcF5tNMgWSoKTbVkBonUpaQoTd8wIMbkL/fBWXEcnrQ09iJzgQgCU4XOPF23eg7t
R7X35VTGgT8GxR7Nuwj8qC/M+HMcTUxIphLcVCvKboIW2WYJekD8uiNWK5DUl3Of
E/xtTF97RDiWd4PLvIVi1WAd2cWOg28fxs8PeCE9GrImG4d9ekYrXlHoA47Ckf/A
RgWn4dpqiE0//p7EuK/4PUMv375BHR3c28KUC85xLSKOh0QnPM1fmjhqivhzmhy7
LmNpHs0iiAdH7Ia+/lVysFz8VYwVkCsjTwC/Xjm2MfWWQsRV7vdEIJRTkA7fLZPC
LBFNi5R9pd1XSa704sj6e11dBq4A4O0mYT5N/msKT3yeSmQVzb03/2Ip4mNPiNpo
6voDfzkiJ20fRcvnW6XLOS4e3HYUdysnK4lAMbnlw2/dtGzj6pc7sPLwcJN8n6nn
HDSadJWXSwu9zsIcIIERLcN9cX+uToHIeHlTXEDhig6LXUWvoKxkFQcS6Q8Ygl8G
aXd2En8A1NrlFmBiEulc3aTvUeG58iEfQdc/AqPeE9Xo58sTrkjmgSzWkS3oDNwz
cqxlV81CB1sh2upqUG+s0A/p0/Qra9SWXCiJlu/SSUyEaSlzd3UmvR/DXGCaFrMO
LfPdzM9kNjSmKf4WzgA27pp9t7sNXdGV7QZuoi4u3h5y720gNxwZ29PRDl/1BDN4
Vm0lsT3nXbLi6DwIRJY8V+5ORgDlTbKdQgLYKGV2eROurMprlO8zc/hNom8nHkO0
ZGczYu4oyL/FiQP3MDgMTxIEvG+EHE9KPcgo2zujuihbTQ629vS2TYpyaVVYZ7O2
ORbjBk4h/Et7YCTiyxNOP7TNdg3uJYLIpoAaXEB3p0o5MaBZQefMF+dgo0YQpLXA
nBFqifs97p6Nyc4KN/Gp41BfCoZBevzi52qgkmJyjlPQI/EcO8bMi35boQyRlh25
vwj/YvXgJtzfoesgIbTvALbYYHOD/TvLQm+mlJrwyXzMN7dypY6mKrhgTAyptUMR
2zRnITAjaV0sATweGt7OqXGAHos0SNDuawE5Cj7sYeLJjOJ+DhihBHr3vRU9ULKd
8SQtbRqJnIGGIToZUOvpejhHLf2wcNVi5cQyrh6OAcelm1Vm9A0X3BvN7lSSiml9
JyW1mK1K459LOKRf8kNuG8sTfRqW8EZmNUKnp9juFAZYDKDhk8RTvXjHzlgOXAxa
Dycs4e/zVD/6h9Hc06qcdrRTD++vhLRzYzqZibwrspo5isTiw8l/Ipa4yjtGiHdX
g5Ul0dgkLE+uNh1dPOHNQIMUijNdyrUoRbJLK0iZCg675BzS8ls7z0rqBxtz7Mnd
9E98g+t2L+SKy8C2lNJaWDLiluI23oXOWzaNFIqRTuCILkENJimihyJ0ZEyVMzUQ
tAdj4jFlNgri8ptwuPzTj9KNL1eDrgY7dfBcBAHXn3tgLbmLYryrqpZ4nVCtFd9K
hoEhQ2Tb8efLmOum/dcry5v/378xlP1bToXpZHeVxbD5ShRmX+hYdwxJ9shxUCGZ
QSUcwZfEr4WX2J2Zpn+o5ezLsYj2lDH61nOQtXfrgs2QxdO+OQZEDEzockWythJZ
trtsCJBzKNSLDJt8X2PxL+7Tfn5ZEd1cNQ7wxYP+EYySv54m5Nqgc/4y30wh2Ddj
WHKqiIm5dnnexQQptiUyUlbDMxQmdjb3a3gkE0OfGw2GRGuthY2H82fKRYaFGtUG
QnMIrGGhKDr296VfjJHcTrNk+4NRfVY6NlOCBqgLBKoDdb1IjOtE+NrIEgaHQrbD
B+ZGPFh2dFjV5qcSBxo7OZKe85pm1sqXUlbPxHepVXvp6HTAmsfOR447vJbF0lRw
SZj5s5pEuvUkfuHjBjK5UjE/xjJmRtZ8GGcea2Jlr9W797+EVr86O9ZJeSF20/C8
R7X1y4DNrkdTeWSlM29lWJg3kcdhbIrGjwkcuyNJuNam+lJD941JeE/De5s04XF5
//kawPyzR9x69QXxsOIkuyRlWI4o1a6vnlXpF8TzoxIK8TFKYrzvng8ForqbSAj3
jZRAuMDwiS6DxStT7JoETtIVVPL0lxqlX1Qw4xAY1BI+/0k9TXGNzONNlVEUOaQ1
kA1XF5ZF+6QJpEdOoEZKoG6axgyCSLkxXSlcpEVZCj5wuwVGpHzai3FFqWfYJDcS
JlRxx1BFbk679rD0ficrTL9toffFRTOIEEYx9yT4wWMT25ynJOxc3oP47dSLFfJU
qbIu6vqnKuYY+cqnhuXI2RBXyq+fkQsysqo2rTzH62c2I0AwCR+PuiVS3ZLXEII+
TmODZ6VltlwujRsTJIBSDKjQf4EcuJytzBdSgHQHB7VQTFcbzQiGUQw2v2NnucAj
1PW50PlhD/7VUMn9/Ct2WctUaHhAmh5BnR7c8E18Lj3HxtgBHFaPr0mkMEpwIT/P
GZrfBcd7sEKIrki1Cq/5I/kgGUYIOHi9pKZm3ME9afbn0A9xSFELdFLRzre0jwLX
38W7uhqsABqoCVH3tw1P5vw/mVY8UoO92Fa85NUrkrF1r2/QIa1j4ntwmls0vPDM
yazwFU6UtLrz2zGhTm4dNQ9DnNk+bN5QtFNwV9XmYziuadzH4lO+UlNgqBKVPO9n
/ojEBQK3PFbuycjTR/qEEVLElz/gTKIBPYBSTyokccJT1UqyBDvlZavaUkYtjCKy
dqel7ZiVsNDefQ4RHZmhCoHB9nfPc9qNiWGhAxaZOSXAhwJGpNSeeCXe6mkHfnU9
XrqxPCjj7YsjMT16n4QG9Q8mjfHTJUkBJpPll/peKSsWh3d3MMeeEHdHXa4s46Kx
Cbd0BJMMfAid3FLwWZdrocKUXLjVf0exBgyrYCP5AoAyp1UivneicBC2oqRAiCL7
aSY798ELJoCSlPGntgiVpdKvqibJOqIIvdSG5wHTSLj6y23cb50zdkVBnOQmzybV
nqPdywBKZN06Gc90iWsbShgZDRuYZbiR6D3unZMAT2rI13mgYNfsBjURo3ToBswI
SMHlNAz8nYvC3+WbshcoTyHKp16CFtKKLHtUt5b5mtrz+ragtmboTyb3V5gciFJ6
qEzGcbNi53dUihibgniPFs+wf7bqoKPoQdkIH7dPsZ35hKGQ8IOr+Xn6w0ivV2to
5x3tMdwJvJYtdncobB+97yZjCRnhBOSupTs67rN0eRzBK5GrViCD70iWiCwoMv2O
oP0UvnutlgxbAbf8d7kDwJzXJu7Auw5IDK01IM1XsigKPL74KxLB+cIzqkE69uTJ
87ZOTsMX9DHuBrDDNZmUETUQ5D5R00U/Saz3HTw0pezueRpUD/ulXfcPcTW1+ma9
wE6fbAbfAEPLQmxik0R21Jss9hfRNguV4RV6oQqDdE/EXiPE7BA94N5TEebOmwt3
hdqJugpKHX59uOwKMnirKaltnpsbxyN9b+jx3X/HR9RV1pzG20Gqiiv4+eiqtQaE
+Xap383i+hIJD3ZBiAB5T/H1Fap5M2jzj2vMAssUNIWb8w+brtRzqccC0Wvpy1vz
P/trB0JRhiLltqVrbEBZc7gDg97fGyMmyp7it231P9MaA1c7AHQQ04iNR+3oc4yW
O3nsvdjbL/cCP1JXjkKkpfmod+GTL4kFODq+BDxfJyQSVokpzBJA8vNm1A7QGSW1
xHcb4On+UeTziluOFJ1CX41sRtfnLVq+geTRok6CYOQYHZoCAZ2XU40PZqimt1uK
yIhYA8W4Dr2/wFuZWrnGqn3l6qsMkw81O73kmKd4ciYhykY5sGWB6vUQmQcUgNNN
dnOGl2TfgPF1nywe6DHPCmH3KzHFM/LEaUUh+dIIrgX52Dc51Sk9TG3Vqa8xg8D+
bZCnhMwOg4Re/d18y60CH2cStmzVdcRxwDdGuI0v6KF4Ia1MvpwzHhg9GOhKJLu+
9GTsEl/nUDHHUos7FzUE/pSA+d2Jo053OQHjMr22+lipoGSVcpWMy6M3xt+SPhk/
s5JA5BjT1RTY5e7pBMKccv5uMX648fN/tnC47NzoGjKDygjimAsoZElzwjdIDZRG
iHwt+INdFvPLXnAbbhnj8UUAvpxqkDSAozEHc/JWoj6g+V77Z+Tn2nAfnLvqDxdh
S2T+urTjyR5F2BzV7QSJdZHLGOlDI/ne4XswVqs+lGCoLqtHWVaSx2iVEYTlMbVz
uN3vn5ulzfQCALBGeCNXeE6ZzuyoVEIWdLbwbRr+AFssistlNG55D72//PhZnfdr
pTaY0VhXfD5pmScfZ8kwStJdep4AJfMaZiMWj7V335lMp72CYt5LLI2iIhYC6pQv
fFG5wqVWa0lUb3MHmZAz0dNShWu7Id6sgQxf56RyQzbXaF9wYbYpIJxZEhLd7LN4
5Z+ejV85tG0FlxmaNZ74saumCubUOFsB4RXenTYKEiJtXuDPssIPmpiSuepQW9BK
6x8PSa6G5JhNoIZH0ycVPMnwaX1n5/T8mYrsco49tpM8NCkdja/oDbe3OWOv+gkl
fVvi+xXcEBuFDMHnVJx9liXA1QZEDIVJQg2ksowjGzj3KnYHS8LCMN7yiBp0atfp
BATu44qRZHAWEjE2pGPMRpTN7SvVSP3NgVe+1ZI4EwJ+s/GRUxO+qgfH6uqES940
gfWszanM1fB7OLKIKlET5qqv/a6fpgi1iJgQrnlXu0gDd67VD1K/Y1F3XcYnsZAM
siUi/dYt7Hf4t5WuNf3uLeGCX9/3ddI9R0M2QAOsmqhukNapg81qpL4t7LmFDF1T
+rzoKwS19/PkdODofSjXzaczGRTfme+5FoJY163sQmQcWYUSFShuu6yfXsSn7hGz
rZ1KAqEzx6VvWnPdVCJcUdcnqH4aloMixh0ZZRxst4zY1M0jnWXaIq0sT0aZv3Cu
VP9hz3ISQlhbb0su4Cmu89ST0yLuQLnY7F6/6aWWBp6Xdxm0tZQSjLUYgoJo9kAQ
nE489YBKBP/6dDiSMM22nXdoQOd9GZzz1b8lcbUws/9BhRQ5tAn4GyA2K/tI+KEv
pAY7hETqnFeS8XoVQBKM9S/O7uTi+QT90dSBfudc6ptw0tigLx6fx1N/CQgkDM98
ogUE9GDCanZDSKr64Tsb8Y7T/wYrFFF6F6+eNfXL+q/wwMdj28iVCJYRWU9KdIcH
DIp0ALZEumi2y5IRBenXOPnpT0vA1shP5MIiC81Ml9iJMIOTSsaMfRfWby+eahxf
PG1mwcRz0fgfOhnl7+/6M+i0kKt2sKUPyVGMNHVzUH7wQUVZU1xUl9Rkmm4LTC1o
52TzMT+xLdLuHJ1gMRe640mvlaZAh6j6HsUpYWoTdtP33O14Qh2Mn0tIYsiuhIl/
NK0cNJsSU176Z//JX9C7kwnvaYB5nwVvxEcF7XE+yLGo45ljgry3TD2wZTmOvWoP
YHmo1x1AWoZmT3ggRgeddlLKX8moXlhEngNXFt0AxArheyt8/XneMiQfNoytScaa
H7YaPzoU+uqH7Veo5o52gmtg4M5L6UrJLHcg8EGJvxcbXlwXLVxSEMyiaQZmw+4U
xoQEw1jMG1f+b/at5KS6cgX1xNZ80I28ydMtTo21CIJTHAxI5xbndhvDzETKXB32
YaoC1Yb55uHMt8M7gpgXYoOnyS0hwIkMsc3GElTyC1da3nCrPpkSjadXr0yj183i
G4wkO39kpwxDRZLJ4e896rW53PqE8uFxAPjua6svGduaJ61UKKac7lUvZ4ngnerD
0KaQRT5HYbrxGvVMnvoJOofVHpSkfMiL8dY02ceT39F3fWEIsMlwsT9AXN6DjNV7
PkvEZVee6ZFD5w3y5hgbUMDop3Xaeccc7afsBlagn+4tATLvYYAJaQjkrRgh0DC6
s/0IIx5AO0PNV5dDwSltJK7aDvM5gaLr7/kkSPv2KFPAIXuuMqLOfx3C1FowVKjq
KwImQwEy0AcYF3jtoJx7zU0gBtMO0Da+6n56tE42tCiWJLmVcDvVk5ycOvrZ/8pC
PkZDI+qQuvlyKKKW2xWb0dl5n2Q5CfhTsoiZtC/v7H3nowRbVcYmUWTcaFcGQ4ds
zaa5SEhLKkJP/hoKk7SAVtPhcQAciY3UnvivHprnwBY/7kB68zxIcAeR4zpbTT6F
x2g1K3pP6l5SzqLEX2o2sVQcUE35EvrH1YkwQSTfJDtwNvaSFKIhIvm4Td54xpET
L8z8ustprkgawtWw6Dnp3KzO3TuLbs6M/hgIojUMykXaFU0eCodeqEePKYKr8ZVD
Fn8Fi3SFtq2BCuKMyc67N0nfmpCG72c5I+CUcNPuMfcra9XOiYpFbkJPG+eSq1yF
WX6oE5pn/a+LZL+t17tNb56QCFg8FTiPtN5rn5+2MAfmMG88bISeslPY+SVK0KDf
6YWR0ONH9ypfuoKvZuPbtGJ7etAbA802lBoWaXFc23KHOrKfRBAJGDi5iEW2j9xy
LMOsAxxld07Lz2uVPsOz0SgygodCnpn8+iQuk/A5IvT88DphvSA0qa4MKw4pP42L
IGM+zQrVe2DJ65Qm5ojbG7sB0ovH4oT5fcIon2ZMfH+0EnunvrsDf+S/y+oIivWX
c07g0Q53s6J6OaSiHF7quKVaMTsK3tWBONeOvPBczrEBD+mpK/9t4CqUG1dc8cYv
uTGptO9ckzzYOM0UyzlOUkqDFy5PSa0OUawFELOvt0IfIoISTDkYwtmb9+8zlzZ3
e0AtyqOYIh9RN5DxHM7xmpPqVLrHx2oUdZeSf8X/gCx/BCGot37mQ9m3m4SAQK9l
82/ZTsE7DXIPCDQP79LDm54vMjoHWESWOnU20sSqO/kUYQNkJ1wjv6cX+RKreKk8
04A3NlUrFN79HDZ9H9eaq7+MUy7p4byBcR0HSASM9S2UmydLqy2EotLNv0YiLrtK
wvKUgnNV+92D3HR5BimtBo/1X8cuDbOpLGgy0mO+mghVvvgq8sGBHxlY5rzQ7Yn+
87qNfvdwfgYKZNOGXocfLXw0biJ2xdtbhOZY1yRCYxqQ69pMpAWzdvZrLy3LiEX0
rS3CT9ReEmcYzt4qFirSqwxh0APZvP6lerbEJE9vwmYpdveSjUqVzBHACSyBeDaf
znc9fwnMDPZCq3+ctTTtm5YaAq66GzX6xyy1VkvWi9ugJ8lTIqX6vsQfYZGN8ZcR
1t00ytbRHxvzt6NRSNcG4rCyl3gDm/ngGHsN0ckvUtAtAMz3HaWV8rNhIYEUXQfc
5o6ptqWd9mR/jxJo6D9MRcviFULznfWvDfznZfg12Q5x6+cE4w7LeEMitHdypuhZ
Wl7WRtKLs7C4kKwYX/28N0zuv53AFq8dlESWlUHvSgElgq6eyWraPrBl9UllS7ms
vJFm6I9+dV6OfW3Wbk9hVGBvTI70coXcmqHkShwsfqvcFUUjl/8GZ1ZmDc09HUlg
/RoMB+Um+CGX00P7GohPnBwKacXortNpalZ56Yakl3MdOiRx9bsat7wC8CmgwXIq
ISzfEtgflxfTY6DdKDMoiw8oxdCcbMBoaZuv5fGZg7dqzF30UMmEiJf1mfLL+/oI
hPqYoMtJgx9rX9GI8EvK9e6CmpdPVaPbH7mVCRjV/SYdgQF9+wcXMTbsrlUgpZrE
jQaajOavuVWX3Dj5NmVHMmBudFkY5mdJo+oAR+arohZeyiQalLGkIiksMMo/f+zM
AXgZUqxSUT1z+8J4izUgEProTMgxxZuODDjg0Cez+noYV16o3t896mDuzBXMRU9/
OXSN6J47ILAz4m1vlcJAYHeW1cKW3iP7/gObR+gPRMKJOFZX6zsFostJiXGXbnKr
iFYxYolJ0JtllSEA/zkIjwpTk2acXoJUwoNO5S2uw0s5zQC1QM7WwdqDortB8lCL
eui8Zbc50hmzv8D8kklTndoJdPJVrkuLugXwBoI/SwXr3MJ0sXeBKsKupBdJGUTC
xqAsPiv8JcrwVfU0O16QpTJZ9AHu6CppQ3R+0gkrvqLUxEqY+RoU6GLT5p76rhCt
+qnevD51cB4D2t/ITg7L+Ba/CkwrbyKZYT6r/Yuelg+wP6rWnVCPH3UN6u4z6EkV
ShKf/elK9UNconF8l0YNoJZqtqAHOZo2zp1RhdiQhu9yS3TAPAqeY0AxhlVYgRpZ
Hotkk/SKHgxxiTm4O8wSIBcjr/n+jFqVNhrbSAPQ2Itdf8Cjg4ba2sZVEsDkNvB8
t/nvRr0DAVHX+KDOXJId/1zeMSTlRCMSHQRnQjUoXVZXcHHB7m5G4JJFYsEUVBhJ
eFODDlnYcBHNsYNGp4LJaZdS3mS1s1v0CRFNAjFRxmfrk9uykYGD85SNTTM7OrKa
9SgDuyIBWTvYIDS4sWBJ+BwFMhX0+wcVGeZ5LMvVEuwf141a+efGwrT5QJEQ7Clh
ld1aVdcP2yWyOQP1Lw7m2p3tjeYxXwlfSs7HlVVYW72L9GC1MhfreQ1fhME+5vwK
G1aoDyESevXYq4mJ8GRsMwq6XPcA7CKc8zzrQawjogNvZTNUWPStVSSV1v1NX00V
b4Fe0uwksb9AQDHYxyQ6ClY9tR6QwphRYWmfH69SsMm9wuHbBm8CW0B4zsmRxKVA
4ZjOWwJyTd5s7+fzAcRDNtSkM7EvYST8A3kVyewsSit1Vb4OPeDwvaeZ/ra3VTSt
4rcl1Yk325jEgFb7a/wI1Cj4uSyw80BjUp21na2sJOiH8EXqp1kuiLrS3Sxqr4PK
3KyXmr0haqsmMCm/yJWlCGEGE1bk2lR5cxvD1gX0LkiNvpXdoFJGlna/MhQCyz2D
2U5bZNsqRSD73yg+9tLmYUktLlV+tb70sgVaZPVcz62m+oV/r+gxEg9e0r7UJ1wb
5r6+fEqG6X3GxH+4Altmyqot7LjycfZn6VRXtVLbejVx4HGf8NePZLzLdo7EghdQ
cEuRdccRTBo/9SLOUmsR6anzI6UTHtakXlj2BYfSwLrmttVtcQj4Yv+LTaBvbsie
ZSu05PxUX0Q4l57Myo+0Ww5pHiIgXoD9RIX0vTtawqf+0ssJqcMjNvDZaSSsrP4x
ZgV2o1tJagqG2Vqdj3ZXVMY2L6jDH94av6xhSnPziXkR88imrI5jiCR6Jt7yD297
3BJuI3zQX/C7bBiqf+ENhveOY3puNzvhyedtyQM+nMNQUrU418GZR7BJotpUowr/
M6XF8YjlOFpQA//FK8qWaVNMX5RHXIesMiusxdDL6Ms2QD1bBs1kahvDTa1OJ3nC
TlIh13HzaV5LBmnNHAVLiZmGf/wTZhQTIEcaa9Fj6p2I1yOiyzy0fXhnqzscFOyK
XcW+EJRF32CKNMSq0WbQZiujCy9l3MVE0+KQy+BWoe7gxlHmXbbB8KvzzeopypJ1
d7XckggQwwPv5brOy1g4qW1BciS2ZVP/Uuc5jgRtkJJMPSQlJQkydDa7J/eRD4Jl
w3Yp/zcpTdxlCkXBAmhC0U18NShhucuZuvYJB7siV0FFrvxjy8E1vFp4gL2sgyTR
6SBBcvxyEfMaiJqqRjJvrZjIE1eivyg3LIt/OFXFQoiTcQbsRHSEX3SMpFj7wQiB
/UqsZODqB75gClyONdHnIyQ0+Mye8T8OVkd5PtSSvlr33xyZ6JKKZ4QRbPJWdVZ0
69KyOAZjmjnYwyHHGGA6rqOeOL2xC9BUJaQJYOFf5JKKx3u8cdm8HTsSPB+rS6xy
dLBN4SeDdCZH+h1pAnQKy+R3TECJk3K/vfg0qXr9rReyC55lZrwvMW433FyOBOHN
V9MWa8NGsa4Dz6/hIziRi8C+rEVPQTzy7j1nQoqlMeZpnk/JsAumGv/UakgjA6yn
XGYOGMt9OF6rUQaHy/xq+LeooSm57sBa8Sm8IK7KFwql/vjL3J3+xnBx6JpHdNon
oWO9WzKVUExRfPMizUk4JZGA4hz19W8iOnleTx/ykLGTv38gueLEJNJWJ51tXPsr
R4YgEJTo0FG0NNEHtuemAQnVOWvFdIM2IXNMKt5JsRkR2kij7+XWFwTACB8ARIQB
rgRty0/MIuoqis4QStT7/lU/l0eetDdAWBdMEtGoicC53BYTiVTYlC9BvbNIDNLu
PYPGtWVzoZFZ+0DKf2Aov6IqIOd1A5U8lLWy++9ixsK1Gh5hqCrgycz9gbHi+s45
XRmdUeUR4kxdaXsu6cxQbJPY+MBuxXOrVLjvL+pP4QLpjJkmB1KzSrhl3/w4uyzM
M4X/g9iViHu7trLq6AVAra3kahrLfwDZKEO5okfTosw/s2/6yStGfosEMyZspqzD
WqT2qUeMLcrDYYUMG/BgMUHFiv/TE7MwamjSJDffJ5k47seGbRUMSxUc8jrEpcu3
gXqv/tMhsOqI/uuyM9u6beiihP3ZDl3AqmQxUl+I2iPQf29WAR2N+yD6kBW5bDUe
tUcFKGq8PdbJ3H9W/hMNkJEkSybHpLvJEvxsDI402+bYWZuRy+AOB/gmjGm+2ztT
bOx3f+zCqvVIE6C1I5sH9KOQM2u9rOkkGqxNtMFrP91zsHD3E+DIpDn922isnBlx
b2Ye6f+mBCmQzUy89CfvBGZXtBomRhFldOjURGvdinb4OnAJvwjyCWIgBnY1F/7G
DiwjxAKvLmmMKyQRcrKh5kTd1ZM0DO7CrWwRFFTsCocImQFaqRvIB3CUYJqOppQm
Amb3LHS9rC3cvCRxgnkisS/gTduHHVuGf8wDSyaTXTT62yUfuU4/QhBPwVcXoEX1
vMCNPjSQRJC9KMM+DeHLOxr3B95fp4T+OFWS0vzCSpr9dIcrGHyjis2PNBdUbdH/
ZLqHyHVQoh0gKI6rWlt6JW/Dk6ihGR7oej8r5Tt0C7KU7v6QJTQSA3aBYxQrg/Qv
W/YGCIj6GtiOirJdeGFsSelOLBrNrnBp/VfiOrffbckWnOdI2Ks0k5t6WxcoUwrF
3pUmm1AUKMc8aZqXX41f+hTGGg6t7J04HE6nrzfRCCTmttdyyUVD7cylrLJ5R8TO
vXAOH9ZNNU5e5gDfyBRgiiIhu/nvKxsBaQ8SFNKYazwsNRnjh5/GlKNKpf/3FtoP
dllDQ23I6+gHMzvvvP659qIDqfdeWQ+QsLRHqtuoL8PXC4svxhX3dQb7udB/Wq5a
uC/CIWc8GJDPMBMn2XB2BmUQiB3jRH/45G/gFgBKnozHu8awoWCx5Et0Wnfg6rIu
f3kqfh7iWHCUGbPmeN4Nx+mukWSKEU/dLQhGVLoVyfSulYz86kXjtauTdMPjNgee
g2/cB0RMLfJV2sLjTEL0539YDfzOok84TEOJEJ0tqNPe+b7QpTCmZPr/rUGMli7g
nG5SJcJ8aHLCwW7xu/jv1K9MdvLKc0PXHAe2gdQff+OA68M11rYEwBAb7dgeb3rV
EskLOKi1shVPy6UIaBdwzs7u1Ss+JIdZzxbc0l+VJR91mvToVaBVp0BWb1Z5jdlV
Wp0Jj7G3t4EMNS23O8mMsrhGZ4AUWoXuH6mbN1XAL1uD1zjy8dUE+k4O7Je6i6Lf
ZBaG97xIsFpkLV9o8RUTxUOSJ0qZLgPxW+7LmJ+wMs9Nl3NB9J2Q4aS1vUwDXUf/
RQpF+1EUUAk1Y+RF6VrBQeR+CjD49Fm3wuZ6NakGiWvr13L99qTNkbS05CqjYCcG
uY3LShQ1NjIaZaJwdT9LTaKnPzIIqKRtPlXkA2LSEEDlO3p0qMTySN5W+uYoTOlb
I7KhP93kdKgt1HFUXibLXSvb33RnMj7FdPUZIsHZaZXKYAU6evzFnhDcbRjQK8+W
TVZHzK6XklMFL2pYGyeXvOcGa5y3ZVBr6SjgP7w5jULVB03FcjxEd9XsqOgRrCsB
gFB2Pd5D2Z5nK41+ATC5qM+yn/sijQClFYSiJUPz8X6kV7KtoQyjofunH0+/J1Aa
UAQoYne+bTaAspWTiSF3QeBONsloLg0SGJktt4zE+31PZON9m5QWKD436LPOI1Ad
UH0k3XA2H5+4LN4+M+unVS0mqTVz/4ixSH0GFLim4ChJK4WL1sYg2jezjYkVpS4n
vfIvkNlfbG/rxWZ/KW/qqEDNQ7l1J2ygHMis4PGIH+YRhFFl2k9mrV1g+jRJcGNi
37Klm3euamx3UfJvCpa3/FzYV8Z0Mgp9L0NzQV6VXHweGpxybWMr2tiFQT4+p9oK
sNniFw1YaTEffbrhNj6EtNr9vjH9t1f5MFb3GR3v1mz1XOj4iwAv5DZT22EbSWjZ
yRJvLPJs0apRRlG0q5LawNJNA+3cGeqhmbB0OJpZJmZxI9ZfYNPtWIxVJRYCS309
h0Huf3tFmRF++Xqjjs4r1dvvEHGQiq0EcSaDKwn1ivX9YyzV+/eZB75eP380/KOY
WG+FHYELjBr8Bt1fQXPvYDitDdFlBJ4lovrtsSItavteKFTvIldAJTho4DQg7qH2
z+a+Igk7lsEfEX1swws09aurnOg6LUxZFRi2Z3ySAsRtpt/Hqevo4QjGO3G6/zvC
2tRXIkYxPxRU5FoimOMPkHxZvTgfLDB1XlDmWg1FcxuoLTEXthTJyE+DYNHMlJ1r
gU0xTAEhltU+XY4PsY1Ll9mIDQ+uGVODHhRLWWKOZiBn6GSkPFgrxeHDF9sHcOkK
nEMHX+CzJ+JqNVFkSeL5e56J8yIH4FJ+hk1C6oihc2WLvFhZSI+9LBo2S0LKB3zo
WHAeBZIiUZvideDnAJdoJx0Po35igpAb2cTV0LeoZG193pKjLp7hw43+ZsUGly0q
SusfoUcZImcmKxzekmeNLVtOeWdLpRmLzFic4gVv4udZLLEEdDSv9UoTjaEwNVWx
OxiqyPLCuDQS2GkKT6Hz0DLrJg+PH+nPDZbv0gI6TLVCO6Gzo0rY0Eq56hYZ7Rgg
3zcGFm85/o78Yb2BgLYFdGfphP64d6MOHAX5W5O+wH+OBtozy6OkXt0Q/dl2FWQZ
0hbWCsaB+Ee26WjTZ55UKQTT9+XsqZW/4/gc5yHA981YGxLl9QdxRJ1hwcpwc0DI
1JXZOoz6Drf7XU0UAZO4uVqH+F2SGGkQpRpWvTo9p19FQUjsDKUoLqckK5HsaFlb
yVIzi9QIwP+FSooZhSFkf/AILQ71Q53LqKluZFCflW+V+AOjfjkPUQ5vhjIRrGJf
jrL/RPm8FKGMiQi3esL9JarkkqPcEpiQPBf/W+0mu3zGY2Ow0aJwIeYVa+ryGBV4
Ovoh+v9ktZBrJJAHmdOeMkFt6ZWGUkXsjvDjd8Kt95Z0yoq1LEcp4bqd0C2x2KmT
9zXIK77KHAZUYuRIzFUGPe6W4kj1gcjFmBA1gbj8A2sohqKKHkiJQT4eTttohPbs
POBuEyeebhgZYlpDThMLXB0oSEUEvQFGGogAHBSJoiVhSiPvAT7EpaDJA9B2a94w
flcxtfXyXS+nAXOelX0x9rSPjYm15VPdsjK1hkweCS9fCO2Ocfkn0hLlC0e3JMr8
kPc0OSX1kVjpgp9ZvaFoPclZvNVJUqIloHQ+PTZwHSSUfjhfWtfK2Ma9GPIQpzLB
cnN4A9LNa4b+uIxZAGzeso73fXbLlcQkxhSVdLWKOkPZDu2vapbytvMUR9RI2XmO
Z9N29uS0JD1a0P7jrPB7X76HdOEBWknBrbCI3GXichP/wA08se5te5B+TFMBU5JQ
PswdEo8RLuOoqOF86YYwe36ea2ZO5m3rWccLLXFySiDimdbsc0AQzcpI7t0JBCz8
S/GRl+UefLZi8UFBaxAl06XhCRQt6Il1Z3O9uZsjfPNSm7LdgLfc174ARoQfV0vO
5hVWxBdnOWO3YN/GfYeetGBx2r1OEaUl2b8LJsax+fx8rYHdudXLZVwdIFAXKrey
eLX0UBwpWtndhhIqy8Hle/VYNrFIf2NKJVWVgIcy1nOlDV2hx7Dc9Q3FTz9b/w/u
ebsNxeZT4AZTC+TcvdPLM7ZgL+c78auzbWDMTYf5uE5b/z9MtbGWBKyJtUiYKDbl
/C33L71U0mp2bt3Pla0vDGADtVxBmcKsI8XWrkEmc5JBDJhQk4ttlkEa/VGEFQNj
l2pTiK27diOoSveahR3cOuvUghOiS53pr9e6hUAVKv+xWc5CyNNlwJnkbdK9/JEv
gZZ447BGdeG1DjLg1gCCw4K6F0SwMoM8BzL1UPkX3EJCi5SLzQWaM0Y2yZ7a6GqA
0NxQxewBAjkdyTvmB5WaOY2MzXJt9Umat6tMlldMiFWSsgi4pJ9TctzBGU9cfDZ/
Rorbsrile90njqqyKWcoFlTz3jMQaQLS2s/6b6h6fsaS9kHvEj9UtJ5LSSr6sUTL
V0sc7guN+VaJcUTT8leQyNX7LlfaK5iEw2jhTe8fR8i5nAVizCKfZyoIy0eM544e
4cGkNVi4JR+NGM5K/svwqpx0zKzMCy1lK1qbxsBtZnfRM8YICYNs30pn353EyObl
JOPRhSj22VBKfZBw1FVEg+v2XTWXxIyD3lK1qsmkqIYEcUTvnbs5b15y1k79kW24
UZGdWyHOvSEk2AoyvR7zUBLGKeQ36R/At/zMvieTrlpgp2lOhugI8U+ux3vUwhsu
/DYBFvO2bka9/ss08YdB135EfBzg6LdheUtx+BzOoiHu1P9HscZo0uGNCGrk6ZRq
fhDoGCdwP12Gbx7BADEKGDP7hZYI5p5tnVmUazeqUvdtksoYRKt5eWNJRZC7J5vU
ruhMIHdxZYwp9DHLWFCrBVTLgyiqqh8S3k4C7ml/RRToCIaf/1ndNzVX1qBSDSak
8gbn6ybCZJqExMm7gcgj3i6aCFHmv9lctSs9uYdyuIZCxtzWUMR5ZfhhgY24NWWO
sZEy4Oq8FaM2qHO4kHgXkSQapE54lHKMd4aiiiczAkGQEOU6ijGT0OxRci2FYt12
F0d1pImTdCS9wmX26N+cz0GHkoZe+UASwasbYWnlxwmaLAXyOOuQkQWMp8e0Y38X
gmysKhTgaCVYvWb4XXe9Nq+e8AbGHAMIh5b+k4i4TXNwxUgqwgG6FS4icyWaFWUw
RBEP+dq7jzA3YfN1pbMVqEE/vQV3JRQnjR2LswZ3grQRM+VMci5OVeFBNWMms2/P
W9EXRHRByvyPpRNiL7fujxwv3FhhuaEvILOjx7MSwIz4IC0w0vStTHvht0xU7843
Dc1LZO3u6NYoh+4mGhohHZwEo30JUNbEwwg00U/8NeY03/fl44T8rVc3BVtsuYyc
lqRFZbr47NItDfbEviHMlzwRxH6mcCaNjGZe+YnO35Ic81v/g/E78BuBx35E+HUK
gQ7Ar3GJ9sX3Eh8hneSVpjfNbtOdz8y5VsYOw8CpYfunC6MMFEFy2m4XmUPLn6YN
VQ7F1NJ/0XNwTRZANZwZ6N//WJaOB/bgkqoHGFGkG61ufcpudeaT5MNZLAfnO70a
JKW48hjckWHIRKUpcYuKeYWHQ2jg1eHsEclkbnSwSk/kclXTKc/VFUXitE6bnMBK
ExdYxZu3VXMVPhARxTeoCXgek78kbTHFVsVTpfb5LMek/LjVXTtQUFCxhRE7KfP2
K++SxDRcMeCAi3SvK/Edr8XGrGAmhcCGFSKhKSCxMtx5Svf4vaQoaFq8NAJQn2mx
8l/vW0AuN1PlfsaqVCmnt9M3fZFWdX3bcQqGqT4tW4+zKLSJAwWRppKlonuOspWf
0HUCzIh448kez8s4uea1ktrkdXg0Zq11qFyr5Qhd5J4pL2hj2d7ffCGRUNrGVu21
MTihM+zoScFkuwLADvj+/zKcVT7QfDgDv3OYC4bk49S5vkVXRLRAs/frtaoqleqB
W38eNCj+AkDsphzoPsdZ1NLPw9WcPK3WJ7pV5LTr78Gm5bkHcncE/RQ36co0sJHg
3bNh9IXcETx2/fc1BeKdlGT/01dzsZbeQJelVGmn92XY3GQ39DOSZu1qsEEIVSQm
R2kiSXaOyyhHvxZ/7J3+P8UPLFdC7/eMXcOuLZnmPCuXgtlxN179Yva3k0kAQnIb
ERoawbs3cdjBJE2Zm1Bg6e9pjYvchRCr2MkjPGGLsn5fCkkqLy7fzTxhYVQgOiC+
QEL9gWuENNG+W8XOTnJ5Gxy+4UAroYMpVYltumAR2IGALRkkEfzzvgSPcVAj8ZRt
2I1+1O+foIPkPGERutNRbJtUOlr38SH6PZSaVANrIvdZbFxI2kp0EFo1z36gd3D5
8l36OHuVkQ8oh471EzSVPwI9WSQS5JwpLXVO4KR/lInOBZSBmyvZU5VfWrMnvT1e
XwfRQfTNRiyRYbGsvXb0oUaalnUC5J0NDLgPpW5+QbqMGl1Qm6NRgkLoXsKgGBfX
08CMLn18cBdtV48vKGf/sZQGSPERWuD6DrGLX1wd/1MDS5WiQ/5dXLg+l0uHB/UV
swzriaWobqZzJ2LGZC48HvmXoV2CM5VY5YS9W6AsptmGIdMZ44vR0eVDRPE+bCKm
drQg9dEGa2cuw87gWtXv3LLQEKTBFDt4uDv9ylX8bydYpq7BAUu6dPuF6bivw8kK
N+Q5Wbj9PYLYSkYixh9v3Y7V3s7K3/ENB9JWpTmZHWuqSVhWcNhrEsgWymKVUWsn
7NH1G0S3bZQoDVKunWc/LsL3RE1PRWBrVFEaiPXBVsBNMvjoS3fIwCj4JqyM/Snr
a+JluEEUBIcmYYXEiLunoxhDILCy0Fg54rvxR5Gn0DL425v3srneR+VAzqsbTBQQ
Yhc+Nkac/gX5O96HlQeyMcRchjrdIa6/xKwzdEJsDrFBj6mmbX7Y4yM/+zFMOKbn
lnl8f0cQTc4eRiTxhuXCcMZoq0g4qNJyN18AAX5PzQxFkwfjpbGQvsHV9BnzE4z5
QAMnxJfj/z8KzZe5zQt/icE5P1yR7XHBePAp0R/xgsYzgJcN5FwkT65LPUn7cs7l
h/7m8vVi8bT+78nSpQ7R/OJ6p1HQnIrMKqNXoJZRl1TLB9GiZ/RdZTYk+1qYGREV
/a4lmNYw7H/7bkUJF1X4w+AprlYcTTq0S7yrYIOeGqAHwpxlFhv+yfaffbk7lGl4
B1TcRK8zbfHrhBSRd64pmOdJ6GX3qMd4qzghb+i62RSfdt7RMr3JyVnba4tSWe2/
u0bIBJYJJgCsKf/rSezvOTkFvgvex1QrmLOLhQY289BUPrcBvczNEbK67Gk+aKnT
6wxyMbz491saYcBS7DyNAgDpR3FWkS5Yjziy4ExaPgueidCaT4EvWhx1hCVx5don
1SqHVnHzseu3hnxU6A2tRefj0GsbzjA9sQteKW2rZ5pWI7zfZlqBFMY/GhbMPRjU
V9qVM6pPJcS85WAmeNig+NaTaP4OIbq/ukRYvDh9h2H44o9lgU9V2KrMz25qalSD
7gm6AsxudkqckyPcotgBhvPphd49ZtyIxklK6QBjvOy96tuIB3/R+VmxLf34yyvW
assIEvfyaCA04gmXaMtGfWHoJCtyY6qBUXtUI7ERW7dlZgHorvF4KJjaQzMAL3cK
I9ypS2mYb6aJWKsEaTUbTOvZLiirVTBM5h7OKesBWAnX59b0KlqzBJe2pHGoodmL
H8Aaa/4s7MRBzSsugB/pETJ4yHnMLbFBz9Kx4YA+WSipsjVcbEUeZX+vpMxFaD2q
1iL9vxcVNdidenVFt4pxgfv9L+NMDZV43PsDTlaLz5JdM2ewTWM5L11aH9hMtQXS
o/WBetwqTc4u/2Z+OObinSL0Fw3YPVn5veCI3bFfdHGBwgGnjb7si83ZRA2VgDkL
W7KQrA8lYkQInYMZUAPN5XbQTG6zsqXI5mUIQLYKCfkwS6lJyhaXraDbpMaOJw0r
wSMYZU+ml6avIBc8uU6HQ/7H5x2GiACWkj27qsAkhAElgQNk1Dhv5EEpQOXX84b5
MqTSmaJ0GphGm4n7G4gwZxlR9YxHPjwc/vbXr6K9BQhiQOEsTHMc8TUMVxf5VWz6
tQ5ehTsgls96lvDQ38lgoeBAUMsuTGmnMK2zTj+UmbwVqNHds5gSpCeuR4T7iuGH
2OmpfNqfdVg0Y72UsiA3Noxgzwi2LwFkwOzvpWyc7pp6uBb11xlFfTWFj5ahJKkC
0nh/A4M6hoK/NhWtZrg57DYHElwE9BMxIjt8Lw+s84N/D8BTNUQUqavcwiHMYUJq
M6UqJPspBVnyBdza2CWmgHUJLbYCYq1npKwi79cyQ1GaG/WtNgUh8CGVBC5Sdg8D
2Fa6PGkl9SCUfUkuwgs9ChnB6NVLB3sP94xsZuByICujktn/sIoTyTMnSJ8irn4Q
+xvX6Dh27U3fGDqNGYSFM00F4ctLC2mT9SN8y9bxq9+nzH3RyChctov13OZ2jrkW
4yRW3yrf7M2oxNtra1opk9uN0zDChnw4GdPAztpOoQ3Z6u/t2GUPL55oBWRUivPW
lqAy3cEWoeN5XwEDc6XEfGYXSjniMqq4R16IZIw0TKyNEZEuEXvwPJy2f1BVYqXP
CODTGYX3mmjqjaiKq7YEBdpqJocdm/qESu/tGWJVzFFF7sR/uRh7UGQRPwuyw3z+
ic7n5188bQ2xfLKlbwxU5BAhyhxDDlCC0E37O2P3dLaCD/y/IA0HJXMdRWwVvjlW
cPlkhocCvB0s0vTKsChWdeEpTR64QmQ0JzB+MivzRQ+GmgmCKf9TctoKnh3R8Kh8
T8ljc4TBC5sbU7wVeIQhPfowTLGPMJ2XUCb9kDI3aSIhjxUMT3NgFuUbt4gw9WFE
5JEUqRt20VnWmHydxe37Fse+bD483+BAymRd/i/SF03KO9Jo7Uja+I9052tq9r4Y
h+57sFWdqJ4vi4/CXTLx03KmFBo17dpPnb6EafvNydDgq95NnnvyuynB20O1/ox6
+hhIhPg/7xFtk7C2jrT7D2mUU9/aCKccZiHmWan3eqiL1Ey+yHrJATi4PdABS92W
B5OHe6JDOv9xNVqLgMlWNRjlJQ6prruxSio3MNorfBHyK88socEnGfak72rGG0Zd
2gbjIEzpDHNNaY7OWOdLHPDZu5BscTOTpyODyAdkpt63yEWqpdNurRmUO25cQz5c
eYFmG1ZlEDV4ecS3uFkV2JOFHsLvps+0etbR9jFJG/7mR/Yejqfoq1xiRDbgq7aA
0BQ+WxtkQUPLWz8Xp7UB+NPruhNG0PVl7Y8pYGGxjHE3Qv0CagxII+H9Pyqfr9Cb
rppRK0H86QCYaTX8HZohFkydRwoJZE8PmLULkcLQ1/vx7Y5oQ6jf9+NqA/FfB0bK
NmnVnT0qkloJON1Zvq5vV9dTzw6+BUMjrPqtSsp5maXjl5U5lH+0S3czU9FyxA6f
jBw/Td2AadvSwiQvQPUg6NWAXr2fVdkbPxXGZiYE98QceUGowdcgIcxkPCl0fUY2
Q47kcJzDQbwYti8AMFEuw53GKe8IRQRpqMgZjTTIwV4GvVoDbG3vfyk41AdNbjuf
SZV6iYIR7HEjTD+ioUG8JPGDQDHXlY2kJtWMp9MdUWlh0DT8a9CCqFQ0VR/6qSyk
4t7EU8jsoqHkFakMORLjkp2aWG2dtDKnwQzT3zJbhfwSwZ2SSqpcaKKmMS20bypn
qL4Jt6i9TvZ3JF03gXa6NPPoKxo+Xn7sh6cA149lFWxuZkFc++pzyEZeiLAtWuUz
4GPR/wN3c5y7989oNF6EbpAlrgpRwmp2UcawTG6FWNKz34w4vdiDP9n0+HIoSNec
pSnnEQhH6NL2i0Qhwu+uRKa+MIDDPXKLADNSVe/+uVyDlkkFykT5j9BABuZChffz
IurO5ZEomF/ssftb9pvuX2Qy89wwIpEZua5AAn9Pzb8d+/TIS8TVp7nv3L8Buvna
gWKCOemFFEUnj+CVUKVqvBoJRROqjrMvg+l3oc2F4JpPtPaycvwF2hW2Gis6umA3
j1WtRu+vBzQ1h/ttPR0RQWPVu8y5nBMU9tFei2vVRZL1qFWPPFVHsbCcbW5HbLWn
HEaYlQCADe35Ls9XoUB/PiCgWZBXPSnWWzvDNMQJk1Cz6VM4liUJW73vaW1tmbAQ
QNIA7tz8ML3OHdH7eR6xuRtgyf37ZQlPy1tAsBGCyHwXWWK8pZPfb4LGKv+kI622
ztNR9oDkhVLaeSlvz3KLfyY0n/6ROhlA937ec8QM4H+xyKmkRJMhKxScI0e5fD/U
3rF0MOqFeTxYsQyXY5+HGIs7Y9E1AV1f85PCxPhOjgwBe7tr0K8jHeSq3WLipjkT
r//SSz8CYXXmFznMgBfU5b7kEOhBCy3tlSZD+U5w5YtPavfSNE4S+xaIZmWN0O/v
4FBZ8+jIDfz/xopji0VQ84WtZyZ+nwtb5hloUsQaBMtHjJjQCCsw7Lll8X76tnbw
3MOzIKoJGQbSD2kJ2n7DjapVN9Iz5GyZRyBIrW1MIhuI71NGIKB+OQyymcEvZKbO
Fmf/d4u429t68dkebinoYmpK8QrOAX13SxqUez30PQGNhAq443M7cMPJ/LlphPJg
D1tCcOAkXDg2LfS89ZFmTa7fl/IXi8jNCh5tQIlMIDEGWQvckCye8hu5bg90pw9H
SuJY9dD7dSJiFZeDSqbQ5iSVaYgBI9IFnn0m2qHDt1/NXPomrSSx6fw1Fp+sFd0k
rtUrTGkMUxVPE5jxorPYJFMxYakFjgAw5KNDdDfunH9035lL/fnjbVxnGflKY/Xp
e6dMdseTUWoTUtibVcEu+O0U7JzhfsM3nzLKD4q72+CZAH6CwzSKDS14vnPfTM8d
vKJxgEqVCkHXq0QgIG9f+Y/+fUCVEAJJ78yoqYrzWqha+DVSFAr9wZa8HiRWstgC
EJan3+FI6eqsUoDsxVVrCl9nsUYW6ioALpZi27j6aH5r967O/Mx48V7dMy/hqxoT
tPrd2yd5bIddqthIPF/qxXQVOnQZXZYqj3BOPQAqp77ivMUSDEGtr5o30CGgO+Iu
Y7lYdY5qu9eRS+qJi9d8hhUyGmd/c9EGcvu3F65aguepwu9N9CGyBcl//Jx631nd
RdEBH57qRta6lwLnG3saVnzt5RIC0DJ5WhRtCVCTdA2vq1bvCvjjys5ral/F2B/M
tBKo/M3AGEov79PpfTYlfsYQ7IGrCf5Em/bFNnwmNrLXvSTW1onGIye3+cO2+Bqe
InEZqiKQUc9utGKsNcwRwH2ludmCw1O3wAmyTeDjH6aoBMyK9gUdoX4WKg2Hkduz
HvfhlgH4aumqDE1wVqH9Ab+m85v8hoDuIsyeaCnOJYWoYlkyGzsxDLmdQtrLX4Sb
2HNWQTZrRt54XsNlkqGwiQ44rVz21vX/x/u+vHKqJJxgIhZamgXD8TWrWofCJJ1s
P/LMmySQ8S0wwxyM9tCGud5mnGD+4Sn/dz1WCpJwYc62zdlwYtxuruwxxrxns4E9
P42LX90+2Wv0dQat1WJHZU4G8b8PIyeOSCyDlPfao5TYw6dEjeLtJ9Q+/4jnsY/u
bAfWPhuW87j7yqYMmM1NTJJeteZ6u29upbeWlbyN/ymN+rf4Wd10sr0VHkT/Njt8
nnCBMuR9oPAZNLhzrpS52dzsNFTuxHEwQ0uZU3ivo8QnYaI6UGzAh9FLl9lc1Ztv
S/eOMk6QTbX6TxVK6WfUQ5auvq14jeZoOqAHBUcJOs4RpZuGs4FkPY7L/kq1hOV1
9LGOoP33tu2z3E9oaIGo1Tx9Yvf0nh8NNgePq9/zXDxpicnbumHKacosnSTL5wEI
IJLmMv1fy26LxuyrnT4xeqD6yY315TgyOjtEMMNCeTQnffxc43woVDETVVuJgm8p
FLcHE03Kisiy67rzPiY/rSPrWlGzlWFmwykM+z4RN9I0JcQ2tfctR86U89bz0Eb+
sC4dix2c6mC+2Xt3G16M2IwSZk0QQfF1F95onsHRXo8/C3GjNSppxt/BIS90GjNh
dm0gt+MrAqfkWnMibHYYa1uNYv1HMd5bmbdsCKGs2sCPTo62kC390z+lrwV4oVcL
Nr4zsHrqQ6XltfuSSjz5F9H18JUeztGLsNJd1oiq+1+Kzvj15nWSbt6Js1wnNBNc
+HKBgnjFkOqqZgw5ITjDBufYVneqU/3rDcO/bpepRPSDst4EUFaT3b3KIPgYVSVO
OMgYmXzI5L2deZhUKvNEjWgXZ0ZwoeQ5TOl3L4Cz9OeneBLvulDwk1SVX9iLAa6j
kqj20d2xz0M4utkRl/AF/A5j0DZcJmTrZQs91RObWc2nvcm81DVRmXsrKlU7JUg+
5wGLps4V4RDR2KCv77hTWd5bxG1dWpHWCJkuttfPAE/YRBXyesQo5a06ZNmgbbEw
t2fFQyabejTjyrqBZ3Ja/W6c1U03mjiCDpOKWQacCG68xV06Ox3XTFDgmHRsDPmV
6K9Fg7bPNZze/1pwQc+otuMl2gSuFJcVAXAECnwYtqtOZDkK/ladI8a3sK3WJ3sv
iGWl7cV4t0h2UCRE2vfmuZ9ORkDzlBnjZ14jArgRb+uAk7F9/4VhCU1Exz6Uz9FY
uliQgjazBcGWtX/6dx9RagArEeK6ukMoYL+8gt7C5pMMdTx0vP1DBDUVDJbM1a+M
egNSRhF0r0cng3302y6xcN042g4uB/V4l1beRzGcVLE7IKQc+4SKSrKQprl4A5RA
kbsJDRAerXS8YzXnhJjFGMdDlA3PmSWQDhfojGuzeK5iKJyGiFN7ldRVuIw1DB6h
2w7lUA9zB3GanlTzJm44WgsQ6XWUFvEYPr6RFCMCuNbM6dx1oV25fqF8QOBzflD3
iipN7othZRkVLhthH6PlbrfKwiAFZz6GiBQrFjPM+IxNBAdCI/6lWpaL8f0XdzF9
01viFhEz6vr0kGJ6s5O3qXNqMO48JDo1Dy9HmsdRrVTr3DsQzGPuRQ2/6st3etEM
yvCkjFgifA2CoRkkgKcWqaEZ8TeXr2rV2LBaGlSAbUZvfwG2OBeXtELJaPunYK7O
mV++33bT1FdLbRo2YtXQl7N9hCCR0thvp9S2JHmv1AmcpK5EM9gtCqC3gLDpm44w
oL+3EMgRFyGz2ATMq3WEj0p7QRDsl+pNczMe6Y0YNFRlHf5bje41cC31/qhcQJpa
FgOS42BhAWmgj8I8QwwvROgbHpI8yrdyyeK8HCFF3+6PtmWpCUTYZY4UblVMPkMb
jMChj+i0gJ/TIyKOh6N6qquWONaEkPN7eIXO5z8Fo6KjAGwI/ZYyWOJxIn0BzRhR
vHAPKHFuOX/EBBumdugPm1TtpHCqzmSb8vO3cseH7yW26s90N7GKyONKLnN3oA5R
ujTK+4YtuCZPcKRFtUDy11jO581FLG6i79CNolClhizNDzw6yiYzA0eF+2VPwIyt
Z7Rpgitz0iaaUN7oBTn7A6YSAhwSPIU/yvqiWszwC74q3alK1s0WZEF1+/ZaFW2A
dxIzPEqCxGoAqxAZJNyUbcMeqnxnHy0zGvqSD4la79v51Vwu/jYjK+nrMMamfECd
bJyMMzWqciSDNvggnVEEqLbNE+jZR708WYOtOeE0hYpNyHfdUj9uWzTDRafEy0Ch
stqwuwm6fya1VLZ/I6gv43fhWViV6jYziAa5a9UZ/7JVPohAYnNeFGgTxfRKMb0t
MJJz3plo79yaKaUdJjeuUnXuSLtRra4BFfuUuotxPpi220K8c/u/2sEfnUwbPxF5
MYmloS9l8Ca7Ts2+XdLigoe+a+bz4Ao48l97BrODqkI8btGRPE1kbea/YRCuANVC
OEVAlAJZGcj+pVcQur7BDY1zCsnUi08wjVhMEogGSkE+KOTfF54woAsiBtewzeAB
bEV5P0QDZL2oQLFV/ttE8lK4XPnkZXoL8j/rDV4PsE69ZAsTeIi30eHti5K6TmCS
mcIXnAN66G7A0zW4yJ6odbNwWYhqdrsqoqEC7wGCXz9ehSoisG3KCM1f33iKBDiZ
+ZFOk0ifTM9FfIe83Yt8ADmUYjtcbdu9kA4Es86/1eTUSwTe8wnW+KyzpiQjGdJF
JWXNCvhTkZo28Ly3yBqYPfMesrse7113UZlhaCKJTQt4DvMTlRjsH7VQlbQtA4ww
wicKE5jXypbIM96TkyXxh1wI/UNocNcUoLmrNL1rfNapv4Jdq7w9TX+EIzj/iTW8
DAEmKzpOfYGa7D+2m2ZTXKxxOvzsDuGuTGmiwM/K+tvpIwsmX3pmyWCc8iaNzMlL
2kF0aukbzMCOPHj7NZ3LRSv+zSl9OzstK6ErKdDHUBLRc8fHGE8iIeybJBv/cW78
sUUQ4m0hpej8OJ/AZDmRgG5FaqY7MCvLXZqAHsMqURUx7GzCms7GD3UugaTJ5cym
ii68U4s/4lXu3q3ma6PnsHpb4cmVHE7yA2x0k42XrvNydemaoEJuT2YA/nnMP+fc
hjM06+G0cBB3vayw46MouhdqbUZTOwU3vGUrT6AUvRJPYhxmhzqch8007oKBkJ88
agh4duzYKQMt8+A5p+4jHsht/JiIDx6MZtZVL+vQXJ2gE5SugFM+BVVefvhHsiLj
mlT77I7ZKnCbKY1LOc5p4XJzL7e018rr6wRFu5wLTr1G2IQbzg2ipVqoQV9/cj7N
eNBbh1Qx9zrM4xhXF7Aan6253N2/oOyYonPCvi450uOO8vS0LmolK3/YgCLp2fnT
imTtuqr6T0W0/cWU0ZkehlgPCQlzs9C8fmx3w4jm7B7kSiXoLe//eBxMs1Bds/NZ
3Q1xAjZCKajdZaWRSP0NwTzRZvYhp+A2Lqn0LzZEgtMTDiPI7fcL7ecc7kTLZBgD
Cypitsbl2bZ2h0cnH0OSt8AGccCh8sf3OSFIr70AJr2dN6uxbGA8Z9IMGUiTnPFK
wleGGpy/h2ScVt5Bz8L2gx6/8bKACFFCidUpn8Rd/NN3yzr1Qo0Yf3FGIgC2Tfm/
1rpRIdpLR3H3Yh0dMcEXSNgmN+rAuJ7gi5xjkfImO+IwiysOwrYYiaKE1xhYR0mS
nW2aiSloSSKTXAai/tinu37Gq4c4K40hlbG/ZjkrDZXiruyWQL6rv22RQ1xYHXwh
lAVf9scPBkr6Cp3r7WgmKLdfArw9gbgugpZsisyax+T6KSF2vLBkEw9JeljUI1aQ
p97q7gnSkllpkpFQFRUQVQdnAeykeqtCeLJ5iv9+3FvUf1VMd9SOl1td8IEDZtFY
+MK7XLACgZkb3dhjsCd5rrX0H5XtjQACWrsFX0fk7Ufi3t2DOaLfjQfaG4Rqs7Oq
0NVrlFM/0kKSNO8qxZTXz4mxYNcuOxe9poOFTHR6E2mJXtq/09FtD7KEObI05rOU
hakmJ3peqjPbwXlBh7fMv/ELBNjWVUZk+2WO7lZYeivWk4/pkdVh+ymwZUY080pP
4J5snn3ym7XnoFKymZNAFx9gnzCICacJ9HV4ipB5mAyods7ZWIjY3+5eEDPbzaph
AU3tou85ajor9dOaOWg4JhR1Jgs39cSKAgmP22LpmcRkfkGMJ/MokZ919Kzxq4r8
Mzm3qzO4DwNpkl+j7v6oU8HMagnutUhCwaJSmsToQg209CKIvlrRF01i4jvZ5LzZ
x2g1svN4MhGIYFM6gm3uXwbyRWflCDH79olOLpNajajUsY8GXJOt1Lujf/pu6NDE
O0xEQhoYUCFiVbzsVCe/jzpIy97r81Kj3gTOQHf+Byx+vOHUk/YkM73zCyUSY71I
zNjKEnIgWROA62TBOTxRNNKNB+bCSEtDiE9DcdVNwlnoeksZ1rMNCvtzZM7xAjze
7NUWnMCHVskLkWi0XyFO57Cka6YwVYsKU2HlhY3Jvp6ej2hQacI2pr4mePlebz9S
TcXRpNw4hXDi9elWWvlFdjft2LfQN6VK3DsagkEFTDETACyxv/TWJ00Hf5OzmONL
f4OGFTr7nIY8QQgFMuYH47ej4SjKB03OeIHmAIPEMeAHY+1V+MdaXN7jS1tvCYIp
x9HkC3slKbQrqwghrLB5qnqeuiB0Go2NynO3DKVevZRGaqhj5LoE5Hdf3JDEHXao
EzM/ekkxbNiOiBBwBOxgYYRWX5i7fwJ3Rgovub5hdCIQSkAs1WtqeFJCKQC2d8qi
I2+ePMGZa5tA0UN7NYboOk4HXAySexP8a2PjYD7oQ25NMXg+w4ag7EgMaEFOnEU2
7EzSyRD95BpBTbMEtMYWFUSwIM+ZUxO2TMvJGRScBmPXLKk4+pIXtHlnGg8yHFo0
uVV5BmS714ztSDMYe6GpDHHy9FyLK/SO42B1jcTChuo31g0nqw7nNJFexYjJCmN1
vL30TEvmye7Xbinc6wRJFTtqUcJSVhrDmQwCGxy2V9Q9LeuB4CUFPllb8rC52cvX
pa3MNBkayMFRPbw5kmCBw8ob9b8y4v5zHzArVdMHQku6vd8e7jS7Q82VLHgD1he+
6TBQyURZfvI1l5liioRgFd60FNQAf4/0X3EAGbXrrOjiwzwjmnpQIj4Up23u9hxv
Xk9N7HtVqphUM+SPs16i7pqEqEx9CllkL/tl5bHT+RwtnrVLIlYFQ1hFYkFYiaiq
6iqkhJexqQIxdw9m/M2yUMLaWD/zsNctUuqNP+Ypt0jqaZblCGzKzSqiFFNqT/st
7zIvrhrjTSxISGDu1CKJ7YeWiTj8FuY7oEBJwYXWv8DbdD27Fk/nbnGaGAaKXwGj
6Q8PBXJ1v7pH8pgSXY13aRhRpmrDC6ERjB65Vd848nVB6CO6NDidDFWcqDAemK2r
PO22QP55y3Kaf4GlCZ5HlA4g85AWGuoLoH6JTf15jqwfnEqDI5mgz4evmkUFBN9Z
ZlAgI5L+dv/T5DrM3oBgVN22qQUvGorjwWGDR39Ss9iM/Hl81f3zmAMFZEnf12vf
67MvbJayjcn8GPmIeqAVWejhDKTBeiMqTyw15+8fBGHShbBj91AK9Ztn9BN5Rzjh
JiQoZ9Uw1jYoJ0LNDdsS42CMyGMSIgmKPjGb0ZJ3XC1sssSwDvc+B1EfV7cozZt+
63PCMNTTBxMxSO9Rs5v3AD3I+npnBLPkCTpghfdko+pLihOFPto2FIaWFKlzeW/b
sF15QbbfeC20i5mE3PSjmrmRozXwXA2/AEygledkS06eCH/VOiXQLQDZ+Yj+db6R
aHGIsAzrJwMT0zMAyCSCovfsVu4ly35i9ntFi+Dm9PC1sUUD8KCQOf17ruhvThC7
TYljVzrgYEOgTFxVPjzgfVp0zl8oboJPzk3T7Axt0XwBdF/6bnd8ztMooQ83NkXg
9IeI7jyKtr77WuBKerkv/kT/7/BmOSbmF0TkvMBMaAS0XoZ7ouVs9rWuZ9QwKbn5
jDkoqCfdGLIBYdVmVtI5YvU5eFkooOqsaYm8TUZbpL/HJZ5crcfQKzkOYUFRpXW0
NXunoyqYJC66bvYBPt5V087q8+kj7xwWjzrgncVYjTfXnon9WEOYMWbkZ76ivbQc
z0jSAKy4IZGVNOvs0mewWZhrOzr6f9IAd0WgOqfC5FnrDGBixYQ/8WDWlW6V4rMt
JTsTs7seZ2iac5t6ldR9sVS4PC/xrpkv6aTxNfRoWnxndWePs3i+d6Lwsl34bCCW
wGvYfNBVTLRKdeIuETNcL57CYQ8kNT+6le/YjiZBf2HqXrkGBXA3Tu5MS2VZ6I3c
I/BlZt42C3ZTQ5TJon0BFTEMBOYAJA/bVRtTXE0s8bQOA1A2RdV44KKZndMDbWAE
pvjI04wSCPSPj810ynQ4uV5sHVuJXcHkU5hmCFk8gH0Cu0g4UCNEdG+ifkaT00Gf
V8/v11LFWZ5ZbJaOHVBdd12rOAZ657rLupPkyKV8dURYTtjEQ8OrjrKUKsK0AvBF
Q5XrpBD85xRl40ABs/lOSqH2jH9PjPiE9rcfRQKrAc+Hk2pbgu6bAVnzO3rCt4kx
5oUoeYiNmKdr72ifQv6obc0Sl0bSQkyyghXuhRKMWksiR1UEGtIASSxB3wY7CyW/
MHCof8FjC+Q2WKAaH4hS0ySHrCz75BziZWy/S5txI/Huf4ND+4QrkNGPybRoBOSI
cH/cH6Di4PoMkitDvjqin7/Pao0GLzUp08bpnKbIfwCJmnvnVdjq47Pb0bvMeSTX
DTyu9oecgWHyEBAHp37YBb7GeVktVdU+tTvRUGT+FLbUTl2r6CHqhFmYxdMlmKOX
u1oNFqvxj0GMqTYaIIBsdUopnodADcOwoPVdIgyjuqMgz3V/D10a8DHbOZmTsvvu
2QuL10FkocDFjHNXbqT9wWJrGNHbxIC+XLy6X67TIcd5bU40AzjjaoviXrbPVzLS
rhIbfQfANjlRkO6zBt+ZkblpG5UXE7NyEKsMWGh+QHACSvCsBMFxk9AOFlo9a+3m
4XdP24kjyVDCmzEhDdJJI74BLvybCRnZEphtNxO768qRcS7Npv10jIiLzHU3tyvG
Y2PACjdeHD5SzzgsfDtDyyZ0m0PjmzqUtGNKkntMH62ZOePl4AjSyJCbf3QH0534
HUbBuCkELC9co97bUVnGQ6pEw0O0RI3uZ++Fl6eAhF7pKksyi075kOhWNsY56y+G
2xUMvptPmlpwqUKqq/tXUaFJnOu+E4jOJj2lUBChUXh93/gKxz6xGvLa8rKj+4GJ
Qgq9u07lcT9oMjHlAA5k0yxtDXz2jn3aScmNTtjkrOPJaMCq3/e1/1sDm29Ur9/K
rt+PgmBqUmwttRh28TbtGjvPJyG56g8fyD+xur6M/vxzISG8896rR1nxHWCXbzbM
sZFljXsivGQtZYunuZjFVTzd+57N8UsCC1k9eZ/6m8c4JHlhgr04G4covWW57nba
UE8LUe4Gk6xzBxZFjzHOVYwvdf5XvtyB4Qiatx3Hui2IbBYKvJxYYz07i2Tra7W/
Xw9VEdl1Plt8Im3ScA1bM5ewxk7JwlOT9+zB/HALcO0iwZkuHfHe9lC/omIeBlF3
lw5TgYk/96BR3ewjIlB81u6ffulvAogcaGHXtvCcSZnM62FBWzjc4KzEwDhY3yQw
P5RiP1o5QI0myLZwsrDn+gEVCtnKI0rcRF57wPU/xX5WCVmVEyTs8BxzKT2JRXEi
x9FpbIMKHOrAiETN1T4SukM1+o1WqjhX2+0Pqi3kdU4oKk4WOkqx3QyRT+q8rMqo
VwPnmP77uNiRMp7q01EOKg3pXcIyDNJLzfu2w/2Le+NlYtf4p6HWzO1sMDmrMRGT
ZlF4NHsIi3CImMYs5xxoE9Yh3QlkgqWPKaModFKc+PT3Oi8W+lrZ18r6zBi7MEas
7eT4pS5D50gLjqPN419DIwCjuZVCJ+O2R71Z+kREpCPQ09mJDKlpuIkmc9ZcijT1
Emt/6SpLxoElXkCbxpIsdULkaznb5Jbh9ARUKgfhBIS0EAPfZYhUyVvLmWZ5xW4I
pqQvq9R+f1Gexkw32+CN5CUYEsTLR6xGNi6NBwqw7s6kL5WOjF47PIg7tiCK8C7u
JbKvJqnEI6+mH1CfWYHp6RGiGKieH23KH+0UB+aULGXOYl1UMwSJMqy7Fta6lhc3
+zEBP2vZ8Ur3t84K4fNl6YlXXPnrxIunCM/+5vYWHwQUm76oJwpZtVI/9kKxIcI+
BGt4WyLvQH2cM4yRrhpbkiAqniIdiyhfQ/sGEbZiTnQGbfgt1QchpHhvCxuem+m3
n2wZlf6BgNjO8sLPD0a4uK/YKyF2r4sQVe8gKuAeJF5qN5CVf+FhtaBPFpCv37TI
VJO/QHStYhusBzLCiBV9iduwSNkHcvzabF8dhQZQDSNuy8YQaqGKkoeog5xicO0x
524ZLtL+JvSJxD9zUy4NvfLton1sI27mmLkYVPKIW+iA/4tA/4vjFcfkIxvFWZRo
n4vhwq5i/p9n0brzThUZAzw1ax90cdi9ZILpk0x2r3pd45CLxtqPu3KxLhR9G4jg
KnLOU5Cds4y5lX4G6UCHOxs6V2gtLlSc5wkA8oyda0IpcscOVkdE/7ZV9cgoa5Sj
22Q/HGUkwR/MBQRkHzsY2KjRQCYvhd/UgUeWasrKkFw8YAETBxASjfffTuR5ttPh
dhA4Hofi3ncOmcd/lv1FgLlGzAOjl3QHsd8hLo7QbXK7/OfPm9ZPcUaI9gde+LCS
7iAUHn9p80+yJATnXcZabVeuBw4e7LtVF5YY1koS4FkOC8L73WxWc5nropxEwIvD
eS7/dMJ53+1fUWUD5LUlMSinUISP+MLJKvUO72nUtMdIEghd6qyZVC8GgqJ9j7qH
r0sWd4TXxql/L+A2361ffMaNiBRouytifvKvVRfc7Ds+icTVYIL/O3oEszUkAWTk
QBUZW6ROC2o/suBwa3kqdtDkAK5vSOjmNpi+/lIC1XFzWnd7l4rjci/U12q3r8OE
weQknNifr1AMXhSa5fGCRpFAlguPsUKM/3iS9ofY360+7OgHPThlm9LhPcCVbH2g
yJiafjpvTorI9MhXZ6bQPgmsL9sJRfdF+3GEKdRRYpBLz+LFUvgEl3Bi2qWlfgXM
ThClu7DskAWwEn390OEpiuVxUrkIFfpq0rinWNcMX0GNTKYiNeoupKezbWW8q80J
4QOoaIQZ4rDPO58Mt2FhBec/LhUqnyfRceCZYWvtmzqS6Cg3G0tLAnY2hc1Z0xnm
MPM/3LykcUizqDgTI2aB7yZY/vNR0QXrr1cF4JB9Lp4eLMWC7nmnaUkG+PkROJR/
hvet3f3TkdpEeAQRRIj7NzL6X4DoYeq3QcXyKujgDbu1c3nkja//RLy4xStFG9w+
+fzhjfkTanj6qUSpGrIXl+lB31TfXOyBS6KZeMp0fxcprNac665FOgx0QBhVhlCO
pVUSHoP0leC7gxGhtQe4p/6vZ4dbog3sIwoSd5NfR/wjciHiZFIzXTsc9HgxRT98
lYL7Br+XnwnSNMaqcjQeiD/F0LC0WMkLwUVR9dSRgQ37WME05eBQvvAznvU+lNLK
ul16J5AZQGOinuGOymignb2xs+M/wvqKMVwfkqkvgadrANDXkc3J+SKw7RjTaYme
8C/PrbycF+B9YPfX3Y1jOW3FwlIUVlMZ7chtOSHrOjJkl4guaCsvDzIhCiNL62v2
JPg4b6dfALSDEqw4re3NCz+a1ATqERCLVllU00EJ4G8E2khkmAsXghZRS89Lg4zm
gj5OsnqbQk/ObGCUAFKKUcBeKNAZrCVNriHffohwcAcUeLIEiD6zS7CHeR+X196M
4I30Y+uHpzzZ1j+tQWbRrGtV4Mkh2idW83+v+wR5hyez8XmYuzikixSQyMGyV/KC
23ApVK/ljh5eFTSgn42F18/J7+VVrbhGqw5jUXSnUl+pLdhQLq5qBhFl4tJnWTFo
zZm9rhCX2HGSmeDXnqPptlxMiQcnLEiMyJHcO/BG2SMqluSE+6Jk5qVE7gQ5b97u
Br9Cb6PQG2sz6+NHEdkmvnGMpJcHEk0xWHtS8r8UmL4n1FVN0ogHOMFPvDyvAtUY
wW6Xi5V3/vi9YLr5lYOlCGf4xY8qQP3CYGze9YdoVvIYFWi0k3zD0yg+O3TSbyhV
8aBRHvlktGzzQ5gZvYLzv20HuUika6ODvDOiETjk9IP/fG7FFfaTkPnH8JrycrVx
SrR6f9PqfBI8+VLWyCYXMfx8fSqlgVYH18tiXURINzKD4BqR9seRU/rlA8Ykc0KB
arzznCG4iEk7a+d/X0vp9KgeB20Lh7Cgkl3INxiHFM8M1cdioVZ0ce/yLom8+ggW
0ERPY71L3sanz+ksoxbMAcIZTbm82FJsYlC/GFyY+I4Qlp4dEthrrd/gjuXP1PpS
lXsb4tEMjKnz75Yj7wRrD9KBx+9XfGWLTjlZNRs7NlXXyU3x4jFGflcXCtlwaqLX
P9+yVFwyF+rFuJhmgbhyXfV4iWIfkTmRVJJKRDtlBYZTfBGlwcA/lfbGtd/tZ40v
PnkgyXWozKDWoVFsl405QR3M97CIH2DOQWOMpw4TF4jl4exfACp7+sCj+/VF7mVe
q1aRe7mKBD8gvozXwPYFKHczIcv6ZYm5DuDMA5TQ9xJ393QEassfMtBYGKjDG5Bv
dHMBMfM4gNQLHLOVn8bhheN7pJYoo9OcHLAwo3+JMQFtPmUFOE+dXSLV1mMURgA0
BqiW+ylTpSnNtNS0Mzt3gyTVgVYXHymvdnmx/EgDyn/wA5ZiuJTYLmGtCHZQFspu
a4QGxlPQtquOHwKCnsbT5Rx1+M/hIGSNUY7KohMoTAYeVOnHu5qr2qyvztQ1qlkl
IEFVsSPvywfzaTURaMDo/EGgyydopw1JH9RZdEXVT1Rn4fRpym7RpiCTkQ2+dVFY
Zj1ER9gsHfB30TBUdqyufE0plrJT2zBK4Gtr1E5nijN+PI+0WM91dnCg9UWXcKjE
T4eRRVKr5CbgL5N0CYNu1yobzsgJau0eRLjfdWFu+wDRSfebWU3psiBV9xmCizWt
tg8PGb5xJGFqTYblq/BAnoQRwYeYX6AN/giL4x7bo+ydKMkca+XjIn/Gmx9vGd2Q
Ezi3mkUHPRaF/xYeEgIjnkp/xe9Q9wMASGnxWeIYIY+Mk/YjCjDNadM2sC84jBgD
Z/5TFwPYd23XWdmyIokHXC6X1sWE26guXKGq6dSAnnVL2Bpvy9FfAcz+gmlq/l9f
/d/xQtOgHtcOoAZ3m9RKFgqCBWq23FF497SfLsOxOY9fkA0ILLe4NPawZiBhNfxy
idVbKwWZXGe78rA5slMSI1FoyEFrGuLrSpW9Cs687Cbb2wpAcVwPqUhi0HPaGv2x
UHhaJBbfmTpS6LvRMuRzhboKATyTRQzSIEFfVB2tbuBoIFcKLf+c4xZhKhNr42iX
iJWvRtPhg0rm8PX8gxBmRzkAstWPeHq6qGdMoITi4xP28EzOTt3dIKG/mbJY1pY7
DkunG6KKyZFz3KQgk8xqocJhS+n2t+vX/WRgszeqATg2V/3XGFIPi3s1AzwpmZoj
2KKK5Ul3zlqpRZ0F2r3QCZMD78E6StK3LT5YaofTwAPQdwZzp36oHeEgQzEfSEH2
oF60c0nilSR4tYXelXL6AElLkdjlzT6dLQH2VME5yPX2ECfme6L4xrt6GbhrVtPl
scwME6BRyxzVSajSjDb129/DRhtgfy1QnTXat34e2xYcwoWlK0oY/32fQ6IOgsvC
GzPiRt0jOThl54VrLvLm9AbjUwxzTjqkSicYUQHIglX17dKiu1vgiQCMiulCASGe
t2KkuBM6uo8SV3gNxCnAgnFbY/3gAT4pBq9kwvZxDlJeHJ5TTW/kSixXJwwHOyja
f4G5iEQaiZ+iaGKuxvKmx2Elb/zIZ9PTn5lIFtueCMo/NwBV/cq6IjS7zlxTyNZQ
Uoz6kOc7TzxWijC2PaZyILrKz9iZqrjmWfYPcFGzJ6j5Zbno7tfVgyXTiihGpXq9
PtOoLQ42LGQKm0Ki8IwxEmwpcIs3PnF2pbonApkrsrflOk2pV5ysaiVOOqjGY6m3
TYfsFDb0X2Ra4MujyPOZ7brSo2gQFnSqhJsNvs45CZS1reD3GyRx5sgM27PTbCta
A94Db1qa8mIZBGMticRCx4hB4NmfuLDnjXd/JRKjQX2OUNd01afsCfDVGP/m6Dgd
nXTkkaJq4ifax+C728ZPZ4YC74KqFbltt1kT5r7DG9dggFrlMipMgCjpAsJYS0wD
xaHzym3gyGOpCauLEAVkTy+pIsCsw2yobWHovXx/6vNOmKnXPmq4AYbguHk/TqFy
KEgktu+S7RiXza649rAd15a7GUV0V4dgPCeAt7xX0UvKGX+xv28cLHmgjHJnprR+
g2J7JrFwwKcaYN7P+GZmXSrlpgFgX0K2a1hZWP44lEz14XYqyrV9iZrH+g2RQGo/
O7GH2Hy/L16IKzZgLWdjptSgvmwOWDPD7wKqM2+qfWmVycn/c9Uk9cMIVNLmzgKM
26jnc0VzDHDduQ/MNoprP3jPVvrne9zoIPuGJcEPccGsKAjhca5jDu7Kp2+AGlic
2Wxxx3qwH4y7WhilJK4iYsG3ja+sBAsqgShcHYUuLxdH8Jgm8LuZWCYC3iwPnGKy
bUcpBH+Kb2/QHfuNhIWbdufOnvQ1SRzszoqooeu6/W8QpEgmc0BIrLmC/xjOobFp
XeiIVrVrEq4juTjEowvO9qAl8Q7cNeiR6dQkjt5MR4NYkMLgfy6yYP/OAcvxCEBu
lwxjcG9yTxtd97HKmxhNPUjdOXKRcjAmT7SvPT8K9Qe4TphPD1WdeiKeMq9eMFWa
ATZB3rItqvs498Rin39koSRpq0DBWRvm/Sw9qMwYsdPuVjcTwKD4nXQE8uE/To/t
UwTdgACCjDMpEvpQzTgic8dr7sekhIGU8d/fTo3zgnbwuqtbLamayC5yiE4kJ/RS
bZ21YRsPMrtimoEZKK6bp3m3xG4k/OSpHTr7n9zNEoyWJxwrgOyGdJKZgFiHlxT5
gQ8ZzWScPx0AewWMrylYzDL/fh5lN2GKzENIO1pU1p9455NMjEoDMfFrmUhb2aMO
gRKl9Upj1MHnJMjBXcyoIw7EiX38N+vw2c1ZnvdCRwf2VbVoKM29ksma8EodaukQ
aNok97TZJFxLFdZPhYWN05YdtKh3fBAJoqApHAJRaqsT3QXQNhZXg9FL6BvWXDY+
+dJdDQAs0KIT9dFcKbf1EygRrdDTsA/W7P23bRb1KOnNFSlSPclK0+kKOxINJxe3
2ECH1uALxRXMonkRMFBK5aZQAszlPCjDLsAY+104PqNbGJtxBZMd1XQH95nWx7PY
1hMGNcjvaPuL6ZPaxuxQYHJru1tJG1K4wvQihE4bVa3Xd6nTt5QKbHekzQeeoWmo
aAStalEnwTIqwXmIdiw2dkEYulGA76I7/IKOZYkq5QTvolWo5skbEZ0l+3wo/SOw
7wKu/UrszG8JGqmVpasImPvabuN2k6Iy79Ggasz75Wqb32zzErP6DKUolzVIyEvh
5hdychCO/0gzkQaGjFkm/UWnyrbfceJXhEu7SvYJjk9hh0Y18gvxWkF8w/bBkPBK
n0B1gDQxcCvPr2+MUCBqrefObNEQWh/DcyWizv0gUgraidw+2X+HwqxI8KGolNqA
95Am2tWLsaQrJNRaZGqcTpbKdsKx53OyeDs75Bv/MhfdNtRw4tXd9Mx/RvP5sN7O
/rLOVgE7sE6bt+rivvReXV2T4l9t404wx+nwL9cSzqGogKTiWUn89B7Ivo3FSOA8
/E4HSTxiTpCxsqKOBZAt7dMP9P9hs5hmEzB5qr/L4gMIQCu9j0Q7b3UOzP7wIvrN
qoUucGKLUL6GOh6NDM/BNXw5WnxSrn4GxdQKHXDdFOoecGe6plkCdiDP9ZoWMtny
xiXhqUbzqA/QJNsgRfVRwGM7RfRjdWrYIpLiA71V7OqKFAuKQ1CvuWsWN40X/eYU
VsY+RYGm8cCJkZ+0Cyhdc0bzoFOWeQ2qBX9NJFVRHiM9YA4T7WDzE7LGlB5Sux0J
wqHZ0ls6VZjQPbD/6Zpq+eOvKxVkRqOXrDS5uxTleZVS4EK1Wh2AwU06E8n8LV9Q
ix7mQ5GVEqbn+DhpgL6LDLgNrvpe1DauyqMuyeZB4Tq72g6cYAcMGhj2fxnaSfXM
CJ6FQI5Jpe06GsaOLJiGnR+yraoVdQu0RocnwpQlV+OY76w2OSEnxNpUqZfbFndX
spzmUCIKw4i/0YPz8ibefFFGm9+wEEpEBdQ+D0ue6xh6OIIeeubj5F3pU5JmilvC
vVAxAieJP4IH4o6eNN676Sn8HNeu5u7854ywqcbhkaoNCLMU2I0RLSGM8yvJpz7E
d7m5Y+apZ5sPmkjdcVMqAZGefmOoNjEXK48iuZIDJ5NPGko26Vs78IxX6TleogUc
0w5cxp5lEaAW9d6OmAgFugwI6oRX4aNjDlINR6TTVd130/NbkYMrjfQhzorAlpnt
dRVc+BU8eZIFGqPJZbGAqEN+vZFf4LCVzAlZDsEt9LRlSXLrhaTfsD4fjtRJDaLA
qI6Dxd7Q6hyXTOb9Z4H0JwWl+ToACG1RFgKwDf04aOwMDC0MwWKyFMiLWOj76D4O
pz+L6yzf45G1tZJGk/cioa37PtqL1V4cR2VikKiydF7IhpR/sfQgnQsXOH80Yfw0
GDeihXgd1D1ImcDVjEkngwagO13L1HjSrpwwk97EgznqX6sG93wg70nViDQxqaJx
CpBCSWiydb32Guov08szZp1vBbyMyQ3QLqloxKbrLNx708kmrKLuuM1S9V4hshJ5
VzA8uNmJyRvKQSmxYdaTLE541GngIXGKc3W8lC0YwZMGBoBMe7LyD59Of0S/cKMG
ikEASmnBdS68K7i5qNmIqMobUR9bLwwuC0+HDfUmw9ijgjKZJqxhTul9sqdxTxsf
58JfyhByf2Z/pBM78L/htIz1LzN9iR4Hsu4OQpa2vAo2xQh5jKbBjmhu92VKduTS
jPy+ARguMpArQuG4zAjMYeo/LIhduKphe95z88MldaTzoN5J0LrKSHB73lEPr6gh
xkqZHfy4c9gDFAZoRDntpaYxWE/tmoJkSVETCc1LGP17oGfY+TJ3lmLrdj97US/p
cDvH+qh8zR2V03f7yMrUeqHNkJ39iO6raod7Zug9Vj4cBoLEM8jq9u0Bqf9A1AWx
4ayeloBXQ/0PQz77S9wGX6l95DvjlTvqQoeF589Cfq6KLXkHeWeSbnOUVF0R/JVe
7h7FntwCXxfB+1bsytLU83nCmiVa30nklTni5PvgUgQrOvneGAr2OuUFh0XOE/Qi
tuEAp1crE6vx8in1ww2OCoWsTJV2ph1Y5bZZQc1UQ0fmYuBPeLDF89jKvDObkXUT
T9h67vNYQSTB8BSMcLE4tXaC5komwUaMxjGwIpf7p15cjOrMB3S4AhWVjF8wePTe
TZ8cVBbycdQMgCbxIqOm1sSmsS95bA0VHOHgG2qmjqNKiJj/q5+H2q720Ozpd4O/
nkPaBV+ewZMCK1/1p5BPttTFNPqtMbULTaZxwgJtNeLv/YUEB3kLeM/hN2n6qpNn
KRfW9OAko2Ey7Xwj1gKHCYICgDz3+OiobYqegqk66kZC4uWybzKym6biDHz6IkC4
Y1WYS23zXKDp8oL7/TBEpw1cJiFtqlPMzCounhyCt6ie+xx1xQ6Tv4KL+JgX0JCq
nk1VP0RfHUyciRpvJAcSfkgaDEV5UUedSbc69OLfF+meAeIfiZ5dKe1c2O82U1h7
Tifpjb9O3Q2w4kbzgLqQNlbpwFSIBvuiCt+d0v8O8D9uccuogDGml1IrOrZUp0M6
xNkwFQ/YpNgUlu+eQqhKgjY9wXd6HxXDG48ACX25jbZmmtbkjJOp/DqAtEw8Qbs6
nN6/bwX1w+FLVGjqg9iuU9Ei3eqt7AdNeFrNZWVjYsRzY9WkMW3BlHKjnjHYzAUK
Hs94cmCBdEpqGv41qFNsxWfOUqo1DjqzV9sGjPlT6+DIy1bygaOaoe7hw+NkMbGz
uq0eQS3Uj5jYxr6CcOjpv9saTYyDSi3L6ML2McOhy/g4H369PskM8x4qvx8Rt6gT
8v/Ns3Mq39vC63RDIjix0CWcj0SjPVHWnAn3WZSOmNrMO8Uufb/qmTsiSMRd9dlz
LTeXvx8UMaYx+eo+4bc08YhHI2dJwx+qLGdoib3hEAD4RrUUhqsLg8L71lsE+0G9
qrXuH8sb29oGntEn6pMwnEW6nnuCbDpj5Sp4LQ3ib6sSG5+QHd3R1jlNsvJ11CMX
16XAWe2KeKq5kknFuezXRuTGSXzqG6Wiw3rp+qezjLDr6KV3gv/Byz8JRUjgGuBS
mzwGp2MnegkMWnx64mkd+86yiAmhtlAKKCXY90xq8CWoPv1o+ifQs2eM3xKVEd2a
sl/soiYfQY297n0jDAhegjMVnlQPICvAbHfkWrSZziihWwb6lCzGISgqn39crikO
VF8EevRD6YIiEL8BR0xLxWPRJR73dQgjGYtd5g8rztCa4FBIcty6idveP4OvA31d
B6GPx2bQA31VouNfV3bo5dtTwuLX0JsFI/HGUicKA7H3z9ZwruwZvdZChvzuDD1D
N3gD5Suf9waDGP2Mrt3E4jU8Cbgl884l31+Lmx971FoBh+egB624hEUkeP0cQlSS
KgziY+Uyk7uSHz3KPAW+ws2MbwiRZYlGCvtVeEmvL2DLyFpx3o/sulL+cnUCh8Sh
yQAaP6ZWBqoiW1S6qqnP+O8xbEH/D53K3pqVv2HZTSuaVoo83nCeyIIPBEjF6GTc
pnu4GxpEeY0rMaKnnyMQ5a9q81b/Ybrt+aojVawrIQV6IEepEaMjTPMabqztcXYx
vHHdCe/FShcRHyDlWy47+eu7hRScY0bTQEZCmOaH6wgDta3vzNTRALFmSCf2frCX
K6hqQo059CXXOisBAvxP+1vPD61zYjQMZJiWq4rPRqY2tNHT7en4qdRazWCAJmup
6HGYjBQG9BBi7nAG/pSwPlUkDHKAFLqxImAVliHrApPzwRANc6WK/j4758DivUYP
6CBCwb465BFqhP6pBCytiTldTCRM6MzvqxYXKbh/G06+Uv2XuhzP1OO2HXy6+sXH
akafEXT4AGjNFS8zgleKyiISSu0x1aX89eE4U9tsUgPQrrz9LKKECPW2HnedTT9k
+fVJ86dbBVvITt0NiFSIqsqY4WeocdPvEEMdQDXWpx12Tb5TgJJPcaB6KxvStfni
BnGJRO/P4LEK3EkcIIQPrJhA1raVKI4pD4M1oEdNTySKdj1+IIg3teu8H3j5gJI5
0KcnBz+TBIhk6oNR84DNQevf4hwztZHh8j25lDtb7rDSKZyxwFnqBIF2vmCxsJmR
dDB83oFnXZlbqDmxIFJ4yGMdMILmhpP7RcJ/G5wT+JyO2PZkbyGQsznKV5FyAqQ9
vZ0FZRFiDIiXyEG35jPX5BVRkIPA0a7EvB3jeUrJx+0JlDhwm+0ut3QlpA6XyMXS
MGSEgMNH4wiDi2kY6PZElRe1FngPhvSLcaUCN6s3+/ndXvugx6VOkaVjJEHbL/15
SY9zoh/y44AAOZQAfPkRrB7HPABKcq9ArMuf3qPS/XMvi+fQb/LH0MGPnE7zfadl
S8w40zXMEaB5HVDXvX4O9oERtVZZ6xPmWnjEIvD78vxjydJoLopAsco9MCNoRp+o
DiHzg288suhjOM2pr3fo9vgTWaBPJCQFw+QoLhbbGnLPV+7ZWJ6OUsD64UgAJ7Sv
xKwj9Kf6UpMp3GYYACY0oouVt68eGczjFgnH1NhH5sZXTpEBXwPBRGZhbVVn5k9Z
R4XvVQ57sEQQLc6qJIwDr4ez/VkTStGENZtHF3i/LLXRO4AlB9LzoWfP7u1KpXbU
3GP4ujYPU7DSeJxAQZ2MrruvP/0x/NdvbtFcQc/e4lKaLIeMDVFhBcyRVFz3Z933
HzoMccFQy09iRPL8TGd2XHQJ7R/y+BQ0eGXUPyhHbGtCkbPebFEGnEUZLk9QDUc7
WU+cwIZluMsq3SfVc4dCGJt4eaVqcZ16ESZT9ikqk6pUoM6plw3+H4aeq6iXUH7r
+X7fxxZZpePbLurI29vSNcABd/S9U7WTevJlw568YD681SCo15hjobqDehY+Ifmk
KnN++GROFiYneIw5YazCKyhzD7hh7jfclOZZaptQjFLQipmUnb9gsT3PR2g5Xil9
ocXvtXnIeLqFPL8RXTRAz6hoYSgFV0Xz4USFSuFEwFsr/R+l/UQBbeGt3X+92L/H
uynvNlXk4f74TLbukoRm1xsQZmYa8foI2/pQkT+k7cgx43bZWswAimGVH7ZkWb3y
5gNcj2cIdcSRcr8gCoVOBjtL7RFEZCeMMyYTN5TLNU3b7hnlC+UqnKcAqv46DCAJ
tquhuFuWGhrMO59+hpmExNNcgLaBH+YwinjuxoNRvV/iMgMddI3dmwXJWYCFer4X
t2H14Lb0l9woXd9cLe5HAwf8jaNhTiVGCf4cgKayI12dVVJ5Sb58CuqC9nRSMgtm
k+DY7TpCTMs4Gmg7tRgXJNbBW+fdKfwlw3HltG44YgJXRs4J+okypsbaAt8syLTx
lfVBUMYz5DXNC7475m7JWF7UaxeOCDrlZc5ATc9zzEYwO+wOG4uW8cD1DICeKFWE
VhFzLuxwc2pBQVNPuMhHeI+DIBmp4oNxwh+l26R4VjpExINKIszqB36Ko7fnP7yR
W7LDagTKZxZBrJ+/499CS/CLJt/mkEpsYJW7vQnU+CuBqjhHmZkxv3cTLFYSbEtX
iXAc/qnSacstEY63G5DE9jvTLxk4S1Y45tCgIqsDKka50ZptOZUIzvcG8paXOQXS
FuwUKxXgRV/fnEJUmYgtRJqWnrN/4BtyvokdY12P7CHh/XPUqQjALyRuwttlzMQT
GypDyqcE0bRAprfLN35R6ZEy0vlzwJ23mqXsA7SnZV8AlbG6pFMl/Sybr6eZkcWB
FqkOlhgQSru28DN2ooXfMJuhxPwvW5AlN7hevojU3OJnd/wybWnY4jt72DfvmxYE
5pGCvf+wpROm5i/Tmyaig/8RMbGaRH/QoDgBtFmrbgzrZoUQKaMaHKHyY9Ji2G0N
o0VgM4/7CUoeMQyjVxXEwBvzK25fq6wfw26UrljWqypAz74Q6D88oy9X0sihRZYk
S3bivW0LfxbvevWBMhKf0eG+y+4bqThMKQxwaKDrSsCjB3vonVT5M3V6UJ7i7wGy
1kVVhsUfxSK3JLQu5Jq50FI279Gd0LceR8wyEw9YGWY3xIGej6wXVMx7pY06Crj1
zi44FCfTj9EuGKbOSPlCzD+fIM8ufo6wAg5Q7c2Tu1tFBLF8aXgCIeC7FnDrg6Bp
ct9xh0ePLF2Fv4c0C4B/VyMy4Gjzt2UZimVF685vjYkszjD5GehcRWLl5/Rz3/r9
yk01HoGh9bv0sPD5NfONlJNvFt/oOyfJ92exXd7ZlFZx+DSaGoi2qh1CYDrPpOFv
dH8BvBYOK1nhR3UlnmMW4lG25/RAMtOnlFC8RsgT+fQZfDsIYErq+Lr5rAdHR0m2
IA5X7ntsUoQ9u0zf3+Pi00smaIR14kL+GzVwPgbqiI1LoYeLxXl27QgY0FTDUsMN
4dPf40nR0IoEPtI7/JkYzsIAyNQX4POnCNJTqGBB1bPCfFm9h+cVj+Fq1pJfQELt
TxW6dybf7c0BLHQdiHzwiZqQYVvv3QpM4VPfX7naDOHxPPT/y1aWkAJCmztLaJW4
hox+PGNbtONK9mYSEP+6d+dl4Po9qI9wwNjVJBf7+6T/ecKkL0+mH8cROP2TTBcZ
mN13ujx7WsYKvRg9qmrS8g1H2UV39M0HQpweGCSLcpUxpjYZfZXnwraUCEW7hlO4
LNHHFlmF89qm8PRlRjlJueNrbUcEB5+yrobN0CQ0KizeRIW1l6lQsZXuv/X5kXif
Oe92d70UoBRraI8+S8QlLMiOeda8/PZ+PIjK8Husd5B8s9woT4eGPa7DWnaYXFMr
oiGzdfaf034Sd980BDj7IpJLYxMce7v0yhEkBbvPXGxc+tKPq/XfODPvdFCLaD/e
RnbzyHUQTk566ZST/+acjsmRuLG9lrN7/NAbyHlt+DlNjr+1UM4GvsbKKGgxFdBY
PFeDXPScdtY1G+lx1sNSdgdp5vrNm8MzwLFh1gpRnHhaxda+T2fGfrozYR5AcGX3
H6qDBnh1400MQBieWiyRsjGtHz0bylbCamLV2EJUWIj2Zm1mNsuWDx8YuHzudvdV
rnivCI8TNWI9+NxiaaLx29sNojQQimuVlzDtvNoaKBDbWoyoJXJS9EP7TDu4Oum4
VP2rYn/oGBdMDEqn5Rr/Lg7a92NPsZ4gjxN6WA0dwFZxm2O/4wpLBaqiHVCUcKRW
imMa9R7Xx0mnPvB6mWnBLZ3Ec8oBYEflFPJTDf2gPCfHGQiI+AStQo0jEgDEmvy4
GSqkQxhiP4/dIG2kTTnILYb/bFyqLPRfzRgSQ4IBfdOLqPyTu7OZUfBQebXM0m0r
LnZv+3OYSZvDIUZYNIRH2vpHnqmDW8WNAGrT5ZbNm19rNxGvEMPrJ2Tp2axaUCl0
nJvgsCY08cgRDm1+PpoYSqrpHZoIWhREE4BRIopvCvUagC+OOFDcH1kbagj3WZLN
jihf/zvX6fl64k4iZLtCEElD/POWVzWiIT32pNV8jWeh3wuYgahbR6J5DY6QmmLO
p1NJ61myFckQUnLtVsIotjaDEg9m7selXNNR4t+EbcacUu61pWadHkjv0KQePH9O
FkQm8G5eSzc4crlHnP21KSVqHrXc5FyeOrtVjyVLfjzGEYrXSWHZqwEugc4q8ysp
b1DCREOzPCcbZS4fMIeFQNES/CNHqMS6U0JxkTv+Wzh0lmP4YIsDcw7b5k5YNSc9
I37SFv7hXgB2Zak5SNrlNXY+H2M30nvgT+9Dk2Bb61HZ7lVijW5UjBCLPTTuBTAe
1oIb1e+Mm/ooIt2qyRl08vI4H4J/1o9DG4biIrZ+il8CiEBqmP01CR6ZQlFQVrsB
F8m4lou6H+w/J1p1c93RX7vjPZd0kQFNhXf1Ot17A/8jm9cKNWKG+bpng25dFSmA
g/gvbzmvWwdDWiA5PZU0lkfgZfVqo/UaiKpx1XY41/Kqs1hG66VmxyuF3zuELxSU
2flcOSn4B1yRI8dBlbGDU5fbXOH6ggw2zNgeIXhNvPkT0ChQzflAKvPXGyeC/AOP
ahhqPnR8FyyzHvAvzbyDUeZpvB/z5tHFqdKVmbpIofyF/AVrOil6S7TNBt8Ecok1
qrr8peeqtwD++lutPY5mS7ttOheU9zGtWmsw7QQgsD7lT+/OaxWAGHpExhnKzTNg
mdDyfHgpFJVYSIC0Vqp4hKaWKHeAw5xc/i0wDnIoydB67HgA3s+uCAjl1TPjt/m9
RwMENQKj0PyELPWKjw0MDTReehpTx16s9X8X4ZNFL+CUWjKuKJLR0h7x0NPQv++w
XA4cpgGigN1OO28T3ulN2+4mmVEeQyx59fhOPE49T2sQS+fsxol8vEBVvT7Fa+Oz
/jaBwnRERU7hUeJ5r0xZxyzamQKZeW8gtpJ8K2uXcVxuDm/lW21VzcwzR7Mvw/GZ
I62nlDKMyWMVFdGSHdPFjfEige2SVLj0yxU+w0z6lope6AvZR18U9YcTSXXG9EHd
8hgW4Qou+TdeLg/ijwf/DadLjGhUQNxhk92Q7e1RNvH0/opY81sGVBubrbFlo/JY
X2QZ7bVmY8b6FwYDBFonMQxXqinfDQyTgkBiK5TGSTn+TUgTYgCS7GiH0cQYsRxp
KT6MMu6tkppMQ4vpIja3ZZaaecpgM1D5m9w5T30aPY8EFLmr5wJ9BnAc/dHpsUik
Wwkgt5FDIWIyYc8geNownm/BCQGrHh6wPy8XUpytD02w6aCxfgVw1kH3w66I+MlO
oGI4lj48LPxpTAmRs6jZ71RkkH86JuVF4EUdnYl6ULJcgk2nZnvQbYuNM1ljcbIa
30hcPHCD1eYzTyH++o/ZBhKA+flElvoVUbxOYi0JTv3MA3C5z7tAPdPnYPcmKNnu
9Mh1+SOLMRsiRThemsBO6TGa+NJ2e1MEZ12+XkiXVLXojQMJo4XRzcYBAcs0U0/7
GkYAusFnsc0rEghgBWSUWpGQT/zt77kzGf7/7bEjX2IcoaQGHXqsc3hPe6zUaSl5
Uwhe8Gfu+XQfpMVZkLB3X9WmAicdCLk0gAbQKkRJ3gPoFSNwHmO+rLk4hn7iDAjl
EUEekiFMAE664rUDBObNx1sXip8dJelY3i0vgiqarF9rB4W+XEHrjPCJnn2geLSJ
igkJUeIILG4CVGqlw9pUjeO1lH6LaRDSauNcSNGz0KLRikUJcoL1HC8RIFQv4N8R
jwsgW3jq56+bxdFaExMxBXKtdC3PZx/qRaKFAit2999tDONVe1POZBRyqVfOgvjl
gDWfYyUXj0wufJ7R0AtbYgOYGSHWHT1w9TsTw+IJhIWPpYmGhyHYRsUtBE0pBwur
01N+Kx4qFwHbKHG5wwapzLX2sv2KILF5ZrfduQj185MQkPDgBZltoawcqiLnJagC
E3cAOPk0gXN0xSNbGUZIGUAR+SAhwE74zShdde917BrM/9ISvlQA9KNhWlrRDgAo
3vY+F7qMcmJmE/Kwd8O19f/geo+DzS0yqluy1t8vVy2tVg2S/ZbqldkKx6arzyCx
f6e/7KfCkQWjaXR7hq/l5/pSldrEe7BzO1Gept+mc6YJ2/0eLG6DoZjHqhMtXzTn
p9EWvHE6dG9+pO3Nh7DmAvDpXtyy4zZFJRCA5Hyeuub+a4FcHQRBTKtEX3LJMk+1
OJKVd1stdMyiovSB173oPqKS19VjE52GPW1bfYkFjOVs64Lxv7ArW2Yl8cl5u8Nd
5d4eahnySLWIKm2Rm6DhqejzHIt1nuiYukTEcXbbTLnj7nY4S3InWcOSwKn24l8J
lAyciFxKvWJCZ4qTEGMGYoIWSMDzqoLhYxX4MGkAFMKdGOdNyqPE2uoe4eidROPm
SqfLX/JyUW3J9kr9K+RNkVx4WaKFOonPpMN7CnijUdctMrKGZmQmHVwuw1/Dtz2w
oTRX+yGimB5NXE75IlNWFZjUcntqC3n3KgoKi0Y+9cPEJl+LM67OInoSt7G+cvGh
tYSJ/hzmVHYGC2S2da8XrMEwvjj2eaxCBhwVMraVLG+f019ajzQOEqYcEVMeMnSE
MaL1SqO1YE38uGBLvQVIZf8ojwOuwalvjfeQ+/d7HJp0QryrbsZDvmGd6fQZq773
lu71bcN15Yh6BwMSImFxFdHpbOQ6ePhh7PMEDsleSVqDx24g1jbEx5babvq7W6Bw
pZXXBMKBlcuXGfdAdo7grXHd+rN/5mdsN3z+K/zLFAx03BOTxi2Y590eaY/NW7HO
UPRkCYg9E9WUwLgIKeUqC0GviAHu7aT8PW+/HgTVSy0b+LGMeFt7fcudOrM2QDzM
7ttEmCZ+h4dpdrgP+CemAJOn1y/PYOIAhL1EOgL9Ji1PhZ9gSb9ZDvki2mTsWftU
alhm3RPmdV8D+19UT93wU8qCo7iUi7SI/ldhCdwb/6GuxRw0SsqMMxTNBcURtZI+
1BihMAn/k+BbCUGPMv4dxjEW2gcyq7/UpPrO50wH9voX45UlAzu4HKdc02brAxJr
kLBEhxNyAMSnKdWin4Y7i2P7PuTTyuBZRUAGUFrE4F9p4pTC69BKzR1SSkIDTlqc
Wov8k0OThp/jmuH1N/NbZAO1580Ti1wh7d4DiHZ8PEX+aYBJL5MwOscudE0qPHvc
PFCyAwBUanqHhtdOMBLF1kAh29MPkm7chDfEOzA5vMIuj2XKCC6X9VKiTbsslOK0
TXs27xmkVrlv+Zg9LaRTU+JAEiq0xbHbDKwE/3rVYgXdnexbpCov00xrnVIQv6z1
ECQn2HZJBc4LwEPlPOMpuPvUSM9HoDnHgPIre4zwp/RCD7uqbdLllmUkxLDujHDB
2bUI0tarFx5s8nErGR5l12/71Ykbjb4laaFWKciRlc/mhYCY+SqwE9ZeTJaScjsl
qPi+iePI61Hn9IZHDbCIp0QIPYtKOqveP0nZTgrzEy5xE4lfgk+BS8hZASolNXVK
J3E6/NBrlhvwFIJGW89gE3bjt4WVy1jONj2x/MaKw7H73bRB5JJv8lX0YpFTf4K0
3SQ6Nq9h+HV1fdAehJE8qzlTOXQiVG8kXAs7FDLULIOpWf/FLjaTQD116BsEyUL0
q3D3KYqKI5Jb0r84gpZH+IxWXS3Im2VBPy20QkEvYmMrbIvlMr1R06tehY0s9AQx
xTN7z9ThEy9He+sIKvIXSgspo7ZWDm3lhAeeN6IW7s3eyHitm5YyyA0o6GzeJZE2
CVAeFE7cJJBxznUAHZ1ir4RhYVC8zSLcQbTQpYL/juzqk2mAqK+s4BlFg66efmYT
cibodZkWBHCpKnICf9POXNrdVKtFtfA/qkLsslSif2/ki5AWA5I2U00qi0wu+tiU
LKNeoK9ID8L7U5TrQuOem0tUiYUnYvRAfS6veUVjRlLnDijYh0osfFyMXom1h66z
Yzk/Ie+ZExZgxLzapg2AMoVNgXN/c8sXdq1DS0ggnY2QrWBjDJ5b5g0lrNq01rKd
zfWeJJXQQ4sZtADs5qJpFpdgDixkxqDeI88df5FLgYOv/hpDYkmLuBF+qMq/GF0B
0ynPMt9b2rcygKDu9ObF8JU1vX/R7favlNuSnGmEn6bujU9nT0ghvACrXh2Xykvu
Tr/SF0MfV++++8aYtP+lCoB1XibSaA8LJ2HKHfDqVQn3VMRIeIRv+D+4C1O8ZUUF
W150VodYODxDfi/mi3E8Xr3+UMdpyRvbo6uEEkKOCFRdPGd9B3XMZ13Vv9BS4JT2
MYK0RmSbb0aaKDeAvsPQ7kFfQ8iU/Sq434gMq5FtI9f3dCXsuYSm1BhVIRNop60h
0RveLFkyrxx22GM9ENM4r5vcquFTmYxTWfExiEi4TkkAvSLOia2vmSoLPDv8Q/hq
x1Jjl4G6SX7Pjs4jBPHzeJbsr5uSekGQjc1jZXw0mV3xn/Z5XTph9k2WL7AxjLuh
lSwJIruiEchyMK+uGe1LIWJHnBb9NOI6Rp7rfisipL7mEQtMeHvTVoZkmBjlwftM
4rzQRszyFyJKteg4CODw916Kc3T0Q1YKmNMuqfWgEPsPap7MH6Epla/SHxX5h5Jw
0DjxdTI7d4z4tJVTQeRPcRDBUAloGBS9OGngctSet6ruaxVbBL2yEQva/lFKWvLn
KEM0BrAboOq6NbJY1icaocHjDeApyWZ9JM0sr6FcnSHGPLWpWdxwoHvuXsVTYUta
wiUU1QjHBtjJYwq36qTfmQe6LLau6umUkU6dIRIJ9J7gucfCxhhfw+kY2BjXHOlm
GJafR41Zi7FoBduQfN3of7tn5J7sTRtgRk4ZKCZ2vMnDJpVVvfnGKnz1QVJRNFc1
9rvp7wFUDg9l5sR26cgvEag3dStAYtsJgRnvhHOoNHvxKLjI42t0Atg4ZfCXN2k9
sFPyHYneyw6dl7C+n3CX1oDzEkG0a9+asCzXz1m70jZHGHVFMjvTqCTlapgeM1nm
o0gvVRQEGeCEv21IzXahn8rkX9YUYoygRtBYs5/gVnIQTGAlh0+VAK6GRAfDuox4
wRfgf8GsCBdaRyY8DbHjDSkTdQ7cxY3dKuT2EDZfqQu3qGaj6tXfm1S7cpTNkbSO
vg9aSdc1KU0+GT5NhupJPA/29r4c8bht8sQDMntLz38M7lLmJcFg1AaiPyEZ9LL3
bZYwHrE6RCB4l9cKRM8NsPGIbjpRAOzn7IlGtRH8s+xOpYlnJ9InBoxJGb9nKVD4
0QjUs4HxbqYhBmfKtE+q4WRIT3Glr1NZV5HGOXcnQ9s5xUB4h5N4XXnAvBx7RP1P
yLbX937XU0BSyNpTpwETZIcNmOfJ5mZgM4k33bzRi2OmNx28ef+yy6sZKmi6KkEO
g3tHzGKUY7KKhiioUB4jOIcBPArOkHZOoqsNsVxscitJJ+eahH+iip+Pp23AUfus
Pb66g/f1dO2MM4JqW+W+hdVxYxjApceV9SQQ5UrSHf4p8G00ZvZyO1xA80/LMc7W
aH7g/5w6KDok5shzY6LcvDSrrmavnyjxX0nzFSQcjPlx+ge63dZqwMg1TI0F9MB0
ct6MZOGtzUmOTu+yX4kGBcfPGvMBetZjNq3uXyG5eKuhPKCx9F0XKAVKaUh2czrT
ChRc1GtEmhz9RrXqDgYiz3lR/dtPZy8yar7KUaV/nLK7u0SLQKqpc8Xm7ocQCWh6
2f8ycpF9ApJEEJ03CwB2WK7XwyyDc3Hrr0hvJjd/+exIihVVlLZJumk2mr64j5LC
7Kf2X1mzAqM69dUJ8NQ4IWwt6sPUrpdYUFOFyhDmmct1f+9E9u3f3vYUx5QqYq/9
XLxI0zi0lmXOdBkEpbO2naEPrHCrtB6HVqVR7T/SejUMqu/QxMIBpc8Y9B/fbUfw
ztbi8eCXH6qXrzAVTYYVL3Ln/S78HEaJE+I2v1GFJZr93+nu1SIqdOkHOJxOvLmX
Inzo5aGddW9Gg1m4MRe4U0RBk5Up8kVEoB1SmzF49h+U0NcffZCZwkjgAbwtOLpZ
UrNXm8d+Q8RqmQcqAbtBfP6OO72bs6LuBoRwtgkrA2BfG5Aa2nylkufhLI9kfV50
+er/rkAWjCfaLjFCma9cdHXkt+JrmkqwxCHgyO+cZUvjxssJjrQuq0B6TE8z9y8n
KzME7aqgTG3UU/WTZ9x3BWt6eiDGiOlJChMTnp18NJjpZK0pm2BR+ETP8cDINlmt
mcjMrMM5rO/Jq5E1xhBDz1SWhXkYD/cbWoh/Zc4h/mibUZZx01GkcoOgN9467z3f
QKTK2DdBK/WMeODnwBP8ldSDlwpB+6JBLeT/3sjmMfWa9CILB3bPHKUoL13ydfJj
eYaZzjo5rUFSN6bc6rHbvJRSuS/Fmvs3l9z+8UwKD23JrbdZVojUZYtIbk4X+Le7
q711RLxfipT/bFj0Hb8pdwktlPmhpdRTMtVuULBnbXh2P4dl+ls4bpAG+zLT4WQG
gl//1PfhqoN2/AGPPS9AkUU/MzoWBbAq7CAPJjRO8pTXXX95d9LfBMGGo939MiqD
x5fsC+e5D6RYbuNnE6tFAEErNt9wWmuOEc1sbNsPj1UVEB1Mq20zb8vC/4mzemJY
2hPfutWRSnkfyoqPDtEOGK499pzZW98XwV/pJOg7iMAZjJlv5K4vULtA8c8yB8Sw
iMbIjUIlFp7N38H9JKdP4QzTqcE+PAsx6eq4S1xKwOlMFch+v9Zk4JsqpfSldSLM
djtpKrPDBkpGKfOXWYdL98gtJ/ZHV+oT5Wkt6Zl6sYHgNw4aYLeMB3QQe/F+xGDQ
VEYNyieo8G04spKKxOVR0zbgVMFLzfMiV+oH+ZCVilLtw4BuLR2enCxkJplxDTfO
bX1ZC8/PDBygv58vZt1FDWNHiRcdQjT7yuYDqZ6SnVMtXl48TUMzSxFoUbav4r7j
YE2YvwVw+Ratoy5udvAlN2Q5fEQGYOeBTkIFi+zE6MEzbrvGbXozceSm/Sfx4rgh
yU0i8Hy+tDOKvHfyS8ruyDTDdckIlt9j0WZgYpeOpVsW0/kNUgrMH3F0JuymQ+TK
A6pzaGk7pwowCKe0qpw6wU9Zf2SG0QEoci4A8Os9YU8kZLyE/MGR0qlN7YhqzPhQ
bDC9LkG0CVnk6qZAuw7F5njk2G7KA4cHKhAZ57CUA+hR5jMH7AluPlB/H6bZ+QCx
QQrqie+Npy7VFSK39+8Ic3TaTYid8w0rydIaT8IBDxppqRAwXDODkTMyqZUuy8d8
4wVclKLodeM0mH4TCYOU3/p94+RkF9yTPF4bLokDr6FoUeOFy3EFvpZNn9WXG+It
/pEQFG2TadqvvxXugZgePtD3WbLPWQkzF5HwrGQ3Rz/+fzWUkcpdRkpokPz4tuqQ
r9nNJP0nQC+Gk7R8fPEh9VQmMByqUx/qu2LgIUFVG/JmwkVUchsAbpAdH09vmthC
x2tHgjEsM5crvcrF2EYR9uVU3q12mi2NDx8C2mf8+dqNJBeUjyO2tKFWX/dQLWaz
YqZqbo2nlagJWuO0xaXgPSLMlk8jjY97DXmS2M+q+cexTDYnFHcbRUD4sUTB1/+V
juHDxdT5Xnco8/5juusmUCUIkgjFG5n/9jXZpy8C9DTTV0Mlr7oKm4tmZEb4eNJV
QCfbkOzDeOjv5I+kDrcmgW6SRedgfdks5HXqC4sKSBTVxxZ/KkSYgqSrx3YxHsM+
dM0ClKD52ilw5yy4We9TIYt1rTHH1VyWS15bKR04EdYTua9MWgKJH3kxW7oZgtU4
a8tjJHlMoTniVMP6GX33Tk3zHMD9/Yx+kHD3dXGvGqeGh1d7Lh841OutdZ5ijwmk
8xbOm3IjEJSrqDSCBh77ATdtkwp4RCyh86IJo1dpm8MBK2+BFeO978OawH9X2Lp8
z+WWtzgKE5bDSU88X2PNufx2njCGHvZRj4rLcNo4jpIGtwIQAb+x83AolRv6r3K3
9DsDDt6tdpr3spu7Bss0dspj5ca2GS5AGt0fXvlZeD18SqxcdRv5kfw1V9F6nwxz
KiXSim7oEzNp0xFQPjogx/NQCSSn10kRqAOKJZWJyjKAPBoFrvMLinoGUXdB7Ag/
7XuUeyjnjxOWQlQkVsJLTwkBRVt8OCnvKYPmYdJvAt113Dcj/VAWp5+ua3R+o1Xc
urga61+SKBQXTaZvJXVyk6LdDqY/TNjNHglvB6qdf2um3Ss8AYiH5K7jpFpYunqE
7hvi5uNO3mf5KLGyc0dVN57MDGmoWQtkOQiqO51eCZsuJC30x+4RIr8LMJx5hPCq
0CPqxdMZIomaQ84f8DEYb01HqxHsGRCHGQtITTnUrR9ETaFPd0G+5cQ80T3tMp//
KYOUbpVLLwHNuE84EF1FnHaFTG6BTRf9/QsLOl5NnKFcG8cSHXyKo9oKXIWPY2yK
K6kQxS3IbxfFokxI2utIQmuPaDQB1vf4WIRaagZnaIjkahodhz94frQ1ag4wAE8L
Xw3UARvON8wAx8zwkOcVJJDWZEUhQsXtw9UxMOyBV22cqfuHteWLLJ7jWLsDT8oE
Mts7gBbP/8kGL9Qj9Ujgh6sSHPrriQUkIfsrYosojOGUAuHzFz87u9b0t7mHr+8K
I/88zAiotnnmmB9+EERBoV/QOXQLnovfrGs0krGBdZMCt2g9psiHOAAxl5ZjOGRM
YuVIR95ouHmXAqy87Vs5271memDdbkyUbV86LqmiE6rdvfUSKNBSnmmGc3lFtCne
Xw+BUPBoE9ejTGaB/MGEygDJwswOQOBd6jl/gpQ8xBJO74XmTQgys+Yxv2QXzEpk
bDlP242VmWy9QQFCYoISZrQJXQtBwKQMi0xq3NBnQIGEhUuM6oSl3+14lr4NyY5q
bni0JLs+fF1W6YEIr3bO+hgbAozpew1Fmm2THTc/5cnliJNx1QOFvlC9GzpocR7e
UhOQkZLf2oJBhvkJy10FUW4omu6oE1gVupxnhh6pDOkmJZNbF2pytTPEOeiRJzmx
5d+1Pqh9B3rFsPmiKYsOjKYNsOienTTTB5PuLQIC3iXXd+OdPUJelAAPVkPm9elg
FYXCuCsq3a7p1wESZrT0lAW7W105doG3f2TfOhTo84tlB8xsWKSRZtXztX36b0yG
IXNEqGuf9R+o6sqoSJZiCgAYBYMYTANQVlUkYC4wERqdCqszh5AqOdgJsW9N+OH2
lUhhmor6cckRJeRJBNjzDiDMKUyT8EYtGznPOWoWLGO0X6J0fM0dDK87W9i/ehFv
AIGgCLFR4+ddQ+M1fl9fefKuZtNXAFAgMdPazH5LpUPhCiAf9MQGjVV3uwgZMrd3
hD4Ykk4c8vW/eyvrCqL5Pz+nxznKive/oh49vBNRY9+LhIMzFt64RtemxKYBvQ50
urPMZzgPlaTIzq5d2gcpxjYbOVpO+v7OSI72Lcf/ipwXP2lyJt6kLF0QSX3PIoQU
DIzrvGZNbBJPgPDJxw3i5q5HPDUc8/Le2Y66STNsbABiExWZdLLeAp7byLQYOcwW
JyLgTOw8/D4V8S2wz3ygUR+PgAFjor9oEMYTkTmR3eZ3bY5pMEwfg6yXUlyvBxPk
HU20x77Q2vVZfV/8AnZIHd3LsqAvmQlFmpkIkAKrkEpQwP30OpJBvpdIACgweXjH
JqFvEFZBu//Es55C8YDbZovlBGftoNgdP6DFEMa1GShdYIBvCVf3Q/SOhhf9pemI
InmuVJ4f5O3PRXGv9tYhF3ggMYpgBWXbGjPhtFoiR8LqCgMiQjw5og7ylflBXF1e
DjOa5RqcaKWQBYbaP2Pd+xWn3iNA440mgYq4HEUwm36rUuq6/NkYUhsRUqiuuiQm
5S3pKiR6C2F87s6YkAql/vYcywCGa0Xcyhqk5rt5tfUyPPn+Fl7EsQ8T21mGeoEC
aOgL+ALz8na9n8wjpLmiuXKrHkfhGCxBQggggwfT1S0E+/bbGonpcbXi/VidbtKL
VBhLVrg0Tw3r4mfIkG47N4dyNGQVl5jNPnf5R2tO71f6FqCZbuPRCVSd9OkqfEer
ag3XO1MqPlFN1WTFu2Tm8tN8/zqFsoQ/4eFLbQ7AMhFkfRA6vWAkGCUI/bhhoAnK
TxrdRj3JfnazcJmLL3v9Ra/KU+/UJ3Q9badouE6vaYABz00czqmIW++hQCMP6A6m
s4O00MhG5Chx8v5X/IBTOZByGtaCiaCPYf02n4wetYnkE/woTem9KghRXQxvd3ng
Zplo5/388s08ryZ+ley9jP4dUGiYWI9XEehuqDrgMmTK1V10SZQGLpHXiKJ9bRPZ
KSbAnofMZYhw4Ar0dE7JhNxuvj9RWLn2ToXwCpRqAUEiKX751NxRA2OY4TAdsINX
VGCcmxUOPmAzwR/Vr1qmAVcPmA8bAkcYH5Poj5T9R+VosoJ5zSiOwk5KZc2BKFmc
K2aokCUxB/T+gLVT/2LQ0AuuLBMHA4DA89Rde1HXv4zvCGX3oKfXNdjYi9S7tUhL
WX+kvYhuFgZzwgDGMnZXkOD621S4+f53pnC3HAZyEl6PGEpJfMq7eSmPRC+SIvi4
ATaHoEMpA1ZXfApaZS5ZibTk+esVC7HJ66rdERLISx+2fhBn6bR0Xb7g5yTRw7Zk
LPQjwUFnjyaAGbuEVM8gar1TrQ8HlxY/Zrybe1XbLdVDkRIVeoVHS1t8CDANHj/P
6i9HPRZhFQ1EfHuHE0pG4xi9Uza+VvumZGYsYHGyXSA0jUvitUTA2Qb1oXzPZijd
5WWpvRkdiv55qqBnkwYTpdYoVXkOZsF1xuop3NEMZ5DJH0nu21WXSiLWydxmfuXG
GD57ij5FPnIz4COjhAsQ9xiOqq2vADzDIQY3fBvwI/xoRHg+g3G6sAPVsnOy65ZZ
n7V+d1neMnSImd+qnVFRPtcZcO/1YBnswTK0KGDAj2NJhQG3ge+pdyxlwO/kGBHI
MU38THMmPDCF/COZaC54RjF+qJFHsZupZghlP2XY/N7TNMPd7qUZsEeY60p9Vuzo
nMFQ6Saj9Q9TFNetRj8w377wCIiYNBhpj+MS0tz7AqwBkx4SPirDgmZw6Z2mzdaP
w2ODK+0mznBaV7BanpOvzgPvdezXUCNe+lXCckYsL+br9yF5HwnX+wwavWkcjvgL
98Yf8GOihpqF5dRrVNpFFGlGOmTw6qROrbiJMep9xKR1bLr4n21TAeLV83dND77p
fOjWixvrK2xB8GYyFQhnCRL5mgoOuJtTxArEWfVU9sy4bZOcGqjT8KHGvl3TWb5G
s9KkX6T2raeMJh5PNbQ0/CvJ2MBrQrFxDfZEevDNRsDzTHZJzD46s/1UrI2340pn
0Mkkcy7WJvsUIx5E8nm+NnP8DjyuBoTdvHWx4wR7tobf5TiO6oQFHA2dlnmCrZsa
EE8OpA3kdj5AIO/cBpyt6TNRrFHn3aGg1OE38Yyc+aBtEvC07lkaukqceocGTRmp
8/bq1aTz7yaMNdyd6e44rPuQJfcCdL+auv2L+qUKnx/pVuBIDt0lrV4ujYdzHAWD
YFf/ghPmG+zLMS9q1HxAe+i/UD/FgfhfBYMEGWdFOqM7Y3w9Y7oTyR2cWUGvAS6c
t08FbSsvX9Tb8zLZBb39NclXq8IZpVzN5Ez4/D+Fj6ZxqJKYrkTe/O7Bd5cThrYh
BZS9iHbVm8hXcuMmRlvU2/ZKc8B0Gu0aJW6fLYxBjhuOLcH9w1dz80i6qrmHXMI7
EX017C+PXXEpg5LUSQKHuZGGIyRRkS1nOd8I4OTSafqz/zYTn93b6LZnXb+lkL1d
l1Qus8UnTMKF/N56e19tApWX/F27VTKw1VI728Pp6PMyiznMpANteQTK/gzBPBuR
A4S6y+xyCq5sdQsdADKOs9AW+z2JIQUdZFOeGFELW7FavSjA8Aatp3d3WiVf9ab9
KLQsUy3+vQlCn6iiL70nGS0d+YPFfNVJMllDvfuZ5hUVGU6KkY6t1bFU1sZ8VuYu
RhW30NvGhb7uNf6cTLegGBikcNregTo6bTWfIs3vlktUFgwFJZlSxz2e2D6AA0dr
PEN55SbrNxqxlV+ZlJ6usjUm+1NPhZsXRTUzH8qoJvXfCPRvWOhkssP454sJtnmp
u1HeH2jHvfS7QFLBX6SBWHLXiBkJDx/AYkrZy9JI5ZbptONAbUE3Q5Bde0hsN5zv
gvnCHxixThoTRwWu3xj+sETRPyjop4mpHjYq4kUbf6BgIMwvTM6p1AduJd6ajG9Z
le6gHbDTlWvEEF0xdrHWvKMj/f3KPnIPwZ6GpBxuwvdLPE5o1gTOKVgKWCpQuvlZ
G9qZoqkIGHlht0OktSG+1SeAkZ9yH9oXpnEaco/WQE0wjr6cIgc3BSfLKErQ5rLT
wVVsfJsFK7kV+v75Dk/LLZbf07knluueIa2Vqs6NS6ueMMYgh1rAomyuOL7VvPKw
vErJVnj62eVgZs19XBq4VC9CFeY0REFOKbmhemuJlnscnh36YIr1ncIrFgUlD93E
A4FmK2iYSyF0YLMn1+CwRkbPaEJH/KnNC8r/qxHH329Un9fkUtHFI7y42S/rMJ1+
rjDpmBmaanLKA0J+Wk1zwTj0324d51pFfrCHz7dQ+dDGfZmSQqtnIZlprCc2ASpo
783taa+ze7ryXl1od7eLtvl+4aQGspRfqyii8IdyctQKGWqWXME3t2w9xGKfPW8e
3/3lAA0Tsx6bMaSAY5Kj4cQDzR9rjrHjA/amgfStF4vLY9aSzK6qvyQ19R94jXK2
5TB8cc9jL75/O8inDz8G0EcO3gyhSE2zB8JYrY4m+bViMeLfwlXsNJDdgPvKxptw
7hd7JpzQJOHqNcfdk8kytDtYgT5pUJFQ/0eRwnkbz3fqxCI4C46AKa5G9yp2w60D
iqhhIZ7Nfa0/YBooOPiKvlczxp9HwgTRoRf4WSkygASz3bzcJ64IMPsmb0R0Pkro
BxGVO7rBPTN6Rk4+5Np8ij1ycfzjRQ5a+Q2kzAcLfFNLwBkxGuj/IiuYaCvm/R9q
TdI5lkqq/gf1+2jJDkJ18N4FdxEoLAGIsbMxwDt/49s3NIgCD0a0dGMyoTHgUSg0
z2q9z4Sgz0YOs8wNDFWF4xM+j4OEaN/3NqnEMYg9S40xhLg242K+AYLpF2547lMs
ILDHNXrFrN89aoJpVdlcvVRG/RTb5DX7VyBa0ZEmC+D2v+B5w35u/ZK+i0td6tgn
9a9XA14VAVOTugfdHjryhnrneW75gjCqamt2HdktdUlLfUsAU/+peg8oY2OBUTDs
jxlgs+0p1B80EsRsid/NGP+fbVsco/DA4dFmPzC0FUJ3mioEAi2yBgSOqxFcqCtH
eTy0FwlyyW5kRAzGvvdABivCT+pX9Z0vh8lFiQrJ1I8+XHuUEyzMi9WOzZ8XYUWl
FJ2NuQ0V73dQCe1Ni4qebGCs+sCVhPhaavx8wPWvdruqrjVX+A5vzI7DKY+35jgV
ph6tQVss6ipmJf+0c1ANdeYVIy0xvTgbYRNBKzhJaWhza3sAdf+OWpdg5a1NOWXF
tAue8DHpJ+7TMpxXW5ykJedaKVfN8NOqrc6H+zOgw7MMutXhwdB+hw1R1J1YsX+J
B/2401SdeIcViThRRGEyiMIawwF+K2ihJvT+S/fMM2X4CUEpDWDvX8fo4u+wDNqA
kXQB9DVVI1a0JtYDGVqwpQSlW8i7bFZL+htHhXK7TZe2lmReT0SrxItSWvxhpxs7
+gI0XHDKvldoFHNTz9VQO9zBHrS50Be0k4pOnmAw554NCmeg66AlVS/tpIP3/1cU
H4as88IgQcmvP+oxiIm7DbcC3mjww6PcjaB7cx0HekINWV2YyUQ5WuhiHnhfwBJu
0q8jdl92XpikulfyVwVGpJyx/VEzCrMDbghiWAK9455oPaaW5Mni6LlYZ19eS9fO
inWkDXQJMiQ7tV7/QT7MYYrXwlrRbASPIojiVQkQaZKtGfI7w/bDwZMgq+gGF3aT
HEtfAd3BIjdtljWbyAcS41DzPHtiLTHZTiZ9jbtqy9JYz1xSE2INFgICpWIrce5g
itnE+9jKEjzPUpugdhQI+4QJAe5WdWsMYLtpliabjqYc554kvoS3Bjr0Xe//2Icn
8jdjKQX2dxfOwBHR3+7Fn4KUWCM7+pzvg5dTIN72SanGrbhy+ztrm+PHPXo+Sia1
jSnRr2xPgvhXfKk3bwgZDNWymGCXMVgYBX2872+SVfC95VwZIEKItjkalUyr9fST
7kWQsAj6HudGQ7RV+arYTIj7w2yjcM9DlvOIZXwEWIr5dE0CYBIl8Xc9FH1wG9Pn
vjHvNomKpLiMsjvMCc4i+kpUUvvQ+IPoy9U2l+Y+cLRI2uYQBF+qRHrReiBhGtDI
yqBegHKCoeVTBSWXGYB/1l99sicvdHA6wDUM+Fm+D1Cm4DFBSeogscSgAQud6BF7
WFzqGsPqW55vUhz9Kc/yk9XHBrJbZPKtA26KJWboPGJvo+mp2Z5os2YhVGao52Nu
Sd1knm0Z4iNoY5G1jPQbFPxSXbRWNzFNm7dNT0K2LEKZRat+EBumzhTmyVRZEDMr
LAu2WvW9qxDVA01x5sS97e/rDdSiElwHctumQF4R4cnGRaZlMpw1WNuV5aR9lsxK
L7e/8b9LqtIblZHxpSTrHTucYOvCfBH5blCLY1e3jk9vGuMMXWm/1JX5+9OS1vbF
90yxBBFfSDhAlUjVsgUmg5q51yjltNl06FfZYegxwvOyPMrupBW0mXnnI6uqRgMq
kaJysIBej42mV6rnIHYir5TX3VS9KH1zfFr/tL4WwrAodGX1Ms0xDF6lxkJV2BNo
LlMcFIfb28CjLd2yto7D6afOqhAcVnQGeX4fnmsRwtlA3xz2Ic/yS7aFGBtYlXkE
DHExPXFoabHHiqbw3kF6PCLFvfb3nwKKjRKqV24qlgUCeS8R0HDNh9n7RKSZz0eT
tuKNsMGCZkAol3yzfmlcvA2vLo94hnrmWzS7DEFcTPub+0dQZnwinyAEwXS0UBzP
L0JBOl433xMjuyS1WcFhgYOuoIYABoywGT9WVOhnDPM0Uy1XekCfQQ+jp0VFLlIt
LAcxEyb6emAyHAoXMvJ+QRll91EszWb/UUXk3JeyUtzKKRSv+NUlk2L6AV+gqa4x
uGUQCRIJGNExI0ZN2pKLV5tyVaMw+qhYZbm9iHKQIlD2kjUHoLMTI5QS2P0eUk8G
OUt3pEy3uUBDm55DsOJjWJGaIjDQCc1YNrLEVAc3h98zmX7MxvoswowJD1B5Ps16
k7bMktED8PL+O5fyF0T09GHlZ2qpTwkv8ZPioG08c6x8zS3SXkCQtdvzh6qr4R49
eC/LKPXhUQzHE384MA2GlcNKOD+HFYr+DEO2vX3TmnarEW4kbeB++cipiKB/Cu23
+6l1cHjqh7rgyCt8p/7lajtM6Nz7PAsn90JBMzSH5VKpcam42bCvGzRkkYcUNSu+
DyJzCtcAbKZ2vvSerHAtgLE8CiuNullY2ZmYGv2CM+gZp3hVdR2+9QULSQm/392Y
zuym1uvSXFodU92NjhI6OC/ilbIawLhhsRmvzbUoiEQEfgpghPoItziJObwbO53s
kEvK+PxF7jSUs41/j+iTSOsnRq3nqhBL6XTy1khsqi8mesQEHIGkLk2WbpUfrnIw
/bagUzJyi3QBJQFSGfzt3PaxZ2pKdN3GuhWIUI5GBFmiB999/fk0682t3tbPV1ji
VkOOBtU+a1ljByOhIk9EZd2pY+o6YZLlct197+bcOTDgD+IYiugKtHFpb0DqC7mT
kWk21blTvsLm3VZzUDhPCfRJD3QYpWfPfsIpj59IiSu3uvKb1QM7TCjMnivtdgv7
ChdqvcFys7xbTLUd0JP7cqu+zBeKuNqdswfZRMWCYqn7ESB+jLz21SowQT0SsswD
HbrclwNxdl1MJzSqivw5zRw3h4PY4n3EyrkI0Yl/JJDi2xOB+io6XxNDP04mTecZ
SNsOkWq6W3YtbR4y66GT04ozuIGbTZTeIKdihPRg7bVan5H6oZw+edyjJIB3h9fz
oTUOV6B/BO+PV02PsYYK11QepcVVb+MhDkw7EePVJ/GPr4gR1a0fxB63d5ec/tsr
INgLxFAhIWDG2Rgna+ulVL2fCPgx0g7wobLnlSxjR6tWWktnXNWd4j05mfWORwih
35iP07+RXSDdpoP78HYoR1G6TdIwz6BzWiKnhecCBYjJYuoF1Hv5gOqy92MAFpWp
H8XMxp9rHeflg3Bj3QYPiI4p55m96a98vj2se2fKHWInyhxC+JXISy4yfR+0cpEj
qoF2bqrLV6l2SLA/kotsDOmnRGS3kEW0p4MAzyNKf0z0XphhawbERMoxUyowE2C/
P6hH5ZA/2XNCp3ZdFkSFDnf2e4PaByxb9tY/0NGfqWxhZmdgqg42MDakPeLvX1kq
UUziLZcOehWyNfBbvKmB1Zuhifu2sqotWhyySv35CbXv6uyo79mjMhf+6xTpupMd
Qk0GEWda8VTMpu8sIcvRmWB1IwJS+9pVxiiFJRfJfMWr3+rIyOL6/FrkHlC9WzkQ
HI6m1sd88HNouP5L2GdBHKwyGW+Vvmkwqd/CmK2AbR5gww/UOciqKJ8t1xiVczPI
bMTd+EOPc0yUvHEcm38qto/AYm+kYpbtokYQI5QdmARHBZTE4K8Bq3l2CAetIRgC
7ITt7+Xd8BxOD+8jytE0+4MfVXpbXMQpBhKa57yh4VcaedrH1BFfvTkSh160Px5j
NBiwfmH1Hp7W6UTK/HoYidPfKHLetEkZ9gYN62lFWyAHxn6HrZ4HEzIhRpxRVEDw
sx6P6CnzVuWDTke17cAivz6nGeUOVhQQg7Cjw5HDaK4ikwT1uNxRdlejydaj4pQV
JikP73HU8a66QClp97S8qTeNi8kfPqEb6NiMqu0c4b6I+lN57wGssMagtgvHfRLt
0fd5OFU1exthUPSWIV0ThgPsqwiFqCdc7JZk1grB0jr6XXf+9LF3hSAxG78jyj7O
UrZ4X+kFxRheHYosYYEDZYiOQfkmA8YMW/Smq9MDIpSlX6KluemeixPJIcdj5UEg
zAkAhdtKQfOKE7xsdCf6dDdpjZG55YHCzw2ccpk4ixpYGtPlkXHFTvetnC0haizu
+QbPbtTOFkcOBZ2Fju3GImmvJ8PH7GwQK0F4epZ/XRBJq7mb84nTFcPFo5ZDyZwr
JwvCpnDM3cR0T9I/hsCNSDUYApMsNzWnC2YK2IRmQb8Z4bObgdEEd93FwY2CTGKD
eV1rF9Mjrm7bcDzeHe6MWC+u95ESIKCDYMYqnbCHVUCRirJICbFWdrSqrjf8vjl+
FaisE9gicXN3FAnOsGRgxSHKFOb6DkMGZN8psKJFANHDLZ/mjiKd2+U8iO6Ojf8B
+cOM8Vdlfeqi8lUdUH5gzcDBZ0/zpv+33uEQJI1JRKL7jFZhHbD8NSGn7r9BHjg/
ELLNIajlxOmSUyqpY3UpxE7jURtuL7GkFcJH8hsAhPmeShNutll8cZUEaUlxuWZU
wCizxZN/CljHKppWutyAa08vJMGZrdRoZ2hBZAAfuda1lZ2ZGEhQfDN2pArw8S3H
H+1cfY8Bn9E2lT3QwNfxKA5nqPpJAbRg4vTO1+lSyWU+Vtwq4DNuRACNryPjf/05
+PFpkoo3EOqm9sRrYWTcpLmYWX2pu6GUJNXRRvd6NzwkUqFPkf4bsfS7Cl1UJWnn
fMQEv7+6qWU0hrTblOtW5N0wkY5WqkTSGzVl4dvRkIDjFZz20W6jMrk0wxSDPF6d
PltcRB0+VQ0Rj2gt6nuMh+5i6OpR5kbBaG5DE7Fng4Oha2MDmYstYV7yND9oBADt
ze2DSjHiudHxvRtfITQcYnnn3z5HzW3QDuC6BydfJ4OJY6B2GQmo5tBNYWKW8Xya
et8epAahp1QGqYKviMSk3MUmGPqTFLppB6WSc24EImPqo589edszA3Iunmww6DQ8
ZydXPy7WV5YHZoAL6xQpUMyUsUdFAQPjNGTJpT6VPg8D0YH6KAA8goRQXCd9BF9g
jf5RF+pDL0rll9tCe2B7vRnObzFMXX0g9VErRIPk98UZRY8UutBDGnkzlkhCtO3C
4bEt2u+zYdOGQZHi5czotdi155axkcXCL/bPzh0XDefxB5zmV990jAez3IFMoh8N
40e7afjK6QVJeSGya8I+gNEERYkt60ZO9dVoQdiOK4vt45WVEIND087KzKDmXtKg
+lxDPckBOYqzwVLraseo2r2gy9RIOvBOaeVBDv9ODyuZvPAIGwRBE/rh/c1nQBNG
4kr2UpKDcY8DQoTETW1bA5okFszfUPzYOX/C1xWhy8fDubIB0KbS/VLzcsmCzSll
6AAct6AUrdHKM7wu8EYRzyPHelQYYArpIzijkEMju3Fp/HfEcIQoo7U1cGF0EGv+
m/m2NJOPlDXDK6Nej2pFKS7hMSwKxf7hdd9qRySn419TmAphRGZeRsh8m9x4u1Oq
4YrOelX8Ih8SLeGMAspIKqT8wuW27vt8JVSJs4QTTNG6wY1kPFJTKk+4XMcb/WFj
qaZBb9U7x8XKcmGGFBcSK+H+j+qSI6JrC3jw99JjVtNtyXWNKnUywcKbNATsfseo
it8j2LC+htS2ttdGmqwM5g6ZRWUqN8vkb+kBtx29sa/QIYcW6fhZl33smvMPyFiL
0EKXI58diUGsze66p2BsxJAI3/nNgh0VeFxis4OEzNTTCgfTifDroFbRFexBeif0
uL5kDzZ1IIwIILtunkI7H2pKk1W1skzxXe+DNmGUbF46xRqgOONCKEt6mWaGq4kl
fpTAsR6N8q92YBfDbeY0Krx8Ul5kKum5jlW9Ir2EXudH2Q3tC9LlIZGFikRPLQ+n
FMrPiOjuobOnPasR9W7a5q89qBUq10VQZrPli68LIxlr0ksGnzoQvutg0JS5ZWgo
NtffMeabW+J4Iq8ABh4ioFUmjohliVlo2dEKi8L442d1D1GO0V5Cw9sv9mYPqHsR
TBnssHBDqwKNWwmIt5FS6wcAIwQ9FWBZmgjRKdwUHYsChyMOs7M0VNGDdVS70xwA
GM9SvybX20sz+pKMWy8hJpTa0dYo8U3SKzYtIfb8Z76YYXHi1oBW2HEQMRlbjid1
rvx0Md5H7WfmUKwPi4TgFm+tmE4cPgcL3ZLiBpgSJbrbN7fw9kmhrKfUvIdkyYx0
gxQelLOHl2vMWNnCnX8+FdMPCKLeV/Rt/EPMhDlcE/0hawnsZlaFmAKvCubJItiN
dZWf3XrbA6CqADH4YUkTe3LdeoM8k6uP6kb4OYJL9TPiZ7XtW1BWlc+2mixPTltS
NqvWUAR1Dsp1MKd+LvMuItQ6I2LcUZr+sF3c2nMo8U/vwlvgySRcM+fVvPDHj1/d
+tug3FFszcn6p4HEc5lPaXTBaWZLnbHXTQZQKJP8cKZ5RUbQfQI6omHjUzL1jGra
dzGMjzM3yllRoQdZMcHHCwZifliOP/ktuxu2r5wckuUBOd6AKk9icu9PrHSugzSO
HtxkWvN6m38vEOQS6WjJXnvAzJE/72QGkXHEKPH1X1YuXbDkpvJwVrM7fI/QNcqX
GqKpgoHdYOmrBzRPf25uzUWaKN62O/GGKwQWzMCYdssjVVigxhuZIKr+bMUt3j5o
Lio7ruaerFCi4jcqJwySf76XWS+kYeZ5NVfTK+Cy5kOb7yOvfkFPFmV0SPus4mJS
2chfyUGhEQTUfU3m5bxTEdXhjwzH7706yinGbrS0GGctpuojb6Cz26CZGANDPPIe
k3cr579Z6iQXfj79VloVrBxrCSb70FhEkRf2VEiX3lFjHqfevrHh+V+0ZLa1SZOb
OCykV5uPsz6dmNQho5O100jEEkZvWUy1/gQv3BO9iGGx1YmtIcQC/0hgB8AZJMHS
C6zpwCSm9g4lyhZ9sjQBw/r6YxZUR34G7gI+ifjpPkqKBiTGoS+IPej9/Uf3uPJC
Ydu7TVKqP//wPCsef5beiz4uvPSU3sbIZH2DISXXcl3wl85q2HYSAsqgZ/2g+fru
v2UdTRCEUsFaLbo0xcJSraLGwxJekecXez18k26fTygrj6tbO/JOhsTDO75rXP4L
y2EF5l140AcLxr8ia19EBcVDS1A11WpNykVBniojLLkmcLly7mn4fb0XznK7h4qt
rNfljbGA/mEzZ2QarzD3jZwpNXm0vI9lQzZTF2WrIv9De4tW2azU46BoH35lDDQa
IXs7oE7o15PgrPDDgbhsx/rNPEK8V48R3m5NrlYK2E+JuCaXEv4/HWSZ7gcmk6QT
VeEWjcQTntAlIuYEDvRp6rIS4lTWWmJs+h4SXizwGn+2FB77lTTbSxljcfl/s0gZ
6weEWppLMDcuvTf9Y0OASHAA7oHxUKr/AkiWRJrJfRoYHMmbAyGEeVFTPxc6KzIF
MhBvixTjLS/OY/VjARbj2kImyO70fETemIyI7SEyjPo5m4Z7Lt77exuEZAfKyeq+
TLY8jFL2/7L3LIPbiOoroBj/nv0gPu50G6oufNOVzKasexS1lygctG9BHgUUMiG8
dKPzHXoVq2PwafxZYYHYpIG8NS/LFIz1zyTl6JfjShLJ3spbhvpjRofPtSTzgWmt
hczGYSnLtvpwTcLHzxvBcaJZzkWSmbi2Go0ZUAWBdv7ZLq1rhLtAZmcTUkERVo5t
tEhb60/xBXJimsGnLNY6tP+hBnFBNhrxl1EmbHQdIyU5KA6QeKetqiKB5DCAHq8h
Z6u2G7GU2jn3sniS11WVFmPdw8QTpt6BthHli3FR9/sXfY6Z3K8++TX3A7uGNJ/c
fMsQMs7+A2v1suyJ1iVbbVePoNDmEh0NCSb2jC4aZT+ctbdO7CmUnxkSfHpMkl+1
Ivw8MRWaPpNPEVnFPTUc5ErbDe5BNcORR31Nw9clNed1a8w88s/K3Ohfzm7CaAOi
UNcbxkftSUM9vjBvuvRRsBOxr1+6lwC0GZmUH4/Y2t86gYK2FAXyZMfSLsODoCx3
w919jA6GuEyQ7VPhthuNLuxmC5ltNVO45i7Fkg9A1o3Iy5HSQB0MBOElO1cJ9s+F
KMDshH7yx0tr9TiPLohBiEUAPCLLfnquYMHZYMDO78AflalPaQYjveZeJe8MJ/E2
V2Qrbct2CHviWe8kIzfK2A9c3ApFk0zFT2Zxgouc8I9CaO86OgmfsH8x/KvXIE3X
aTqM7TFIPP5UXi5N/s+yR58r7R62BK2QDQNtDoZEiUnYk5drGeAptE8SN2V5Gx5u
9nDRhVP3k1S7QsLzLDcHvsPJs1w407O64WFssvIo1UQao5TG1bJT9Eg42W2mnMOx
v81f7iOOrDCluwuH4NntBVLyAGJMZI3vblS77V1PHSsFDmNtSMPDcPyY2b21BWe2
dRLRTax9yDbzq+K4tJ7BKyFUZKZpDJ/ckenWpzrFuQU8hNISSrMbZW7Ufv/yL1kU
6zw8s+klq5x7d+Etb7F9LU8GFsMR1j6MDupTZOm49pL02IOZct3UrH5McfHABVDG
A4tkNdEDacuD8DQP0cZ5grZLdpBL91pZIs4KhTerJPMX9bZIfIsMV1r45rmbkx5/
wb3eaj086yiQducxwjSmiFSoPyh7lk0UBQFLNOJ6tlcragP3bkEExAxcKCnNeC9B
V/CEG3Mk/hJduB+lIHYWkLUst4Hu6hSDl/9A16RLt1gBXuq/FbLcCjCMxSzMuZvD
H1uFlFqOWxgFFVDwvDUihhQCRpekbaqi0D7hMOwHeG44EDA2sBkCG5CEk+IzSIXR
/sTrhfXHV5JOO9QmkpAoGr7AWaki+31mXN8nqE3u/UgS8t2729gUBEjBnEMBkx85
EB8ylJObx0mCE7Rg6NqNkIOZvbVrjPDnvysFw2QjfusXp/jYBSy0g8zqD0CXmYeY
Fz6iuFIvIgpa2vim7zJFOsaoTC9JAAn2cSjKT7WB4N4fq6UEJb6YDW8QExrhCwfz
GGloEXhEAWLbYcGBS81dJFIChLqLw2EvULdXA570Y8MW5dxvtLSwyE/UZ31G0dAE
pZF2ksVvq6n2LOInlZe2i5NpoTa6RLjyIAXfU/7fOtBhq6unOTm5B3+X98i22VxD
IBglCuVSfk0uo/CFws5VFPfFmOur7RckgkqnngN1tCdU1w3MIiILH5ysaEgzmSxw
wwow5V+I74KUp+imOB2EF1vmmLOanEFRDiIeuKcMWQ/L2BaXBtM2pbCXczOq9cF4
iDkjUIVS4molIy/pgIwlkjCa14524qKmX7IZJBFvHbfvCpj8Y3MwyjjPco516hiH
LnvMDwateVZfVLX13GXeJHIQtTkP9TpJPiOyLCNRonFD0ZlcWy/HQcPSlOUUDouM
uLoPdRVH/CLeKW2/s1rEapmE8xSXPho/nFKovQW0FgteJuS4IHjGeNUoW/XR1+uy
LTkOvoqdycPNJ9u2DkqCinztaRDeaTjJQ2lP5/QV7zuU7aecrzAg82Ppf1NFY0bz
CCrVw4WDjP3opL9tKlXZS5qBbimuRbOphYFuXduJVM8Vko/7eoxc7CYZgR5QPaqW
jGnDv2IN4HCtYxT/4OvQRPzndy9EAYKymabCxOn5HhEG1fYWJ4roNZ+V51q49Mq0
Yvj+FRewVt3PEINpKtC+aYjNwdMXzYnJ1UZaV4WmPnGenRAa8XZ/zoTGU2RQzUax
NSxnSse+4lNazxcwQea5+npAkUfIj3Ef4091HwNFl+bXJLj6J7ftIu7QEpuMOwiy
qbRWR21ONOjmva83zm6nKcb+/LiEhHHstJYbIcE4JUBc55f4gYsOjcdfXjDCRgZY
Nybiew8Jf/fsfztYBIPACfFwzE7Do9k32Gc20Fi6kC/gNHz7c95f4pNoe3hGGQIG
YSznbtMGqv8UiEmvj7DGVMzqkcc91KDPsLEikK7g4jehC55h97/S8O3O2jk5lbN7
NUd3K6PgLCmu3pcBA1iACJwdSHdKsHlF2ZCyuRd/tHtSf3qbWSrOcvMVQnSAugA3
NB5AXMXI13WjiIxiKho33KUKBSdY8B3czhN2PHo/8WAVq3R1xGRzHOYWG+Q2Zmfw
gfkmq/yceoRlVqkuCmWdHbmbOcikox/el98thribHcQ0h8SuZGpBfaDfGay4xqPC
IL/HAl7MLpvwjzjs/E7kyPoXr3DwQDL4SzB6QmrZ4fGKw+S0A0yplPKWi8+TYpH2
GNqAKcLm699Wh9ixdqotlsE1yrJv+Brt8Cl3A97HSy/egK/Cih7PeDRfD0tlSdrw
PKUZu+RY/yPxPq00mCd7TOlW1orcdWEmYY767l4f2LvyVRSnjaNLT62Vj7E3IJCI
hrJ7zZIZBpUrtgX0iVsC49JiuJgktyLS8UOyswAoNMLNJ3TejNnisGxqQUN5Tn3V
tZ2SND6WjcHVlgsciyeKsAsee1UcG8+Ysx6pjQAALPcald9YO9iGQVpDFFIUq+t4
FrZhveCHPko1rh6rWVgYIQN6AjJmaT6OFrPzoagZ/OrVOV3XU7BwPdWFQ1AjZnQ+
UW4Kp97ybwoq0I88A647cB8RnPqt1C/Lv7hxr9KK0LWGq0Lc2vULjHlhbYx9YxTg
mu4zMjkVPoSE6tuMnvC1LuWFKSfl+syA3bRWfij/Hkdwy8z2yuSm/NEbkLxo04eE
5y33rY4bx91bjHKTyvW5cfr6/+BGaTchbfTxY/jr36EUr/mX+Sd1yHYu6MLcLD/e
g88K5vz34b85BsKOnJHVvBJX028VjP6zln6ujoPnJSmOJ3jMD+evJ3jwaHyW5YEi
XxF7hXbeqlntZTEt7Qx3Kpgdx1Fn441QBuS11ov0mv12p4fMFcXkxZMwTqAPNGRu
DWkMZ86X/S+Ulhd5zL3G2MudyLKbgJx6S9ICFMI122YIAHW9PJsUBaSRrTzCTsUn
JrfsoHr2VYZXO3sgewAj9DWA3BEfX3aIZhUiBEgL7dnN/tHQOp8NKVVHLfRBDfZH
FVIMgAhv4UjrPzls/bgVvQxeQ3OYMV/sCDElI9HT9ud131QiA+p84HHnLM7CBFDC
WxS9GEAIqp1m9glNBCtj+ycRhuhCLXL6L10GcmfyoyfHM8eH8Nd8xU+CLPqBs1BG
bHdqbpqasz3S5i3v1evh7S4S4nnxoKFIRcE4ndj5hTwcpNfxgywQ9gz+/gWbq2EQ
KnOWiRYxcNry9u9SyjOIVbf3cA3TBAhWMRBD340AvCNkIQqWzwtK7QIBuyxCfyGq
hZ+XqMXTs7TdYjaKNVGfwfoszS6WshFMsiPTgY4wNDttgbStOgktQc/a9XA07aBC
7Vy3AwUifDDXycaBZOvazqKVvoPZeoLxqhIUt8yIryytp1p7NtXd+NxBMA63jD3q
pi80LTFGs3mvcVd4TU8F0lm5VIXPDaaIQCt3t5CuVoM5h2MRO1INxp6hs55Hf2hZ
KnNjqiK/KIloehGvrgDUCsh9THu2rKuWgSAcPMjivRdWbwGowPo8nTp5R4K1Viwx
Q7h/drIc+mxNfgFJX1z9pEglXJePxrfu0cJlKS1e9gNU058L9zB+nD7NMOm+6n5O
76AEI0FvbJqMT1P9o0yx1ElxMLAk7Ef27phKI9sElm1cQOzWZ3xKdJKoBiOjgeVa
Uoe6mpqsWbIT4CvNk9BLCpp+6+mzU7/iE/E9wuJp01xfG7DM6XX+hQJbzyqj1x3T
yIKbGqQ1+zPmfvHCzt/zxLqIJTGrFLM7nn2dGaakcAurSHA3gEhR3zvQfcr53bF5
pA4zhpPEtDhUHDrfyYcKi7dwWmPaayjeZsKTioEbEDJSv3085vNWkFf/W/ZienUN
+9Ui2/mvZxRaGnK/szvnGjZGZYi9xSGsqTVXM7u6/dy1DZJSjpcFBTc9pa7TPvUv
EYVIvpnHBs5i7ll/DaVlKDzPeRYRHG8a12FttprNKaZnhxAYF/6Tk9FrSXOmPV/v
L7D8m5yvrDZ5s+/r5m579ERBoEWi0MqA7LCqdLv+tKvw+QM/9MvdpwX3gxcG71mh
0g8Q3JUZlCm7H/JKHsU8i/rO5ilbqNRC5Y88Bm6sA+hgmns6Zf49CKYu3lqqzz6Z
fADRdrIOw8eIS8BVjF+Ke/cCh103eg7i/aIQSX4H4uGh2ArGTnYxw2nWA+fHZhgI
+eJp0IURNP2/kclz+JPeIB7kgtMx55TlUFBwk269AfFa59t2NTCY0VV07ZfhkgX9
m5RbjhBMtXLJVP2UYoSCTlz6Up7bdrpULthSi1E3DvLZObydGL+HOdX2nmfRI6my
DCzsQoDtG8BnYBhZMG1OPb8JMWyoLEWJTWfIvDjxJDGWadmcrwOwpzHm7d7nOef5
UX3RsPdgy4/tuDMrsUIcG3y8cXkcNQlDfzvj2KeIguY83QDcXyV5AgoC8ChVAWMW
mVTmPqRe5qqgmiA/SylFWAfGF/4msphgVfNZloUGuGEjRp197JXJe0Qj3A2gsGjC
3+zvOOgH8ePMt0rJc8bgi2yTtmH1VXe5ekSBlHDVwZ0lBnSFx7msqw03p9QGsw19
imrg8gazFpEwVeITc1g3ApqE5uFwZqXe3Ary6WGFgDBVQCZ8E1u2GPNau48rOoq+
PbTRcpAVdThGb0CccWC5k7+IRykSlikmGoan3+3QebVYXgwTSCZLn9eC8bRwuGcE
CAcYfODQ8J+lgO+UBMuALBYFttuNLY34+p5uu/imrLQbjstrKeYLPZ2ImpSP/xFY
u2R2JLnFSNmmnIYXu4iLN+JP3tf0nqkrceubgpXV86UN6FCsowxLdkS67O4NOpCM
SR4puXSrWhlup21v2zlJXgeHUQuMf+Sgqc6EfYMucMGF6qrewZoEzXbPlHScj7TP
dxiUofuwY1+u2lPor6NXZoXIJ/XdX6Q+H+kKDV95e/6MYaWfi8ZaET3wuQcUVUEs
5u3+xSNp/dWJ5ya+FuXTZ2ddQXNt77pjTAY0+a7INg7iZzmYxzR8FVgdvOtVW/X/
Wnt3pOQEVyrvweKiA2k6xbnTiKSJcB5j25lAgChedEn9gWYJYHpdy1CtPP+51yw6
/MOgSOTczyUt/FnQoF0Wc6f81OfIv+5bRAE2vPMeIe7jhA9OVQTmvrzxmAa2EO6A
tY020pmhfJWpJvEQ2HH2DtIG+UEJ459V2+JnnJu7ixI3ox8LaiczmeNeHvKNIxUW
LpEOJCiaeiujXjstHrYyi5f8ltCGQsbOZNVtnZWpZEMtTQTsDrFuEtuo/YAhJaJs
5I7Hg0AnBrDZ+u8uK7WsuwgJ4ZHWJIT3R7ntwsjmfhw52UdX4puxCsXqe8j8sq+5
NWTzeqAW5rzDnDJRjWKquSDEGad3l77Hm2F+4ObwScSdfV9CVbNkIc9YuDC0OqKb
1+OoOODZGoFF3GGtiVm0CKgBFeVB7jekwMUEU1H8KGH6xTU2KaWaSUchb//uBBPV
IIMTTvioWrh6Yb7mJF10nH0rj7QI6R9trg2bIsQmbUXBdtpg284ExP528//VpRsR
C6PTeVQD3aUH450Hmu2EaQmKw3cxtmo7SbIzJLT5crpGGhljLvfUh3QCDqei3iLH
auXjXnKY+/7TS/CV22c9eLNYz0RA+Zw25ubtz9LIw4GPYRzofau+zQ+o6QgBvCmT
ZOcMHyA0M47HKKMITrZs1UKiSQMnyiD2wj7xLYzYEtK5EACCOKXDVfOo1PWrB7pg
Mg6N/voxcIk+K1Y1acOS+ohMrJh5A43lDGzH66yqHF5fhIMGG/VdbIz4ScO1/tBH
HdPHv0+EaL/Po0GZE3XqMSizwOgm5p84d0sD1w3zJ3A95VwCve545SH5PEk/r0Gu
T3snSY8Bzr/OLXx5xo79MTr1doK48E2siaihqup80mNY3pmiLysrq9fB3p878+xz
cB8cg9ffnc1wO3E3VIet43mswYx9sj4ow6Doxh0X0TGlFaOmO1eK6MeutStTB7Z2
HwD/BXXQ8bhomBVGLuckKYOZED6n3gq1d71NgElV/pTTDEggUvgfzu5axCWMH3Ck
EhGDWZoWyWIisiW9HcNEkw8vXYdH+5NrX7B4GPlq3VDfCKKdVhe+P3WFx3SCTE8O
RnbIuVtcky13ueRzYOBSpYHuJjXiANYzNMqu6sK1gg8grTqHlvkpHTM9bQYWHlLQ
kvz0bdnROhyy/WGqEPnk5O4NDtBsuwGrNUAZhuY+0G778LBX6oDA72kuJCEjpnj2
pjHB35LB3ptckRzflboRMfAYs/Zva3eW96pJPE3rFyzKAQwEBSw89p8WlWwSnlyd
IkA+XUvRJYRJ2US6Hz0+PY7zuFNLeU9m4m2DUjX4Be7ICUhBDD4LerD6niUAm/pM
AbdnzmJIUOwTj8YgGa7u5tE491DdkbqWFhmnO6cx/W7xdtBSb8tES6snyLxEFUol
IpbBQCACcz4ZZWvLPdemNt5wCOiQ2qzWF03dA5uqID06fqUpnLsJzAHtg7ju7EEj
qVBAASdvUY6z8Xi4SfZqksokrXN9H5CtSl3JAzgczuc6MxRoMkIZzn3fN3eJdeSz
4D5fG4ZcgxPQIlQBcb2wGIHIogq03e4BpVoc3Q8CXXRoDvBTntBG410twdBFTXsj
qFp023twDNnr/yEleknnUInpZO1HBgcWvhaHnnQb1dqaoaqHhWEIs9Kzx/10k4+d
7B2HKBala5qp1fLAHbh2NdIpyeKdi+o1d75Q/2H2Rx1tv5d10p5KJKNxySLAdEBv
9Wd+xO4wPODycX47lh2kZGlIP2XVHCsElLiWRMcOYf11dXndksoBYf/GIKMCHN+I
IfSU+RDwWG5Nk9G8g+4IMi1lLb9V8HipBJ/yHH5GFpHOhMEng+TxelIjNV+kwHUz
kkozrPyF6nWoIOiXFjv0nZOcf65j5PvF06IFCb3gLczajiR3/Gb/zLfE9zc6Ri6E
UabBtuzy8CeeFB3atircvfQwgNuRKCJeG6Oh8rBrA6C9/g6mHNVb8zF2IvUHgTPR
vZVbSDKaMZrofO0t0d+o/W0b/FaSoJrwc0bPpXOkWGLhf83lVBRxEg5Z94TMnOM0
lUV9L8WKXIFVZuUECiFpHzGcjMpMnT5zc4O5C2Q/GZtwbQnzMxDK+sm6uKIyPtPG
eS7npOTrv37t14HISf9eh3USWooH3SY18QIyCUqKLqFotBaUofu//bPStptTPmc7
ycyuEImtjUCh9hA77UgnKHU2xGGkCEumue1Jz/3kefUnEJawykpmA9qk3TaZxElG
0uP5MkHtq/o1A3N+/KesxLGL2kbduFBgU0IiGvtbFDTLhFDrZZlzD+dH9uOHqFo0
3sROdU+cxc/IjkRwTp41mpo5766ggVsasS52wLFFwZe4qbXZOed6Q80WbAA77cOO
KAHw2hGOsUdXN1tClLkWL63TRmp0K3isNDFKPg5Z9KAVC61HxF50awJZOL3iUzI0
BddPm71uf77hLLam8eL+FOLpLp4StTtN+koUj8yt9K8/QqF7pU+IJZSHBMjUdd5W
Y1orbeThaAkMc0uZpgr019vsPW93WPizxpnLGPaXAzeQRm5IDo2ijc+H3y8Se8EE
dO/IHZezcK++dXV//5cnxiHtCGkyAS/TOFtMJBnJ8U1Sb9ZPAxO9X9MkOzrhrZUh
/KsMiTPiJm1ejYd/nstklcIlPD/MgTLbtH7+DpCePoaFgKAZnETdXVj6uP5bzpJy
YTuRPaEgNsaZyHglZeg1XDDz9z3cI2jRM5KR2xJIdPswYO2dM4aby3hTqtk6dQl0
U4domLlnFbhGz7UqUphpuocTgSMUFaTy9Of5VE6DDB2O9CgDXGV8yDqHum4iYob7
yjCWHWKGWGbkpfcsfKId50QgsST0QwXB9n0kDNFVaavu0Oq1tH07EPwVYtPQ41fd
KdFTxTWvYPro0tn2NXNlk6H+Js3Bo0RV4Hltdwm2TWSpCfrhZ1hDfwYKz9guiaLU
QoiZgs8PySPDVEoOOV6p6nhfsgNBM0P3MbErmnQE4mYBLAGo97+MfnMOtWr+ZZ+X
ytNjMO9xpvY1UUR+dMw8EsFzHKzrOe6qVxr32lgW8GylGbypdfcqDmdiVe5IBSMQ
983Fw769Gia4MJzeo0TEFbgpfTgHhJWD3vmVNmfHr4lWGfr/jsYiy+h6psBQ2YBs
0lK8Eywgf9f8K8WqXKBdMO+llfIzLapOwy35afZJafmbKehwJHTd+RjmXYFzzYZJ
KV/gmb69QL7vFG1SP9Ju1ghoXlUzOsCh6tJLcW4Z8P5ERgRvo2h5FRtINSek8/WY
gikvQQmc+MzgAoApOm60smuNJ7tzG59FNFpNObxlXRAumIf9WSulhONIIIwcK7CN
xcMABCH5BXwDuZtRx45B0JGhl8UUQX3YIEI9qBwoREPKPelIbFC7C5dXNDm+X6NS
YEmlTHhFUjCwWAMu0L78IcuqSfXbtN7L5f0JYS/7WX3YsonbuRh0049dHCCpIzpv
5/jdybdCx7w2k/JOIIEbKnOJoomSYYuZNZndlMaDq0P6wU1ChydBaRPecnFFOOw8
naCsnOYJb1CVuYEa/6WCjIA+adeenwx6BKVXwcnCHWx6azvOHFt/qvdeeXTUo8B9
6ueWTdm+t2/+nkRuTTRDxzQi65mSeDd+byTC0/pGhMeaIx1yiHB6tv573lWGKKtw
0vDJOmgS1K+0aWVnP0iEUSJYqE3+Tr1dOmVTxN5fX71+3IvGZyAucNHQgJ3puTbc
AzYlSP+csckRmQ7hmyUkbbRKi0Wy9G2wp/IsWyzh8DVaiSTltqCGvkP1uq1zjI1G
M1WhcWO+H5rA8LRjTDE7y/UQtFCi+HTID21gCNbPALzyM11yrIzbI3jOTdGsCTfT
RIVjGhyBRmsyvoXu3g9osF0BUnXpuX0sum7jTDIwg0pln5Z4YPs+g4mU2892W8Dg
XIbC32r1G9XhQmTyzGEWtjCvD+EF3lQMRpZePZXJy5XWednXOZBJd0jdE3D5Md8H
3RKtH2yxsWRvI78Viu1YeiRug+MR70W/l4MSQXdE9OIn2K05x/ATUQKXGgcC+8DJ
90GCWuexgmzgY+h/9/UZpuz38V5NC42Ok8x7m7DvlJmet/1hiSlKbCFmz/lx5B9S
pLAv8XjNw8jory0OVMbTCWcNSSe7jdG0LVmXuwXo/5YnRVUMnt3ysgqjeQZO4cpZ
Z/lSEcKlblMunON4R34uFC10tyNaPZI2eP7mZr9eVNJ6tsf3Gcku+DKSaA0VKxYz
XhxrVir+mlXuY0yUbPLtKCFxnUCaAcafYslcNQ9Ej/Q+8OzQKSX+6rBhP8GY/Oax
4gUkWBVeynfRVTuofQOEdSntaWkyXCEq6KYdC9Z8RIOshdaSwbnjavC5bxgQFhlJ
EQX3WChIpasoZX86DQR5DhfQAV9jAyJ01Y2BJOqXipZ9tofuDCfeCokL/r/iPEFR
t5/hmufwE0+MpH/OdBFi5l41GXSCEgto3pUOe416JDt2OywlHsZ+MtV3C6yHGYCP
LGjeQ349vMXWIN/keFYtbfj8crCBe3oUFiOk3Eix+zVEZoEVYTqEdN+ycJb36QPS
Yp/1kVnqik6pQ7fHk+JQvQvD8a5QpBdzVDFrxpJGieuCtafbEnOC48AiKjubbtlt
4zrYK0nEWDYOLWpTZUjheCVrm7yruDO+yA6dyxL6sZ/FHkk6bPKcHkEAJsRlOgl9
Tv/6C8b/+EwgO85OYLHC+ybZ1OgzyT7F8BLYiV5hqrPdV9Bq3UuGCcSzdksQ/35K
SkunQh6MR9/xTLFpvtLGzQ4QlshQKe2qCNhZTAqRTruUI/O0A/DTFB0VV+Dxpjk0
u72NYmjHv1NDnt2NTCx3+aXkGBIq0nhDyeBfwXuEbT+QK/mDb0QqYwqyo/EonoLF
jFpEt6Z7Z3I+uGd0VkuBOzGzwq4oES7C89QGpz716Rl0hsgayclI8AQph13kvxai
pHMBPllJ4MpIIl5Uf4YIaTAfLvwk4nvJ3CoWs6ubypkrhsrbIgqubIWURVip9Owo
IzZ2w99aWAuHfMw11TQJUHisFqiwN29AnankABxu0HoIwtoghVBPMQ4ralXMoCCK
vngubOJ+dXSRnywx5fnUU+yCb6qvMR14xfEuNin6hgxxPMisUyp8FY+cSq9xuIGR
IBPYBfyvkLN846gVl99LGePAHhHJRyb/FtYKzTyf/WSB0FZSSm+w9RkLikxJYb+J
O0r1CZr75i0/AHoCHKs/W+BeXBAZyKhzDf47jEcTXD0w+eMkgQVnGZpLbzbBxXZx
IZSCkcjcwcd0K+VhcjLrGgADBBJ67zF8y6/vMqxDH/ioRh6MwmbFUojBbaaAtLI6
ECjLeAzlWJcn6ZuINSFcuEJoUwwlKdEWNtTrpKazahMQC0VkhyTORznuLWPq1I1r
hBUi8OY6zByQaP9qsn++uZBS1WN/Zy5V5U7hCRtxm2kbjXEZ5+oGyghjfTai+WqZ
vNp+7MFpCVbyoWUasL2a+tZbwP4H4slyQmitXOvJlnFC6qv2aCSVYULFZ3RmedVp
zcamxrSJ9cKfHtb9FljfQ0FjbA69j/BB/hTeusDaSKIYsBelfDOwek1uh9VQb3Q8
tfdbBzQQG7PfQgA6E1mZkzL56VxZ9rHyPODkErgwcXfDG8gdQOV2x0stDtTTfDon
FE0FlxJkAEnDPdStwaUJP6OqokYR40UW7krvllvxATsNzQuuwG9U61yilkQAk1P6
7W2dBM+KZ2uMJdfaVvFq+k0NJdIcrCpnJyxnK+j/9q/NbZRUm+iUPX4MPrMwylU4
zz6Mgg9LmbzF4WYEI0xdBxjgmVvvQ6KQ9VMAON5aZDfOAoFiBksRnF0MffarzWI4
kBJjDWktpf+BbnJUoGhCaV8arKiQLeepB7FQoQFfNrHW80OYn62+Ht1wHUMrUFBB
D/WuOVsGM5bL9TByGfc7EVHK3RrDSO+EslkmAjXImWTcvm2dIDRCi/28wqkNdwio
atYfBu9ZpJEuqJu+p0IhHSGJf2nEyVxOF3Y2U6G3SWgTFHhMa8G6PcNCN1mJSdoB
Gb6CMtibJ5ECpA53FuhK5LYb5vbUdhQoNiDgmmgto7cuKAFcbe53fsvZIaWpltV/
s4nZs27wiJBuiWDE5x92KMw7IigXWgbJfpPrJXmz37Zay/RTNroqJZvHQ9X4JR/z
FIFl5GTF7t7V24HKXu27ccfTeTeRHG8M9IpfWvCezM1jGGJl+Jl5hGD/k7JGYcqm
q0tcchf3u0PAlfw9yHxsJftQk0SDmRX08dhAPYBm3qYOrMTOAFoB/Ysovda0mah9
+0n0eTsyc42N4yVVjD4qEZ2mvVZAetgF9sJrFikWy4+8tkLiyckeQJK/TCcK/xXQ
Z+8iVzhbA8xXBAc3vSXqsXzpIcvDHPrHBNySJ0Ztz+tPhFGIhb4nN3q35HsK3UUn
MJX1FTNwT8FsCRMeDEZpdwcn1Hox8sfRTqTkaqUiCuk48N8E5xInkQoHlNKP0rrL
XDQlbkoqf7K7x7D0Br/FwRkSYtu5/Z0AULPdQMhgQfcfkh7Hk/UCu0g7gwgk4Bt9
mUybtZjsDxQbTLztZSeOrgytUdru3Ri6C5vtLkltYydqhJP7j+evKi7NWJ7X15CS
UaaXxVtqYQhYX74bJrdLpB/1bifmd4jFhCADhGNPro2FqDYKeXnhCAlX7KoI5SWM
0cSug8NXcKgaeF6UCF9NQS9ZWfXdjNAJfGAHw36uka2xCIIkXUARs35ARYgBSI92
mugsIZUlY20Qx9q2yAEWRDlHPCBz3omnf/3S+Ocf5VPyehjkqYp38Yp92dxeIISu
RGrRO5Z6W+oXyA4dXnCpU//6en216ZRnNAg3ADUdVcKzRpJg3huuojJQQsqBOGLu
NwtHXBG7xzLqHAHunA1puN+Hx23pnPLUeNfmFGU0PoJddzTnhqvDuLT3UVJP6d2/
SmZQlp1V0OTWXAza7HwM9jlMFWLJgk2aZSlIEM/3eDLj7OgNvkQ8I5th66ls/8fa
7y2ZpHiQ//iCAkHozqY06T9anv8Ysb5CrZIfVmu6yzouc/u0QrXqDktqo6Gm25l3
fdDbOY5K0CbmkBjC0QuNHd8DZbtXUw1zBzCDk/QnaXkUAVHhnQt7sydyBzLiBnWj
D5989kvrAuqC4IzAi1LjMVt1hF8cunQb+SV10/6OlLieEQJkSVm0meFTNd5obcrp
jBNKkYLiebLwFHlixTeM7RI3+GTUl4DOoytzIZPuQBoMEI2Qp/RTTtC4kVYRsAxm
/ML+ar5Rk9aggY9hxKXrdE4I4a9hMLTLJwnMnQkaMWjHxN6T2iBo5WMaCk4mPaR6
30AM5UMPiyIYt9YjeSnkXkEfwqroFgdu5Vdr4hVd6pcd0g5G8S2VpCsybGOGFl3d
9kymN5RmS5L8Ot8dgeByXLRHrMwqVtfSNQRI2ZtK1tommanEvPLK3XnVvjKHOfVu
nzNmJo7x1+4lV/YI8MRFXbBXEV0rToZ5+OOUdQ2Uzf91ul8r40R9bNMbpD8kM3Lg
tGGAwZQund4mhEHIRkd0BcgkzaJW7ih/0lR4zpayvz9UaNYNy20WUonr1mQ0zNcD
0f2Fr5/jT6H/C2v7YRPpyS51zr9rhJ31Q4A33PbdHpws5m3VJJ0ekM7YFiuIqZ62
HT4uXl2l99fEs2gXNZ2KMFh8GnnlJM+6ekexGObgYTcEZylqh44co5kjxpnFozN2
U8bWl/6/5Gea/qOq2AgYOv/uMnRA35tzb7sUe17NAafgtgxk5z9XU0xqyght9J46
JhuHL3lGUrPPCbhoHx3TU39JWcYdIRECz9CAqTiS3x+PnlC1ZQXNVekD+/kXClnw
XpxRSLWPkYnX4o+hwSit0G3D2KjPgbLuhHtewt+oxataekhN4fprWhwrZ1+dfykY
2kJE9+T3CBOPUj/P/tMbbTSLD8S/ybYMf4X8AJuKAhC2RjaAhKi5iCFzhJhyNKkI
psGNosluQMHxR6TRlW+j875KhqZORUtPZ8jFwMtlen2dxhg/h530ujREZ8WAeVdf
asH1SmZrNyzK4l5V/3Y941Hr9A6xn7ACdHZVXw4PxNYBjPqqSmnN3BraEyIXPKo7
JaFAR3IS4n2xDpOIwX9rSpaUp1kPrv1NlhEjaJb/+gaGqv8dOhw6nVGgPmBlgS6t
VBAMEL6AAj6fCkXbuZmCG/ZRCe4p+3shxU3jN50WfA/Z78779tASzGbjCWmMnUyc
Lri+TN1XEr5y/NiTM/UtkgwCt8drrUrQIqVzhfk+x0nYe0ekf3+f/+M/ZVcCYBof
nETcM3jAS2+W5YK7EvtqFrsw3fZIOy3/iVdKj5CXhsqUxQln9Xzm8UR7qTx9Af6a
y5ktAe5hU+vGnPcDlYmU4vTmnupLNsYdRwg55rIcrUpPcoUEtfIAJe27ouIc2QgC
EgYoZe+XXF3ubf+SmFU07fKUs1Sht0ja/meL+xqH/A1NHMuUWBGHBWYigGCRXRfQ
QgTqsj0Twf4hsOOeVyP8iZkBPFbp81vJv1/qQE2eAnNJqRbG5yyO693+m+naz60f
F5t2csP0uXW8RrjA2gWqkl+JeZCal2Tno99d0mB7T1zrh0LL3keo40PQgpWAIaU6
ntXzrmDWigvGYY2tC4n8RqoKWllitCpB8UhceuiRWgX1evFpB1z9zAjOjScfdKX2
lmyljwwTJCtjv3BRpK8ydIPMDxTxwYHDqSX9y29XYGSKm/djD8u0xtzj+TfUNB7a
LpngRW7w2pXOiLSWAUET8nUtOMWYIHwvJEOlxKJT1fnIYm/lCMHKeDgLhuqcmcus
zc6wKir3RRSlKVS1hoO1btCt9A4mGDtcNSBLMDVLnLH+i1QrUkxBx2OWFq4+/v9w
gfLD8TkwVsx8j5FLEUUPr3F5/gyo6x8iNZB9jYud3OUXPLr+6XKFOPuaaUCDYGN4
DWDdjGU+cjpssTeYEyt7em3qoZxa15RvtReNNsWZDSx/f6e5bbyGqIgzM9qHnLoS
nI0KfmwWVgxiJtvl3Qvto1YiruBZiVje5nhZVRt4A7NSkeCbWwyqDkNS/AXbxeLG
4eLCM00ajAG/zo7QjT2IwbYG0p2TV+BSRt7FJ2TSyv7S7R5P7U451UzaW6fOF2i/
uSzYb9qjVtZWUE4YFEuquMYlFGp4ddVW+UBJXaaffWQcaaVYBJhf4IM6UQ7pbFie
sPW1A+8zpS2tU31b1/kdaA69UeP4XVMNyyUhjLfKjUUvmqmXGFc0ryDXp1whyzCa
BGdCxtdr0OsdJYKY0eRZ3oqsq8KzVJ2SZse7BcJD1fR5M5dLd2YQr4rwTWI6K4On
XOdV1+a1gVUZroLxiQGTfsKV69LGAusSrASDW8nuSOcwlfANiYmSDhW6YKILsXul
C9/x4TMjIP1GJAdGRLgTnXTXinYhnce5kYdMTsmmW8DNRbwLr+JzAcqDxRbXslC2
+eWg6GKTpwWc+7LFYiPEY71f+LQcujCqiM8NHzuSWzp9PcuihQ4GxomeYOcPzgPm
mpesuLbxJ33sukYcL4PzbFRW2SiwEp9hTwXWIZVdJBxFA+38KyI+TLm0gDujxu1F
RV7fhSfIcRoXDTE9NCiHeDNnl6klUHZWhfvYcX0FJXmHp/+BhWuYbYETH0hR0BNY
qnbhyrCFILv2wmTQ1wIoa7HbRb3qBp/zTDtrpRO+TU7LAJPyz3M8ahV7QTY5qFZW
PX2Jn0q1mbOMkRndN4g0O7u8S5+K/QQ5GDM0dGQx+LbpfPBaYoUzBCYtO8Ol1IrK
hy919hPaEaH8kdd6v+tMsvaqe3zFBfzA3cu7LvOJ2zH/neIfdW9QiEXl2/yl7L02
7y43btqVQ7zFLMS7+Q2uDA0YTkQGr81Kh8O2yfhyCZliqMMzQIFTfg4RBR7m2nup
MQb/ZC35uYCpFFzqj3BS6LpoN6WAmLvkSfFBuzdfSmgiwlkwep5Bn2aiFR9rd6rU
i6S2UAiegiWp0MG4lvMYtY2SsHwb4kc9fX6FIe/Mr3BOqGr3JJnlO8AS61/kCfCV
kq8MlXf4iZwSil6gD04B9PSAHsYNXjnyQGEdS0fmRPS5r2kG7thMuA6pxJAJSv0N
aXqlYXcl7O+cCD51bxwBLJdAI73vzci3mYI6S96yNC1D5tzHubAiiO1BZOs3GNgu
iU4sY/ue/+lUsYjCQhwAzH5Kqz2Aw1ChSWUKROZoWSB7qdKsWdjnFaEuqsXra87L
6LeK9gexg8GYP44M2eGbHPy/FHEGnLa0tEqTQbCykYdiLYGX05oob6vmVU0FRBVJ
4Q2RLGz1ZQaFc71XMYcCma7YlIbyXZ3EFlQmMW+1XNlfE13cEA/asm3i1P4GMmLG
V1MUBnZJ8Yjt0qA87w3O8jwGWgEoQWG4biVdlRds3XSUKPFRBEQyit+fCpajVMSc
fBA6pZ8NKMWpWBmiFW5UYfR+qCgz0yg6OQbMFYFEELiRtdJAVHvMH6y1MHeu4Luw
LKScq5H0TX8RKLA3OBbXmzPQPuwLi7b5TMo85DlGRR0D5B1oxQiVty1J1WDjkhn6
Novse+GIQJuNHZpSdF3nwL2J8EAL4cNWRw+J4PaUNTyR6zatdSAvqUpEO9rY3ofo
FhyEMm9NQAFgLPlww97j/kaztrW2B1wlpHrmdNt7XqK8TjRDCoykhA2e9oJn7naH
FGHMnNpAfjsJzY6Imsue8vmi7Q0x4fahSwqoKfw8PXjGZL22glUj3NyJVobSfbOy
aH6Xhi/dcvRmDD8CEW3vPaGGlmTtZSzvi5ItUmSbnCnZpprBxYw4MeGrMcyNqljw
x19HkNrBq4/P6wsTsL52P9loNoZpWKIE25RfLRwF2jqw18amTKXC5ST+kH12FSkx
15Y2aJJBaE5f4LSJQGSD6ggX7k0eVWAZ9gvUA51RQYVxwZM1myaLp4NkiaOsmecR
HCw29gRQaYOXOJISEBt0sxcwpMzgsiPWmBaY66RNo/o5gN0XAX6wdZjxlsBtVthk
aQ4rQRUXCsn4VA/i9yydxdB5HEir9wAgP6xvolPllIRm2KxqBVqqcY9gSnq13gIY
GAorcoMviPo4AK4TiLERzKipiRUk9zrJrWOH4Kpc75Ku5c6emdNR1Ojucax4SXRJ
OjojOVlI6S9Dync1CKCUyn9n63aiqQpR32Ivh64UcQ0ZshXHxZcrJmo/ZupqtdGS
tzzh9VjuFLM8lWnWmm9dh2wtixmUpnMkEKgH+Exq8E/9NvXpmjmNYRDEDiFjzqjP
O0//bzr3pyY5jKRfjpeoH8CERsAjT5qzls3AMmQ0G3qBGlPUIMMo/Io0SFLv+zhu
Kq2YI3kMfK/KNHXeLsNeviUW/9Rg+qOh40JQ7LOAyqdwATUIHklrj/f9XhO6op17
/LJ0MFTQio6l/tgUei4T85WyH1l5AsMouoGZI6swXSagk5RCTeV0B9xuyZf9/nbx
xjGj8kFXHAR3MDbP37z5jt0NoLPUl0/LEu8mHTGZvPz8Q0ZVHbXcOdc4mxZiyQJw
yj52GCXdvtCr048eGSQIuY70yggdZn05CZ+mIv590m2+VqzDskzs2E9FtbqCTxuS
3smC1czzi4Hn5OW6IH032zyGf/qn3b4AMqAW61CWnCYomvQn60RdonOqlQM9ruD3
FbhIsZ0eS51JU8lypuulDMQDNyBndKXk81AgzIpXoBrBTyxy7ntH27Ju/0obGoxs
j4VIkxKHgHB0BX+xtzTF7m4pLrLLiQkv+7yRW5suedJ7gnmvyelMTiqqpjSfvvNV
ZWLbvojboU3lKBqp2A4TocPLovFKdkb2xOc5uQiGxPN6MIJsYl3odMLfhj4ZrSsQ
YqEfRM2hQ0P5azen6uIKilzH/9Ro4VMkyEFa+PqbPAXQUsqokxZl/AttYfXhCMjF
aaNd3XqQzF1LQITd/f4jrVXfuSF+NzxnWvV1vwpBIA/OlPQXzV9v13zsMR0xJxOg
lWkhiNvjipnuUgrNOYjVih5B17abcS34IcLxsf/xqF9L1b0rYzkY5Y2vuaf25jcT
2efL87h8MQeQzqBy51QBrHkUk3Re30r422vrQYi/SwfqzGh/YDRE7jvR9wgZE5iz
IRxkci2glbTBoTgifg0HBYYDM8J7zfQhQeRtQNG5DvKDUTEOhBfT48hdpp8OlzqY
qUgw4dLYrJFttyCNvbu1TDsi5yZorW4508IaX2y2bniitVdUB0EQpftjchkRQcRd
aX3Ygx1oWYZ/gx66YX3ql7PzKGCAFjpi80zFBFsHdt0LYLDOlaORgfAcsBGaVwmK
f2i54zR60prZgcrcis30smiIqO/SSHg/6/UItcR06nqAbFD7AU6tSfp7yq0BirZs
vr12TXE9VNVPzzUbT1TSdJevJqHLhqO6NuMDrHL1KKj12YeuerARKJL+1i5ouBum
x+7Ljiog1/i28lrBhU9AscbMJK+T2ol/nfaeFfu+zR8QHbQhmLJ93fsyVLS2C+PQ
kVlsDxVCVp+OF2s9nwlye2wxu3JrIVPpty9/jsDeb9pDgPuDGC6ee9mErMLGKo5g
tEzyiKNsbJq2jpf586BqTnQ7ihNPhV4Cv6PJ33gR5CZj6o/MyHc6euf+lF53nCKA
Antcam+1DZDeMV+EPpMSjl+dGdFrG2bYjvP+pUNInEcz593RMwN//JXYy4ZF084C
f8b8kSVCE9i/6KtCdhELKV6TuCBUIA4foxOwTyRK9WcEMOGxT9bGqBbJO5TCotza
/wKtZUcoCSRM6RoXWzFywqiiNXXaMuMvrEmVBpAAEpXh5vHzREZ8oSHELbjj+Y8w
0l8aUubW/j9kY4keGJQuxRc6HDX+TgffYVO9f1wUR/WV9GiTHWaLaIhcVF9h/c6S
fl3Rad8pA+XQuVNw9keVmkkjmXkuj1pNL10GudvdJVjevp6KZWkbWL1X4CjVBFU9
oqyHAMWNz29n2saX9WqEx+Z0RSWWZh/CYo2JJKo7IQy4tq1F6r0DGJVuDTjAbkp7
kd5AUkBB/leHLvGpBCuf+I2j7SKkPpzDoBO5Gr2r40SaRSYvLZJXs/HDFeF9f4ku
bU1h8UC2IknsV58P8ddH4Cl2LwPpDbquZoCgTiBqLpK99EOgtIfz0vFPFcol+4SG
xxsAxQG48saO/4JA/17UIBaKk9MjUTSAPsGXTBpMvTT2xnxxXWI7uEpwW8D1Z7+v
Ti24yIPiMbLGugHRKo0h4FjBmOkgpKhp7U2Sp31E+sOQ2X3Tg9QhEMjQZHOsS7J2
zTXpp/DLgRTq3hx3S6rO8hCtKdL3SuZYZAcLOIl9rufxeKwhvGPsirNISa3xAIDH
mq5M8C4ZgyvNEd4x1h3eBfC/ByxcJ49UrTfsqxTruv12kImhjZJkV/+S/z2r210x
Z+NJpwhzNEYTFqUs1JSlWi6N2vod9SRRd/1w1hoK6fcMgwk8WkoGofOGe5jee0Qy
vGSKcckeKRq5iaYEABmd2vYh77HdVAKAzFDqBoXSZ3KN7md8VlmTio/nEmI1mrYU
71CBx5webddP6nmuSN2MmpGN5WxC/Y+BDRkkG67Nc6m14JeZ30Y7GqiQlzq/hq/S
siBhIzrbnSv3LKdXsKovdLZfYBFDoNbaXrQd67+fYdayAA4UKegb1Xhl0QUbjECl
JDxIu67m3Pl/hsTkp/U+GF8SUzZ0D8ckBiJq+AEhg59yPsqpLBCUND3koJutZDpd
Ok9CJMi1BFy9LN6vmBe6zPi6w4u8OD+WhU1tEJ/m/H3AeVF1KDVzHOmSIcCxqITK
6rL5aW3cJd5Eqfvu5XQizymRVTHx8bPTkfsk3DmW8teZnQVKRQmCWydnFkbdEB0L
KAHlp0f/vt4SDx2+gwg5r/hShSLxvgcwyDa1QnnTY3o5ogBa3homBRlr0MCeT3kX
OqPSnlSHXTPSyJkiqp1QhdtKdqbOtXzANQBtaRmCYfZZkfuMoyCTEi6wRY5lbKtj
1ND5YL3XZkR8cZkVKD0Cv0NcSsfGdEzUto204tOzxBtJNjedsnNCft0CsbhdJNWS
cGV5bFUBNzSQW5cN2vJ6fPWB2IlPKLELAWyc5YpYOUIBLdWj6dWU83rMk84PjOGl
oV0zzrTYUfUz72yXvpqR28IQuL9hrFHtgg+826vf94p4A0s839gHpa7hmkrGYDRh
pJpPvbeLdKc2yOeWHs52dSySOe1ZeuBjL7UA61NJhwZnf7009fF58y/DgXmtKE+b
kVH/u2HZEZP9mWycxj9HZ3Ilcny/skyVMGMNitTFJfXCxVvZeXg4LbMp6nZjvnoY
l04UFfq1+geJZks22q6GOzCU3nI7/JHeEncA0gPxHtWEl68s3Jruuqd+LjAk6Gou
vfwWXmTJzxuuaEHVq+r+xT65FFSo766FN2CNTQn+90XV69uOFlpsCSrFG1XLvSS0
3oUWsxsFq/g6Yb0ia82u6AbcCPm+0/BkVYPwtZSOaAOSIk9fH6Bvyt527fSc08AN
TuP3FAYaDYsBNvX9tGTNnzJJaZdGh6LdoTX/J673U2Fh+1fbGdQQFIUh8fa1t9e9
X0f733KM0acQ27uDQst3mbfvj/+QnEsZe5KjyVp8S/xrKDH2J3Ih1EY3dbuxxxrd
A4H/TPoohu/419H1KCyw/scjGnM/V97rrUPdBxZJr//oWsDpd3Oo8MKSC6gv4m8i
EtxaFWm1I4LVbKHoJ1wpnSV6CjOtU/tiJiIN0lylwbwo+HEyyVCk+WdrOD3cHCGV
w8p6NuznreHBVSttzrup3yfE9x9T2piPPBwKpZ5JecUiTNtWh+OAPUwCvP/LdUA0
yGpcuCRVxBNfXNwfBHyt1mR5QNu8Cs3TJOZvsZ7erXXleCI4UZsu6AvXzk2ussWs
eUWzhTrQYL8S9eu+0qqsBzkqvDsWtukpOk2RbktePJQ1VumWm0vjkXrCKV2rWKG6
ucO6Qhp6B911EwNe516kCIhVOIBO4RM6POvpRRs2kxgqox7ZFnY+vd2eNf9o95lX
8ZkARjcD3eMJ2YIDTtIGuiMFc4Rmng3y6Tr9xZ06464vISjJgBb3Wbbmx+UvGWH7
zPAVti6A+ftFRfLjtq/aASuD5xXwhfv/KBc9+xiKazaqZtXqKb8Vjv9Lr8ewKggG
Z2s60cxMEdfT3pxEcvE/gWvetPDhbidfTkBFkW066gVAgNJCwXSdGXoveEAHhUk5
N/1dRTR7+9c3u/7orkD4oPgf99ubiaxbzP7BqyWT4s7zUsMJ+OI2okJqIZn5SWNx
zvMl6uMQQ5eMXFZWq/YtdVm1d5No46rACLjCszwtmwylprO75UYfHfGtw6NDyC7s
8as+XOm8HOvTOt//4Ufih0G1DksdgSwyT2K6sXFaSTA5GcdCF9ZgI+Eum70nFjSe
GL2Zjs9+2jVfPDl6Jh2xXbHuuatqBaH4idHQHNrdxAPPwHXZ3tKV0wJpxo5geSaT
q36BCXJbW8/z8jMnbZX/WplMMiMi6UO4tWHPcrgUpKX0h3KAwmsJbIpWu+O85BTC
A/9rYA4DTKoVx7R46DRwJf4C4PJIkf8SU3BoeOonkxBa+LH6EdK7qIjjQWxh50mf
bVoCYFRdBN4RS1preaHTA6h2H5/LhLWcFY3opEwRpPGSUE2XAKfsXVaHb5lZ71wn
EsJCIoss8fuO1SIyi7eTUMs69NFjMt0x5Mn5QG3AfhTHoTo+A7SAVZHxHzZpZdel
5V12bc7rAxhfY+HpgpwEnAeyO3x2Mx6+52qQ4di80beQrpvv5FYAvv3CrimhF+01
9rNM0Yw7hG/Yw/HCDlv7ihxNGNeL3X2efd8qjsPxp/sacYLRU0aYxXGumcsjD/Sg
ZbGcrHkKdKRYDFik1yK+G3CUiZNIk0Rc47ZO+EtCOoGteFh9YGW9y8eUC5QTiib/
p1Tfiu1qqEDAWkpXY1JAPKtLNPmC6+fLaERuqKED5FwVKcE1hXZy72njRsIBIA5U
s8YyoHz9CiHZUFa2wjFwldyoNh6QMP9h8xPsECVTwra0ACi7zW/XTiyVL6o99SZr
cQ2KLCVreoJ/y0vbIF0r5v4X9E3bF4geFJjdjw8a0uCemwsOf7MHqHrrLwIugUS6
OoApsYXDqBsfvRHoes3tPCFtLJYgxWkeaReo/7krbW9Z2BmnSBCFdom0XKOIzxSG
fo6AWXaTyKfuruseGDZi10qQDwJcN0tDVE+YJUiQdeELftLsauvx3dZ+mKuq+AfL
kV7gWg7GDQJwiVUq6d8E7eFTqKu10QsfG97XpIaXQbm8D+lrV6IHQwG2RIB9lT7c
tOmKVdRdvnpcRk8CD2OQt1tQtaCZWElP1ASNWwLUqQDYrjNBqbL1iCJRhJLgb0Rn
PlhTy7iJZX+6ZJbYx7Xylf5R4SvqepYOnmPlsT42YfYKMVD8EgM1DXdiwqwWSBfk
QjpJBwRHIdkzSAJcUpayLiXlIHZAQ1Gsakg1/XPMLv7CB4wf/MEliNPm5Njh1iPc
S6dVLDwIkQWHN4H3VEIAJO55zTzNv90/skak/ksJ+xcjxxkm9W5rP3WZoqjW3zj5
u31I+mMcTgeUpZq7rgTTrNxqAPd7G08Frlhw1vaWxu/leeXKkygrGIuhHcyfLqPi
yr5R488/5sbw/i97+k4NHCirOUImpjEISvzhIO1oHSWr5ZXUX7f3AIBotkvVpBlZ
lxkoiZD27o7x22wZWC1w4fuQdQnLkgrCFBgCeWR7Fp+jUm1pFIdtnVLGOJNr8VV1
INwMeWg9ViuPZPGej9P+39lAxNitEfEjnbU04yFKqi6vOIKmKHoFl4nFC3x9bzMN
eov3QyB6uOTqf2S1Hd0/F+Raa7qFmU3iNOY6TrwGisQ2OmkAZ6I63Eo06AqvLC4d
M7/swfu/aGeTn4YdNDAQb56nt3DnySWWwBL6NWn8DORO63dx6rO5lVBuEVcsweBa
Raz89fBmt2Y33DN1Hp9x4K3h71NsVy4//6qh+ClHCe3r7qFQWnVHCM41rm/r/jNi
np7A0qfiXPNZHRfVAx3/rnwH9B9LlbRTdJXc7U2Xr409YysvR5fSCwdEDNJBP4HS
d5EPfT7el40JvU1fimE4Ql39nAxCTTiJ7mCWrdFSmvq1jXq5UXS9CwkLx58G5v6s
JN8ufFoc/u3Bj3n0wtZe2bG6Susb0YAPthSf46YJUTATgaCvYT3DOMBjpmC5ENYN
rxBF5iNWI2hwEbq9DIqV76Gg3JYPrzMbVi3ewDAxmlTjqdiH3+TkX6Z9yR0BmF4N
VrOW63YoQ4HjgtHCN2pX0MAokY2iJu5OUsxSUNJUj5J8Z09lvKIJwopCsTWOiJcG
OVLX0cmQOd6zKRZRxy2grDCIQZkniGH69FBTSZL1xVjoQwLMMQv3WdvBU/J0ZSrG
5OOhilm75QqUR0kl68PyjduLhvhk9UQBFuHvDzKmR9CoSowENflPLo4ihjfddpBr
iIUca5Nv+5hRcia9g1lkZZkWZW6ldSMvTFs2i32exHW5hL0oHHRUvhmC9mPAR/3Y
BMxOjUN4s/rkdkXfhEh+gRE/5kvHBIyi7SSVLhcs3F5s5kOGTopa3gZl3vVTkz01
LEztl6UV8byd/RE1YbhYw8sBaHT4u8yDg2IlRE67ne9W/I8BWygV9NX7UKgb7lSe
E500WNRme9klEki7VC9eb/hBHL5ndyVed0B631Jqc6lRpqf28+H9aa6kxQYNpVKM
f+Bkil4cO5VjSy+yDPqfH9JBJ67MuTrVhzQMG99H6mCddXEe/upGVbaCBsz5OIjP
9mMu2O0l9GrU8qzDrez47cWq+Qeb9Y8cg+ynl4aZCPefJHYllYw29tvmFymKMrnr
Z/kEFrbv2vH5iowmGeBA/LoCHOoyAZrlxNmrWRVqIi5ahly5sD/+h2mLXoeLLumi
vNgXUpI9sQe8RQCsoYYwhB0K2ig7UOVcfGpKk1WdZQhryXJifOxWZdoRYq+V4opc
PZW6//h9s0UXtuPTISvO/aUOgU0mCVwCitpFcq/Sotvkzla8W09ByvvycKIukhrH
AwJ5r1YcS52NSHE2+nkx5w38UfAyNEc0M5kDB9k9DHiOiZmO1LdF72o77M6fG/Uu
Se+ooMCDnjdjA4UP1UY4F6OQ0V2VqwERT+Z2cj7BOuJ/laRQ+QVB7keBvEOe5SAV
blJebZOueNmBf4UwtiGznZlo/MKx7D175bSP1t6b4BXHcD8+sSfd+iewMo64fH1v
qxBE6pi5jEzQafvz4WhUuxgWIu/SNzCRTzgmJZB1qlMJlQwVIomsNsCfBM089EjG
YpfQDUv3elsyXy/P5vqDS3Cbssuloh9zrEGI8vSUVIF/hnyL1ePcVJwgNhcSWv0k
PIGOd2I5zdI6E64cSPJfCavYvJtCQmPcDX0JN1HNin4KwhqiN1H0EW3Hqxj/kwdr
igGJ290IUsMXSbLTW/UVP9/Kqt4P7E0pw3tWcEj2msBB10FtmfmF4MBh4tc1lkWV
KLmJEhSGcUxjDZl8lJxAij1WWK5mYu6bGkpr7fvTaqb3Klu238SP0EQyVkmDNzVo
BMvse3UrXKVj9WGiytwBpmy+i9S8UrodZ7jcN8Ogr1GYMCojoNTDN9sC+gIUj90z
TT/TaKBXe6FbhyP3xk3RAvoh3q0xsrcNaEvyDe8HM0TbgMWleo6SaOMEy/WSus90
OjD90WamfMzUd/fUm5EhnrDp46gRAVc7C+Sqao3tZs200Vq3CwZx8nt5XdD21tQg
UgEQZuqABl9UsdcwGEJl6zFe8rIN4tHV8FpY0u8iojRHchnv9YR0VdKMkqNLb2z+
6Y4wHRGRChWtUM+9Xj0Zn90UBZy7Z6S85PtKchTb+m69oczSPo4bBOzbVrTV2rcG
jV9IBLZW+/CtYz2vu8icatWbBCYFwaMdxgadaBf6R1XSnSnS1v80eT7xIr5EDk4o
RC6+kFpy9LO8txo1qSWRJ/dcjqg30vcZQ9MQkPzbTsV/kvtl+KoOQsIuJ9yueci0
Iq/shAiNZm0GXp0lxMJTZcAm/nrekiIbeJvYvXy7W5IwaIuoY2O2e6bL6cQ/65Ks
CdVv4dxPLUwDT7CogGZktDJHcRWJbGJlSjCAuqH4pnbO8WC9fJ0vDfOggtlZKo+b
kcT+7VR5tLju8I7X7TAdN88AY8nXiyPjx5i2Buon2ac1SLBBXJuAH8RjuISr20oH
89ZczKOzwKInjSvLywN94DgPXKoU73aD4WcI5glXo4or/XFVrKcMClvWMNw+Ltk4
7xOSJvt6qizTrkdkdMz/tyFLR65YhRYWThT5EdKvtBIcY4U2mlqCnKlIcVnIFtIS
C/Z3YMLtZ8zexR9cFfxOl6B/ljTv5xrDC6MoUo9DIh6UM3J2xUgvEcnm7tKfUozO
PlTIgkz2P60CRPp+HdxbjNDx7thQOy0NWhB690z4Lu4Ud2p9PIr4/RHOpNMYsGeh
khkYftvM0Iy5wUFkaZkFzaq6I2wfOYnbB4hpSgnyBSKwiemQC2d8ZLTSAm4CAu0n
x/SfZ0QMlRftvX9OtRycKySkwkBQNM+FkCN3MNITBcxS8jcbUiwBki0c8ybneYoJ
12PrDnJIkRliDWuiOYWFTSzOjSOj8gWXysxvPXgE+7AFy6IKQdAnRrcJ4aYMeAlv
1z6fxRw7NBMqomR44aOTrILRtUtZgVrALdHwZpvC8JPSI2TOiji6HgtXi10wcsLU
wAIr7+48jfZn4w+7QF2/TDAHGEhn/9U2JA0h4/h3lhxbBONOdvUHo3ltt91oqXdh
rLRs80C/pLdwF7kEDdizeMhyuvu1K7QJwTTNi6EE8MpvDGUsdyIjwWqE9WpzErNy
FiiyB5HDzz/VNS6CphfCJQ3q9jfw2Qv6YDKrhwA1TltxAPjQu4G4eM/3knpSHvnR
3RGvW8Y1qEjwza0BFZQa8ztk+dZabTbI9hFXcKge1H019Uv5Cz+o1Wo2T9Uc6bZU
aNJjKmSs6w+QIpCZv4YIbEUPFXO4Qao9u5j1XIGn5EKuiHheCwJRrSoTtGxxns6g
dUVYiVsI8O+Pm9tK+fFfo410tmZAhRyDsJ46xP+R/9dBxaENoCBpZbp1gp/dmgTA
raimjCcdssOO3md2cPR0GOmq2fMSndUH34Bmaji96L8/hyUqsOQznTWIukeNwN+t
ZFuefuGxD0ik+w4g+eyJRE1Y/q7SdCkiCWIKAc7omwLeElTzqiz1O80TxsMCHf/a
rRfAqDfXgbpvgH/nueOgVG15imFgrcGR/E/neugKqfNUIQqw0j7KialJOIsb/+lh
TYlAjtuGAxukeNcjP9Pob3X/ZgxIkjAcg8ZIQOFEanUZdivDnnf8pwg/Stnf/hXW
KgA2w9TOFCQ/1NgJTel+S1p4Ct9SdDGTSO0VVYDXqEhEqcMHuiSn6eZJ6oxdhWk9
RePlpivRoMKlFR05DklX1Xcda9D1+UmK5Zc7W6r81wa81fW99tSwy2YYyya8g4SV
7cNS2iAWq6uJAAqjcD0YArB6uctHhRpj+kWgJsvCXh+8yaFEOuMn32mBFb5GMENq
tbN6J7aMr6+MOeZEXfKrYE9ilVgTkR2OTNrdGM4qMDphQ1y8lx5oM/tIhO058Kn/
LdX+Ywjr0tQSrZgudnq47N6xpYaKkZwiK5+UT1MsEUN3xB/zCDGnn1eb+rTf/xQv
ByDWqw+1GMKhSftx63X3AUWnmSaQ1Bji4B/wqmuGfru/37VQh6pbFcYGK/MWQlQ6
BCe1jJ+zEYBKBniH/Euzu6YKc3w1FuRFFB2QpS+D9xWzf2mh+a8G5tFLMNNDgBSx
xsFeUecQI0Fs7qnccRfOdEAQKLmVUkEC+SLVyLlKBGuDlitJBW62CpcOmZ9ZlIGZ
R5+h0qiL+8oDmJjqUlUXC6gzfXDFs7A3IEinCz0mBSfx00cLnNQjjHTb5QoYCvkb
SY7yNGISyKwXFXdGMJf3vP7NrRp3wYocn/sygthwTN9sU0DF4KdEz3CCSbrgJQon
j84a6XY/Dd1Vv7E6Fi4kWwcDBGPdYfJaLegmLGfy0yV87b4e6+iPI14QS4SKvKwP
0zzWZxoQ5znG6ZsajttOFhRPZKc+1jO7FeXqIXmqhlPNZo6jzxcXaXvfe5O2HZir
NC+H3CUlRtxGel7Bq+ejyIF1zWGn13NpOOsZAm3zX5YheVZ/SC4nhORezHVcUyE1
n7Oy+HJSTd1GAyGllXViggklje+zkrjLmxO6Co5mhl1swULF1KoxF2gqeYTn6e24
R74TgKbWRx085eA1+4mL+PPVpJFw2z1ici1wrvW5sFtX2VBen6VykInGq6UdFAUt
RaidICAoBoCiUw6O4ZjQdZDDPVGNdKnTXUMBCBaTtKfz7L193rxww6ALEzs7vgYB
vOAelOLgboWJSh3Eeo3rX+BxYViatIyyKGKpisK3awH3UNaqKPmEBzUGFb6malxN
w/VxMU6e/Z00TWYv3wKbQcYaCovH1jQcGGi69kyOJ54rSJOrTGXnJBM+XA8Zht0f
PYQlWEYS8/9iZxMGZ/OifnM0s7R3cmJy4YsfW5fJEkWv53ZKEIDE8YxN4TMm580x
TPSYhE0jWyV+afsbqcf9qRlPmG+hbN2+2yXUGeRtdp0wjSAKBEiwv72ZodPD84xn
rhnMX0g11uCx26GNGrLtilcTF9lUs7JkF+nUKztF9Gfc5EzkMFHwQVkB+AetpN+U
erYWsWs8EeoqI4vpKf3UmO4RkrUOd/Uw5PnAi4Lv7aaymTTebXvu0Kli6BXsVheH
Jhr6x/G0bZPcndnrMlKdGW1V1Dx6SUnlOshheIMB5XhcxbjNTzMGzYxayHarV9pg
2XSTVDAuoi72X4LxkhbhS1VxDEh1Qv8zxc1jl4pFwzWOQCyUvSFfy9MrwAZRqNlK
5N2ogMDP1cCu+QHGMV3Bg0ltttHxNPHmMAYsyWy+SDBDppEiJUm1BBGFcRBBc6My
jSIYij6tUu3sBdpmFEoo1YZCHizzk3a7fCNLtGXz7AI2N8cxsXlFOyLcp57Ob2Vw
SIbTbFyuLGTqr75ppfcKRYOL4ZZVebTjI9OpdpAidDrlC0SDLDvtjB/E12ALDh2U
nEzYzqe6ie4ogTIQKNTsalGow3cjLinvXTBPZWG8pPol1rc9o3awkaK1VkEF44nm
OKUNA22/ebTcFlCJErFGBexKop+sACXu4q+S6DD9qNStlcQvYWUjsxT1NNFC12Go
Uf7Crx0D9grxwXKkK8JJpWa5Sq8sYbI/oi8I8D+vj3GxgNI7Gk/0ogkZ7sq6XRJn
rVru2sqXVsd3Nwm9YEYRlwpkm51igyoHLfInkV3Wq1jHrDFk17lPazRdP1xCOUix
5Ntf8spKsMLmLD2lwg75BLqTUN96GXxA17zIfIIAZQ2pbJ0ZA6Pk6pHNEYHAgMV1
sXAaVY+O9OihjPnwlmv4tSTIrX4LzVQWukfUPNF4eOcEpWF6OjY+E2pI/XBxS9MT
/7ckKhLpYwNpq9qZidVgkTy6xLxyIBQOF9xAu+IMUl+XLvPNPhhvTEBJhvFqlLK8
Q6IxmzDF2Xtr6mytReQwjn85NWgcjj/5X9Is0XsFXqUJ96UC58JeS4g/pCDb5vpb
Dw7NmTuL1oWV/yRljQGOigVefxtg+BvGZnjpePA6FbMgpNd1OQ9zLOCmOfplTIsI
RZswNxiH2wC/tDRlJb2myvy7iIrQjE6J2KGLMn4SWgHk+b2sRlFYKGvYdwC7Cx6m
q07ic7nPXD9txyYOS0geuYjo1VIHcsde28JSbogMrKgyM5y/dX5nE4ViQOjs0dPw
P5UQCMZBcvr8pW5Wm2YzoebzD1giVUS3U9GLh8yGZ9FrsWkKImhW8SR+qWGmKZCf
8wcDLV/L9LYqOc3MSif+Pd/gDt9BsLB7RvQTaqG/rVhTAO3ZUmvrYj0PsQKFX5+L
MR+uK4QoPFWhAOcsDCLXZCS9KuMG9d9qQojYQwr3v+qzSNj0WImGPULlMqnmtEOk
/TY+zPoZS0LRgD6aZD4zgjyPzmH0KAdmZYvo/BBRK4NCl1oCW8zzchyfngFBGo5t
VYgjukbPJnydLtKdJrBt//p4XI+en3lrDgrEylTVNhHUQAuvtNZUR01pyndN01nY
nhi75CoXriBDAoh2Ypo/NO6zjhukNQ62GXOUgxz4ek2gMsDNq437Xp2N2WY+D28S
sSPc3KuXHb75JwUfjatsHvM7QkgfZjex23qMV8QF62IU4M/wyQebFBeJTLflhyqf
CuHmwM/gdQji0Iqx/6IRq0MKjAx9ZAznGXzy7zisklfjpVNi+OCGgy9p/H/XE0z3
vN919IXF1ZCQmjgSMsIUXZ0pNRN/qKXj85wNlpew/D2n1Gh56uSnry2TMYoWyya+
ji2JYiQvIAQ8PgsUthyCwmgUxrxL9grAmA5dQdzCikpj75KzknfLNFnMA+Op1dtY
ztIl+m4C3Q8/mdX7bDSnWp55KIi8wSoVKw4hZVCfrrijgiYDUGaLClgiIzDR1Sfl
RaVm+pMvD+u+Y2S71NcqEWhwoTI5+A2AnhFs61uly37hUd1Q3cGh88gtfd6ctlmi
tIvk1ZjtVgqk0OUnGy8z6/z45K2JSFlQ/DmG70XaLITzBPZXai3b1qjJ58VVfK5b
4jzEEu4tGcgrEFLjmHYE85kbUnMPp5MThDT8gDCd4lmJ7Ms4B1iWCYrEMevFNeqV
D3LK8zOnTRCMzQ+s4gFHPg3tbZSVzX70iwC7HiGFc6x/2zViTrpzkR8Syzyek1YV
Le3Qoo+RPfUwsgKjVQ6wTDyAu2iebLxQsBomggRwInc9r7E1YGknaAwnMSRnSYEe
Tb6XQZGFJszyTUVJuurSWckAE7VyD20oUFUq6Pp7LJ5juRyw5MasBupPj/zKXdBz
ILCBvAJPRZhCYz+ZVcpzYgDNcI4H7m08mDONlU6Vo7U8SsRjVOiirgf+s8ctUwnR
aQL+qarXQMAnQ9Ue2v7aO1XAz00GecsHqIVY7kA+c/uW60Dt45V335UL2Kp1SH/r
aV9EY2J58GLJNunNhNPcyEFgXzcykEvd6TkO1YS/9zbxrfDCnKUWz/wLL83eVcXi
FFNOhU5ZiuTfzDzE1iDTTkVZT4xiDhGJTf11A0i+YGDHJjyywoNhPV4WjiqFmLqo
NgLkAh8c3UjYFsoLT0ZiehYrZ0NyyvUDjoJaWRP8ZYgZ/rkcX/j5JcrDh6SmJJ5u
9e0u0aWkw546T7p3PmLd/cOb9HGtxyRFCZXZeMnV3SdeIRFuJbNhl91mec+lqe4o
T0VLkUcQpC3SYtxqyfkrMzgZ/mROwjtHfgR+97wMVMlkU5FAjX1PA0FogH1jRT+g
dBnLp4cd0MxkY8LIp3+GNgofmuRYSHuFPB7lCptJg/BDFTFNBiTOYq47u0Ksf9eu
iuPuLO9dMamwMYCJUnOUXiyxNINsCicphCnJLKzUVcrFiIwTa90W+l25X1nRpNPT
Pv22zTA3IyF8iKnbMpD00Z6njyY4IljvpDEgpGLhzT6ubnLNhSasNIcOVJm5nDPc
dyOC7D7zSCGUuZ3BJZ1cnQL/qL5O2xMk/VjX8TylxPCxpv7dI4PlP1b37j8bYTid
GcoHaKIdLCUhcMB3QVdGI7DRkinHjJTU522TY1EQ5FtJaleLrFjuJ84r9GEE1ba9
s6irx9g+Cy0eMRsW+NNrmGRbYBdEqWnR+n9pveYqECn/VYmoT/sDABNtWe+5RFNv
ewM41zGuFMcm6I5SfTPa2xHedpOpDOo+mhj1nNImjF2ZNB/OmZ8x7xYX18JZRGSK
Z0qTz8dcriOvuUBt5KcscTx9sZRqq9yZPvU+twDD4DXyixSnSg1US/HUPBkRfOJq
G0gsR+7kLlJKASOZng45CJfSfQl2UtSWbodeZy33mtmTLzeO2iPyxTdmZGfa/vtJ
LwNBzIx7FCaXx2t8MSTvzPGPzK+hjgIZzQYDqaUjb5UlU7fUvZUpDpKKKUALpAso
JpBWjfZRwDzG9y25aqBmOp86aCogHuswIqlJibkF6BrNyPbv8DlQ77bugdKCrfop
myXesG1iALyoAlesVBD7+8zBjMRtUVT/N8wfVXb5GSYaov85RhzHVorH3o+UhtJJ
6rVsAP4Kbhd8tu99a1/54UfBBu3mBjh2lxDelhRLdl5plhxIY0KClO7kr1jUF/0f
rdFvshRbVVLqJILT3cbvwt6w48gCbxwCShdvLSUzLSHb+bvSaDrIjoJXr9q7yaAK
bK7Mayf2RT2nsvgLqOYo8biT6HNVuNq66DVZxQ4qT2sAqUN9GTPi/1ASLWkaQamv
FoaICMi6UcfSaPcrfd3OaLfcvfDHXrHyVmPEmnWpt6JLiSi9Ram3d2nfzwwLLMzS
oq//DYmoAEztp1gNBCUfD/PNAIJ4qf7sO+Q9wuqbGyGAi56eVWvTVyPQ24K3v/hJ
iF5Q1rV9qZL+xAVeh4LE0HDjs8txym2EWzFJl6uxjaS4q0UOgSfQhd+Ff/TCb3Mw
ojmZuipM0fLWnIIa/I0nH7ht4G8qkQXaucF8l/3FmlGqdWRYSXOHBsicSiQOMjHT
RJIvOXjZYvZVPsV3AsqhiKBiWueRZnQePCyJw+3yXpVVmhcf1oCGTIQyJqhjFcDL
cHs/Lq/6S2ooqqYpafAIylscC0KFfEX4UsIWeQVxaWL8WKSMY+dlzjuIMebt3JWN
A26aKS1+pwSO2voIUiPcDDeCBboiE9/XCQM5t35XNBv+CDu7S0utcH/2otVL8Msb
47XrdssvcGcr3SfiWUfRDXHnSG5ysUFlVXahrEzIpEwQtPsZKTVn333jghnxJT8O
6+KM2MVIpQmsxOmrx1EoIqOAFS4m8lUD6pkbpeRgvcqj4aCofyyuMRL7NEIhmGtU
xY429kY6zVUZpHozQX6BQ83nsKlO+qeBECjSOxsqdfr/nbA8BKIwE+1QYACVQ0xi
HThzodxF55CwkWiSKIvmjPhT91vZ8sRh0FlmRlACbmnq5td0BAyOKPFkJRXgRPZt
6ksW4gzBx7KphcsVtWgV9KhKGtiIpioGYvXbpdEM/CrEQubMw5vKGzMVdGlOrHws
4ln8YvZu11fK2JVmSZr8Fj1OyhNLq/fyK/ungBGHaXnmg/QDJkUwVVqsoeDsfT8q
n7xtgCJ/ccDJaTKroIJ6d1/1v2SfKomwhnA9xst84nng2lxm47C+WFwVIK11a3LR
LfDG2b006uz2v53z2AUKBI4x1XqrdLI/pYBy9RiRlMfOxvs0m6INgE87Yl60VR94
gZZyS1UHTInFp0prX/CwKWfjP3wPz+xk2DYyEOIMhfO08BLM1beKGN2sIrRrzLpd
akswtt2R+7A61U2pYO4IyuXLy3e2HbM5l3dzPBlFOzOKKEWVxb7u1tSiRjV0cyWv
PtfgNhgbMGG7/ohlEFHn5IfexAvtLhu5Q7SZHQ+9oSbNzKG1eNWO8CvFGBr/9SzN
WmNnjTpQVmuW5nDEzBxnXAZIzvIf4t5OeYh8PainSKFYMJn5fh/pwEPApOypeGMf
aB/rgEofF2hHmCs1mGFCGJOX/zGC6VFquGxUzpfL8T9Dfidnlq6+9X9YAkyydYSj
gH/69Poxw2KgL8fUmBs4bApq7jjFQpBJbGi0GD6l1Adf0litkOr+BdJI7w6+DOS0
dPpd0irtrUovHZX5wwiSb56XR+njiYPyx4u/sCquQ6YqHlk93wOX9QGnsD4AcSU2
xeDN1LY0tP5K/UUkbhQRQQ3BOjHlUqnrwVrt6ciQjfTZORksUP+BTgCsTMwttJ9r
dZaFFg7Y2oxJf1TUI3F26sKm8E1BQlpb5aK6J/+yxSGb8z3QqFLAva3Nlds5cU53
LA8Y0OvbnU0x0CMpA5xGxc1wGwJC62LXrpvUc10otytYnHkQb/VH/Ooh5tqqIrtx
SV4uXWmFi1lTVQVqnRXz+CiQ63PBI0DbJpKI0bTIK/i2wTzJJfylrd1OZRCehSsV
u9XSnreyK3y7V1pjODEml5ThaNzfr23JToNVG7m+vR7SheaAW87fxMMqjHe4WUqe
WcCGUODLxvGWX6DpoS/Nn2WNijqsIuu2ByLW9SviCrWVWjCN9u3Wt8YMd8mPaW2a
vRBgvYimo8yzO75V+DHrTwSlz1lTWzVmGv24NEkmnYpN8MTE+y0o4lp1leMA3K3j
XSiATFnHrJyEpLuhO9forFpfqyn+zvu9zVlr/vihcZg0xm2hM/LqN1QoWt0mQTbK
YPG6cDF3/14F8NXg24zGU7fU9BDjKS3vRqZnAkUe53nuTGW5jXWq/f9bei9fWxcr
VjEmRAqKjZjBYTSMMuIDyl8GsGycMexz1jXlVWGlbk2t1BKo5jIE1AtyiTwWc/IZ
uCJlgEfactsx516ky4rCoEFidmfeZPVPjeGfPEkp52Q5HF45huhNnmlQtCTCcIcD
gIA4eHuxo5PJ6SkjZUkatrNasFuQdBu8CnrsCzGzKtG1tXmarNKTQrA1ggzalkXp
NBFFa5cX0Npxw9eNo2Rjb2CRuehsb+7t4ZD3BKKp4EFsO5SgwLMhUB/OxbcJFmee
V0/AEP797wWoaUHHAOee0ZbuD1II8fIbxZm2liyWZI26VibgB4KvtQPSfpfofU6j
6LtugiW1YuQmD/B2fzOeBPTCru0DdQ762W1apTNN2XovQi2DtLbpC/qEoeUxArnm
kpvuTjx91ZekwNDltVgduF8nYtsaZ3rll7JxIg31Eh5RS1dpd7yB+Nt+kmalz1FQ
QobcfuKMBvY7fdGWNfduJ2GgI2fVtR6Jz4/4dxMAqhH/aw5kFZpj4OocEGF8+rQx
TM58oD5yHLEQMipCC0jtsxv5eR+kvYDXkLcqCdtp4f5c0YtytiBmG5uamwn6VmtM
t0EVLHQ+x++Y9xW2Jf1yT36qYsKcQGBhgoXhgEjXpvQhUYYGCr7a/lS1+quIAUMs
qchdMGq3k/fg4UoSn1kBKOVbCP+MXkPiM+q6uZGq/z7QydmEN8UGPjc5wmmyceAz
sTVft+w3m3d8eadTPK5pdHGP+trfdPL7TBUg3NQfBvNvge3KfY0X0SvBV9NJisgO
dDAs+uNlOClXiMczjO1Ary3fjU99ioGgBuwGwnW0FjYMiAyUJNvrPCOfv7h1ad0v
n1/dnHavDHmn1Gxh35Ro7tuNp6orDNpXNnhlGHFuIUwuZ5xAgibn4vYBZJQ6EIfk
Xp0WpttIwIDOqATUEmUNNnNWc2L8egKvPjDO/H/UX/s6eUdx2cDWeHVdbO8VIKa9
HvswPpvUT0NcrDv3wdpqWzBgO2h9Ga6qtqK97q8wk8SnjIRDWHRZ2Twtw8K2Rzib
h94GWoX2LMImIXO6mr9zsKSLsORBXDDjsnqexLizYeFs5fanzQ7FtZo9PSCJtqy+
FJ86/D+/ZuiNDbWOZQRlc6FAZabKmnwpGZjDuUDf/M7JBd5F0kbF94H0jOfgvoyk
dhaIoPchS0Ggm4xDi649zZMfxBAdO11rcWEUm58vP23URI9KUcjG5JDdqDFlK5AK
ogKajVAhsaVpoX6dgP5fqGO8rEcBfMu9AWJbBD/XrNlSeFNuY4dFfuca0lNaE+D8
omtcgmbHSQTzID5cfbYS0ZGgwCzOJ2NknFgow4lgusRvCQzhIj+CMQyOgNoCkgrv
aufLw8XfFJt2O1Y00tirVoIRdfqe0EIS67iHAmgW+QhIVL7m37Tf8ZABkOC+APvH
ajmFN4axafj5FI58M9Nu4pXSErcQstscCNiN1p5txS9Ea2hF7ozG5HMlIUF9Rvn6
sde6KVu3OefjYFmW7Irq1d61seeWhs0JXHJPOsT8GCPsNUcw3IjTKw+M6tzmjrZh
mWDRgDTCmDad+zIZBzoFabxWlfEuGxqSuWGHtcq21D7JymHm87zIWtpGnYtRV3um
b3Ewv9pVTaz94nE691uXXl1gKY7wZE+6DElULx32yCqOfjlralv3ZNT7Y+T6nUTJ
Lddo/8vWJsNSZcUxy7tXmVS/k1/oF+DkbYstp6eiuFjjkM4SjdzMQNRpW6WBWG4h
4vJJg+3C34SsFc08cnkuhHukbeEky0HBqKcDfvD97gaeD97JPTJFYzYQUWtbSqig
xOKS7WVfcd1b1sleUwiVfVLBlD+fAtEBAyInlrWevGj6yjczZOh7DxBJBr5AGrOc
aq8Nu+mc68qOjBwwcBbJ14H6IXNwstptoOFZNR4woa2AqV2IT9D2rYr3B73QH/LR
xa+vgDLUGdgXWIQ4POvD4MEz8/DUuAVst4w8A3CTsP8VU0zvH+K98JJP5S66bITY
tzKuOwX4rZQlT+S5povyBH7lHkYE/psIclQeWX4J3olE+9FwbDV4LHRK3j2EhMcb
86GAETdFJFg2eVimZvtqw6dM6ltKceGNYdi/Z8d2n5zbeaomwap8nVW8RdSNl+03
K3hv5rvgZKuKRf1NUGKzf0dU8nsYC71rHTIlpKW7c6kq1fZFDDrL+Txt1m6ncN4L
KQbUxp6zaYeBm0/UcunXka2FKOLYNBzsHKD9bymqQKgpbnmx67dRiOeBYltjcMxv
EwcJ3MyN+MSLn+Kre/reowar9n/c3BAG4JABh2wcjf4U1Z2CG7g+TKFIaBPc8Fki
S3Sm7QQ6RZgNr0+sWnHXpxJKSvSLt59EfZ4lL/9qeEIcJjQIbqAOxVNAzvsSiu2b
GBexk2Z2adNtqot424r5rB7V6gcs1o7FoKM9Ar5oUoGn6rmQiP6Pemn91+8o6gLF
wyNsRRIjmdzLiYsMJ/AcqW4R+W7BxKkDLjhQChZ43K9uxphveesGwgipUp0VhfbU
V0MXGjDgRX2T33+UMyDzAmLeqV9lngOo75K3D64U7o1cAAfGB8w/Mqwm2uKpajFd
+c+6sFuvkXXM5XGTFsbGiV5ody7JL+S1wFQtBUKuQAnXBe2Q+fR8cICOAcTNS1RZ
MXeUH43QaGALer4622zZXgNVBu4E37+GNgNWnAtk743Y3r1N74RNQjgzs/nurhB0
vfGTkQx3+AsOKIZv+IzpIHOEGe4HW9NlWpLPvzWKshQnWCMxyPGc9+n4xfN1/iX6
sD2He0cc13Evnw+O/Qtn8C19zx28z6ebBVY4wv2lnhQoVJZe7thApobIxn2UQ5eB
aALN5wzhdJ6thKV4M3QwJRr979JKT5MLTKQnoCDSBgoYCMIz2iOCXPm6srdf1wR/
A8WbdG6gbOUX97X3C52Dxcjg/x4MeYR7qDXAbqoc+QYVr5R0gnX8Qdkke6xsFRw5
HSqbIHTl0kB2ANH0n4p/E9Ke+KVPEcpS1+fH/qsp9W128OGKCJszHGxFohJM6SxE
JGeJFvs+XZaZ4BSamEKuP9nLcIcjo+CIBZ1HNVp8CdtSxOzgZ5Zhi22rt91DV2tq
hGE/7e5evjL5R6NJ2PVzWZdqbmTDytr0Gd6WFCvNmqOBvH9LYLNfL2r/DZmHU7ai
y0nqOLSmcSxJVoa5QDMI4/y3ra02mzKv7JXIdZdZ3uDweapHEhWeU6QxQhjXyO4T
e8E38eKt9QZ4vXyPDQJtw8OYqO0IL7MCW6f7oLuDKiS7owfo8Xq35jk9HOeyUOPu
e+h6qXsNljLKHsRQmACmz16H7wYzf1LPcTevpRV4JSSDg08sgvBEGqZxZs1HRBAw
JxZ3qG/HjyIrCMwLPGqKAa9GIybU3ukx9gF7iOoJtbM8A1cupbHXri1l5xQRTgcC
zPO9QWiZNUASZeVxbcXy87MI9T8bPLU92+kxpuBvfy2nbef74LZ6s/UGeIhj5z6t
hy8PgdQbPS/3z7Nb8L+csutVepPMs+UFgUSCyEs9UOTzU463RACD0Q6d+iR6qi/J
h5TjmXTsyDv/ICw6BXDO7QrpBdF1urESUOGgFDMnKotK3tQkB92W4WbuuF2gcl03
skR0P9UynPKgvJvga2WlZrstiW34EhsT1AU8FgyAbsDilXjdb3+70w2tOpgwYSus
jHRn/iPeMbnjx7GwDfWLwXUWPLx9hvR3RP8w8JRhYut3idkYEXWfw/r3sPJcaGdr
GMsUn7FHS5KI4HtgXQN2h6vGPaTlAsKRxPRzDkPT3X2NP/CSHdo5EiiPlmiZUDFm
9BTRQjA/GVvVu+FfkffOrzlk8dA8Slp8QDcsPpPIIOpBkSsDmO9LfZAzVl20qeqp
NQigy9K++OeONnuGkMbWmOPHch7Z39zvihJM5aFxX3UTJYR7It1RuTn103JhuoNw
Ql7p6UrT0eqACCXZGEnplsbl8ESP2IlTmySnUds7VO5GeZaV8WOxM1DK/aArirW+
MiHlZsBl5sPQ4x0UmWd1pa9NxJDgJy6+be2sLoxnWmF55nZqwcQ/9OjeHAmql8iH
CNYdrDUFWWdfA3T/mHHEsQt09NfwnZ5xb0vcjGWlca3wjwDZnL0BeN8Uo4piHvyS
KtfcMOwlJ2iboojxGg3QndV5whignGyo82u99xLiCi81xx3BZg9X2bw6Rj7paY0i
5RcDlDTQdNIBNJ5AHPedxBL4x1pua849IupGrWEZafctliy+ELPDHbKkNmuXOZyd
kiH6KvRQl3hTz8Cs0V3flE2zGBOB07CkpSgS6PmmG092fqWAFhzF17ONzAG9dlYI
058/NnhiunJr5xa3EN8Sisg3QH+qNDoyLqV69A2SHkA0p0ml7t6PujORS7Nes/kv
B81rByoSa5DdoQZDUjaDY5D/1y/7/DQBI3OpvShX5GjEVJKq5J9cwPmcMRNNyD5g
hbNaztX9fybrvS374UBD/g4XR8wfWMQFxf4wF7Fl+0vXfFmNOWLWqyftejwbiq0g
ZP1ReNp/FORezjVtvdJcZDTvU1pKDPSk8f/TdiEjum73PmalHsfyx7ayqQdPCCTM
lGBHmDqPZlyK33CqdbasMqwGbtm6qHZKXmHbQTsQBBPKeY1+Ouy5VUK/4JvjQOnW
zIXZWsteWlREa9YwYOwELuqb9ze2N9N9yMup3SQMFxeuk5MgYym1Joh8g7cgdpQD
tEGloC64Jn02IZEqkTdUQeCr20nndpbgc+UyzRheoWMvJtOT9zhxJhxZvs1yvqFi
jfERV9sZpZ9nnYO/tORiCSE5zm98AhA5zT2xCMpQynpdKemes9JMaij1rcR/946n
UKZV+hQ3VcO37/yedNkCxU8uzUSpIgoN2fs0MsvV2cshDyhZNIS7llPwSqbFYNpU
PO4IhwhmHeZPhbucrBS1Dw7+bS5AG0oKA2zAF5Lnl2lA+ZBKadZA1tyZAq/F0jwQ
WRgEzlRYENTGxixSMF3qYb+3Dtfj8MChSmB1o51THd0liwl+zeF//LPlcDCiX3dQ
/klB2QXtVZaKQz3BNfauyp1s0wvqOVdUMbMX9SarAmnW/8yiossDt7HrwAP41OLM
oDoM/xNsv6spVvnOtW06lkOnCkkYyM8x5gJrJPKgrM4axy3KOM/g9nzWSbmmediM
BCRLZKnkaZ0f8yxDVgHrF3/C/289kmaJREsHcpGQzLeI5s5ArT9EmZMLPF1+iuA8
otAItEyfYqws47i7I2h/ojiOc8ug6Pw+I7Ek1PKce9Zkzp+zL/tb0Nke8P6VzS/c
KKDw/5Twipdzav6kWlb0dYvbTQaSYBvclvyeY+fxxPkukdS4OcFijJcH79ylj1th
GlHApMDeM8pNfrBrBLYHqnz+zNKnT4QI7kL1XOJX8Sg/qMSlaqMpB56sBiWZWF8/
kFYbezwT4ZgsEN12ZEnEKk5g8SbX6E4Mj+q0obnKOI9h/eiUp3slfhZt/ASuVu/u
zo7/RUOIIeKA/5nPKefnBLfZK8C3JM1yinyA64gP9AWzSpa7QsB96DwoWicUdZxv
RUnzlFkPt5B9o+t+Loe5Y0Q2Ha6ZAk5YmUWyeT8iNYlb1y9Awcycm9tkUk2ckt25
bl5gzW9H6txpe8P9sCR5EA3iBBTnYhs8+W3dNs7siq4gVaKaDM6FQaAdAEZ/Te/4
LpSgG5AvbWSS5kTrzK6A7juF/ruNV21dgSTfTxSPfapbAdR4jTPKdBzFVVw4nHkK
AjsJH6qfgz6f5O0qEwgtNJ8NFuDJwbDmvhihCY+rfK02GpWbyDPg6uFDCchFe9Sj
QYLYSi2ciSi/Xeyh7Syg8RKETeM1huCWlMk+IzOLzSS38pgp5gkLJwf8tR6hvAsh
2Uu0hVg2z+bkPKSfpimQkHg96QUmBLRS8S/LtOO1Rqqdz607pqCEMk5x5TuuJcw/
lxhpS6Ae7AXVll3QWodVBEtdMBM2Qx+TN6915vAHKXHuosO2DwTjpf2L+ETWIsia
D8P+P31smSI3ar3ZrYbM3S6NuK3lCnwV3oN9Hy2Rt7b17HxjKMRDO+ryVUbBHVAP
AV14B/3xDa9T5QVuc290Sq3RapCsUgmrBLBZPA4nH17g+kwSXisvKN98QvrUqp8c
N6HAMUe2JYyiA7mOWeZvi4w+nUEkQO1oYoHn+fetP6q1VMp88tXAJKNTL6NIha1n
+P1z5WixEgr+22Ekab7qJNJW8/0lhLegwDJ1k5kaTuO9ar2l/IA4GktCQq32f2UJ
o94IZA+iyyRyje8AL5h+o9x+a2xHsW7idtYBRJg4OrZ7dSm6bctatNXiaU3TND0v
7Qh37cQ4kJsWjmzRHxrGkQQREIxUWgy11npEi3d9n1/l029/biUulgYDt6/CthLy
y2Hkvt7f+Y5ALKIeBj4LjmXqIC6argRzu8rym82tP5scSXhdluOa9G5GLA583F2P
L/yyUb2UEhI6Ov97zyrwvEBuzLsQ9SFWUuTHAfaMM9WJ1pU58nm4FTLpFfr+BlNJ
wP63Skp+t79veYZQ6ADxTWzJKtp43FT2IXmHG5JM9qlWEm5jTRB8HQDkE+s82GIO
IyyiMq4Pn76r7wlGYBpUoBmtYAtyFYsaatlumRNNMNa7xYYi7qLWROlPbb9bUkia
yUgBm8iHFg3sSBt/S/0cf3VGgVspX8RHOMTeOELu+0uRhEb2CZvf3gbrfYa8x29L
oNW6pO8Zp2RgsG6k2enx3vTH5It2WhFVUtGk6uAoWUMTSuPwcpItGopYkYs/RbSb
8swTaSOZuAcf7pJJ7fMxO0XG3SeSxE88VgJkelx9kbhRCB0NeMu67412+qHfBuo1
5dkNZxuC4vofy0MoXEJlGfbkTL/0mzPlL085FWwCU3O7aBglwrvlqK+WU400YDsk
fWbMARZVUp8zFccCpm2lMrPw87mY9ITqN1dViGQ2iTibS8s93zDPtv23qBkMQQ6D
MxvNPK02Mpy9SQUai4+H0t67027scuQxAkWMSKK41t7JkPtE7VtqVK+1jSW4fQQq
WNDAcckPxta32p+OY6jn+6dDilSP83lOvryuoeGfDr5Arz6dBQSMSoiakgyKER0M
kKzERkYDShH2+WfAlq6u3Rm8ODEPGhfo+cNtQXX00cLqG5n1+E39WQ79fPHln4EP
MjjLT4YkGoOvXihRksS0iekPbaqMCcknU4jCeEj+OPsj5et2xYeaqUAwk3VN8yOl
9bTbH+FvPnIS3z5RBqMTEFc1gBIyIT0rgu7Ci13dv+ZZx9ewiGX9XKyY6r+Q8ckN
8exP3HPjGdzpSxUWWD1naBEnxbMmigup7gQ/F+itGp3fqe7qbEQihN4ubHUnqcm+
u8gLG1/XDbYCtWEp401DSHzhJxwph9Q8Q8OCpd2yNs05y7jfoN6RkgX/BfFDHxQb
pgvzyjTH+pthEnnpbQ6Yra1VcxqBj5ZDot6OccKkxNgqVbmQ0jlGU/no6O1cOKMa
lApZwdYCaHHmwn1nLMDGxW6en9Ko1mRRWhJ8Rorwbr10/UMJ5xouBXsO3Vmdmer2
g8/a4Rb6BBSvplE/yxa4sbnbuFRaBFF9ZdP0rs//sZXJS+cS6p2AqtmudT9z9moT
4XWeyiCc0+NmWvxT+dWeYAD5KV00CurODHxC9G76uc3K1WTxlBS9Q9Zvz732FRfS
MPsDkWQeUQvjBUcrWrMoeDf3GMAAYIF5pvaG9n3T+uNwlTN+usnEfbAXGouAEUEF
wQcm7u4cxeZhIJOkoTDgCI+47XcgA7bBBOyx8JO1vwyJLjNHQV4MNE1adK0ypnwv
g64Oek8s/d51pxmwxR9Qm/L0SQRuUdSGI61JTYPIpMdCKPI2ci7HGb6IarIgtJ8e
0kmycT7ItGbbrwbARon78s6I+FEJbQnLvH6ocQpOHhbvxcLT4FiBlPzOse8evDu/
rHyHVYlsT7WUIygzAUNnc0xS0cAfvVyQGh3F5RzJxN7h+C6rfZ/U6PQbe+Rxiwg8
csc9f3pro857K6jMOXzU7xGmZ1TFP33k8Ggv9qSyjAl8CrLhbKCarICUxVZfj9qh
4JsWizC6caXmKnpGS2LGTPeJy/H5QOWVNSWx8lP9650JTMxFUfmTlE5csRC/Y1iN
tlPgTbu/sspKNelgQw+PuW1uOpKOUMrFNQbQTtEeL/sTkZVeXDGxKa9qg/Z5qrbR
zUQFCvyTd1GHMyKG23xeGCIrnHFln0+G2962OQS0NEeEYMqN9SFQ1/bN9y1ewXWk
yFJnCcfkRO/PgboL4rhOM62SDDOESaFL5deJOUO5DceWzWh+8Ea7rKnaz3Xg/PHl
YWr94WT44bE8v1+6fo8Qy1BZUfK8N+OyU+HtonZO0q6hvZyzqKMYkm8Ad7+5b4kG
+y4DS7n6pRnjJE/DRKc9VkQb87TUO3hJJXlGavLAyDMOTJAWyoLLT7odrPYjQShf
uM1O8Rd+PxIAwMti8nUPiKsc5G/l23D6zpv+oD8oMlM686VwzolYpSGZsiunPiNl
R99Y/uLl8LWU1f7bVTYoGTBoEVxuOYOtcqHyieJJsxyTxS7qNCrVf/Zm+Djkt4y6
YKAtiSWT1vOYTj25z2s1kxcO+frF8Thw6lgiPc3jkiV26Le9MHf6oYWRNTJ+H6pe
7ZCVxUsyvHQp0CChwJEBA9nUoCOR25hC4jlb6Nn9eN//yth51ILayNMmL1GbS0Bw
vDmFiX34r/ZbFH28BANqKb/QUrjfo9elUZoMJE1O4neiTNlRlGgpV9uQK57IP0B3
9SEJDNp6A1hTz7x9ytVnQoYeZ+oLHCLdUHs8JjxMTKboF6mLJbDu1FSSO8dvr2QL
O/+CMcjz3t7yxpmut1h18wmlqNqXSseGJBXurcxUmpTOADPzzpoFXUGgzMkTIOKg
HG2sM9VUwFJKVPLrT1JqYFTC3xosa2qydcBHxO7kvxbkdarzNk4SU1XO0ohFKRXG
5ME6R+giI1JAE43NEJpJelTpLZp1pDlvXOvkZun1UfL7GpxqW15IcAgLzr9/s3fl
6DzYUDNQCTovrWYBHJxN5IfSTDa4wFzL3Epm6Q9cYHnMxsTxKPRJNXZI3CVMrvnf
YY8V5QWDDdWfi+B7yge/zxuXxpefwxsrkL3XhFHu2nPZz9ul7n9Oz6ccnApDtmTO
YKWXXUu+8V5KmgFOuNvMxqHO7ychPjN6a1McXLWKA9U2MNxiRcVvFpKj+3oevqnw
qdVypRqdkzVZAG/8tuVTlIrMad7eYBhOGuPLb//zYL6uw5gJGFVafirNNm8owPEs
79CqA9W6jWFvlxa4HNotsXUqs8BRO3EKsNX28yj1YThxaaacg+yl53Muhq/qufsA
hPXBBqYHnGA0Gr+ARt597j0V1ekY1EB1dJJA/0z5hypViJmXQyc/hryjGE9GH50G
VydyAhCtLeHBbPjJGEFRWNsG+0npa44IxM7xjO87FvIY6e2njioZbJ2FGqH+UgMj
93wLBmIOq88koUErz0ntKz4kVdbjggis+dCgFB92j6PnYDdKc6TKDDP6FZLCHvzY
JTKph1oOWn0XtZw8sLp6OG0njhbdR2+CZ81ihaDY4Lo7Yn3jcZFW5WDEt9ASaqQ+
6rzkmm1p3nDIYGpMZHqMKjSPf7r9xxOdn2tRv242r5yD5Psn2r6e8ZTQD+W+RWvN
MDab0XS87FnBsCDMkkNg/ZWZQc5Kauh6+wPftMT8tAMtukWdvaxYSvr8vGIdTR6O
qk8miRlrdxDSaEcX3WW91qlUh8XZFcykpQat3p3IVFx/p87NOrjLWMScyNW2TlFI
63OanC/tmA9+gY4XzI5/VxVfFnAngFRHzdpyfHCxjKQIq/VzstlovkOlou6JL2wA
5wAGykEaZw4D/o2DxjlhzH1CaUfYIZDMHY9jjc0azT1bA2JZsc8hiUhRLrOdtAwe
7II/NWuGALu4ESI8i5Z+Cy1iqf4e6iVdI6o2IMSav8SUj5DIkicXXkJ0KIdeHJ4/
akcP4FiWpK3v/ZJsSXq+mIjHErbVxejH4zl9w1lnoNwxT8OCe1iOsUtVSraHdwEu
gTvqUeJIDy4dIjVDun40KgV5Hn287nID0lJqf0C1eg8lKFjvFqg+fVWeJNVbhJ1u
rra6Cha3mtRVRQkABJ3qmtc6nLpPDSyPO28XPWvXVUV2n/90jHl8avqYMFA/F7fY
W/l6AMEsDW+4WYaMSnURY3nivggN9ZYbqk58IVEnel/1LvioovlYcwK1tTLsaw6/
g4KcwZY7dJnbjUY85ZIi/QWyJU9D+n0IXNzWs/+QplDuqYzAkwbO0rqKw7KCHWh0
txScAlLjN6nWmv3MJkgSFgR2FkIvDCZGGfkA1S9eAbddVAfKR5ghO9ptDjnfHyee
+0NBEvJuqp5Eaq17Lfe630AYKRNJ4+hJY9UVbfnus6rgyQ4+B/GDEaNdRduvRXux
rH2nYNUAu+cGdaId+MMQbNI7N7e3e6j4Nz6hi8Mae6xYaJFXu9030BCH4EyU9Fi+
DDZI0ph3SLgQuCwf+5ROENuqNF9KyNj6Ch/CCE73Wcp27QbZshxcntQrda4j0/Ie
JFgNS8BwD1zY2INjrS33lNOBJDUoYdI5HY+rPBd+EwmTbOtegVNGVhRqFIiu0V4U
TI1xbID4ohgNp3NwOGzM1Ms+6qHRMdqdrrFwHVqVuNs0J0ZSNIduqzB96YOeZ6rL
p3n6mNpL+EGxjY0g97p5drDj6YP1FOSuAYpg1pKL49krU9mhb8g5H0FmpuN5SeuL
RkltI8i1XGFnETQok+iE+1ebKsyoFM7a2pwkymAu46umwg4CCgWNWA2FUrMoSxnT
PEs+h90YEaKzojnVDj9PBP8H2gJskl9ruBEpJgu1vmMauJ85AKacvPV1QcgzUjy7
FXVu7196VgtmBECfYNuykcKvm/Kwt//tjuBiFj46v+wfSLiHvJJeUCefrcx0ig99
RaawH3EnbYionVpE8JNBqHN7cpjAdy1CBsISYe0K0YjTjdzFGusd6SQI7Y7g2xUk
9QpRqGIAKZ1dA9XIhMfeHwHPXMsAk5tRXb/jODGwKuybyWCxPhpIpyztlvN/huTl
2rCZ5azT7L6vc9MeTsJUWYcK8U5j0xEk4Fg/VkDm+ZsK5Nl18F70ZSpZzBm0MslS
J2DnY7CS/ltB4gWTgYsSj7h0b2hA7yr4o3VnqZ4Lip66jeLclPX0/wzYGGf6zDo2
bue+Qb8O7agqLYI+z0+QHZTprepJEMR+O90AUENo3DbrEr25wwufeJHOfQspgRw5
p8e43jUMwJxUIXswrHBwf0Dg/APR4v/dBhHZlUgWsa87cUyJBiK0l1dSETWrEj+r
afAf0LjeIPqTWJLEICm7dz93c/WSFafPZfoV9Slh+tEAHEjzqTq1kXtCoiyWmpDk
SUseS/oiMBuROZm8EGpsivP/n+YX5cNa20S51ZxeaPpKeevWgvu/JU2FhrXs8jr6
mBBlg0kUVUetD3A5MpahP/6/C734ms2gkBy3Ig1haw90564/O/pttQO3QwzddO/Y
cU+AQ1hGnpev7GvDIs8ykQTXY9CHsPSfqEA7fSCgYBtHTb77NfP7FO+EHfcNiJIh
7qF1HdpIcNQwJ0SbecFBCBnz4TOszuy18fSeZRa3APzV0ggtgzn/QOMBdD3xBjh0
83rieAFXVjIEl38mibQWkm5bR5CVJNDnzXczFIvxKWwyV4U+ajTSx4OwnrFZg+HZ
sj9EF+bfON0zRwfU3FIhrNVLQsdC+JCGTwkK3HcnRBrC1vBzztfdD8e0YH3Qxx2k
HRKV/gCQ5G+kbUtbMn+79x9afxvK6p+cLTtP9C/me0T8Tef8WYDxT2QGxVMPZiku
YiaDbQ0cRNsjMbwasoG0cZCtQAF0EqkLncxoCMdFYLmdCA6tfBmT1r0+kqmfssXJ
o9sE+J+X+wBMLUTp5/qNLLegm2afLE+B4s/H3zwEI02CZA6GnOUttKzDH9vp5Y7Z
CuD0JFTlEBCuzT3o6fR76x2vBWSNxtNFLZ/KYrUu44pzTGoosjBLGe0cAL2C4l2B
g8bAN2XBH40qRJQ4Mel0m7kkFeOnQziv35jMoHWw/Vaghr/KS5qTttloHa8CjQ0u
4h5I8gTLSTGp0DVyPjfwWSx7GMpDHvw04Wdyq8ZokzSP5ZxbtivjrdEIMrI/EZgg
MkbAZ1zE63JlFoJaBSCMW+XFt2VBCsQwtpEgHkvXQqp96l/wu+u8PVRDuuM1Z3/L
0xe1Pl8d2a4NRy7/PlOJ8feHU5F6TBhcqXzCxrQvF2EDrWt0q4Nmy9hwJqsRHuDp
CJlVjSOovMchY4xw6wLQfDhBj+8ewgKb/wMWItFvofPJFPbfm73BqNfSkXtldJno
+FZyenlU77gSothpyQvRyPGLTGf5Q53rHY6+YsAH+fGOewhOTKBwKasFoE71JKN5
Bi07tp1bAnLzWY+e1yUey6xa7GUIipB/qb6tpe9x/UCy6i2jQqjuwFdOAvdXSQid
FcPA+gO5SuwbB5D5TurkbQ0QkYaF7ZYIVm9S6Ot1Kt4/3nIFVSfKuwDYYi2BG2DG
tkvPusD5T33aGrLFqUdaqqE+tnl1GCZk/xMbSTywJTXP96+b0SpoCKACrwQrfCOI
58A3zCQHnJrqXJ2OPfhV43wrqVwd5cc2E2mMYtVBhRBt7svYGN8p3DQytmg6ieAY
qnM+ZXZEr16KWrO/BJwDhgHnjKW0zoupP6CQdvwXmgQQ5HH4W4ef1W637Pkol7G9
8ycPjUaJ0bC9x9pukZgb0HGgIXF6X/loZNO+qiVGOuZPnQ8Ux98G5nqsJkMuacfW
QZnNYStymXJpQ0UQ9of60wixY0lgSrLkNS6irGVsnfoCX9il4Txv2bXBF1ZKHsHu
Cm/zJ5uBj/zf8c2ttTJR6rW0yHo3JJDpMOsI1r7rRoV9WqANgSduhh8z3pI27NDd
0RhGvmGTDT5l3g1xCpNYSsDTOXDtEehkHtRjC8QI3Zp9IhyEjsy9x79d5piHpLpu
THe5Corq4ETJ5MWyw9fX6p6XKtDgQow7jftxRoNCojSM0sm8dCR0SiaymITqC9mW
q0oYVITYwqppOU9N0RTT1b2yRTGK9p0/JLxlI7tpyGV1VXM6+JOTeEEgK5MlWhkD
p2ZCDtSTOjEenOW9WhuIhz/dMY0lpuVBxw3ahqa++h6zb0W77n3lUyQYW9Oo86gH
ETVQxBCj9qQ+eBTNSrx8EUYXYhnAmooO2vIO5FiS2lGyfk1bT5Vh4JWeMWaQPZO2
tMUpvwUK/tdBOt7LwLM98gTybBizLIQa/HkPIQnEGnnxXEY44A3VW1kIYkroll3O
dbDglN2lLgYFOr4gy0nW5ktZXmbd1KBubIsAjfLEBhdnMymW14zXJlSYnY4ewPKe
uHFL/yh6UKQ7f6hj3z9JNQ3kvn/BeGWe5nmRD2DUhYtWC51RnWVNabv8fQY6lzUC
sx8maKRi4cEbB6X9I/rHFYcTr8poULSfj0Dfr/8voMtv3/dBtH9lsKvBACVNoZ+u
Y6Bl5ianUFAG8vBskMgZzZAuZTIjLxZlGcWhkhFhhrZXVVu5ymBuzKs059TId+Yq
TNmVc7nSy3cUyD8XwsFI0enyl0LgFnaPToVoWVY+IrU90mIIu/s9ifBgPsSNeJTa
5gpKTHhTjxBJ5cvMICvP/VR727KtttPgAAsfdw+91KotXqVM23/0R/uX42XWuQpZ
mSZvRun8IPpCHKaB1R7fKw8EczaXYVUAHDJ7boFFKuo3DyAqgTggfA5D5QtWPeBS
82H+ea87VUV0oFnV2nQXtMcDhGVn51KG02bbVG+oU7AWbx75rUjR2yVLOHnZmoqZ
devdEJTuaeRh44oWGq0tZUUJt2qvhIVsrH0/cOqCuuqMMfEoplNaRwUR8DN+Avcv
mpzCH8iZr4odLg88iBXMxGSIXE/3HlPYRJV8HN6HyfxP4QN2XcZDi3i5hOHG+887
WpYZqwvn1BMYp+zfMSkF78bANpLqeD61namjJK5w/b0NISBfuV8WpB6ozqOzRAQL
cOmmeojBRxfILsKHnaGILlz/+ur49n4q/AnBoEiomPAC+xBI8lGfp6obViRznbL8
1k1e0gwyd7XAuYzERjDQAOgzMhA3VQurlC+MuTjJxTKwNGa15Dd3IOrPxBvixYYB
T3VgKkGrTqSVITDo5LANV9DMdoxa9xLA9fDgobO3q4dUlTZAo/GZIw+dz7e2u0wm
z7Nys2V2i/OiNMqYRdXhGBGFFtFWNBApeggoFXQ+MXYIGeaC9J0ZjCeF/2jmaR23
T6zKlqSZCRVKMmC8mB9UpO5DqmtB7xiLEi5jwwZAz4PNjyBRzJ4criR6hg9CwRIo
RIW4nfy7vg8nvmUEx5LItkc/mQwSBG/cD3b9HR3sBkJp5Q4mMFx/xikGGPNJa+1Q
uoLN0N3QUlvOPcdjsItQT2+tuC3tCtMjfleeoVTs2IQ74GK7LAoEpWSW8p6++ii/
56DBzL1ZUa0FWVXT9fiKRJYJttERQQJueIoG6Tutrcw9AMm9gZ1fqjXFzuo+ErBh
7fY9ryhfkfoUT/BHcHP70bPWMF/2t/1r/NpyIe0BbHYlOOnWiri9eGrfJYE7BZzW
DA7GAUZfUYM7pnPP5LIE+xeh1t3aKyGzwI1rDbqPBv2Fg2ObLX0WdEOdCKYz/gVk
zhZtO5/PpjwDWwu2rLnAJFCOgpKWPygW9NnkfxjX96veb6V770CszaW+NwzvJp+G
h2Mk7w+XuLg5nboHgiPQz9NjNq2LbH2Ro19kybFMuvuBA7Nvn/u9NpyqMtpgWac0
R+jqpRlnUcoKsw338SiwubGQmvexbgtrivfInK9g4myqIwXYPdNoN85onXtV3smk
Hju1u7l2AqtUHjXxh9BnGJO6DMhyf1dkpUTuzMPZhProuefnZSPiS0nqK+Dj+Jcy
x7tvGSI/S92yyeIhPkrWomjtVHexc8lErWakjy2tdRJs2NEOaiBKVhSzJ7zqfxuz
fGiBnfsn703uBdPH8f/DUGowhpXtw60Gzy9wWz0UBQMPx6k1OjjI8gsajwOEkUaz
GdzbdGKSiGHVto+smjX2UdsjVU4mcGCLWlROJOE5zHp9oWmN690hRSxx3R/PqqKP
o3erqI0XV9cDFEMbdfZySSSMcQ8LpF1GoohLN7etyndUUWA/QPpQUwPUFPuHLF9N
nCoPWlA3KbyiEHJme1hdm8EyLYdurDzakN/XpzFwHP6jaKNcb2APZyuO6STvsa2v
H4oBq6vN0rJXO1wek5HoU8h7TgFWSK6c/k5LGIRRg+dpVkLOD+0S6G0iSUeDhx+o
l37AgtLkIHmAsZIk/Ih3TF52OLE1KsavVZjLCPBEGLjl4KfEHwDFzN4JwZaQUp3j
250zCEaeDdeuvZtXd1LzZcXP9n+DBldgwqMkrbA+sdEEawtlEvgtXOz15WUlQdml
LkUiyNNevh4Lhey/5Tr4WS+n2YgulYVNAWH0vUHGCLr89lIjPHX2pM1g1w0K/CeO
9DCBLjznXVty24gPm5CSoHUlRCrllOEUZTJKCdVIkd+gQ04hUCnE23hLUiHq1KHh
k57pgGFxeTE8zotG0jGbGHaajCOS0w2VAi54hWSswnhOiUJZyIubdbBi9sJH3Bq0
Fq0tgmioxH0pX3ZfRtk9QyeyLpw8Np+izhQxEvWbXseP9qLE3MU378iiUZUBcrqe
rQwK8vXwOf5eAnKI/BTgYr8IV+Hii0mJOnn0kryleU+njF0CfjZHq3IkiZrF3Yzs
jEolWr2DVImBGvN6A2wJZCoSde6Dq/HlXITPOT8X87XiJvijT1LVPE1i+v9dJ18r
YmQh3Xeboj2XXTuiBMrmFjQEc7M5ivq30oQ02iMQII+ffn75U5kMyNccvbzFTw9S
CZnvesRbAvMDVtyI8l4HqSRFnv3HXJbfMQwEIaV61ps+upVwpKUYKKshP5Sp3npd
Q60HxjPkq++Bm27BQioANSjzNKc7bc2b3L72Y8fDXGyWPrzqwu6QqWN/79WTCiEc
qm3ZwQlnE8A3jvq6hZbahq+TjNHErzTVMZan4fKQp7R3zDbtwYsIY4Qn4k3wHrmF
Ve9GIBcHiW4VfpWP1H/QX/kQTiLJgQ3EQso7KQFAIYeLlooYR6m56fLvrxmm7zfB
fdcOhRT+/rqjEzsB+DA2ukRbaSRYphOh+nbL55EO+MD8klo8wumeRwUf4XhSSDnY
0AVxa3sQvuBsyDIUHW6B8h/VfHziGxUHwQ+6IXKJKolbomPJuXVk4hxp8TOi8R7D
/eeLwbSZ1ukj2/DGeU/DNXpkEh4IUVJn/lkp3zDoWM+/jVXvdJgk4L4H4P/l9kRw
nBCTbTNugqsUVe+D5WmxRjxVpmWwZBzvg1JfyCDmLrTtZzP1gH0uP79M8qRt3Oj8
V2QSBEOuI1gNo5vIxkgrPF2llB6rjy+CMDPVK6vhSLbPA9QZdNuIadLuxGtzVUMj
XSr045RuNxeEfTX1zzJeFRK2TyNrVv0c8ZL3dzNDUdTp4xM7P9cRIrkFQYdNfzab
RsfD8ty2Q2kP45fLQfjJ5FfPP3eyPQEbyIjT272sdj9d33rCttOp/aAInR8RBp+O
ZKPAwBktlmBfDfHhXqBg7XyxCqnWzpyzXtQs7jICUTMNJlxSbSSv5F0Cl0RrrWBr
EIsumms2LNoskBUP84Wkr3fMH73CUohtQYKBpJzHbVYWkRB7V15Pypwn6RE3EA3U
WCzpHjWguyJp3JAW+FFOo4pP6pZ8RQuLcjN3sYTbIjCNwjUWW2ZjFPTAVoiewJaB
U5FO4MT6ZpoVaACZVgi9D9svyejNWboaHKbZcXjA+Mz5phDo27OszdJYGjsSNz86
4wxwC9ifqbz+XGkLvx2dOe7xrhy9wup6LKO3g4S3d8c23prlGCwahO3Rw1kngNcJ
4BS6hQmaOQOB61PvqsrU1C5T31sxRqlmlqKtj626vB/F1cf7ZqZwLwAUGxVrGTe/
SMuddDJX15B7otgylX4H2Cm/WNGyJbns57+673N+vSbF4L1mkt6NIYmQfdryA1Nq
SwSxfAn5pSXF1hBnk8Zs1e5X4/jjiBRximMi8NlofrOZVh0gOW82WQiiCA+wwc6K
0PerwW1GIjQVvXsXrBuGBc+8to8d5CHpVs1gHJ7M0G7OE6/aUdP3zys695MBSYdg
dvk408Mg9Y6yZBWmuBS948j4nzzs4QSPZ4IDjyE8F6Hgf72GJuMKxXeOuvhp5ICe
9uVjH67AVSSk8cw1dZ1xhAhr4+SPuK+12EOmF0+Xr8QxXds5yKZLDU5lEXkZ31eo
ILX/juKiFaX0z02MKQIcTHZ6gkuT0VVJFFrXuKi+moYXfW4CVz3L+5qiRZA8FJCt
uMhpYE+uLmMNCLEV7mufBgdbBvkigItjeRvVfjUX4DqmN1UbwhuqZ0CgihLnbgyU
7ffqs9xLy47TTMmoC94GYzMv0VWnkinhsAFQ6no2DKFipfPB9wZ7eXjw+yi0fYdT
N207ADgm2gTpYrz8/Bf+b9kKv4L6azeC8Fmte7h99FpZTSnHOKFBzBaH7ooz4owv
MblMRue6ilPy32ca6PXE/7nCuzKuL3PkC/ueIWd0e6sXW8kDW7nZtjjyHXbgGKSy
FhujBRheCB6Oyy06ioqJ6h/hvIbfO73e1dcilm/Gcg52Ko3/lqQPEUhNPVlQBDRX
sLskXvMgwq5cnKky6SdYXJasZxYnxmz3jJMai/OLSmCG791vwQOaamv71rZ9EKA2
7u1Znk0ubOSJ8LimCdDQ3Jz/sElld/w1LBQfhxVZy1+bOie4CuIt9bgHWWIGApS5
Wa0SmnhYtvFuilC4F+CKJeDvcyHIXbcoIoZB7/S7n7umwS5VJovPXWINVvfmlcKa
WRZfWsEEjKyQkjA/aJh45wG6LUof5omFHpkJPoBAUiRjY7pVHQPrOTieJ8JMppVA
yFDuQ/7OL99496LAlOqTaxXGoV+/WNYRBl/fleoE+G2Txb9FvXHDD14VUpiXIL/Z
JcgGuwhojgPsFd3zC3kz0rpm2ZK/NTZudjoKHpuFjkmX9SYqM7tXmDsTO6ReZHAM
eemn6Fhyq0MlW6McxAbb+cdjis1Lpp7LgOu0htyYErbjF5OZxWePUcjyfGDJaUqU
AW6zpHaX+MqxVTsQKF7LkVsoN/VEaNxgVwBRA105vIbTcgGmJJfyk5kUGoE5cWEg
NF9RqxYPDSmYeNPmefy87rbF6zgN6l2kyDvN++0zzUyQ292FZf8WjPP8/kaWzIJ/
z9re6f/iu04u39DaOrvbQBbMDD/hLhE2mHoXW/mSZK9zY5QyKNsSPlaMyPz6XUAf
zGU7GrsrziY6n3JA6DraIxkYeeIqumiS0P02oBYqdTuUiNM2/xYapwadqkuN87Jd
rWA1vDcqv27RCxu+B0CT7tFdGv2vvRjfAHGriO8sMiv4hWmFb70xhHG9fx10SMfZ
TgK6WyB09S53h/F96l9GSEDvpd0iLVdwM5RyK7GzEJ1wDthwnnp+zOfmBjZqXsvI
2DsLaeTKZCRsk04pE+ooGzpsTpxFRkI0JIHp55MdZGx7RsH5Q9sZbJS/3EuOgxgc
I0Cj/V/CA4PusoMM8fgNF1TMNMW1OP37cAoopT5GRC++c8yuL87qfynQQSpeZoac
hhIorISb7Yl959MGSSDnclK02GomMQ/Y5aQO2NAfZUkqmXCcC1uXfyxR72yWJNbB
ca0/6Iqz/3sVkYv9dmMWZvY8HaTTRownyhjFPfcJ4wkDHV1SPk+twDJR4h0b/S4W
j26ByHCIGlJcc+EYxupLivX6E/zNJr3Y3qHEUsF/3xOyuNxfRbcXJ/vpg78UT0R9
GMkUNaRI1tj/hwsRj5Zcv/d0IBhQ7UrQxk8nyACmY8+3884vkQbn4pfDYdPtGw9f
uPhuH8Jel4b8f5wd6/TJi+HhextFRdeeLysh3H63o2DkRuuzanvrkILtBbhzHoLZ
H7JuKvKB6+Y5K/EbadjtlBwNJ86nvLqlKKdsxVce3kECLBZQ9+8GYvw8sYJdgmnI
TUcUR6j3b1t+4y09QVpX101pF4NaledmrxN06OXxsCxCGag1yrac9t6eUSxP9MI1
5q9wzV2di45a6aLLhj5qJHV/DPH0gRgI9vb3AxcJJP7pHO5qR1DkzG/RPllNqW/8
A6522ty5cKebUgKpWpQX8tC7kXRBUnLgNaEA0KOmFz0PI4eMz2mkYLZNttxIiCv1
rbQgvcFwyLpYf5ovTaAOLGqySOQ3KQzGADu1KDHyymCHUmG6DX17O38rg5D4zkIZ
b2ro3SyqN8ZCa0XP2Gq+tCh1MbYH3kmsGgqaLL6AcIUKghz6vaQqvKixeMZiuk55
JcpWzYVdxe5Exk2cSyvlXtAF+AEJLqXE1Q5VQNw6fTMgZBkIsPRfLxUGZT53wCuM
ff40LFdRGrD2zNEa2QWLhRPOVbUrcp7sQo5gVjQs43F8k5/2QtUEGCY1eLUMem7N
VIoiFs/3F5WzobYeGavo/dzyJhOfL8Oywcm4CQKzddb4LmXbOt/IsKyjWvZr5OOO
/BMhF0CyzSQ0X7lNcou0K827SqmiQ3Fc/+TWF2PKzdEKY/8Jvs+9bP4l9HOvudEg
gOo+lJLB8OSL+1CttNjkccVhxEcgbJ8lCMOLZB58O+Ivs0GgLdOZRrY4VU50xDH0
z2XFwwz6WmLO52wFQIgAQTOTm+88IijPKM+LEVpws3V6Bcgm56E/0pBVHVIB0DFV
Ua7hGKmSPU6Bzlg9dyrCISx07Og6fbqghhvN9pDkMdDhLsXsFO0m6qCohANKt6+e
+fB4Th9mYxuxCpgAWOe9JuDGRJAMRkHx2lkOfFvAPMbBQB3ZZBU2jbhqhm2mm8no
uhupmDEwZym4PUW5vVGnwpi7fjtsIbNoTqjhZ4YOui024OcC6JYz/LOyVoLyuhsF
ZIjLC/47mFeK3+eTFGkOekyYsuTn9nAJ1XqKAG7oIhs3k7eDr6pzuXzJh52U7RyE
aXZqTLyqtV/Se+z9vkKhvI4huyafSewIp98T/wggoq3fiYuFusZEUyiehSqHDnja
1G7AxgE8LJBzQafXPlCmik1VxkAEnSY4FbARxzF9oXbfc/7Pol7QEKcP5sHQuqBM
fhoyHngTz0tjRY5fzynbdUx5wM9VPE1DDcWZxRzBxYV83pZ10TjMOqOZWGg2UV6v
bUy8VWy5e6cjK0+eA+u4pZuaw/SX562bMwrWaI+w+5v2BvjjW/YghkaG1AhBqOe2
ukuncN9BAjSgqz5ysnRSCBMmP7+GdR3E4BibyrxEPpn9tWnBD23aBFzc3H1bTpa3
E5RNFOvpvLyEViLKy8VVx1hB3B/ldD3On5a+rNbFF8IUJdjV1xkw84dYncFL3via
VljlwfP2OSNEUDIQplf9Ma8Y3QAPf8F3WquN/1XIBMHhUWTQ21rD3ilqLBNxiAT5
0v1v5ivJQZ1HjTp3pDKO+fXsLmb4qpi7/n0xv6iFOPOuyNDNgOMohDhGG+c+VUlq
7lNsIPgK3eJiHChX1wHwKW1nZzQ+Wg7KmpHdoMM3tkQ5VSuTAm4QPijqp9lj2Ns8
HV/IOLlEtDjV+sShVlLO55ASJw94BuF8TAp79XkO6LdPZCWC11Ck47WAFqJzhZpv
pZh5a/iwiLF0khjYXiYxiBLydxHOqaD1xCm/VAhOJSvH1VaGC3bbxjD1K5avNSyJ
Pycu55qu2agvWMlpM/hWIAzYADbRBRfjJaeEvCclxEnyKSRODz9/6U07FeyrRl/q
oeI4qlEy6AyQ38DMnaaydXIYraE3y6Djz+sA8lkXbgE5DDxFEf3rYgbSddI2ZUWG
UeFCaVa0MIGOefU6Sqeb3AK/LIfGeiuOztHENtvu+z5XBjDArtLKV51TrqqX7BMK
nvvh4z9FDUC7fVLeS4XP8WQPLbkCdv5QujtQC+QYbwUu8SNBs6ayQSwzXzJXILQn
ZI0p54prsY+bO/qFEaitQGP21VhsYOg33ebtVD4C7r7aX4AtMvGiP6JLlykkB7wG
K1sqU1j1ay0aStChaUX+2PpkJwpzlzZOFohxJk8f708AjVC5VmwRRnZl+dFvh6ex
4QQUwheCaqKLKBOVQOTFjq08m2mQ1rOFEsZSuSs7uj6+66hqUTHnPq3OVAwlz0hg
XiS+wNcC3I5m0rW6dddB/KROvXHTFPGbndCvEe5HSsFH0d2eomcEMDDjrobf/Buz
aHwK37qyRiUkr9EUEZKmxqs9P44M29CQENmPGVueatu547roPo0ObZAoByYBOVqv
k5ULOZuTqcx0Th2CSYGR3xx8MFmXI3YLpI0q6C8vkNJdykzdBIHiRp7puhryPy3j
8PXrUTJt3lCl0AOAC+e+bu/7XypvCrb1tAryKx0M2MaDYpsbNuYf5repf+lvTAIC
3m43cWf7fjFVWtUUHhy0jvokDE+wiSgBnbCLR/SJg1q7ZFTcm/+suqURtjUWsJJ1
YfrtvrrDH5RHlsLa3mURIdhLa8wW5M9DAlnqKC07JMjEuNpQ/rPfja8D59HNtv73
gCWG41BTJis80euyeN6uuGWp0CvXevc0ojJUWdq7J2OjfQ1fgZIzSJkqmD08PzRu
V5s1QW9La2YFfZ/oBFkV645uMhbMyhArZy0zafeuFxbF0MUT/cEs+hJlhvklwzma
oz27Jqy97V17tpxdVFCYHTxctbZGT2ktDttK3NGcfuL+B3u0+s2/vIQz5hK8Bs13
Fq7QXDTtpISPItAWmjlb6h6ZzVaplO/k3ehZa+d2fA6S4gQ5c/jU7Nut57aSnCB6
6LimhTBCXFG4wOo3EVEstmfl2qDh//GPXj8WFQWBttZFwXB1Uzlmz6MeA3wRUxBV
a6aOOMf1IBBWq53o+wUeaN7VPJP3YqbQn/VLzWYqECOXqjJ6xYKOQ6V84mxW3esa
FQq2n4FXOLm7M/nI0xGJWfcFltIXVLCEmeWp/sMfjV0JsJ/vxH3DF78dIAv6KOVT
bvVMPiOzGOnYIug0HqFA+IJcTch0Z7MEiWHVwlBJ0PgA2RtuV9b25TK8c4GEhg+A
AGcKJF/vxx7kcijzXRtExIJ6/yaUkeRqC5dfbBzoTE4tNvoB/ZEM2y7wj2wkVUEA
qnrgCY5AOAKI9qiIWBsYsi51p+gOJ2CGQKRgOHbmsGmwZPhDXGhWBYdz5OStDeX8
H0G2HEhsrZUQ6HL3LPaeukWcywEh+QJq2Wu3wTnJJCWFcR53RMysG+lSk3pKGapO
hiYb4GfUB59RZRNg16vhFGLPb+qIt2Le+nonTUeehSQqXZNsRf7CuFiQvG9h6lHn
Z+Ii+HSucoKnpKNYUCjP5+cr/DpZkJICeMXQ7+sQTfIHzs+z8QVmJctpk4NYD+z7
Y9zjJMOtZgMk/MdWljTjk+iREJhHvFFHqAYpmH5t/RdFmdsFa36RgxHPcIhJ2yMk
zgtG4PnyeLKWn23UCfVPAIeH5b23GP3j5tOTcdx2hIux5XmxVlUZSQb47E+X3vm0
/HbUcuHBl5YkgvyrosCuE3UFLu8ZMcyKRkXIXAKBnUaSstLO7jx7zguiviu4iZpf
zVtm6ZJ0fxZicnemQhZRh4p1cK8SZYY/9LV76JBnwkBuGkhbE0B0ezlgBdmXlBJC
wbpQst/10lTGkIgq6AIW7H8DPpc2Pu44Ae6SXHX25cZlwzHsSPzMEg2WurJehBv2
mwgxR7ejY/ole3GLz36T3qJ93HGHVDs/3Ruda6TyEplgzP0/sv9Ux+HlB2mo8W5t
MjALl60nqglzzWrBTcNMt6xNB+eWUdh447Z8H/cEvYPbBouq4Z3xVleXxhwm+INE
JCwMXcav7Yt0tqbOIXRIdNk7+RhuaeGTz2BVHpzLka3wuiCQ3DwAqE9LdtUsdihQ
iEXxCD0elx2T13tRpzpxDvMjnj0q8CRSpE1Fuevg+1UAtF1fXmTC1RBwN5tDJLgW
Cgd7V0AjV7AQwwy3nZ6TnboY4A1hZM6eVwhmu6C+35Yb6dGD9khUMAQ7rz1HD8jJ
gEdnMjJjsXOEkc5wiseRk/zVUr0kd+VgnLz/46KAQN7xoz73ZuUSxCrg6RL27pZz
R7K4GK+D1MVG6RDYpRG51Op4i6KMIt74PIS0b/fXL+iwFyfE7IRCTWU4YmjYypaZ
N/rlWcR4l7Z73RWaNP9nSiXGyPXOhjYpqDl2ECj1ksBs9S4eXl6SJj+0Aga+/Yc/
1WpOefXbTcOdxBs21s52njLutt6JVd1T/lpV52108phpmq0My3yw1trv4GV3qEjf
7E1rac2B9y/aFkYv4ykwg7/MtkzZczCD50x0S8qtPW6iMoIt35+zIcvnWSxx3365
TT0S3OeJNiA/O22VubT1R1ayV4texlceUUcCI+sF0ubEw9bInxtowWZx1jzaazP4
oaN3XOrb2GYremxoOlLx2JCvagxPo1YbG7zEn4dGBCNRL71vmlbCBEQyXxagTHjq
hzyl97A0qfMcbkppByfjUm9IkHNVhL7VEW6ZiOIEwPTB0UOCWbnu/SxtaXNIjVJb
4v8Jsa3eCOwMoFbZarsWtG8EstzdkvoEiDYf2WluKL6L9+ZIyXkgXUUq//kop99V
39CEbE9hg9Gdcp6ADqPwVCgwJ3LiK6iyW7aukW0AE6waqu0Xz28sUnV127WXwW0L
g+tziKQrtFclJQ8fRhSlD/MNxN3pDZRIrUzjjv2LRLXkhS7STu4UGG6Y6fMWw7j/
jWO110Hbo5lf9PdrMyTqOw92da4tsdARWW3asShw0ULJxgDisu7V6f8kPK1nCzx5
rVbSjwgnfoFXF6wbBNJJgQpEbEwH9mRTGtOOrHUzTOgQStnKTW2kNNQ0ygPczAkY
argvatHWXY5l12xQ2fYHYBT8yft79PcE2x6hFG81/yn6FtIX6peJ6xjMGIOtw9A+
K/5ulGjU6xRvk9/qrIUuyO16PDEyFmvL+Lw47aeT7G3Sjq+kbGa3wIkKIKqKV+Xd
Xm8aekrl2tPFmgIn8a12Jep6M7/JKyrI8RCjOpclB3T+LE55e8lfMfC+nU7ilKRb
GOeXWszhTSlF2YOJ1dO/egow2PQ5URmBwnyx0B2HAeQtqu0a0EWE/Kt3q5q+L+Gq
VtGJ4KMI6GPuzu1ljoZiFiqFeNMBJ7Q7sxVYHVVekxeKewXn2PdO61yDfizQ4VU6
XmJHuFwNWs03ZgN1n2nQQVxh6e08mggggIeBquMoBjwXlSkyEpVoDylnCgxLFdoT
XjkrlPNu7lA16tA9nhczknLQMDmduQsHjKQ0+BvGk8wJCbSYyrP89WsWpRBO/GfY
gJ4HXg3801wLwxns0+E1aLJEftSDNY0EpAC4qqKeAZ7dgGIk7lFSfAAjKbVKNYPE
5ErTII5vV+kie4cnQGullacgxF7+iHH1NjtNcs62e5WPmqbuNETCIEInXd36HN6I
SZdRI2cJxAhsC1NSeQSluSO7+swnvAPEQMsGFkkq/DAwXQqUTx5CTi3QULXPP+z0
iJt+JKgEVbUKwSCJU33jnkR3NNqBhBji6ij9ioVlfVmfViA4qfIBGULPTbVqNHar
G840PtqG8HC7gXGhXKeuT4igTA5R3vTddUZWWezVxjMo62VUmxa4bXOlCURD9lkl
OvU41M3WbDa9Q7+bK2jFBRKT1/BZzehnnZJ7qQhdTofMMIEgTOBYTgS96ZkOHleY
9ZdnEede0aWKaMcAbSbnOnjBrIriqejIOjGDEwC7cx3GKH8tL+tJcKL/KbJBDGHZ
H8KVMJWQWQ74CBbhu7YyAf8j8Esl/a4IgSepFz6lkyFIagUvHwNSLpgH6an3vJ4N
ujZHMdg3iOfFyx5k9Puqd/qSpl4jk9LwTQwpLhVHVgoU+d5uy733/UJpqcUfQkXo
cYG1MiyzwYFPH+6RWqkEQhaF7WdKZL26RaqF2wuBc2JaKTibwwbQegQM8OvQMbvB
ZvVd+tdRrJCMGPJI+B9TsfnMWSzVUz7U1JkHiqErMJBSxWw2nl5PSMXHx2uh/jGL
Jy7hX5x5QqYT7POuSPH8Q7mVziqMUbSL6Y2eGJELhdmBcTrzVkNJUfsmSZeHzCYe
6esiiAdqmkVAunTVGeybG5w2wfgTbaz262xKbqdiq6dOThfk1R147F6sgRGFpfnC
sKfIcjhFG0ziQ4b4SdU8ag4+FTlW+/6wGWIFdQeTkw/RJvBmohKYp3l1sORkGn1x
smZoaZdOQcqnhz77Of306MtGXMma+Hlm+G4T8S1WSX5gEYC6WPU0MCo74EVkRH96
FnTFvxHdA1K+qXcDkqMhMNoZqs4Y9M5K1HOFV1hU4qcmmWwXOrAFzDR0Fq0F7Ndc
T64GmjBHVvijldLCfoElr6pq6ImKB6naJcJ+u4hHZ+1JGmReOY2+ynvvT3t75BGb
H0SFMFH82tkORLmjZkOOVqLOvedELQxMXBo0Ztca0DCVdT1GJfUoSmcTj6ximhd1
PJI9iIRW19S65TjBP5X5fyBPv4jqfy9tOV4G6vslzkeAP4A9xbe/nbHKJ1AIcPKj
H3OrshmI0oA//01dFfZfMoSnrbW+kjvKJlXrWV5SR/9L4SWB9GTryV7yTN+LgGJL
vHgVVFm3lVoUMwisKdBg4lGJYouHE7F1VbB7/sFm20JqsEILXD9im/stuztD0Rac
/NmijFkvW0nT1Z/xpD0Enx876vBph02EfeI+TrSKk7uqGVZrd6TxRe2Zu1l1uVDb
1OTKH30jXP5IAXmgCmmMCjyz9Ee8w0R3Dp2ypBCurSxtAN1eIeAES71+LLR9b67B
Z7TwuIupgN1T6y6u8Y3mK3zpJiOfToep/Q0frIDrHV5U0qgkOkR3lbeX3YaRxYR0
4D6JgFjWY34xg8YoUsKirLRWvuoF8R5NMgn0GEeXQHygQppJSkz3lgkwLN/0HuI8
ftxvb0jCtTiTniwc1oRyFIB+aBRiPlaN6Cx5N6R/P2wE4QdBiIB0HCw2aT2qAAg5
X9TCyrGxwNa/qsykUZnv7WpvEZtSdQLl/pkJQrwtEYZfON6gRoI3HwVy3+2LQQwB
rOwPUGI/11UJc+YyuAkXJhuyLyCTAbz/Y3tKo14NvxHGYRPsmeVtcMwLU6B8NBRb
CET2fyIW/SQTu+hbiBB0Tv9ZVVhjJp1qi6uBRzKKuefdm7DNj3ExGmKDU+vFSMAi
yLq2IXMb2bXZf75Ns45XkDs35S2RpP7k5izOv360D0VjivfZD2cnetPLtk1ZaMUX
bVc1Uix22qa5RzismcxbeWJVuHTiFaBxbMfUFWeVXexovY+wcNpKQOHpmAeAnqhx
6qBiIri2yRptKgvX6XA4v7RvkdeCUeb4comgx18CFNwLKTREGLgldF/qTdsDY7to
k5GWmGaMpH71GfvSqICv2aLZn74Z3ATPLT0/s2b21qTgKPy1Eu77E/uar+Y2W04w
zZYgczxWYXuCKFhuiuyjE2b1BVNDkdzgztxaiwqlsSRlm5+zVs7/NfBMMNJf2Fpv
ncY4gPMzi3rU4FqFbuie0ZugtMuFrEBLHRbqzqdYy8iMnQnVRXf+ea19W+TvkcRD
HFRMQIM5fhTA+vL+K4FSC9YgI31ZKAjhElWXv/AJAMhjORicmsBl8Yrzv5ffkPyL
8kWmD4lfnVU279C9XYEgxq1NWRcEfeuEGdAsCb5RreK1ZoJG8VCqeGflBEhZv3Cf
dV10PvjZJdFrvPLZxWiDY9ZRF9CNhK70gDXcIGvSoMMGAi3+CIV+deNsQTAsxClh
YjEeGRiqZudvGfmjPhwVt2EHLfdiKiTaMeGTaGUoWf50voe+lEsiCZ5kwnpD2zSS
/lsVMhLJhMKt4MWMZtREEyzEwS0Lt2rXJRM5oevr2CSotsD55ChPJlmcTSekK3SU
hUiIHg/s/2cbso8FYXSQ2zRDJVi3+pGVNgB7uGgzPHO0ZdjeVR4cDt0pQXyOw94F
mqWeO+DTC9R3SKUtlcX7+DA5qteaMOEazlx3PWV/CxeDgGsNSnOCtsEVI38d/n7Q
kCL7E9WK/VLHcAPL/M1Zi8CNbtdW7OqjPeltJJf0HVg4m5EhPXfA64Dfsa3W7yZb
851Clrk7HjsgJt0wtmGFtKctoUVKSdJnuAn+zfEFN+6X8VclilWfu6qdNSl2flOq
gQ0g20uIjMdKwYrxCLGw01EHb595Ak+rZoQzz560ZZCtKMwRVJxSmcZO3Tt3CNUK
7WsL/xKsAA2dJuBr8Bgqc4prO0qwkBP15N8wFkrxR80xj6MRdjC0UlCSy03V1blG
iJU1plOH7/tlJU4ku2zGiYZrVd1F/CyVrAcjUf7Yt9rWjDzvTIXiJNN+T4oGcMNc
RpW6WT2WWFWjI65/vBnGCJM0SlHY56Xfe4SsOIF44scn8RX8Nr7VJSxXueHoWtsc
FanSPEaaHNQFfj8fawvxrrnEZrCylYBxIEStLIAbOZ46+lZbOnDR13aYoIYuMOVj
ArnX9u5lgeD0arSR/nW0Oox67Jna4zHsRc8UvVPCGZa/jQkfywBNJrdtACsdBL8K
jN7MMphKQWl4xXrgiYKDzHXn00zpfHm3SUCcdqCxIeTlLQu7jUAk9aaew28p+cS7
IDuZx9W6seG3HQfWhw7dQd5tw37R1s+gtn7TKOENuoSoPa6NN5rmdbR5268JSYxY
bpzs92vCjqBq6N1ZjhT78qPi7XTxdeUa0mfFpgo1NOSIc3v9KQYIPQEUqUJoYdYC
tSwaCcFjAiKIpZULYDZGY2C/Tij3pHJTEKDOsP/KlvyPDej9u8fJRtmMkkt42nvh
w0tbKujDzGde74VY6sv77WvMKpHP5t27h7pxPoNLObUuIaY+n1/etVBmNiOL8OX9
QYjAAZSZ9lx3a3+VXGrw9qEJGvydmRKZk7Xl9rqqi8sH51mR8jjkOWxXVK+S3trI
jLqggnFp+vtwaPpqJZC+oGFHU+xlNPu5uPT1Kc+Zjh0iRrrCFvB9qPWjqZirek2p
Hh/xXgggzEUE8Q1eoIuqJHP88PwbNJcJeLQwnhGAgwmIuv8Rgw5jExFrgazqC8rv
vuxoVJOPqkAEkBg+x18mkZQ43RowAxaxPunLVq4TKCy8U6CxPBooH2rrPz8sUsEC
VUpZ6Ncc492Wiz6uh5x7sxAUfQOLuCJKpY+0uZ7QhTu8fv37p7jGDjxLS5kqxuBZ
3muTO778DFwZAveQ3LJ7rsb/gsnVmrXqvzVQs3TtaVEK4aplrEjOXRsOWYR/Yr4p
ag0xTCX4mW0ClFD6Ims4jZGKNgAqsDb1IlzikVsR8NNykbEGdYjrrFbyjTaddXJs
Nk1Ef8oXsUm3qikXR9j2h1scJc20dtodSOmRjs545GNPr/J7tOT/MqB0HXzriXyX
hy9lPuWwwoE1rPBFRUs8WyQ/50TonG8bvcvubEHBozqdmCw8e3AkTUyU26rkvLTV
Vedmv5Tl7webxjwLiKkTyg57tqTfBDUD4tWWCzDE7V68q4LHoazD0AG8SWP+UZjA
hseCqRuF1peoTCS5aPC138M12Hi5plNTn/7hgNrctE5BHmdcoSldk/0Cpllhip7y
tHt7zKuI1ApHuqZupcpcARaazIe9cRsAAijK3YolcysW9PweYpHo8dzPtGcz3dIA
yBvDNhmppeQq9LhObPdmWOBSn5D44wXAQDH8XYXzJEiumMLh2Sd3nOaARy9D8PBI
efs415MOtBcs4x3vyEeN6uN2cYfdlbyKkj3xHEjiKqoHw5rfzkx1uLNSHGjwzlKy
jAOH9VHk62e4/n4LWDCZubRoks4iLkztJs1k2Xsbl1VsmvwvrX0rg3mXY7l12F3Y
BBhXpPA4CqxHodgiqedvJVr76AFmZAy9HOm+r8739Mw1OCC7n3ZdVh5Vb8LpunYf
j9ulEBF1DW6ZKx1Bk+e/xT2WaBre792FAi04LtBk/3BPBPlhEwno2vOTNfHzwirm
4r4uX1dPqYCMGURlTrNpu0VGajb3k/LpYxXrhR2Au2rO4mfoun02VlKyLPKMr/Za
2HT0P0Sk4FN/GNgCG8OxWSA/rhyOMVp6+xxz5JQsFhUBujE15ln0PRdw3ftQ3TNQ
YlFcAChjJ8U+qIVn6ER+8NGhoBPM81bO3mLSi0FDSPejMSaGSdj5DOjcfMarm9e0
fuj3r0LE9FcqC0v90Vp0Hv4j658QHpaoygw1f8yNbpc/zAQWJoNN4+wrO5F0O4H3
YJ733UfQT7k+pjqQqNEuvBgNL3slv7PfZZUL7mVyaEawq/IL0EyleHI2IhFiO+NA
eeQTnYEii4kSE+VO7f/I7geUS3LEJLpAloFagmy08W2RnUCYfC2AVc5A3mTLgrsN
DDdPkLyGZuWelh6NRSGl/bc0+isPvhr2puEyV+g7JUW7F2KEokn4cWV8V3kXQUfQ
gE1E9l/3RTTh6mOZYRwqORRK5OwhIn7h8uWAN3DphJ3AoxWSnn0PWP/INw2Vr+rw
LPwG0yjjmAh2Y4Qp3jzLyVuGvx/4/dDUjQxD9s8+B+7zjB4wAgzLFcukwLvkI5hm
4LY9Wme1NcXggPo4+r04/8tlkW4Rlj1UeE/zvAzpc618jB6+zcS/0JkHP7j/ejSG
XKhxeO89qEkdESva0Z6nIOYXLtemuUa+Ov8c1ouoJdOgb6meBVHOFAbuc7AyOa6e
+jVcWkID3r4QdYvdqI88Vt0zPbenSXB7wBxqKYnIwBSf8g2dNmyBTm24n24in0yf
KdlXadY91eno3zN0MCt4mKTm+mIYNhL0eXGP5WzODp7ekOJoHonNacMHNDBJaZUQ
EWCEEEbQPGlBNYq64MJrpLxT9LxrdzQTyy9HbuiqXF327xpko34DGuJQXvxqtms8
a/6Y2y+DhcDY62hISf5cCnHiPlPUa5W8sswNBnGRgjkjhLgk4+Y1yvnkjGDfjMxf
GLF72b3sMlOCkaacm69Ps7mONZu1FISU2EMcaiWQrYUL7MFwUJOJlahLUQhwVMgI
ndwbLJyPEUsUy43EDn16v/8z9D5tanWbY/qwwGUH6BVGEWCfx7aXrlWGyypzORPO
Y1VZ0MTd+eOe/pn29/hz27BLMDIDi1fQftnAOG8urCj8BAWluARMO47qgEwcAHP/
LWjhNHWXpa3xKemdqB4svoK4yekzh4ahkhSGslobeMSQqGUKSMuyAz3OJlkd7jeQ
S1uZuF8Z7rE/z7nt9wFKRPryGtOxOqd5b+rJycQk0SirWgVwIxHuFV0fJqd+L0X2
WQ7fNM1GlkX2LW478dS9LVVOZ7OgdgaO5/gWwUCz+NhB7DvVJHHcYWjhdQrtEcGG
JXIkJ14M3uYs2/l274gHgv97KEi0a9ivoEFhc7QBeckREvyyFHv+bNqLX4NyQ6ve
7iMxEfu4/5uy+E6y/Xdukbmqu2ljt9aiJNWFLe5LS18hJhBdrUeJpyZu3ZQq4Wvx
QcQ4ko/tvlIvbgM/Hjc26dXjBUNka/IUYdzMfE159w1ikJ0g1YteNKVo0aIuS480
x/WxCHtA3SrF/Pc4IN8KLhJ45MIs67vY8Dseg264Ug7mXAEoeuQZjZUJYS16Vk7H
N+2EEddJQj765Ac6QEavN4vsl1YsYtUtJjNs5tcwIoS7cP9ltvWePfaxLlcX8RK8
fi9M4bKLjr6jw3En9ZDXlmNLcnsMLAaujnK7SOcBfTC/EE1BE1W3aub87G6p9Ltn
SEa+Kwj1BMk8pIsM4Y9TixXA0ZtiuHuVEarED00ZCGklzhFMUhwkqNiO3d63dW8+
eHgJyxF12Mbad+dairIvOJtEompH0yptLlBpeD4uwtDE4pqxL8Fmgar/xhMN8oHv
ynNPG4KsZjw/TJpSMhxtXlxshpqXVb4pZk+n1FAtxApJeTS5rh5hAvenT2gFCWSL
Qz1otyoIqliraTOVTulk8Ytdop6Wr+bl56YG8dlDZnGG0UGogXPo+CDndnmnaUOu
+zlcvwXGv5/L0xPItKWiwXDpirRMdh6zfL9B5rkBFRWKM9xJ0eBDKI2YHox9QoYp
Cr9t0P6xNsjiN5laSiQMRrjINgArZtyO24dFAU1rSq1C9EfjeX4shsSDI4F0fkPK
dRxMTrWXEXBBjpIc6DcT46tVAU1D2aD3ppa2Bn6Zd18NrOVdEQKQIok26sc3HJ5p
tE7xTv2DO8einIqJ12Mgsbv2SQct9H2zOIdGQdHYRKwYwZccHWJiIvqeTT+OovoS
y8V3K1yVdA1vPQrY9Yg0LZMo9RW5LgmQ6pi91jp2m7CBQJVu5g+NQIyL+J22XzLn
3jh3qEjDEzlHoOaCqKYkynXfJZyCnN3f9TnmYAQOqoJD4gdThyjaX1FIAENtYDfJ
9qhZqoIO+8+UpbTOYIi5xkTTpLPLZn1vNp5HvWXgmlXT1O2PrMCRlbwy39tl4w4P
otzBOoOSFZ/ZCw9jtWyXw1Fgm9GBLQqGwZ+OY9isQpEjiqevraw5iLXcO9hhkxvU
51V6z86F3KYFNAedu/mLN2F1NTFPeqXDOF1z8E62Z6fgrkLOBvBgjZ9kOwyXAPJ6
NQHSF6IG9Ck9ikS/vMKTy6mDoYzmY93TJmdFEUxvhJWiz53E7ZppLxMHxCqSqvxf
Ox6CwWX8yS29xXlE0ScZBn6c8lnExTF3tXrEGYvFpeBcPkriMCGbXVDYacQrW4+2
gTUoPHnmr+qQ4v8QojtIE7rNBcbt6hMWeEUFJrBFEXP5c3pyyUE+8CMfy3npULrj
Jn+/ITeUtozJe0GHL9ko+P0Wk6RT+bQ07XL7F1lp5iFMo0Fbo8yoz9H1NwthYpEP
+XtyyPSBkT46hV3kRkfcy85Yx/y2TNJjhjQM3W3QR0jukwE6SHpVNpZdXzGWeVvr
IdDucfp6i8RA1b4VS+BflsAgxiN/Upzx7rfqffE+ViSfSBjjrsQbGCTAZvf05/sz
RRRHBbq7QjE9VGk/Kv9NMG5i0tNWN4350rc9jFM+8GVyoqkSg4jdGz+Ysaleu4t3
weQkjzyU9aFf5uqdOTRUstjuSZ2Kl56LG/y0jk7hJ79lJKUBXr8QBgNa1rF8WbQI
kLR7X5mNmztRKSyrt9pDtpOLDNNFhPulAteSyla0El4PYA+4xAT2b+e3TVkQBfVJ
+aleXbyBppFOPwIrx5DGkm4TVx4P3BFI14tsamymdMyaEN8R+30MswrJl/SFZzoo
FE0LTwlYdneTLjstHJYneNFN7bY/liLjStLcKkMstw1v9oAVhWdekyVlAfsYG+L8
Fz3t6PGVsCyGHoaoFgUj08JDos+AsncJtVc/6E2d6apXMgWg/9lBSQ4VXTpDVboT
a6AKhE+Zk8bXv7W3MRPli5guN1Z42t0eDap1CENZ4YQj1yg3OpOtzbnpOAmvJ4+N
iZ2OeFWr+E7iFhn4EKqa9Pq27n7gfjhsCExN+37VL2DD18kC0L4NTct7zOSHIrQs
vdNp4/07AUO/Y7Rt5uDRsezbr1lqSkuzvzdKoz0MqJiTThhtIw0wP5r/DGgNglHi
+BlquICNtoWaqaxsmEOIVmb5+2Rlk8sDVe1xsxsi1JJJciEJWR4vlolIAgVm2dMI
ZL/sBsmJx9x/eV/Qv9+DM3NVO93+NyBFc//tB5V7MGHcUVY72aSONNodtFuMIYDe
rxkGtVaplbTWWeFzZ/9oDzdiOU1Vp1XvtRdAX55LaUQm0z6iuCDiinIrWELI9I8a
3StATcbyib5F9H/BD8FXf1yPzeuD/ttVNmgh/w+GGvpcRuRE/wDimS86WOO84HnL
vxKftOSf0hrZLLR9mHNn/EX7sPBClEpNaYtRVgY5NRjuIoOuuz9a+wLYsk0jsZuz
OflQeNb/zxdxodHJZWPVqj4kIG7g+E1Pfc0TKTVOeirh8OvE6kjkbmskTEWIg93n
lo51HtKXIdmGLvvgSaX9GdD9zxiWb0eJtaNGizI8K5bn26drPVR9upNTYDwdvYce
yRoE5N02icAZfKVd9DcH0IbJDKGTg5oPEzuOImSFDIGReJgJtgqsAXuh/gCYxNPY
AWlLj18SYRqLzPX8GnkxncEys/K0SVKHQn03ZGuD8Nn7/GIlO2hKNh5dTo0z37fJ
mcIhVoYh6JJ02SfeHNbS7QzBKMFEmc9EcbzLkOuXatq4m3shAVrHvB8mORepihUv
Sr1ZS+fq35VuxGC6SIx+dHDG8GvZRGLkPpF3Uusfo96yWK3S2G1S9Kdt8p5vvYGm
ZmK34D/3WRyGxkGfUnfg366N9FTKc9pxGUWUvTY57+y96nsPBgkm7pc0Jn9zGliF
3bHwjXwR5x4a5BYjTavYjud9ahT0s+EnhCkGJJCS0f4D5XDFDU9QUdANixH7pvrl
Zwq33h2Rh1JLGGnWmCCM/lyr+V+AzqqqUehymL9PS3BwJCfm5aBmHXor5XP0Qk5e
p7mkdWfmpHVtEPYs5kosdbvMxvD2rWPMAgvHhtJDmUarGJXutbbVm2OYzAdg7EKk
pGp3MJ6WCmp6etMMJ+wF3ZQxZ5LF53V9rO8Fzhst5bbEEu5ykmrTchsHUmsKfFN1
ogF+74POTUGucU/B0JOk9OrBqu1pq7pk3kPrCNAJ6R7skU1dunVp1YM65NBqHMSU
Yg1bCKg2KNF7aaT8bhiOiYJ/XCNXdhWKShFoIFlrjiwxRY8zNM5u5o8N71Aq/4bT
CA7EPWZBHjsqV6wE6goKStmYCiNZuSX6XmganRa8LjsflNU3CLil65qbs/tk9rsa
7OKg+IRUOWXQpMCEMSNviUNX/7k4RrEFJuBSL/V6aKkzvxsjCFBCvL+ptpLe6C4x
pn+gzmotOiD7MuQ/QT5/cTDXqqJYcdnq5ozTB3fBJBi7DAJgdjYcGVcTJuyAHFaC
cTayrr/kK86bfhiIvy5l8DageWsPBiSdGekQ/IXc0zluFW8/g3OR51jSjQuMf9Gw
nIGEGwGWEhEZXpYAxfx9DYApFAE82HHuJgBSGWLXoBNI7BcRtMDyY0U1JfHB3Ouc
QlpHK3KGJD4z0OFdMr0VhMrFK2aCUW3gAGZhLankwdH0ualDZmUM1ReCyo+ZMLyS
5OixzIwmiOS9CB7E1VySTzMrjudWKUg3Ge7shLjXCKurDxntmAzMkhQ4N0abX3va
uPMylrtBaIcDGFg0o9g5ARkXb2FpJiaZ8KemsuUIpN7VA1e0NlNNuVLR0X8TeoBu
R7Cnwcra8CTE5pXKAWPZ8Y8UXIbcKPVgvrT5B9ytbqe/yRiI3ovV1pPEgfxxWniN
LHedQt9gXiqJRNsyOL17CIDQ3GhGNgs2k6l7J0jj0tlU2azpscs0NqbKzGXh6Jut
QO45ZhD5+WnasxtzoXjPpOK9BGZ+qDtytJMAgJlBdTxOMAVOjeeMeDy3t+d73Uw8
bRdLfxQZfaVVQ79SiQDIOFJkWEjdBBKrIQ/nWoyDltxEAPYC7+3sXy3IeHV+GKB5
MWM49UT+5HatOvkX+gf+QmSVYpQbyxHGr4gTqYvEGZ3sr4B3XsNb7tUwtnGQV/mp
yKQdOSdYlZHL9sQcm4pCS5SGCx9Dh8tuVRYR27phnOPKKnHebEqSsv7CgMvXBXoL
hSfBRlu0i8QTORNgHn4Ezw3CcMF8MWeVpWizcAZbqh6iJYfLn10qYMTRl4dVd0tS
vjSkwjFgy9KQWOOW7Ln0/D7hvrVlwqXDU0tufLraqZv1eArB5icBuG0cdkpBqghb
GkpbLVEoF/BrhGMWR4TSTKjL5ca7whAD/3pcvdOHfPjnjZjFwLp5IyikI+L9QmiS
pvp6EOsa9N1KysvRdZETfZg85thQLFSrnp4SjtygcZLiaQaTq37+CcIcnNwxzeZ6
pA/AnwgD7wdrlabQSi4Qt/XGzq7HzdQ5tHuJYDmDlmenEF3KWNBVuv/j0cvVReah
8EWjq/jJbzS1yZp8Vqkr0DUNK2K05wb+7Uqhljv0S9EC93XKDcjtHrFa5xWrrC1c
QDcxuGlB2gSLQFiuyEHydrUL3FJ5ZnZUzMVc33rF3EHvB4VNhgJcCU0dhfO0xlam
GQ8oMGuFZLw2Y3Kv9GDFUxP3GKBryozd63yb2D2kTd6cYg7NmnM375Njfngh1VOj
/FkPL8xazkwH1jh5AyWMlTJ4CzbY7Q3WzEb06YmHeZJSY7CCwFvd8IipEZ4E1CD6
vxSUIvucizq1N+Zy8iJkXsBN9s6fJh/r59zHJ7oGACuJzUgw1DGs1C3Zt1ZkvQp9
OU37d1o145kUTx2NWG1jnM7v04zh9iBiasXUVZLYpk8QVo25rUS4A2iV9VmIu7wz
YZsSUjzafaDtkYhwAbrJItPsMzGDrpocQ5o7gXvbeUXHyI0wJsKDkgZ2KKNp9C3K
DnyImGhJRYt2+Zr8LeUhRj3Vh6Z3c89a9TKp96quRIbf046vwJ8HP5XUZQNQXJaq
oKpPRDoSj3f5J6B3w5mQO0LFd6C/GiYX0THpeFZc5/CqnLJvR6i4YkVyfl7jyDgh
+mqHsdNnNdDRhKcogaROJcf5zh5S2b0O5WyodBMuKsQ/AW5MEjUtwNwKW8Khrk7M
chcdm4m+7ZQumcKBzKMXz6cd/8N84REviAqnfDswkwaWTqZaWWx+bO3tSENPslwS
FntloUE/civkE2T7CjTMWXZXY/yoycgJ3Tt/nOcBIcJu1OZ36LanFq83k65ImzT4
dXtQ5C3WFb/btk+GK4O5CxUZOq7bWZAAYxxXsRtsvf+X+kkx1ui+dByHQKWsPB5U
a/vbdWW3d1wtbR8vRlzs5F65Z8tJqbxLgCPPPBEduy+OfYMithgK9pGV/DfPNJ+v
xzeqGjJse4UAvywxrzQQp3cQ8KAc4IZfywurcM/jndkMzhpSRdRTOehQ1R+UOdoJ
CCwadDNdg30a2hO7/0mrMPFpinRbhMdrplI9GlThTkwgGhG/ahz9RjicL6Al04cH
DtuplVMcPQxmReTgcDjPHQ0K42jhq09bkQSw9DDaJgVYwgHOf11MQ7ngocno6Gee
OFIyz7Ik1iRMu0a7E5+6DhEgO7+liP9efCkq6/65jpbUOjEdR1Gxsiy7dcJabwfJ
fJTXoIAw97Ni/xhmeaPQl3rrlRH45F+NvZGLSJ+kSg3iosz6Nvfet/COZse9JVPI
H7n91NXEHhkdFzSto0y5x8uWX0celnv1FDjnpp9VweTkF5+JzNJZmhaI+Wv0fP9F
+6mwxlut4oG5kdPtOW5FP7lUeZk4r95sU0H75HwdgGj5LDs9n4DDqQt0iaXdY7DZ
11Yxm7xNl0SgV8YdlAcfao95ulQVErsZut1qloNxa3zkmbuMJGz7envTUMqEv0Rv
xaKjkIq2O1bskuO7GbatAP8YjoDct+7C8cGTIniIsvfopT1NFEFwaTTmuCNMYpz/
BCEmuQLUWfpMQgcDTODm/xO9FtMe2d7ajxvYoFkj5kCbfJlFLpF0qVrObrVNyw1s
gbS3vVDiToJqO6AtxpeG/dmUWmjQtzvVh+4endYe4aNugQCUm/6J/VNKP0knsnXF
OuR5GDdN5QUput+PtDHQU8qUAjboWpnWeV2/ygo6cKnfHlXN5Nhnj8dwEU/u7KSG
zhW2UiFhzuhbZGRInYQUi1fh4jpDpWfjkb6PUmL2d3VD35xzRDp/zVz3HDsplhuC
PBZ8iLmR9Tro+Wqh2kbh1yRWhW00FY4XAgLWl0uZUX/KSNYadZB5a9Sq4Q5rpEyZ
p4Az84QV32Vcx8GdXMEaOwgsjVtRh6QhxOG2bV6kyvRvdJh29g5QKf6WzuY2SlBm
upshkTMi7vh5D8WMNSVaTySfKQCHNpx6mo8opx4dTP+akPc7KVBCM7AmiwJQ3MIQ
GILa7kqtjZJUmQ4/YirlaaerUlfwJhjn1lWlYAxYvA4tQkvtYzTbIQcW6CLz8EU6
qs/ug5UYbj/LSgzmxVf5pRzTC2BX9r04VYq888vBPaJNKRaTGcAyPK0+ilq1d1jM
NIeV9tAQgW0JxTDCgFHC+dBsFCb4eWd7ko/8hVKZ1yrJvWugWFb1FyU8UOC0JkU2
Khq0zBbhcAAO0E4u1Sv/1sibA6W2qpNj2dseXyovDMWs535WZrOnJ3creSsFc6dv
CSiVfbqJhq8QighQZ50h8OzawwEl4TH7CGYn8u87AZwML6cncyUnV9WO99gd0RfG
CWDmmxM1nezCvy2XGch+fDCQGlWaQH/cawoBoyS/lB4Q0eWxeZ06bN1NFvCFvtKB
An/olPtSI1ORoBwZPUrb7ckmRKDSpd2zZZJUq6O8HDByrFD+azqKux3lqSsMpfoO
F53d6oUmD7DMIJwYqe72cpawwMKpMoGKSGUmPTqPyTa9UZm+3FZ0p3ZrcRMMrZjS
JKzqpR4mXm1vBzx3ENRVc10zOb/BZqd+6h5ayIAgYfDbORtPXFjCjWS7SOiM4ngo
zzbXaqNMO5XP7QHB+NTssdy4cBsZe7aRyBbB0FqUPMW2vSiOaHAwqjh2VotWCEuJ
6yBg0rHDJr3Za0FLURHeSRyPkRh94WgoQB+quhYf4bAIwVR0ft9MhIs9u2b2oxpj
h6GaJufBFjOx587w9Arik6EDtobPbtCbPbnhc+zSjcYevVzDn3YoRPlgfnfVzENr
Kn0aUpEpNVgDUldGwVHEL8d+q4eFsd8IcRO2LLI77yhSTqK07BmQJhW4EoG5sppB
/DZxOraAekU1ejr16DbdHSnmFWt7UBHdAX5T9/ZIJ2OrUxHX4Lg82hpAqxdN/O/o
J3flzzCBe2hIpYTDDrVMRY+YkZxrLUhhQdjH2bYLyp1zTJgr5LndVTeLpwn6wYVt
cproX6dZLTk3+v5q/ePcQgPmu//P8TOMDLF26mregFaQNg/H0UmAQKNaxYXS3CBF
rB/xmfjzO/QSO5ASexdHACHF0FGIM2Rb+iAwRygPM7yHvbJi8HYQ4GmZU9XysZEh
O3EO7QOq9BTnhAFPeH9OKf+uoFRM4PBcHHuix1QRKtIlIQ4QR57MakvYgsN+8J9H
QPLz86v/zFkJK2U4IKC159Z2TZsSWdJMDI6vGQI8P6IiCZlAKAQbzN3DPwDRLJGA
W3yUTqA37lgnhLzuQ0G8omAjkKoIHcbPNXwFPOjrw85WNbO4SooOt3WYwHXVWAQi
q4xsnQlp6KSyw+p/jZgBk3m7gtnYDzmuHcwPwY7dU7eNehuOi4xWMrP1obiahddR
q/6zmfKYX6OgW0cP142n+hgPMQ3Mn1LC0Cxkezfw5sj6KSXqpY12doHqI19+iQtS
nQI36uElbfyzCslmahjFWR0y6xko8De/VkVPs+BFoM8dGaFbtpU5O5NC0/zQUYeH
oZS1smIHLgsub1oeCx5bG7rihkHoabI3j61vR8l8HfMkdpdqhb8WnmCZt3vIevQf
qGcMGG0yCbU/GknbXKqxUBzTyoXSpDz2xJmcd7EECLp3vI6P/qXfeQ2TfK9mkmM+
V8pfor8ol6KqwY8hC0Bgy8JXvyebcODgxQQhQFiUmkLuB/BPnYKWu5HU9gOSu3pR
IhInhf3t10Cm4vPPySHt0ir4Nga3MelDXICMzx4LigXQ67IPXTVu6GU/Jc6lJT7L
qLcdYbszkHIo+VRrT28gLKYY9kuzhmp7w9fOOsvawUC0KIzn7L8l7MqGB4sK1c/Y
Pxrk9wqBbp1SFpZa2MTBUfdekyY10hYmKRWl2L9JznuG//oPGyHbgeHEqNGMXgmK
PD26saUSInsRGw5SegR32yoUJ758J2KeieebothRt+F+n/ipVIRb+zaF9yoFu0U/
/a31a15x64WYXRewSmkez5rSYY5an10wo8SiihFP3CdZEGqUxt1aa4riXavD6SZB
2o6YOdQ1GaJtwPdymjacnp/m0VTatOnyAikD/zREud6b/P6vtiNlZSAPFegH663k
jPcvcqXvVAocV89Jia4HDaE8Xgg1wAAY8rjdqqTQokxEqCtPeYc0vQP/5Hi44LCq
v6IYz5iJ3Wbozj44MPL4/EW+TfF8es8bdMyyh7QJYaNy+wCARVo+hGpgfUCeLcEr
OWUxeqjjndxmygJLxjCNPXm1FVwclmjx6QnnMkmBB3a8wT1hvhBVc1R7gnA5RfN3
+YHTWC72wBVAjCjAfpuTGu5VexASVwf6TwCODPcgUDYg+QkGeuSOF+iO+1bToPFk
5OTqv/57jGVrnLIMC0a6VWKAFQGh9FM+tSKv0PeDHtGJ61L8mWnMTTttyNwj63cb
xuUFmYmBFNMXoJp4kn345IjVeOFaFbediEOkkm1zPuIM5U1/9ZawZK7H2sIlx7jM
3zUgFjaocEl4RXtbB+E5dXNiVWqPaWADvjc9vz2wQCYMSjnd3s58IUzQbVfUs2n4
r7bl7RYfjzO632Pl6Bt1aAINqGK/HMVeeR5+9qn6OVkI3N+y44usMYOizG9a5ySz
y04k6se3wvsHAzsG3pbMo19WXwNwu6nXviK7IHYveUwK/yX1AbGdA1TygPS5xvX+
a4lab+BnAmroGnfjCLsj83cIWdu8W7t3IsRV3zmAMYDbtu28HG24GIfhgjGJaHti
WRQOeRhijeatflDL3Tx3oD1/yw2P2vdh+I2zFOd/kFRHLGFmQvgXxFs1kOU2xPQ1
42BZK6MHuhjw8XOQYOBSd87kzleq8k+ImPksVPpZNjjOB/TXloD8bvM2Ht8mCuMN
6haDltoyP4OqM7l057yIzvQCcy7NuNDA+cWn0DAfGeeCQkrNfSvNjRMYZhk8kEYx
7Tx2ihLxR0/N2SrbnPAkoXJ1bmHJ+iKqhSmbTu2dApNIeQHh8ybJCgRPJ0/2+3AC
M6EKJGti/zQwFMFBGWBUt9xxzvSe1hWfKE8tciwFJpPNeo8irRhbtoHujniwyLYS
nJH1KScQO32nFmQDLv8FBPF5uMKye8E9QLdezVhX1F0Bo2+/ePbFyk7tCbTgZ55N
zlbrw9uozetDveTXmbOhGY5PvGZNs4P0VbdTYddl5n+Bdrc3wyK/qVqOwh3xfbVn
HxhIEn1NvYn+1t/5jLPb0ulsDaKDnd0PPpXoNRIcF9feuDrn2ZwE2MwGNSPHgRyb
THO2lMH9t7vsvJ4iKJuJoj4yL73wrGM2qEQvx/fMEhZNOQDUoOd1OgrUhebf8xmy
TFGlwthCQocooL43iuNer1aUZPFaUa+xMpt80LIpFwBaiZgvXlrbM48JZlisVJIa
ECZSxbfmu/BVW1JDltO3nzg9JekXnVdkPWHb+fx7qWi0wouf06gCOTP/NGPQVf/e
fHzMqhGta3Y38gBYmkjjC4mzXnWpD3XXToPX3sDYLqBb20+oKLDaOSkE/2t3LrCV
XZMYCKO411e5R1a8CftCKCp+iwYcPlMYlQ6ap7mNjt+uuPSlVkX88T7syWlKOkYs
UPHpg42IODzk3cWRGixMWI0mZIOKbt7flBHS47lsJ7rLsd0GuxBL1VJitvXhYhQ9
FXueU27efV+08hGrrsyO0e2yOaW9B53YAI5vMEF0r6wSHFaRbDtx+K1CoTrJJi1Q
2YtRFuXADuixovFqN/xXpaiV7rI5oKw7BnC4OeTb9NqimHS9KuWvs14qcQ+azN43
N/sQD1urgBzfW3Fm7emAOWFpsxMWmwgJ9xOenRsbQo/Zzrz+G/IoQARPyzZP9JcA
+nwjNEicOFiDnVMyuN4BbxKUS+1Q4D0LzHzKcrSv/hs7KMFAmH6IjMetNIv7OTvc
oICvNIWmOA2ZhwLwMcll7W9wpPDTiHoYHffcbvQwhGUJYoBliHDXvzL5MZPO2Ed9
n99DgoOthmne778XFCoPAWAe3LBnIDHSwifTMiORyRd4eQRiIljWmvo1EzWUjjwF
xtEVnk3vziI+ZRbljSJKHJasCpqgy0rHrUSc4QoPQQ4CsR+usbdwk21TFDPuBpg4
11uq/G3eJBbBIJNrI+hKAj/3mp3bfjINxcgD+6UnS2733RAaph7dSqXysmVRHaFZ
BSy5QscHtqOuZ6hLwY6OfKc+IUwpS1h1Mv84r9kPzHv3t7hm1VjEnIcmZP07yVCd
9I3IXAKbyAqX/wUg5/IiW+Bb1JFVMqm0155M1CayOPV4tfemTBU/zsw1GggZRBtH
QhTDkDcwCi7FVmaMm+Z3aQ56z1cFEgG+FR5OeaKvHnnlsKgaGKNMIgiyFYSavq0J
MQeGoULRW2LvZCkCD88sL6gH7rMoMZOSloONCcDPxB3itVrmGKxI4uTVa/PUoHgd
pKKSZwn1O8eY0igMQ4JbRz4ZMIp5eJfCU6zDDEdGzu+fWzkaAKYun6Nq5Fo0g2ax
zJWrnZhBfsc8W5QbplTX8YO/0PbWme0dMtd8os2XPE00QM5KS3qs6S4aWHJQTQWi
w2qqmSAoLKT+OPnSy1bpqfPkskHpQTD1Yx4ZWhiFRE2vMYI9Yqf+RzxS19W7oEBp
eSBJvectnStgKW5PVEiiYgLCtHqxPE8lUnFuPgJStSsxbKKHm/sQ778rustO0fBo
3gwGJbyawYoli8AT5PTZ0xJrVHulgN82SBgtj6OacGNfnB2AUUeG5UKeWGVj/4yY
u54tne5YCTM0adBKEoOSuIXO+V3YIZCd/T6pqv5CDDl1ZwiUgcXosI1p3vonceNy
p7UJoGsiosUqCxWTLx8G9TLf5A1uBu5WForLKb8Nx/jOMjZ9+lTNiGKnm2JjRfAL
HfLTcoimh5s9PE8hu/srw36FM0abkgxmsGzacNHZtvHsUe5Ed7Z9VlJB4euY9GK8
LdPJGg0eTZbWi2bVGnOiPp6Q0njPIdJaprfEg8TBolgc12I2lbbKaimcHArNnRgb
Ld5BFFkZ6AWVLIQZEytW9jzlaY1w5NUBJKXlwM9VIo8Mvlt4Qui1aZnnLihlgD0M
oDDh9+hy2pWx3AHdmlLGBsJRqU0SrYQFpAce2KiW2/fdipp2u7Nio+2tXp2O5Tj4
snN66o3WETLeYOmOTUCQhlQo2DTs12g/XwTo5JEiZh1vfM/TKmzx34VpKCQpHUre
wwLRSogUK43cPLbIhMeRWojSnhh0e9SrptwSxhaRVQoWsGZXegHsc5i1+oayvCuH
TS8HRj4mswLfjm3ZHFMz5Z+Ea+G01kUl15sbpOHkyRyLMx+noFkVVErzPboibFEX
nJZrhIgYjq0ps+0Mx+8jRmC7wMUE6ldYPYRkeeHxgONlRkX4eY6Rq/0tj8GKaMtE
bAmzGepqNngaoRBQlQpndQw19rkKdo1MzBn5SbJ4+lPw/s0g42t1yz0jRBUHYi9v
EmRTA2Rjkrk1jR7LbMMZGnwcJ9p48Kj/35HapTLVdpp9o2zMowTYFoajDay4zgC3
sEpRsn4umgGmc3sALp12Psa1Xbm5h35kzNAYqoxk/4wPbA1JhwvIvRVrN2yeZZH+
TY3dAvOrZm7+IoPTCpP288UnCGIZpuiZAvGqGWpkKsXufoWYComNBHN+93ui/eBt
tKm+baK8iaJoh/G6dTLwzNSrC9yCCFxZGFB9bYKUicizOG41W0kGKyOSbGKS+AP2
B8zcAbs+dCDWPbIshAXJxKC6KhO+mizbi1KZpRb/t02sOp/qZ/hgzI1nkkN421mY
MFIy18UgMv0T62NaS+afhB649dZG9T8+jQ1uBikTEaplSSVJ0W1kuDgAnQsAoYRB
dMuz1e3oLVUSyldlMF9Hw8SvXrZvYRUtHGC3H+6dvRjsbKKI9onHNxuawxN1BdeV
01vaZ2UDmf0UsD18FmMH6yDyGu7PchFNlKEaSk8Eh3ETlpKsSGIQHuN6dQv81oWv
756jxduqKo/A/LhqftLp+CAz48mgGZFY2cl6cWog65Jzvqrlv95oP8wcEWV1gEGH
Pjlq5gNtPSlbTYvPH3/Y3RGuHP7bP29UStj+UKsOWExAHVdU0zs3IMJtZOJqBKHQ
3LPhjvsgeDFfy+56a5pn4ionnxj1MJAhzH4oiKCLhKi2hP4VPkSUs1R5kiHltCQn
j6fnzRVz0OqvD/bUDfDS8Ear/FDEMUXjWHRHjO5E+sqzuNQ7q9OS5ckmYE824ES0
pJViLkzzVUWQ2nbvNRisM9gquJoNS+EDqh65MCZKKsAGvRwbTxd0z3C4263GhJbK
c0OFKRZQKf8k3zkSFKnudLnRJ+zVA/035ZlInWSchXdoF2N4bH+Y+z0jMFbdUW9E
HEY+Clp+P8DC1CRobVYYjiD22++N5dnpNT9DRrzYRf6GiSIeW447ADH0WiFKEPtA
pBwUrRkQD1N4q56Hf1fvTfRVQEMy4Pn19Yx8H9NVOl7Zj4PVtjhApWdu4OsPt0Bd
L1wpzDsw4QtLxoV3SJUAqWcrrJ8Rx1aJI12xNik0euW6VxmwtXHN5A3dB5MkGWaG
6iDA0NhXKtvYOd0BQfK7dM2DlN05pegO1RXSQnsxHzwbH5n9SLLJdipDOqmXTmzF
IGNVloXCQR20eFPou7XXwbgMdlJrwxF7nVbxP0dps/vD4lbXkuM5mRvXIOmmmM+d
6xFTuuG9ddi3e8nP4IgHa6vI8Tr3ZUvkfpB3N/f7sReO8gt5+lM7ZHky4IJeUorL
8JNi0n7Rwhh+u1OxiHg6vAxJN6v1YmSVbea9opXh6Jlh3UcV6IKg0RFYQ2ceHDgX
SkHjPJE0MgdGdZ9v90uvV8ZMnFYAFQPTci/vP7AYzZdJivoZZW4MR7F8eLGZQkvd
x8FJpwRp449sPoI6pvFnaphnbzUEmbvCi4lqSdVVQdWsbO/aJcJOAIqBiKnk9/MZ
oAqaKea5km3h7Yb4T2ifuOl6bc+9PtpjJL8Tp3VqUWnVB0bcQoPRH1PyRRVL11mR
Pkk/fymn+hlrvmmEcqt4yaZaW1YTFFBnRxA8kpgaP7IOlSWWz9l5MBXH/QT+jHif
+dDOuRomde4F0Ak69oqtupkdwSXf6TOfD1RKm98RUajoDud/55+2AWR1gCY7eqPK
LEkxU2xdslEfqAKTigCYZpkcEVlRfLuUHGYjENAK6M/i1EHsBTsoyxB2P2gGDu7x
CQsQ79MHhgAL2ONaYYZzfxiX8ZW/csPxzrobvn9E3Mu41K7pcMaWaZ5jNCHLIHKW
1eA6sxi/n7ApG1Zyhhua29MxcfhuhYDr+w7isDlCvYOtA8xfTUsq7R2+rI/HUwP6
nOwTEh5D0qLg3n5ErSeCJesQd9qB2ySzH1ndlDjbmAGiEwaw98jwoWBt1iG8QQeA
lMTtBzAL7MTiUoQqdqiSUjNaWqPhfv/plI0AwU4nDacvABw6so9Gasa/5MpdMmsI
q8yG3BcboGLs9MGmS6IKQ5vCerKv78O57kfQmKEVrQblK2Rjgx+3pqOXz32ti45g
meKkR/KrGr3eNVcX9tt3mvfC7otNkfKJaxA5+nIBoENhFsymSKEkxZdv995krbE9
VorD5pmNWxzHCtMC73W9Q34tfveKTaZ+RhpuHrm0o+xMlndVyG4+06Xz9lbsF8jm
quXO9cy0LM9adrh96Gc/G+lOJk5Dx7DZJgLBpkM2EYaC5oVpL866jmh/C3RRYKn7
ua2ojyO6EiY0tYuVPzY8gcLovxy1iwkaxCZzF5+MduaN0D30ePwS3agdUhaRajmT
aOXq9RPDEu7rj6Vy4PnXDlMWtEs6F+wPs+8UBNDVslxY+daIhjJvPhHDckxDfrIC
++3rinFbm8ypwOUS4WgEf5dRSxzV+F8RXFE5lEKe/R158+L7N0Ni3/jBmYl+CGhj
l+gbAKDn3ZAje7KjTvG6up50FGh4958OSeDxnAu36eY+KSqOpncrom5TCxua+AmW
i4pH5Ggunm3o27jm6L/E9Fm4UlypjHqVMqk9AdZoAUksqln6vjAvw5X1SvSiJ2ER
aoLW5jPEgmQUjgeLFV7q99rtBDUBPqSn9hbdaTM5IAr7mgYtLubk33+CUVi/y75Z
g4vJgyTQZpR4g9Sn5PgZnwpSn5maxu/9sZAGvlK/C1Hfro2CyLfw9uH9Omd1aC/P
MDOHk1otCuSYDOlU4z/G54NnfUKwOawLeKglSXZb4Ulj55sMODVvSGytAhCPth7U
JsSShHOT/xIEh2+ROWL2g3HowblGi+N+ZkKYm6H8eE5f9/QhTU3ReozQzQp0+sA1
ldPqmayxvvUPjEmnCr4eP2jhCMpJEvHC+06m0k5jskLL8sS74QiRAsgAAkvvFlPi
YpWbcAWBintYKeM4s2ExdB3uNFGynmqCbqtTsi5g4yQMYW+K+bYmgQAbjW2Shpgr
CPpcXnhcGlrwC3m2LRApE+9VbP2y6uf8+OTweeazYK+vuIMZoFbrFus8GSkVbV9r
76iJn9nxlnR9OBNy8ZTanTA1hyBox/HR/Urq51PaIhvkGg1LCCmNmAz8Sh0I2WZb
7L2HQFGIhLS8BXLN0+/jlBbhBPfkBSDXohGEnnZqcOQsJYFfjIuNuI9x5xX3PVU1
tbBiT8eciGlvQSFMEeq6EYmO0PV25bF+KvgZI266Pncw26PmOGB9XWdb+MNB6niD
iQP5s5WTX9iuzCJ0Nizd92jhxjy1XqpTC3bMeGc7QARDnmdeuzQw3NHARIFAWAlO
LXGd2Zf2S4uiRwdPArJMgT4zfNgcxCU2Y0e83N3h0ELNUPTEVaw01Iqmp/mRgZhi
T0kiHQTbM9Ie8td8oqmVzGFjMXjIt7ZCiySD28/Thq74nxhF2Rn9giSaMsHF++I5
wT3ZqFaJf10BBg94FJGZWClc4H5d2cDRfdGP+FroQzfVvHG1Z2Vwrj3f2DGuQgn8
Iog6KF6JADAe6YXAMUmcEj3rP3V0nz7iX4Ce1WI0u5kmdXrtwu6rUrmmi3zBZ3oq
5Yjm2gML1Rwg6kGNXiUb7wfvSeuSM2IDXkFSmAZ6wOpn5UmIZ1vkzT1J8HEHzrfS
Yy3WvK4jTtvBDXsCbJfEqcof0lt2rINRFHNpVA18AzKOKOsqOgMwSOwHumH5kUiq
zZDRNIywVtiCY0Ed+7XUXoO5QbZM3YZyVQl9ktcBpEd4HfAAkkbEsuaBeLLcOhZw
rAZrph34VD0sSzw/Mky+1Rn1zaqXJKHpCH8+UVcU7n3ovCjGU88ETAzjUCeSph7x
A4N1Ym/trfovHcSbOFMWjslxZbq1T/hR93K0qdNsufd7rngUivLpaQyqP0KbXeft
2QG2SPY2oQQYk134fzppB8AegfFWphiiSVffds3qrJ32OGAB6/QnwFSUqfw5ym7a
Gkyn4xdaPqwQfZiaIHz331O446grvnOad5+i8bqCpcihAryb+QXZdhJ7GuTEQDy6
noMJnBNZy60Y61BD5BeFXpuJWBNF1jxL4gM0AVtFVVyimlRw6e7uP+1gF9OKCXsa
zr74slj3ZOyEvIb+8N8h/Sa7x34V8dSyeZBWUAP3Ph5/ZUDpkEXKIuIe3zMNqFtG
bgDB9spQFFQSXxfxVuVpAhE2scx8otNs1ppXKufApRdTjXu6hHmPdKPQTFFIzaUU
2lS6GvSzMbc1hxkRnlAFztzY0NWvlyN1YNZqn4VzLxs3eY0BIYZqygf7WREznfTQ
5XjMT5fLJk8QyVSo5t4W20v5acIZhHxb7vZDxo1ucSjAwkCsbsoGfXoy9g0MRN0K
kBGfK4t6V+VXiJ32eyFWkpZtRiGtS+u5N4q+HBLJDslxkyCxpMmtIH90FcAHTeW2
61RkD3j7XHc/gMHr0ezqHCS9rbSOv4eiLAu8dpz7f30irDVLv8Tsbnjjk43TjALn
ujpUWQol03nv8Y9Dz3RrLhDjNbYX1AdSKaDJE0KnyTaJmHEO2KqRkSFJea8U5CU2
SpzA8Rq7DNTso0qVg/4aGAGQTBEB0lTpsbR2wEdN5ob6Wo6DO72XxkP+Ck2/K3gw
6e1M9J3dtCiJ7rKyB+S9AWemhENxm07zh5+ueuoo+soQvcb/LEEcJxSEjlaTxuET
GTwh24fA25zFuyntCso5yDnyOBaAvSF167b9WC82MZe4aAhSEoSiOe/z3EjUgX2g
ix9Cqm6D3IHvcWPaQS2PUSQIBMNr/d6i4PcLp2wz4goWB6k76pjXBsTve+SQ5r62
cmV7vPYrYRK6SNkoiTxX9BDNa/k5sNQGHWUv3sxElsKciZC9Xetd8+G2rprzxo7+
U0mlfa21iOLtPMDrsUXuRXrrT63CCt2N6aQ1vlPa+hmCpRaoYOX3n9XCMGL3MfVV
FY8YOQDVEz7Raa4B2RcdFVoljd8eGDwZMZyPDhOz9g7jEjeJhSx/AI9hsGIRM0B1
jgfGV208OIRlqMcF7bUByOL+5KpAUL9kbJMetARAn8S7OOHyIxpe5zIzhMRWphv/
vYCxXIElHSVvtgEl3YLkRc1adK/R0XBDhJ/4Ek6Lj3d3xbLFcC1lrXzKZ3LNDVGx
oGCruJFrt4L+mnlt6tU1vPpscMSF/Xn/bViyaWDotyqFkT+Z2mwjgYc/X1G2vJgU
5bwZ2PJyheFhocm/4z5xOPapJnwxidV3edeFYJ48JjWoRLtBkgZ8hjtrRJHx7cyG
RhRUm5wWaU+A7wPOqY6NlCzE1W2Txd6Zs9w57KNCnFg4fGfS4byOZ/RLeN2jKdo8
iu+PPlWkJkuETN2B92isX9fLhSMV6oXOyjhzd/ptTqaWu/NflX6pO226KqtvF2uo
7Y9fBg77hHhD9ijrx/VmU8Jb3e6wMFJeY693IqX2xYsxyyxtJ9Otv3a5M6skWyAP
7Gs+BfbHj4fOuBjgKzQm9nLPBMLWzVaHm12I88AV/bBDL5W5j73uzIdaOkUIrPSb
NqK/Q5Cs404/nuUgcH4MPjrc6D5P5ExGQJLKdDJ/AfWdFdmWfpunsjhwlRh3hQum
L+fp8nm5vbGugEsmuZ3SRyU9YTwccnJntJO/NtUS589GvLy69J+b25lNN2sVITJ6
78pqnvxFnHU5UafsyEoK/2+oJr4JWJHlVjTOuqh/oSyN4yu39/dqu8iUnW8wJXOn
eYX4TSGCc2GJiib7ljCy6/5UAXjnr9OC02xDZK0EGHARhRWGydnGT8xc6s2YIzvC
OilCgtoTk85CdbctW32Ejbco3Dd9ewf11sbcwbCiYxgWBZ1xfsVRSHebx3PREkvA
hhipUBrQ7CI9YAJq6Ml1iWL3p0aDuXslEyntTdB7OT61lf9+0liXhGCFw/2JhVvt
K3SbkPb+C+cMp0qGDJ8dspmS5u7JTTJnAGzYbqDH1X0BOoKC7qJHaIP5kmkr+E8j
zG5t2molGqHHpsBrnuHedxA2qef8oe4oYdK1Ef7ztb6kugbxysFQLOUitcQ7U1O2
Sowg45amkpRTLHoQQQZ0r93mtK91lvWi0pEK/T/KLVSOwB4FIeDHy3dQEChlgOOb
hwcXU6oNVVOYTS/4kd/wIUR8W7CbtY9v3zH8MM+eXjZ+8zwaOdNiN4DNNWOJ5Mb6
EdTaOBMX7Z7Ly0watHWGVAr6RoOw/2VoeUF7Mke71YXx+qv19Q9zdfVs5i+BTr8s
NlXoK13nA1C1U4WzaoMoRWdX7miGlFflZ1cVm50Iu29h73UNd62w4O4bi6HB43dB
mA+GDzRW+h23et260xgbQ3jz+4jfCEot0DuA5uS/+xjNTZx5gzRXF7F/qcl5+fup
CpRGgHtA0XkIXWkFo4x9UjsZBGQuJu19IdLJFAVMY0Y2FHvTxLZdtJtjLJVRrybB
D5kjht9Xb9uPX3jN2pUwEx8g7vW1RLvX5kJNFFN2kqhVJdW3yONjwMZxVewUcG+G
wgSjEDE77dXeNay0CjDz4a5jO0qiUAHlIr6VWj0Fbh4jXiy9Pq1Hr5higBB86Mr6
ZLeRiSbupiMzSfUixQ7J+VYlkE6UHoDarkeO3mxwMOOv0zU41KAKdlzC8NmdPDNT
pN/TH5GxMf4blndJkNgNyGy29xXzLWtUZgToY97usG5nP8BA70kBwFPHY5PvfSZG
DIGjH81FQSDx+8M0PG2Xe8RtUYwx/hC7cQwGBjMYCD38FsLALqE/T+M1BlTDXRaY
AjvSmuBFu96mZQ/ZW+zetRmdc1i8Kd+wiuDnV0q2rxLbAPvAuKllg3GMcHKEipO+
9l637IVEHcImZtCS72zpxjKMzXajGWCDayGi5MxSW0haIWTMOGUWowgXfSnJUIPP
r6XYEqFtqYozvP8lm00ZA3Lx00IHVpzHZ9DTsT3bCCSamaY5fR+UIGL8sZ3GSNmk
Hz+bN1eXuFIIBxxVW7u5aqM4FGvvigK1u9m86PIkZudo9OqMc6fEH4G+b1DuGqmA
T7w/I+P+kc5bDOK6XH/GFtZ6KzJEhdOHkpjqDepkd4D7L59LdQYEsKj1uaxRUUI3
jC6NsF9+rL5pMHVuppZiXWuGq8QJfICK+6aFSDasOIC8ATNmlnIpcW6GEUVza7X3
b+X8FSabEsAlfLAbD71e7Ebrp40y4Y1VBM1ezxqgLXOHHdhx+bdUws4SFRUqXlp1
ASDLB1gCaDMWM914hH9w2cuULDM59gNfZFWutP+TSO3zjjPSaFuIzDbVrhPFPVJB
j4XGmofvvsLEtEJzz3o+5izy3XRRtmA8E6g6drJOaak+Jx08GPwVtTQIDwjih5bn
6JQdjMLDJd1OV0EGxYD73QhnAGzoYqrQ5w5Qt1qHcAmtrvidzdOOsFAwU2UkxfhN
9LX71VL/g9TXfuPMFiVixosPlx5SPt19Y0ywCthS4LYquVYG9l8Oidd1CKmr6uZM
lICiMTfDZDMVU4xZO+R+kABosatT4vrIzcairPXaS83y6IyhsEahcSSI6w0NeF73
XOSPe+e7xZw+Amg23mZ16xuBV/ZeH8HQekFHmEEheXF5c9CJQkpY/ibwj4piWpwo
rZRNYGfUgtj9stxmKt8MdqSRYM20Tv8oUCoSvBA0mti3h+VdjOQUBQ/EvtYjzz6L
c8FUnhDXwMMplZ5a+sizRIAyc4rTLMhk9Y4gWmdO4eRf0JPB82tX3Q3eTzNMvqU5
P5la2hZmVk3G2T77xiqJCfhmyV6Gur5qa3kzmCD2E+MFakC1/4C97Iw337o4/UUm
CMgkNCSorLnXbzj5IdewAARVooUxbOfr/3k3U9/vVyFewSr0CVtj1X0ungPtoLSb
NWsRjLoJr1vFhn4ik5VnHa2ELfA2G6vhyqLDn67vLJXZDCEWAcFtKW+O8Kca+T5v
ZOTrSnZNBAe7gEpsgX4gqIU4+alsOMhOheyoTo8BhrXjrgBBP/DNmvdp144obobt
E3OW7o9311YWZ7GTcZqVNPqyqW/UzxbEoN5dKXceXIcaIYHxCD6RrbSSnsPlzaiH
r822iu+k17N+RDSytDzfLcTjbhEdFhEUxpQ9yhNAmhptZu4PCAvKgA+CCXF8fDLH
nPdxzCJ+uqomACv5/IxlErBamEl5gtZ2XaHALA+H7wc3qgbpBa0x/GQrDnEJGOqW
U7OCJHDOCY1+OulpOklXedMUFzKd06X0yFhacCe9hLg4m6s8OMftY/ZhIiz15I1B
5pfbAjuXLPfA8THkUhVC2Ehydht9WB4IHS0P5IWUElRIDieARNrscSlV7eoWOlQn
1Nm1qmudCRxBDULN4KrXkkt+cUHpHKhGbe3rjxQOHT+351CBva8N8PcOhBVE937x
eSVY62cEpWvEUjI9TWO5Uw9N2SK7DBLUS1md7R/kAcz9E2hlNHd09l0KItTfvnzn
wNGt8DZNij0i1zmysx92kRNYfS8PJaAl5zf1o/Jc2OmDEv6IVtIkK9FUooD/5vtL
3iUnNqq/ngUuZko61DTG2YjWmoK+Ot7hFnfQ0CPQ+a/ty46dAg7lK3pzG7Nu7HLl
plceFFTPOvpAFO+Gh9qbot3RH7kv/YLDWBJrWDO4SRkdN4YeUhcddF1q1elVjNwz
jg0sUkRe/HsDlCcPx/hQxyJtG4Tq8cJGS86fUvcs4oXnDVwELbkdoPDhqdamXNKE
miTrDIkwyNPxlVR8xa6Ee43YB6lLi2nk7C5cR30q/unTIdkbr4sZtR5P1OEaqTz6
k3QtW85B01oxSGwBmtjHR6C/uSzIlieu0V4DB2WXtl4q4V+/9RMp5v768Ivjk74e
HqRJpGPnLgYfMsPEzFzG42g6aYy6Of99SanEK2+p2FVXgZBL8HMGZBGncfZcOhri
pTPspYYrPMZdYfBl2SkI3c/aWQlSxydCh8HsfisPjAKlot+RpIhnmps1zPRCbOjf
6Wj6QA9aSFCeNnSW80CjA5sctNV3AxhI5vCIDY1mLSlI7/zLOYCHKTGVZpqR4ZQG
MBGljcT9/I0Udf5Wc/IdmE1YIascBwUfZW8oXSfXUMCl1VPxPqXhvv4zZcYt2nGx
dHiH7ueaNOi049x/AUq7nnAqqfgdJg0Eoedw1FDx1+BaFkZoWpiqNVUKQH6N5g3s
pYbRM9ezefkaq6qWSzKdRs+vkf7PAeSAhqSXYm2z5/pvNsuhF/klPvSer4H7GSB5
1/L98Tnx0YvWk0cXfxLuqs1OyfZ1i+IeZUcgV0b2ruHGuP2y3xdzmvFjX9xPVSeS
fMLl8AkchjSa9jXEUHT293friTaezIhwADkvivRDSiu5NJBi/f6pyL1gYIxf6YJq
RaLNNpkRTlwKwlTZOACx/KPi+Vb5S6xTHqbN32RvIDnGGWZzgjxWazaJWX2Tz2YI
HIWVFIgqUe+UqcjBFianPuwuzXyGOgwzvFefY9RA8x0EHzQnLomAk/zsy14FJVHi
NxNjUgZ8Q0j88ivFEvKHiflDCCvTIz3eXElxoc6Xij6mL+6yOINivRs+E0uCBvBb
qHbER5XD2Twj+8IvJ/U8qsIPBg1MuUNGvTDszxe5A7+8T0pVg+YPuFU57hHWlYoP
R5aaldEJUiG983oMK7HcUWpzDn/MByz04ED82vOf8CJXwEEyw2NYfXX4xLmd/xnt
k7ygLwMmkoxN8eiT4XQqV+9fcwpjyKqHRO2sl+FHxHWiPpbP9acj8BULNOjlXLaA
cMkm3MZyEroWqcuILtoYWs+aSiwz2+LBKOzg9wgQntZsQk1VdC5OsifIS9xjGjf5
KkxMbeOi7nyvWD8vMc98xI4vzEMhLmIkGCo3ZmKsKpWFR27uAlgdA3jTPQgqoTOs
8euDHCA6nFjG8j155x01bO8YWux0yX3QZHOVxqIxH3huEmn7y8BJvna8ppNoe5v5
DkI087Hldg8EF/aNmVd0J6jb2TmtJoQ3ygJcX/bvVomyry674zd8Hx9FDcQzDkFK
Qyv1HXXFvhXOPvd3X0kP2/i3C4uABmyH0SWwens9UnzijpMVCmQnNwzPO8QKi0CO
88E+3oq+SW82Ll73pr6K7KmeL4+eSnazyfoe/vJtfhxiPfLC/eDHYSa0V2hMEIR2
WCB7+pipMEcKeAsjsC81YM9V5ZoHi5d30r3zYMpuYWitVBa2UpK/wdRFfFQCe64w
Nv08HpjHqAd58hnYcXhtM0rMjWP+q6gHIhFY5sDPhG0lVe4PqmcmgxhvcKI1P2t3
R0hn44zJTkHbV9fHwNJiYk+FbwY8+iXRmkYCN+dCxsj275jS/a7I0kjMeBpe1Cr/
KC2zSvfjHCRTLkY4cn7l9SCRQIqlJvsb2Fk+0b0PGbIkrOvXCxs5dNWe8VRnJUq5
A9tGknYIA/xx5MKS2YEA6jFkIQgym2w+NdobEkRwZDu5X+9rZAue6gFSK2QWhgIB
R8Gm3JfOpI0mR26Qpob7MuNt3hk8f7JEgEk1Sniue3opib7KHXacVee84mUcRAn+
Sbh/0JdneQG4s2+m74JgTAD8ZbI1fn2UO7bF5Dfxunq7i6EdIxCX5uAbAHFc5y1G
xKBrWwGBrm/JZZGS9Rmpu9ZkVsddN7XqnVbbVeWmQOL+ttkdBU9cFfx5Uu20U+/p
dy8tVu1QVJFkq8FGK4mtjY/eOGjqVaKy8Tnoj5boMYRLlbAolyJL1sxtNm1RFBCj
4v6GJHiWGOqXfYAIZYCfim4fZaCNYYh559DmN0ruPDxT/4Vk7mT5wXQntdq8YrHq
tei9wcAlx6iUQchNuCfUc57O6Sg2GdSEA8M690yCKmC0o3HCVBxIuHteITZVQBro
QIr1m+FWMgYqEiIHmVUsixGzUgroV2HTYeQdJDGr62t1CXMmKUsq6gZnz3PbHSKq
iDsHe+J7Zw79tpwIbwpn5kGcXYQdCiwYOYw8zAMizx2aAUyRKBYJAcSxzcj+MxIT
mC7XIbKxoaWUfI25F8W5ia2A84AgFAB/AuB6nVPxHdeGSC5pAHZAlGNsDO3s6gss
5TiGJXuBOOATWkotosUiQgrwTc70chTwtIKdz/UpFaQ9fvR2jUv01ikFc/MphVY4
Ud9+rn/i1VL19ib4EfAN2mcaADCYTKJjxYLWVFt1qwgyjxIA5Uxzmiw6+Dsp5Rrl
OBFowO3PEuzKw16h2wnOsCRMhJ3uAvJ2bywH/fc9vBhpig96G/VkAtGj1q9rqavh
IQ6K7Pu0gOQRrszl/8wgxg7k9MOlTu0zTwRXdpnaU1gp3n9RvtbtjFkKs9fHvndI
LO1ab5onGM0yK4SWYGwXc5zEG72RBbOkLEFkCabngxvSjfPXM4ZXcfEbFo20gWN6
teupgbK55l6lJsifFdgxpj/m5E7Zv8KOArh38mZPUJBtlHmBuU4OfAeY6BFSseLz
Jl0yfmffKplEyYLN6r5lRg82llujCY68y8R27kCUt0wWwGkHXuzvXwexyjvBVDBT
pPN7jGiW8tj7PxFNvNBssxmKwJOK7NzmDrd/w2IjRw1fZpDnHUo0xIIUv+DftRkr
6h5wQ0LJeUt4wW2Az351jlCqMSuGQuFuxK0/omns7hykpJVC66Q5nfCCjaLa4vf7
10A+xHFwhxVTOV4Y4qc7eNPj/zaoFgzPNIcvrPMJu3pVog4/ysz7qPhUlRpcwCxc
A3FoS8HAhRnRrETtcgebdicgspAAVPKy/hqCYbTPxl0lZvtkiH8BnGyiKkl26LQQ
kWPRbdey5gUlgJqq7du+A+o+C4bH5FnE77ioQtw7AJok0nryZIKLxJZ4ZswL7kx3
K7cW7SPHDJpl2sD1gXzV7WTSpL6bW+TSfjzx/tB1R9ChBn3UkjRyqtf45sEK1GuF
LNy6TmFj1rVJwO7yJqsIA/nz6JIVjQoPRM6YIgwQBtEhOLEEFWLeNTkyo4Cc0tsm
SdJOS/Jm/qhAXOl6SQ1LtQrfph9wzqOiCBD2tyR/xI9YH8Slgat/myIlJ/3oGe9D
zoaWeC8szH8A8nIUenOqqNs4upxpyrMz3EqRieFASLAEogKsozqgJmRzy7iqgU7a
OfZw9kwK898JH4VkMO5/uKL7LFAnaLNpj3QSuKRG7AiXlQOYLM9oRRvHRnLAJVIg
qygVblW/iApduU+kf3fLoAtEbagjsEGKxBUHtOQc3T4CorX1hOexnTLcitB8/U04
as6VkBbV53MqJ8LrzJjIby/Us2IrYWJtrxwn5FOwRxgpqqg9RmCwBThDOIBWwm30
v9Ce3tiEQINPpYXvUO0VWhwjF5WFgC2YP5BgZ247rBJ1TZj71/LZKCpoOJCMlrbQ
UbQrdevLebOi8N7mMAvbswWj0Hum0a2ZK+b4zugpZKNbE2rKvU0xz8sCyVBcUoer
gGHNjK2WUN6qrkvZM1WqCOTqsQQl7Lmsi3lV0ZPjTDeb1S5+9VNM2LjpHGRpdi2p
apLRKnsTikG6Qqoi86XrQhjoW40A61Q5Mc3lQBbZXrSqx+mpS1GyfwXJDGHXPIVs
jf19ntbUgFv+tLSsFocGaqZ/R9XIe3pXIdIlBltFzaTRb29OpeuaI643Ktj5ACPw
TL6Hcv12cIKLppXzoMoobEbElQfEKK3+dYbTxTixL2HCX5oPcIR7SuE+Hx91dEF1
8jkxo2us38kXRjxDI+QYTdHd7AXm2IfbbhquOegyDBhVgHeFfagbIaWWAspVyyvq
C5azhgToSzuSw5vHb41NMn1cQWQYVDGcFv+sJpaf/oT0DwC/W9uf99jip0s0CPCE
95bRjeOJwt9QZSxw8jRGu/SjOmM6xRbZMoLcbRGhR/Y3iW1cTLAPBDeF7kZJix3y
s5+OPiargdAj1jpOve7h6QKsmZY7gIAd7rp6O+gex/yBERm/0rP0qCI5OCOK/9cH
JpAIa4zqJSiaa0qeb6CAySA9PE+m2cevs41mgbKeWke/9R1OGwsSL9eN7x1eDDaU
4jPo0HZdjuqOu2/a+XhxxSk0Dmg5QMtS1vYS0CCfbbUc59YIzeJMb41HREVc741y
RikN5KGEsl2uV7H8Ctg40seuLMa0rKtmJ9fz2rXXol6q0aIFUvtwQ+/xC4EByhj+
z1rDyZjVO6anMDJoLnD+LR2Sgk8JE6Zd2dzKojbOo6PpIWlqjbmYre0hT7u1j48j
ukFb4jMGoWD4NM+M1opMfdmNCh2On6Ucy7eJDr4pZ6cCn6TCXVweGg0mZFqsa7S9
96xTSC8IYCnd0Zv+F97Jp9Lpt0ygvVkIAeoojrAdOOX9KmVwPc5pt0bVdsXUXXfj
vYehYZd7fYWJkhiJJKd5aVgSCbiEW8hNU4VeQuZaZAubj2GlB7bgRZReVDf+hSKM
jxpEcjntqiOgzD8S4YxZL/JNEonIC2bXnxdHv1s11C0jGM1kUPt3QANnzHbcw9gF
8z7PyLhn3OElnMHO9EIzQagMb+iixi67w8pzCcMoNQqi2fngZkusnZ5lYC2Y973m
4kcUsCW+2V+D34TZQEGg/2EoMLqLD4PRzC/EM/ENmoG3pSz5cTvY8oCY180q+qP3
SNpDkuG+Hm2Cd8zPO7j2JVG5lBkH4GlMhyteyEvvhpRShaGKlpaVok/WP/xtr6Ol
s96pDAjpuBsgciD9gKs5Ut2z+SxdZOzQoFWjasZaX/rVfMJuEkt6Mz79ZSO6KZ0h
s4Mih301FSledcnTpFldX3umPAjfCPSz0mgojUaJ+gwmdAWJdohILkWozcMNXwLy
daxAeFPs4bk8UPuzJTCUBGD6uV4ZAk95/GjOiFy1S00cNJlGWzsgOGOeFbFKsQrZ
nAgeq9g0tco9RLcE7qrxOd/0ZDSeLFysTE63MreKwl+N4uPPRfJTJXaqyVxIFtsx
zw27w3UUv3O6uYJtyOqBFZweiq9Znof9EuMGUxgCyVcVInhVpkLueOG3pyEipTIT
tjq3JR9ppbKmKHz7kbCnMxMjPHuErnmNwS/BKrcRgpO4pQIBvJZt4lXAqMn1/YhA
C0pDiOOKez06XEkbUnbxQj5M4HsjaIbRnGoQ6eT8fYXQzQJdzZ2/DzMIStNbyEko
gExv43TMUwFXbaKVWxnR71rHKw4/p+oPSf6zV6GcCpaGqbdQ1iZkgINmxjALWQCb
xdw3HkQ0Ie7+jvYUc8V0dYXihMeAmv7HI9OkAqaa97usoGn8S3wFApWkxEcIyzfs
PqwPlPyzwSh/AgigeVm/ulY1b0S6answl9n0fRgeEcuzMl/VLJOQ3iNThkKs3jg1
MgUUx2TgVgQfO+fS92LJnu0/TVdNB+GL6uQuUn5FeO/Boxh2pdjDkj50N6dBJaoT
h325m4EVwOT9kfwRn1zUOkpjxcqMtczbOI4YKoQoVjtWp6XgbQEVe0WH/Qsg6kho
rFruhRVFBThs9NXMqqCidPiN/js9lzDAMvmAkBIcV+lZ1f033Mb4pdDLsbYnQqzL
Jk+Wu2hy7aks8GLfrI7ftNbIrAXX1LspUrekht5JBNitXWaq4QxxBSajeknilah8
IuHQWr82xIBjGOZ997rel2Q/9BvaPfIq/iSOPFz3TBeLCADUQtmyi3CSCbJY0rgX
xwkekyb70ooGH0CSPRaV6SIvc1zvlsQewklOBkcu4fK+otKaYA8482xHqwQkj0Hg
ctqLqNbACcFo+LR2a9OSrewyRzBrQ6Ou7wNd/QASydzsXunV2NS2NMShFIPWfTVV
Kf2Tu3orEKlNZ2vsm02rjIEq/XXNX8k81jNb9lajTmyd2tm3zEftobaGyejhBqsC
JtxEXNyxIGGl8UpkiQb/Z4GoP0QUi5e98jnYQ7excnHbNBzRx0Ea448/43x5l+AI
/htscRtzzTyT0oTA8eJ81ypCDioSWlBslJmNZd92Rq9SnsOgljVjbKETYoe6yV6r
6AYX3W14PNzFZIDebKrbr4KgF6zZM56DoTAdPrOTaCEfJnFUwxJC9XtUOR+BGrj5
qeJ0PgfI6hceD1Qe30+b7jfXC6n4NmZFdsYeniokdVeW+Qyq98rI/HqHcOEzrCJ3
sXZBdKa7G/p1tpAZkvQuU0jd0I8wZ7WeI+H48w7Atkrktm1s+1WE/fppkird2JqH
LAhXAOKYy5sYSse25EyorzKLW/oOLZqMqwQqGwrt0RyD/3Q5AcTHD9dItNRv9/Gu
MeqKynJ1tf/b7joavIWbdSk4A40E1XEClLGtyUp/C+Fo3U8AWdH5zCXx6QkNRz7V
Kz/urFOtjn/TE4XGC8tFBo9KQFnLl41XzS0sUoNpfCyixIpWPqjADERVLtijgK3J
30hRkPR4xHcNh9gyrZ+WYWrxzTjyfS9KKOzMbrCosbd/5yqyYkSaKjgU39IFR4+L
Cd5XVAfUbm4ua1jc8sTz0iBnltW9npcf04sVLdQgH24zi6KZ20r6JJa4m90k5DI6
n552Ug12tq/D6VVHtyKEjHqLrfzWFMWJfQVE6YyDxeG71bNR6LXydkJoow2kZcw6
oCPs6UgP9j1aJX1isug0Ud3Rw7BddtH8pty0bQEzGMA0MqulOAMXzBFE7tomv5lM
o7JZ6UcFEUn9iakVEXvatjkruLPwcMsVp3c/Yd60ZhVQpW2KUr5+NzLWjcWmekXQ
D+A9uP0rBC1ac7yS0moWEYZBlxE3CKcIzin28HcClVzNRLuqPrrGmHiezbMm+l3c
//KY1mMMk6/yKQLf7dD67rHvb/pkTv4rxG7Wnfa0VOm8Sd3CGjfZ0PI9YWcSMLTB
UX2EBXE9+KCeyfNK/zjJrl1Y0V921stftxvRtMbE1hyfIGQ1MrNkUvNmIgck83b3
gCQZ6Kbv3mbjFdanpjFgxzCs4+cTjf9cGzzBXpeb/mtSlwGqV2OJX5jaTZbv/S0c
CVv6FOCnpuzWSGyGxvTE17Q28JkMucyqwQAD7DYmbJqbi7Y8Jb6bXOikC6nTBIva
k/G/tvC8+ehGlGrm/dPcHV5ZNvYJCNRdmjOAIovgAe8EY1PwjA7F0izh7+Zyfvh+
GBV/hLD+Kfi3oBUp6Tlzr9rcL3jd+2u39dafv1h+xD6p8opaJIEm6rpnmjHsBwcn
USxJFtxCaqu27ldQEy37iCAiKi4vE1CRJShRE0EPZfzmsPlDWvlsE2gPYLrjSu4J
+DDMQ8ruijDmaPv6J/en6GOIDW9chbs5jqj6gAvokDgd1558HG/7XS0xKyNfGLkm
kxxWhFR8yZPJd4yAhi2qbRzZNilj8svZwfmvAAvV21ttnpWFiVG7IkxWRzNpbkMB
IkXyDqnFRHkjtgUxcGvDWEIQcIupjuceFiKiAMkpec0d8OS5eCxBwl2ymXZsfkbt
NK/zWgWsqHO+F7SRNY58k52YDYKaWP9s+CboJck7VMRN71lzxupqBO0ST1YcFrGJ
YFRJ3wYFVaWt3XCZeXIpkDT2HbLHvugEy3daqHqINif/0GCu7+DB17XLvAX2EQNQ
oK0Qnn7h7H+JaCzcN6fHrgkHMNHRZC0kN7yolFmTN/IR3FHV2bMcLkvxPOxDjxwl
tg08lTNbNmU9Plr0Ns6zDtfjx93mz4h8n+d933amaRRbSu4BeOuG0QLPFxaDGglf
Dd+LAiDn7ALATjeDQOA5oeG5AVHl2gwNk+lQVHBir5JMYEU6u841JiHJS0c1dj6c
x5oxisSVYwUXbznZyBv/DR8LwGk1zLViuKTGZtpDt6CqZHhfLNdjT57mQ/LZPHkF
ATlA2jUXnJsfQQbbxOvIwkptFPzckuYf//I53j1JUSU9JBnza8aaV9MduK9fofOy
rT8eyV/u/uHSC+9RdWoJQRIah4fQyZ7aSHZbGCGR9y5DmShoaepW1jyiIrrZD82n
oKmlkE05Zg1nyD8Dd4oPrePRYIxLWs6H8jInCRh0/rGJJ+ygpO7ygrdNP/rECR4+
tBgkLd+xAhlAqC1ytHz68kAnDKxclxqZUO/snA8YnK9pCnlq9RwyH1/yjS+WNYe8
7FPVuzDx+lgodSDTM1q8jdiO1pyPqjCQ49dsre8T4/3I45V7wRYvc8Qw+zor/Hnq
swCTbF06QB3avgNz2bELBDzTD/2Zww8AuhFoSIlOrXOVGukGT/nbvhCQRL94Dv8w
+jES5n2aZJmLBwfHCnJ18TWdEJK1ZPwnhO1DL9LLC9ozfExNMkSnH6WFk6XFKdSL
ug4pkv55nKRMmsaoh4cfFxbvy5Ha7RSocNSVLRvMHgxJdQRPTEXYDKnjWtlDbv+R
VvQ8YLJUPS+GHo92k0qWPT5nRoUu8s4TG93fN2BDQGN6ncv9BxGFkSmonvDazaj6
aji1tNDI9J3fUBtlGYk12lvoaqcvxVhOcF27BGuAdcdDqoFSVva1D7W9a7spAyQe
oCenATWixu/pRVyAi3iqfcI7d9gM5t3Fh1JCveKDDdgzQcDB7HguX5FtRXUqBVYl
A5swkG3ROzZ49NARyGpLMvtoPpI8+E04AUXacLI5IOh2q2JYU1wMlaBdV5yMbr2g
k/auP0J8kF61/UM1ePe6HmP6gLEYmWKChvZbJd7p6SQkzOmLNDqPWl7+OZmbNCSM
9ZwdKRtVT5BCJDqowG+Xl1g3HIrvXy+4AzwbXJBG5tH+fJht4+4WXk/gUNGjVcm5
Kl3/bkoucfWxsmEsCfgWYf2RCYPAda+WoggHIAMsjJeOLK8dhXyHXbyAQ1Aqp6qc
eo2YTQpAWDZ6D+7hOs0jalwvRD+ghkuTSq2dtDjMNu/9bGbwU16b1zBUq7y14VHh
NBt1zcYz0TzcRVt8q0S0KPupNX3444VLIPdofR+eWcDMph3sc/stVEVjPYqKd1Ud
uYv4OenOZfeE9uMqlg5I1bwWK+/PTvfhI6rGi0opGu9/ds22NznuD4hwgd4JPltG
yFFA8QHIh93OqtIP3o7VoTXEavQNcBP0LFLE+n8WIg8lTdEiIvtsaVvDNrAbboME
kCU9AOljDXLXO85JFWpdpzCf1PgFAfLsG6/dsmMc+tR1ANzRvLsbNshyCovQhMcO
BtCzzfEn6k90wVjIMAIAOJ1JlixCTvdc36Dexo+zngJHUyIwDJkXn0WFBDIjfDwv
njwEycIEsuBBGnVHtEzNaaHFQS18dF5L/PPv3Qc9rKRmyQfSlb88l/P6BFu7xhUA
GsfruwCRpV42XyU0GYCq4bGwGA0zZfdjZEwxpL0CcOLQEAr+MhdZcPXlDl6XYZXd
3yeTIpaAHDftpDTwvElTQG8iPnA/7OatUHXE8OOQy8WtK0ywsXo7B//4SfQxLRk9
kToSkCcYLB0a5zG214hrES3slqU5PFjrZilzGf63IS6F8tzyzso+zKkELeORFt2T
cnC+5rW0HQcn6onx3vQaWsyk5Fs6Qfa6GpW5hnfiQZiGBIf1zR8zv6X+ycdVcrva
53Lta7LcatElNd1tyNhFLpndeH6dwFZSO1EX594gJhUetPqoaHmNT43C2RqUfBVj
5VxNll3RqKrosa8Y5cesX5pZmBkvtJmRZb0AOpme/soEOtaUjV5ZsPD+iH0UWBKe
4IlbqoggaPZHpgh6TlKTxAYfuRkUkDwpQ7NM10Bg+ESvFW1CAU2DJR5hyPTDgkg6
Z4bEIoM/1aQ/4260L+6WkOX6pE7SzaEudUHKDpSQ0MKj2bGiWWhDFcLBvEhGmaeN
sll1RjXsaPCzOBsCsdI42XEis4dez0ptNm88PdLLoex1+9WhrE9a5kt380k9psHN
rTMxTGGgQkzL5a8BA2puEt/+o+KWjON9dPzhrZjYLRa89tVohbfeglMFWH97byKW
lUddscqk6SsV2BwBGmYpa1blLSxqrn+3vI2FGnFN8O41Zc/YvvH+4F6umyIDg66x
UTe/nsFs1OwzI/1rXDAyvaipLm2ANlw9Mwl5iZXqlFLyp4UgcUy/EqKdkKVdBZ5y
1stiFK/cEZNfafofA7PPwgyHbngkXxkDan/HrhkJxB44aBGWHwy4o8mwLb86mqYJ
+iGkepw3egtYFhg3YoBiTX3LxwoL84JCwoyEGLqzIN+zuS5YWB17zKSWOoDuEH/O
4Ml/FPnUigDhRKqLR6tGc1YwcDoYa56tttftV5y52T/QcodA5KgXQ/zhULpxQroB
huUgHCau0ksbqLqhhbj5yd1wb7D11nFxGaXJRQPK2hFUNvdP1XC3wbPILYeYwMvs
7CV2ell97qQcI+bN9VRvpBObjsTz9aFFA59mJRsgxn0fUuJMFzaLW/mwv+6YpM6l
MnnFyOBkwTBrp5BGV/2aV4+Rlg80PYpVH31xUBa77/JjIFiSOnTmONO0f9Dg9wpa
WzM7CU2VpyktZivbismu7B039IwuHQIkgtOL0VJYXCoHHKR+dBEyfaoecPDh60oz
6W0+wPfCWdYqSrl6ErsgjTuUD3RJsHZLq8ZTwmh1dPuPpcNeY4QqU7e1Kl+HmvLu
CXX9H0kS6+YKu2Y1qk3yGCWqGrdna9U9AYCGj4blSD8VrBYej2XeUBnmVXliEqW4
1e/xaNQm9PAnvlEwmPyipA/kVSBJ98ovxpprieskR4Oz/H5QfJw5uy5OykSS4xhI
pG216CD1DXLSY9gWpkWe2Zg60L+1C+Bgry5pqyjqegn7QEomXdmoZpl4wM+5MLb/
yuut05JIbc5Lt2bEO9B6ok7Oh20wJpnI2OdAJOkKZzxHX/fe6Uy5t1NXA9KWLWfe
tmlOQgHEQO7JfsyONVmZMRH/yBO7aSFndo6ZTDeIwIx6N/GB/Uu1RHHbigN4wN+S
nz027IfugRDURhQiZPSOSBIJ97ByGOW8cs4Fhv9JLXriekB8ip42a68v/8Hz26t1
4tESZk/bTNA1v94R/RFNupByA0lIkvJX8sTQYfU+DMHtEFB3bZQSea66p8FWRFnU
dGpVD1HpfeTKidMABd4dd9iQXEMrXWQN3X3TWtcrZ5dcY/KeZo8eE7sWqbGWQCbq
tx4oPmYEf3ShgpiePUKfU3BpY98JsCNVwSZ0CUHkxYBI4icGlVEOdvUvoGPyG8XL
ukDhxJCgVdfKMna7vyEuls6pZReohig+BqqaT2w4r8afCcDMkxO6ZrQV5bo02t1G
cAGq9UY5KWKneXSEjQqoT3gX5IaPCuuiXJAFZZtnwjqg+wE6nx3INMyzQaHQ3d3q
68sGpEwRizy3KBkldSJMtpaxM+xLQWQXsKdbkYztryBVoyygsyqPsAvDDCiakEbq
JNS52EL9bOzTDlQ9ODHEHEViaGKowuGD248QPskpvDJSXEcT4yPJtJgObJE5BgWm
qg+zWUDdlk59ETBlzFzX1BnTm8QyX+dKv2c+YndM4BwjjkvfvjA/Y4eK1hN2oiMU
IH7wnmWiYby2SuJAuppBqSSkjiqWBtHWgdo6P9vTlObsenY4XZ9pNIp8Ax4I/1cs
JjYVVTavQbVGIZ2yDrYN8FxEWxlQs2qYOgbn1ryr+v/Ujppzck8bZqqBL4qlVdRL
cDBPUz5HH0Hk8zmuk5gepjur2KKuNTn6O2X8kQOpBZL0XrQfsrzqBGssmcU79Uzs
Me396IUGmy48aKOoClNUYiQGg32pF4Kxq5EEEW/v4W0vXXLxW+d7e3jKhPlQ+3tu
TMExEt0Othj5ExCIs1ehIxOEW0hVNJD4iIHurvUVH4Es12Sja+m+BjFN35pVTSJq
bbWgNlorMJ5nighpmb5lPRs3NCJRsRpG1tk5P4r08OKCsCQKOYiGrtcwrfoYqh8E
3W5BCjo0IHeTh+PIkCL9YvwFRjs4nXWf9rtbpU/AIuDJJHs9GcR7z7lBDTLX0cNt
dyjY6HWnv/VTGBSBPUd4tGPLV+yd34V6Lt1GF0AkQ0f1iyccLjWcSBw0HRJMQD22
Qw1Opjdz1aZLJ+YMXgF902IlEKnAN+MsgKBfq6gdQZxO7ZlO9+jHxPgEGRj/QLpf
Bd8H6S3pk0ye6v+Wa9MC7QMly0T3x3Cca2kPmosLvHySFpuk9SXohTNWlsGcZKl7
aGXmnk9/qWqo98KrQAn/c7HeWEYwRIWGoIt0B5wV8jHNsouDxa2p1brzBNGV9CpQ
Pkeu4xYSQSDiBcv+AuwhT/YrPuD8f7/Xe1TihL3kPd1uEgvyMCn+kITxvbz3Jlmy
4Q6xVJp57fnkQdaqpadooV+AhySgcJXlksFV/E23Wu3pjBxwqqYLD4QH/j7pvLuk
moeTNhIwYAswwzX7eX4nO5gaa4mF0AoFifiq9vFmPDKwKIvVFvSYzn0nnNstEhmY
fwoSmYOSSZ6v+T13+gbCOpJB/5SxKMPAQLO664wfWgD94FKl/po3T7bwYVeg9GOO
BgQJIOs7wgeZQOM8Fh1CiiKCovJtRmFWxKPX9ns9KdQBP5EpmnEd5iozCfTbtkCD
LPntkLvpb5VULlkzDUMVpoV22RHF2y39ZXjlQvHdOZxhLHCPIHwdveANR76bHzLI
ojuy87xpGP99go5StGAPlm9NxYTR4YzGOs3qlGXRwyC7N+PhX5guYS6IN7EMo0f9
jPKi0kaVff//hXL+lP1hiA/KdLEpOiIg1M/Wrro1Vuzwvu63fuk1O/gG5QJr48FU
KNyf0GwyFMK35z/t1onandr8EFCh7EEN9a8nC5lLv7i1bfV0Q3UTY+zdtpVtd2mt
oiBK5WAbvVtkTawBHk3hg0AIh1/L4s9R6gJs1Po83MiHHr7/GYog2NVmgbZ4OrG8
RjW/FOSsqErn1MziRWeSwKMHV0AX7a5QViFKTx9jms0SP7C/KP+2W5m6KwqC7/R7
tBPiIL26tNb1tJmtBSKaU0k5QwRUabxupF4XsF+vW/TvtMEgDVD2d1NsoekgN1v7
6/gp4z+APO2DS4hHlk6zCK4xg655d3vs0mZH0LO5BJmbNZUPV7AcmxHCWWOCetGg
tMsn9uAx06eXj1ASuQQh6rJMxj5oDZN/C8EN+Kidmxo9b+yjANAJFoCNIBPO6Ed8
joVEODISXc0GrEfXtpid9JUIuZdRElW8/h0FBpmHJa3sInUYVEdF9kCG63k87CYL
H9R0IB1AYRK1LNymnkM4lDcj289X0+5DVJOz2tetYzEx7ZHEToi2rSoifXUNZu8K
o1hy8llauGWQY+qYwnvtXNgSC0Mh3GOJClQSAwLjZ+7z2RIcWlk47Ud5wmV9pkSr
UeS1vD8+ER/hPlDpY5m8ZW8Es9fow3XqJKQEU+G6FSog3ZoY+m1RdRYrgaN3Z/3Q
dbKoyxOehR1lERV9pRcure7TrnCybovO6bSz8ngk9G8EoDPJnLvQM70Fmsx1xnhb
GLuOK9yxhz5fIddMA1uGwOmqxQOEnpE3ydQF91zAz22+/Zwixq58JEG6UfkRU10k
S0dy9oDXfplOOqBBA1GAvho+Xo9rAENXD/MWnqTfHbu40sut4NCm3yfXuXbSLbAI
bpiexHDoXW9F5vn/IIT3Arf6Lp5w2XmlI6kEZBFTB0dMxEZDae1zECfr8W3kgDJO
+SxoYAi5/glsLnvfjbAI9A6POp/PUyYqvtKcYUT3O2V0dqkaKiVOtyqAfpNBDad2
CydtLelmoyl6mR6LFhhwWbCSPSUnb7ZT/HwW+0yMW673y5R8v8MywGp96gWulSgr
yujovtGCK3XpnOSZeJX8XZ4Ab/E364S/qCIuUM/5brcsNVGJ0w/pFvrVxIzuOR3w
78k5qWQjZ7CuJbBSFsrolHgfuAoEM0pXzYqDDMQ3uAOAgVmsJ2xfr+YSRgYcf234
u7ihJLrf0mGLn3vv5yuLBOEjpGGCwMQM5BjALMkkJxMUxhCq+oOVl+rfFoO7p786
BoLMK82HnH8W+mpXTYw1+JtcsmYokDngtpszyLRbvd0ANBjPB5TirblBsh3JoVaY
Jcc2p0Z0kjVUxfya6Wifu6Fjtpa49OsMwKB9Ja+rCfr3dnEjA68n8x31Il6cjgxM
wyXdA6mHeOAS1zrJ6EWbv3h4Z7FPUZQzU2d92vZHIyWYljPpr0v9Vz7WYWon4QIL
Bhm8qm/qViSFw/9fcQMY6tz7ccZSU3D04JpTOAy3GwM+kaOFyKRcGM5+/wqwev2E
7bLxVROhxaFcm3oZNAcOCrulSybI6UXZ8DlF67MMnMb9z9QMGSOaYoyt1ZRGkst5
g0RpSW43T5UzF9kY4WzQAlETFsOdoX8dDee/QEVVeMUf4w3m4d5SCFdbjFV14vEf
A3QyacaSrBqoCkMov+ef5J7gwjyqpLHO0dq5T0wx2z+s2jlOdD+1oKr5KaBZfw2f
dyo/BA272OEra0VcEoh6lrxGm8ybMfDATXKG21XGqxR+nLtk22oPO6+5ZzRZyJL/
neE1+LGSBzrNvKMJ98EfTI6O78X/A/kRZHtLDV09NtwRF1FmrjT8kD44I98mnT3P
AeJ/KNHRSjosyqqEgwiSHPiKVLxdBMagvhI3zzKO/Adjwa1boXu20ZIEF3PP4jHH
JYEL+xzhN3SshY6lz7aWm/MBkd0riASuGfqPRuw/TP5/57TOcariZgjCD+SllOVv
pIl4jUElAEDrhqqJWdnYV0FACjme+MioWKKwEhgnSFPPOKGBVdBkGG+qnGtO2FyH
iC7B4FiHBQWs0fUJ0vYSUSrpBIXFboD29q6OxRMTaGAq/2D1xvgIJPBBzaOIf0vE
EjoPnL5oNIpSH8TOPEUEdgL+PNbUnrpGnfFChXyN9o2Ux+u0kVPugR5lOWAmQf/G
vhpsnih8PvaRhvmc+SbZQIO+HuU37Ag4PQG0Fi42TpbnypEtiIff7LfojbX9Dy3t
RoqJuLfthsmBRmfiOfP2pLIwzsrFT7PhnpS4h2biU53kTzL1sAUER1mJJEzjPg5U
NwncZpbCEw3BPWC7+mjZKA5dHWR5kryPjEYU3Tl4KgfZFY8z9btVUidSs7cBJN8n
5gQ2I3fVYGEnfOi00XT/Nd0CAqc50DfJuHuKJmC76smRoa9w9em87Bj8Y6L6GfJK
41Z9s6kzJqBEN3lIpI+ff6S+f9MiFTujMhyKmqixMqD+YspG5/ei6gJ55QFbssmS
+VdbTV3lD/r01e9tE96qWlRcKzG8Z8eYmlXcBXxWXHbti7An3UJikF4sXnzg36Fa
mu0KFX0TMP4M0I1pE/5bGw43JK+B7rz+NbkgeOIZix/85QSO8h+XPbHvgr5UW6bT
nzeCLTmPrPLLFuklmnV3A+GFCBCSz/EOWJ/SL68ybYPT7/qt4esh38yyYRLTrep1
flAN77mHIQ+5G6j0nnE17g3B83KNKASELh7zKslEsPNBvgTIYa5HsmXObdP23ltI
qo594biMFIPucvRBRGwEmCMcPrafcc6OuWDxf/YFmX1Wm+uf7gp5iXArjtNhPkii
kxkqiHslL09acbpwmEDdF1+LVpl01dTFBES1ewrkI/zgKVXp+wMVclAelwLZDfKk
3VQFT28FHZsENlh9W3Y/rsJtMFoIF2WVUvNxbGJr3sXPKu2B0/W2vnzeacqq7I2f
ALdgyzdbUpTueSCsGnKvC4ihsXPwC3/lQZmwJ45/r3BsO6hxuZHuyWLgSDd/OVHv
7vIrxrqfo//YBGnZy0Br0UBsvKN6AXC8wOeymakm4zhWplkMCxLG7qyaTS9svRpg
4wbBLxd4lEnT1njEOKJ32s3r7fXlRj3kU9lQD7Bq9fDl5QYrGEmUa1yXSuIlEYTc
uxxrDiIXsbub3AvBDA5AWPzQkvCL0ZRGbDnYqAy/Alb2hKvz4ovIrxNaupupDdRP
uECRZn0XXwzTp/VapjYuq1iQZiysgutHw2ao8N0Iqx2YnAnI00Ane6l9C3k0YEp6
5CtqaZiRAp6vLkt1v7jfRK5cOdRUbtNMYgk4xXIG1PxpuQgwAVeJZok8LqMYOZot
GnYBXmmN2RVi5JYzpvw2/BU99Uj97YQa6bbXdwF3tYkvVfEg5btsForp2MWpSQ1t
Aj822DsneSjBcRSclTNcSxUl1wD3pVSnjbYDpd0oQqa7G20vuOhIPsXLbooTZ1/E
4Ze4IUhQ3GEloOataLR+q9S5mqPwXrF2v70YAcBesgtja2nOnnbTU+axIKZYPVvx
cJlpsXgI6EWcN9TEkKr0t3v78/PEO+DMLi9o15HwOD8qxORhySFCpUeUMBURnRKr
VEnCgz3IUNZu7Y3ezHDfw48cjTN7MZEMT1u91S2jDvfv7OaD0eZzOceDAEEUC22z
HmmU22ts01e6zaLt7XJmRnSUTqIphl5e2s2bVH95tHZ6++adDPEL2n0y8zr0Nqt2
JqwkDkGlgqb8QKB1M1+RnlYNqxlh1uGap1yq5pAiWvFVPuNq87dKLLCG1mRXdYSx
flGv0rbnG6R7I+Ea7ir4TZwGIlBPHXob8eM+sE53HF8W0NysO3iF2fe9qm3mUIts
dUeX5XK6CpZY/aMVkZzyebHbk3KVlWar05dn3uQH07ZP7lW7dcnds4/+FMZpG1Qy
p3TPgJzwCFmgalvAo6NEOZrMm7wblVkVoMwj2772ok3jp4N9h2aulvLhn/mrU6Us
B/f7LnWZEXwtFV3IA1UjUFZfkPplyQ7n+Py82qEMK2a5U1mEBroaRwMmJbSrgQGA
4OMIh3BSqsIKGSMouaoVgY8xR4vgsIdGlDhe9U8s29nwE+xsx9sEYqxX5Cr1nlGj
vQpUub2iwOGMgQES57IEhh6KSZD8QJuCT0ijfgtJ9Gu4L37dAHOT9pf9YlUWypkQ
2gzHe3vEW+7/dBJIr+IsHIOzlPyFp+vxUAjAwmN3LqqYbgX6b+vqqJve6Sd5Cu1v
qybxUapLOyJZLJ32KLQ0ZUlXZ3kW7ej0UVyfvbo+UobeJAcV36RJTlvCY6Ykj3cI
3eo4IpfpHOGo9F1LznBA/RFfwQl0J2EoHoA3SR+BrgKcu25Uj79uKg17j4boDzxf
2GKRiVexeH3vbiSIn7oNV0JGn98/tFDINL/rUg5xrP2xG77JzCte648d/5nxLLTf
SG4dI+13mmvF2/BTV440+NITMn+bP0xVT0WS9+yadfDfDHF3EWJzJAVRDgBAu6O/
Dm0xq46kJ/jfNbh4ldwDbErFFFc+RtSF8/H5jNHtbLmnVWSxBdJA96VOAz5nD2Bv
xqrvGoD/IRDNbHlGH2fyaF5ZAbSLBXPBShkkG9T2b3wICXlHKNAw3LtGc1CS8+/M
zI+w0JNYmWFpFA0vBxnJfG+fU+HK17V8mbdWal5Y30axQKqivlMS7mJo4R8xwCKz
eEbnrNPEnRvl72fwYtGsBpy//Dajy/vAOd2JeXhFkjKQw542yXdTdifG6/iCV7wQ
Wby1yUWfwpmACPWq+HBoIvSxXtdNXLqaJen7EF99M1ZzVNiu5wwJtEYQVOiUHJif
o6IRhQL4uc0eHTgvjBp1vE1TdW2Dya+we+BzXp7SPujre5Q6jBJW6wXYk9fNLLpc
yipF/wZ5YK+uqib2iTIgfaumgShAnebcyjBTO5LeQbYSyay6ZqUcNiqsTp9WtDP5
sa7XcyJNJQr0rsNq+QUZD1nHWbKGgFS79MByWbExkZT3IXn5Y7CaDJdr3uo2MJLI
8xzyb3Pw/wY51PowjWZX8CGdDCSlTcPefPo+PfegMNiJWf+FIS/ANZFl988b5hlr
/AIJxk7iasikzSBQxh13kPxHZiP3HkcbeI8X4RCiK3hUaLYYllZg6cfH+vV55qJ3
sfb7KHWOoa58jCroAHSVze+6yPFQb8199HqX3N7VM2nYwMzuZOsentEJcsY6pxTI
Zh1IRvmULj8Q7kcnsgUwmoK/EibbKnQ6FFcEGNijh94UjM/AF/Bk7v34mpwO1/g6
y3zwZAF8UKnBxICw7RTjJoDswrRtmkxMJmJon5+WqGLEkPo0ZhLrV0XETgpCe0h+
tICJVJsgEdeC0RpyJmQ6xwljUs+pgPloovOVrZ2POq1WX3nFFuR8ucHIdMtoeOKE
KTpfLwB3h2cCzSNYw688fIe7eDwOFbM1UnEqw1KF6yfkCKPQJkrE3AWgw+58ZDru
dBDf2ad2PCIQONgHZvjx92ApxMr/4DL/LV6SifmZUpwhwm3a6AJQ6DzoH/UIJmOm
RogipnUvzQCfoXSrISMs+FJmnMKBx63ha0Q25Sfi5Kt78YiRA2xtyigLO6j8zYVQ
m3EOq3QffZmgdlEjxnGfm37MXSLZSWMuYkeEHYW9gs2nVha9k4pjFJV/otI1LIbx
Gd9tFMdUAzcZX/MLwGsTpAp8Ps8X5mF72Th4wya6bDO7DRB2hUHwZlkc48TsQXoj
IAo4uIIJAA86BXpkDG3f+YynaZXVxxfuUt1sOoPDPjLek9iEy8vCP7zZI8XpoklM
Jmx73Oko+afdb4SPqfEJ7E65v1r6sLR5jTfmx8lll+3dLjK+XZWlyjI3oJmhbQMi
WNQ39VicFQKH9nQ7D+QYopEmQB1iWzR8ChovvEXKNCBibuStTWVTkxhvxF6iyKhw
PRm7dfuIXliVAM/Vo5qH7TwspnzhH4VjHDL8FvLM2gcu2kwfi7lGY1FIrv9acJgJ
xQSREtVvsub+n+Kxu97BzBA+I3xG/W+EYgllkslghSsFyIycyIItxCTD4XjK1FDE
VeOBunubj8d/lRM8lVrpASISTN70L0B4kCb9bhTh1yazLUb1XkY+XZZuAreosXPW
NbE1QttmUIMRO2GJsTIacPegwbYY9dXJSdAEALwb6pyOC6NZ/hSJC+JDgfUv0XF4
nKLnmhNQtc6j2s4tFs307wd3aKSu8DkBPL0UroauUG8x37hS4hm+GI/mfTQ0hU8K
y+zWrf+cyc768aV89sT2Wpi1fX6hFTVPbuhdsdfkKTbmhw4pdD+LQGUjuufQ2iXy
gLRIYd3y6w9QyWbahVWjzBdUYUsnj+NPRuGnoN2P77fwYCeboJukoh2mv3y1gEmP
NSpTBC9Zv90Otl/DF4582cYvkQqRYhaOYcVqlTk26ZpPTIgA21jCs4G1h8vuRQ5v
ZeSPOeS60jp/Ly5Ubl3vM1vuJJ+wqbdiq5APfqrtu0q6fZSPCLxrZe/tSyoUk3b5
Sd2gDQrouIMzcITa+evD50/i3B2mp0BJ/GNfIuDXPYxQnAX7w2VnID/FGJC/GceF
aR+tgcp2vlmSotVMgmdIpDRwW9K5QWWYOzlTzoTT7pD1AIE2rcfuAaW9gmMkei2w
6yRRzrtIsSNk6ecpIQ+w4mzd7GSs5OQS8ORKDexchpb7A/VumU3eF60tWrNztN96
+Y7dsb7LrYTtVBkJRndA50V4SQTNRNhJTcDv8WAGr5RhfpHgQ4G5/b0Nwah2cQfP
zKMh937uzwHMeIqs9GdAW59Q2+0kdBxs2cuUwj9nPEfwq6hn+z1xt0KMopWJ/ldu
h1yaDdLZ5fY6fWpb5ZANKoSRFLobiDC6jZJw/UPnyMBu0wGYglYS3IHtrg2Q5hnq
KibrOvc28JyC9Gvszjk5CjL341JdCfvxbyF47BH8ovnlGvJETOV5MBwFmsi0SRNp
dE/ASxSU0ICvO1dT/c1/Z/+r3qCCadStJ0mP3OVKHNCq7hlRDydSuIJ3H16xLzni
4du8XNZjq3/hmlOUK7dwYpVacFRsu3zBkTJkyQfQh2zSHgVBbtmzY0xvKYq7F+iM
J26mbk4qtXq+SotXOqvKwE8Ds0P7mMqaevo82owLnRrX6WWbuu5nQBfBwm6N+tLB
CIhLOVRZ2KpP4p8gWQ9N+pculJqR3Nx2Gug1aGt7nFtonDT3mf6YeOOXabD4Qly/
vFl+EF2HDh2QdOPVpgofFDpGaegadx41QWvFw/o6MHd6YtbspYBHujgYUzAjRBuR
YOqhqW7WAqcBZQNDgskkw/URO0xhU1zYC5nlnTdmwo4SKNYKGawbfwLw0oHldLmX
rSBnD+BTe/v1t/JFiMBNKnAUhbiJDEfA2zu/Q4Jh+7mEjkB+3iQsd6KY0k5Uql7B
nxHgcf6UkZZNYodsWA6Dlo1WMtJBq3B63eWGV5kFvyvB5Ut3jWKveAOk18F/B5LV
il33gVXLCghEFG2sux05MdThoZAXv096ziQfD1+rgOIM9U/J+3FooYqqmGpCgUVC
Cot4MYXIyH5/wIxUnCwmDsyQNcmuc5l2j7ly13xsFZLp0/pcO84lmvVlCUBOTnej
PekFisoNytnTwVIdfBf5Sq0gT6pUnX07GTzfndE+8jGHpTCLq8//GI7WOo2Tzsvj
TKNiybnzsjGcTD5F/fysWN0FccFz1DnYpDuGPaTRYyUcjfRSlEofgZhiMKOEAKfF
yG1XvfgHVUOw8sIMSnTbMA1cvAAexeB97gG8//YuldbcNqmNO1uh34s1jsEknk3q
4bi70673RwsMceaHbai/azXLxhHf58cmAHLejv4jOSfatdUUjhsMjMY2JDcjZ/l+
jUhSZCPvMGnupgaoF0oXOrvV3AMetIbkHar78ZUdaIq6Nnsp/i1YL+ocI7awSVqj
eIdtOMVEnsRmOL//dYn9OVPRZkJH2yuSY5Cjw/xnViWrjTsmlvfa1TouAzGP9kZj
MdT288bYgiI/MBhMg3gm9k1dKUGRvNiVHBcCQVaNkB9KEN9/BpgEY9FsucClgDFA
7Eq5CvE3DncHIr1/QgQ3uCmuMjmji85nZ0AvImSdssVGKlRnlns5YqhyK9f7lyqc
X8JY6r4GaUWshQbap7azIxuMHD4wstrJ9NofhGVZ8sPFfTxw7RMzPkDVgpLCfrMz
fMTBwnQiJ4CtTZlUised+ugtKGSwN+o4fMZHurF5PTJb7N6XkNUZVz1GXXHs4/Rp
9Y2f4L+dlE8+spEuIOL5/HhdI956+vnV/EZnikcHnk6Hx/1XCke/9sxe+C2PtOkh
QLP/6u8eBYk+CV44zy7NU7xiz0s6We4ct0t5CB0Rt7a8jsjBtfK1F8EO7yTbzqc2
bHzq8i72kfOZPOVjK/tt/i3Gsikoq7Ezr+MUTp5sfb9sV0LQ71C8bVlBBIjMMTvP
9sEBSkcJeLgW5X9CiYCWNKeeNVjoNIcHfuQwY5vuFPiZs0X1ArluixxXVpH1Awc/
AEiUegSJtI4AtktIlt/7lts6E3pvbCQ64sYU5j080ouciKqL8khzCFRYjX7ayMVI
3n3dIytfuQtSUoe6xw9YT7U+svjg1gmQvnjO+jEbiHucY3Lj8pfjdctRPUUdlhVi
mPT8/tIGaloJQu2hEoIOS0NCoLprlhxawMNQIIwzR19KgOfwSSlyEyqo7NNca6C0
yBdwT/8Am+8GWdkNpCjN8UQCy+lvSGeHJUgXXhgy554uclu5bSPht/Zip/ndbmqz
67J7o1nUOFXnGUzIuZtVR/lqLLkV/04Ghr4lUnERxr4x0TTv/RR/zLpwYy8dPoUr
yTu2w9WeUN+KThW9JjzEo7KlL3RU2OQOwcthAc8pv4maF9yvat/ZuWYyjYJ2XlSg
LirJeWkoisKWjgcWoBGxJcNy5h42qWZ4XUDjToTsChWqxHoWAbVaCQFgMsjxzfP7
p+oQGe8sFMILX8P7Vde4gXTEKOCeYSUa53g3pJAaDGPviCqgzgscGmvcMh4oCUfX
ZdfTJcetz9mKbuJpWZJZCpgppy/8CokRBSoldar9/D4CR3lloZvHMPoHxdFe/hrC
hy1af3K8cNPHV8CCWB7iP4plhJ4IQgxQVbOOBB3hu8Zy/JxJlR8M8SFF1cyFFJ8O
mkdznBpro5Qc90qTdHs4/R9QPdK9Ah3ckELxLjV4NRcAgVe8rwY7peVhz+6ZRS7v
aOIo00hPsZq0Ie4GOACcXENuFxdeLZ2C8lITG/1kFrpy079ka9262qxpD8nJCM+E
giLjMupDX6huOzQzsFoadG2V0w/Bm/S+uoHRa5CxjR4PbjJkJcrpciNHrpv+QQC4
U8YmkEP/rXpGl9XNuSnrXEo9lIh508oYsF416y0klxahwwKwNhQUnzpqSP0oSvgK
G/htmWSuAMMi3zuXWuPRuiPhC+uU+9RvW+84ojinsUk8NAFTjHwwc+lRBISkJyUv
kcqjmtTfF0GGYxbglm9lW0KlCxRcG5m5eyVTR6YNp/bRsr9iJrHDII2UN7UwN3kz
NuB4b1tyzDBVV9+N7dYCZBQo722jEuNsNV83LCL8pEyzwSKkxyTf8g6L4jPoZLaB
BBQ35ssv3VpS2KG7wsqH4RXIvuzJdctjj4Vya/PYtf4vjT3Q/xhN9TYO1kyaPWM2
8qZKkMVE4TEy54lkDuls0157echeXMRF+naAxfmIOmu/Nr3hZunKUL6UfPbD8D1q
RbrjXj3AmgswpJ8liZ0s0toefQg3wNEynTSaIXvzSsMrnovYhb+0KztEGSCh4Nem
Ad9hxm/El3Qqlt6O/zXTEVdb4QmJim7a/aYwOEODyfhGmsgikQAdq+zahbeWnPnv
fJyy+lh71lWN2h3+udmZbBwtx7HivHKjZGG5jLXu6vQbI9ThR6c/hRPQjIpKWtoY
IXFKWocjhSrGk8lrn+aDDl1OBiE/lMiHGtvhVoL8XENEKx2INzHKUuX2JpcDwtzK
xXJiTCozgNRtl3/xTTFLVha+rK/zKP348pf5yy99MKF/jG1zOs+fw/bPwjJ92Ipe
cV3ZszlAtrmXhev36BdlV69aAvKb4xio9KBFWroYT9CslvnriYqLj5Q1YYKYL10Y
bm9/4rlRV8MluUhDfGrRUWCbStTYfk7M79zCO2tItNuvWUlDkdlzGbJMBfmblZ4z
648BIWTI/Ac+crN0VGk6fiwXk7841hFKkoj8qy/Des5qAYlnQ3A0u6M9UFWPMfbR
wAfjKSh147/c6TfkX3ydLvnfiMpCRNbTk+NsN8yl1Gj5IhAwR7Vhx5rvCE5LojNs
7VvQPLefpiPViUkZXIEvedaI4lqROfB8xB6SYo9EWsZBuABq6MwrU2xPA1Xr0MB6
3AOt18CwWh3l2we3tzqagVUGWfZ09enukUtBGjkM/Vsoc1oC6VpoEDlBIjfCqoDe
nrtfBgfbjRQjcF2IDfNPD4AmiqJ2q05vecUiBUFBRVbgl3OujP0n0jPzShZK+LEb
dLfidFkAw58VXFP2sf2KyBephhWfCfqNyaWMv6H4q5EsrbjP02GyG7keNiTDvYvW
OM60l49PoB03kyL7ueESHrHf0nDfpVgLRcoFI3bCSyFfWfV5K61J+extmKvjmRBE
hhGE/0s1IOaGrPYGCc0y1riEt5xY7/oqaFKono74xkzo3I1cdnl6aWB6uHnJz88T
+wCLTdI0AKzlKeglljr64F1imar63SLiHFfgGAurDIavZOiab2YcB/s/B/ZCe9gI
fxb8l/TsxviopYknGOmCoajf1PBFU3EP437bCX/xZtUlb4IwDgD8BafQxBYaRffW
aaCDI1bI6ltUNTIrIZPCmpQaYvLRjz1JTa8ufjs51Zgp5rG2YAPxDvz7UmXlytLQ
Vp5pXhPoSU58LEj85dsgpWHsVcUmw2gigdi+eOmv8YRR5gT7PL3FFsztPTlO1dUK
xs4gd0u2M6oVkTrwsOAaAQ8mmDuNbBtzxM/HjwhQsXQvJdwtn+WwL4ZkN/IOlwwY
E0RJN3PALU4agMA9rsZWHSbCyKRL+nPMju4awXwyEWqC7oGm1JZS7u0xRrcxITLr
ItJSWWt/1ZK8QqAP+v1iAMm06zdZHJd8ZMrTKrfjvGTbs2E1T9GuxP+mRffPHXJP
4+fjGGwJZNGMQofrl+wnZ1DH+EDyCcXGb4h8oMe/uJ7ZsbaTfkYCoGPSUVhWg+5K
IR41P/URJtaANDFb/GfuWGd5rxpgnjt5qgefedaCVBom2zkxXZPRqlzSGCwkWtBf
E2BNntAgzeQAL18VHzhIdBv9DMX/+sDhr6FTbehveHLPUwv/ZYcnSq8Dt0MhwhV2
I2RCa9rF6lz78V60eAE7VUEMVRJHOH8piUHqZgqMU+LrNUeJaIWunWfbNLkGXfFf
78rIA49t7W2u+QYMEHFn5ZQfbZNazZhGmcxiQmpt1rrKntGbaNoOT8tp9oT71auy
wt+2lyEyL3DUSTmIjpUAqXvWe9l4qAg7nKzOaUNlhKQ/9kvrt4Du3p41RwF2x6w/
ZJ37vN0ANkdWz6GwxqberjpOM82PXF7ZsVIgUkelxIAMN0sQ/5rYfsbR7Hwrb+QG
Y1ebQ6hEvco5u2I80VE+vBjRt/AuC10VnasZmJeo7NNYxSqtiD9/b+h5vOEsQH/o
TUCExy7VFLs+Vd3y+9cm9HmzhGS644pj7WnRcDk443oMqu4S4rm0hQmC5TwYPwQ2
KVQ8kDhjMq5TGTjeK17Gmo58ktkiF+rGlM99ul7RR3TwRBx5fnF9XUn+jaiHjH3f
/WQY2NFBb6rvaXkF2tJx1nhUnjAB0iQn4MPsCImI68PmyjS6pTp6s+WawGl7Llsy
SjQjFV/2TUYQWhW4wHA1bSUJ2EFj79YMH9LcBZR3/7CUt9IzT8S8I9OEsM1j955K
wOFGEz+AufkpBfTx/PAZ/saJ99ua9rFzdCSkqg4AtGX/xQgMQA85SKAc9K0MhIsX
HQMKwYYa2hyTQfg37T2DpfWZM805o11q7Q+y1Dpqh3e1PRtoJY7GqiLGGHFa8Xh+
Dlc1MnDpI1Epw8rJj0sAzrPyGU/E7c97gbChEkLHxeNSVtGM5VmVIUJCb+qd+Ky8
fxMVSZERS8WQmNpmiREZm20dmJt4SMi2fBnVzUS/poZA/uWj2ZZ330+qweBGFi/t
BjIAUwTVHwgJOT2HKrsI9XM/sdDSo5fbhyHAkpmLPZC8lS/qtC4Y1zYt5hDyAjsg
6YF+v+P/4tgRodKXCL6l/eJCPZY+EzSXuD3rh4RkjldF4ua3vM7YZWs1sxOKaGaU
BBwuKQWJ+2kPDBfeNunpqbA2NhU0MjSKthkmBMYfDKrw8Q/QdHjew+83ww/+hbYg
ZsSRiKciKemza1sICEJGimD59v3XiUX6qPnEnviL4oCMbrfu4EvlzGPmonBMmRBy
iPEm9Syq6LK8waD+GESAh2j98xKcAy2ul/nQuZoUL7iKy458o6Wrq97Ol6DEXLLj
Hp7V1svpRQcdqOSO948jTL74az13jeUPxh8AL+4EQYnB5qpzPmWENTBgF+ltl9ZR
hCwY0UAzE+nwur/OOTAhZYVmHGbKLZc2gqEMHFN62FAhLYIezatK0Jx+Lc1bVcN2
SJGB4XLfsZuCwQM7G2BeMFItbyWWmInGTUc2gjfbkIqwbX107MO6EZYgaX6kgBNi
vhmmtft0lDM9OGo777+coP/vFGwFwnDTeqp0Dg95yMEBoPSknUlXj/TjnXxD4ib8
06KhwrIyud3xTbcyf2kbnYs6GDhVjBaUydCxMHPNZjQtJsO7fZZ7Y31hFrvlzOdT
F306q9Cmpv5KLY4v8dZPnUNe4OHC9JqckX9tGXAuHz7/QglEitFSgS7kva8fdTRi
DDy2in+NLUtRVd8DBv5veQMD+JzEn56gPD7Y1jYo4OSNT0t7aicHplQUGths2SRv
AwoaX1qIBD66ntcziHj7/c/eDJYw8eILv0VepyKenEPOoTxzBFGNZ0+kgcZ7c/gQ
HUAvj1Fs+38R4VomglurSmyj1aqUej1LrMmxyO7c62Kzxb2XikDG+5NkgWzQv99Y
81wVw1dvLwKh9qbNyqas2WdmlGakra/rsTBFFdyCpFtSkqocyMO6qJEa1BVSTEws
Y4h65HNoOzQhuAumjkLIbPIeABf7NShpGkznh7mgdf0AZ+4HHRAEhnpytbU48zI9
pPyUrrus/tYocffWdus8+3m/ml0oi2XYF7tkyNVwRagfsVlw1KJtSRR/+4lBMfBx
06wAUiEpbhHzKHPk5+zYd/SLqY6gH94mtTJgb6VDmhzPvz2+v9Gfe+AytmOQ0BwR
fKaO4Z/BzSxQK7mx4NGf+XTgWl07/NzMo6L0Gq6bWlHKXeWPPgIycCPQgx05f0IQ
07tS70eTBQ/gmfeYZZuw/yJ54JEV+WahoKeIcy1/gfDwzK3fTgzYqNbPlg5Ql4+I
eWn7L/mi+wJ/y7SalRqFKGnugKxy7/8ZRab24vPvM6bUWgJc4Zc5j1EnVCAcldFr
r1HL4rrOgjIi3bvIhVOT6ObhY8EAT+xZ3utIfKQKyCdDCZG2Z8eX72Cq1FlREhBT
ySFFKdpK5zJAl5gTTrxu5r0H9lWagRPAHvJHQtlunZb1PdBKWMRoU8N54iPt89QO
ZKBpJckd9FGXP0SsD/XBbRenzv/fVd77UkG97hb/bOnvFXTxPeBX/U93mRfcX1Vr
aHwivTs3oOkY6VhmHQorVDhO1C+/Y58zqUphuM99B/ev/MRgI3E1bmLEPVBlHcet
bH8UKqskK2ap1gWRxwrUmRcsI9SVgE1y5tlFEJ1eSd0rZambLe265NlxRq0o4RON
41jp+6KbASypB76Jt3rd0vow63FWzwlfzxMZwBvVQXoKu1jv5dzGcbkv78LUiYN8
0KhBGBqVRgz0VBPx1Yf+U+TZGof9do5MZs4HbZg71/yDnhBh9YeYl+4/gllG3v5/
vkc8jfzaoewGOt136M6bOigYrUxCn+PCQhBU1GSXrINWkgmo8TELo+GvM0toaDu/
mWswbXpEe0guY6SVHw4gDZ6NQ/WvylnWf88u7Xum2yZ75XNOmMXTyykEWwQ2lJWT
gLJam6/TsZzVaor392gx3mBDU+9HfVDN/OqxHrV7CVDm6gTElYj5xUg/GCzwUFKZ
2fMMqfu2fIs5gC6jcOeYDMGYXOh6WidaNRWDwY6H/ftv1JzlZRApRRbaCp7cUjYv
G3w/PtNiMPFPMyzLYEBOWsmTYHvdbH7MglFLBA0GaahheB0F+R0LR8Pfh/c4ays9
3sOJxGIymdKZVWf1OD2EivJXadbbaoQYfHlA45qm3w9yGVXizEMBqrTbPi/w7knE
RURNh0ykYu2r7lgsgkq2PUbhaSCWJe2Jp5ev0/rMzLRuXibF1/LIU+B7zoxuHoLx
9MahVVhdoGVfJPZnd/ObVC9toQlhat8w4UPU1Gw2+lJ1g90MaMFgV6uSd+xFO7Ae
B9w8WC3SEvsi5AEilyi9A1VnflDI+k3GVWNYWQ4zrKZOXAISIZnC/ENL75+HZhnT
6c3aPvxGX8HSi/A0MjTxX5+qOLonO7W/Uc5MU5iXpM4pJ7kGkoRtZBrYqvYxat4e
omAjJFCvUVndAL/9d4uNt/g3aJFqBl4e1Zy9TVVtQw/KN+ABSUVAKAacRLdUu8nZ
ar/jbD5Gmv0lQuSKUS5o/BIlbeQsX11jmtFK1b2Hcjj+ki2nDYjIuK0iZLSomX3X
dZ1d8WEcqdeAg//nsEHFsvcTaH9HEBTYXXnl5wkFzwJCOYv06b0hVfNhGKccHPEU
ZV1yRS9+IDJ/pfxmZvx+NbVJaaTaNtdZvZQhPCLGrcYskpasnyF49f1r8j2O5f6j
smRwxUwHtRBHzhDlVekq1JgTdMe18kvlY8h0pmvb2e9PAol2h9i8ABsJZk4xWC4s
tt+FkQU1B1OPt9ldL0D7oFd3eu+9dLT10D8BgSdVN6GImGDkgSr+4cNs2cKuNh50
5XLaVHQvh2StXiTbTj+9dz1LQhish2rapmCJdCbZEr8bBXAl9YoqAyBT/q/MOMNh
7yXSYXAzrXEoTQOK4KcBRJ+462sEnxEHZM+e2wYzRDQJIuHxMzS3tA4lObCIfqhw
tWMs+/bMqVk090TNaqmZ9uEeTm2LCvTyN4cBnwbyH+oB4YztiesGCIABdRIQh4p0
DNv6SSMVreZJNmhBmqwgggJXyCsSXXMXIaACc66zuA/q1FQHfqvENY8T4kkjHHGD
7GL4QucHMTWVwf/URiip6Bc/9hgfxzwHxIzxhuFflna0OHVrwggeKtGN6G5Q2Wrm
I8kcZgp5VkW234+JQcRG3glC7eVOwHg1u7OShpYy+84sA+pXJOzZ5mTcIv0v1t+k
5jd3gK3NCyRSUlff9vNxP1QafRfANLvaD9U9B2rgU2wAi4mU35sVyNzLN3PEWt/7
oo8mksdaFsylC1ljgP9tY5e6JgIkEy5IBIQ7nfHL4kfcUcvIB/PkU8SBgIDvz9CQ
iZbz0Lp4S2toKXlY3hcvl1OqbIRnccWOPHBI/szOe3Y8hrdJB5oS6psKKZlMbqu/
/XBb0tS8fbj5XVWLNIleldULQsiK5mgsyHqhQYM4yyiEymM5Vi4vKpNL84erFDyH
gk9al3iQyV3ARiBzhS3771QYZ+CEJUC9aWY5yIDjF8Z9OEj8TtMnoCXJdXV90873
IZEB98PYFGDpa9b0+M/YChw1sVcXp5a9FMP5gSX6p5QrO4oKqRzdL1JdufJ0O3cH
DrqGU2LgGLycjSXANz1E4CEThc+3UWb5LpCPwIM6Dj/VWjDGoTAnTloR2pbOGmZV
qDYtTBmOftZaWtV7yRMmRxhzamp31ynxtSqr/perDYS1sG0/LHsWGBXBohzqTPJ6
8YfIh/KQNOoZ0tq3+92O7YG/4ThnTuyHIRBTVguoDU3NA/hbjqnCZShQmhdkXb0D
kAt2aanGKnbWY+H02cWNWBtfIaNakPiTjC7pSNu9rmWGWtBb1zNpt39xMXwI5V3H
brxLdDsmcXnCq/W8tDESYGqMK1WkFCHkM4M5ESupQj/j6/DwKjrYY4JDk9elxsz0
FjpI9NctZtuLexS2/4VNgBeo22zPI0OTsOd/d+C7OcvqhX0JKsoy/DF0lvOyN98e
+xXoxUQ35xh5FX5aEKMvPjBpKQwIMhnDBFah+RqC4YWWmtFvk8Bj/7LKVQ9Ob4e5
gX3zllMENE9ENqdjP1dN3Ne3jxSqt+pXa018qlqtPATEv1Y1SsE4xcn45IcX6qCU
LJ39dZm24v1CiO4TD577c/TbaCry1rWMOj2Ymu38GNAkdN3pzaJVETr/HH3mVPuD
1yVW/OGLjUk2MK3I7LsLQMrOOVo9V7id5dqjKAifVcQonLRNHH5MmNxDpfKYx9m4
miDIJcxQr1oGqvUi2N+fYk8+zu3fT25MOGIAGIYDoPiPnPv9Fnyx3mEuXVXRzJP4
viksPEvZRV9pphF7jZbFfiKcmqcmRB7MZQ9hcXYbBpRdYtZKY2ck83dtqvLZ0iNU
mKobUF7d0zl0JpmqN6O9tE7k1Kk2Pa9oHfvmiI5bl1bgjdtd/f/2RlcixLBnn/9p
spQnPdvBkZbreobUkY2E+4g94OcRyVejgffPkkTZc3gjOoeZplYJx5odrupRFab5
WdiPD093WOhGSS7h1HQj6lt6GY43MXWp96l4nlPg/T/S+tG0vYsg8VE/9UECgJfZ
fjriDPtVNaRSEOzegFaC42ROkBK+ZYJ20jZ5NtOuLkcWgIaHFsEEldGKN2Finy6+
qYN3UHA268I5PM5yedJYh1oP9CGYclFDu0twQJDivEZNXaRVzZdb1/ZGD13AqGeQ
cX1fgq55+D34vffMabF1vHqn//vof5o6AMDoKJFHUZ0bnImMJNcPu9iXmlVAcYs9
0hBCIIq/s7PbrW95KlgpX+Ljh0lGy/m+jW2J8M038V1z1p2xU84VeB0oysWEHRbo
pTH95lRx7tRKHM6PqjedM3LvJKO7p51duN7+31KSSH77rdq4Djb6nii5wk2Fa0k+
MHzEO7YnqDcY3djjuaIlkKFnv3ZCVI47dhPGECJygMeeRR+/IFEOSss2wUL0nFdf
zosrphSexL6sZsibwHydTJDiETsbRlOcXUpeW+l3rql5/ZgsYChELGdjdU4KVPX6
/E2Q0cXHRuY/yOrkoCrKFKOcGE/bA7DLMv4tdYKwyQmKAKTt4qDGjs/GpmKMeWf4
n//lX5GYCxP0bVjy3A7ArNtkFehmo+2v8B15tzcJrJAwW9hxiWRKDjKLM+qX9BaZ
XHAhPXtu5n+LWtcun6XPoU/vSv1GUOacIXGrGQJIRfaJDc49ySGnWddk5zKUH6po
BRMO+XXgOwtNkw7qy4coxxWB5rqoMRTHIuPFT6p/zrjRm6WFo6Wn8ZsjK7YCVLEY
/2heksCNBN9jFCyTgmIBJBjxaAC3FhoYjSFFDQ2rWPNZxJVyYOHlw0XvxFSo/2UJ
vBIh3YIoERVQbQG7zYqBoM6PxojsedAgkCf5n7CpDYBH5XegOl7HVBNZCXqiNI8t
8KiqW03Wl5UoATO9vxxZMiwXiE5eUhu/EhPkKuHRNC84ukjl5drVffc5kuFV6M0u
aoqxL/f7io2TPVuYQ3XLgxbFWkv+V7B8G1TqWC8DtJ0xGLixaWRFr7b1fSY2hu32
R/JRJlzT1U1jrmNQhSqPZSjxXq1q5nvHDAOLn0qtj5RJEnCwSfNa72e0ZhuDfD//
IzRE9W8luUcosAmHLIe+TM8qyn7l9IN4ZPuV/EQ2qUYDm9orK1w1x6ThvwQpgiXC
Vdf5B61iH2OXVwNrbTaVcNJAyyACOpBHR/OtPeqgVXxiubIegptLJ3RnB5ejXUbp
vhePvjiF+RH6JK3PmML+AUnJ8yvvAl37p6qjIells4IdRimwhujg7hz51qjNGT4Y
hGtWY/qTN9giAFumiDm5CR4nbTb4M4z3CZzR7pzh1w/c0zzYVLlmggKHFh5kgsFJ
s+uu5UUZ57ekCu60aRSyMSsSDuHsu9QJQsYPAk475y3wd3c+aedUMCDxhiBIfNO1
GjU4pe8soo4otWZSIZIxogZzDyiKWb+NQusjF4sUNnSbVjT5l8y0LQcoUyqWIn/V
RwKPdwukgHuXUdGW79/dbrReMKABxnChG8s7xrk96nULbFoDArGreIm7u7e+5zDW
ic0xZq2vhLlmaATb9Ync+Caj0orc5IAxMOeBlKzJA3WIRFY3zarFj//S0jds+H0c
9PeEu7gCNXmWpbctYkK01gZZvKrcIt/HtdV92Pofg0pQmfCOs9pb9y/BcCnrMs/R
5mZTzvDPqpqFDQLCsqVanwWUmXzg+k2DtqMoa7YpF0Hs4C9ocNx9xNYjdOSCRLga
kzppx3G9yH7W+77wfs5qv8Uh4c9DBhsV8iRI5/l/OkOFb/5xwYYH+6JEMLxf3YrK
e2og8XA4sbkIRCWpv1j08a+ilzYjyeZGX0vkXo9lYCfQHhOD5yw1IB/73QLzQ4Q3
UH1+qbCiPKOb+SH3GXcVxgol0h0/bKofNvLkpFay0ZyqVVs8sCy7YOT7k1cqEqO7
sKyFMrVUNDZKEC0JA7Xk5pKg4rGgF9EtDswD7ViRsDhR8T+ezuaiH83VPC76Ki9w
FrQ1drKcprtEKl5V3SdRcpSmwMSCZA5K2zEcgUA7leR0k2Ca+v2z6I8IBuE4uW2/
Zyb16/ffwUjZchlTi3mODZWhfjRA28R4e0JiMEw0C9EAOat0ikz8dg9Y1MyLjnKE
iTCJ0vu80vcbiyIHnU8L1HG/srCHsRZjg2FsQ5EStvwPdNfInP4m53WQIgwZb184
oWGRGX4CyLQRzLEy5ZWV63efL8wiuUxHgHrC38FqOJBslOxTct0fRe7shBmUwSAl
BWs9H/pJaJP8ToR6/YQhFfWfawd/eLNWICD9oUwahHMKr9Mg0nsJ7/OZ5sdBqbJx
NfEQlddDhOQIh6FygM7SFmOBuYlg2bG155gtqB763Sfyf146UefwnAp1q7KmodpB
dEVGrqYgecqv4yFqc3/T7Az2QR08Q/eimSfQio+wh5WT4Ix++R9HO15eDFidwPCx
Ssuitf5TPvDdu5W0asqeh7xQS/Z3fgj+zLT+jhKFn13g8XltD+M1Fu/UDgBCe/n1
qt9YSHGXRGTZXnHVdrB5+pQxIzZZ3xlG3Z/eX7nQEr/cmeB3thLQUz9Trif7QXLJ
NBgx+vaeMLZq7CQufxYoFM0ayYyLLHgRZCdtKyYDN3ZsB6Kxm+GG2TWPnasA7tDI
TBPgAWq9arYGJruyZYrqegR6X6Q/c3DD7ILpAVMhPZoJfogwHW8NeavVnfwFuOXx
d6OpQbJr5913qOBYSH/ffLqgOQLR5TIvZ/yTT5pqq7ETBANGkVkqwYDWsgaCvjUy
L7brVBC6s3VWxufGpLQ+K4a+JApFvaZohEcs6HgMHR/cnxKK5CN5LFMu+oftM754
EDf2s7ootaqHIvTeMnXte6xxrAiRdl9XVCb4X1lbjwkyItdVMyG7m7nFo2eHMSPx
axwjR2ZJFjy87tNMkiQnFxcYph4WnytqB1Gbq3QJr3ALaFqZzk3Q1C5PkTkwpnWf
4ZOl9nso5Wdd4B/OQSkW85MRhaTRncEyks46q1nwCp/rV+8i/AFraj9WHXP5qAc1
f5sEJssudwJzZnSnOs4lvm4vka/Ml6dwLemJcX5DLvdSjacjJtSZ6Di5EmcKqFX4
Q8eVWa3Ollf+icJGLrcrFZBEsSm1frh/AOIEted0qEuphlzpy5Bu6M0r2L+E639Q
7Rv9rUSKhmr1MEEnjY92gJ42VzsKerrco50pL9CpVk1UNkri6SOr0lL8D1ExShjx
EHnIsHG7lva8grnYkg1Ks32qB2RXZBczWIDasgJ2kXRhJ82yR4HKOPG3fj/sRukv
ZHwEVSJnECbwsHtkMI3eojnHggOS9XSmQtQP8aA0Jb/vZtVg60zH5DSQAn/3FPxa
K8F3eTpQpvvTQTpWp3thrfrywY1OW9SNOoUVJhaADi/hWoiaRu2EEIS96NQAS1rw
XRRFH2eoxEvNZ9ikfFrbPxm9O6BtCWHPQ8SJwJlb+IHfB3ahtSRYdK501ziKrubU
jyL5VKaT6fhX+nu4zNeC7Wbu2f1QK4UDXfM0xOa9sujzW3tADjJ1s9ilMpB1vFYx
oeEIECtwcJIDnpMTZgQProNplBrJkbyEj6jjGtR7kb0OmZYi6mndVAUEpzPeXChH
V9pAR8B+FRJizI8Siq2NN9jM/chbpw3aFDhv6EyCA3Sj4ijZNiSuFqjfO6UAoXBT
c9BRVQD2Vre74VPAIPhLtVEyZNBcvelMhPYGDpxRM+RNqMg83l083bHPctZYIGN2
aDNwLeIaxXhOkGXASwEk3WRyUcxbYCcvt5WM/dvGfsEntT2wdllm1SkKr6S6SYqK
EIrk/lqeCTy3sMH0uGaJbokAOunxYWB+LWO9UciaUfkuRkxP6v5r1asqG3hp4ozy
KqK2rbvy37h4rHuIXRlnndcbh5zWCEOKlaQO1phy2podLWIDU7VUkyIrU10Aqp68
J+SMr8AthiiXqFl6y7j5vSwfTcrTHIHGf6ZZQb1mALugXcbM0EK44Z2ANsVKtcqx
v8Q7klO2frs8Rlr3stdVAgHmcd4rO81G2nEdUNnIAG1ErCrrcba2yeIVVL7cFh52
YPJqGncejUjCD5D7pRVY+XNQG2AIwiCeweFYb6wfhCMAlHDWLfzYBG5a8jQ78neI
p1rJPpnW1U7hGI6oYCFEk5P2+1YhsJquhJ0LX0/OYeEHuOh42C+elGUu8XViXINi
d1cbBnm86KQJBRmPGA37i5F/WC0MVbLI1K5xKoXqtlCpSjkNQWSozBTO35lJ4RxP
1GiHbV/O02W1GU8atE5XzyFR5IVFbhI1hy3qM3M5gAc0gjaQpkZed3GwAoOR4Uv2
HatbDWs3KqDQ6YSJckl1vvc/n3VgKbofLqzjDCtegtFtouIcB0paZQdhfrsvm/Qr
eNZ3fTFjsJ1+5H1Pu/cvxwRiXJ5e31yyJscHwcYyCoJIy85zNSPiE0pOMFK1KER4
+ATFisG36KP116hmj2YSN4jTGOX+XkNsumm1J0Xd6O8A4S9fEaXxx8NWQzfHwIde
bF5ZaV5+etgbR0jG4Jw48F98GD1MzSwEjLTqS2RC2uQUJmhICjgjtPhjGY8fU28Z
92/RAweZ1BVcqDLknujBBt09vIezoyuq+V9yelT9GxGQASbR9gucTg6sMa+Gh4Xb
jkaQ3gbQNMJNFKpdbEJXv0u+Pi/lsvOqOEHmn0udZ9hU54KRk/suUiUQzO5xvpWL
wicReMF82HJhY1ON+/JzViwGYpyddVuZAeRWyfC3ui/z4ECoTbdxfSC8Cl3QBQMt
/VYU7SEGEUSb23XjcFlkQ94p3qzvZa4qLP2aqlw72ihTY67QeiEDLKCxR1RgLmHw
fSstuuiWvOraZJ3b93PzuxxtCX+qQ1YviGHTTYrl7XFyR5/LNW5YgeZFijKNPo9z
YAhNZtTsglihahn1iVInDYstPT07JG3xz18DzREzqBXFuKOhHgny4pi2LLq5NYB6
2z8RSASbehsGdSjF8/VR2PVq/csTK2aBOQwIi2nIJFB48xkKqfOlrwn/YobnbNxQ
l3PihYEXqcWnhtHStYuxlxqX8yBwOBYQ+95CbsxHcIav4fh42YITqynrLTAZJGLo
FvCw55tnCn0aCSLZFRVWBp5FkYD/o68kbHxcdCmzBIBbAyHsRrYjinJrP7PK0b9R
xLzRANInbDfkOQTSkv2MuP5ardQnL3BC9mLjs9LnbcOoWyJc1QkCtvmK5X35Vdrg
nlB4oYM8d2l2/xkxnagNfrIpn5EZJuIyPAuxknUlzJi5AxdKC1jReRW43oSOF9eS
38TNU6qNlj7MR2IOKL/xwCtJT5gfMq5bJ3Vu8kPWZ3T0RiuJKwTbZCKvQUnC52eM
YXDXXdBMIz8NTRrjvUZi13KslKmo49z6BM2eii8eN5SYXZMVj5uWTUqvVsonHN+G
/pBYr3QHpfTCovpQiMdRxCvz9L33E8rRDXaS9VoAPSUKU0q32rW+Eir+tzu0WiLD
8LUsYpJjv9FxZrsWkdOtNC5xyivlI641VTVf7clvNM2Smznb3s5UPdda2S4vRI0d
tWe2Sobv54cGLfJwYZs/dfj5+3w9CS++jcDc5i88MOqP/lxK20FFw2NSlZ7JNlp0
sdQAbf4g6s0LskzZb6SmjgU0MWrIOXThKifjbCUwgIlpPpRx/buEDPbVrM3AqBFU
ho9qzxV+gJgFO58/xxkj3nd4U/9ETKdNhAJ8HwnXXMKojpIFM5DrXqjXgLmd8AiQ
ha8Bq8F3UVRN+9ECfETFHD1wGFJe18/kgCFUYKbKDLC6yWDagwKOsGKXgMciQf1r
0BxxehAu951ZWlpFh12YE11jyxve4Kqxry8FNqDxhtkZ1CdwhVkB0H9ssgyxAuSV
5fekQjqBCkcFe+Ijzy9BHmjlftIVlAQxYqvBhxEX3F1WIew0FB/XMLdIIuErlgwQ
cU6v1oSkDv1CShI8nUEIC/SQRf0iXJ8oe1ECFQpARByeH6G/UvQRb5KilGRxKGTC
r+mVHHai1HAZePaegp8nHfMMxYY8R6lSbpMGqfhKcgZtjQY4i852B5UAlMx88pRh
scVcNaYsh2rutP0bkM1MKANeWVh2IkVRdFXx35/JoaYPjpkZXdv1xGDIeeD5OnVq
M6K3sWuUqyPR+0gBCTD1E/l/mOqAlqajO90wfr1hVcGkpJ4iCxTsD1QciFu49Rnp
4MF3ntO44dCmGZvszJMXhOklBfAYUU+EW3khmIPFeVRLwTAqHqp6/aapS+Hx2xIa
T88hC2VgIlGaYcMx0lPFQ8fa2vTgY1r5N7UvqgBe5XjyRdOTXmBjNG/a6rneBkkH
ovRJBpA5yOGLZ2kxS0yNkQTqex9Xz2PXs4dmqRgurrK4VPW+wY+/o2sToaDXf5IM
B9X1LCMHB4CPLG7vHFslmRchtrkeuxBM4oujabbK6vTtnClRpd+M069ozGJQf7ki
+yj/58rG+rgG1EU+YCYrlYYkA0j2Mqn3E1FzxgaGea+QQX5UOwxXYKeFToaEfv4o
k0J1O5gdIZwO9+UJaUNqOscsdUAMmsa+rm3WEepX8ICRgKFkBVklP7Lp5c77xeCz
6r7V5CyGP748cJPf3Ttl3QqxEPuZ2pGSEKV2sIhoY+jDrFsHqfc0dN3SxkKYKEem
yR5HsyAUjMFMtO9O9B8DERFb+FJ7bU7pgDT6m1sAD7nzNZJD7BNlSP795uxuziJ4
twMfFyD2Pl0rbUAOZ6SVjf/OVdpimRsltwR3BZGJFrLQjNe1NlgGZPnBJk0AuPTD
qDzIozpawp9Z28AL64bjq2P+AOdofkrUKu/yyeeGxC7K7C40QeWSZQkfPEiUxegY
q8OSyiXjwS3h9AS3pDnGBiuAgutOPTrCg2Yqf+XHFYOWTpmjmCpKKGzRJ7bCxqMD
Ej2UPZxTNzf7Pd+hrpfGK7XaSrKN5xigXduEgjq4vGzWAvDh89eWXcNgkeJ/2XD4
8xq1Yn6tOjjdfo5xDbodRAJlenD2ofTdAoOBvuWKlLg5MgeUWBKeWtGilf0Da/8v
/PiOMwj8JBXp/DQbSLnzvNbo7nEXIXTBCDTMGQkb+koHuMWtLyrr+6jnqv+bitDN
q4JNyDmHHL6McsGCa7RvfQ64kniM6dT9kVLmD2cbimVsS0PCE/kpZV8QQxRFUJN8
2DdcvtHboXXgaDfEBfbwvh7CadlviTBLtXWM/E+6zUS9fJapTOR0eh5imKUvzDGC
+iFz/xu+TZAQmEvr7Dn8xZQTwN1eIdo7bHYqaI31CPMYUq7I/obeIHzI9fTcBwNV
nkPr5m34SQVJQMEQucQKiCsK3LoisIqPmJrEqemFjFVb1Prv3xWdeVAB+TJMd5eR
5NUSvd+kE/EJSM1u0my7ZMKC8G5CvHP2xNyWstLVsujzKDvsZca4uZ8QGq2PsS5f
Cy5feKNz9zQhkMJYLrFpoHSDxRhpLuo53l+3Tipr54juJPygVquv4As9gANfzBg6
EPVGY6+9u9FzItYQkgL/hBvIKt1E3JrE828IvUltNWaBFjswGi8Ue0A0QHRILQLB
nv1sqLgsfDmyAqAZ0uGpRvtASXcVwRNfgMHcxhbmJtXjzonMfsrLvh/hHWGagzGe
oRboupQQp9QustDz18L1ibhkjNQpNbP4b6Vy/Sm3T9Juo1osik2zl+HJ8g3vFwGA
OxYv8yz5NXPhAZpRGD6KNCcRHrrN5kEJtdEVCBKfNADVOx0jKz2aBESe2j3/ilvH
2NNleawI2YKsXTLpEcGQmepuW+3uHwf88QLwDqoj9D0prIrNm5qrDAOHyvHhDtLH
GkkJ9Q2sAqbz3jpjHzwFsHZf9fqHo3y3jW5gXqnVeNJbDhYRH71lG7573QVu4vux
xCK34Cv0i6GQEs9xPUP6aZXOdH1I5zoAH9+6PGZhUuyDcFbLQ06ZLeZgBhFQEOfi
OEKFyK3J4HAvtx4hCfjiMGtiLkBplSYlwi1KJxX3xeuqnNVm+JDDQsxQoc6vbiIt
9ZXHsCWcJXMbV8FdatMWeKvanimdGL2ye1x1ghpzpz3EM07c346T9/mIhOGb6guN
uiMahZykIneCBPd/MejsmPc25uYLrWuPABt/ZSnGOqt9apUcGu9FCv496ALhvH67
9stB6/nFpD7fWoBIg/8PLm2oI9lqLPRflN3XBRq4jB30MuUCcIHcJKaaL0nq/XA8
DcJrw8HIDezgIYkExSIMH9hZpf6RYWk3zXQfIFrJsTffIGH46pHybv6iJM1eVdUw
+7cjHKg6tkICQnsDs5tPlExsQHrPFkNXtDIdrX2PGNqoBQD05x7KWD+zDNkvW53L
IAjBsrHLLVduDJIBdpGS2KX63b0NHTPqMCkBxGl7tBd4Z7KJ25ww/ABuskiklzeB
M8GCBnbQnERz9xs0283C1QWjXyn9QhzzYaQDinnjuuKFWocMJZMw+4Q2dRa+zGXL
WWjdcu5DTvaHaFHW6KH96wp0c8bc1DX7pTLUUDmVNxGCMMnymEo2D+FmBgBKrc3X
sJZShTLSwsLGPTnYcLEShiruCti7r53/IybWfhdzv8mJmJhxIOqygbchulRlFOcp
DzhqAh/EpuT72xPNHDo33yIGoNk+20HVlGYbZ3J4y0bdYjm5uA1wJ/F6yXvbPH9l
VK0TltpF8ApblVVKZ8UGUgWHYtnDBcKN/1s1gJHL/yZ3EPeTOTsQ6CJRyMemHQEF
wQZ3PeimVdkbRe1jASqt4WTN1wZp7isd0G04Dg0ugHAMVg4uat4cQaU3t1bmuv41
4fXB1aIsuluBfteGJB1tNnteld7KCg9mQWEvXvT6wPhojLckQ9cViQmwtrTjkHuk
U0Iw/Y0b0vxGDL4QI2X9zXtY3fOEZqc7K+OnessxZwub8PiT9ysYeYmh5xHWSRa2
nGfYbvkgEmO8pcVnokqvHGB/CEE+zjBQc1NHLh3JDaT9TNMoE/4wlzPlnw/bx65l
CBabDwpEgxceCDYBLELSdk7QcDHtwO/MYGtd3gQsh/+QZt/4YdRoSc2+7Om4/ddg
wbzzMB6OxtLJ+IG0TD3jte1pHnWiuxV5Q3Q+pI/SRtT1Yx5iAt2dMjNxhTa5N+rV
45v4jcEyLjtd81HIyWWl3rRoHniOo39QwiiYAWvrnDsR4ZG5OPcuLlToGXenm1q7
B4Joc206KLnbgbV1a0Qrfd2Ol2/2qIKhzpnIJEdb/Au22zNNzy16aI9vzjrqe5Ah
YVuIs9FYSIUauoI+iM4Zpzwyfi2U3bor7SSqF3akpKMgqIq3HHsAwpGnZzMI2dMt
Li8ngw+Kz9TBZYguZxKn+zfvQEBHWdWt2vHJ+m7X/gSwyJxUZmy4qfoJQqA6v3bh
ajXqjVK2RBXcwqyAh0FWeeJUHAnRWVmHpJFP4f3DD/JQ2a3VkFkqaBIVkvoXnTJs
QQW3yhEqycXMoD+3MWMLyAU4xc6xB6q4sljKEaVnFzQd/W5tfngYq9y52/G6WeI8
usuCqjqicovURZdlPF+8WAztHZGSqwHCuxrNrm2pMf4umIACTNPSOUsnWhMnUovs
58PlzrHBO+fi26CEV2CzQT5rATkDO0sVXh28CBJf6RDLj2nPXgjvLkSkW8C4g4PG
0UNh3SDTBEOK9Jo0C/ALDpoMbzp2FN/o8E/BMkQUvglBRnqnrMp7yMptMrO7/0MD
3fRogqL3BqMW3onFwVcR97ixUhHAEBLS9tUpO5DX1wD8BeI/b3YiSgH8caXyrK6C
r43FY6t7bIMfYn4XQCSTC92qc0c3SdwjraXEsqyFwJlwTF/IBQPI+c+CcokiJefe
oJDcXNz7eMyRteK8gNYuZEK58ZDyQR9E5fm3hlT4wMZuidc9iXApUeDg1ieovn5R
Qj6e3N8UC5pCJMnFVSHFoR2tX5eNqZrTtXT6pCDDSOh0/mJfzNy/FSTm8YwqhXkD
tTxzifXL6dtnmjeMHQnoeOSIieYHvhCjf71u4HiBM6L+fPCuu0Rb0DRLBlegddZR
6ZbDhGixa6gWTiMBeUOgeBYI6ulP9ROr3+g+Yog1JTqKbyx8G/p5r6NWk0zQDnI3
gv3xiqLrv3yMSjTRr9BYEkftTPEFqt/5H3ADijWRNFYudCNy0zvA4ARxSZ3+efOH
1ovxYt78yAgRy2oghCWx/RYwVRVt+qiO7Sza61OBSKGCv9zNoBu6X8MZQjbE6p/o
AJjcAZhkipxyd63X2IY6F3KH35jPFXtGBvpjGTIg0WP+tQqLz6v5EFV44I01ENIm
pSeWfHaV1q6lZ8EV3EHkF2sQV0LF70mEToyQBdXrllVlWL1mToced1fWJaM5lYYv
0CvsqbGYqeoyPBSyapbO+fRocEhYKIFVJOA2m2CACrODlkwK7OPCkrDBilDJ2/+O
bNioEB6lI6YO0g3kuK0Aof+8fNLuEEbZCQ+OaeRS27vJlcABRO24Kl81Rk9R9WNQ
0VmqgFyDW4p5sHxYroIBgKcuQHhYVUfpLGUDVWADG1O9lhJUTNFOCWxHZu0T82aT
WTDQMNUo1aECcV+DEej7Zz3heKtcu+aK43KvgJvPVoPikE+4QQrPQiM1CCEqnndt
9zAHccPoCwxxY40X4MY/ZovI8sp2IaPucC99FZwnHUQf9QNM14SwawG9QiZ7zVw/
yjFc+gxlKldoT/f/KL8SdzQMBsnMCjrQnqRCy6dRTRy/1MEnDlIYTTussAD474r+
bf0h7wv9GkIitRqyGcJ/vx2R+1HfyTeS27iyTv+unkte6WLbV5BD/1YvjryGYbaP
qtRuPrvaXKIk/boMLBJB23a/xMEh2qV2/1UQj8LOkpHTgAR9Uc0wNfkWtEIBoXG4
9cOEFEtXYBZ+sWFA6Uu2PUGqKVtUznW8BO5yzdmwRNPjG+oXaVdPXm7vXqyyl0Vd
KfJ0gES11vP5En9GUyI1rpe1pEXVmeyXiyvHb303domnSG17W4xT3hC1gcicyZkw
DXa7E6+JF9YI911Ym+WKkxqSa+48ciIBntyeE2iJd3VCgz0AH1C2sVq3/zRw13q5
oQa7sLvGAR0WZ362sGYza4OTO3L8EmvLsmjxVOFKMxNXD8dshCZGgjpuoJy2tB4V
0sSs1XfXJYzE2og+2yHim495UdAOCTQqdCUTrX/AJzuE9PZBoTpboYqzQqwQVLB5
aN6LQemJEDpJc+vcgQiDSnqjswwa6LgDoonf4u3lR5oWh89Y2W7wcnH0nsDpGg4x
o78egYeXINi07MXgMrdQl8vAuYiRJskqccX9oLTfTFgKxelBg7uPXIhOz9V1jSc0
e7NYYnxnBk7amcznFQjNKMew8rD+VpeF5pZ9+1CG7Zp6YVwUKL0L4jTqNfW/9abv
p2wSlo72X/pdnzBz+G+52MP7AWV1fXbmq04Yp463UrZEnqKWYBhkJ452AXmdOB36
r9JaHgiBQZOZMPA7NuxepvDOC1KSkLsViWgcd2OeGY/h3Wyh69olsXZi2VoQSJJ9
2DjGWx5pmw/6KLnP+vwkzTnLJ3My0L+gFC0DT+HEXNRQLoWes6Fl1JHUFFgfkIBq
m4odCWRqkJpf2FvpjNn8uepBuvoceEUq1/04v2JWqtWMNzAsd7HMfC+LwoSNoenU
Pmz4YlYyEFbR9NNmNpPEpoOm/zzxgZ7U+OkXFbTstTgEPTtYxM1aQOmIdSIoeySV
2rCNIWb+Txxe5xb5QhKuJG4cPJR+YAeiUuKl2a4+ZpZqCwc/9HEzYoTribcXBK87
jJyMK+N5sY7BJ0iwViUIQNTjSPllBlag0w8ulMGwI2ePtEtL9KAwBny6Ey9pPgHP
xDk664I8WuvyodoOGEAnsuRKEA+VT1EsKlmhhMXOsAA0FlUeiQQ8zRysL3RolyfF
gNcSV15H485ADO6qDw9rf+sfS3YI9FcOboQhkzAYuUAPYiuvFsekeei/0NjG4amz
nOYe/RCsZVejux7VMuKSI/HM+XRFjymDUvIT+MUQ0fNWO9nZV1dqz1TdumQJXnlw
dJ9SvkupRlZrmdwPUWMsIowKmFJw7nhM2THIRdgsc8SpjTs40k3kdI5+5skpFQnR
AIbF1nMr1b04vIV5Sc/SHd5B9k1XF4oZCk0m208pX284uh8iv+3yrytl6wAaz3i3
Fg5QJJGhSiMyCSTF3+qj2wpNC/1kg+6/z8DsBJX0AEgKZYr2pgpFNKxtk2h1XbZJ
hHUF9EdDBwkMWMpANlNxKpKHES/nrZ382fcEz33AdGibUF2+m4roF2IPOpaHwIRn
LUnDvjRK6RiY0PjIO/axYC8NQRFlkkDKFEOwQJm0mjNDcDrHDV+KIyCBfPf9cm33
GJSNHyCKnMU/yReXqiUN6z4p6ZnX64eHFxOW8Iucwb+Y8ac3lbGrvA2j2SpssZIg
CuDeYJcUeiiB7v4BrR8TXiKNsDmigVim4sl+/oRd7UQVK7W06+Q4vi0TIjdj0G6h
Qe52aWlLeGLVNYv82wGfrqw93R6db1ofQVLJU2K88+pQSLhRBbxmUWJDPUd4r308
M6PNr8oaWARB3ddJmsYmtXm/StfiDC086h+kBBNulGXaL9SLRQWmLCPH51vJGsT4
3OhAZhNZ7HfDo5JWd7lMRFsqzmRYrF9DrHWbe7wtXC8P3u/99PhlRPeFraw1LefB
jPfCgTV3v9hIYfYuelc4k3zRfqLxDSX8ZrXDcXAKYT6i91LHeMVGMV+17l0sfvo/
jvaFJTMH1PA70FcEb2dpIPhz0g/8pSETZksLbeqthPIzuz68xLQsPVBsWWo7OV8J
iPZl9c4/0pXOQxLFhxOvutt1gbRji6KbkAjel1vTub6I0nNyYzzAQz0qx/LcSvbS
44RpXB7q/9ZI7Z2Llcfltf1PeWdFg7VtF6meQMDiwFZVfQlSmeSpQx3XNlkm7vDN
FikPe1xrJ0ueYduC4TdEVgP695+AVu4FnR3nkPIzoqPRoC6jE2NJHnzirNDOsEXL
DqB5d12bnJTQqDAvpb3MRgSx98tQhKspkNDThtRAd0Xx7PKvL00sDoGIrKHjfOzd
9xz0Yxo/v+M87k8/W6GnTosURvpHsFfpJ9cW7AQO5uoqsPyJG/8DMwgkXbxhneQj
VS/Jjhzxy9F+d2EtEMyEYaWQuGv7O8Ca2KxF24J1SP7cfrSgaRg7GOLh6UtzqBjT
j1I7j8ODafrGIlJjHJJ03VftVgxqO4HIKrMF2IrstTFPPau+yhP/33UtMs3/if6X
P01TcIJSzOl2qUjNCrjIfoV9pW733CZR2tmzuqQZjj4WGPxIGBcmSvjr/haJ2NdD
hsyCK5yHqDdwjSiA5tUviOusaXa4KiYB6rM423DkHNYdqPUeT3dBAIEYHf9VlITz
xhsnPa6Abkly+v17kX7uD8FmwSP1YmAsg3w5hLUO0O9iQqx5J6/hIhYJRROwIZ8E
j/C/H8V0/FbEiPjS/hzxwVTz6EkqoofSvXS2U3tAS0X+Yvi6DC4qs84APj/QSj41
Ugx4ZD9fOzKYd51A5VSi4aiETwOYGWawWbrWzSEUAKaTYuTIfQUpNOQSbw/hq4lL
mzXUm3lyvEevpLSdhpyAOqyPBQFLkQ+9gsfMceJ1cpFrl5jqBZXda+jy6K1QHJM4
f+QHUio3yI/UP/J6dSTplmg6BB3h0Gg3L/5L8RPehQrKgxf966osXy9wrq28YHtb
QmB/4DaxRF/gQWAGa+yT+K2fDbzPpQDQeNLEPTVpvXQmrFPjF6rJeEvta+9L5MQk
7MJQ6zcl/2tuIqmwmsILSiz9IgTo/rGoK7vy4nCi/V6Y8oIk6Oz6W1CW/JpcmDo7
3qfexQxyXkT4ZwcL3WeXEKMHmx1ueNU383yB7eeLO2BxoGRiyy3YaWtLsaCyXYTT
YkY+9/uPKOYhQyUlP/+s9gJQZIXTXUxEtGwoHahuVstV+Tz04hEKMuIZ9y6Bfs1X
xb53znAOUZ4nIgvZzPxVLIF53zhpJjlMVsZxrY5UaMn1tLcJA0mbIeZ2JD/ovWau
sP2BrBr3G1P/VbPB+QujoGrp7OGv5hpYUGN0CFU2gDP9bC0dB2+F5IR/yYdSE12R
JIGPOGEE9NXuMfEtQ833munxyCFpXW3AS6CXAqyyuPXXSX5o9dfaNpK0LY+3167Y
UPFYh1D3RGimCHKLm6uGewaDdCpV02uDgprPwd/CsuYXQDhokCdk2H15M12tCJHD
A3srb1MXYucgYVLfsRTFjiPOZ8tvxxaFCPlq+dfwdm8qalAV6DmPlvvYDIzHu7vR
a4DYBJYK8TQp5XkX1ixQU+mRzDeaXaebLUcHQe4Iv3qjOH8KmZt6FdYQHvrVqxrh
tkt2QxcsWl1OzBqTm9a6g2ywokBMt8Vq+iXMyh6fwVwZOOGAuJXjmo379bMqjecl
+mXEGAOIeqDrDy47QlBs8UNivbQ8H6uBx/oJrPhMy//3uF1/H392rFPWqbt23zlq
RXaZ4OoL6KwSXEMX32cDgC2zoSkluj8Emrq7fqjIotrxj08YEL2GiesGM7uKs1pF
vnUIy19oK7axMlQN2QAzTBEdgStN0lNRcjXdkcK45UTawgLqkHoAtbDHWXYDleoT
f+CwuQE5XLE49RyXNA7wpKRtJUY6OmYFUpurXNh5QL+c8A0owFcE1O9O8RnKOrtY
Y9w28n0xzIybrMtJSxxqn7LpdX/ichmAKgEuwLc++BfEZzislYdo6LEaro71gNL6
IlW0r+VcEPvFaTcq8e4XhuioXVLY9QNtYEYNJDs0Gz19ngGsCK0O/Ph5fG1RCm38
yenNZPVuU8c+dSkZN2tKGLRhZDn0A1ENI88b0tWH+AwqsQt+STrWPZYrHUyT0rAc
WsHeUrRxG3FbSwBg2pNgquQqUYSA5S+iKlDrCk58O2YZ8pIVIPZ3INVMnI+tooKp
ehFq4fgda5utWva9gaCD1UTYIYAo9P8X7oHW9V3mHcgA4SoDawmuqR0bBzFtHmI1
lfPYW0F8bfN8rD3gfpfzhLotYieK2ojoUvudRogkufzWo9/2Y8iZx4Tz5Ev0SnIg
CnOO5WPLNyZP36dFH7kbjY4ZE7Z8f95M9CoBuo8HXST8fl/wiHHt/UnOhUhQixRv
YZzxS2YaI2t8DSu+Jy/AAjVLqrtMYcfBYpVFfBrkbyDtkNpvBUcvVMjjUPbkn347
H1ZXw3bxHqdpHoAXUQ768+fsE46PfhI9q/Ol7unDCblq1Hq9TTWY2NMFkBCuc4DC
goj5YCDJ4daQR14iGha7gvYGeqJVfL35PvQsJwSBpRZLm9lZI5spXkE8XLFofW7m
mJM7uzjdvPIOpBpDlUivYLe43nJmP0UvMfcYrc22lwPjV9k+yNm6rZkK9oVeupNa
wLRlXwfNbs7USobPQPMNOA0PeIkufhFOtn0/FUPq3D1IxecRPq4BiRFU6CJ5aKJ8
Tk9sFYNUgrG4Qi7hE5JpeS9WmhQg6/ui81nu8HZcVVHW15pQH8v76zx030OaMAgG
P53uMs/IiACkA41ljh1MB2LnHH2XP9EHpxDij3fx64ATcjwg5l0rEQqH5f21ROW+
M8hXkdJiW+xkHUebXS4zbszw7APiM8dR1jlSIjVcimQjLYYHB13yWNyYYmdnO4yc
bUn8fetKdReU6xE6DOFiLQKboDXgcbTvrbM0cN2KGlPxvRci1dCCjQxjn4+sYlPf
mReSzVc7Oj5/0LpioeCakWUBHXZd7YO+45PnUsERo1S1rK9Mw9NSgfoRTl9mltZI
kyD97rrh66B/jZ0tfY4xSIn4LtTlIENV1Eb8p7dE0nMJy8puSXcKV7uT6p4AfecI
m6m8ousqKpvaeMXlRH7W5+VXo3mDmvgtj46f511wlh8draTxecQtPwwqCFam9+Sv
q1pZd2Cy2pxxVr5hF2CF0X+isRHiy5JXfvyr9jzpwL2lzD4nZcAOC96bPROtlCAH
THzCQYJUm/zzuTNIPj2igRjbWQxqhULDJ8axhtck+IxBlVDH1DbZWb2r5j9OSXAS
BlbFb/f2Rdnp4w3UPNZZi96LVCsMYOJwJvmTPg6x6dXOPv3w1avrR8ripvLh5EXT
W7yAMoon4EFKDujDjLjNVk0XzDUkLcEFUKROtqLUhE/K0O4LMRhl6FNK+am2udTR
6r6dAf43Bo4Zdk5qC6KNFaOUip75TKkJiZXjsiKGKxyaj8QQ5Gil2OxurDNoAPoy
JpHdVehycxRLRaIOqXKCHutj5snyuPWeP2O+qiDxs1BB7C5lPLgBI05tZjmEkjqF
IR8sTQBKHsTD1AiazpGLY16h5yX/XCZZSkAaAPQi19JoLqPIH1oAILVBx7mq2bEL
JtvBhPONTyPWUsr1tvJrOipkaJiFbK3i4ig2ak+/W2Jj9bkKyz22LQpDp/qAoy3C
ah28s21G22bl7hOQLsOQy5yR303h04WzXnrA+dolDpkcRRSr1ONpNeDBTzunD8xn
Ie14/QGSz3i12PEvn2u1ljoHymwng09lPcPVGT8aIbRxkR6uInosNvJQjvY2LZQh
akxI3UIHgHMXcu0qdcUX0iIr91f1JSgbpH9eNETRDNBs+0S6nBi1DAXiCPqYfEcc
7Nk67lvJW9SvHxi7ysSf2mUwq3ycKzmLa2NshfusmIU7pVaPEegWMXumd8Wiwu4n
FQj0gqSNnOyxhzdQ6jr1Q8qZ9XoXg+hm+OfBeACM6nyscF2VHnBAvVpb4NCnasy7
6HuEmWpVTfBT0t1yJPerZvWGAgrYZMlpHXRzlVSMbjdiAyjIVQroADl66J6lSJWN
E8xLn6IuRFtGZJ6N9eczA+wabe8qekq4nje6JgdDDzpzy37JfIwwVKvIChD7VXen
8OWAYfForyvjyHsLUQfrIMMshTek9t0ajU6EYV92NJ4J4GA/9IbMNtVITTmzUtNQ
QSb2sTeoGmMM0AELLXdeo+nMBJVE93+gjSq8sfkEEStlK8jSZU5Gy3j1QNSpy+8E
z5qOR5K0UahE9TJW5PkdhlsvKtwlpupD1O7xz9Ffhv2CNUrC8wCGZaLVQuP/KLjx
O8RKLAmPo/z9foKz/zT0MawSXW+JKqPsw2MpzC96KvYXmV7LBrY5elKUtDOxaVWE
bFtha3m+1O/7nfIx2fswJVM+BBSbmgM3QyZ8/LlyBa0+bHgJN4d3L2KVSM1YMmpL
jiEHIagcQgMnsTdoF5msvLGGatchhAKG95KUX5fNhA9DfpbJ4tQ2z9jP10QiifJ+
AJFOA/jpQ7LTNjXPFZm2FKGAUxU9j6+ThchFVs91N6PlagiM0FGyN5yIlITmFUAJ
nBHIHOsPsk2kChPTvlBxgsM3f5d4OX618vSpjlmWnPyUehG72jeD2dL9303d3G0R
SMi6wPluJx/YX/cOumrw6K9Q0GIZYzyQuoAaVOiQH1mmXI5cU0+znLKumyNel8fy
KmyHBpOnD+Inx7QTqhGzjMNGpfnTxynjdZZX41D9ORsrlBD/E3vDhzIY2bgJyL4E
g1V3pSrHwFe/cpT1M6V4SJjMNr/K52TdxR+Ae/V0iBzEh9lGEJ99w9jDRygf2Tx1
I3wEs7bdDnPc4/7rwAb3P/bMYQ9ZZMKzfianMClvQWLLQJDL+3a6SlZCaFyLFYtM
c5NcKINolRxGzauSNcQ/PsCJlhbbKjg6A1e5e4fY+5sgi+jEn0drBIZDzdxPBM4v
XKquTSbz/P8BFRibE+NrQZd+sNDvn1u2pne/AFW2xpu1GavCJUWqKPMxPiNl3Icx
8x/X1VsUvUMaU41hHCWzam79D0OgMVb6ebyAYhTc1lnmqlHRk3zyMuILpLhIKGGN
vgwpSQc0/IGn3Lz3XAIWZlUo9sRiHjSUJ8Xe8AYquAr3nWG2xEShghvf/s4oI1Sn
JZN75cQLp+lY1rDweP129h4NEDN2ojxlpF9xIWCD00YITtkkY1/L/PS09JXTGy/8
l9FQu6jKuF+Xg9jMFuDEg2M8ngQ4ET0c4zU2UcorICAmvB8Cw4kshWtR0t4AIJPu
9smTLrd4w+0IItTNTaRQVf3P32AIiaDBxht3TgjJxMM1dQwF8V6+eyfD98jOGRjn
E5SZdHYZPtClgmNcRhoy2Dj6QVPH88rTf8vZxN1tjCWPZVAz8nQCkVPEsPQayY4X
EtCPFzCuzzVhmKhPi2kRZv//wJvDTFExRr0kjbVvLmQPU89uZrn4QAo4KPduUb/Y
Di6un/hzhtzuBP7FCHZvpAXeiHdRoU2CsCa7lGmdQ6MlqbpUTA7s1FZWLkHhkZjD
GZU5uqUFxushlbvxq5Q9QZ8OocXaAeh1eU+hwqrx0gMfclVPchJuRep2LjgfQNpy
+1+h7bhLOcj4C5BOLDvUChaMiYU58YqDo2CPTW/3crbgIW5RfVd0y+pjKKtUMMzj
//v0dAFC0XuXvEGjKTvgIl4mD5uOhLqPTG/UhRoySWfNc1zEuycAfgAjGEg3MY5p
P3u/dVRjYgCSGbZRBAP6ya+wz0KHtDFRiEMhDM59TlauKmXpWpFkcDRrsuCFDxWy
ZvyUIQMYZ07xRnu+93upADdKG0S1MshdftSV7N7/7hQrgJ4OzpySUpPSEJ5GhUB0
WMDdIeueS6ClCpqvH6q6gXjAvbDXLs/BiToW7lWyX8UqMa4rx5/rUQDyad0X5K2k
fXDLavMtZRSgCm6O7p0Vg1CpWYYa+hKzniVEWO6OGOtobwBYWtmic9UcTA8ri+4X
UnE2yK1xGB68OOJLvlHVxlvhO/i6t7EhXA7AN+T+G7HN9kTuYW5HOkT/2aFz7lCe
tsGAE7398cX+TNiWsi/bYb+y4QBmizgQ7woY0FNOxd9gdI6kNEXVGt9LsG2t9M4R
v3Mt1woIQobbvi5VyYZ2YAkwMKctwSh890uDb3XQlB0C6d5UJTUTVvk/r4SveZSh
p3h+UMlWzDfN1KIpUv+kMLCKuoADUfydfix64oXDRDFz9tFpGHWY7ctngO4bTSM4
ncb2nH8PUt4SOlA2ZTeYDiJ3jAn5D/RlvLyvJQmNlvc83/2YhySf+hkfGO+EfJVo
oqYFdklU5JVfDwqHPfpaKINUXZ53mkKhlr7iEbSLBMNJP2BL6ZLrjRUCBpq+Is2+
RGRF9EeTTfi6CH00UW9JF4BcfHcv+Cc9en95gFFalnr/6wzQ4OnmCSS+MqYfLMn9
1Y0nqRz+5/okiSZLAzN92iiu9M6whX1dWX55lurvwOVypA19Rg9syxEy3ffYBzQG
4tlkwFHO0Q5NtPOW/w7PvDh5Em0Yo7lQBluD1c1JaxrQexVwe032JLgFeDykLSqY
ZLjr9tvltBcG90+kFpyKgmfYEdT0zkOKUjbOF2GjhL7J9zUj1vhPvoriYZ2i+ZXb
T/wf7OHki7PevIxkO6FDlfu7Bnqp4/l1OdcpVSX9Alci/QwCEXCMiC3SOA7oATpe
5qOdt7TFUJZncifkxFFZeLDkHMW8zzkZG5Ch5irCXLNwP7Z3inpmpkUQQA6UobzQ
Iu/7wFdsKndgCzNGa0nGeMm67Wc2RfPDdErQO5vjNosNzLvTBAU3o6jy03tSmbX4
SUl7KObV8oH1jwYdtwI6ImgMP9HTJiI2iZMI7x0YuRgEYT03x4xteUmEngpfndXi
wMDKf2d89P0xIq0HxVOfeuQLSMntKz+TDNyX+m7Gf2AjH23KfYlDINrggptoEXQt
4BEEAS9ZPSJjg0BBgaaP5q2xIemjefk7OWlnCIHpu3t/rLm1HPKb8p0kXkdK/Erd
RP5OAlbHI5Ff5qgZjS9sJGxM49hCUpmJEW58RTOD9XwE5BnqTPzXgSaLO6Hm9efh
BhhC970wPNeL5kUEFjOE5sQmTstng1rI6RBrFZTNm1u3c3O+zja3Yf1g8f9ZCtre
mlR4tmx7vieE6IyQbI2yLETnAjvpnu6YageBQhZxNggxAagzd/0OTsoPFi4Ol1WX
kYoOOu6zCkDgSRImlT+E4+4ZXqtWH7bxpdCR0WkyTpTbZv9+1BiAA8P7zA5UTWlS
NalFNY9hI3a9F062BbXwkNXtfoM7m2xcb01f/O7Ez0qTIF/k7qsGQzkSftzGyEMA
r5X6/HUXMocz0+2WUuX6Ja1EVaoPi0R3smFKfCNqW+fdlh3PaCB7o8s3dEOPYCyr
hhhVIi4pnJBcgymPARYrBrXvd32BwQzCMIJTyz93FaOI1HOsSV0yEjVhNQGD2i/A
GV/ckzb10D3+QB0gR4TvEHiB1RlxjmxfEv+JtU/NNVrWt9JiEB7LOtRtG/yDg2T+
r3UY0B4Ze7DY9NkLmhXbObA+4XAWEROY5OT7bmK2zOMEzSSVYmkHDNQv5v6/aTqp
4UA2ZaiIkJTfkh5Lp23KMGkThvDerQZzWSUT1VSRlad5Qe06qEfCy3R3b/xoOd6d
QiTWE5e2zkh0lIxkk54wGkf4Z+SwBNV0uCqzyDWSosw/SuaqG+CFD9cjb2p7yUTM
OXvKX3MEDZ6CsoM9uFepgAXyxH/D3UeqOXWSb6Do9NF/9GMFeUOfClnd3Q5uNWku
IqXTd3mx97YhL8yW7dG8strbEI3ISWPOSNj2p7j5vDyAozWNckKqVsZp9cOwzZWj
GuJlPw6TCIERU+1ZtL56cQ/AYwlSMhWdQnPWJjqFI5IxLOnF44VhhUDliiAJsj34
S4yl+FY05E7aNtlZ8ivGGHaKrI3VfSs5rQW/jjAIQ4KPtg58Bi5gqWbpLcdJZFAi
+Rkx6nJdo5dCB9bF3tyb0bIJTXLjA++p2vz5yCJ3jxVVa0q/g2/QUUbqymmHIyGP
SC6SB4un6JhnhvA0U+kIMnT4z0THAuORaxWMBcIrJ0ZX9H7ervs0LVgFtyLNyjF+
wxLtp8cQtcmLiLpCmi2MUZAaxTDTPM7VHihf/hhkR93ed3otq1w0XQh6JV+TEfLD
iUFbEfxTbJor/cArveheXsaafRuLOFGI1QdW5Lz9p7S4sOS60RVp9ciqWEx6/Ejk
+z6+k9hX+zqyqc+BGn4lSudn8cDn1L71HETElYHpZIkRFcLwda6skG4BDRRIYFgR
6XBad2q7vWd/V9D0H5nChejLWiRO5Aya9Sf40QaSzWlxVUQh8T7V8gUZ4e3OHKLf
RrPC4i5TP4Ix3xqoMUXHoxkTKTs6Pa+PAE7vqGvFWCW6VMHVokmFV0vLllEBrERb
m6PRfMVBdvccPeseHFPi2mi7ivt0NV/TJ0SoNdfnyjJG47lKLAXUYSt1am0LqjmL
2HZqc1CtJIYDgMQB8KpGLqbN0ZDwHLwEhxt5WcxwcxDq5jqC2WwMKayGcta2KSjE
RLKRPQxQWRKUgjuOAtV8GeJmJhjWsjcIhALp07IAYDMO1QcuWwzJEHJ2dM9Pa1FE
sUu/cm979jGLDYgEdVQKMx+nxu+o7BWRyfsecJmr06IlSwCmcnP9eLKmCpmzZPR5
3VM66LUl9ao65uGiOrJa7bR7YWC/NyTaHDZ0/CqWgl8r+xBoaJQ3b75AAxHJJxZq
YMLBCJlLJ5qp762V8trjUDUhwSbfUWPVEjX2h5YNF5VWJ97pZMMM99o4ErqPS1+t
GmGNzsIWVUomXne/fj3NT/AqaKLP7LPXc0zqWwdY+DdGTiocbDqhrMwQcmHk3Jo6
mP0MigPojc5fLomSOlgQa9WlE1kDwYKXMRdmhnriciVxtlLPtLgbYkmiflsoVvle
Jbk+KYZ27tC75LKHJlnqiNeYIfsBMYS77f4eeqqwicOqR1pLMhb9z5S9g5i+BG38
9X1a3fWeKKuxtdLQymghx0Grxf+/W85wubhztkxnXNFKTJf+zBmEPAP7n2l7mKqs
esJzoj99FKHzLmyMYQQJKKK/Ajp9fQVuNPD8ya3IllQfeRRKN1Ll3SzvD/dP9DhL
B5Uvxlpaqftgx6ncD7mhUkB/5+RklLS3fXwzTqNaPRYYI4dJC2Uog8qd+wBhAiOz
d4qH3B5xTwtwzn6WecSjst8z/MbAItGN9tDXsXm6QWwk8DwNLY1KPzRcOWwa30si
r+hiWH4wLSzwq7z2em3wRQtwEv6wg/4Sd9vAOn0OrIHJUBCuLhDoFEeyaAs2vMoR
+DCW6Nikfc0ZSPUbfM98uCJPrQBJHlBkVVKLbZZT2JMZaxmNYuxxpNVcJmGHg7jH
ZwUlieFGJMfSzdqGgHXNxWaGtd/03mVE8w7IlAdw9Nya47Hlzy5vbq0+02eKbbHq
vIu/zD+13h/GDgUPUistP1w9nR1U0cOBg+I+WCUhiBK4A8ipzaQcjLA1N2VrfZ9r
/PajLjXJF01QGhrQn3pKyil7ql5s4osa1QOo3AP4Wh19Hll8C67eIrW0g++164ND
YuPoRpLD+GKVjz9OI7t9o+vg6pO5QJIybPITAtGCBNngjE3ofwZVTSC5Kg5dq4bf
tp7RsU3OdweCDtloHSuH0GCNnxr1igUJNMgR3ZazEILkrt4oHTMclXg1gANOSyCC
nFy52MgezKz40AvMeMggklT6vNtliZ9RBD+c4w58Ioz0RbTEmQNzPvBD3Y2Y9zQP
/GP8DOvOSVm1LhwJpl0eaBZx6puWeDCn+jKJUAHctlpzOICkWe32VUfrIqU+aCXG
5/ndh/eKfuHKVNZCV4+gHkigE78SSmQ7mHUK75cemYJLKaBFpKY6sNPEXZlH82n9
S6ulFlwg14H1iEVf8A1SyYq6cN7VYYYO2G/HMBAxQ5lppo7OT5CbGoSHhCD3HTcc
+bgAilFD30quHpgKC+WpM4znF2dONd7IUj6D6gTNgxFVCFLFXUrSc1qXBnvDTyca
HhkZPKBOtl8gruju/dYeJwYzf8RSGkH19dHV26iW14Gm4Ag57qYOJ3FIUoYmNsYF
poHH1vOTYR6GDOgGsxdXepEP/yBWXuKpb5L1Cd51EWMmwB+ORJS2b+OKhUXyM2bC
1eb966EPy7LjN8DoKM4KDVTEI902DQoiZyfB6ep4XdpN3ioErLukia8ExDClZXQn
YETXrVqWKPLD0vXrv5eguLwz/O5xScMeDP9CwsBf5+98gVJ3jzJP6NRKYJLkTva+
j8lVPji6VmG5KiGX0Fzr6+zSKNelNG4pj80/YsvcXXLSM/IgjVVZNy67YPdf4NJD
5Ce56+uO0H4nEZy3JDvdrEtBcRiNJTdAfguf7sRfP7JHOVpvZXoY0aueSm7cimr8
MjXtrtCPVkLvQHQHRVJRYFhirF/2fqjEIhhjJfnWWGGUohmYFpm1Yyyo9xUZok3W
8QNh+r8VxYOHoDuNI+hKFCffTeSLj4YUCGO3QQwAVv03uKSM+FiQeDExRSW3Mjhl
ZIs5+OvXHoP8EFlSi/pfIphbZQ6ATQBAeTqi/9Z9tTf77tRf9PxIvwxmxJTXBCj5
GW8LVzk3OeVFfraR6WLWwllMKJ3e9dTwnZy949Mpu7ApDlNztNT8nyMwGcTEFPik
YgmtPs33AOvhFb0ezLOzcSxgN0rQKtzX9GjjXu7R6B0BJ6yGumSdCECd9M080VMh
+Hu2jWQMP6VBYkFOLgrFB5TSezEQNN0/LZGQdtyWxO1RgPzM9s/015OO+Dm3l7AK
/33RB02QunKYrxdWa1dJWHRJK5iXeaJb1zgfx9wts+LDnNRI0qA8VbuSOx0sIhk5
fC40LW/tk/da7X60DiNuZH9PF3tlqJAoOEF3Bq2zMxi97kW5qeMzwBFs1S6QfXqA
9XQelLyIHmDTyYgcfdJZNPc9dPr6ah/Y176peQl0Nbka5drbaIP7XygHzA6s3UXQ
aGE7RnqNTLJ2R6I7WDuqGhyxzznaTH5j2nN1KYAU2QvtvrUL5EoqaDmRvCkOxlXl
oMQ7w4NMYrbYHGD8oHQwaZDauFXOulqiaUC4iQQKvwGHCJgT8SO09mffkqccM6I/
8LHT+noRUq960GCOa8j5OBhN3kXuyFubgIyr5d4MQ0P48J6bT7k6tSu55hBALQtV
1v1YFUc4LDjsoQJ35uD8yO2rjfsHIECUmF5GDcB4070MbUrvqhmTucX0RNdV16ob
wVzaqLWfEzei+UFNwtaatE7Nv3UmZT6gCugXhkSczMJLDExv6dgu4PVgRpwb9yOE
pdRzbWe4X/O1VAsM5smcdMLkwKeXO0mLre8/JF1s/CRaSwiJUT0uMfHfzXPfsRCu
C0H1wujrLmjy/0iuDNtOqsIZ5HQ/t9mUozKJIwa645i36gWznhUP+dpH9amDePQj
3lgwDb/xlFdvR/n8XV3Qb1x2FVlGw+BgsQt6pZrNLTzEF5y7cpPnUC1NYv8fSnDI
D+H9zSY7I5woQrUwX2hFmRIlmvEjbeSJWopPNcKXUqbs+ETyEbRVvceh3s7jrIoH
PPUNpAf6Ax5gArZhumAfO4551yStgbQEm90aN7xnoycYkIgxPpDFanIadDEN2gF1
fEtWXQWVpsKajneeGVD40XOJo3DescSTUlzLzYMrUjuodegiH+OiF8FJakEkRClF
18tb0VL7O+ZMdP0uuaKIXV9yhr9Q+VhHzExgppB6rutgPqZXozgegIoFsdklznFb
DUX0lwwy+BYFHI5xd5LSLLc28NjSt23R9gIjdHEx39Znjn6WOH2SNytRxho+wiSK
5Avxy7XicEsruiL5St1AJ4tlI0rWK30sbju98I1/vgaVPVJ8eIO1jlyzefYl6867
2bCdi1E55W5UTEQ5DQRiU1zf0Z186J5G4updYpAZyTDQwIwSaaGhCvyGHiLojxVn
Afm/KcY16OB9sELspCC6ZjxOE5ZMPwJj3ANVoxrcBl5D1SLJEvBc8I4QH2xvA9Fm
k4RGYi0izEu4Zq0hiFJNvQkx/D04mxR5LtEqBjV/rJ9t/prfzuN3lxkW0Bb6mePu
diKy8cYiSiXAuC8Er+0F9O7nPHD7m0owy2A30C4vKmxtzStBqCVVckAB29bgq9A1
vp570316pPJevF2o6/zqf2B9Co1eedyERQphVeYyaS7sxxHxeMmeFZfc09Vhjtdg
s2hQmYtm189CPyjVP+M31iXmVgsRx+UPzu4QYlbjWqKAEk8O1HAIJ0Trjjm6S3qd
kw8CKHJuuZousYwzZ0A+JEFNsetDfVVq9pXx0FjwfKZp4I/u6t7tPtHYeRYbIEPn
IIB06cF1ctodOYuWj/hHIzDat4ygSItlkleMhXGohlPRV/PQ+eE8lQxJe4/9SlV5
0AIok8eHxm+ZtIuf9FIGcbk90XCkBlkZnyN5au/Yvz5X2khMhlCC0s1YL1xtyXGj
lul3NBRGMQa+1HY6GgesJZZUcfkwpEy2BjFW9PI2jdpDW+XKugWQf1PvBV5XDGR7
kxgwUsJBUQ12BQaKbJc4nbUDYHc2+4NhIJL9BG9n/yuxpcseRCJkbk83cpQsJkyl
fkNX+XEXFTDXQWje78jaJpy+dzV4RKSO5ruGyyAvk8KjjmXW1qycBjq5n7E2Oj50
gHoArX0F00KTUEnGfRpwd2KV12we4NBpypsbWHWbfdF+MRt+JJ6L8Ga8cD7wWx6m
TfR1rhbZbpGTiACQx/oqrD3KZRGfGhviYpmspibQpcbrLe+SLxgdu4/vWU82c0Hh
sHDFjRx5ZRgHaRMHW12Z7JyAmaDknGVxUCpvhvJcntlsD5+zb764obXpz2sCyGjG
Lr5+7NcpAX5j4CFKWLc+Daw86yeewK6XOWDl9wqVJUWhv/a3GR/I3CPQjcEMTuIL
3xe2IuJirgDK2vIAL9CvUdwJ+Cwr38n1O+FPWVR8OLWIWIfLWcyOsTQS36Ad4sF8
riDwcKdLEf1EP+RU5BLSf0I67RpInenDY5pNCcQPKBevlxho6AC2XNtgB0xekSNg
Exgj2w+BBhbZoyr7b6WGIMkn065L52o34wsuYQAB6y5gGG3YjzAYwAwrDhOEdAQt
kBYIkwxmUPW63ir7PlR/CZwX/CXB1XG+Ncn/xl7PsKWRCUjvUEAKuLDx0K49y7gO
5vu/UCeaTACXUwNiFwVQwfSrInD9P/a/sNtvUXTAM9OPC1hjnL/0dSgcMhtKU6Y1
ynVSUfCA7Mumq5t5hvVmYiUbWIa76zOpIZFmMVwkyCblMLRaJBPMzP94AKGNCEgG
nDdftOgO66UQ1Dg5TICATixfAn6mzQoWYnhnkVVYoqoQhZm0kp25ABt+rbde5xxd
g02NCCpb8r+nzN4+koPKOQAfWuwvvsWilpY4Y2zHZ6hO7fYRhJ0NLQQCvtHqsIPA
jSz5uaZEayQ6eQl4potaSI6ypAWSrJhwLHoyMLKdv6jfqcGtJo7ZsMQTqYf8zp3J
CHq6k9BDLufLgyARiVXHnfVxaublbfXGxBl/PiVETFyt2coJavVAJL/0o/pCdTfL
cnfnKQL718uM/yfn6u1IaBBmAPvxI7/g9G14yBJWlYVhoYbY2YuBqcciw+/b6sXW
3oE7m0YKLrbeZQhRJ2ac70NTfUdDOKCBss1gBJ1YH25AKNKIelRtPwkOPCjcdGXe
mu8ZY3ht6JmjZnMELJJGjMP0qc5XdhS+DUNfOhjTx3kLbGZ1TVpZ6a2x0wUf8j3U
9zr2bIMjUPJ0RFi4LflUoKv+U6DumJ4qrAbBb6GYyOqe+jMCoixifYkGochV4Da1
N9dRE/oWMxZFQkJfwb+7Kcd2ZWOSOgEY0b44Q0DT7MgOvT8LkA/u4LJWX9QILqK7
dLk8qrQSQOrt81RsUaNILjTgWoXZzp4IfJRh/Dq3ECWGVYt1uJNfrHChz23xePdJ
9GbOS6nJCMsaSGsB6+s+eFos1XL4rv4NJyz4NEcfNU7geNdGxpN51/rFiMwXvYkO
EAa7yFSvnVhxM5CWd6Qlry8pxnp/oBz6M1oLjc0xLKv66UMWVzxA09AktRFXURX2
QmSUTjXnMdPiymGZ8QMh3VdqlQZUOLno1ynuvoWywKNZeP6pLOIu7/4ngHxs8K6b
hnu+R6TMKK5Ilhq28g5Kq6xWIicYHn5WZtXYq6Bh+hJd+OWfLRbgWPPEQtN0dZZY
VHUWp+YBZfPUBDU6Ry/gkK3TaK1DwzPg0sg2lDxAcYJN8HXVWXKjo60kE+OM1MB3
f4p2xXKv+WCCfah8e06D643Vb5cEjDvjrbcFVY9J+u68XUg0srpKYTQ+VkYdh6+J
BLuVZpwKnZaI69+fIEYXwXQceSohf7D6iU0BCbzb3YuFdvCCy5GOWyajxMmpmX7n
UOih0YrhutldmJ6zhAyn+vw4xTXHUlq69JLwDC0q5HQUvhCZiO9MCIntJ3L2N4ij
+o4Aas1L9F/QMfmO9W6/1CT1AMYFLyB+zbxMiEu+gsPi6LHNEBCGdvg/f+21iZ6Z
bLaUJHzxTfG1xl1bsRE+wzNuRVVQK+Y+wRRUWnoe2vIbrhVymlPSRv0QTTHsapo2
vWU86PWNys3jWfZfGEkKXDWoLsgZoBVt+K74DRiIPGJ7PIfQit/qraMF9MYPh466
JLAy0ZcXHuUWnKH12TO1gQqrWHuVhhpdc+XjZuJnbtqoMqKTbh5Lqn90UxIZM4ve
3shbeFOkVnojCGBshhSnJi9Z3QbWmn2Fz27/lSkGG2wzhn5mIVmGDBiIsbFkzBKK
qhTF0kOWRqUwYzG1azxLHH3BJG2vTIFTGQFXKauXxfOiot1ATpIcSQzairTyQR7y
sQU/YMrA5kkcSC9sZhcdapPKBIR8gSPWxaJDZeW9IDryrzeuXpYZTMRzc5ZaC5Z3
vQMseHuCqcHC1gJLfV6f8rZc/dcxuQ/zqMxltpDrZcWuAtbn13rQcB2EFTwGNDvH
6qWEDejyrldQ1ARpS7Cp6sMN3Ed3FhQV1RpRrw87v4D09pqEqjsMsePaFgndCbqD
ml2Ptb38E7OoJFvB6HryPKhPfQLuXMC6rHoY0rmnFx7Sk2Yl5DvAFpt+tKmkDPxg
WMrT5dewBzPAY97wDjh2+QOydEk6fLGo9ijegzpDDpv/ayWPsesP1VEh+7/VwnsG
IhnkLTdsGkFjPR9Fl5H/8nCs1eNoitnNnustz4s8nX1IjGyAQ7dzVaqMLdhVnotQ
hpdvXlW/UdaQwPPIFXbhbReyn7OP0hChEOTa20E/tMGWE1C0UkpRtHhqoPnC2ETT
03ldi0nmYEejQe6aTlR7OvGirQZSo7EP+p+0TQlSlN60kh6wVmnf6ieVigds4TSw
S6Ze/gvZnALlAoehooA/FpES2sQvD7kHWyL0lnGNrjZsG58ojOInknb2Z3FGbPYs
twp7gBp6Ux01wnK52LwCuXkPCLY4D0umEXS7jbXA2zP+1JNh8vfKMuEd5WV6ObM9
o0zL3jtSyaVyK74qYAy3JYyj6szavCRC8mmflS9WG5fDNSmxctXZWRtOipkDdAea
/DFmP9Ap+LyZOUb1r7Sgib6XefvEDM1mTEK1fPGbh80h+kMgs04eCXXsmT9wMalJ
IeTRXcAWoRRt6yHPKKhfU/bJyuk7Gb7UFdsXuUo2eQz3xi5opAgGThonQrJPw8DZ
88nm6Afl9bVuhAMebqYr05McK9prtp+Zboz1tEfzA6OAciHJCCBm9AjAwFwLj81p
qaaH3K2w30cKW3q4GUR4RFZ6oXBi+kJiUyVqy/pVN87k5eyPTU0bCQVKpVhQXwBr
7zb5w+9AePijysQjUAvEay4KmlwEaEaDOtuuTg044P0YXUunUwKu9bIzfg9haQpl
lwyFtjVKz7zBcp29WwcbbjZynaZAgpNN/gX0LyuZEY56/R9ImuVNynPxOWrOOmKa
t/m5+EYlY2PQczVpfVSKp/LpyJHvm4JN7D6Pcbtj8uWBQfNuY0CWVqHfxynKI9s8
/NGMryk1003PJ7I+1b3VuGQqWgVOlhZ06bnNQ1zY/1t4ATZnWCOXV5necHN8iERU
+e3hYnOQA3XhRKvmVwaV6phL6tyX2sqBweGtwc2VhZhGWzeMlhuEsazxVWwmHV4B
DMyUv/i6gHQbeA5swaY+0ehb8rQlf1wc9zcD2jg6nxBg+iXqBvn8Mokomrb2JUoB
2AOn80vJ2OmQNDm/HiZQ3+9G84+bxGdSGNG97Uwg9pCuRwOorXZWk7MuTFWzjV46
oJeRIwpj4XmoBS9utuMCi4D8Ungdz40UD9JFZAxwNstMftZ8YYXqDwp+6MT7akGU
Pqs/lZzf2xPFaa9XQPA6S6+HLApmMe3FZvFz+WK/U8TojpWkzNaH9kqicSO+JlZv
bPOcj5khKOujTxl6nfQ6MGgqWIRyuUU2e8Tu1avB4gGWzC0SPwERFMJyM2Iczgpr
BCG+FS11neMKTVddkd6QSS/Bl+aP+Mko8sllE8xZsMeOs3fYkFV1nk1wH1pmmm9X
xF/o08Z4ge77eVROoLuKExFOAo03O0zPs+8JRQx5prX4ju/95MZA2xT4DHzROqZY
XPISYVrmftcb2jJhomrg4TW07HYwa/yOsEDb1SvM1qSnIWYcqE8SHQhajcpb7iwc
RD+ZLx7CYxtz0tlIK0KiVNdNQDQeYksK7fyfslDbCkDQRE3C/HKF0LbY3z5LViO6
8Y4jTXEjZ4kQ/NqkKuxTw9MDt3wsCYzpOAkoMEesm8047+KhTAWvkSwYFqSfNOO0
9YGytNOl5AGIzaCTD1gNo8YKYKPgqBTkYspKAtQsFyeCgDmK8qmu9+o+pd7P7vUH
TyMdgjUrPzG0sUScDRod9Pc351Yn7mkkxJ8y9s57VilDkU0EDWNArMl/hifaIbkO
H53RUqG2ZX/0EPWjLx46hUUqf9s73PdcFxmb1A95UX5myOrqdQup2eC/hQXtGeKI
ENXEJBhd1oqey9HD+uOgwrajecYxG26s2/yfv5zoGaTiVmLSkGXGx5iDmwWW42Bd
rNmPD3DWyF5/DHkd3FxWIhZqIJF449uvZzEMd/9eOi25JXAaCetRsTtT04M0UbjO
GKOFwpO81ntH8CMbSJbdmJgqiSxvapyj9GzVeKmw0JUIXUr868obg7TEAv2Zbhhu
ounsMOEUWs3AXyZ9Y7c1j5AvcCIjxl4sK34MYY/ttGhB8zjB8xXQ3bv8oWELiZqX
TtRatEMs15ls80MFsZ56uGa4sfcjYL+rj7rALP5u/6mTT+ZLSjKKhafGqiLBf5GQ
pmmEFuXXX3WCkjakKtZ9lnSNFBLSLxsXvWqYU8CrBLGp2jvCp2pj18tzIaD8mwAw
wHnGIfcnCjFtZgtLenl7kRRW1jToRVH1Anr7gSb8oHC8pb+879t82HadX+lTuEEk
f0IhC8DQVKeOvuRiazsiY4WjFtnKNi5t9egezsbKUz+6eqN2SdTPtfabJ356JZ8i
0jMRP4aedjAEX+px3dMtLNvbqQsSg+qg5m44JFAabFbLte9DThQTQqlaI1msEIbF
BwKHvtUbSjvss1sl7t7K/9OcKcOwcij/O2cLxn42QO3m5jsfHt3FumZ+U//b/74D
RDHFNhT21xtrOZ6zrKdaJrQInGbNtQiLhTjFpNowaHUCHHmtHSS+2VE4POHGMBjH
3hVblZxIYLeGQS3F/WigYcQfvymtRV458k2k7l1BcTZL6Mnomf5AhsIMzH8AOv0V
OfSL6oRNk6s190qhgw/7wXMY5nuNoXz0SNPXhhPCiJpZMnLQF/MkksmFbQamHtaM
gc4jhcSe4YspgPyN4msmwXQdtzPKr9W+HYu+GmIwFMg8b3osDn1kLG7Dobbdctc0
BTVllI1sls5HYgqgPHGiQitOTf0MZYVYlnhBwK069e4YVFn6cjxp/fds1UuhiatO
0a5xGyKndDeFXvyyEz0ce+MiQK954ZvJKtvFyrlFq53us7Rg95swSTAEM1tW3Ypj
zTI4OsFo7+eI1nvDDdyIuEZOzxokBxAe8/5rFGAGXEWN3dIiQyK4DtOWF7JI1qlN
cKGFahgJ6GfZw6WEUsiRRD0Jm1Zh5JqMRYX7gDDaGhIK8DLvliKUiOLoQCgu1rmG
d2SC3kLu70EKzEPsCh4BeZCjT8lwTMjQEiYHR0lYlbtp3gGS5SmKuBdC98bMNimy
r9cPcxluPijlbidW8RmGkgbqll/zOAIqXfUii1qg7J1uqDR5jTf1pOJZV5MZaf5d
RS32UJoZNL4/aJOSyaTiR8fU1qKg3zMS5RCC4ZTC8WjUFoD1fc5qKVqxJWlMZwTL
4cze1BW/jlwQmbza4JJ0MmdQTc/O6+W4ZAwhBkAj1l/90PrHYO5KgLUady/1Dn6l
YCVKSsuHILW2cG9AawqwBgxSzkxUWumtDkm+PH7SHvXSbuoHyuSpfhPMCKCbkvii
FLonnMMQJaMq8t2tC/uUejiwQKeQaFYTOwIBldCsjVj6PCziqHTivFSB3D7YbylH
fMwFo2tRP8MQmHn0E4u2GSlamGx0Xhtfvx70UqGYGn9O3v6oOMAuxYJpU6wJPl5I
slIQsAlsXIxn8HCYwDrWR3CpdvX4OH6HiPEtUU+BNAtuwXDbVZ/WRVS3ATrBWQ7E
Qwg8BKorjb5+suqGWfg8gdHTSWO9pJUuRhUYaWo0uUelur/juy/MZOgOb0jCFFCN
htE1VGZRWvD3Hjgx81iOZVZTbZ/WsN50OjmSNTPYJNAEG6BPA/MqMPKWYA5mfvGn
tvPywh7imdTinNWLea7O6SiTXQFJ3lNqBVZA06Mo/B5RCIBU784eZBi0P6R7v+Kd
HU7MF8xmxou9vUvIF2PyOH+3pTNVAndvswppUqpHERwMdbk2eaLDKxrBs0p1SOew
lfzHBEZbPaf2br1d6E/zEOtHR3cjVscZ3YSMl/n4VI9nORN/SYswfYVgTC2ovu+p
Fkzg5sG1cHtGY87VVssUeq9SUIs+CnQ8T5T5m6Lpo3NurVb/KoZAdaAVc8OE7xV8
lgk05YDZsfN34wKEy5uGZlb35C0PgKh02OmiIrZ5qCK8yOReNRDCBTjzE9ejUnUP
kTM+KUHxDX7xCwiLB8PV6bNfPRGWhlPpSIU4JfVyLBhJnR2iWvdmBqjwhiM0h9sf
WDTg9LsVWvdkHjrkhmA95N+9a6WXZ7L1Vq0q1ww+NILUPu/zM1g1L/TEZxeazNP0
dSkvEgeKwlfIe/6PVGNALQ6hX8EyjsYFQQ83+ozEHYYsQABWJItgmvSFQ8CfUSlV
hYXkWLCqd6lDAGnqB2XuB3xy4Oof8D/KgzJmnyWDI3y2Ro0EgKKcxNsddAuVu0tA
lv0zYRmTuTmr2Kw4QdNextObH3dQbEOj6l6dr2NmEgetbw8mzuEWmLjEgQPZrIXK
pn1CrDLU04vaxXoMS0t/tyTYdevXIriRTzU48jm0WXsDD83SNrw9vh1Pd3RPBKln
HCqaGiWFMjU9m28XuRsg7NWck280Eb3GI1DPL43pXx3DvoqI12l7qKe2H28Bt7wy
X7vCEjk0SUy3GvFGxAsbTGKkxjB7Iq9HPBXVnk+ldjXQ0+VIJbBwlh6Pi/KIWy+m
ZfzRo5OJNdaEnqPxUHeb7bbwRZMn/u7kp5xplTDgAK7bIr5SLwanRsgAxlfCbHV1
DUbV7Zj0AqBP4bBWyL05ixj+YrYamUWLDiKyccaQb1RNygbbrLZlQ+yNC8uM9A4r
726oTxUmZH8lvIkqNNQWnK2RAdU3sYhos/PGAHYrVmukBQsEPje1X4D6dLT0zYqu
Y1N7NfTVOoVlPQ132vWFP2cu/k3Se8oaysgWKQv0OOuhqQDepsMOS01yYVzPxtU9
nJQkvg63u7VZJlgAeJUfS1Z+jJjj+3ebsw12hW1DQVucUPIlTfg0ViwdOgzgnfyi
W89PwOkV6GU5BeoxFlgSXwzkcyPRWBbutMHwg49q57Z0GupbcR1dD6ipjoMhHp38
SQCNCRX89jOlxVpthzAEWC4N7kMbep50VTYjp5EYF12GiyjHreBKVaC15SPG6upv
s6oFI3wizVt5sMF8luLGHuPYBppdZ0PTir3As6X2raKW5IvGwrKx9+DmlOky+++V
hajB52diNcCCHGRn7UZNKV5Fz05JzLnx/raXlAgQGvOnuR+EtJZp8xGIePatWRTC
bssb7VFtBuPp8YviMdb16+rarb65jPVBA/n2K7OgKRW6PZmD0WLaSYE76+MDROwT
eMZ6xene58gsEKm6nta7Uzkv9Ihfz+UCDaHfbTdgw6G4l0c/T0iqrjmoO/SEF26W
cO3p0FicVvwQug/M3lnntDRwm44oBXkbcB17wMbtLrWJJSO8IK8Oh03bHMw7KEE3
ZE2uuj3edGOyv3273g3YSpGez9DkFyANoFcAAO6y4i38Xo5FdNB3H7rvAjJ82ZHa
PicSxd/r22FRcJl6nYuLeAJV0EPbmHm5rHikXX5d9kaU/+kJBneqOfgXcKC4RFpJ
oq/fgQDfVK/+ETt2fintH3Eyu20r96qcYnDGW63a3rBIa0HIGNY3qjkQA9xAf7oL
i9bGAbpgbJsuM+G47KpoJOdjkwR/q1ik1ej20TB/E8TGMffBCrXAgvB0F3FgBbIR
aWHcpqaR9Vc/6Hs4ROJ8kBNpXtvjgyJlr6qgpJpVT1mxVOlccSkDo5R817NeA+La
xh05FQ31hOCCOviqwC2I9K88btb01qlfnQ0N+kXpotoUOsFR2F4D57CvqthWWjOw
XkFKLTOHxub75MCDawXzo8gt6KMX9dQqrUw4Hq83hBiJmifRvhQfN0OAjLrlLp+0
r/hJRJvE2ejYxKeaaE9F+0vIbo6iH8zpEjHGR3072oXYFku3F29nQ6Cw73qmDn46
+E+ICXHq/7YjWA4NK14Zz7DQrQq9NfS4ggf9Zwl2kH+cjWbL4xbnaHTQelIRkLOG
kt9rVmHH0rxRu/I9aKCpbg+BOQisWfdgIvLcSr0Kt+WimRjGuevp7igKAiZSeVUq
VVGB6HKew7ab6YKCvxJLkyE7bRUF04viPo2p/KVfE9rRX+Aao65vN6LFDXGzLVXy
K/Fy9gnHthZUMFWXOAQm4RVNwav7V+HXqgVf/qgwlFUP82YjuycEekiYi1yeiP2f
5o/t83E/LvP8VmjnpuNCEW+CQ0hBOxWyUFwQse1bbcFtmiGY6i5FkeWJJhGmpxgS
RXXudRme+0kahCZX3sDQ/+x3RdTYMSYl8pQMDjcDjL0ZvmrIouPqahkh/BbbTyx3
PRduy2Mdb3elmsGjp4tmyz94AM9SnstSqv7E3S+gmUc9g9OKM5Wnh5GFj7/ddKUb
rblthhxrWxxD1IYeRJcZTp0ZgvsofbMNMrWF9pRu6hdPbs9wCQn2FV2Pm7TJp668
D4j9pzEr6eSIlRF/AOrTSy34FLBf+O5z8a+crkFPNmnow/omrcmwmq+PA266ATva
U909Jf6KkTukTCWCSxaURFu8IKg69pcLk2NDRnhFUSIxASEDfrRLLvawjMlgsdX0
qarDB3v7SkzqtZ1S81h2hvo4yKcW8vANASz2ahPkpgB6mMvZrrWkZeyLntIzueFJ
ZvsNtbfJQeJhLLVkOwLJTrS5roHNMTJVRrJrODWZeggos4KZVeLCyWJVfZ66WnYO
sMGIGwEI/6Hj90H5eWCrZrRXym4ZV/xfWruPWLHNd0MQxX8FBU+xXEh3KEGAiSy8
ZGKwBKD4pZSciC11pDB+RkpepE4eKB73UuyNmHVbcU80wyMzA0WOlAfvTJibXy+w
nbsLPdaWm8vLaY8zfdMZsorg7Iuv2Y4v96/XmLAah6otfXEf9m3C8fIOMZkioAz2
7uNwMrJmnzeTRMt1LlZIauYcyL1m+qbhhOs7X86Meqew8OZZSa4PWCw3DWiAURqS
YReSPKbElv+DmMluoQfgBmjPLaaQMkmb4Y/je9aDEUX63ETP93gHCOBPwoQt4hYe
w+WZXNaYvfrtAgzXM8xOarG6P+QB6/J+umQihA9MsPYmuPWLXt78RSy4c3iNnGmn
Ar3cZZVWdm28fqXCyXhQi9ZeKhms0wK6IsVNTH3lwa53c6G9tDD1nfSmiFHqDYJk
QXSUVE9w9N1WYPeQ8blRTMESJtugskaS2UDFHxMT4uMyKQBZ+/bqTwxTHpAMFo84
kqJtFLeOeZU7uGXBWS3u+NcYPYnUnDNa73VQ8rM8zWQ8p62PmLDSHRB/N4WitgNr
5Rb9eGTyesh2ySHlyNoyluNygJKNl3A44p1ZwM0uPbxZ4IoQtCeIBP5/VhBW7xvw
ecxpFdUGEY7z94dHmFpZnrzPCKVdmMQ7vBswjBFMqjnDS6NDVp1Hpcmzq3QzrqVR
wCjt/DdYcMQpwk1slkVUCrs6jSr4CjZmG1UZdP8ptoXzW6gPffiLurEbXYbwrWqH
cyZ8+0ysdFGEbGSrDUaU+PVuBP45QlncFoCdkyyzheIhtUAWHKspS363WBEqUTGs
qsxXotm4VvGw9eq+INClQ9iTKfvgZIHbJduHFBmwPckYJKlIZvH2R5gdwCdjKh7U
ZqrHSlxLmjPXqM/4wjpt3H99CRSzQ7ii00jZRlDIJ/D6vOrrS+W1yWe77zfZs9Uv
TM1rh0lJFMgepM2otUWqlRwl/UzwF76K5xas3VaUcuuMYZdn7zPVfo5V8KAuMB2Q
sPZnpVIAramMgrnrLOSU+YMusPXLZGa5LHA8T/9NZ7wpw4zUPU755xCQawe19UtA
vtW2dqvKE5wnsSCZY9FC1tXRZD4iRsesFzH2Jbsx9pKGluy6yRukq4I/lTbPixVb
FuzFoWn2Xw47sQnFw6n9SM0Y1uI1OGlNRvW+E1pU52+TlcTZIm+WqWKSJMgrwBGy
ocyphgXGAkv39pT9eaAK63CeosTB1UKBRhONuh16lM4I3X1cA6YvleeGgooCil6N
99qnYy66txj4t/DPT0iIdg4DDDUD+T6FwqsGtWx7ADZrdtNGGTnKOSUjZa7touDd
jxo0rTPdzHnqNLB3/X0XIHkLVWiLxMIb4rd2oH359muVOC3tag59fQ2UiGBEBsZp
o5G7ar48FVwLan6pmi7ewtCWseasLWAgMfCCSy8mK2ITdLDuMtgcRGGfJGqT4Zjy
Uq8pOD3qoJJMSyQPvgqz0q1q5jFNc1BJVO/XxPlF5kxbvnIZn9ceoFFKU4UZ/c8S
DCPtGpkxYi2/EZzNa7ErjiUVbmIxNp1FlXUNJLLmPIG+U6YIvtenfROcvxEoHcSV
ALb47AUKoP41IyGXloDq3C71uSKS4Y6tvVXIJY5a8XxRg8QNXhJrQw4nBbkK5KLd
GjRhg1YYvmtkw0ep2B1qIEyf4BfVfstLaz2/UjrKK8vFvVHe4ZnSWl+1oKMvLjAt
sqiiUzqfIRpCFfIMU7b/WBhs0hu3n2g3CjDGW8v3GF3342YoNgsLW7kcMNpdJBqG
AdoPPc1HrBgLH3SPC5BaCYW27hGutXMWCyu18uvwHSxl+NS+d/hjn955jQrpKlGJ
Sb8N2Sm+wsacDczPU+N4aP9yIYHAzFmH4NCYruIShUF6heSjo/cc4e2PNfYn+rjC
xJU7sS2tiy9mcDFt7h2jFs7gCjZ40EdPzKA5x7/hicb4FQZ4Rf7hiPpNATb/vB4X
qpWw8E2Rqg322pmFYzxYKu1iV75ath5WtIrIXqkuUm2P9qCVDbOOg4mwQIC5S6n7
sPt3fy33FYtdqgLGctUON2G5j5MY2v+q6aynwpziT2Ck6OlY1FWRx/AU6yFDSusa
xBOdwCsqgwuYmGthkDB91G5GO7p7r7dSRdRkdXfZ27hNy+Sbj2eddQPUILpdAKDq
m7lt1xQJpEOAtuM6XUAEx6ECMzo/2E4cZ7g6JiqKddGAZjADcYkpfsMW+Pc5C3yW
PyYZMrDXm/xXNR8YPLrdSqqR41hhwwgyO5NsHfnnPdiKgtDgmIuARgUbJiMT1QYb
1zT9yz+YOUHqU/+amDqiS7jTib8KeF39e8yl/vJaBsPYX+gcXGGhAtnd/oAN7n5N
GCSvnbVhX1+O6sHn7omkqWUot9XBbeWzoZFOpH2dfvAjoYG3Ela9EHN2lbE8F6tF
ABLP66AkMz9SkLhPCgik5cko92/VdCVAcQmci0/MHIuCuptvL+/3lzznGiMb2xwX
WHO973KEoOI8wSS05oQIHdt7U5zg+vWMCMhtIBg/FbrHnXqA3H1v8vqBLdpaLMon
bil5QGtdBRumcn7DpLbYszdCQ9VxFh/mK8EGkUsDDZ1v/tniTlxg8xh5jaSJYdOV
rT/BHi48L+aatTBv/PLyumQhtBE6QMg1s0WNZ3EKZ4NX1nlMp7FSTQpUygtfFeH2
ubiYwTE0KyR65x9E7Pfef42l1rk4ZZooPBZOB8eh1NgglkYZLozMifIS4TT96p/G
i/9m64S3hl7dFBgRyp4UuZe/fo0UFMMOA8V5q9R/fPIK6RZOAvebArOdPrCRq8jj
r2ygPeehIXJZpBrUy3rhA/Fb7dI6mcHT1tM4cW5/HwMnNniZ1VCnjf/iZZ0LEm3t
nzrCkYwjJaYfDEOhvMrz2BDcV7PGX8CSuu4yzf00auu1qWbNkuUPRRk5CEB2FW7s
5/LAByDnQOHG/4hvgwl7eipKy8Ab8AJc1uQrwpFxcyxPDSCLhmtnjKXx7Yz5TesF
oBS8YAnf0PuITRdtfaEr7VvUCoALSb0m48Tr8s9EorSqT4itKt26rc8QaLvaM5Gy
zrxqMYMa4ZMr+Ag8UTneMwowaUUuZi3MdhQQgisVUiMGTQNarGEcmUWLtR4hEWAr
HY0R16v8wQRRdOU59S+qQEquUp/i734c5V3vQV2uD9ngByUyO3WHPQN7UOw/8xI/
+Ri91czzy41lYQ9U29Z75ZpCfnSXDwoml9BUy6EP3B47KYps5ImE0lZ09mKVVVcY
je8qyogzPNePu5YLldcuQQgMyOhpA7GGxTdhyqR00thjnlBB9T4becoOuh0eWBlq
NjbpdCMayu+NyEvtHH2hWCvNRuXdveRreowRYCDBVo07hZli6bUIOqKc15NrDoLl
B0Ki850Mb8uxlW7wbtAZLDQOwbW/IMrqfny+haFxHf5kMP/iNnJURuE7Ww0OE4U3
iHKqAr9XxtBb+XbeYY6BlOE5a9WnGeP9HnHz3k4xb+QYAapi3+X0kQy7g7k5XAbg
L6fFeJ7/QGkIhIBYIrbffrN+TqmhavnsLSn2xgbPqfUdW7uPxLBwDspZ5/CV0wVg
DujLn/GSmnnRuJDChOb+Z+DPhmJTybrspzKH6bovLsM+KvJp6S4V3DywYonC3P+o
8fInvkIKNI4wZiQ8If0GF/JpkM1b4s0fA0XOgHbXjCq7iDnr2RaqYstbQjFJgnwV
KlUbi1MzdhgXKVZTDiPZYytNMrnuTXHUjgYcIbwYWbDKT5kuoK4LTAP3JMBrFDMQ
NGjeXwYAPzR7RYBq2Q0OTmsTa9XGh0mr5Tmi74QMoEpgB4DJsXPWx5xoCXJUb6So
kTNSOpxgYuejuX1mobilTCjYyYwkfMaYfMVgJUchnT1wSwShI4B5lhKJho36Co0L
G5cJCnNsTWiR6X7ApyuQEIqNfuwZHtVouzX9FmjoKDKkL++0nDCEw/UU3AqvYKYr
pAHHDNHAyejU8n+fVxktKC1VgZaA2h46lF7J1s18hLEmFqffllSxnt8sHHuMa8mc
2jYhQChdfv2YMPqTfjKWFqw+HPutRnjBqR7xejH0MGs+vGuKcSy7SnUyO0c1RsMV
07fafLtWZtKxBR3YczNX8kVeC3qdWUPHEH+ObF9iGKpKqpllP7NB2HaIqsSm/OhR
dagHVcNy+sFObwzdFIbswOoX9blLr0rNVUhHLAtk2Q/R7qsS7V6Smbe0cK0Pa41c
2wVjJlXQVflLNe5uvbvdAFxgRiCLmCdco4AmBtCeCbe40vIrZZw4qHVlsGwPzuOI
3P5cLNaPohisJ1NH263FUj1TXIxge70vKcPyomD7SJ15xmB7EVuHK+xW+zG2G7zc
Od1JrMvgXpIxK/SmFFDJ7xUOEzIrtzYP9RteP7A6ZV0X2XZfAmomyoUAtnKZWnu3
FDzLP95o8yi3Xcw1tZDdRqHjSocydbFdadWCJCoD3CDNVVt8iFxPY9N9mcpjevXz
zpTtnW+L2xRjV5inAXMVF3T4ThstR00pm5MTwWRbOneE+4AN7A5m7FgsCIVYyMhF
OCug7eEGk+9RRW7xsHWDWm/XmZVjceX22Y0d1fuoKKGJsRat1iVygtECxUjWN3YY
0KnXqtSNA5Ns8e0c2pR0x+hw1KIkLkmg56L98jSfxrwPfE24ziVrwUxzmY2/UI59
UiBfYLWLdEPJGHnhoHVaqLJo6VJV3QVr0G2eqofea8X1Pv0FzcO3GFJh2ESrZ46E
oy2BrrZRTIo0Aij5FJHg21iB9D8l95GB9Ne/j7jeE/j8gU4w7zIqBP3P6SZZ0K76
eoGjE/9uJFHyVoKmH93Zc76lRedV1JhISkks63YY4EW08RusvjO4rvJocsPVNMI0
IjgkRszpNV6BD/N8Hlyz35hxBBeCKjgJ5zkRMA5JP34RuTW3MWCngEkM/qsayzJE
0gMl+iv97GocE0azraTmpdkveTpxtLJMi2iSoMyGRy9ndbcldgE/6pWTd/p1gmRw
pCAZox0zgcCVNeyhv+9tAwfcxWV9nLOoSWVhYYN383unzxmyxhGqsbZ6D8FxIPCP
wYSar4lEq0Jrot6aKi4OjvMZqeD3Vv+QefOQ8dsuxniyiDoJkFxqCWguUruKTOBj
aH5xgIlZtHQEiBwqYG6lj7ZkgN9DWBhkusQ6+3P7iIKmbLvadhoBhdLF1OEHWDif
PHEnfi6z/tiqJoBf+I1T/dYLeNUEgaAT9TZbnZ0SgFZNhxbcafTBB18CVID7lrvz
7VZiAeJNXGhoNicvVUTD/v/pxvROE5ad4ARZfwAByh8EjSegeQN2lxJ6i0Hc9hFQ
c785pXd/QJp3/cBWtxWWIZ6DlAVZfcksPQRX4G//EWhsfqKpbBAJc37rWtub8ayZ
WqZf8r9hAH+If5wpr/s3asgdoE+m03BitzTQuCmUlpxBRTpd4yoGleaCGr+j2gZS
rFFjawx1oclTpqVwecqSYANh2wAUUum/NqrUSGerXTrCwpjX+90VQQBkozJG1S/g
4BNOrCLIJeahH+/bhZ+cuphba7xiTmSVsYMEKbhI7XQqx8Ep9xmJSgSpoUJJsprh
0hQGhLbDMd8zSV+LvP04PpzK22H2ElSlthkVQqpcdOw79Qe+G5KIDSCTC0/zpJwP
3ivYdlKeaGEM8DPhN0wCwzaHvuFIlMGBb6DJxujQoAemkxyWvlXPtHgWSP7MaYyV
Pj7QoQDgYNzKu7ymbJIa5PmibkpWhUuo9WOv8+sMbZFeUg4SMn9vhcjWAVnponRo
kcvppbX90T4Xn1BAqthJsatjG7CqF5REEjFIc4TzjwbHkYOoyyIhCEob2ez1/rW3
YnlFJVeCkv7Nmz/Xi7sqHUBjExbIa0KAHVZNfphK4Cxmrm6kOINtTPp9ar99YVhy
iiZvOmLEBr7sriIHLfnGfJEj9DrfPNhFQcr1htpOeuyO6dvzER1XNJDtVXrByiJ5
B5sQoE2Ns5D/LAzo30XuIsaEbw7pc3glOYBnw+cvmhOauQkm5qCb0Y5nppCaUE3n
Vwx8PBWXNEZFRWTbJnsFpE5wV6grjUxYhGAHviRhO4o3Sg6cjTb4Pc1TQKuOYEye
ouHUKbVFoytYP198l0d36dmF9SVKSjFeVy1cd6Pw6gglU0ut0DZv4l21Fk43nVBW
blDMIbqpzTH8jwo/aWG41R3d2GbsbJutIVEZaP16qztmpXusea8YNneD3szd2nec
e54Ayl6tkqVuYdTkBcpuIzw1RVwdMbSC+n9N4If3UDa6/nOVuWykLc3lLMoxmBd3
w2WuEvye6vSl21E/RmCDpy3onnZ/0+OWC8FyzbQ0AmpRd4LtnEVhA0ciXgjYD4Wy
a/odcozzwLZ1ueir0sIK7lhk7Hjet2eC3vpCLjhfuUYOo5Sf7cjxisZMh9nmpDdd
aRPAvP89zOLkfULUetsXo/VXXohckBKm0l8AjMm/VeACxEtZPVbeUm9yZZikSomT
z8lJwWb/SrtNsnyiCwfTaA6pLy2+Ppe5ROdFThHoq4Y9CMkmJMMVyF5CqS5HUWFk
OIMRLdT7YLiWkAC78SzdHNHhxQ/CaPiChVT1Xxi2TRufxQ/ky/+WCOVhcbWipwle
V4RJL3Z623KWDnhyJs2TWb2TuBYjsjmj+xOWZwUGMe6vRCPbF8pbeUHiQhm65zjN
UeZzmBks7ZNN+RxZ1MTg8CwfqMHsujbMKPVSqU7+oMwmbiagfLxWkqf9zVIHhasd
i+L56+HZzUKDTFW9fTfhiWG9YjR1v1HdZStYRJOYo2o54q3V1mH3nvOmjUg20a2L
USUK5riSuUcr1qteQySai7RYG1/VZTLgSGUjznymABB8dfGyJYSTisaBs16lQy1J
a6m2oNV9PkjOFvRh2xU8tuJcHotyn7i8W+WHRw2YYq8n4PCW4M7Az06diy6fJWu2
diH8rVoHWRje75xga6AavOJIivaOKKh9tjEae49wbdy+OaVvdtNKbm4ty6iKcZ+g
8PMr75+TIhcCncWE/J6IN60zeJE3FHcEJriW9QMYVsm1jkWj4rZi2Z+xLzIeIcx6
b2efIdV8e5ArzmPEhLAyJ2i0OR0o1RQ6oRmWTPRGutku/imZfndeHT85qiO7CdVX
lfxT92e9gZO4s9iR9GSoCaoYu+HqitQP+X6X3PPYnl3TE2gXyraqIbBoHs1qD9Go
2qGexLmVPsjBolLH7V4JfmTFLGnAzBQftwVI5Qi8/jIxmnM1EyxGZWvea9WGc3tp
cxsA5HjXIO1jCztYhe2CB9MNBy1tdjpP9zqLBYWJQ6rfX1qneL136H1C1F6nHIqQ
Xo++WFwF8cNE7ps2an/vdsE0HyG38wlfftd+iiFFtVU0oJLhv3b6GnLx5lP+vri1
ZXDrbZXrHg1RIrdOdCf4lQEcSLLnID8lxf8/yuqnbhRtcwlF5e5TyTQL7mnQwzKU
MMshgdOOncl1nCmcpM44blDcs8NTuDrr6ViSnLtiJ5n9aWKlmb952UkWM7AK9J1i
JBA/iBYP3+U/ZFvvvDSq20xhPj00Vl8eWVjtHOdA0f5CovYuZcE+8GTTYIwOHSc6
al68UjU3GD7J3QpD1JE6wbyfIBTn5ANP0junEslP+E3igeTIsBB1LGZ5tccfgyW2
hE7acJiElQ+1lGtR7W9lyyx8fy6uM6SpRK2sFattqikbc4/du3AnWoFJCXWIkm4q
qINwqqBtnCTec3ruQRNphxMAIb397ikNW/7MnYB2/78DzzuTtjLDZkIzofhtMM2Z
uEUknIv+q5IPMiikUgujIyouKIVRx/P6LCiRF7mkPOtx3CuZUH0bStSXvO1d4HLa
4liIYWO0ZDpZ6cvtY1yjFKuAqnaeRVg6JLxxu6sa352kR5LsMsUxV3zZpJIIKRuK
IN3hwYY2fDchL8tpRH9mLCSHOueRCGLE1rhzm3l7/VX67624teqi1JsWEBgJiA9k
/tW13fmOD4U1ZqA/KrrllKhjxXQCXp8AnqXjUUJOXfaMe4UYtfiVKtXHJlOoGYZj
ksVW7v1pV3iNRr5+eHmYH4uxj9CnQIbNJ7OfEHJvjBJj6z4PSk7TTWdyEbJnZ6Rx
mcaI5/aje1ZewyGXbn57eb7LB3tKRk/OdkCUgBVhhQW773LCMzAVWdtdrj7XHgdK
IWD7SaolWY1FPvAUFA/goVKcVOOwRnxptZmqhUQ9KweSCjV64jm83RRUivvwzGZv
HT35bOF40v0x/D0EwHiTOajUyuyfXNV990n6LOr1YW6AnbWxcIgPh8mAuKbNz3xx
DFDOLTVdPNtItm3lDhCh5CV+vQm8V1Qn91C1E5YmIa7gjcjyDi0aqCt4qPXh/PII
QcQfEUYA9JCMpCa7mT5ahADZLZ+J1RNCvjmE/i9SYaFER9G7KeWBF4Gsj7avHh0Z
C1agOpw759ilHt94iKLaGmUKO3sdm5y6aUnGy4eAKCeb3OA2mzpCAEiMGIeqX3pl
LKq8BL5R0/0UWwvBC3kexOnUSDFbygvPB+ApKWMjMCWxJxESJEmKzZ6xMaeTsBhh
he18LbkHbgyDBkfKHKmZfaOqGvnB8oBdWf1O7arb5OA74uNxOvecTf1E1RDHPlJp
gMq+2rt4iGLZAeeFtjFlReuhQ6dhnf9q+fWeGWB9m+D77o2D4ctwvvx8q+2CoXrd
JHsuRl20rEU9J1eHKki+o9pv/tii/MzemQAVE/wIZkmk1KwClaMq/Ij7smyKlSiM
c8v1dCrA6aflKF5xJfRKG+VP2hv7X4mTsLpgZVPsJ9F5Pipd6FrN/oBkLzlvzdk4
Zijncn2hvo3Ce+F6EVSdnXCrR95MJIbnD5Z5Admzx5B/JZ6/N9FoqjmXIntCBOul
fbQxW5h0B4thAyQH8IeFTB0BGK+QEEAAVoXY66bE8eAE3g2hRC+8eKRqjZ+Q75Qk
j6LXcgupS3wMdMxHvBFq6G8oTsKnmo3S64TR3gVE5wYIsS+CAfEyro3XxoukfEFu
Q0GGNNSSPCt1z2K1SMVjaZAQcQMryZWLwc5z84JVfi4v6qNiV25UAbCy9D4bDwWQ
iVlgabEVIdY//XNrK37R+2y61MGkloenibcKiomnuNE2Vorf4GrmZWzXkRjZIr5V
93g63iKhrODtelYwMpLV0NhUiI+T5z7pvtUxM4cMfuSYfJYemLfKOgIREEd26K91
n3zzkQKkIyCn6q8j31aHw80K7qiw5FsUS3oI1DbKBkN6NzagOA5ydSYK1ONvdju0
cNtEyWpSAeFuR70B/K/iO3byltV8gm9DXeMZlUJg7gdtPz0c9YtHWbKJXL+Nv7Iu
XMVVHm7aJvwdwYpanh16IU80mPYCORkb17ErJsxRDkVaU3xauJeML1pjgSyrenZ1
ftiSwK+WGybESu5v1Ep9STUefeMrtYNoFhZ9CNQuOvNp8C4Ja1SyuyK2VDUKX5ed
w7TZ8PavlC70WN6EoOWfwf70SAjZX1/RwMzeYml4AsCiZhcBd2lWBZE2Nmut8kg+
qTBTK0QQp/B1iZOZ9cZtU2dkEI7BAZfxqCHPdpBUITixCSwHof5juccX8MRRwYmh
8iBhOidv0bU4uVAN/9/ez253wGUQz3AZQUKox/h+KwOL5nPSi9dIionmos3QUZi3
Ng8aA95yBmC4pT9WVVmrCuHJS+ovyMKNPmOHqw2IBV2+eOlsi3sDV5f0THPRWF8V
hYeKFNATyqXTERrxKE17H+zh/Ou145ARe7+5jOWW2V/X2al6wzCLu/ly8n+9R0yX
JIuAl53PHHIBytTZisA/YeQU9vq9kzZkfCQPMRxpOwJujaWH9E/k2NsYxiMEPFTJ
MoUSih+lV83fUUEKYf3VfVVeUVLbeKNP+nKNqYgMad6blvonJonwpXUi8hiDgVPe
etuF7W/UtvYRxGMHIXE7kREi7mglp9nREYAOEEd+Er3UghB7y/Vi4pNr8LY/xPOJ
xbKXbhtKpkRD1rSgdc2ixsxdXqN2HTjxLiALdHyhyvwKnxOpkPOCHWB54o9/33NS
EFJ66hxlqcHRzouckk5LTQiubrf7a2aiGaQLJ1Ln8mr8E6o2hkTbx/DqlJKQwTvO
seXxPul2hnuOf3ilJMw84aTLQgRNdmiXskbez9rREbZKutqHltQBL2fE9NvUDZB4
/TCQBtyC8izfOspuRwh5i7q/0WIGw6LQKyGUDIS2BY/9UgueVClOqCN3GWqG/kwn
fc0L/uRiAfNGp0R7Aj8NUUzbhTRkwnioP9jFRtbjfzMTr8nQ6wIbUIwCykY/YDwh
m3kozofH9wsnUgYpph6Vm4FGdQSO96mR0PP4iORqUywbIa+cxtmeb38XgJpdlxBs
GbVIvV3ga1xFRCGivrW0o7I4QQx3uJAF2z1vP9Nl3xugOycIIF0B1FFd9Gx0TfuL
aVQksyU+650j/GjdhJNpYGgXOfGyBhHFGSaXsOJbvqzAtTSjSFR2zYpFRAOLcOZX
EAlMUtCpluM51bnpnTYxuIaOp3x7RNutnVDPVGKeIsoo8abXFnXYYyYunIxlk2Fp
WI0ccxLwek5pWJSSJ8PnEfrJ6YaROTBdGXzA2+bZxMFx9CeGJwpVIi1mI3cCp5dm
0uf0qcsXpheK+t1I1g6EJV5YJ/t3NaXAzEmt9fXVmfJxctEteaxRWMoZY0FfqMBc
EAdZ/nuMiF64MqY+OrZzHsiMRzh6p/Fc/26zZcT3RRvcdru46NxvUsXNDm2xcyd5
C4/HnJZmXL0dZVN5BieqejhAg+7R7xfrwJsKed2tYYlFUafKFH/tkwSCbgqpSshW
S7CByhpvSK24jlUpvFGlg2Qb9IeCnpYlggb7EvylvpwEZ6uKPBQIAOoUcs+vN0GF
ULI2JcLVHvW68LrNHPJ9O2XBljaLSFvwBfWc/LXGum2h2AlW83qCmSGecR+cf8sN
lDQlNsXpvgpWFzQYRGYSWpEyqgwq8gdSIb6grNJ/kp87nVcDyj0ctrefoBmlh6J8
rerYiMSK8eexQf86oIBhtNV3BeEsCTWt/dBeJL2XzCoBC8g8OAMWRdeqYT6S1fvw
4bU4wwgOoRlhXi6NfNFMNIcC1Xkoc6T1hW4cCemSvGH24joj5wQRooA1E3Acgh5H
+bmIb27jH+L9Ick847Zmlz5bpXbWYaxJ4suxaHOlEesPOfSMDE04I/AjbYeCbTAj
mOt101tCSH0OM/3Ucey6uLZ0D+SL3NEtdc2r+IsnxSZt200bK1lcYn2nm9xOtNhj
CLv3v6h3b+KrqzciWXuIlylGJgPsdiwaAyhIh1NW6JK6ql2uor4OvAwB2VShGdUM
7OgeAYaqsYmodd2FWRWCzgL8YgIEJumfk54FvFBHHyK9S2JRH3S8ARN5xkWUAWMZ
+1neQ+2D4tsDnzi8uptg3QcbkN+K33j5AgQEsKgIlBo1xVQ3FP054lgquPoU032k
JZQ0TjHr8FjBHUAL9t7YLIbkzoVU+0hHBx0bDCZnCH4O33qv2l2D1WYU+0h4Xmmb
AIpdR/7U5SEXC29YibV6xekSY+xLPCuTzadhnxRCB5yC2OcKnB8Gpen5yr2hMfkK
jnrhXPS3dprdIycIGm5FztsSsgHX0SHibxJN+suAqkKbqJvYiEUFu9GcvtVWj+Ug
cnCdHprIJm4L6bJTZ685uyDN+KcFpgv8ibnMbvkDL5RqaxEo6Ioa0Ionx2pLC6WM
PSk5LzeKHDMVKHfGoETy2MX2xK4QbPVNkZHhJERRWkeR8WuCFDZGJ2OrjBR5Nxwl
XFuLx5bnmKctjTcgjvp6+/ITddoKrJYe/sH0VlMxhYHkVzUoWJlo0HW8In1OjybY
xev00fa2I9PpPPNrXpb68vS1gPLwPrOkzpK/mmcdo+rV1oJ1lBxOS6uzczwr1DNS
84hJer+jY9LIo6gOKfNWT9SvwvvC4RhhCLExhqe/cWUbB53R9BjIZQvgEY81h3gZ
CHTH6RkWGWouGExHbDMwUpV1prGQc8s+dj4tkzGuye4CVqPrmOpsWpif3zxPkesC
btiwlE1Olji4i96xpIkAxjXl9y09NdCnDDJ49CiHVZ7QxyuHYqd14oE6lPnn1+j1
GPCYBiBQpCifdKEa4wF3XXWm6iIb0m6l3K1NRmzMDNhaoawhpMPHdXno2AEGDLLh
lGpRx0OdKMLPV0p7kBqLCM+Av3OXI9apGbcbhcd3g056miIcrCiMjdiEGMwu0Nrh
Jx4Ekp2WDsUsNERfIJP7o4akADYagzJtG2mCGkdRSrUJtg6nKacdnO/Mlbgy9cce
bxY+z3W9x3GQgBX4y3jyG1WUwI4W2iMoqkit6+k5UIB6yNLkl9yqKLnWmvgiRbYI
2zTdJPlnjAFjb0a5axE1nUbFVAg3SXQb/fqHhKXsYZco4lgQkCHafo9RPQ7lH/BC
6xgPBQhQ6wUFLOTTIBqMLVub2Y4HJjHPv3cdSxZnE+UzObFEoeV90AbOCx8x31Oi
cylAiB4GaMwW++AFpk0GtioIs7KTIYF4C1s5vFygxBdqCXXQ8XCRw6BgkrfHn5ma
yuk0TqYSyGTLrjxE/M6FIlEcKmjlOaw2OHnrmpmzNle6XN4BdAowQgx8hzr3McLl
am1rK4GjhuCRwiy6OM6O3W7b88049xJxpYa9RisIjQ8OVrk66p4Y6q7a3zNZ/CTw
5/JGd0x4XfjSksJ3utZdr5Z50EDr9ODevy9ST6TZ+KUwgp9WXFi/xt3gitG3Al8w
zAgZhmaDc4K/1CS2V4FxLTce3wvPxCFZUubkzM/fHZTTsOdOGmqQO92D51XTEVoo
Yn25AZ85eiXx3NmTmeceUWMPemZlL/NUYdp2+9/Tt3eTcsdvOKGRA29g1hZknh5A
khQAMR5BUpylY4Zqqk3ew3ADcpGp0wStckUDvVtdcPcwJhLFU+5Lj3ghHIXi9gnG
FSCZm6k8ZYh9KOqxOZteXulPCtCFuYMjjyeVLcCfmkXpM8UK8CUdFnY6TykBCd67
XAnPkxnDfZJEXFguVMjRizlpP2mHxs32hbcHvvSbrxaSC44shGN7cVLbCDt5ZqOA
x8ot4Ar3PG7X0dLtWmmFojwC4NKpwv7Fwm+aIVnnKaxjOS8pbax8TcR+ZV1aPDAJ
ENAGBPor5aVc0XD+991GEwpRamnGuvD2FzW6Wo+Q7atCDwfWB0/nksDFpr5sliJX
FUKAEErP6XZvsb9kmBNNELDejIShQYi62bhdA9dovPHX1i5pmItqY1ywFArdbqtV
qblI4CyODmuS/arDRtt2PCPWVpTX1J/az6S0bkuHIR2BiGzg4R3gVbKRcJcVXyeL
1OGSULFhe871KVReSYhRqo668PP4XF9lqYE+hYkm3tH0ISgZCjI79IBUyAGGdx93
jK4ws4xKwk5YogjTSbSh9yPwO1s8kHUnwNBALdLEFksJuZXQaGfZlXFO1Ju+51G8
qoG3BiH+gsR9yLL+BtuLElgloFdK+XqbntdHg/bWMCL89YV1IupuPMS9SoCOuHV9
2cVVgfNhP+c4C3/roaH9As9jbN/HdwsoClsjMB02OmFh/Zulzi78qCwO8NGLh/1U
dvTbldDY8A+ElR16LpKfiiM7+Fo++Fl8i4DW82DYrEGmU52y6k7c/zL3BDLoFpFc
C/ckRaMMEKWN8n8jTZezGX8GiWWQGbkuo/dYjqrbjME5gV/i524XSF1ntnVkTnR2
GsmCqFjguj4eHhzlYETF5I95S1/+biwSsyjSXEFe1dyt9tRY9N9QwebfgmoIwoYO
Dh52cN0tadv1DE/Wx8zJfXECyxDkHui4z1rqGMdg5Mgn5cVe7MG8Jg6MO3EuD1rs
wCfKW4WZ8JFYXGTzBIRSA7T/PB1W4pGzovpVSQTJ65zvqRCHRx57wj5ZwS1wlLno
8XTZkP3Ek+L3c7vhwGORyYnd9ptnb2l4PrLXfMAtVdDRfE0E79KU36a7IuPkdNdk
ike1N/M2svydcJrjs5R3KKBph/9T7XnPKYkBU+KlsCRd0unBCr/NBbyO71SgB9Zo
HstyfXOvj8ItB4ULDy59uyGDfe9UrYr4TDCFZ1DYvTcxtZmWyJlaD631W709j2s4
HB9LRC32OrOudgTUi0nh5PrOKbbfPjEMc2rD5+kKAN3GeAIGPvmaJA7X1euMhTqE
i5sLrv58+uy/pmjn2oZKwea8xogB82cZwJ40/6ULQidG18YlxuqZynm2fkKyuQNc
B4hk65/WjBZOcv7jioYPDUaIipzOPEa1aUwutUEvDxDDCx0ccuphfLu/DdxZQqeA
1Y/fIDcx5kIiFwS6NGydv39LCYq63r+TSFOBOhEc63mSNpdJ2u4VvVON+WsCgsNg
dkC/7fIVh6GhkDaDZNtWL3uavNVfOM6Qgr18xYrgV8BsvaQRXfbIHw/YRQREPCbM
0b9FOX6JuPYPUPdPsakXCImtxI6DxNvivLAoDsyC6fnRtD1aU3kWxXSFNcbeTyQl
qpMrsLja1kAbh5HOd4Kb4kqQl10s9+aiO74Uk5ou/wZF3Y38A4g5CEsBXmc3bWZS
fcd8mwS6R5u5WF/j4DcimL+NwxwTy789gI5G5vgxH6/j0ezhfAahl4cB+p5RzQQb
gNdTbtThFjmxieAZpvcf/sWh+RNRp9eyJTrkHrXTKfJ3P0p2W8LeUocz4S+107eG
840chdifXs8yoW0AuR0dD72xHNTZ0ptKZ+ZClygyV1e5v9b5HJZhx192fPn3dx4S
oHhZvBwAiiC0NdQ2Xmk1MH/N/Cusi9CJY9E1HzXrfunPrOPPN1cAbYAZKjSloUib
1AKZtYm7QWooT1HnV68mwJ3kRgKvVK0V7v7JTvNkIiO71mAA9Oi1ZoyDhKd+2iP+
kr4joVoprQC8iUaAU47cvuhlHf7ML6buljtUXKk3N+Bae7vVhWiN6LQixuzycM1d
3EBwhQh7VVThVYJ4CgDF3zqF5kaTkA3yxGQXVGnEIhEwVC0z9j7CYZFKqjzieLUH
DwZtNpRWylP97uF8Mi1L3ePd5Z9GeakDc+e1iXEwvYTqvc7+j+XF1ZXMLK13Eueg
x47SldB9vuTcV+f+fLlaGFBL5nRkwqdfhYhV89h9ysLM8LwHJjAX2loM2ZeAp7ct
+hmwr4kvVHDdjIcDM6hii5ppm0C3vKhwY+XyIZklHYDMjj53fJFYWYqefiEToa4I
OaK5m0pwRSJ5oQeEAUR9Z4GgHU3vboAqdzNiwcQkH4K6aL4gb7nrVAQeMQV+BTrP
xfHKRK/C3N1DbtB1f+jJlg+EWyQZn1MZC3itagrkAkjMFNptpA0qgC7G2yTjvR7L
FgVpyTCkW2dqBg47C6ANbPfHdRKe4x4FDoSew22MLnZOl5sD0DwkkW7c4WF/Ktn/
HyEJ/Gsg8OjjrV98r2OVPBf04c//KrCaToJDb/DB7I7b97Y1rCDA5qnqNHACEEuG
jOrly+eCqY7YlseJqJDgzOxOenPEdxTTe5I3DmKU9n4KaDLxFxOeiefhmJFRTk9A
6wX1zKbx2uHwQFZN0R5FBySZGdWLFa8WNLa19jw/R0aPdgTfBeErqhyWs1hj6E3s
J8i6GcNiI6fDHv73F60Rj8Atll83556pd0I8OZli1DVCRBfcZJybfg6gt0KZ+Q2K
0EQIK12gWpOQdz4Sa3rrT00BcRZQHwpqweKcvppx8XYEv1B0Q1dDoun1J7ZF7BrO
AymGvsJO/nBR4gMLYq4APzUHD+qrBfpoVijL7nGK8Hpla3D6lM5zribJmiJ61Vwv
NnFsjsiaOCeY7n98vxBJfzkwpw6rce4M+ZUoYQWk5RJNzHdy/uRNH+hWcR0uGA0F
4FiranyW88DT4brl2BfbdmUMviumpNHgOTZufSqaMyjhQ2hE4Jl61gr+8F8IYJ1O
0E5Hl4uA4PZKM1b8chG3FehMR1ZvIdAoIt0f2v8YPRRF+GjdNRMsqo79dcnKOMHW
d0ZI2YAr7wPVhV9ferrhLE5/xkYmqwdI0DikxQmJVROECWFW+u0C4B55YhvYbZZz
7i3IOz4JuDz1N0HeJ9SR3gVAiYinU6E1hjOgAtZn8j8RJyquxG3ifSwqtKoH11zg
A4se22zWE5QMRzzFWcg0/IryUwOb38/89OguDnhWVnm9tFp96lop3VNpDCcZEgs8
gUtnxlTZzxz+UaX1LQ8lcSth0TMJSZrC/KwHIwtnU9r53+K5IJaOZdQdJYU3xNvi
sNFdYH6oVKX3V1c2fgtuJLmDRN0Zj6dTOzrTHbnSzR8EEerSVTzqcT9C2NjUjXID
sx/R94HIwPLM4NaYpfjY1GKu0RWAtFn7AhnvKUYUVvYHZPjEIWEmpCki+wAeFffm
gpqVwKtV9sx46Oqv8r/HBoMV9T9mkRA9KHgqLmfxySJUMf0s8v1zdfR7o3CWLq62
HmK/tJk6WYTOrHY2oCMaHd5WDG/qXqj0V9HzVdpU3WGr9ueO8SKs1rMhvXK24Yam
GJauHW7eduWLckPHTBGyN+ZDooAxI3Ue2Rf/py2Lb5+W+5a6ABVcrB/E6AK8c5M+
ZLlOSL71yaudkXVCpxyQse/etoRd9aF8oW2tVcRimN8xbhpjnpn15gtDqYEBBlCO
5RlvY/d5+mC/iLxsxMqG3sy7h0A/Vb2SM9Skc/b9tdAoMTq1T1OhHDl4ctx6EPL6
beR6a3hPaos4QgDDWc/tDz+siaQ2kys6C1qKTyi7yDIMkCzahj8DmwknMoroOdhl
58nDLdEI7DxAPY358yeADjU1hM0NZbPaHO1Ct+oGcKO259ct+jYHYcgOK5cGTJRX
d5697pNNFYP2/qun67jBjS5yahy5PEZS9PlRTOxOQnUYTqcdqA9CCiaCN4PFHBGD
v7x6ToUEvPYZdWJBXgpDSFjOiVZ1zpI5UC1romgzdXGLD0qZDF3RUtkDxHpwrbgp
6wPgNDGDtPgOvKTBkHNKOM/gL9Z5IgxFCo2+sKgHOiA6/TlO+LE/6FCiLabNdRA8
TlOgzBU48ivglQn0E54V7zJmIr9MtAns/NXU5ZP7j4FcO/JgjfELmaRBzj3Llbz/
GSbECBw4h/usfe85d9x/SBptVK9ttfZbIs5DIYuAJl9sO8qZc46b8z/fRGIv7CZj
/K6bw+sOGqGfEHB/fEC6BsPppumI30a5Jxg6OuDqJEh/iMSsyO3iF9F2X5XQZ1BU
TqzsIlvOjAUZsQuaTdW8Aw7XcR5Uqo9AdEs3aveg73RbrdPM3vpvc5lK3A7MbtOp
NgSaI1W1W0FJwQcIkTl6xQdOdjFajSuDShsySXnV7UHMWIhLSplSW9EWUlWZcZdI
FxEeV0p22dBYSMOK/0jKUP1I+aLanEzmEJbrPQedpxllqINbwi1v7a1Kt6F+0e7o
u3Tnk1PYfmSE/R2qcc728orhF9Ez7knZw53/n1l64Kugp5WzA/LzbFDNEPlpxUcu
dw4L3aO878u8JX1q8vAQ971IRiskgrK+y5dlMp8MkMR3dpxfh03hr+YA8cpv2cxY
xCa5uGEcA+QVIhvX4cKMKpuAKGPf66B4uSUJp4XTs+6Qes2TyH1j7SV+vLFDX5cl
gxqNJT4uXg4aTvGKL4B4+iQxOrxkC0xfqTBzBIHb4EIII+vbTTSZ2OWFj0Y0UhNA
NjlLDoD9DfLRXMKCmo2yCbuf/lv6f1XepkX9JqO3xOsLTjfMdrREJpaId/xyd3ak
IC+rXkZBlLYcGDUcj2dfk4WUxYmR72BsVGEt8S9h24ZkRvUIl0Riu9nz8BR9qWhS
daa6KddGTUNtQtkDoUtUvQ+lOxAQ447N8lFHLvW5FGOA2x1hkFha7ncV1hDS9++k
P8GFaTDNDKOhvFa5opuUGSGUzDg/prlRhmw8TJr+VwuX44CKN4fO+vGyPwQve+EU
Kd/Ibz3CxGFYQw19tcTUd/h3osSm3QSwH+btsuwq2cfbHOz6t4EyYDyZZzv5nX/B
85ZholX5Rb6Mk2dBxrCrTRD4QD2VYwbaehkLp//lZbqtzeISZw1EEFDvWZQ/DhVk
SeAGjS5s9XuTTEdhd2lHGUaQ3V56oL5fox4HQxNMw0FB/iChtJkaW00ZHbcwlH1K
B7eLOujjRe0XX4EqMqjXPXNnpUbQzBDAU/zWJJitHeHZjycSCMOFfUQK8oDZauje
CnnLrIbmVbEBCUJ02lS0P1g3f8OQri6Lk/y38lIAVYKOEr2hbF/GrXbJ+TjP1VmJ
3pbyQ/lgUXZ4CkRyDkWgX9XooptmKbltcO4YrfXanCLbFtWc9zvJlqn5BbQnxqOR
rrV0Onac6x1rNG+SCKwIi1bmUIY3ZDGX/ahur1tkCn4UtE0u6uMpN2dL1gtkbKSq
tKeI25kISZUOfPS75BNG7/M1svIZ3om5R/cLg84i+j1WunoiDS8aCESle+6zx44j
61g51Putzzk0UWSsjPhU2Rh++X9RRBc08hXm66G8+i9fP9G8hR+m5rvz0hCW5T4P
++WnAD5W8nzfs97aWhGRB+bpNMHsHW3wmbqZM972P3Zszc3zyCtdz+vGGLQD2WaI
p+sJu1tXB+JMwLax5tnWf8G6KMWEolgTTNgKaUn1ScXY2UPm4hKDZauezVIwgCM1
Y8SUzo4eJCCczGW2lSPFqwksHcfvNnm7fXcc7l8pD0oZeEFAHkgn+zuHHW77MD9+
rUsLR+/EKtGcwsslcdpLwMLvl49mBPBt0XlSO8SYKdsktTHMGbDyfmSfZOMDgdbK
lI9s+sytCiTUS3Pb30Q5X1rqGFmT6xHyCQPlrTOIM7HY0btC7NmVEOw2WcGbGXhR
Phlz06Sa2K6IyhxsxkCRuJLO8XXyqMwfVUAd8SyhBXLi7GeeRj+ZV5sxhE/5Kzry
irrDbeOp7m+y/4slKQ0Yt0Zz5zvjk6QgJan2zoTKulFk6g/0qArrJAaDhVMFtcxc
t89pHdPw9c6vhUyZbkJo9yOSKkX0RsTa9eXHUxahkzQK5+33PiCWuiivqA+lYssn
+hdTHZHMbimYwTa/c+KIULOLxYP5yp81D3N9yAm+dLOvqD+s8VvznevvqB6oj50p
OqFcJwQBDaY4AgYxhbfJ4DWQxhuiUI0bOcROeRBL8CmjdCp9EAmLBoOFhACJZYR/
bwgOEsHHjNnjoc+GSluXoWCCGZzodgRWhKkPWNmRPmQTql3pS10LcI35r9H/luw7
OpqfyWkrqY95BIxNCiFrmxhapSIf6WmChX0cMeb+MdFQnE7guxlivGfczamSqbUc
KkWhmdVDjP1pS41Xf6qAI1BrNWMvyWhZgsuG4m33iQIARWYvYGZGkjy1Y2N42GQg
CSuSuhpE6EUHYsWCXj5R2U+am4IkNUR0IQ+4hqcI5PRcNRtKNLObTv66d8OSfqKU
xbGLKyRix7EIz9+ubu5n/Tk9fpu5PA9kfp0SRsQeLM4AfmMp9j1V4tbsNf1P1WRK
L+0msk2fefVsxeF2IlPLKUYsecAzyCVF/yNniy2E2s/IwdDUVIwJHNAOT6g8o3mE
MkLK4yK7L2r3IRCVGOAijOQmGsOqqNbXVqQQ2dxeF06ivXuaUVUuExt8bGvt6cMy
3iODC0U0zDT3yhmPeBOE7NtmAekag9/ygUnCwiFX8KTM+zMFXJLNdsmlqdIapSln
+WlnbjPwMiiRkonL67GF2MTeRFq6rkxvPb/jkbG6Gj+mCjJNePvmQOYGqGyWLpzS
rvVc9TCRHyiHMiShLecjZH3LiFxlzf5Eel1cOrvJ+O0ElARWgw2lTTp6THU/cZcJ
RzT3J/GwWxCURUYA+51oM08McOk0a4w9Lu3hW8X6GtrVwLhGmWfxkiM3q2IFlKV+
jWkDHVJD9P+QzTQnGUR77ED2i5x0c8zceSeWbGnlY/Nqtzz6Ft+6qo6noyBZLkSD
Bf9wxJ9n/gY79WKhTTbHIA6KoPVLdtTdkoqUWZp6XRCSD+TfH6cksgo1Q+FrZ3zX
6moA2XbjeJtSaVa/a80LQPD5NaXjFdld/iP9ZPL6w5S9LQcCtZxSvagZr1sYJm/J
ZEIgXIUUooj9WQ6U0G+FvJQthby/sGxWSxSlmgUJiy2euJbSHeMSgvtAo8XrI1G/
TQguOMA56O9NZ1zJ/hDnRW1SuN5mj40XDJGSM8PNWBJPyMZsja/+tUaYkNzLl8oE
nPjSw7gBbSawTxZitGWprKtPBZOtyOH1rGIYqVO1/Om6CFVJptBqLZot5mXmMztX
S5kbW4HGEjkO+g5qltNiEoMZN76l+15NpZYfCPQHsvY6gWxUyOX7Fzmx6wjMcjV+
GCFUMn+Zf3yOFwyMOl9g8aC/zmztqQc+fP/xdTlDPIWfMFKR1HlmlV/0bKlCCOQ0
VcOp1TFCOMbJfUjsLf7OIrJAgvZCBL26SbFH3/025A1TwDvWa3yGKI9Evvv7SYEt
897Vx3NKqIdpdXtR0VKHF6Up738NRHHnV2PxHudlWyDJ2vN7h8Jh5VJgfDnLQZJC
Hw1ueUWJSV6WT+c24kAcGrUp/CA/+gpsIOAbCdesjVc7KOpd2NIFfWY2mjFYoLO4
TW0lQF0US2kFOYS9fPlbIle++a0i6WN+0ZG8twRU8xz7u7VnwVigM9/oo3HXS4lp
ZY3u+dwOO3Jn3P/MRow00Qk+Bv3+Tme8uUJxQpsoKes9PCOmNSO2Y28rx7/hP0sW
1YlER0cyfV5DpUhGFs9O9LWWODBL+ecKaVrc3T/Us/va14vVdA5QvL2PEOQePJbN
I61BJukr2NJM8uD+ibmW+majLjox7AGHpVgHuejN2cu8TPBWB5uc4/UpHyFrHaTI
zB4exkELcYY+r9lhgCXbF++GIPMGfpSo7C2pOIKepTWNPGa7u+hbJSD22plSZbay
ZWDH+E0HOa6ZdAtD2l2I3wePFkzOV+XU+59ZyfUpsf3b2EbhbeGdeGP5G7S/Jfvr
DA4V1kFWsMxxemLwarIpUlDBcGKr74iP+/PenzI8U/WfQ8NkwI28Coc4cTsV6uv2
tiBsZI1Yrn4fgfzMERwdJbOYGHn8/v+8dJsSVOhURJWyI8E+ESY9ZyxLsz5jrFnc
cgz9CFx2HdKWNAwEzR9xuU04hS7J1OaWWJbvN/RZVd6Ea9sNXYm0G4x6aUhmp/sk
DJNN1lMr2Of/Bf9Y4XNMSsQhjKvm2BXd82eFTRkGAMVS6uCyhWz/Ig5XHjSl+W3F
GK35Jikk5tf4pzkM4rxjgEtDQn/v6wmDm4QyLCNHQDY1V9kuDaMzaX+xXnkAaZJr
Yn/L2XSgsiHebdXuanTD3ZE8CncaFZvuFQzpoHuAYoCmKWEWsfpYclZ77wylvFXx
iEDK2XoIGSHwery06DX8ab7f4j7FNafDVziI/ehdsQsROeFOkPvraB3w+ZpdRsys
ZG8p7zAR3r2afUvD/AEftg+7ZmkEgvJO9VAUI0Ud7viy97+BztXcwprUuk+cCWww
XyOsGe+q05cYPjk7CxovH8GmJ0KHqAG9X3X9O69qo1Um0gu+Qte/tRa6a+xWWXSr
WgZebdavK7Y6DQ2iInKkdaqsRVkl8lIDMPBsgQQHKMrmfjsj6BaWN3rPMVF1crlQ
gfJR2V8s6y7ImBQDXSgL3f8dp+/OeixPgzMd7K2t4wi3BEjPnn5sJiGMdjzVWEyd
UJjZUulH74GjBuMfORUJ0AuGkuO1JDu/KR14QjmoHYgMpDogTmV7RO23FKr9Xc76
UMNae/pZNFTMKfPXrwt3G06kVy9zRWejuaA/XuP5pDuSkBKMERjTBXelwUvBHvdr
1ZIJW8o//ViIJFw+dzMyBiCD10xD8xUjyciz7iw2ssJFW0Mgu+9+m8CpcOSUDhGf
N3o/AaxVGwfdWrxo4srLIlCctrjYH/7iRWRI2BSapHDWYvPnWT9jnRiX0cNnFR6J
Dz5HfwdW5pY2HFJcRDC8gnjCh7KdFOV4hGk68HEUwJ5yg0pxRh53hM9990ILmOOX
BzR/AHNp/0j6KG1Ka4+r85d/OAdKllzLtMcbfhiikGo85CYWu1qBhiMqYMhBSBWh
1qWRWiFgKv1BUkuqx2Re+mD0jS09PPGInhn6meLDQ3E+gQa52sWPJcwnAAIergbr
KDsISiWwMJI8o95uODzPSr+k+YtnCBxllZOb0BQkUo60XrmfSN4Nd3r/JcAT2NeZ
GtmJtC2j9eN+iRxuBcuCvNzyf7g1oDulPo/zo/5cX4kqXyOhuQUxd/HnVqluSlS9
hPj3xKzd3x0VP/lqW3Fkggp1Ht8z3APb9iqKi/XbCb5PkPw2xDKFcNSzDYjnRXkG
BfRksNlhqsVbzXpUdHi0qfCKrEvPrcdhNwUxy3dduLw/nWFeBsa0k8kpJ6Cwt9II
qaQYKwBwsVXH4p6/YnqwQdBh8Bbih4xZnhj6Y9XWxOnxrYvcevllYhauNgZDxs8B
WFfaSBuqYPS3elpvBUxLjc08mENUfF0tjlaGDjoV+riwSoZ3A+jU9tj0QgbUvh5n
FHmlNNdQNe37tjcIarZZPQh1fiiixQYEsyWWHGN/VnMVzCV/iindoLldiPrz2eve
W/EbqeL4seaG2OskG+26ldfTUUmO41mmJPBphqho4K4kjGa+I45otNn9iy7Zjepm
0o2TkHPfId+y3Vofc2NEgsHb4i1p5h4+0/8kim6WMVoC/mL4Siyym0GMncbRkRC/
4KCqmWS+pgFuw7DRTwx2aVo7LhS0QadicbhmR7Mo+TypgIBrzPWSC8oi3TL0Gw7o
RXXsCzPJHX+wWWEdYD+UUC0CW3FVGw88NSme7zqBK56EFBdqni6R327XR7gdGMuI
5c12IRKu77YjAnShmdagH0rDIa5kwLGla29XddxTgqK05UQpZdvmai9J/i+/XjbF
EuCgR6iOK0epda4VjSNqjrM+fXh6JNlAu7xAAMsp26poLXyMVrp4jHeSc6Uaslpv
vRPHX7ROighaTxYkmz3DkRmy/YnVdQOoAyhyZeUjJ1w65pc2BU1etw1qL1G7x9Rg
fO5rgTxPeCcPZAZcRNVn6ZNTNTMeFTVTi7jDZyoFgUHHVPWU2WkV7X8S5lE+sSMA
Gve4z0Ei8erNYwFs1KnPGAIM9F2/nxB7OjL/EFN35rxBpjlHQ5BTXXzboCsqp/nu
V131I0UC7o3opr7QgJQQAZlng3ViBhKIPN9nG2THbv3rG8zMT6NHx44EcRRvrr3D
I0J2ngv5keBT9aweT87tP46ZzRrzMKXdutro0M7m1qD1rL3Mb5jZObWP5Kl7OjCP
CNM5GMxbs90BJvDq1jupH6upSiIpg85RZVYhrlbir9PItt0CBJHbrYQ74IfG7awE
0fIemqz3LbeqyMIRZ6x2pJAikTk9yYjU5cBwhSBAzKVqd4zJl37CVRA6AFQ8qB/4
veNy6RNHkdEI1lei9NcjGCePye2xNGmROzX03Af33bq/ANEbqZtrqjr8TF4gFZmH
8JTrjSlDnAnRAFyS+bvDzD+fAwoqyN4HvMJ0CiiBeRhtAdJXcRXNiIICzt0+LKw2
heiwEyYdjtJTviaTuZuOAZ7en5+T8tRWaycSsYxbevbhAYSDcD9QjRQfgNyJI+l0
GKIE66+8iQUhbc685Kjvx2q5dPki+lvb/Gr5P1CnNXlLvqBsbeOBnOVMgSHP3FIJ
nA1VslxMeBuv1HbPAWTL7aQSqValOxlqAyAMykHHULn/rmN+lq5lvpZtiy7gMZV9
3CTm1vFa+ETRXkn+C8utcJIkTx62QwyZ8tDHwtq1d9gy9VK6rOyeaoj6l6hM5F0c
efRxSJo7JmhqR9YEEDDm8jm1+0Yc5DECZBTPm+LIgpYTmnUZ9MuDkMUbjn+Iwrya
p0BUFfa4nSoKCpJwvob+xBuIBwTmAvjqQA6qstJtafL2vQ0H8SDV5AswRWBynEEn
TE3sLZq2Mb+LUl7vMzNuAaEu0vbFiuQ++OfV1m4d02WPzSrU0LteSvmy5hRsP4eQ
oCF/OMmHMSd8rmM4YY8fafC5Nh9lmUUgqezvmcZaaN1aXy0mYHBNuvK6pzO6xudr
KFYIqK428g0TprczSewtWksa+I2YGCCm3xWzo9GDpnRuquXO0jh3KEzCdIxrSoov
xCZAbFDDSsdcOZrxOBKgVbI1JnntVOie8K3DqzDOLuqwmwBR1HMkS9UbwWh+12+b
NoZhNolHq13dobs+by4l/Zh6sUJxj9wgAEgrsTaL9TzyAHM8pHxVfNCGXokKGQS/
I1GjjCdMVA/lehb52FyKU4GL2SB+opIjkpvoDyIjlvgrP2HGfno/v/SVir1IfzR4
/nwJ30FlM9SpmYRfVVRQTLyeaNb8bss2PPZMxnXZcgV27FIh77x/y5fA0H54Cj77
bohJ8SCyebgswnZPltF+t1+zAeKCkEO61WpKMqm+khsfkH0cP5N/rmPn8JajSxwY
tzOQ5N8OoTqW5cJNr2sxAfNpTpl2ebohfXzFoujLGVugauwnbxFL0kRhWRPcC3ll
LFawBreTtFvqy6DFIFyZLhG/3gvCtOPWj6sb8Z1sPbMujuGTFTnxbeaiOhigE0UB
jSh4Dqef5XSYqk2GAGxdt1jzmi/bZyDZiQYPX4OcFN8MYb/a2s2ph54Frx4mC2iC
q464TlBW0FZNyTjzEQVq7L9RJq5PGgFTTRHL9xtBiajuKJ47bd9+QQCTk/l/xCX5
Oj9N1B6tcMh/9Vlpw/+Ff4PnybNxRR5uAzQc2CtAngn4ApbQyqWY2tk6x77IZnyS
D5EFmKwpT/M4DMDHDP6DYT6bxx6M/xxgI/vjaFbM3kHFjPs2m4Aq8RlEcIOIkp7C
VmOyMiqBb1CqbF+/27leAfpERjVeqUzOU/5QdfuKrhk4KhtrmS+3oIrrDBYagKFz
QtMmcIAPaFaGENTX8SoAa2lvKJB4yTJUG8gez/qz2DLiMD94ihghUlU2rZtT2pLP
ryAze1rf+UDe5ULr6TqGR1i0sFqLkFNvADcsHHvc8W6b+/BPGnZzfO5Dd7L23jz2
d36BAlNjwq62VMTzBh/lUvlkOl0HlcAMlyAcEoDeLn4v8YG9XPdZ6xlAk/awuB8U
2zaefAktYOEZAW+Zi5vkWz2+II9t+SuXZCaUEwqR/P+6SxDn5HVIn+JxQDxjDc6I
5US/cXnrXHMJ/Uoq0COxkJDl16K5h1q53ZrruurvVpWYfX7akQWpVwgbE88znY68
uMmbP6R1hszEispPBOGNhRDMe0yD8VOZZTTix0nDYxlNhJZ0tGOePC848XP3rbPH
7goDF0Xuuthdz67IRCdWsbyampyrY4m+UgtSOjkaL6dczvZQsN6BYeqKg27TvQSe
ALc1KovP51fm91F5EhUNMMP9q6SRC+tCzSsgCEJ2fKygtK6veoH4oO1M2zOTxOac
rHAnYyKlOGxTJmIcluUsb9JXmDR2s58YIgOOXdd93hR9Tqvj5QrD11083Ja/cVGX
1DDb6g9l8mavQ1vVGETZ8HWHeEkuTJrrt7WU2K29xwB9SiOJiZITGfD+/POmJ6U4
Bc9YDo3viW1VA2B9OUk+iEeA0RO3/dC0lGjJfo+Hw7V32M1YmbVrSmlsrGGmUvQH
aGfKLqh0xAYXnC3s6fO0cZFSmP4iDeYYzCxUowWzF6L2DZNuJ7cl7q4UYKoBTBF6
ZxpbYkFzJzDCuMT5NarXezP3GOwRS7OiM/DFpGTJv0xu7W3d9FCrMnx9x4UGJr/B
Ln6KHXM5r7I36HbT1UGw5BNUfwTx/ictjXkbCJLbJZLBlxOGeiTf+yP3LDbWRKXD
WHJZck6tV4h2hz2kNIgFsY66+ZdOuadGYnAbOVTKKRU5VmYpx7B5Iea4Vqbwk80s
1oX6wFIxOPfxU8j+LKwZYGTjFDNN2UknCtwfMcuGfZ2GkPQ9bQd/nRlwto3zqQVm
oYJqjm89W6GCvTm97/t3hESG8U7nyQiCVNs2YSkE38GAd/1lqvIkrPu5Ai2DLTNe
5Yvt7KURiEjIX0P8qfrsLysiu+QcQ4Dn29E1/9EKB1dBkanb0xlXSCWV8ChSYt3M
3HGa9qNejeX1rRpnvDfUUV2H2YPJv1sSiSVnnL1joNoFsJjxWy4/Uz9AypboFDNb
g9JBpApIObGSCfE3dL9xYNJteEMqOKFuRezgL7+3KW1mdG4KCNnSQHorkTJoYPDF
6qavZlThfwZuTu3LzJFLGobPcXkfzRw5ZjgJdvXDhXY/dmGdEBQkpELRMOilLaLJ
WqmGMrlx37U9sEg2W/kBke1g4koXM63icd+id+OkUYKh8+Q3Gu2hfjK/vmRwyvWA
37lSYpyHlsjgsMJU5brz9oTfkGe1cWY6K3AJf3DpR2WF65vSVhdnrshTECT0dffD
Aydopm4CJy43dqIdQ77uUUxfywBgxDKgW+ryExmoswQVTFlqk8x/Csc2+q1tcwX1
nmQ0MBC1zcihpHR+5/gTyiJazn9UP/gD4HagaVA1zS2twoWandixIVmOPw3Rzv6p
5Gn2h7KXbLakd19Pb3x1cXHDwfTga+p8qr+HmQIUmhv0ZUGJOWT3rTIaMGsxQhbp
2nIdCTrLxjVvf+muTWC8JElT/ixHSpAuD7f/NpvCtycGneZKHK2PD2/Sgd7IR/Lt
tG/Cg/lOvW4yKXLVXX2LIM9LB/D4rtEkVSDHzexH6pTJEmXlxCuujRxPu92cXOyO
ACP45cd4CGpfM1TxRwl/5P9AJR+Vrv4ZWgN8w118ckDyIWSRCkdyzX7Z5lQwMso1
agjDoKKblZ0yRcOzlfO5jWBZ5HWcv8VxSuuiKnIdrLxQytnaJqP2VGcMizel7GkB
owK41icccnyy5VBKbGlNFtM5LkhXm8YaDQh/rXrkBieZHreWSFTriikh07ispb4n
kxX0FwaCJJtKHi7kHwDNxJhfsq3C4PqMvYAbu+E/83kZLgHQ8hWMYFfpYNztICaK
ic5/1SR88k1SFD5mQby1LnqCGWW55d/lndBWQcNxMGtogAK94sGPcnhmCZHEkdiC
KRZm8deuA2cRgFHZu/rt5haiuEi9d6eZUwtnq7UP4udRFMqhhziUcCay2PtJ+9rV
RNpmAoI1ZHGMm/9129q3CndhAnPTGnZOmpwQlmK1m0y+fEZc4rvE/kKGCLiqb2IV
HENBbYdoG2fj7O4To3CyHhRZXWNzCq2SfUXw9rn4QFXlagZaZ0iDGC23sKnpHBrt
YOXm3di5iRIuVwr6MSZlwDesQ6oYyVcxmV+0zrHaUsKC+RK+DNLGdXBxghidK+LQ
nuv11KlAjpCtRAvpv5rxRQ3sM0YRNz5h0uHe1RWN5niRpEgZA7Rqo4faazfk0Z7U
kUtqPrC8V3ig4NXYma1kT9XZOa6c+QvA4iwjLH7vZC/C1Gd4UVUTLTy7XpOfMABV
RIlJWVLmCUIPCztI0g6uahH9QP1UKQYGpG/6aULotHw3G8W59i5wle9JPpXMbR1N
9ClS7K1aaco8WaN/opBmAFje8nRLUQskpBWVctcAWQpGhblFJ39FzMOkSgnAxGMw
qw+y1oqAE/uCnhkHtn5BsvuRLPd4mSeUaAWlO9bz5CvwAIWG1zU2i8gOMcVYARIN
UMSky8ak49526Lh326/qTrRcicWvk/cgwmvrp5GodWIokFCp7WJ8zRIpBadab0RM
D/MG8na31DE1XodRMb0qfey11K2HNdtK+0KlIEHXn0OrNWwONcEr68yBJbYTx52k
0KY7W010V8zrsCeYrIqtrJo2ygXlycD6NznGK3DDSlLp6fxiSEmYBlLYbRoObhnF
n0l/LLjwao0CUDxQjPV2axCKnw0dE1PsUweNg9P4VfIXW3mMjzr0B9moIqJyc/CT
gPbmfpyqkAjIVuIzl9gcJx4RonI6gktlkNLQrTC3TDCEMGD8abq6b2IJ1lYsmmac
Hlg5uy9RU9SxXOzKQcRknSW4/NbuTLkc5/BOriUJgJfeqABScSG/NcRsFbqD0tX8
BiwBKHHACEQBpZk+BkKCwk7B6SEtVYb7BRu/wE1xaRW99XUi/kcVMPVHem/guIwR
Pus4qyiyRlbKln3TlmCs4TOIDTIxb95TBrBAJE9tH2lyS59Q6PMPPVnO01TzDtrm
xtbLnqH6ugrKilu4jnmm9j3sfUiAeZokbqTZFtbBvwPl4sW0oQliwZd//3AsmeJX
s37JutZJPCLPXMfPtzifzX+q7876TFcBLV+8jCntRBqszQBD7aRe3yvgpnJ3Hn+l
adUjMrhu0lU+V2Fa4F7yImCss/f0cb47+sPWSxtrVNt7qbDqYiHxTatnig4ROabL
974UI0b8HuWoFO+fHdpwRyk/uA9rzN7ILE41OfYLUA7zLp1a+y7o5dTJEprKGcBn
TAQBibM91vCPqE+MPjqtseMNtK1yWZWatdQZQfXbYfDQrNZZn8AksWk9zCF5KoFb
V1bkKAAo2BdlU7UwBau85wf+rSNf4r1EJdANmKcu4o3KEkQ+06Z880jv4x07aZUw
z+UhxLniGpAPYf95XV691JaLoe5JkiRQDBBLGjlMz9jp/cKi7FdbAF6BheotZB87
hweb+fSDj6UI0c/0VV3AvB1rMrbxozMO4WaHy7V+xkd6d4GnusiQArYVyyQO0iW4
yVtejhRtY1nCABqcob0EqNbjis48V3eNEe8NC/44Pj7qMZQLek5IyfRo3LVfM27l
pKE+bx1bSpXhn7uTHeSM2OgVdTJxsjxHlymrTMHiC/3RbkLe112IF1shjwRi8JtU
LQZU+BWEu1YUQL58DEg0/aDJItRSgwDJK6SItfE1YuE7BugnbEDqZAU9v55KbhOG
Fmb3J4G47GJnrktQ7RckHmhV0jiAH5rlaqP0gjAooLgzfI72wlJKOaZknzvGq+MR
+oe6ehS0NEKMz3G17irT9RImEUG+vZ3+2pnodcNrm5+L7TfOjMpeRDld8HV3/TLv
eO9KvSoFiYCMBIZM4ClT/HJcLdOQ4Q9smGjVYUvwn7BidfU5fKo3ZO0DayI1ChLj
X6lIi3sArlkirnEzRK4tCAT+h1wfUSnuMRlqfTUzgrUD7H21Swyz1WAa5pEiwOJl
h+/FTolrx45BtcA5OEAGRVaLxOjlJVqrgjn7uLF0Jp+h5ten/JN/G/hl6rB9uSYu
QhUzJ//I1nKVCxqnjTNVovKS2INlB9FFW86IRz2IjRU859wi9GOjdC4upf1KF9oM
KT2ARqtETXpvUJBrZH2DwvpRRKvw8vmHiq8Ehpb/YZU10UEH2B32UGXovk9ES24r
gtv72dPzRLC3/6rcL+apsMtUDTbXPRoFttZFKerWptUxXS+Js4G6xzMQQKXsaPGL
BHAhdrd9O0vBecuWr/C4tC5/5/nxIJA9fSPIgaV/2Def6OMKOCiY5dRQwNHI1utR
W8rxfs2UIqTnJ45Nptc/mS6clwbK7BLuOn+rN/VXFPxys/cfa4r+qbZGaNevy86/
pCkAvoXkJ46aBzhigJHefvWwq0oKp7ySOaSM+IEyQ5lNdPFUhdzBGJgFVidNdsii
mF0i8s4oU23vVP7haY8h4AarbrgqlEDW+I53h9AbODm/0Vg9QLjouhXrnnLX7ZvJ
kws8hZqzt9pawByT2kLX1xEf/FeUVSBkDMS45Y8vjZwzE0eQvMc54glKfp2XZ0kr
ja93aewlFmHtOCUfPqR+2nFjkg/nh/H8MwG9rQ3NUe93HN4ppKwqiVxu/+OEKz5A
KN4xrkL1CczTkQhd9LCbQ3LS8SrXwFjJr/EdQ1855DR7nFZz0fggmKyVHd4ggF+R
/xDUKSAGVI4o+oqTC5oy6JWpN6Szg04EkZhTQ8Sh+iqhPfvRhE/SKbY02hmu7GMS
jvoe/dNgRhRihluUCIx9jfUyKraYlixrBaPTMrJJhaZsrBqpId3r+zU6CykKo3PD
OZT6QjTO04XtD+s3NL+9yY4iYcEFHLPR5JYpwweTSS+kijW4LvzMLr/4QSJljW6r
RXeaSXb4QIbYXBohTTmmBVpE5BHZXOC1fvPcYCexO5tlhap+bXogIFvgX1pOqffE
HvErEYCXS2t8tgDHWNBssvPN7o7QZOmJTKFtdiQgFLfnWdS/ocI84gQ53p3xIcoW
1OP/mxTxmCt/L7Jf89nA0d3s6YFk+zEu61gGWrg2NkqXDaZ3jUFF6o/tJlfpUHF6
D9ZAzfvPc/SkILbgESwfTN7cnjEczKUTG/24h7djc2vTSp3ZGwkHoGYDxdGHqBHT
3daUPUXS7TJZR8gJxqU976IR7d9DLm8tMaDfuovz0nxNol4D8711dPkdQBBY+T3T
/MJXGvHOHj9WogWCwmnsGD/6oi7tLZk7cYeGiPQRegBM5AA4bNX68xREqYa3gHfL
m43TSBIrPdRqSreg30CG/XiSxwhnRbj6YExOZ4HBsRN0xx+mvVkOV5MwsW87eUJv
ImasRYbxVXX2rxMo0r1asq5mgDHmGrCbvuy+bG0PR8T8gpzBnD6qbYneQNNi+i09
Q90UAz6NBS02HWN5nqiohUIZJ1J8CkfPHCxGnEvPdR2PbMyppf7y80yNh6ZNqCBS
0L9hwwp3buCD8ptnJaPfxIqFHPQvOiZq1r53av3BCh/mFn82g2UlZLCT7zSXN0K5
SvIb1TnEJzzdtVFcv+oEZih/AnQ+ls1iCdfXnOtV9PiXrT5toxVWOUw0htpCGoDk
NP81xZiPqXMhTdH3Hugut4IqEQW3exzRQSLRS8cdZYkhlAyiKjgDDMJVmMEv4w//
MLGxfQ/FDrFltMuXOV4D1g9PtjKHFcvgJemYd5FNoKNrhKc+KXY0sOQJXXhizEFF
JB4+lugyUo114yHusRcxiz8w5qBSUIN7ID5HqAJkmGnHGs68o2OUV0ueVs3HxhSE
O9JS97tRLBXlj3IfHGk3vvxiujucYTrHelFZ72CDrmY8Kdw/hECcNe72Vht38Gh/
uZ6vuJ9rkB96/zuudvXGAYtYYQk2AnKfyLPXNiqbFe/NwwSIhxHaMHaQpOwI7MIS
tQGl7WklfT87gwBMaimVW8tt8td0TN61Rhjky47IWH/AORHq/89ZK/eJMfuj+534
2jBIiOQYsxoIDoibr1qW3Mm+uVZVyvnbiDVFLVzrTRKUYpP7hoJuaUwdJx0AIYQl
zOEbNl+8vqOQWT5g2xUQEqUaxI6Oy+yvltxLKM3gr6V+YdtGBjNk3aaLQxkNB4Bz
iIsuM3CzO3qvtrw2exPGfURyet2ZEhL17lQ/dtzIEy7M6SALTBRtQh8voriaJMwx
yUe4Xk13//NqlpbSgHJMRnxZEx2E+o/O5I+QtgECulOFQOECW6Ybg2cggl6UkVcO
ma4vkJd7m+HJFdNV6HVZo4kp0PDeP32+HJGTjsmF/nB7XsKtIidfKDMDd4nkW9g6
W1miBctV2zNMkLISM4W0HFjdZC2egi2KGh841heQi3T6478kXg57yFM7EoMuZQI/
MjRF2+kW+Q6iKiMpe0jk78qAL8oxnzJXOgKO0TrrQ2Jx8z20dYa9ajqLtjhXxFQf
A4J2qt+ydeP5Gam1sicKxRPrc8xWnGKAt/2hNPLcEfpPUXZUxiWClnIGqbyARfVI
lHhUzvxSEwJzfSQR4Bv2hGdEw9HQFCEj7PvflhXkOPh7uOGAwQ2TXkLPtqc2XabY
cEjiCnidzXnu9mJZC4XSar74ST4T7MAgYpmFTiCi1fHIJBVn+/s8DiANbfne/jBP
hg8Zqh96PknaU56lG8FvsdABYsOB7Bk/dQnpQWXAoAw7oo4ZVUHp0D3YTfJbRCDK
yW+G0OpiVUYWVKx3wITsiT8UQNEENSYv8yY7xh4WnNt3G2UAphVeK/3HG8/l/Lhb
5UY7MKlzpkkMFTjhsK3yKBiLGvSKXy9Alae6ZQfrOAozeQVVWzkd1SwEkF67WyFl
Y2hWnSLJuUmaPsjFfpHRAFF+34UUWp6kL4D5nJyNNnDddbqbKS+SC+uWVGHNOyry
kcP873VAB58qRu73HLveauy9O2VzrRQHFtmWRyNz2Sx6s0eJiGSw7efzhMeZxhK7
X6T7ZFzLhLUDSAmPHfCbJBrUdAdYvFWlOVc4DvkeOxt0avCEVLCkNlBfytrjdoZe
/Jvd/jlZIrm7XE5bjW6PYchNkl3oYU+lhZD8fIbifQhMmjAu3Z2eAu8aM+Urq41B
J2tWl3z0CWN1MslBy04IUYGLZZ18B/mLDG4zvHG/8BIhJLZOm5ISbZFut+LMQCyG
gNxPcHhoEHeEVK5hCKvTY42B2xLjw9OquJgbzVrCsTWdgD3ZFZoS4KSFNEzh3Fy+
pjeBiAlMyztySAxdEaEPOOVagJPBlZ3icZW1rCiYMYZTzYDfm3QWYfz5gmaE2l6g
MoiFA1bvD3qQ2k/CEPWRdg8V56F/pg3jXK18RDR6uIWAgH+QkmtKcIZJN10VjrHn
B+ZfLgrRJUmevCY34h5cBe6PBI0nIF/69Qbf6pS4anGyY4xublXjJK7eDbnlhChd
100KlV9ODKtYoq9rjRFY/WSWMDwaVPgTQM669AeXp59U4p8jU/2bzNz0UiHIORil
yvgEVUyGAHm6Yz8Kc8/F7vPV040N0Quzk6SeduRRAVTXTpp3yqvFCM0Dcbd3UHNs
g8sA2XCtj81hdtYXDLkqdeDuEkjeZOE7Oi7InNJGSwf3GcxGu0f/HFdHEEtVlCWV
+EYxpxHkdrW0X71Gm1iHcyHMXS+JFiJhumc6oNc6IvyT48OwSJJYSZgWahzgQ6s7
Zv6LUtelZAyqOEikrs286M4ipZ9LKeZHAv2T4qRDpHo2JPxOj/2TxeBCGf0YKY1Y
eqpeeprGMZ1el3opOqi4Bzf3mcjDPVh4rOF3B+McbelM/WVDsBLVof4cCI7Rzdhj
M8bxjfpxkLS4Gow0hHBjwGqEiYL7DKEIEtMqCBsCpehk6OV8mTso89Fhxkv3+SOc
Bd84So7oI4XSaqfcgHJnls+BQDDukeE/hBAxbfKMEuTdK+scRHdSOSy/Bs+sMQu4
j2D+ruEEpAVdHi1NFpIZOsW/ltRtMRzc4gSaizG4D/gb6QP6LT4YZkdxWl4ietXb
D5wQLxpWCPjhWyysJs9Vd0w1JUmWQiN3/YSeqwaCZ7yTvsXNOPZmKqfU/XiMTkvm
kisOrdbnmVkyuAEINkD4oreUeg8NATLp04+4cUxAuOcYHerZbBCoCPyK30ZcMFTz
oTdTyAwIVy/6G3xPzHBnbXkdUufV5nhcWE65LeDSjvBYuIJsEkv7LDn4fWp10zZl
N4hH5u0mAtp/HFw0R1wZB51MhpnDijpzfvI8AvEauHqkClsD7ZkKDIHP5+V8zKxZ
YAUT485CM1I8GEVMSxGqIOVB6ZfONepYYwCHQxZuqouev29fp0KFMuvHDELKYbE9
XsEQlnkfc9IiOuRrj/Myfs1PBECAlE260UXr2b33KKYPjzHdQRPikquhvXL3Nag4
Mr6qTFc721mNsY/8n896kaKwSD/Y9/+fntlJoCsC6SVK8ZzPwTaxbJgTItzPo+X5
eNdaECOoGRfHQvcXvEc1gV5jATWmIlRdMxAYg2gycO/39cFD2B1e7MnMbb1+M97B
4OZXx/x5OVPC+gPAix9L1dUOafofHxA3BJx0ZkaIYqhcolgV++iHttUPqMbMOV+u
UwYenTgST81XwJ0FCIk9lddlp4w6juG9Mm+zQpT2SD8AqIHBm2jH8KvqIDQSO7uY
KJ4ZprIdNEFlP/BpmuuNahe+jWE3kvdNd1AFi0gMRRcVCbINAhLM+aQ9CdjUWUuE
u5vXccrMVi1ox95MCWYkAPMzqTH5Xt07+6Tk7mcIINXppPXH7G4VZFAPBV04gO0N
TleJD6/Z18m39mWculotmrzsrkkR/z4Tc+bqhQv+bChv/Ms2K7jtxMjzp6l8tdTt
FiSbLnklmZCG2mxLMF626rT7ntXTaB/e9yvAdt2urh5qcx+2Go9VFp2LbQ0QGbAC
R3N2Xx4EwdqJMpWdHxv2Yfe11zND6TlLfcKq1SNs6rPYKcsRFPVjqUJhG++7FNWJ
4kQDnQdVPp8pxXM9baHr7XugAmksNL7Y9TuCkIIRFK9WJDHluM4ay9rIz5jx7I7z
wOqkAUtanN9+ZyJmRBuo0qT/QjzjXEBKRYRkS2VO0PGkTFmbV0tMk1iJkCYGNW5N
MM9KDFIC44xnDIGm7YLy0P+k0N+KK6YdLij4R6YgM0BK5bUkFqK8cWwxGa3MOUiB
MDbwgPCBNHqlbJ1QlVoV383PjQ7do2zvOjKuWl+1gyO+d1Cie/Mo97wddRgwkXN0
W9UrD2DrgjL8pBR+9s3Tr+Oc3NfF7JqLGzjj5vtGbp1xXxcG70/DFTN/VSVxYEEK
/JQ+h4I3wPALdCeU4ueUOqtpIe+me1wG1nwdd6D3eeUgT+Eob5VYo+HBrrDXNUuD
/XUp0uKHlsWD70/KRY/a1NLyrc0kMIbMsHcepr0hKRYkKStqEbwbF23CitVF0keR
c4R4fCUrDITOdmfIkFckJfTPTnrur7PuI8O7A+awQrR15ygVp9G0uOG1QPFyGSX4
K4CEzDTp6ptRbenhGVnVgPXxGeWwCcfXmtL9/lhy+uH2Hm1rhKlBIQel4axLzUwo
d5RGVveeNeN8VolsnKD/n4XoQw4EjhCu6wo8a4ExsYHR8BCWO6inzd1MYzEQZH4t
CLBsoABw5JAMx7S5lil+dy5eKwi3cXRJyUH4FfAqbMT72pEJzoVJ5I3X1VbhQLFH
QUrltsCO90qn0tbmqqB9gaaa0l88QgDwN2jKDMf0YFAzgtgotOzgbFbBc7Q+oS9c
sEbYFbgRrMq9VO0CUo91wEpsgUNkOtnTCVj3n6+/f9Z5hqpMMA3k23wZw4VcDhim
uKco1QyQO6pyTAu5XTcSnpz8H45hEYkrNgJgkSMqDpkxawwxdeoXCg5P7FkvKFuM
mr5ciTJ3gj37T8PiGTksmjpOhMqj2a/53rmsdfdpjXltz35GamIx4x3lqwjEiPJ4
O/HygMPlEHRpfA6LoN7FkZkE/ivRF9mtOd8E7es622zQ848zU4R3upjBdyZf44iy
rsk846B6NbWmZsG0Scfgzk/9iEOa/+s2NSAI4rUMRM5euIopHDuChPw4VGrSPZky
hVr3Qo7qDOoqBICAlH9d4b6WLfyYD4M5SZQQ+T7gFnjomTEoQ9EaFBIrNqyIsffs
53DSksy8+tOclcOVA/0mR8XSnxRHGylcB4j18xxr4VXrmYFeR0m1g93+XyOggcl+
ARO9DXBZQqRYOX+cY8xl/n3m0+brpyHbyuu/eHW51gUTIgMhkShNRp9fhBIuuhQb
DH6xtyEFAZ7A6SZmLGkn0TD30y7sc1VKaZ0piubnyH7f+uuLaH825w7W26pzB9FB
Y96zV/ifpP2kta+Qc9YjLUtR33MJ4CdC6PDSidpbnhLqNMV/Gcx27vEivjp+d6T+
Ugb+dtxgxrtiHeKI/rvpP93DUAlbzoLIG6vShgX+ft9VDuHrCLDtxx2YE63NHtef
I8VOoFWsOOLXo+27QkFLNm8SS481Ykp476LtzDYnhfvWF66/qcWIKccW78E9yXYg
fbtHP/ds+oqOmFdyoRjeqxYcLb/JLtcLM6t8y6VSVK7vqt8qtym9hIXdUdFetsHs
sKZrAYDgeX7UTmwE2QrotR1OiDjRK3Y1EEY1vlSibM/eqbRSf+nZWQ+FRNHLv86z
GK4NSbXOlTkpnG8w/dZiSjvUyW5pQIGLG1iEgGBYdrVPABZAJh7zNdvFuIl9gQNU
9+eM2neDGnpl5EFoCkipA+A9iAxD/GIMt/fh5+KyS66OduumzztOn3ScHqjG9Vk4
XSC7aN/YYdPpIMJDHKcnhNRK3LRzQJqvOsPRl5tu72TVo1RvWmGBEN31DNKAVOcC
tj1IuGOjkvKesd7VCXe0QW1e746NJIGLmUNzUMsvho4tUgwUokBaDytxfQC0CiPV
yxQh4B15nihoCwTeMel2Di0yJ47obLIzS7SYDUaBv37XTvhCSkRy+QK+tmN6R9Xp
FZEbwospU8o6BVy4t55Y2fkwJ1tkRewNNDJt/wNcA2K0z99n4XM3zLSGqVNSywCU
CBIuZpdNQ1FfblfM2Af4dOsSPlbjdbr1idizozJiKcZRppiKe/SIxDZMapzRHxgc
zlf09us6ZTHUyoNKzexWW2575b5Rk6XHl2i3hDUetVMRWlhyl95IZoI9OVOrkNwh
l/TNQVfVNabKAHgwUckhpgyaxMzyoTyd8c5vH7DMGjgafJU0y+c9gL7GyDeCBTwO
3Hbn42iPVvANHpJheZtunLzNcYxRjZnnMv7qFHWPtiFbzyZ6baLKv/7nvd75N9EG
V3o0IPoBQJf7FS/63C2LPK7T1x2gETGZlujLXEpiOKwSsynqJFxzwYAA3Q/CIU1a
yeO0VOce8850xHLVytatUUAfZOMR00El68Rwf3VgaTdh1fdwgJCFH7Sjjk2NygT+
jfUtpXNwr40C0AOLfZEH8SnwFfEBiPE5r8SZXjdeZYciw3DafT3I4foavYmo/hgO
slRGR4g/jmdHOgaPYeYUoNsX18O4HXIpRG8+WJv5a7rVMyh7+Mdgn5z8P5Unhohs
ahKLEonAmZeOzO/sXFjlPy8dXQZX11t4QjsN4MwpQfQu92GRWMVVWn3VacKVLrll
y+l4ehTJUeMA8y0WRnN9eZzd8uLzlAT20xGqHLx1Dm7NVM7TINKaB5+u0sj94YTg
5nTAghjDrfWb5y9fbdlQxpycIAsQfgqlxyjILBNmEK/pRzryZH0z9WnJBbHgxBk3
xUJHCqOarhT+bhEHiCqIynktd0syx5GVZ2lpKPykSkgTzsUZhF6/A9QSojYrAB6t
/kz6nA0wJrTsIbCHXpCaNIfV/lt6Ce0SYxflWWnXkPsxwLrC9eGJRLLgFUXN/KdB
yJfFTGETmEkOcPKxQURKJKt9W1gIazcoEfuzwb/a6JV2vsrucZ325PS4xT0dvZrR
/VdhBEG2cGm6NjJUD/MctTaBUli0CNmZ+unGqk3xj4tBKk/eeIWk+2xKd1jjkQgz
JupjP54gTa6SKp2v8Quk+04shfVMhOcouq9UEr+8NmvNNMB1EWqNSFi+gi56jWpt
rAGbTGctVGeU72afx/bKEsBsmz93JAJiV8gQs15ni0ryKFMps0WA8q+DsAK7M6wC
FJMKRpoc0zLdY36U/Ni8anqBJGULazS8lW6ylVl6jJZ0GRpE3IV+NCDPaf9sLfxV
Y04U62+EOOeb385HM8F1D00emvp5Ew3ExcM3IARMxIq9T121Zy/e52l1nhjD3QmD
WkCzZC5NmLB3VQc3fzWatE8Q31CfupDxxWUUsVVsRr3/RvQvbcsWjIDVi99uZTgK
Sap/i9zoZh3FXQ3GG9dgiz/2rLzVKgk2KhhXq4ZcvLmNxRL5RjJFnIqu/v/QLSCT
W6C36H1R2XwjYGUPIxrX3euz0DxpHvkyhbsdtzC6g/5ANHVo3+s97iej41mH48ax
9eRa7cXLRIXOGCfjTMuNmdWV0BI4MD0GBu+YxMkX6NihjunSBxzV5qpI+D0U3Zs+
ja3TXVZC2MJhR/BQxEAx/2wwlZULtX1tt0H+vrgbVxVYjRdYS8iCvtzMnz0Dj6Nn
C5CZ23oFSIDCI9EADpwS2CoUBeakqRX2YfgIvw6eI7rcGYBaCIPHtpV/htVWaLGA
8APGSmDWFbohWcTQPauieq47cwLFTMXlOprZstOWNSYU0pnffyPBubOqTPZ6L4C8
0ehAggTImcNxX4YS3RM6tWF5xVo2TCJHzFiZ47DhDbOOSkYWFZnCkDOqveyPIaor
CvqjqJgxOacZ6FFp3+YaTQozK927T2fQy0u7wu5El1NHx8nIZkvTHULRp/qW3PZo
zB04alULXzTaOffnQZnahgg1BB8EUoQFhHwSbOZjR7ZxlGj4V7L9FKjKA9Seg1AH
YznTh9hq9EwM1Swm5YgS9RCR4j9+5JG6aTlSqMRrLdvpdU0XBWQBUxjRk39QXDjA
0vHkawTKsRx4mjaG0TS/FVH/bqM26gYaHUAcYvEtY3f5ktEyY4aYD0XtORLmPGGJ
zokNdraYUtxXjtE5OofbLuCRXRgTnYnNlRGewcxAvpSG8FktVZk/wPSRX0kQSCwZ
Mc3r/IU43Fu99dEjM5ws97v1txILevXtThGOptLxnLUK409FNkOUDVntA6OVF+Ex
iR05XyNxi1I/qKKbQQb881GzveFhOrnSyAgfrpXjkqlFkA6YugjJquDCp/fC7F3i
0wqDkvPWXwZ4x5LGC9MWvNKuZZcIXIpiLg+9l+JkFvUIuT4f4gkiAyqSs8Wu7UyG
qPijT/oPK34ne9/mgNkHzRAWY/nvuKRscSRDuX+8lXWK5iRb7IcKvLTrcf2ANyQD
42hhind1VyQobQpb7n7rX2M2cPwA304ECKxcXv7VXKl+ER+DXQt5LwNjM9rZsXSX
vTBYWJxz9XCm+tP6+Bm3PspXe33S/0bTawF3c48A1Lf5ptoEc4E3QGNjGW/C6qEc
wz7V5HELNjp7Y6pNI+cgSZ0WZClkGe3b1C3Z97whJXEUZVdB3xLqme+BUKew/QSC
hUhFkQXmuEw8SLADm6GukTxhReINDKlcNhe/dVhF3y3EU4jXMW/2dvUBEopC2k/C
C0ufLt/qOlmoQP1nOUkd7ttj3IvVA6/a1FCjm/dvRSHZDtWPto5CJe3aBsMD1f4a
rh2+b4+rxJr0MZurCaZpY6NqjalVZfTptMAgPjl6QEVqUEFjKrRzC10JsnheRdEt
gUHLcIGcnVBvTSLXmTbxQTyJFsIlFbJU4l9uJEus7KCN9slqv0LoOMQ+NfiK3fTV
ywNgvaFStSwMym3hRHhKTsfDWW0cJH1EtMEMpfXRHwTQyaG9CjUfIWUm5tqvBNXw
ueTZYsl9F+1mAkBY9NwH/oGpEmjStAlAayal8sr4vEfwKvKbetTUsI4avkZ25346
TsKknQf7uPgb0z91+k6Ha41A/7FutqRXGxhejKftQDaFZRL2Et7rHPRY0/JdyG3R
JViLnmc+5gW77ohglS9e8TaC1vD5zuoMmjMlhstzwr3jbpdU1iNNnUjje4E1M91X
kStsxfar//CA+lydts8GPVGNaNdpr7gtVsu2z+Td5xE6NAK+MU6P1XwL21emJRso
Wg7e7eA7FKukp8YGJVYFwVLHlbuJr1Xm6wCTuh5Lud5WdHA18999msGwk7pYdueQ
n3nxKcdXg0AgDrpXX2fCNFyT6tpX7GJHdwpgAvWKeiHc5epa7DV1Al1nqgbfdaCv
Y4uctw3XVgYrnJ/K/6qG3inye8QkciQFqJWUo7ch30s8LwqKs0inw6YoyFBFAnf0
DsipStBWWsGDhQIvqYhZOqB4egYZdL6p0j7mS8gcmj7PB38DmhLaByFCI6TJydzz
kVTYN1be7a6LCNq7AT3H5jt3T0xt/09kO08ZM2WXpKw5rG51IJXbgQzTnIF6RifO
ZLSGBnxI/6x2sgf54Ltb15R1VjviNaVUWVr8fP8cgYQaIPLp2bD1I/TnTCyPiFct
TtRArAf3ywbCkNHhfdfDt4mt4eA/4w0s7SmqBTfrxTyohJr0X5DWnOksxPfSNZ+/
nz7ZclY1GnK81029LQ8M/wr/qvMpbP2NIVlopYwzplOmmxRViVPzAyG4ZT/jNh/Z
0ZdxpfnDMJ3/e23otOt3Owo0pygy/79JYg5Jon2zgbTWuIAoyALIjgWKaUQ/8b3N
Ht6UOrYvHmnn0xQGRLuAsCqmtTZg6yyqIZeqQ6J//Tegvda4RIklPwiDddmQSM7u
ZUkAYevJDQjSS5ngikSC/KTP2JGt7agr3RiqQPeOWPBkxIKYCtBJttVRLu/MhGml
5u6BP4141ZY+dbVCT/OWwFqewyYIc21jDDzmjqhp6zgbKq7DHG3i8wtOOlJ4KjY3
qXcCLZb7JZ+kztLcA8v6i0EEdAdHTJIgmiHQhUMwzAtOy/9pLPnj1GlpwYdNZ2h7
wgeYiLItVXNYjP/x9eei4AuYB0W+mhSmGrC0tT0hB7l8220j6eei/w8WMlMAAxks
Bq5U9eyLKVT+WAG1zFrVuCDdzG2BSa7TUqvaFasTz2XbLwPGCokI7/BtAlWUdWKU
keuhXmsZKV6fliU+LRfDMH2UdT6Jeky7CR8/qeBlXtXstovJJF3kg3+5/zSpOke5
54PkYSlPv+hNxe752a3LZiQEfBUBC4Ryn3B2ezYhjQpy2p1n7/nQR9C27hrker0O
NPj9QkBP3ZtVY3Ierc10SF5dLneqJkGddydL4cgTiiCBs3q1ysDZM3bpQQ8id6yh
UKMGA2pqaYqZaGOgvuj/QpXzNxxrzGqq7o9hXGDPi5h2rAEci6tDRGWP13kRQAXt
NjRQABD7+a9Rxmuan/pYtJjrJKbZT2ccvqN19UUufvOm37xhBtLVBIpRsmuvGlWu
HyprKGXK7V/9N0QAoTPN7FRJH5/lm6Igd5+2Gu79eJveJxJ3JPHqG5KSZC9xr0yL
HHZGIDgcLNRvCaptKke8IyOu4Awh5AmgDiGvaI9ROD92GeDHEDd4IWBKtGGxp138
7CNv6TlZEuuKPS/XLMHXLHMZ4AcTiW4CQetGFQwR0bhk+9DfqszFzR9e6By6L6MT
WdHuhTqFWlNKw0UnSQnbLsLBYYINz00mndLUg2N0K8KfUo80Vs8AI6t2ykRb5SNn
y42A4zGONsqqdraa4YhytRiQjtMbFv/spZ6HSY45So+4QU27J8fOG8ABWPIxsKTE
Xit+MkOJ04EUVqMIMB7ixPkc/oDewHLmixfmziI+Vf0WNn/rNRzfOChMyx4ZTdR/
lSFao9JIHg8vV/UZCmwQI6pHoMFQiJKehhLtoU7L8oke2ccNBtCdajXDYn77UeHi
x+QUSEaZ5y24Uvv9jslN5tUk9qaB/ttaT5u/RWgBObYY2S5XZXU3iOy6nONmB30J
DrdbTrmCQgFbdpOw/y2Pvf22lYLu6PgRvvSCQgzh4nDZhldRaX4K8//fDilQ1zuo
NOMMO+MVrO77pybxZR/rH8FeAZLbxIMjH3aPA8txdDDXOGxavqKSKwJZ7Yk7Zesu
40TUh6KH+ypvm6qjQpMrxFys6G5JCstEaBxI05WG9/MiD841ZKgNDScKjdRwQWwi
ZqEhhVyoh3TZRdhY5ab2225fHQjbaL8WdjiGyGzaQVFQ5x00Rk6RaaFYNhamy9Gf
QkeWG9wvxUInxRfl153j6FTMKN7ZV39exe1rIZo0/ee8Adsuqk7GcIkKEbgKfIDp
AE31/g2cMe0bFmKMYnmdSJQ2k7pNNPDcf2GuDEKk6lKKkLYwWEn9xITzgagT4YOd
UnbziOyo7VF8Y4OQUAbitjfksJrO8rrO6yjr5CcBQP+fQes8LA3nZDPRADiu+0Wh
MfvpPZPq8dF2Ld7eIsJI1bB0nf3hpJ/zGkG+t+RAlv+iuwLAQMsGKPS9sT217iRX
GUz45s6VBASKgwFnLoRx1W1t73u80JXSC+6VJdxfEu+nXbYlWkmP/tANOfBNf5di
FS2bujQgGK2S3rHqNYMofbBAPdZiaA9J4DqfaAf5MCbF0r21gKOg9Cmd+KM8waEm
8YUeCkcPNbk1I6Zc6/cg6lkyH1SxbmVi9AwIk5O7TxE7AJJjXounqnYcvn/yT1iq
k+jFzIHDlc17Q1ggA8Qw+eR8U0soxFkiuqbf6wpQY65Mcdy8CWY3FZybllKx6pqP
oJFf35+hENHZ5xBNFbJRtjrXURrB5smwp8/tJ2WKFpiixs2bvxUfnBxCuDgn3OT3
cADubq6EVA/sYdATbLyhIO0DxLOLXQFMnqj4YLQ9OiXSWG7FCbk/LM7j11gmuHtq
pCo7PA0RrWNWEmQREnsqVMooJcFIOVF58UNacS73z4qT216mqrEMec0UYpmMJ7E6
gKHm0Hdrd6WSFYz80lTu4elH8wMSmCE8ClPoxRPbxvKHThKWCIOt+BFf74Dy8EFe
y0NHWOyChEOu7L10hHG8z4ZWVrajeiLqwOj40yUEz0mK2I8s8yahZtykSIu9WIeV
AZrjQ1v8EOykiRBbq1SXemGryLSx0cP2WiON1dUhBasrtHq5oRLRzVlvZd0XF+88
KCNOwNYE9j6sXZXW9Ob3ie5ebOUvQKcxfTONryXmQC3oERHmhFpn+VlJvIkJV+BM
4/CqU05wvF1DZGCBV5JU9jSGp4k2BPoY1DC767KpM1hPr9xTzSKfIW4GQjiU+BAV
BApA2pndPOHWyY4Z0nH6SjVJRfb0kq1cI2c3/bCTfYq03o5BopEl4wBmN7PaVn6C
82rO/csini367T1zKJGHB7BH0HZeyy5IS1Qlj+FFvXG5MGX6Ns1HZ0krdQKUdJ1r
i3/mBUVMMDqHrAA0TpJb9eKDFq+MWLbgVP31G26vY6zxgpNbzf2IhTq9hduSAIrg
ecHbkWlzDd7J+7ZvvognpOVU/xF4tt9wUu0pBiMNWFO/YqPLPsB93ebM3IcwgHtl
XZ8t2RgaPN7vCqyTpeLCRGjPqwb4PVejheTVo6zIz3bbdL63et3t7NHfOqHpCDw5
/8IvXPqMR/GRyEdLNzgA6+K7zc3WowDgBnnYRjETLoMX+3A97KxwpefjX1FnIqFI
ZnqlLVc5H+GunPQL2cPYZjXueF4c5sev//10czMmpWVeWI25zU/Z030wIo4xxArI
0em5TBwxFGaBk+IB9Z9RtxskM1OLiMusWZ6qoE0m9m+lnq3YQQwhYYRM1EjkiNPU
1dbuyTNShMdUiVFu1+HFx+yLQC/D/+goAjXwORkLiEtt0xHjqw5aEmB542gwA7Jn
E+r3fnLAU2EXz9eq0uUkfptRBuEoPy7ysWwdNNHDaD+jaDO8GYU8PAibXX721gMj
CqVoLQ7YttjY49eZwRKGA0XBOsZVrMSXyrhv7ZPUBP328tMmxRpdv5T/FlHh3RaX
mql0P+JuqcwnMe0IpQFwNCwTAcwjUghkwiHqyf3HIniX+q/645Wmhx87MUWNNa3n
82/yYihqLGaQ3DTyU5cSEJM/+WDIfIdRdUgs1ibVr4+EFORBoQ8YT1m/Hj3cFd75
lZua5u9leM4+zmZjDh3K+QArq26b1osBGLmzLQ7xB+at5urWjVXJKJpYvla9egwv
1dOG5gQnFwH0v8CHL77JObpeCnERkPRSjZXVLNZrxmcaPHQ8fP0LOoPzd7rV2VzJ
LPKxm1Q0nCO5HBtlJ7Tz8Rs5RRFtIaTw3u2/LRIcRth/FZxQ5P4ZEen/XkA/kTxa
ftjfQeFxfWfnACuRfb93gGgcnJynitn0F8nxDAlTGKzcXCragjBgYGFHenzITHbm
fSU9r9HUL1VgBzEjha0bnvoqxFiPxft+RIWU04R8hGEDZ90TX16MNIitz2EN/EeF
guJ95NJjhWULbEnBZ9VxGvjpxUb9ZEVDP/Jn4iZDz10X6JeslAjAc6igWETOHVLt
s4tKquH3Bplq/YbqAzW4rYLdd6XwNqatbSPh3KuLWLfKKgUogbQ+Zk74BaaMvOYP
6NHHwQd1crzDekkUEJTQvhMxTewyKd/rjv7jqVMb88OELats0l+a4DbBDb+4UL6S
YDrkx7ZIW8M9kz1bI5/Oq1enHzn6fqlmh7O/11Bk7tiKdtIEMPP/Lb1tDZaio8ce
4yiy9WCO6k9neBGIBCTsoZpOuuZe/nMUSiKfLupigsGkLJfo+im+L+Hw/Rh83jVV
6wCbBR5VUUEK3MyYNqwFEFMIPIMNVooL2PIqMhp5WApQVBDTjGwj6V4xDYnZcXzt
QU6n1s2MktPTR/4+CbBeavXTRW4+aAiQjg9HZ8yKEfXPzdoBhst9/6JGzbSyBf/p
wg8nvCLGwo7OJWeZvzBkDzmAc+3DDNlFgZTIm6D5z/7d6vjnAXN1Bf+ksZq3g/lc
BCjJc0cQUv3XgQaxDXtUQoyrrCUiIykJM3h/2XSb54y65pgwRafOjsbDTGsJRJKb
6HGmGkfPREJwZPBnEUJhqmjlC/rVak9OnqEiqD6dSY0REl3UuKBhDFN8pUOdwJvb
yEaCg0YkCnmVZXy+aUuWk+4Ybs+r+RQ7BoaSEhZT0A/YQJhFxSuIhyHxP5a2WBr2
JMUgTdbJ41krJODtejaJQPy/I6Ok1lZhmiQabP+3pJ23kyjJrYQ/Gksk1eiaq9EU
Lu8ADeolOuW1g2CEHeO2JwPuBOI0HFBBJatajuOEIibuuE08pyG4SQOj194v6QZq
fWalcPqYCjPGtYc1GwfzJtcBeEOE+BlDkronc/LQPIu+6WZN5DEOAWmXiDJh+xyH
NQSSbYnDbkkk29+wS6lNkbyvqrgOMF5pY4Vk81qoyQkv6IP5M0NFlTSTnk/tVRA1
XSE0C7T2oD0swgLTVWtcGgHf1BijZptACOmdODFcE9JWVrDPSlQ8hrLZNmj/cIcl
UNQV54tlIiiePgXKLor3H3dzixwIhf+Do1JRQFmMPtpYGIlpgTroeB8YRkfKnXzI
gh7PM7cjN7wFFWVDOaQHvGZsZ2dYUnhUTg7fhQEgJkiYqVredwNIhMYTGKQsIGHX
1VmCYy3dusfpW217SOw7hkM8KnUC/qxaKEPAGskUkaYa5VpAX1K1zJhq4quRutmI
ByOUq1HKUp5cgRnsEbPoeGEt0qg2DXjSIpQXYfEwVpD432/ZIonDQYlO8qvmW3Uy
SptyLNegTnCXDiHIydgR243CP791qOiwwNbsSmczefuVY1u9VHq5Z83o3RqKezRr
TZhMwTGkbrLUxLJae5YHDGVR8f7mUCvaDOuM8eOcS1y9uZtaA4WL+V6iw1z7w+Mn
9P8j+we9u6AmPgMnSkdToWSuJaCjNEt2wV2+eVlTEAmu7id9Bvr8x1OP7/EvtZ5O
BPq4BWpwknf44SIMhNlK2jdgspq7NtiqnPDeJGdSEAiPA3AvD2RD099Pc0JgbE7q
WteKEavCqk3qzSQbeedGoIc3liCn1P412gu99IP8z9J1kEvf8sB8r//2QN9pLr+N
fvr6N4uZVwxBEDrVThJZjuSngCvxXQXemB4BBbVbP0S+cSSC/8o77kYNTertisX4
sPMbUjRbdj+SVOLt9829LlcqEgAqLgNenCV7oYhAiC6ewaRdaalH9wkyTxvRbPkE
1qNLBegjCzOhOi0wbeIXc2KV3N/Qm7eUds7iAWEpW44PY9aJVPUwTbaHTJ1ZVPW8
pVxYaiKPqhIAeCI5CRJCfczTrCcn14N5ETerYLcBzEzvILNbMVpmC4UlLuV8c1Xc
4hPKGjCjnOgIlksC5r/oKbfOVE6JUFKppCfgAxcAQAjp6cSBtE0KDDtotbm5KG7C
70cGVHLC5djPMWr+85RomdlG2oby99cjzyynapcHl3gjQCkHTTsl1LDLAUZ9TMo1
wCOOM76Stdmo6z1qCHtjiRhy0lku4M6fQmxWUPNkYTMYX4Btdn01uYbFLTDWISxD
J69oTwT3AwguvU2q9iYysZRSF7OKeFAqgmihv8MTsv+86EemG7Lml0lT2BrF0Kni
GAS59hFU+E8ziiYdC4HQXGZPUZLIUEV9ACss73RwjMQmPoGJi6/fztAlMdbYceT/
NO3QsR26l3hq29q/jCeTwWg8qUOzVDX/dLscCwobyrN04n70iAttlIpSTnZVHbVu
rYnigz8vagKwRh0VZK45lDx7g3Z0OUYoP8tnb40kl4A8mfVm5D197kcq4npmU5RW
u2at7zs61ZxTbDVIg9LeyivQA1P+MW4C7HUymj//RJDGiPzSy3S6fiLDKeI7qXnv
bFAAkVFZaZIpscB29M+AhEv4LUzWdfDtYcXQvF8uuPzoBo5oaowcEWvQ4uj4b8k9
F0TkDSPX2hrdXbsCzhazytxJoe12otrCnaAirFTbjVlW3XmFKwudkC6zspy8bXX+
5eu5RkqzoxadFFzyOjm0F9pm6kE6e2ED+6LNn49e73TLtTPdt8oRP3zB/MN86vIQ
JZsScW660OPuFMMBYeCHss81SaTFVyUcqWMkdvErJEswYppSUETwsGlAek/i51Hh
ZHBQ3G4qHgfsho04UhQddeXtKxnP953aldmhtJDZ8X2VIC5hd8zd1OSO57xrm0MC
wnNcDEE8uSRVB3FzH3RHfBMnaoBJFfoBWb/Xxm1JZd5l8ilq3JZudrTnzaWgImPD
HzoJNInLua7QkMhGmQftPi/ZEjEwN2z2zk2k6wNjRmWpG/gL/Vk1pkp6Kezr1eOO
txyFBq5+F2PDEWAk7pyLXe8TQZH3q5f7eSTsUnGmODFqZq/JaPuU1+/k3KsDRocg
J1D6o9cSGS/V11mfaiu+5gesUnJvwQuU5ZFgQ3SzSNv63v6rCaU2DwY00a/I5XM1
4T2FGEcrNXark84E4PxXKND4ZG3BMybERfiFHeWMLILJJo+xyWvYd+pRCnY+Wx6F
1aUSex97EEF1tPZEiSDYhpvUP+l1rgQ0i3Uk9i1+l5jxX0Bz1rLNWBiG9ZcUDrWx
QCqeyof1M53LFcIST0Njj0g2vjaeBoBDSff5HcnrQNZMFvvL15P0AlrwXqtx7D8e
nJKO8z/u8pDobAJbYlzol1HF9Wt9KAyYqHN2UoPchwnHsnFAxz30VF3eO8tHpJjf
hFAFX0IE4bnYiARLa19TX/V+jSgOX8XUIuktDgVNiQCZagq3NVpEYuHTuFvblCtw
YVWBrtKGdpdvuIQpyjJ1zSOlvAObpXuIQDA61R45gAZu+qnIt+TRvwzVDmowycwO
HEjn5lVfenBphng7COJPZJ/LR0xp3IkC5AMqPf5i5dWW878wqRnMCgnHACRti1S0
eTr1p1OgNwAmtCjnLeQoQ8lLOb1q6cDKG8TPr2Q9u8E6HuX/nj8UYDatqCFbmUHz
CUTzQRo/LUIaB8lvMdZaPf1qYu4YsCxDVLckaOfex09sEIj/YSXU42I6OR1t0WMT
QFudzihD+h87d+VSKXuWgQPzghxHY1iYat8nf8LCg/VLTHwiEmw35Tw2USoJuZl1
wvJib1AvCcD+7aSD5TPxhx0wu7C+02Evq+Pn0TxKzLBGV3sC7WqHL+m3JyG3HN30
FQaq4yay1tfM5GrqmFhNcnB8Cmb6ubBSAIfylYpqLveb9zV5yp7E6cbiRl9kqigH
HPw80qyj5a9WoxCc1twchWHvSk2h1IsnKjDPX38SYThUNcDzvLs7NL1EaS4NqRR0
2YX0JhjPWyCEP7mK37562EFTy3Sroel2eW6/iaixgUEgqSUzAC/1/9JCDRLQ6zsR
Sltgv0k6KP7Vw9dwinPPq+ARaqsaATgV0iRCsShY9wcap+zaNZZP4e05iYcT77WA
GGZztY9yOE493VGg+wxItAXHDrVyjoCpMROMMmV4Kaw8LkX7SOtXhrnZXJIRvT3u
ElE8j9QwzidMoqtsb3UfoUNGj90rS28KufOS4ijXyWiZ9zALjDyVFeEoDBNKhflc
ge3BI5I1cjTspgUKK6f2u7O7HixvXB4KiVyPKIlup8P8HGFcdXCmjxCvTfln3tQc
Nola1TpdY9Bv7XhRinfw9IPbJU8bm3Dae8ZoV741MKFizuWYOvIZ6JQDxnI/Tjz0
Rs4IYyWAByt7UZ6iToazJwFkabFkHhqXLw09q5xNjm1GmYH4b5lh06niXFcdCPZC
Yx0eNt+IsmIJPb5BJC+CkIo1tB34m4eTgH0ATf73of4lFaERbE85MQjnOi4swYog
DR0GPSuNyl3uF7i8duXYHKJSDJw1vcKb3DZ3yyLK+hQiaODINXKv1D+4enpQzd4c
6EXjKE9DQz8fHoMMYNj754bYmnDdeSav0r6OCzja7eQEIpbuyw6aG9N4vPBxCOIx
ZRtoe+ND2bw3fQ8RjpUBZrRDsjemruE4HzHJyv7G4qUO6VEoC/g4KVqoFgszLrPT
Efwkq+vtnt7F2R53Bi6xWaCFUa1b3TNJUfTN++BlQr6tpay3dGyrO0AtfnSFFLMB
zSUZisuLoLuTfUjOR8I2aEdWxf2E973Yc6rDfrzfxa0c7kuAEoQ3SKFh0h5rsPmF
0NKtkQrFjpc8zXq/xUsDuCQ9pc5dx7sJ1NHCG7jGThrtVcZNnQ/SMywV09iLhRwP
AJ9DiHza2k0Yf7rYgW/QA+4LzOH8XmQolTgSBDJLABlQ68dJWAw9c06XBpbtSmF+
q69uoMp3nBYgy2t+PktAwt8rNoTSm0j/eLnPtYG7Tu/PCv/zcn7V1E3QXVHcP1sh
cYNeXi2xpvzn3533wu2ALUIogMGq+S4IgwQ+A2q/WTawfJDYWaaw+yuxGhS+RqZ8
ZhZP2Br9Rs5xSx0KkWB9+ixn4gz40JbxvpFrhgGq81s+b6XkxbH6GmV0P4TeG2dt
e5un2lZEd4JfdUODk+rnYATTE3F2d2owtugfCCsMxbmtUDDlUkIkh2g+EFJMCWKa
jx/8GnMLBWOXrsJywrpYxsEHafS4QOvb3LmTyzVi4UAA+mWflQSJ8Ys5ZZDoi0V+
RjVNFhNv68d29yxv1rtKUrfwxmCUtw6+T7H86oqzcmeRCgvflzrXsWR54moDPw7o
u6NMxXsckvV2OaHrM47c74si+eNQkYPEQSt5kyScIc4F6rqYzu+R7wrDowF2Q0R8
OFeF11ak+4ToIg/SKge1IhRS6QVXTODLg14DIIPc2kIXi9yrZaFMJWcE6fsTbtEL
Yz52NkgI1kKGNfwh7IbtyZmUvVh4jH34zeyhNrCT1Q65TyJjo/8z/Wr8mE1d31ZZ
bpL1QQpefdr2JbsrsaZMqGIG0NhYismH4lFwM5jHayZfIz58r/tQPIB7h6viNo/u
zzHgSNzQtJbmSOpAOc2Z9fpQJGC5SrGjApbXhaGrnWV9RQHHArEovoeOobFYEPWx
8b4VaIBCTi4tDY36yuelUOl+CIqfXvSjL3vkK7AI+hgxXs4C4HVmPSDTuOasj0HW
4h+At9+InCDO6I4FNTxu6aQUIVi+3paflv9PgQKP9vkmcfnLJnSQhElWceaX/wxt
uc3kxxApC4jcQ02/nea4lTt1ZUs7237HfCJh6TEbfGo3HOqgu5WMpHXol0dRmvKD
nTnkjEc9dCTPr+xUP0B4R+Za70qP5n1czeDYV/ePK8qdDwykxmldOffGptDj8/yP
TsVbH9iOWN+3eJaJZIfF/qRYjZvLxz43uYuUFHF2fqm7F0Scee4EVX7SE/WK7Bfn
6/J366+BAETsOuVxtSFKrI9r6FEYk6e+SaLSaagcl1on9cGH/UzH9QeIADsOfIDf
1WVoVnrnaB0zZ23nZ1BNXzzizeG8hI1+OBZjxY3im4DttkHRfFkfua0ob7DfwV29
jQcOq/PPVrZ6XbUHWSmeHiRirbOMaDDu+1yPRtpXiOdXMplfToyqn4bA+gM2cs8T
Lyub+ea+WfuIiyQ8FO1hQMtBHj5+uBnBpEafu6YoQE6x6WTPqihBbZJ6KXAKpDOp
3iIlERf3Ph0a0Cd8k3rAwLu4zosj9bJMt6ePdLJDiv7J0Mw4bfPnvoBVy1VttNC7
anUIYLE5UsVGLOchJsv9c3H8yXwEi6eWNSz+UUc+oOohvEU6bTspNTlCtoqzeF5l
r9YrHtqsoV8g2b12tqOzD9OhJx0WIpp+J/yNZD6R9jbQlCSVCtkjxFk3vsb186ul
hn56Nc3P4mvDkungmsadTw3vH3aCphfbe/mi5j6gSLrrqgRsrHGy0xSDjAlmtJzC
97Hk/1ytIn2xVa0tBQaleT3Wwxe70WuR0uFmKQKnQ6g/wFXnR9yFwM2NvLXd+93Y
xLPcjayA0OThiq/5kx9NMih7Sd7MJaPFkhDXrSR1FlwE3Osc+xayXNgmOQfEDGX8
a+ORY3Ls/SkoDJu/quoS9ckKe6q5hDWV3RuBC7nzpzpUJGCFrp9ZlWrYrkZ3Kx3a
AhnBYEqvsVOm3LOpZdSLgbzyNXikrVMPnO9nTCw5vS/3CByrIjleolu2WFjwc6hk
Ubl/dmp8vKmTCHmuFuEiPeOrrJUNAlqFow8hxIza4EnjnwS2Hj8swFdzD4HYnBM2
vCl4h9RA78Nh1tAzRKg7GrwA3fPQqmWeapoeTIYAPmOtMXa1qQPZAvZUCxErKc4R
WEwDjoJ0UjDvRDvLjios0+n+RkzdY5fE9CZxpgZKYT/ji+2ijFoM4FVdnce7q4zo
zCwA4bvM6ThSiFKj88dgC8I7laiZCODwIM8dJy2MwX2yoMQdxNJLDz5e6NrxhooK
GqaDl6QrESV9BlIC5uyT3U0CWHP/HpTAURW/RjjjBP9h1BllIJ3QIidRtyosOCKI
9aSGebwatR25iczXWXjHG3aws7VBQr+0WxbtGG1Cp+pj/5ytD6YPuqtO1a7saGyq
KdDm/i7huqLWC1pcO9908c1A3q4njwjmubPNyu88qVAXRs7MG6X7ORel3ywv66Wt
yKvYKNoWSKcHFlXHFW80w89qcu7mP9b56M1X7dzdj3B1SyYkxY+/0M15ZLtAqfIx
HzmBRHosV/ITQfCzMBOLrRWuRyIi3PxxkA7TtKJ201mWBrnR65yzZQKWpO0wgIFw
lsX5ZkVQtzrkd+gCAyiJO5QBOyrU+hAJ70UgTSGIpGWgLjiIPy65vqMRChGTJ9uQ
dJpmO/Rnl8r6JmXCrPv8GkeZsFuJ52RKnrxJ9+xrRdi+mi+/zdV/MN7PBwTV1ydA
ShseOGXn2e0IZzOGknG+PNX8w5YwcQqRFLZphJtlPbfHH48PA6/nHlh1/tKdMel8
RvgsorX2WShBoE4+XhFes3yZY6M3NQxtYEv2nqGXka+NeRsDFQ5Na86/bbOVfI+i
kXEZfU0NU8JamlC6UKHD4jayabp2t8sPPKfbMaU9MUG22KIFJ0UUL88l545+nyKF
6ENqUFD4kzLJFE6HzqbSVP3mtAboEcvEbrpL96/tODnpsPyZoCcS1IDzSJNa+f8/
kmIwfCB9WFdlAcuFuAZZyxH3N6LWmRiL98+zTLdol0FNQL2d+RMoNf4hUAKHvDwG
an82ilG+66c+xwjOacxS8P7pyxpEhCXUoiNAKpPLFjUSPM8AtbIpFt/CuERKhGMr
BB93JSXBF3onwIqmHOo5j9zYTQDhsLKXjJronWyChXQcuCSy63aUYCSfeulbJuBA
oMVsqen54TGcIvHpeMzRfGnEw9OEqvSZrlgYc0sUCjfWIccFpPRM+EzL6odaVa7Y
NbNXoSzmdCeVQulVv9SfSPmpx8rqWiV50X8zeEy7Gbwv8qiHfa8yj6Ks6nlUZsPb
eT5K34Tgo0sFABbJg7KkW5YjysUWRybZPw9lAv93zNuEvNWgzw+XSVVqDJY98aAw
WW1eOinru06JZTZgIMcTzDFQtKHG+e2T+aVihTGa53p8AlzM/GlKbWC5kUxAcwlD
fXSjmdHsDoHuPSDJjfqQSf6/YfW1HDV0QKYCYtDK/OYiTRk1PsSG5kPAYEEy9eos
992nwAK+k7ZzYaB3602mayMlFWvlEHV4Y+TWteBExseNZ+qvaVYJEOs1rP+7x2ui
xfm/KgFt3Y95Re1M92/hzL2msFZYKihxbPp9KSK0UHcFEaKHmHcG0jagDX6gt7cb
o8U0zMGi04oGuxdO5WnNsEyxpdaTejEZtGb9uqkEmx/aaEpQMmqU8a5CRzi0Akko
qkVlt5GBcFz6+UvD/UyM8/uV8YhtUZAUKB780fgQqnvFeFRwMhYBZcJvwaJ64C2V
k1gdDzgmhqDo1ohAHH+YYuOwmbGKs3HrlZjX1iyGbNG+jU4dTIeyuu/5XtwCXpsN
MtvU/Kto4Hvhs2S97Sv/YHbc1LGuT2NAcdWdcMqx6W88SCpJDD2a/hr0Dy+B2pyC
B8cRyb8kqVYq2xTW3nwPX3B61RuWO2pr+7VnhskziMeUORIGHKvMPFDlEsibHrFN
MjLhSz75mtzl6vOtXcux6aYQKkFZE25/ehFs3lTqOi3rWBrtjBxRgpZgfYHkbYwm
+P22bvKzJk+4G+RUIWq/zQ1cvfKuT43nU3tuxQbIMHumiOaNIHy5HkhuTz7hJjf9
tRYBlxssxevhKrJSH5cx6bx2AvCGbSL788Sa6Ffio4eN47EgkPKjk0+4VDVK6IoY
MRM8wxtmuiJseOomRzhv7sKQ7OjdIChm4AB78mi0QF/QBFAok5mD94HiWZMqa24q
98fl/lSrsPaMFfxaVYCWQIMZIy4MZIIoCWlxkaE6pAUgj/3xl88DlBpI3joI50S8
g9NTjib8Zd9RQfOKx4ldlFgTiDi31e/BMS3PpH9hJVu+5/Sb9zkoj35Wle7wXJ00
uvmfSOeFc58HSlqSV8trZGxXmrJz4saN8uZwowie+mZY/0EGlFP/NnDU4N/KdUBi
8DYS1OraorMLTstGHwl2l+DQz5o9BUV/iDgLY4v+Wampl7f+tZT+wOBfggxRlE1h
eakVD0T51daxA4jMFADGnmx/3q4Mmfx8oR4dZ4pDbdl2E6IWanGAQv5UNrmRBHQp
TWe58mbkZVsbvP/llSg9Se+9ZagTN1EYDxMAedCMmhF/FIpEbVEp1VvLvl8S88N9
3qsSXozdIj3VqLKlFGwsYnCF5VYFq93l5Y4y2pqITkaRF4lcMcC0UL/eXNjitlRh
uZ1hhJz0ArgQeKjkPl4ybl43bGqISrxOJEcY0He4vFCN92RN4DFJfYVVIiVXSeRf
mCEAnqvzNZ3HuuInulpgHwXxSCBGiUEP7DJ3mCIw9p1pBlHClZFkm4uLFRw+JlxS
D2WRrjjw7c3RC3A/7O2xUUz0NJIMund11Pb6oee6gYaD9IUkz33FgUzt/Swq0M32
m+RXmsdWohshrxT6cUtv7iV+CWOdSCbEIumAUyfgvrZfhBngDkJL14xcHYC9bURH
oARIv+yDAFnSuVe7rtyYGVrSYX2RRRoGRX5W2FHY7kEdpjF84S966exsZV3j3weV
Hu58acImL5LQcL748Z3PfcHO3Tjvs1WAI2tRQ0Rb3pcbv2p5AM+ABJ6wqvXSzR9j
iP4p4h8jF7SF2cFnvzLFT0oAZtHKe0NZXl31tLuPcPaEwyvSoG2W4uZWCjGDALvd
f0/qfObK9Zecliw0aZeTzM31IYXlLV2nelyJnM9IJhTh7SHSRVq/Zjq8ezkL/SIF
QmrHAwpHHZyDVOJYoOPqrOyA9+hzXwn7511DUP3y+6XDz9hn8asoVnhykGBfTY9x
3mHkqZYm1vCU2uRupHvw7UsKkJCvsUalGNE3f3uEij9s6sASa4Cc0Uyh09CsuPcQ
HX8AbMT6hkaZKksbgsMcl7vXciXRjbJTz86n9NsWtDOxhKDyBIcVq8+03VoCE1AI
tkHcFDdJrYSkpUo21thRiBaDlfgZ/6SHAjVmi4BBvXqu0xJU5RjArsVTC/gkKZiI
/ddT+yi7ZzIt4PL7uCc5Ub8059rWqC4Q5qTvIr1BHl8BuYeHy63A5foHTZhkFypz
KSKmg8bhHyFhjYwg47m0Sw+nI5FAEZ7o7QppEa5zepCll0xNVtJPj4FaMTf5pL3c
0sZmW7gbFPvSgkSsKVlVqOzYPCIPsRbEVzk8Xe+GbTBKae8z2IH0TPGosEtNDxlV
5+QFF4JVGnZcCcgjVi2AuWSdAvAkz01R1Vkzg+bVyLY3Urn/9QlBPTWwvCClr30w
9MDTSZFJb6zIiOL9L1cE9oTH+syWtJqot22upDPcm7CfDdNfk8fSLmOkJTDZUXjU
SXZcDxFrRmqk903LvZ9IYnti0qQeI8acLT0yGYFuVsbHgITsNXJ0Ji4vybaVlU9t
IguwMpR/a42oe26+IxvC2JxmtRqLUDH/096+9XjYJCI2w7u4Ccn9bARbehNKg5DT
IDqZvG26w2ZvgJ6vf4RqnlebR3j2tUcrS4BcaMP8fyrhgm1smwfyP0HEiPniKnjf
7Qs+8wy332uWz8hfa2AW0hoG10IAMrC9KC9Gmm8rrgSOCMr5gT35KKAvBZqndDc7
7jHR21tt0vmqYwWADn4AK+h7mNIGxw5rlZ/X6+K/PHSkuIM49NS3ZY/VAsV5lm0n
8Bg4kscmplO2JMfzVDfuupGZiO7MDalDVulov723yUXDGiZewdQMlogs8DBgU7HX
qFc59p1/rw4nXcc0OiQhvEXfHwCj3RkTEEcmnh3pdskgcvTbsQcKZ62oSOwfif3E
CzgWcPJ8pQU/FENBA50X7AT7QplnkE9sfEuTSB0dWxm+dKk16A7aU29bu0ibLBFr
jnDZBsb/K6tNAScpCFgqRZYtPXqddpeoSHPQC595On3wwlrGANnCtB2GO16GbQ6g
8d5Nmik0Toq9biDjZOIu+leHsMgojUAa/U5NRzm3bCia8Dtv09hwbTj7pd0vrPJM
aUv902lnsSxXiXQnvw0DxI9MGgz5+XiB6D5ioIqjAg8gSwsTvo0nn4oqOPM/TGL4
PtGCJbfg0y2VKIWs9S0q//6JX1kyflXPuq/rEZ1d92UCxTaxXCna4L2OJCfDBnZx
jcr6p/KZwe9uirLdwbdHfwh9lX4CAEYl2Q07c4C4cc65pt4KrNi2r2976u652Eye
LAt6sbaTs1EvS2dc4cBDi6yGrg7v/keOkjPubM8zQbaWmziaod54OI1u+9jvbuTi
ILvmQnpaE70YkT+5aQKz/svL5fj+xfllUroBzFWYcHHvGWbgNQNCY6b5wtphLv00
xYTLX7WGX3QFxls6i/r5/Pryu/1ZNex0bEbsgJDMDd8CArF0bU5CinIDT0N7OQ2W
BAq7dd8GULTk6SuaGStMd88TcGvPrZxvItWwzJGLkpJsR1bB9kNS+JFwHCn4U3wN
stWxzdYDuWPjXWTupxnhlYijHPV+XzIg1J/O24uMvyE6EEX1dbA4s9rp4LZau/sW
kZ16ODPQMELtu8y28AFGdeEvtqWL7mnVTk//Tz0fIm39t4v2IMKVd/SopwMnYhaV
PSNqsS3aWbtz+h7vCNTL8YUo1KW7tqKjz2rg57iB1nBNWTb2WhklfUpXN0rz2mvs
LeCHnB3QXsy00pvmyc0wf0pLsheK4Fn+hHqZSVb9ecX6d5kDNlx8xMVpT3SJMFIq
1PXrlLkii9kTwZN4YsDjnOXn3IF3P1TWb/Gb6VwLtdTYmR28vcwtCA7XXCRpngX1
PqQJdMXJMA6VlMYDxGNal/9KEvDBOXOCDNzCJlK6EtnDoiRbYK62z/6GyO+IDlRq
BUAjJ5/WfbeAlVcW2KXzwj0i/rXnIAihFCPcxK4JusKMnCdQvekJA8LwEadjnF8c
R2rOpKQI5wER9qhwNIKV388gKT7k+Bv6jELCD1cY179p6pkZKuNnZuRvLDW0D2BX
ALIlOgFc2uHCYrgFCQZ8IfffbAxg5MkZgsbAYwfupMWDc92ddqPXslT7q3JmT3az
kSb5J95RMN6ubQYebDUF1NKVYbSdxQRPu03tbSAHdAt/20XkLMLS52AO6hXEQ3md
GWnyvWK+0CBMJUnQqbny1htZqYHuS9kKvnV5jaIkHmMbQtf1l5J0TJmN7sUw28yP
UaIRzXYbEwP0S91Kcs4lpGqbbfYdJmSB5BSau0HI0wc6E1AEbq6q9X7Dr2q3k6Vz
h/uUYm9q/UekQDTpPKqWSwYNluO3DHAa5uDqLKuG+whkXVyR5JDWQsnnOw0rzDNs
OQkCdgV8TuGKKz24ZCOvH7f4g4HRLIWG0dUPGyblg/SyEZBzh58dj8omTLRfI16A
+/rYozYD2ztNF1qBNc26cgVBZVV7MejOqKNjLcnqPpx2azfUOAGYAldgltb/16+f
yvh/Q8wxQbVV+Qk9HEPj9UVDoBmsu1CDR//vYzvkyV1z3ehi1lAXKnRZ3ZJJUkf6
B/XIkf5Tfzlt5P//bKFkaUfBDJMOlSHHoJVuVwBcrXub9VcoanguMmFqR2wF2q4B
iwl/GXgJDHUoC+u6aPDIjEPgEZ6hoZnJi0nds34CDh3UxSDVEu2tsgFBWF8RVQ9w
ZeGRoobszHxTRzmtdoabT10tI4F1y6apQaUJZi9BzB7VT0Xpi6Of+UqX6iPkI4rp
cW1cIU73G32rBHg9/wit21/iDqzIW6ya5BnltviIdvJIe7qzpSasXlXFV+/W4DFr
drd8+ycUtmXO90QbXwpxlJrp40TXncekYiTOTQkMnI4p6E5rF+khf5M3zxp4cFsd
L9MA99VUHrpBVSOm6GDsZyt6Dsl+uiY11OE/6DGPqwBX4AyzO7QVqlncitmPFPTm
volkn0kBgHc8h3SuoAKNQPYkmABZwpIVpPI5S47y35qblbWw9wVLS6wS4CRXHAUd
uEYTQYDv1QkoxXtB/lhfBf5N2b+3T+VHt9jzrv36Oo3IxGawmgH/uy/SmbE/+qJ7
FQ6sfr7IwZNTx1wp7JjmaZgrcuc9mTzo7XZVsNsFcTEYhUwsBuIFfgVD0N1s+b+L
T/HSqpI8V4l+t4HQ/UWwsrQ7Y8Kp66LYdlTftzXacGmojFQtSuI7wfqu4owpmT/L
K/Daf7IB3qg9Fs9XFgOHdrWegDF3UpgQYlH6Es2Bd+MUDcfqfG+R64ebDaH/c/en
/U9QnfXxJr6BE9y6sMTJZHSFvp06heXqz82yuqqnEoShH1vmpsqpSsunmR9Cfjqo
MRv2v6tx8GD9EdvQU6GwYQ3jie87f6l1+BC08x7tyhqbJbMJDqhRx7eXB5xSOxtR
8pkyHb0VsIbIUgG9wYUAWm0q1y5LKKW/cwO/WFoOuVxZua8EdAJ4muQfsWeBPpYT
JON2Tv/Ypi9p6oiJCJ1Jb67vOwSvLANlcph+2CND+Xy6cfB78RUQdtJXOUC8hLwU
WWnixXnzmIIzy4Qb5PwwDSpa/89zLBldMglUVPrloMW8ADhcP4Utk5c2uZ3B9y75
e5IfJ7BBW+TnPSxRWmWpewLfmA8wCUrAqNHGlZUIjHNrJn8VI/Tn9ZY7uBldzpn7
bZwG+mcu6jx/jlb1P//7k9qhqhlIw9FyDlWRQv9ZMFcCF44j4hwXEmxktcJXzuP4
gLg/bSit0UPeyo0sDche9pF+F5jcpbGERinoAuAXviHpuLpQeKTPYJb3MA/jIG96
yIEXKVdzAV2EhmwMyqbvA4/GfP/HKPSIe8QMacfKzYwzDfsRa2m3vo6K0PxnMaJL
7oqMR1BfqEqdbc84q7ww/YetfrP42b1kOjpwbkSGA71B0gf/Edb60G8fD3bBpX6s
Z3t1hvlVJJOJjx6y3qMTVSuO5I5Xb+MrpOWLHlIAwHNk0P8G+24wXlMPRGCRUCnv
EqatfO9KvGn7HxVCwujVrYHnQrmoMfuK5tRsKMzcFZMAz0TePBUb9Ixtmme8k4PT
5qQHLYk34Sp1SgAVdEIT5HdrjkTCJsmEbrZz8/1+xiUYHDnWBgP/sF/DDP9aZ+mu
Zr2RMZ2AypVHlc7cD2iHiTXmc7eVw4QXJ+JSm9+E2EBbsrbMBsVYqHU6bgeRdToz
BRm8XcgEJ4pEPk+zmhRzZks7Cp4Lrl6E0g3KEdBAw4gLo1E3vEpld/LIEL+KWMH/
aZgN+6fFg2+pObmtIFxWjAwkJciRlmvNy41eH3rmmBLKe9vP2desVxY8gb3C2jDF
styhKbhYpfot2PTvzT2lWaopgo5MSyQebYawRCbBEshYq7yEqFpIkeZpK0Xz1Iz9
Og+/hLNX4oyd0s+RMf7QT91yER15oJ7XEY5rf95qTJkHD4YbgGkj/X2tSLGeb4+v
sk6u4P8+t0J45pmBFYkONP/r8RAYuLzCoEzphafNVLqGOVK3D08fr4vNSr9X4xru
A6AIu3tHS0veCscJuFWKxWTrakaToJceqgDwuaxYISQNSD3Z9BxQNUn6jzEINHsT
ubasIp3BSNuKBq2w2Ke9vAkT4BUz+svEP904KJvPOfM6tlX6MM+xbiItd4EFX5SE
OPZgiC8luBjVASRWXMthAzPia5vW8Hdt0hS8hKtjdK1Tbn9L7vrCKiOjGML+lV6b
bTHigpD1sPZHtrj+d+WjW6E35efH/35QgjLGzVQVUblKb8eSLTv8EbtzymoUNWxX
xfM2nX85NXTZLP6JWA14/ulAlN3okpio2q6tlX4DdNwclKQkSrHz6fS7P4f4SAva
7L44WvSA/ijhPXLsPwHgMqVvIZXQs9d94BU2HxJ8HM1yDwGCfhpwwEiplZzckKhw
Y/xlB4dhy7BCpLhmAGkI6zqXjnb8mbVeZpzf06DN3qoVrJ7w+5ucH747QBMLZX+N
eLnzVCQmxJanHB4litGJS3iPThJPOKFaqG0CN4nZFBmjNYg6PyZHZN+zFj8rieAu
6kVVne4MPa4RuzzcLZnLudS3zMb2Rqi0DvFvuEsa3XqTYMMn+Zbn9nkkOpTsTeSn
ixfF6KbYuLI+x0mzbI7delA0yq5hMdyerGWgq5v/jnXu2Vq20/l1iGGtWbjJAXlu
q7YahW4VTgB0BFbYVDaaBSW9Dr0Ncf1vIxJmKZwK5zrqtMy06GCKfzHagw/WQZC9
28F54GIb84f4kjx0gI/bX1jQ3GUwnyhPKdACZjpN8p3Mc1Kr15/fvu0xyUU2QtvQ
wgIkJMQN7V/tuLZ2okSU6ok96XM0NV9R+scQINheUf4MpFqSKEx+UgU+47Q8gYqN
A6ufu6HEtqJN/xI5KrRDwdaK3ubj1DIHT/5o4CduRxQ9wfYkBhAlEQrOSfsAbJqO
MGEjiQAtdTTdI00y56dAb44BdHGQ4mlnF4hfxDrOVy33rCd1O/1pajt5fzfxz1S+
ptsM6rvsXgY4lARGXBCKOkzsJYnZ1s1EQbp1sG2b/bXTzOknIqt9hviNSg/lEtFr
xfesoNlOOCYsEPAo14w6+KaXrZy2aCt4xaWbsV4QAFCF6DL7a0F7PL2SQYFpUz+L
h1QZ7aALTC98YI6hBvun8Mhb6zesaBAfhMDjeK8LXrSyjrRAJt+9kbcgqyw7zfBh
u0cMjs8FFbbtAFHqkfGAWJsTl44Rp+/x5ASl9QJbyIHrt5bwM+FtZFmq3vN/3a6X
7TXp41IlGmBLtBNjANhwsAQyJaw+//p1yzq6p9KoyQUzMdFhiU5SvBtb1AqJACna
Z+bdX12TrO23zdvL1raBaZcYYfGLBbHTqVd2SGjRR/vcTDuoJEmJayj2VXH1H+NH
8hHlPkxTANO1chtvDr33vgWEfi97z20nbcDXai0Vclit+CXnCWbUp0V6EkfDBuWr
sYNUvjWHYehXw7ChEVLMHhm3G7S9+yuKifCYN7xN4cS9NU0l3Pv56q2OjnHsFvBP
sc7x4+O06Br7vAgs21DIBttSS1NzeC6P/fDHeA/nEy/mhVceu22XVYBDSjNVoHDA
Y/FduZoV9h42bx+/VbiAbG/SUogwJBjf1ULlRnMlsVxQQqzrCCZ81t/WrbK0z91o
mk4s4bYw5wv8z3svQDbpbr4mUFtSjrJrKmeY2SyCdGTEK23oFNBawljLOcrQrqBY
X1+qJimobxnVqWBKt67ojU1EzRIxHQtw/rKsOy8UC3Aq9GL1qX/mFQbs3eYznYn4
kN1NDj7JjhZwXPHuqzfPD+QX/1Hn++4TJB8B4h9qWUne3UunphYm6Hu4ZUEcfmcs
p2f2xkULYmzDQM9CYSICjWhpuJKKYp8z1jOu1SyS4PLyJXecszS6aTTWNNMigeDx
y8TiuoeX38EkIFsjy6NyW4mB7sTr8p4GRFQ+FiokxBtN6AsLQC5ovUV34L/4n3HA
13lb02w1BJlpVr9HuMgvJ8NfNMH9zphexoSPSDPH4X6oytcmcQM9V2OQOHqRjSVA
MtFa+yaXZsdXXxN2G2ZQaudraSQ+F9OR29vwEDHC1vdjw78bc9me5nwOX3aE3BIu
dSb6U5qRC/0jclhQ8vxnGOpoMtW2WpPycOJ70zAOlLSXS6IWuRYoQJP1UkOBa9oH
lo4V+KwvSODPK8jNpe+/pzwmuiwzaT/J3urHqK96lmBfx7ZhsB8uYSjX0J93g18m
mhFUBeiyL2Rc/AOQXLCXfQzY7mkpqLfPTZihR9zc7CkBj1AxoSk8oBz+ZvzqS2Wc
ecRMpdimg85uvDL2W3tZLQwx6DWktJSsRpE2Q3DwPquXd/gpbD2KXgj5voOrysEL
r9kIeipA3B+VTillozdt13ElQUH3ZqbgIH26sAlnomzXSBk/3fu/CWmxkQiLEK1P
Yw5E70S3MhCvL4LyjTNbAH3L2kyG9hFktD/1rdawMnPRNOT/CJnjVnzfuDJfoAHv
ZiFta2aD9khOBiPAAH0k4Z9hcfy0DhE9abc2fOcDf7Vn6Z8sIUi4jEDaxqtgMH5Z
NIa4k8WtK7eDW39T3ZMPG3WWAWcRH6TvXSDrmyLT4gHIySTXvegg8h+nLQa7n9tp
aGj1g/sLQfuH0RgEo/d8ZvBgkBN2iAeFYWobRCqUaMFqvkau8rpr8eXg6N1LIdsx
H/yd4G1lYwVRQ7fe8dBTlFPAa1jT8oIw9cqj3JfGxXvnYRTS8I7z0EU84QguyH+r
S4EZmmknTfwEKZhf3apj6fzwf4/Dob7RM36caeXVRTV4NauW4rBkPEFJN7OCUloM
tBVXo9ROXPyn2UD3NUXbU+LLV9IgPaLNFfQV/KJPqBvXQB7tL2qNf0EoeMgmZu7k
wSOASWUE9HhnVWg4neDg95+rM6h1f3qDeIMoQArjB4rnrDE0/hJ/uNxkDY96GlPt
uE4SHxw97507QS+nTNxLN35xXJoR5WSfGuLCms8W5ufKPYasQ7UHBegmSDThaTe3
T/bpX9Q72W7r2mUJBn4X+PIUADyWZZ3rMpSIc0sgaNuPg0sAEuKKf4K4TtTVjnzJ
CGrMzLM0OCZ14su+B4KzT7h8rJqF4R9SQxPZ+paO31v3xCNxbXETsBzO/jPxIq79
VQnaAI5o+QwbrEWZIy1+XU9ao0m2H8ATAkRf4FEJFIV0OgdibPq8ALLNZyoyBVhS
atYtO8lVJqs9g9E/ADPf4kIygBYNTtIdZe+/SXwJkv6PTUd3ACKqjlKsGttc7ICE
CY1375N5Az61jNSBWJ/p+U8NkyqgIVT7zilrRxrUZQs7f+5ZmV8Ftblzs61wBedY
zQUfA39mx4ehd6l5hk3yJVJgWZhBv1Ivy+7SGslm383TWM792yfYiqWe6eNF8Iqd
Ie1Ptrp8y5BYJBnOUS2JsnhDEf2jkuI7L6heiR/6LnxhppsN2vuwkP/yfATjYQLA
Ejn6jvNMQB1l4dKYhw5a6KNqUsr2JNLVBm7X0fQymFJmkzt1YVvtXJjbDxNzqgfv
dHnPjP3Of76ztq95o5xloeCBBo3YzmMQ0fLYUgbs7DKqWeUZkekock/JVO0mJWYu
wUpCj5+fpTxnDNzTveW/mEbzRwkheufiix5uqMN+1EWqKn7ALxNp04mrkgwwuVI6
txQWoVoY0dqanwZRwJAwZjQteYl+ZBcGSz7hfWrP9oC2HX4HWOu0mKh4uMS1sIYT
2cD5IB0fH9lZkyfJ+jwyDZTALI3ji7fyoKJTAh8klX2/+mF8DEX0UiOMPB0siN2F
K9GNl6ksi3ROYbCy41hJ7GaT+gHxmMJYaG+ZmvM9mOUq8Jw/yM9ToO9nuDu0ILT7
YOn/7mx1CEkMDXlDCmMfTp1n1O7MMmSmufpP5zxCUXuzLJwuspGsPtUoxHXwCDO+
KOtyYgE7T9BPL12C4bC04z9UkjBJlL0Akg7UCfoFppG3ZJOw2c7KpchrdH7mDLCM
9z55UdbN0o8IE/w+EmcJHEOA4vTQxJbmsw9bvZ9aLE+OFs0X6QsPweIPHbWGQ5xh
sxwZ89eeXKhfyIEADmCn7jld9VVmcil16Gm2l9Wo/hEYAb17g0SY99qqWsU5X+9U
W9EVU3KwsNSfBiNURIFc80UvFyH06NEYOu/NmUIaSekFJroSdbcUDtEgk0fo/8Z5
XXzWvmSC1Hh1fxyL+2HeaxT5sBmfQqoiUdKwZkMcT/cdHKTIcbvqCIOVG/vxYZ0i
HprMnCMVoNTp28UImbZg4NYypM2aArnOpQCkIKieNMy/2EHDoTMvjxo3NpHtSvAa
ety2ebA1EtSF2DozFF5Y7SYNKQVzZQO1gwYnhdsKVqDG20MmH2mmhSbCsU+ExRp9
3+raEcPwVfZ2aaOfNWCchN8zIrQjyKTRrBIOeNorxtYe0MI8CazJzg88i7oDzF5F
I+rdbt6MLBzJR2GIDV2cSYePMv0JtblcccXXdqxtWdyNsR5/kS5C2tmaHk1Ga/Vq
Y+nPJNvju9xs0Zq0XBAghfhMaoC83bKdXc3yyYisrcdDPNdi2LmcdEt6jRZi5iCP
DTNlYbIyQoaTWEb35HMiEBVUsy7b7rBFgX1GH3D2JOR6DwVL7ZjBNSYmSEi945Cw
DXfqUzWAzF0VFjDAktYaQe6yLfTqjF+lx62NJ6c6hYFTptn/omRiCGgy/8SISbu8
Kaic2PE3LptFvgJlU/sHQLiF8McNUVpbt9NNNfSBWTBJCWh+UIlRq/Sn6p8O+k+U
pJqOQPXL0ds020aMoCgUM04oP4GRRdozc7wfptvJZpVnsvmToh2iFpbGKPU4TgYx
bn38UCjqNx9O3F6Vy3Yrfsd0Uq6oEkSFdrkofY8Gml2nF8zM7h1ZZJkiNGXcO/wR
kzovKZs29jFjbwl2rUebNv1NLbKSfRWXf1YPHzG5HWxoUkHDVafIvY86r8rib1Nb
TkE5RRBe7GJzWXJLN5BNU2d2a3kUhx3hi8T57Z7E1hztRCwFnrx1O5vd8vWL3OOI
EnhXZ3QExKDbyLNk4Z3hk3jZVGNkGV+QS+JWiVPJwhGxfUh52LjKT8W8fLmr0yhv
KpE+tcHJ+lRkI0ePsmdh+sE7OvLESxmZKnYxk6jqDIxGfxk4zeInblyI6MRGUYpW
pXgBJ5CRJBV94ml/mkftcueTDsephlU6CUzGljcS3ZP3j83XXoNeaMrGlTUhnIMm
Svr+tXfWcY7CMEaCTma4Ef27AxB6obZS86lA9DrAfaSQ+8F5f5gWkbihBBRq0T8W
7NStNv3HYOzPaSeUVbx3TmpSwOqcklOYADL17xQbvGZFgZIUtQIsY7on8eeWYhOW
RjLJj4gzwmM8HmSgTPY037wBCFwxhVfMne+yhjNGurQrsOQ6AywqQZtx32ri8jlX
mHyj8GiexwpSaHl/QwwWFqSs/H2FOQ8hxy0NaozfOXuV52AsTxJIQENybgQeAeiN
RqmcDhnN1EcvbPJE0E9+rTnfU6BWH96h7iypU0PYZHjSlTVkTtRdCc6ns6um4XUc
5WilghyLz9cpm3L+xLAG0eVuiwpfO9NnsvvcY+Ht0HdQGaE5CbXL37lOqUhsgZLa
dT3Ae15ze+IkN2WFwVbngWTnfPUkhWp1RHzS/5GSDnzGE8IdTrpa43s96RlYt19o
lOPJLjtX2nRtSwAPbNMRpolYMTXHs6+kfgaFAqjcYWSq41fIiQ+DEvpeVGqtT9tK
yAzACUzotZqpYCBkeFT/3oezAvxSgivPTYRXFegFhWlYfAJlgvfJ/izWezNnT2mN
EjOg+ZQdfCpVvWIG9jucZoBv4g5Fe7j1ljf8VALiqt3OFQw7+o7nwgo31ggBWitM
HyU4/fLo1vCb9Wm/VvJAvHM/hx4gJeQoh9RdnH6xaJeMDOn0qCDA5kUv5k3uNvsh
8K2fm8oh2iqRTK/l2SoByEP1lAiJrMANjFG+K9YURBZG9J5QU7pWYp9AFowz0d4F
RctkW8T29YBRjlasiXsexUNw534gVACqDZxkVbBc/V1YmUTxoYZoJYGyHgruSR2G
PbrmTrgI0LHn8cZXmWmWfu6jDK3RHguMEN8sVsDe/Qy5tht5l/2oxS+C6LianDwz
j/DXgSFaxUBxL0zL+GSblPe5axXiPJNJGtTyg979WCKmH0/AqChehLAU/OmitCdZ
agPgfY2hg0o3fiite1tRiq28qQfbG7Cuge5u96QBKnOlua4vqvr27M2qwMaT2e3I
eTrjvop6zBo5aG8jG0CuorkEr+7sMWlUC+9HRxeO5YiuiNYO/T3ya9rH+DHwPV3i
upGaItf6RLANoel27tmZ6RlkxVK+zbJuQm/co/D+IOfZGy44oBVHfxyIVNGhv3Zw
wtipT24bfCMizkIx+t52F/eGe2P0H1gVeigiQ0fVjO5YTwANJr55MLr1wf1UgXda
/1aBW+Pfec3I8rxg7dOtEUCchvCyOM1c5iGCU/bBzg1HTAE82vfvWBNVdqunFG2G
mm11be/T5xRoAjbdqq6FPpfnFlnRr2knUtIcXtrDGisg/p7WII9ihVaUyQOwHj0v
edyMDZSSfDpqYRy56j+4ua6MtZ4NP1ukuoWRfpzzWwz23LyPiIhdjb3B0gH4EKLq
tL0lkuTnvCEf64rdAs8ru+4U9YH/Eox4egzKogm5daKSPUbkjl/rq4t8h8H25LQ5
1Xr8eQbQkm3vVqqulPNEZphweJiMfCugmxdHNF/ivpP0yucpF/cRn1oQSvG9kM/7
ObCu68qw9C2SrbsVKjCyNh2HRDcmg3VwBt5qUtgaTi9x88KvzCVGaLvPI1ITT5bJ
KHDBeD0ekYI2qhk2KPb425vBA/LRBLNcxL0KQ5uJX4jW84/Tos4Sd+Vz1HpIZDXc
UoQC8V0vpPnxllpOq97YYg7QNEi8XPE8hCAl6cvUPBvsdQXV6HCXj7tj7+QCJ09c
aXQH8O6oGotK6ZEyH0tl80nj5mXU6hLuG0FwgyKe4gFuprQgUw+KMQaICafLE75a
sLnMJ0kI0ah890O5Pgjx3k9VE7CDzlRwlq5H2Uy7Nj+5Q//zM+et4OQbbKB0YsRe
CgJwP0i+fbmOegJUtaHL7qO6Zjpn/rteDlByJwvemCxNNFg0gdReIZHf4tJoByZW
soDccvZJbptxJA+DadrNV7msQYbiHxRMqsYX/3MlWUO3i069fkjOd+KaLCK6byYT
ao2z5KiwtRRRMrsuvTfWgFPD43i+dvHWWk/0NhccFJdpcC9yA/sOyNmXMvdL8Lxq
gwhwReek9gUvb/36CaRrdeCWn2hK6hG/C2ZYZc81UG+S+FJVek8NnBZDKCFGd/P1
f2ELXW1rNuBSrZWpdupSc2aKHfrB4vXZmiMrpRj6og+znK9V74ZH4mdCUDr3jPww
JUHQExFoTb+HNs1c3RRRbvt2MexKZkWRE6tLoU/rNCKxzSoS4B1dkAR+waJsWEY7
qDt3iWMtI19H+8WJi66nmcrEYzm9/toEE+foFKQysk7j6hiEB5H71xfa53JboqdX
q9UUdANrGLH1glWKxJe5LwXZvpBciPwjNbrCalKYxMFK9giT7RokljKk8Es+vk51
BCvuqJeiU+AibfRadx2YCFQYgqMoXqHSh8HZdItY6B4Sk5S8VFzTcoKFYwxyJfNP
ga9z29OAiTRCzFld0XNeVY86QmtZKmZYB9yLQC9JosOEJtR7fd0Ny5KYF9TcgBHv
44Iu7CaSoYWud4ekXR5wodNTWde0Fk85fLyuPf9Bt/UJ4Z6+J+B7wYg9fhGsvy2v
mDMEmp5lyGeN0qy1DZsbXW0rJo5+L1Jdn+h06hdfCyGI8C2dUq/ZEPvg6JyIJviG
3CGYrVunQtWC4w/4LsARsmrNFJGMG12sbBuaAtP0LNUytLcgv3c1OEQYg0mzMdbD
DV9HLSIDikyy0u/GK3jw4/rQ4roMUPGDjeI9LN2gaY5XAyQEUJqfSFUOQSc2elTv
QlP1MWk3L7pE6O9Dq3vVIjYe1QWAX0BNXrA8CjLrv4qqGn3HSjQ2cqv53EtevD8v
t02U0B18gPL9ggrs1rJ1OLXrjimbz+Q1zElH39S0gnJtJCe8U91bf41zviZ6Ml83
Dpq5ufUG0S8pl+UF9ruGnRAXe3AySg56DOq2SxnBb54Q0cuzACC88SxrtgKkoWj4
YeXm4+XRhgG4t8GJfienqYmy1esVhyYlWuHVqtCbno7v7DnFvJ00vG+FCexb5Jnx
ePL5f1NHxZK/ZwV7dLlWwjbJOYrj9Edf7QaDgBwnZryNJrXBWVP5Fkkq2Lhh5j6d
aUgUS3IAUPc6GZ/z/XleaJ3p3k3pQsVYRdwH8A3tZ0SoPyG58H7jDqABmZlBDTSv
17p7lP8/qMGFE9XyboiHkKCbqYuEJSvKQxLTIcI36VH4Vc3A7t3ChWT0Hft+J2h7
dMDrIh6TftnYmyVU68wGwWGzuwvmnkieIvCE/0sCHXC1jxhkWrSoeQVi0ullDLR8
KahJ2L6NXFGdfyC8nUCw1VsigBNGLMRbNAzRI2U0DKc3XXox0GjBUOX/KomMYDoG
X/KYZD2hbP5K2TYvnc6I+qG+jmwThgZaFUgDPnbCE+MTm3mUYpoRvH5rfaDDKsKB
PF18YIiFC/bnhM2LK1ABPcjejD75csl2HNpZ6HsbPO0dd0WD/qgl0NpViLpqxU3s
jQXducuxqgnOZ2jjEUDF+3jGXmvg8+XbDf7ZRmcksP7yD1irEhbvLLhFSz+ByYkb
9NIcPQH0jgaJWunZfNjwt+d9dTQsNAWDl6cU2BtZulaqKN8Qoo0tvcArHo9azTGp
pzSUAADsj4wYAfDJQfPtY4QRfyg11D6PsrYl8VSx0I+of2h4QMUWXeHxQwgdcOI0
2V3FFTUhW+VIHBQlKSzGsCqedOUQdHybCy/8M7FYurQUrCmyBc4NiRb0Sq7YIHS/
hl2O12Yy7Snd2WVSHxGh/oTU4ITZbcfxqzN1/HBb270WQngNYmP1Tfdt/Y70IJc+
w7DKO2kAJz6WXhXQhxcqfk7wV6wMoJZubuy723Bwjx5FJhzDuJLj2K/hMA10qsPf
npixtlykmnoXZeidtOOXsVOZ961PQs0s3faRTblj4WUs6lWv/MJLckHKdUJaEPQ4
S3TQ/Js1T1PMABHFTDb9xnfJ6IVDt/vVJYRTQvQtgrPpp5lcVhmAjRp4+kcziynA
l7I3NXNoGrTCQN7eFvu5vxwuBmnYEJnN+APCDgirWs9IQxu5yYV7v6ybt/6uebiD
FQ+wTJ4Vm6b+vkdOQ6qxdG/nJP8aFX5amYv0RIOjhctrsn/IxyYSDfHMadEz3GKm
SvuoAEypCi7fs2HO+AXGlKMNe5B8+moTV2DP/IkKDFIVfRSYUuARDZR4R1vrs+mt
wCWJ6OBTrozQlUSbykdsaO3yd2CKgCHUiBQ6Ig0C4rH9nnKFYpDvG6HRojav8cKX
+x1jWa0T4ju8zB8h/DtYMkDcC5sdDAoaYypbBZUDMBSd4KO3NXSLsoOuZnYva033
KX26OtBAtMxJ2WfxhfLtXXksgoFHFwmYx6tpd/3ZpitoRPfIFTPK7A9qLTL7wN/E
J0GxquvhuEBLykEpSpdZuTFeKMFzQXOlxYwB4I+bsNtnvR9nqhpoqNZLgokWtzMF
uDZFK7PuiZXHPdpoJzYzOn7FLSAPhR6B/NchRJsWVE7hce5k1fuQwieDLk24Bv2l
g0dKmpjbGqRIHhvx5U4k6bJjWI9Ah9GJBPrR5N98hP4l+YuDIYNde6uL8yqHuznQ
b6mu9POglMzgeqXMuSZ5h3HLRNlfgJtv8Y3eeR9Ry6tpEftkRPx75P9WqyZs4TCG
XC6RrQxPHqKcGYGufugH6dw7/f3Cvs3zCANOB9kSu+cX5nNvRWsKjfPYBoCF6RV7
QoXPzFYDLIWakYwjHs9ulqrEuRUkpEzvFqKDrrDMKkTHNqDE5sOpx0lmaj9OHG6C
Ga0P3gO1CGyGwuxXMqEYUunBni2oBMI8tUGI56bGp4IcletNYDbIHKqMcwZdAbBa
zrof8BpupzICx7tfySTmIf2ZdkQwYU6vUWax3uuVnJMQRX3avTI0Zof+Moduk/gk
HKw7xUsr6dNNjwCEdRYrp3skJpMN1LoEeXBzE0o54vuBLk9ecHM833WVCpECzY5g
O2oxG0jnAyRlWxDyNLYoCMzP7MkZHrT2oJ3o7U2eIDY/1zWF49zKSV3D/BjHdtni
YCVg+J+e8Fq89OfF4VZF0mr+nHkcWHgkV4qw+RGfTE88Pbw1MVCuVPGrKd9bD8AV
55jlBXSyZ4msRSQiKZy+PYb71HsBbioxiqsrhKRlBCenftio7WZKq/SciK2HgKVi
h4JntZTMTXG85y4jnEYMABgsfe1lJ1C4surg7vuN66SyU6GlLvwGNT6ctIU3GzVX
S2xUMup/4VEddcTNZO8DTVTJ+tPsdE8+TJSFsx0zft7jHEcAENEiBX6OJbpKwOPD
3FSGSlX80LkMxVswoPK6CPCVoRUz/hJm0HnexLV3/a6iEuPlC4M+Em3AJ03KQ5SS
tvkz5pQ8QKpQFebfzPGaV5UzEsf9b8kuwEubxc3qs8BsVfnb9OlrxPfEMdSWlW+y
CviAzh7oVw3n9UtXI8o9ldVOsVOzECFZUFKAKVs8ZygH+KbpIURfvD7rENt/i1yq
IXvZCEFBkd6xjbjNNlv5J134RbLhe19NCOVDAd3fCXNoSmb1DHk5PY1Juc9k7BC8
w01CEt04490V5mRCQGeX9u7sdfIVSoRaQt4jVlc34fU5zWpHLF8scIgLwTSSd8jL
Zxq0ANR29olx6cWHQKJrzb1DkzeM6jHkzxWXxhjrC17H5wIJoWDoQXYZpk0Fc5S5
7DyLa7up7n29pBsR+iX8orPLLXXDNgeRc4MPGBGAQrr4PBggpoSo8GYp9xm/vyEa
gQ8JpKkCFc0h8POeefKW4ZrCs6I5wS8QM0ep7JIioeWfDLyeU64EMGoRrjpPtt6y
qwitgHp7pd0jfjBxtSqZCn52gWROOUqx3b6wReBXPk4bxoqU5OF7M2QB0YfYbPtX
qpGL7ib/e/SLAz0m9abBleoQmX/QdeitHMdPpnfmm5m3mGp8Ij6kNIuWiidjKr0e
pF3z9UljQgLEto8124+0VtOworK61/vTskQQAYxwYLBRK3lqETQpV69EfGQz13dU
wzK3n3vmW8aqT0k7Q1x+P+CRUToRpCSUHBrvLAkMikMIFBc9bwwnNkqoHPWxgsO8
qfQs792GhMgDFp/NDZXaMt5kXZBkTtiNuz+6WS2wQWPwHEXkU6KPu9stiNHpdEi3
yo7zBSQjKTtvodJAyrJYCry1h8OiGqa98H2zZO7oqMXKgl105Wl5UJ0l+WqGnk2x
vJSfvjhpEM0WxOKzzxGLGbm4wQvxyPyMePcjNkKeHmwTsuYLFwMmn9YArQ5sL4M2
BSfEsKQ5dV5n6oKEzToyaP67c+pnaaMF28KBE8uEDlh1aYpULZJ/Q0kGdeJIa9DM
u6eVEQdLmR6nRzL4rRfrgt7NQj45FXA6Vgh0jzHr01r/x6w+hXVXibsJy0U1hXde
t97QBGNvOCd3E7tPp0WmxJkrslOyEe3BSjlQBGirEYfuZRKBIgy4S4HkircSgnEX
FTwkWaxQ4OLIHbBd7L/Q9Mxmk0TeAzW8n6VOUL/sjjr0Ha1wuYh/VqDVbNAhInMf
nvQQSpHAs8JXs3LDzPGq9QJViIvJeAZ4V7wp+DqlCX6rU8nxIFVGvRHsC5RMnV2s
hI9FhZhQjCY5vaR2jrExz1mntMOvneGrpoZXXMWhhvHtTeDD6ovjaX+dNgFPUm1h
B1OXJ2SKvh9L/A8AXDirunDh8/JZRBo1UTJp3x1WbHtbtPIvuWh3/dNW7O+zs9Um
PtXU4/1r7YRkmt3Q/QbknCaekbQJNZkupyw+ylVGrYo0x9R2HdWzjlfKL5wqaAqh
sPprN3FqqxeMH7bGdbzVFeE//DMg09wtrbaF7tOOV6I74Olf2fQ+HduoSA1xl9dX
mj3gw0B2JAVeEdh/lfT0/HPuah+AXiKqD4DfVGnHFnMrGr8CXkMIo2dwqtb/1sEW
ljdF6ulAWRwIZGyBZ+jtGp5Lw9k/zn/AMCYfQIrF3yJhz7Nid7kGIz8p6m1OIlSP
BIZo78J5HyGoScjDsVpgwFhg6HaZxvHe+zfw864NkQGsgF2mx/ZC8MQeAwwqsJis
PsH+TWchtDI27geyX/egsA8zIbKGxl1PwAmzdRA1Pd+xUUUs7tGOiPaZNGt5/+kb
u1NEMXW+KSkCp3MjUZS2VvtEpY+iOafRNyEBfijX6NEnVbJmyyXBkaHZDb0A0NDO
f5cSc53tI+GjiypPvskxqMwJNx1MNyvgBirQ3zHPSiWvn92cONN+1biFeFs4kt+J
hhRig+m4o0JZTznjJnveMwctv75e43f7uuNFWKAQPnsTBP/YbgxYurFnjv/Wv/N/
mm+PkpVMJfQCPZGK+w4xoVGpDq9+bv63rtq01n6xSzEIFw+5iPUO7LHTwneSt2/S
dPakLzonXver1aEY7u96OIRcpPOwbhcEuZcVJa9YTShEiHdJB+ua6EhhKKwkd63M
JJ5H51Acv8ekFt2c1DYBMOETR5ayT3xTwOAGVlXfTf5oWK2nfB/GN9XMUaBXhPx4
EhI7haHB8tOOUujbAFQCvWLd9OyjkLeKrW44VOkhpbqleyfKO4nl9p64b3QjYHSe
4amvCJLCIOwUA4OkNpRc0evbcy6B5v4AWIalJw+2qk833fp2bd0b99zQNCvJYM1/
d5+SbNc5PIwxNviMFsB1TbnYAEa+LC2gfbaudzSQ7oKCdmgYYvPgMXgPCGy8JxTf
Gd9guPRRRrMUxO9W1c1XUnXe7eZJs2R03fa540IxI4G+2RO9OPL5JacuPeXmXrQC
upPZcsxQgz2O81Qd3KLSHDUhwJVIrLRihzUj3iXl3bBIofIo+9njoewodejYrsU3
4cUpfcgUzR/kFPTUHfuyZ7m8ETyLn9PXj6mkjA6gBUKQA7AlufrmrETziQFbVi9j
vMK9kcEB4UapiBrtIsBqwX3TAu46rMNAm9d9SM2pJpROOc2z3fXkN4wrmtrviRUG
jJ5AhtAG4RhPUJY8gDox83RSf55QoEBL6htCX8/kICSut4WrbJLuDGeQ8srGtppq
p/0SX7lhPuMMEIBbRF38bihRKJuHbOhNnsOPHXAzSK2QDTUhDhHwXtqpTScls7Qu
k0zi7Bwquq+Xa8WLBDfUGuQ/h/Fy8/ZpauzEz3PzxrOB1tm6TwhoX6NedEQAORC2
Pk4/QOT+xv4MeQEYsIN+j5tE5aag38XqPXQ0BfCue3MiuNtjn9HrkwHmGQqa8m44
O/19s1kMnLL84Vl43NifRsHuaN9n5+PX9e8mG0oXMvHbu76pzJRA3S4VSwKe0cn6
JWG/dch6Rb9xXv1yAjpYXzwC4gVVVBV/MeRcJIrKNNJp66VUvqAkYE7AHhk8+PV7
4Hvgp8bOWgfHSLjbjRCuXScsVIcPrpzD1BiGt06Nr/nX10rmHvKvGjMZffIkQQJm
kxcHEkvIbjJZMaTGLCo2NSwpFZ1sEAqCp9NNRiEk3XAKtqwcuU9zbaKTkP09DUGL
bVda0Zm2WO0jN9A51uqlDtY2rvQiiAx8jd9V6NikePL5mSGdqY+vn3McwOCgJvwW
8atyNXAxkyV2/NcdW3AVH8vGUmRbmxLvuoT+nZEUKt6iespaJx3nWwdxo1MX3Ssl
PIoGjJHo0JJEPy+3+k5Wdr+euPfoLNwwWsfdWZ6tSKG8W7MtQPQFF/A7PtrRDmR6
q7H5dF7Jxte2GwA5MGioq4Ldoe17aE585MbKq/Ygs6AzVyJ2gwLulQW0s7AONccV
G1sFHhUlGegeIUtNzaBQ2dw+5zAGrWd/WeFHNrW+7Zm+Pr02AV84ODCE97etX74c
DtxAQgCGGQ8WPHfDcfKUJbyMNdHRRkYau3tmhlt41jkB1j4o7juz6oPscOqdwjaZ
3mWI8ll90fy49F/yK+zebV3n+y4WPQRSuvaHKjmWwWkfV5dhNv1eQ/z0+YYpHKbI
DbEa4jsqeGWw8abrzyVEdIly2qBmLneeznDZYRs9VLhyG/FOFRVxZz78MgzJWE+H
2ZZeWtosIH0c8plEACPNAeivLIuYB/0+yhvGtcv9mS3F9OGUTb6tHuH7nlyse23V
niQvmJZN6LM2Lfg9mryGtlv0GCyfTC6scYCpOWVGKgwQ05ES1NclsgkrtkSiAtbJ
xlftHPaMzAV+/lwH5cTztsaZP9vzueb5/ng/SYjVxWBIoallMMBiobVSB7DZvF7E
7oCXc33tsME0DzCz+PJf3dri0h/3GWT65hyIoE0X0mPf3XKXqJ7PJf4JZDB9m/6o
SbUz27ZzKvo6XHW/HZSQwSAXLPqoVrM+zZjvv4iFM3w7YYsuKjXsdm2luByNKWNM
6eYnH4Grsm3ut+Gy1+h5NZPm7Cn9b/AMb++TF461zWRkU0CwVXZHFPAf4peMuj0j
dJfRx5MDCpS9NjXXuF5tjqyZkdYH8OrQ4C1PxTfvbhu77VHgfCq4OFakvWfVIII0
uEa9F43ud2Xu8WmrMnvJ5PcKdUQBBlaAhx7MJiH1KZ5ScW3YxkNECFRY9Bu7VbuG
ithow7CoU4twTyeR+d3U5XsEKb/1IdB3/DyBOoT/97LK080i9gWWxuVpumm7m3Ok
dhYfrobs+zNfsaGW1QJuNNIkbznVi143+1zBgJBRFvfbD9sHrX9hFOUUddMhTOv0
LvOnTFX0LgMSdD9EYra4cwZuMU6AZMIDQ+hf6L6yuiEy+9qZJHJa9fR3bdSbqYTP
i5H9mLr1BcMEhS3jqc5pIY932PevfF35iukwM1jPPApUoGVpIIDGd8Q8vstH+W2G
bHoDP8etKET1lK1Zbv/YfKFhzxV9oDSeWiCjv+0Xs5sF6lwbzXW4t7sTNa6Tl2WN
3Yr3+Ss3rBtb3I6eCPDy/IrThDHN34m9iopGZUiRJDkSpGn3AIXBIZ0JKVYO9fNe
6NPv2nVO+yWcTLpok30Sp3e34nJZZDOl1MWy/DsipP4uAbxK7EQcaJUsCX77wjLO
uxo7Y71ztXX7iJy5h08xii+Fun8udIXE1qR1f1cuLY156uQuvNvxR57/Flwws8pJ
6mC2H6BLMOF/LaA/SbLb0ZXgLbLagvlq6c9iQn7O28xkkbad3Hq4qdNikk24uAqQ
Pp1J75pI+BdKrCk4SwqI3nXVWLa22TgpVsC0cmlM01OwZ34jmy0tNIRDSxEKc2Wp
XSPPHBuiEJtRoRqDiTdHwBquvHvM+tkawA4iYnFVeQfGwIeH+6tdUVfErODyMmjK
GblgBKKNmAk7LC4SQrQmGW/5FZrsYu6nfUwTljM3WRIK6fbk9XllZYI/DcW67u4a
78KIj8zwAEDjp662HJ8HIOol0IuE2SVQN3Oez3JiCAv/VhEJHXv8oqRmYdt/8Gle
W7hb+99x0kS/4bdNFqdRFoORA4EbuglWXuZ90sZedYNRNUrChdvZHFVUCYSMNIH/
iwowKuxPaCtl1B0PaHgAqqN1Gc394Av5eiRNrF4ShAUhKpIg4CP6iiWbjglemqAN
rJzNN+bY4VKycq/mZLVj5VHrv5gB/qjJGVql2Di3tHgPHvdbE6iSeCTxkiUPN86f
FowyWUaob+JrsnEQWS/eHj2zzOyKtuxbg/kuWB8HqSOCf0yrTU5W1SaUOpxwxK/L
hYlBzo7RlxGOhxJXiGIKHu7qamP4UugxfUsVlzmG0uNLp0TR7rpcRephxxiig4Ky
fd9VCo/DOb3gt7rX2WhgnsJ+TkKOOWkUpaIi/xghl8BXidB+fgc9ScjVy+T3zGOT
MRFQJnZ+St+8aDgUAh+PdIFgynSRugtmlQDuSdFYtw6sAtrrEpNbExp47xGgCkdj
tnkVio0pUiRqUDIMdzVhB3J1jbAY5SW2xsUHK5uR0RG83Gel+V24nfh1l6coe7ew
Fhq8LSDzPW0o0pLz22CE9zvU88643yqgJ+Hax8foXcWxr2yRsph0L8UbTPl5vN5g
pqU9P9fXdBprTkG5/q9STRr2hmSn9h/t52m2DMzbSwkD6n5FMh2ksOEJSLBLAqUn
ssGPMHoxkE3OU6MsgeIyQ9Q+MsMMsv1VrWNyKwAJnb9iMOle1oZ6TuqoG2pDxKQO
iverk61S118IIKYzbesaWZpeZYqfj8+ojF47T/UbOFWUBHaJFCq0BkKWnTA9gJhw
qUzG+TvYoH55yA+vgc0cands2updA3DO0ZCtkh7sNozXb99y2Hdbzq3zc4DSmks+
wkAxa9FYjCeCqdNUusfc4Kom69HNPVhxaoKNqT1zAyIkJpQJcPdWxS53IgHZN9I5
TlpmW0DR6WpdCPN6nYqaLKT3nHHr8FZ8saFPNd62J2j8L5XaWKEHZtSD8X8AzYJe
Nu4ytNlsTvfEVdYbeWIMS4/lHWSrRYC3PFDi2aHknbblHeBJ6lprKD3HCXAYDXqQ
xwfAWV+bAozwiGnesEZLX07Y9kPyjXuBiIFAOXsN8DSzcAZM3+E1sspAxfP/iV+e
74yaPkrRVy3da7cMZoQPZzv79zqXCfhmNa0Uy+wi3MgZBEMOm1sTMQx0A4lwWXV0
U4Y1Jc85Y9BiwMa6pVzIFA8L1biGs7LJ6lqof7IA/xvm+iNa1YE92wLcpezspOZy
1YlvCjwuSMAy0Wxp1ncdynqmQs+S+PJ6IlpZo6DUCoZSOYEYmfyBP2KV0BdAMkGj
5eA2347Pvg2ba0Y0MgZPv8PSfHvXuSa3ukjncG2Ud/S/yD9bptLeYPujeOWaUIUu
xlcBor7M6un7Lif/IFCw5rVRJSEiTd6fP7TsCvXf0aVJc2f4/03BPHQvpqyRHiMF
Kg1AIH7dsei9Lq1Z5NJ2+GX46SHxOqcKdg2vjAWNQ7xqC9X9Q7jEB4Eyi0NOEzJm
ADWXz6kKkAAYU6fvitCiYo1hPUgPKJkXIHKCD+JwwWdvF3vXlIhMgA6cVOKJK2M+
3y+f49EtMFypFlXQcsmp0eqkxoL1xSoBJjDLnrWaMEZl/jTPLv3QjMi8XKdilNAx
sP+GO/32J3jIWVWzPtagMijW1KGEj8UJTCmDSHwpk771p3tUQnjelkejXcQbLa/6
1BctjKhm3C+lHmtAANb5RuIQ8w0ek8m/T+3vQZwKjBG6/e0J62zVlKhp1TerGb36
zJockodhqu6pgU+//ajl/gMbXG+wuhyLYsou+2kGzcAmHag+e1+K9dXXRtIfdZ2W
i7ak00ZnY2yiCY+twN8nHrnw1qpUhKpKJic3rEM+NGA35ID2jwebqv8j2wyOD1Vd
Wm/Ui7b2BQeRbX9n0eS9blNpcliPTfU4ZnOzwSkYSnc7lcmQJJSwSz3/kmobp+uS
JGvDAZZdXLb/joarr7h2OBCsSWluJt8arwjKv9Inh+iVT1cqNOeQM2ix/p23HgBh
SjrOPmQp4MNhtY88y8NjNCqqlLjIXqSBVXOyF3jo6dJ18xkQoVifrsJpqIzquUjZ
P9xf8qwXVQqyXmQ29GIvQv+nm0WM7yveDSua9qpdE+IW/0bC9ISsCwnQdALl0Agl
pVWIQrLqpBg3GUUYvSpWlD86Q56rtK/BIRM400L7+leQlby/P/R5Hbk7H45tg/oK
fmrv4K3vSVNAnt6wxGveLmQ14uY1I+RjRCBWAWSunGG/5GFnFim9Juk75tKPjWQ4
7OfT7J5VZanXZJCskQ0rgmcC/URGQXze9yb/d9vFFtWCc+oyEXcmFyVzwlVY1a9j
9CJx+6Z6+AVzLBsq3NmRyUYB+pVxHgXKeGjIdXYv83I4JG1TAjR6g01qcI5hUTVC
jBOuLqFes/nB5vthnbx5VtX2RvZHPJHxisJzpXayEEAFdl4RNRczorFM6CsZo/lw
6q67NZ4Ml2Qlzj7XdlIkiMIuZ8xL174C7AhmFWF0UkVzSiaNqw1jmiSyklDiXuZi
FeP82yU79vIcUOh8+pCnE1ftLgZfeZS9UTlKxk7IKJuQeIwb40/Oz0N8qIz0yqQ5
rzn59Fum4I8JD2qLsLKo94eX6Lfpqc6wX75UHjQmdxwjLkd80VuwM+QuJZl9fgPc
Wh34lWDWMMSeTKGm+iGTaZl65mHAZWelRJvozrtflqtAYWYvyuIy1IOhxG6I7bJZ
6O6aB8GAOVkVEle4RRBj5bCmTsyiFrs6qHvr8HEIg/+K5WnIgvrgwFvm2rrVJ1Nl
Io+neQ1RZDRpLve4fgJlnfikTJxZbExz3rPo0ViusBeSiMnCeak04d+Y05/dOrBA
g7dX2XcqVEJDr3LB7uPqGYa1So3HYkPJmxGl6YOrGQp/pKUdZaMtjVxRcVuv8zKz
nv1B6KUkqhufSK0fywK7AwVo2Z5ZKS9u5HBZayFWQ9z2P00iilQQl+cjjt0HfQqb
3WXafmPhE9POWO3LAfkLh3Qiwvd7kexyGapk/bW1kJff2RRgJKdPmGmkAg55fLmJ
VyjfhkxgwS7d6VWas4EliyJzQtcp5hK/fwsVwqo3NAN3aeQNCs2WPiCTyx3DLlbJ
hSVGQGhsIdggqdIMkudQjh/wEhjD1oYI8RD8Reocp4LExlvvcPluVhxhcN3bhPWA
pNfj73NEa8n1MRwFcG4uLM1DrDGg4u8nwvI5dTJ6khleT9iCSEN4Xpco/lgg8OSB
+ZwXxB1zbe7yncqP87usOVXrvsS70Up/dpwK4v3v2XGXLSOxRLaTJ6Zg/63AjcX+
OA0EUX1RhBbvPO3hKJwWW7F3BDXfg5+n7GMUR0LOi9hrv1anndEaUloFdoH6lFBs
YQyE0zuQQVEjifqLShKT4vsCdv72pID46NWWht7Beb9Bivzz6NGv1HWd771OqWG9
cgEkTx9PmsNh4Nhv3VUUYE2pi5m5mNN2+AJuAJDBCf3/PkXovpYSsBeeW37xlg3l
82V+HdmlbFJQYB/Ul4/nODzH6dZKv8GD5xlA/TFiEnY5hrpXc8TnbXZ2GwL3NhG0
Ex7EzHnN8+mg3iJ2YhZW3pIolbuFiVWg3LEyRekVtKV2f3SVfXsjsBTVTu8XGeTo
7ZGDsTRgQPZ7fGWblq1Fh1m3tQImUxJgZYlbBWgvnEkJY/qItEtxJ7g6tt5sStEz
PD4I8UxwBtfPUE27Y2tpu/uvHhxDOUOEnx2cErqPWh4Mg2OxIcDdrvJOhlrmm7iC
OxRfclp/m5PTJQyx2V9Wps+ONcUQ3PEp5BJvYwVN6p1xYFv6UWTTCiJuoWCZE7r4
YIyXJ9sLDBas0ZGEaXk17+pFR7l9DKaHPU3hyztZAfFOdaFXmyEyR7oK8hZXF5me
PJpm1gJFlQfeKuX+r5d7U+MBO6PXTPqaCSgp3ITDbC8ycl1OP9VtGgu3sCo8CqSa
AJRMtiifn6wWvwyZm5FRV+scs/R1eQDkPqjgoHe7JnsqyzeaT3ITgvpqdD2DENBS
Xyw/kEqCrOdZP+qjhjokpepHexzn0mPFVUOTzeUDHlVUpQPGhTSdYrZllqbx/GP4
hBqSDG7Ap8Y+YMN1phshipKjLXlUm6NObZgXMlYEO+rZukbicT2gd1ck29m20t4G
osYGsGt1arbz/8YwlB3ilYmNZZmDsmZav8/jFVfkvcMdeHJdpAkhQxr9D3jzyWtu
b0JjF2c+zfsrUqw4k/CX5GWFrO4rfkcVJKPanlRO8cc2/bMrlje1AgOZjhQzKPbN
1QeqJoBGzZ9001llUomjNnUdj8PbsYWPn73w5jBa1go3h1Vt2xRlLhNrmDuzL/kA
P4Mmx36Y1diKqDCZWckqwZn1jBcJozo6o7f8CMYpEURnKVmvoJT317sbv4ed7iXe
2Cn90CkRUAgIN88Rb6se4gS0ZDHoA7ImvRB+1OHPCTcLcrbETVT2h7VQCHBqf9Lf
R8aolV2tW0jr4IrMdUlaAd6dPW+n0Mtgt876AA6W977PTtvdym7cSFxdOPAZ+cfR
nU7vqkAo6E9uNXn06olQoopb/88O2yMwRAxCeYwitOlf+uzLch/iv6QLSsa53bon
s7pgWCU9h8Iv6PSsxKOdTS+gSFPkMCjnRhrUJh6URnbUOUguP01rtwKZ9Gk3RLIT
G/czsmdLoSfTaKtyiZ/MQDz8u/go1FXqUqID4ok77j4u81pXAAa5FH7Qu2hPDqAd
Idbrw88boIHybQveVKIZ2iIu8i4sXB8yrfyhV5JkxEqpKII2v/6Z+Hgb3Na0I33O
CF73fgF5HG0JI/3SyhmpaseSv5Q8CoQLY2fZaKM3uTxQpV98FwivoO0FnG20YY3B
Zo7osBG81Y/22xJt54lV25SNWGpC5o90u7RVMfkQGFeeqY7uD7DZF0+XI9gzIvWk
+/+7ca/+Lis0XUeBV0zN/ntFmj+PiDPsSAQ2/jZgkOp7UVM8fXAZKmPijJp+FMxh
slxbjIx3Ie5XyepUibTLZcT3FQj+PsAQhpo9oJ5qscK6g3VYtkTYlwMMANmeFPry
9jFH85FWzcPZ2GTuYmAg5mKIutD6haJaOEE4qCptkqj7ZS2OElc1ozXemFTZNQhm
UQ5p//hZcm/8YbrF2AO3BAavIlpdL95pUne4AbMDoC2IWaa5vD8CAWr4Em8QJSn2
3QMhpt6uEajWX25SQror274m3pfphWTUpMLNOCIUnESE67GVtj8xwfVX9lzzAY2B
nuzNhvAFVtiCq5wehrVAVo4H3XEEimSMUlAZxlTMczaSQEQbjsxkr5Ynfh3THPFK
vO3G5nTTSaG2Lltf9VYz4+IBuvNPs4UdWMgUwsz7nFI3iX6gs9GwyF0rFK4GqsMo
sfDGvR74ugpRF1lAouyZc3zN90Ow2iCeDRLMDHZy6zJKM1Dsmj9KAFG1Ab/o2v5w
EYY4kXElkocogBLWCZGuUhlzfGhhaDzDlYNCehHbMrqxwu22umjgLGlmnO7LP+Yp
HmErGG4c1PKU3xb03pVgXMMzxiuQeIZzfQ2o3R6PBNXRC6gP6Xeu6YL1zbBUP6Qu
lv7bNEAKktZCLV2aWcCs4/jL6ulXrFszFdwCvr1Z7QNenREGh0Rtfkk1Kl42Y7Jt
iy+ZeanoBYrkz+xR0Et+ak3QsonninyHtYGoqMK6JT5YJKfSZkLM5I2K8UY0C5dA
hkgPnRp5gAjuQ15btta2SMGfFdDHCallNUuvhitA3yaIvUBAXWNrVnmb631jHcz+
za4c5KaORQXifOpQZInOLMini7sf0ExoI7RWB/11g44mlSv/u2duQ1sEdIaORTLM
7AwVaaFCZIWwx62a17n4YCtCiX8/o62pRnjEXH3m3IM3c08o6npupvMe7XeGcx7a
SBkp6eWkXNypYRQlKIPpHESXt7OHa6u5CUMbTZnRdIXsISSfg17jFQA+dtEWKYbg
UUMHrfvGMv6nweYb5osKo7TGkn2MmU8p3w14XqP7U0nT8SwlYMTu90rsYQ60Lnuy
2rmCCHb6j+o6zVAGZsLuhFk8XcB3vtTT//YuGw2s4bti5BRFd/eoFZSqa1eEAzr1
YpCpsj9E5aUZGBAALA2y2eMsdvpTA/g7Y16kQ+RKf4wKWiv8RH6J5u0zi2mYOdVi
/QrEFzcSKDBpBOjrsrU7nFX+Jkw9tP9ed+2ytA4nKKmPH6vDyywPpDUlc/zSvhWZ
cho+wIrMivpVfH26BHNywvjxuQ7Dj9B4QL2ma6soVv5hDo74OKSyBj7NUJEgJ1jI
6jXDN4zj5wuJmmXYprd+4OslDa0wJVfPwGNiIiZ4Z1pH4Z72AVfaJAOepL+N/rzZ
cd7CH/pY4L127YCSl7qIRmn5zD27h+WbRCE7mABkBZJThMqI1NYiJKonJr36Qh3X
dC4Om2g8IXuWJm+6A4bPJJ7uE11/mKywna32uen3c2Toq/HIQKQEKSfoWnQfAZf0
uGp4WGcL7U18zDt5WiUQGYUs42yGad3XGMaLoG/uijXqM+/gegqJ7TWEForJrbc9
qlWVhMWJPBOspN7PfPs0SpcragvZyqwpmT7V5klZ4QYA5I2umzXhqth4wr+X+hNf
dJqv1UUvOrFZzZGbRYyNhzhKqDsMbIGjmPTPRyktUjlSPZ15LBSapdJhN1luSPpZ
IyVV5EE8nijifICWI6Gkv1R/uGwuYe+/GH1slGsXgH2ienvnS0TjYJZYGb0sgZL/
xM1ag5zPeRfeUfA3WoHWeaNjsmAYe33HWQ0IPz893H97D9I+chgmo046VI7SITyZ
5xZNNCmcvXImmZg+Tc/xX6+lxQPYmopoHUArmzndK/l85EIxtaUeMwAwH7sGMPuv
qSLBImKIV0AzJ7tnddaoqaXZyBRBgpEvoT1NV3mha5nzla6fuF4FS874Lmgp8H88
OLiSB5xLpPxYSZ1xETMoNsEP8cfDCuN7SNP/5RRof+cBe5jCwQQeTBLU8zmEzDnn
lnKap21wjAOjyNDJQ4Zln6uvbDnvZr9YS9/P8eUjEQFihDpTJEy5SZ1IV9aV/o1/
rEm7yuCbpNqO32J666ehdBU4JDTIcUdpkHbXAwex8Mm3KY1XNpHWYjXEj50T6iN4
oum7S37mDcqvoTiQ4/TmqGsHgclWKkyk7brB8Vzj9TGK0NP6QMYYdtZSiK1e1ouz
+Ie7c3CEJl+3SMIsW3VEwulELObCD7y3idaCzyP3yoLbmzMUdIF5TTqrcD/usnmR
B9qc0x9TagGtcQbLUr3r/k/6H9O4/VkIr9Li3jzXbXWQ96f+g/C1ES40VZl+1uFI
hZhneqlJyT8iSjqBVau+dhn5ydD3q4o9szzexzbqnWYrwxGc3OU46xpHWUJr67b4
Jo2t8yiL1QdFOu+3KoBeDQ9uGYCQpgbGJlhOW/RCJY+Eyxj3Jdt9Pn2jioGbvqYT
xU7raepO+dHO3e/RjAdZDcZtUR7VLXAVDBjIhK+wcOU7WirZWsz8qOlFGb6X7J99
ZG3Z/KCR6mHaRgnsIHrNDKBaZwLQ/PKfIo30Nk19P9NhbvuMivr+ZJqoiapKaiVi
/3kTTQdbQIZ5LzMpoMzJu9wOiJ2JGs8Uhbwb7GBnFxFCQXxJZyoJQzV6Y5C86xv3
AywcNtjg5/P3KK6ksjf9n3ZTP0+mHjNZ2QECRKvXxGgW+zdMOk5o+ie3pDJmJTAm
d/yGXi0SW+83nkAiCnOo0Ijsx/1M5dWHRBFsnIB8RoK+voZEXKz0wmDM05qX/wUq
APTOMNbT3CcAiyj5Oqvu2XZhBsrC06EBZpyD+BmDEuLf0wp3SjJFTYXCeB+1bb+f
XKkYM5dbzwEeUTeyiqNHQo+kgwkJfxkRSEDlZOE4tWupp2wXCBysDrlaCTi/FA2q
HLhnp17YfiUCSPFEprSWNTa/9lseFPPmr2QMMczlutNaO41WrIX/zkUs2PQf3alh
KI1wEodJby92yu2RtF/hIDRgN87zAmzeeoAikcN0A7CzAiKC4lX2ADrer3d20Nmk
r+G90jD42E7Wo1XUttwK8QaqaDKonqjujGeQ3Ywoi9ZMMg3MHKaL9j/u+MqgCPP3
MR76c0EuDnH1/AqN2nj+zBwwEds+QlHNEq74fY1hbDOInUKB7g+oAjuywq2AWo8v
FFJpCnr6S+N/pfgIz4w5qPU5N7hqfFl/q4TPu0VRXlOp82osSTvZGL4goPZsYORF
63Evb4H85vYm1q21ROpAgVZ4ibhfPEjfcMgLMAjIeYZQnlBl6jDTe+bmwarlcCry
xFZpFUZa45C5H1Z9+zKiot4PTqJS/PWfbK7uQyWw4NYtBF8/W1YfVHs2xgigryd9
uBI7U+ghK0e1WzmoNEe+hy+4LADshsX7KCAfmrBhGrCKWspMKeV8j3e+q4IwFoJ1
9DwGJVhL3Buz218QXD0hP9GbdK155dWxJwBLuOg5IhfS0o4x6sFT7b2DFqYstT1W
ZUkuZyl6BKPbbqAIHnO3cr8KnNydqoGDXM9s4OfPXAKnTfv+8g+M8sxYY7yMpxca
RptspSUFxaSDJqfjYn094SG4y+avuHPZ3NMKHipF1zH0vpHfubeVIn4F8jTzIGnw
/0SqnLJyhvZj4cCLhwSCyARH7hQglNotvk3yrfEvLhmChQuCTE8NPNO36kKAL5Zd
51u0uRlDNV+rKZ+L6SmvxVAUv23x8S3kKsFJMw5s+rBoft8m7L90arvZCULxNqVH
0D8PK2FcMSudC/gbEDur91vaUwQVYedAeq4LUVJ1u8nZhknGKUk/fMmI0fJ4QXbA
nmgugvbZFYP6cUdWdU9vH08y/2zbnIsurZLfCzIoK0ECW36QseMvyuc2zU/XFuhB
KtVBqScovt48C3bVpHCq2Q2Aq3NQ4NvUteKui3Yof0uxvpu4ARC0KBG3Ww9kBrXs
lBSO4xHa2sQk1DSmsELPPnhykre7oYhec0NtgeSl5ZgfwehAkD95Ccscjd6QxtXS
oNoDrVGnw1WU/YmKrdo71thA1tQDuXlwORTylTYQqI6SHayK2ucRshZvj4tjaBtp
sMOKZ7CSKQqwNZRuWxBPMt0VjuFH9NmB7IKWzcbypzHykHBFMPqbJ9M3xI2+1AqR
Tfp9Wntgflg2VkkFJTsE1kFo4JyyKh7kkohMsm/xV1t2GNP5e3FaOwmvbd245jPk
p9cMxTsq2RihLufST4dwG2zfW9HXVe8df8Aj+rzIvhoUngGU78ZU9GG7OeiQtvkg
JxeSY0OOS772w0DKphGtglJZ+oClvQMWOfO0Cc1k4t4thmumxj4tocwsdYHbU3xr
OlmXkxBYnD6i/bTy/UyWL4zAQdxkzJRLP7uu5jEq1SaDcxmjJ2zYZLEPPP7sEYHr
u5F2+h+2Ar3MATVY+1yYaLWItHGMc2ro3dPQThzJoJi1OuxaHezPhBDa/M+JRSLE
ug85ZRfdP3zX8f6Nu8zQB0i3vFQS6gXHV4TjuNSq0YFOTKo1mHldEAYpGSHAxMYp
QjPNGguZQgI/6qv0d84sJ5am9yHAOk6JisLrrepUZfHvHeJOP4FxJNU74wnH1YdW
NylMn4votIgvhV7C5iL8BVTkItLxmSqfxrcXlibCzu9ksw4Px0bA2qQFUqRrkq/T
2jzH+icT+MuTr2qNkBbV4Fj7NdVnHEXOdDVdNNmcylHva93oP4Q9U5LSWgIGaKUk
RGHc3DZVaYdvdf+sjgxKyG0has45NpzOByaglJNmmHbMmgpJ7/pKNvihHcmPNcYC
sa3SAauP/IG8q+E9i7AGd77dmfzN5FGuWznkfp7GgzIv0DC07Q5hrddhw62BdaG4
0raWL0m7lIvp5beN4OyO5VPet+WZHrVEjIjOD7taiexIY/XWbW0rI9aCcdrEkrX1
YrSHCpgsIrLYEVPqV8v8m4tOrFZu5O/cH6eSqvTZMlfdaUhVNfhrhEsqbVb8Hk9d
qcc91p1g1jZ5WQrvytxfMbcPaTaG8C2v6nKRk0ZXgOPewvvj/xmyXmYBpwbR6n3V
zgZlE+kXy5dX7PzV41PKF2ID0jYfSzNROEASa+TcMXquUebuuFITPm28KpQn46d9
+Hvk1YgufIqODG2ZlNwodOC2fAW1c4kDB029VPuOIU9lfxBbH4R4DiJfeYwroZcn
AEfcmwimoiRNF9iohbQiu8ZcbfYCePUxHS2hUt9ROVUw81hjK2KoVfrjwoz9fLCM
RLfqUvwynoW0iJC9u1S+mWPX7ocxb7sNvAMc9Qo01s+SgOxIgRheNHruMf9zz+oJ
3tI8RAjcCDOg3Fh5x2ykr4og3mm4vBuQJlv6+31l3p3Fy783eFJoqDrn1DO94pdh
FstihacplildebdY+6+3Cl6TxTt8EiApOYIcNECYsoLmWrueGEfdG2uDQXdbpjGS
lbgjmuCIaZANAsCNDJMLBsJARC/Er+CcvNlUIEFXYfQXTDjSsMYgxDuZbBmp2h6n
1qtk+mKCgTYRcaPFcdNcJveGke3sDSqtay52w0lX8SMVpVcxrBMNV29yy+VyN+Vt
D9BmhEIgspbHmbGDXuyGWN2rCnG+vATz6PHNsz4D0H2BbqyxgiNFXzi4hw1nEyr2
IqJx8a0Fs/Yp0b61VtTIBMRCkQBZ1UkeD2WEz4pmsQcE0upGJ6DeCc+QcdHXzM2f
D0TVEXgZezjzG+PjDImqP4wWcAL3viBnAERpgZ//FgMRDlMjfPRZEcrfZbFyhrsc
r82Kmn4txAa5CFm1nJ4Xw+9UHOjkXdeYRUq92nZf1ACGUQypT5IutTiBY8iXFQv1
ByN9qMrPKVWec/SZmtvJLIfbq/e7YUsKgu31T3KDpeCBQg1/N+KzRKND9bgFkv78
laLhN/JteUDn1NOddvRvZ5LsBRObHAZ4OtT656XHmzDY7BshMTJ8/FnIE8GKcZhB
dEbWMdmRzyHZrSSnJQ7MXUyGjF7B88s5bCY1xomgTn/huUzGFcbKcjgG9OHSASvX
Gc6DXgZOmeOKiD+FDqv3nbGGOu5QnKTllt38CoEIDeEMeF5qCLZuU0ZQhdxDCTFY
lHJHVwKSXcU+xgOugu2ZbFalotF6L5KZ7o9wILx3G4cycWJltR08UWby/mT5BY4i
2TJ0E0kEarBDbfVnKgXSlL7B1EvWPFnKw7G+F1/L/Xmohotxwvm1Cvc8DNMT9NFo
ngI9EPXRpCwW11UCztCXqMD0dk6eqZsxc0EHL2d4qf28kmYttbj+6nZ5bDcY+o4e
rylI0D/yws5EJFlFt80TjKSjweRdbqH9qqNtEVJeA9QHC0E5KvrawdpaLGWbUqVb
fbm4BkzND5KBW0Tn/QjKLLgFApX9j+f/epAP/Zo6eFtiUR0ov1D4i7OaDmRvT8Xl
DcjBn6BlHJ10dy10CHS/xQWUWntNmYdXzNebrgBoDagZ2Kbd7KQKpPYRfIiENG4K
+ROtDOrXBejVy2rW006cHlhCCBwANxDFYfnVAPUQzG+6CIdxfscPXzlneskEa66q
T7zw8CLHnLnSHnHLZcPWrKR90y0YUm3KqU/thkR7AoEGlCLFze3K8SCXTD3/q0eG
vngvyOxSK2GgnZrjhOMmGhKbI5o+g/RW2z0ownezdxqn2t2PY1SHuCYVGKu7GIvt
6Z9QCRICLNloErPYZCR1XxOSNTdT2y/I3MALmsY2lRXVQrn5Kzux0UhlX2kRFOXp
6nAofPyHYMq8g5yMJ6z2MGbLQokyhy/3fYZfKpkpFbBf346I/nftx9kD4oc30+Qt
MSmvQXRUmLlwzqwwi5KSxzSJidcDfjgbqQ5RqU6tcfA/w5ZPEib1wYwVCdl4/lEg
El78n2ybrmc/GQIMAxYp6N1XosSiQsUSSm9LQR6lG+/Xr78qiyINqivRkPaDsEa3
LTFTfZqz7FpAyVV5CyfWSPftWsCJundBWKvsv33SBLYtuefDuMxTxjq9Zy1+xtNE
vf+3kyPuWjdVkHYZuVmpcfsPHMXW3t6VP7NTtXv7zztsv1yx/3tf/dQZ+0ZdosIL
Q4xhG+Nn6dud8b7/kwd5010q/LL2AWXC0Ok9r2XWo94P1usjRRS2HpY7oAzqx8W9
/VXZZ+RIDOhhhYV9FoC9p8vVUaVrC55SXM1XNKLAKeP5JsFkZIIIcfpdObhw0t3R
8m4yk383iCzihFRJeIUO4PI+A/ahzKYnrggwI+xcfvP9ck4bEPpDj/ZkJNP6DCXS
h0IsgfvUCQCCnvhV7DatsINDPFQ3rXZzZlmxPs6XE4cGQlplnuM42884HNsiMCqn
UKFw/hel1tQ0rtOnVHrEyJcXstRAydLPvOxzRTokpm0r62qHILsj607AokxJL8bJ
JJsPW4MDKnh8ESBQv3tWG8HtaV6k3iYsrtQvQ3E0qDMKCDe6cpC02ypdd0jmxMgv
XAuQIx4J/r/jjDF7qyCx+1Ijuq29K4cdUYmwCpINdykIsjVZj+Dh0l5i+jS9Z3oH
B6pnZh11/9g+cWwh+C31iUm4sC3J8NJCof2aQ7UlPNs5pKV2gY4jl7/O4oaz8dHi
w5UN53R9omQoiDKSEaVc7PfPRLjR6iJbvEbaHl4se8of1GA850t81xDR4dR7t9nS
9uOalNuwbCDr2LVdsFt3gIXAvOvZCV2E35c5lAjd6IgYkrCotYH5qdSxZlQHQwCm
dS6xWHNiNq5yakHj/XxA0g4m+gcrrKfRZIfDEGdlY9BGY5X/4yepVQ7FT+ZC3GCb
jZEecjvG6Uk4RXTAF0LdgmqONV+beuBuCusEoW/HoG4Y0RFNREcaoJigogBqe3s0
twI3FMsK2y1p4ucDP/BGpyL3rltx6msUbupfvIghXTdITlPRx7Abiw5gozvSLgCs
Y6wlyvOOQB9ZYIViOH3hvDyJIuvAkFJit0t9YpZvMzPYXHnR4rBMqZK3EtRLMFs7
6Xnh+D2cldJ7WNJSXONod4q8UxLsoHKjmhNM4KngtnUOrhaNa0V9Laa4Kfkl33nF
f0zJcETNPTtlvM10kqrjll9fxZVN6eswlu00T98+e7GrbyPsvgCuKlZz7ZQRNbgH
icFx8UVSsFy+mUSPViDCVSJLfrAxGZTWrny8p+QK5t3D3lEfXEbHo7Tyy2T0VEEn
5SCALnX5fm+qjbEWSG9svB5wb+Rb/WNi0ET/MlZwbsZVWVbZXWqxKjnFNmyCO6MJ
UsjIt+DBz2e2L2ThIKAEiV54AMqSAT4z+yIsWq/HBQAWsCYhM3vTs9MRVKkYrvrg
RrRnamFdZ+m/hXNAxXwQ1Kt6PDVpyKTa4k+x9xPKXauLJet75BQUFWU/Gyo0fObK
M2YjBn2+AoqJNHWpWxMH17KsDO6bkMRr/Ctb+XzcuZ2G2XuNIpl1fgUChswJGF+s
PcOY86rydWratGijcktbqxXCeB1E5TGh9bMOoYOk2C/F5RChuU2N4hqVMFxMS37F
F/V/4oXz5iTjM3x1DMOYyiAXkbw0D0yYfFWImQXZmfk+O8YDwBRhtRrpP1+LTzI+
T69rLXxXxa1ovVMSfUIOrk/k0GOu2YH72BCg85W7hP/0IMiIKyFoW0FKhM5kIVb3
/Av/ainR5S1A331zPVXKm7HHNYo4fEatR7NJe8AJ6YmC5o6C+xGWLc/dx7oDEzXY
wZZuIueXL+NvGY0HabrEG9NC5/6xcIQIMcvcBMAGeytxs5Ecg91k29bYJ2SX7tds
0UFrVbLhIEEyglHfEIF8ISjQyEbBL/kCuKr6QstOWO1hz2h5VvDsqMRrty4T50wL
A0JBZg97F8bHumELbiHaS0tp6N2HGs4Kz3iO+vieC5M+tviXO3TA2Ku/Faz6CMVV
AO2xkJAkac/kcuQkn5iKKiv63+Ki6fbIHfKOflwUzn788Amni+GsM8j9I8oRbug5
4a1WcxAdinltXXEDkGo7qsQP0KJkCLqQkyOjdkn+npY7Mj6lk6/9oisWtdSNwRuX
fBM5Mj/NrEqFRms/EffrT3sG6OAamK5ibazhFWYqwKHPbRYyrTK7txoQHHtgs/Xn
6iBbGq58bf742YxmwGhnCkoXaB6bWQZPMmlTm2i5Uv+5UyPcWE4LFuxz8+DlxM4q
wHOhKC0cSq2Ko3p49Z7aODAKzJg6z2NFYsVC8nRs9TwShVkWutzINRhxpCCPWgJ3
BlfUmwRgkIIIzt1z8xLe8TuHnGNcvJ1J+7HiIGFKPBmCfW3tcmgzR1Gm9nZuxQ1B
IWRlRaUjSb4Qy+7Q1gF9cR1tPKIOZIrei4OMr+Skaex5IaW12m9TcBzQSyhLdIPo
lLPHPg8vm/2JX7wwlGT1uQoHWHVDDn6u/2FOV73GC8VpDuWSWEL2TyS741ALetDk
8y1acJg0Ds+ROmaS0R5e2gL3EETm0KWISPzs4TfqAcewKk4Q2h92+CONHdi9qEzz
Oj3U8xN+qe6tkeKM2hOMQYXBrQG6guXII/nH21IJX/h55bl0874JZZuiOdSADne+
VAqNkE+twihlzIchxKzRfhV2cMQeIjz2z9aCPf0ZP4S5fET0JBbaLXHuo7NAnztc
gRdJY45TDmpdfjnDfUZQaoA5JbIwvs/MyK6U50yKkKytpYZHyJMGMU9B1njiiXCB
E8rkj84qYx7ZS/jfDHulXW3S8OhaYhN1Dmofpzve4IqIO7FptcuiODwt3i+3KMmO
euFFfSvHf9D+XtyAmjPlgETKWQDYNeiL0aVLAsGTZasoFIJH0nRnjo5Vt6KU34Jp
OSD0uRZfKbEchdmBgMYMD/g78RmGwxiu3qAb+aVX5IuEorwDv7SsfVuI9RyWtXXL
ISfgpvQcpLgbxSJzmolny+d0ZZBcgHZd3kBqyf8resC/6L3fcGEShBSm50rArg08
tsGIDcbpwPcvH00sPEX9JvlhHBYV+WrwUTloYLYi3h5Hnu/Wnrg4rTa8itU1lRkD
YO4E5cRZPCkYvoNbXPu1W8KrJi9TgRvv77m2ybAzdJyYlw4Sh763urcgIFQrnzeG
doG02TVKHS07XcUvd+sl+eSyWRi4m+C6HSDY2njGWz/6ggJBQOWoy8Ypc/0qVaUl
r20KsPK99uDFqY7Fi2y/hS9+ng31jMMy1nQMWmY03IMsIhRnZGG2xUGx6kxGYk6U
pdljXy1kx0S7dCJZYUlICi9hl7+zmVI31o6nPRWPr9u4RLCztkGZ3no3QvGkhL94
tdztTnql7JtYX7pBYE1g00Ueywrnv+pymlw6MJPggxHNAGFVORQfd2O8FZUWUARf
5YnTSQvACjx3ywBsdKwTh+n5Iz41prrXcnPDBigCQnbfsXCtWDFc4Zw5l2Mm9ZXa
orenZkQcWqChodN+xh5uwwADfMnnQ+reCfn8KvyhK3MKWpC69rA67Yj7ekNdj6L9
U7TXvAQESK0hnsp221hZKfeqVynsUaa06irn3sla0GhkXSGhfgimFBdpmpxcvAcb
zu/TQ/LhY1dZHs997jVeOVub6d1s6kxK8D2wdFkEWLd4tK+4mDUgqTdGQpedGDCh
ZTk2SeSQ62vThMeEZm6kzCGlrk9nCP8oE4iJmGtxi7sSLBwzro8JeiPIPLQQSEHX
eBypyn4hhTdau0P2achzRviWLi7G0UIqv00SqIlvXwyzeFEOpk+dJStuC6wHRopO
kP5790n0IfDSjeAwDT74mCdZWW2obtlk+9WMhEvOrY/HyH2smTIvTw+K94G4a5xr
5WOnBqOMtAQR9LShVXjQl5h/ShCZKfFAMJMz7bnZpgpJi0iPDeVCwIkDHwvNoBfc
QU1yqXHYZMMUJdDJ5sXskXBT/CvgyA2sILbgsf5ArkyPgHbebulUOrOlT4JDUUot
zrJ5c4iO1bCe5B7Ss5k6r0LXK2e7Mhjq9wSCuIpdH1qENWsVkFmTJh6PpuREeDox
s6r0HSRYqv5SAEHiBdyj6v0xrEbWfLy42eolpYhDb3+yzgUzcKQTh2RNPFlzGvcl
xBimYOU+lenqOQtBLsLRo9Q+vQoDgUcaWa8jOiPR+HYSJ4Q33HTKkcorUgHsZ3yl
qW11fWY92667pqO52Sm2ZC4l6ITA9aYtB77nbVT5QCgGdFX8OlvLlxGf5dS8AafT
Xk72frDvT29cRpID0KFPPRPrJBjnCTlGFS62GMPROmnX2JC1XTqzzkGMQs6nkpou
r3ddOewBLcQRBkiSsNogieUFppu/i0eKBqi2WtJlMqKMwLLrFMtDGE7TIiTbG74V
LpeL5rTfsfi24N7fZUqpMkY3AveqqC+zrjeeM+qBmKljhfa8i9MYq4LB+awqjlFs
0b2hD94EGcVxjPj3A8eg2HfmevbMnfC3a/xrdzfWMcaG3qkfBGIw9a3QJGb43nGY
Gmtft+nqxdr7SU8vG8Vl98fo9E4Yk1ysF18G4JMijFa0TKuR+qTwe+YGl/ptpbFQ
aKzS4pw8Iajt1KBXcMxtEYHNb8H7TvO4Lf6a7OuV4fPAfwehPuGJ0VakrQPeUWc4
YAJ73F/QxQqAGpTLReOEXxSOcFleGYWw7Af2JEC+u0yFOMjfiWGXTrs7fut7GJmp
aM4RIPj7Ls890Lu2I08ZmX8BTn2JXy4xx8X0NnTpdWrYmZosOOLmc/81BSUuXgJ0
xneEGyyvlUc6EwIkcWAOCsNIKtsTRNvgf5ooLNLQt96AdTN7rBkgUIqmIcR8n8SK
vrGndDvuySSI6eccmVRXP74jmnA6UrvC8tWidrb/gaVZDGivLkJbLiLWx2m/w3uP
EhJ63GOxtXvB/UTyuDNo4J5mdIS18lmTw4P65j1qeONPNNIZ2FkpaVHQop7ORw9p
kyEttJvjdJWYOFXx8bBmsKIy3jMwd8u54hrESFsBG9DdR3cZJW3Ei+0REti815Pf
ItDYGwh6dx8tI/nwGWWB4vFJRZZd7RyIHmZnOslYnfFoW4j9fwu5GL4opEpQ/JBC
MRy3rmQzd6Cku4/xJLauTJ++O+Ot9fAVz5EXN7t7RA3j0obf3gdO6URI/Yt5yz5s
ux5lfgR7NqIv7b0/FPH++xun9qtHoa1uHnTe7nwmWs1l+oNpTMAN0YnkcSZ2tzle
nT2UqkSGXboT6n2CLEJ4IbLTlXl6a2jrUSlykwQTHgIvQ0HNSgTokeBgrEOaoFu2
gFcsvFXGCd0gtbx5cNHR5mIM0oQn4ko0vqIL/TX7qTG/qrqgssYeWK87IF2bjLdV
AicISzk7SQ96YDxKQ8wdSUi4h/76XIgixaPSiUQfUswE/pl4JvJ6BKOY6umkmYIS
UPC1qJVJKVMIaE2XDl3lLcbhVXjC1LD/ydweh4FIg4FXzYWu3Z18mTUkTfNuigU5
+4Uz4p1I0scH2hS0mtf79wPopk7yxpQgQb5xmCDjByIMtCydSetP5R+5KUqIkP/F
4yV24tt7ZtRI0x1R3QymvtmZZDf++qyDeRtxwQa0L7qLEdL6vdKWKdWleMw0bTsy
+zEU6EKT+YeEA+ND/By16EwBfbLHQxtqwdTUra6PrEmxGLt7fnYv7gDI/nX3flHV
Sw3sGkHbahxIQMPSDofCHljHDz4MQbH4RTbCOKqMLUGAT1wPyMg1x0HiUnNnm//i
1BqQLpoJ2J110QZFpv/JgLk7jz8Y5WfW0j06hTNoEOCta2Gr/vYAnkTKFXWhBJaC
99QTLMVbyY/z9DbvZYaiOIsZk+TdqXr1rwm07gZuc4pT+cbxkm5fA0ilXFxVugZl
mQu92nxdSz1TkkUDYu2a84fnhTSL/jvaH8UneI6QIZ7KQCWgsS1pQpKOVZphTB0W
9rgEJPGLeYCylUWQihUpyCxksgM3W5OBYIC/zXVmeboU8CEsgyOFBvLtFMUaEq8F
RQBkzW5nczJaORkMn1wRyaYgtJGSqpyRSyRiktUjx6pv4IuryC5AGsCAqoRd7RQk
oMaSNsvCmVjJfYPQ0DMo1VQg8TZH7AmpPI+qh9oTW/7MQPiF8p+K3enKdYTf84Pu
7aBoSMt5s0I23+LFJKbUbsLkP2BKdgrxJnQOSlutWUGyRXxDpMAxh/udey8Tdh2A
K79WCK2EL5Z2QgeEgFB9H9az9WMACpWcviM8WBWjfZwQ0UzpE2R9VQrEMpVlE9Wx
BoNIjCuewx09gK/KtgZZKPF8W6sFneVNRdRPhUMNF5nKjczV2fkqNnTqg9zGXu/T
6j6t+GPSGsX3kPOQ57/Bbyo4isv33iQq40FDjgtSY8TdNr0Q98THn1jHdZW46+se
XQu3Qx7xcBEg8rOvt75384STuP2Dr4fqi0nnEjhW17fC0s9V2ug8Ue9KWWztsu43
qw1EeSV4LeRLM9m9XlkNgp4eNTzEpUsZiH3WAvFUZC8OkIs5pjyq7aSxK2xLTOea
DgcUv3B8z2NnPu2lmGtWweKW2Jy+aN6Dk8FP5WpVAQxFClQz/XMnaz0W1ywL4Qae
6hWNmXlAP7Dnk/8X7It1EhgF9OPHhdWjuJCpvlxMPxfQcarOYvjExB3ZSk4M4puU
bQPITmzdkPjvcZnePdfw8yRL3XwCkMCagXX9Ss7STa6C7zR2n7Mn1CQDxglvYJjp
w+n4dVyRggtar3nqVMh+aFK/9eTCINfPM6kGGeeNUjxzLZpHKbrLgo++jQDaM8bO
smpdyeFd2gfUaQxphrJCAfq3QTL6TtMG++iUfCAOuZUx0eRDCkD6xLYUZGu/mDlz
MSfhdGFbh2971T0DgX51uJ7NhnIyNYX/vJIhPzDeJMkK3WEv5H4sQRJ6CLgoyOIJ
sIJMx5+UC6H6Iq8CLRpQ053RLI0oJ/MVyYHm4vDjB53DLujk+W/gbaMVwx+wNzoR
LT5GCfkuG2E2fBobIv0g2N4hgcUxWWDVA9jXvG1uEpe71FRZ0kErXdlI9fYZ2yHw
CcD218jUyB8mhwMpo44C35zA1vTMtdGInT22jqkvYegXfmXigEuXT8L0jOfVItUP
jzyJS76NhF6MxjZGKHELgUpl2t23H/auCVjpjl0lmEwMmciy0GJTEvDcBRjVqdFu
Kz5ptIkXczc2nWyyl9WxqTwURB71R4vGyXefBj4OWnlaY4ufDNcUDEgNpbIjtzKp
CoV/feGWz9KzhJv2NO4oF7A0AXOPFm0P3vJegZV5f3RjKcpv6fCAOCxrmOhR6b2Q
Lq869MqDujCw/+SzJCAzrtiX1VwtZI60xgGg1v1o66AEF2JdpA6bSo5KGn1vzeOB
BEqLKF6trFcPqWRqzvLWWhvA7Tss/CVDgLCjkjPKJX1xt5qt8eRGArl441+Vtd2n
nsgCPqcPURCSE50f3YF4L4BuvJwxuuAed3IRVhd52b493ahPXTMJVWRr5kjVwFlD
N4oaKDPFuS2ROvCU6l5TGFJVFOZMQKiD/cWowjtU3eio+yvOTjEnyTqxNjUvb7oO
D2gC7GZgpua/mHDHWEiXDRI9rQPNywu4W9F97gHpLl0fwhbMNZOBm0nF0oVZNEIx
x37L1+c18NEV9TVEssMDUGatHFXIzWLn4qR8pRCJdDdlPoF2ULZpKXW5BC3QfCXg
XWs6XfI74pjDDcKoF5NQedRUI0czn67u906BEbatX2GYCywHZ0Xrb1c1/7OlerEb
gqU7HlRI2oiDWaZAQJOD0gbb4vdB3LClb2EW+gyvOLCn8hkniOzY7nG2Es8DYEuA
IDALQl1UEbPWzEezgs/0LN6qPtQFGiawcpUjjgnkO4bAXbrdt6RB3X3/SZIqJYTr
8Ez+GP3W/9oPkcQv+Bv06crLw90bRkBaU/tJZV50iTaOWGez9N+ybBrFYRcUklvC
zScSOEYLRckh+MBeI2EKiJJ0NB4KrkeiS8quZ3Bjj/6bGCNEI1QLTzrOqaGSIe9H
1J7tqwIMDHIjiwKC9nAVPOdOtlDcoBEiUDz5L53U5NvhhEk+HAonE17UjQftLUJ7
LuLceQuFKPWPs0gTaGJVys3dQP6RNXmHjHpEuLSI3cTymNxwEoNkRnYvlet+heOi
xbSBsOmMdMfG/snOJqAvpxNdsilbF4235nNIVIJB0S0EbopQPfAq/3zD5ASaOSck
30C8tUvGf5Ot2c9+ICkM0bZsCL4toOBTiwAeuP1jioMlffXDQbbvmCwvsGA28vBL
nN1PUee3eZVKa9Rb4+p+UjVrQ1IVKffGZTHx7Grw6jV4DYGYQn7ENpe4jhX4Lsti
KzIfIp0HiQHayDcMfWJZehggOhO1PGJF9G+a0JSZgAH6su/bQnbvswIwegAq2WmU
93FCe2Ugg+n0ZMPEs3vJIKUA1RJ43fLJzRdvEQY2gM9ptI1u5h/07eRKUMo39Hal
Nh3h67oPp6EB/ZHJNuOEHpdPF8zfcBHcI5FOBFwYolwafe4tRt6L9YORejs7bIBc
1aszV+WAR/SQLuqNZfhPz19i3Hxq2DM/P8TQZPlN0aELSxJt/nWZIu9Oq8iN+ufz
dAqzoofUN465kpXT3DetbmmxE+1UaCYIR0YAfFNFTnUoU4B9nWMYDg3mniaoPfgJ
sr7z5ww3jP7EkhpCGu8nskjeh6kQUoi+Nf+ibHokNFXw7UYQ8VEkC5ndxlF67rIY
JkYNOAmd8RcsPk5Cx1yqlf4VZH/tGx8zySJo5E+ra1z7zstYiviD7w6UqONp1B4O
TVWCe5NOs6p9CIv99Uos6BLclJq9m82yVSTe72mtB4tt9QU3nPgvjQ1IzQRT0YM9
WrHJGCczdJENMIvQd8a+EwO4Kg+iTY8/pdJOZcsHhm/mcS37wrcpJR0OzDg21BBn
qdmFeVQM1epWew7uQ9CAnwPZ+PDvbTbqP1UYGWh1loerTqSTQnbUzZjLmS3JAu9C
Wd+3focQ00Q2Jz/fYMzwkjEyVnvq9Yr9L+tT8FySWIQQ1flVttpm/Es6LSo77etz
FrJJhyUUcnBuDIlZrc4NS6YQ7FU9mRqNVmSIRPme7YsqUGd8kLgW2/tXHZ4S/qWy
qObfEGUZLsFq1ESyYnqKtjRkWxmHdePfhtB5PLMtMNEUR//EF7Fy8cUIKM/h43Br
i2cT5TMijUsKxV+9XaMGvvb1S5IgGv4b7tqSjebmOGei2TbAI1C8FJoi4l4BB8we
NOK/5aHYKedAb8s35wJyze1vObsI6jH+t5/4eyMEU6735DALStjuoemC9hNFgUOz
rGbGCpECkmIt7oIE9sUf86QPaKxoXP9Z9zlCgTDKh4epeSsnWK6NZf/T3ItXYXui
rhxAJNZ1PnJ/sjRyfqNx7gAfu0RH9FGJ0yG79jXIpf2XK2ZK+/9cr+6iC4OQM7Oh
OJwr+PWz+NAk3Ig7GHG93hRKE4DZ1zYQnVCpaWAFLq52LCxOrAYBYcm+q+wnUNze
NBvPlz0ax33bkP6G1rLayNqPDkh5NuU2n4Q4O3v2+BS2D1IM8tMaqlnF4pRfCVNZ
vc4VJXPzC7YT3kFqhm8prZFK3U+/b/jeDzM3XFCQ5DVpbVW8M5Q/HZkE8FDB8D9a
AE3vGp1E5KSBagzdrAss29evL0GRUbLWECUo/aYWXhdjE/m5NTBWF8k3Cf1rw+eV
/cvdKZbBygSPRqxPuvYpRJaSMAPE8wXASLEkdXvlybLnavnKAxYex8HUl6RbidsN
90KMda6tNh/wufNx5e9PIkeGvP8mPVPvhJYm0I68Sp3/g1zrbLY/eo7lUzfkseog
55U0A8HYlq/syknqL5yW7BXO8fjM0HVUj5WDFOUmQ2oDZ6UvETIzxyHa3QsMPvwN
JLya3Xx6ipvQopqW+wefeGBSRBgl9W1LhV2Hm73z5Gs4ziW90MamUoz2bYMN5qFe
042y6sd/xVTai56QNPpFPL86CBzFwDYtR3B6xS7uMXS5vimHXEFtajj1hGESW+et
9PrzvlHe1RActLXyXZ/OO1Bv3NkQfDQV7AHyvNtzAN6U6k2DyeksKmbo7wqrfbep
NuqF8L6CdcFXyjCcHbMdvjq5kGtPdeUAaNj5tFN2nG7fagHL34214cLVjHZQsmPm
1dna3HKRPa+BT3S/lvHn1Z1SJJtSrmZ7V/TxW4VwcnsonaILz+0qQzf99ZIDxG5n
mpYQ7Qw1w2rw4/376PojpCPYebCIuHABRkKsUBpmw2x9uXt6PGtEwfycP/icB/Dt
LuIZhsgRTUWOWyOvQ38wXgqmuBSBOO3m5kMtL7KzCFrrTDBEsT37LT1aPTfD1yoZ
V5Z/Yq+jPORp4X6gkfjd/dTSRZKCnMJQP7WUvhbQ3doYzyQhH7736U9QvkwQH4Ns
GV/pkU4jTBbk6Uy15edgS8x2kr+5W5bW7wx7UweyBg01NhWbRKWDM03ksI0eWjv7
3hgFElb8HmFxY7srlCzqA+2Zl8qGb2JwP45sGyBb3emGJM0LY1v0xYy+qeyisIyh
zFagrL9V2qvBD29a5kC0lHcUmGaNejF0dC95/52F9PaNKqbkrJChoEUZT8yqO/1l
7B+A+hetUsMxx7oUgVf1MUYFimEl2I6rMbIyRHoWzel9hxVqv3XX4Zrt92WAfw04
215gsRcRN0YYIRAif2YY1E7TT5d6qj3FBytYuNM5pWBUmi+Iu5UENt7QdUnTPgRR
zSy7s9CmmE4cbVkh70ZdHeV6s96VwUuY1SoKcSNWV/izR9wZJcsLNH0Fuc7+gLmx
5SDcW7r440ZH6IVUp1fiovJTNpjc1Px/3iIQhnez2T7nZPI6JGjNRjI7cBCjXc5g
Y4w34HR0Y2IDICeXRz4lDVCOtXtoePyhlifEYBERt8Yd4J4mbdb/Yi0xDuCDQcjD
w5PMKqjafWqAauetan4CHQ/ryGExMWfAYRlPkYkpHEa/grCarXDO9E9Gt2RTrZOV
kUSRVWVc8VIMwI07Tcn5vnxedk2T5eoHUdmM0+vOYLAQneS5TsTJLpBmeUP2Mv/P
iDwN+yfy2ZH3gUKyDb4NvHm46PLAlzD7CF4MYQlgFEkrBHnjnHL16kfWeWnB0vz2
MjtgIddaDSf7oEOzkaZdXeu8LoRJ4+9TnxCqdcMopTzWdEfTzin+fOCz74mXZ1lv
2aTCjhwFWe9FYqYTyOU2Tt+vHEqNE51r1Omjj+tk0gLnwj2nEOx91+e78UzBrnDG
KyyJGAlylk4vTEJ5x3gMm4aEavWexKpAY1SH8Hxsp5l3Ro7LQs5yUcM9hUsH2lSN
ZvAAj4WfYJZXe43WBRqc8KiIykcKUTKbbBxAgoa6HgmA3FRMGaufM1StldkR3V+R
yqY8HI5RVDr/zTM7sg8MsU1ynAdIp6/JUiEaoBH02otsMBAYHr5Z6t5++BzePYo6
BiUqJhvEdu1JALMlNCxlBuuNeWntIenAltQzFZ+h+hqu2KnVS7Y17hFAibMsrz14
FsLeKgXGuQvk4QUj9hajITYc2HWUvilCx1hWh7eJmfqLC3NIz/bxkw7nwf0IeUtv
/WM1anvnIV6SoxLkUZgqCvTeZsmCfP/zzWMFscoB4rzJQY6ySNKuhNvblob9r5UK
9DbtuMwrwOwVfm4uoOyX3Ut8fbVB6+hre1AWwwUFwhVVr9G2tEnhwxKybk7BikaG
GwkoSmq3W/LIEWqU46VCuLFxBZpZn2s27xOOOrH9gR7pmH8ToSX0kgH1Axmz5rZr
QT7SG0rKdbSQArAm2Kc32wfjSWNcq0vLbMaL6btvem0JIsUuy7GDTa555ArV7vCN
g71LuyjGVzFoPpOWRfQe3MzNQByjPw2awjcSaa2CYiSAy7dGKmWH71exkMikVn60
e7VvErv5hgjX5LOJj3P3z6n86sb5KRsBpITGxuOvPFx+rresRWypxypwXnYR09Ow
KRG3AGtkH/ot0VinJtXs3KIlEo3ECnva1gy4jqQn1wj/uZh8iqOtPEJbPSAVc6GJ
CZ0uabfs9SIKdcZ/PKtdW5q0BZhsgAy89R84vZDdQlRxo1ZF49qjI61VaWtZZuB3
MDzpPqlib6gAfMOE4hX/b9x/DGGdQUGfito/Ppe0oB5JRAeCRFD3b1a+D3u2zVwO
jxiem81dxEnnELwBT13PhclijdefWz4XUobxg+0zuQhhwNC1oPLzIsiAzc9r2wS3
QG/RXwFjrM9h/4KmlOKXSr0nWUYPHyCTHzqd0Aqq0PAs1ZtOrgpoqwQoZNk/v0fk
qC2h1FENorh7Ll90womPTKWE2In9RkjMwdxaJcObJspvY4j+kaRo3Ydhyzwmq3KC
z2vxaxsHdBLVklsFtXEnaIuRGUwJ6gyOtnJXychH/RtWyaVAlNNNAMrfxhbX4p9r
Whht4rpWo73n6BfW7dwVvcOf6+KvCcA5vk4BzhX0yp84EIkoLQHjD5BjP/YKVZ+C
ZexL46oWE1NQCNZYe+zpbjKWYtA9MBrdTzvunq7l0JIJmQ6Maz8KbwvwO2WiiypV
oPv84BIyPTUmI3jIMkAmuJH+qeyyExjays27hqLwusF95xYr5nVV2jAEHj5vCmd2
tQnVbluV8tf/XQ0KaTS+jwv7EOw6gnsGs6ENZSmzLNv6PDyndW1ZVpakJYW0e0IV
DLfzOjjsdRaq2vuxPah5g0MaVedMSHzaaXNrUob0vg6ykvDzmeevUC6zcaO5ThlM
AZdCnfbe8pbX3vLxI1DhJ4TkThRNK+ya+zMednfhJRAC2RCdIFnXA9UqJ4ye2DWh
iWGsdL+8r6bVRbwzQ2f579pUbkVf/hVQ4WdVBC+LxLuwZEodGQSSKmBwyK3yzj5A
+drBoVgTvXk1tyqdyCb4AiRzDh3XZ0JbXKJQ97u49vfvAYxOaNgb+n5AeFL3eRO5
85KnurKo9fh0yUj/9Ut3C7XIotDexrn1KEs+qtWXp1L8g6KW1mRflTHDBjma2iyl
UJlcXH8SAKi66u6VzmCqY5MvXpnKslHUbe3kZAmXRzzqxUMphT/RtY1jLA9oPnPQ
1JBmkVsiTM55bvfEzi1N7kTa+p3S3hgydj4sA1YgdyaFdJ/Yk0+vV44B3tN6DWI5
BnUDs/xW4T29be+xZBAU8pfXQmb2qLP/JNLuP6UnbQ0rMrWWRfRpAkVZ2+Cf+Mzj
CIIAqiAAPwINpU9Pc1DYpW3ms+/Pm1vCTyW1g1n7xUmme8/TfcH4pGT5uxuAjVmi
Ci/0KnsIEQ7qvQ9nZ26N8Nm1Hw+AOVe1aEGbgPkPTIC14stVuWH2dvpqjrp0SAVn
8tuUMMLz0l0OWWz87uohIqhLFeD7qSlhDPEEjBoImecg3l9OxU/StIjH40KbuAMU
hed4VhQoEWy69mHVUjDwZupTgd4qZSxI1ZA7YeIBL684Dyd9ENUlbCsRcAoETaGE
DZVS+NG7g5Bs01VZv3qb100naRzF9nfmqcM10YP6ACkIBo6JjmtSYCUeeZiSL5Qv
sLT6pVqHKkEwDx2R9QmkRwjClYpZ0AOP4NeaT3IScMhwx1C/iKla11+D+bumpzyj
4QJTwti+YksuDkRZrzACy97+1/5Um0Gh8p6WUDgaoRvXDpvqqJxI3ttykbSTdvVh
xYgp/bCsVIJEe8tmXjunSC+beJo1elW3et1sPmbFYY4WLUCat6yvSLb0fX56Nugp
SdgMjQifAvXD00NYUxhOSKZXC4Aidqjf/lh+UWGqWClRpXt6ayc2M3dJ77YB0e86
0DUM1yso2m3SZ6jwpCvjeQsisznYwzVBYZOnEjVZZa+V6cyVoVLP12bpPXHwf3/R
OvhIiruV4bul59ofabuOSM60V2cBjLjvsf7+QUAYAfFfixGMSumOX5AAaz4nwjJD
p+bB9quAjXrd/7lDJPR9d56kujt0+y8UkCygsDWhSDuqZtmBIlLshB4y5alEoVdm
AYyfjkoQIa9YXlC7LUPC8Cmcb5Yb/HGOyEioem53w7HsVaZAZb5VFlOzK1v8ZfY3
g3Vea5ymZ8FqYPGzA2aQzZ/R8p5MpkzBNFQe9zsQsWRT88mOr2fs46KGTBUCjALw
O+y2j++eLBWmX87j5MNqY4I0Op8u3Esgeaq5l1nz3R2AXT2KArwBEWvATrU3QYEB
qsH8hR/lPhDoapG5glPX/eFzq1BspZkr46AJBox16/a8oPgQOx0Z3vMJt+GDUojf
Ue/boXXdWFApeyGDX3VtmWIIo/u7plATSD6YMSUF7+zJwRFzNiUTKiTdDBKLyJRg
yGBL14u/Sb/OaCs2xMv3GUw/rhW1fGUqie0Xo504BgVjJM24+ZmfoKvvNY2on6Zc
IbRdxLIZqvLu1eaKlaRy6VOV0x8ehb+z1/6n09kWbw5HzvzbhcHLXFBmz5Xa4aGl
ueGARcefLPpGZZf61i6Iw0sGJIHOVWUV7G++kKOcZQXwoX0gfFIHYTchz+E29lfY
U0uK8zwEeRL0I5clS5UpbuKHgI8I/Xbt52atnalLp1hn1DTQoZ4dGapgQHrzn/C/
q78Ic7lu1RSAFmzNZLhQ1LOm+OeC3wIE9lizg/gOuKU0flPx8gS7uKK1QlJxRqlw
WFp1H03o2Jm67BOC9qAOuOvJV5eZyVHMwvAxEXEseIaqaQDE9g7sRIHnYgqJkbW6
SawdYeKjmAskbKBdW75G7yubmKpcewkvxmrY0uJy4OKCMcScZgrE0QSA/iGvvSsr
0P4gbgEFXPnN7jnBg989uIpvXVOkEZ8JP9rCrXLou/ok64qEFnFcpt6WM2qCJd4X
8/BRKgMRLh0oRiuslxhKlQFyZYXkoc/gmcttjIEND5FkMpJCJqvKFSkhWooi2YuU
zrj5aF7hBynlD0mGqifpBAfVqm4Hy1LLisn7hgkAxZagZVGSeVMCsIXv3Y6j1l1R
90rWfNlHvKsUhFFWUkpIfVs82lXJJ3BpKxZ0Was30NBHulpT3q0WLRAfDeZYGIl3
Rwheq2Dy9Ictw2PzQ9XCS548AB462pzKlfJqY5vf72yyrTzM0WG5vs/EAu9s/elx
VSkK2HRGSNn8nLCnCex2BNnbk3K84kiZhXBfEX5Gi02MlTHmhpChKSmGTHtTuDe+
lZZ7cZ1xvXW+2UBEoOrZKqNSr1W6PYAkdafU3DJZL5mj1Gk1xO+P/NO+kfVU8ZrR
vJHXjSTmFyOPQgYI6OBwikiPrIHqCq+9iVo9lSThWk3dUZopSg0C4L9UM5ElvAoA
CGGAHJYIem+2ipqGnGl4bFV2daVMwr7SqAeLm5BhUr3PxYrUzP0Y01s2K2JLW3c3
BSVMD6UDUB8c76RLEoTjIsSnrxaANrjpf06mnfaL4TbM5j2oFnJtj3YHrY2HyJh8
2FvkxutbNleAdY1rzanffV02mbRzBhgK029uoJFd+9F1m1WTT4+1NpODNFv4ExoI
dv443BwT6pcTSgTxUyXt6+2Vo9G+HVofNsCJNvt63Hu99JKL5y052XYmwX2TEHiz
nYDoh+1TuNa/9rZ2L7gDol+vzo5cJKTOlvLST5hS/X1hAsEzUqs3HS72vDcuhcXB
6jxt9SxzN8yg8JOynILwbC6nUSqw7AlkphmBZd0K6qUJE/SgpdmcqkzDkIsHKm6s
vLZq4AFCvyRgQf10Uo5UUPbW6UMG+3Z4a2sqbvSpxG+x3pirR2hXQCl3B1QFGoNH
OWmqRRMKOap2XOkWlFARXCZc5RKfYUVLYtFj3H1mlsXKGa0TSmh1qni/NrKuLbzt
r3WsxQe0pv+yF7OIBoE9h0V6hL7cs78xLy1GP8bf0rdW+Ho4tl8gq7ZyRjfP1LV7
VCnKLEXPjwj4cyYYZr44Luunt+LOcFfGQeEgoYlPz4zSoAVt9q8cuscZHQzCJegW
tm8ChLaeLHK7nTHyYQiUO0qcoAHUdOpKU5lsUVIq/Ki06KopxvybMjAHcHz0bOvW
DTr2OVtS1kMJLkrintxiCbB8+sDR6WXHlkgN4XC5xz3SnzYGl8UXLDDtLnk++hF7
iddeZl3U2HIkwPjcSubPlDMahbgDQCe8rSt3fNHT436Qb8yr9cEnlYkdvH0bQa8W
if2RSn/fTIph2zDPoGzOsr7RNSAuH/C4EP5198l9KxG6E+y6g2HYdFJBJCazYS6B
DTBwLIKlLv8os/p8+EEHvarfUfn12qv0swCjljcvyWQ3FH6YHM5RBkkh4S0D0kAg
m5eT1FgVyw8SWE/yfpTZ+CfJjrYmOlHHJ+923xEZbm6IQ0tZT0BATzYkuvMqcANc
3fLl086j09z2TCTFd+19fxCAaZgTgMkab28gpHgxyYwqxnk7uBMsQR/oTJaVbYzc
tGKOrz0FE6XE3xoJBO/aO4yO6eZVq7/UewW6Jo8HTksxln9dDTKg+c49RsGUtIXz
d7kKP4XS4UZ1j/jiimURQECGWswp91XSMpkZNi0RBT1UODjOUKbnT5IZlrKlJ09j
L42F6RoiP819YV9U7WcpkQdxQxEqMzjNJwB7eS6gp2u72T1EFhyc15YJb6smNGuZ
6T/MS2fhHdt4MPsI8FPhT1iAzHxy7QnTLjy6ovBDwVOEpCmeXPcO4/kEtyoryjhp
TDL8kavr2+EMGPUrEZuN+hcL0hbNLHpBUZwsO0hCqVsTvajB6XIrFWt9QqyUSe27
5nWGPBHsWVGCeCye2gXqKYBZB0uFRHptuug4D/zQ4ZvzAMGcZ3ZPoo9xdGBJxvUz
dot1lxGT8/aMDYcN2gvbSgaADY9e4Yz4Qw9rVoSYAUcZcgqNF+q1qRE3BZPt92nz
uTHZ0S2Jw6TvqQJjfqkVRB60uy6Lzp8GHgCGvtUd+PUDRE/6P5mJQQYjXsnUPpMu
aA/TY/1YRndore4mf0iCEJEwgAC7ZxGtzsffEEHaOWvGd/GqLWT6XE70QfEq8Mok
jqNPyaFuR5a8JGwPOiTwpXtNvjFQ1VJeZcG6mSZ11AoxxoIJnh5B1+iaN0CedlD5
NivffF2RKU1SF/3sjGi7k+0sOjHd6NFfbKRvwCOmg8Dov4vvPYIsUU5HqYHqLPgI
xMeDyDAZSXLKFMhRddrkpfOcH95qthzcmMC/3aieuedQV+rJDa1NOLwKeYMotLzG
hZU3cjf4kcdo6WrD3Rvmofd/bv91x3vtoHg11lcBuEMAwN5hOz6yGKYW4hN+C+96
8/F4p7r8wKhLlSgTu/gTeIF8wgeBOJinjxcJb7PLTHj26zse2McvB3EE6gYT0n7a
mznCDgGgGajFAzak+Wl7VmBlPSu3hxxDMRYUnJafszTxFgKvPBbPH+SCrnk/aFT8
pT5jzCxZGOQm9LB0Jy0APUgneXeeuKqPobPiOIhDLqXOlKkLcu+2WxdriNCzC+ct
2mkULy4u/JV1lY51IIzIlOnZHIyAVU/yifyeR92r8QgfFYu8z+zBl2u2sbqvmw6l
GOpCYP9/XfF0Y6ZljMxsy0PsTt/4uMCqYd/qg0C5AMeW/50CErlJuSLLIpoZcgUo
niAH+dwPFUf3W4R1RVJCKiYckn8AsDjuG58qvof+rHVfKhW5L3Ox9A/ajGVqbLZp
RDW/xk9Tuju/kSlDz3Nbpt2ZQtb3ihQOsCkZUqMcisE7hpOBWuXxaB3/klIqd8YV
wAKq4D0Cu0itYTOhAY041rR1TgJCbXlobyWOlMzOKvSC5338Vgo4kxUfIKcLo8a3
ZdnoTrsL3aWpQpvnKdYsAa1+XTOOK9VEVtqRkKjHt21/WRwHdYxifYr+4EJEqAJz
9wxQMypHiHEFHSgW0zA8qfY+PQkEZU7Ubff1YSH0AULmDv/ZHBu7YUjTsnbYTTBZ
VSIjDrc2Yi7/51aarTgKXuidnnwf35+fe9VKl5CfYX+i6lfiQVRetIJLnlQFvJzE
mDLz5pRlsuWuKVBxa8vrlmgr1cWLEI0mXKgGz9feXjttXOaXVwDTVQFsZx2IBKrG
N+FDwNi/heGZEMCFbi59530/R8xL8y7AZt/YZhy07tgmWevJMX9Al/0vjC84nzOf
5T1fM+PgginRwvLJ6cSBz0xJBuDz3HVTxIPG1ang1XRSfD45h2uBUKIwmxnbDRQ4
7k1lpaxt1hAxL9nHOhgwzlIb2T0+MApbAUKYezpkCdPndz2G9fWpRtEmZPiSAeEa
+Dn+DertXXbjUSqGgc0uZNoTHvESWhbzcux1oK2iXVPGDMazaEzMta27JBHRiRgW
JCikNILdQPWXOsyePxgXn6gUxtFoO6VP3qJeDMXVCMJTvq64RNZUYD+u1LKOD+LC
7OoDE92500ZU3IMvGvxi+R8l8FkOkLKceKRaipAs0xUfZLqWBVlcuvkb1BfBuG0d
LqA9fGzNSGAouB1CPcHJDGPf6fzLdlvXw5wswh0TM8zU008kQeHh0LxubojDfG4u
uN/agu6+ub3pxupjHnsIJ05jw4Svx/0fu5x+pNgIV9xzS22+mo6jwCQZSz8HEbwf
OF190iEfWBXUU99Ul+6VA9exLZjbMBlKBmQzs7br+ToECqXFRCHZC+9QUhFlgEws
QyhWUCJYHPuVTiECHGRK6ORSA2dc6szyu7+h2qcol92pYM3d+3kTzw+FTYxPUcI8
eoVv3m2lktlJsc4AwGPsJeZi2Z/wrAbq6nIUYsfJMbv6H8KzyKlkMFIHJZmTtQfo
KFevlos/8yy4zkJnpq61fhiymNrPNk8dOJmT36caR1fJM6C+kuNOLayFPsTl/6Hm
SEXFIGIKaZFnHa5c61k5soOyI9fS8xNh6f4NldOl6HquAgxHs+M+jaySon5/+H6A
feVTZKJM8u/oplkiH8JUGHMHl96L7cNGGuOFhheXOQqlmurTJXNRed+COKwGY4lf
9ubk2fJWbr+3BSwoL96pa2sE0mh2fA3hhCj3Vq7yib7tP8hHcvOIWOqGvyVqhpI0
hFi6/d4W1TOL+fU1/Y1q9cdWfgYkM9R8AbT4dXn8lKV6VkJMNr6MQO7XxSeL04W8
jBvewVlJ2MAgRJ0l2hmf95qSP4E2I/3AKV5YHznlEgYKMVOgCZybqn1snN8l6Plf
vzi/iz8DaFw5hz0TsNN8jtU2VndRtJGwqRYZn8mjuXlGum6rjEeAOC4sMJ4+B10O
S1K7rYsnZ0K2+1g2ygiAopXtMwGLM6b45IPsl1FhQ72weURFDv/OZEKtGtRvDjAo
EXE3w16Je6Xp80uL9QxWtY2tcaxmrNh3RYYDw+zfkosDuK6FbacA5nSO18Rmzbb3
YpplCY4f++eC58RgfPBySeUgRPYsefQvNUm5STlQInW+UJNrWO6yo+9hU3h3Akk4
Z7GVhCxcJzf3vTBfEReWp1Bd43f6s2N8azULTLtqZCLFiNjNYojkYnh2rH6VxtAD
9UfO8NL4U+AhKvkDJhKCnj1BelLCc03qCv83/lMhcrAre0tnIH6fuFmHTIo3QYcA
49nfY0DfVkl7daOIw+o0TfX1aXCn9yRehprzJrcMHlEfZQAT/WIQkG6Nrryru+x5
R0JQvhloLtk8ZauPBIeR3xM5z96v9yurUeRmSUtGI6xYPgT/Ak75vVZlAC4+NVYF
m8hNJyueYKJswokYXLk/aRI7KNcH+D3wcSiy84Qby9OHKWwmBjmB5w0xDcHuQKhZ
9RsZzBeEVC5Rq+ePNj+uSOo9OBrFTx911GUhj4ziebUPm1V5KzVEK+rNqwVNytfW
ykyR9ggz/iR4RZZONor2DlD2pVP7Hgm9AKJ00ovp5ggjme12cxQM2msFVI47PBJn
NaV2+RJx40ipfq2n3qEe2ZD6gGrmCTDrpF/xz9Kj1cROx5ZCdOqb3nS8yELeBmM3
Pdkl+0U583AgFGYyS+us39bvXCDLUTxVT7rGAt17h7j61i1XfDpf6HSCUHOfjo1l
IU+pfUWDjT2BF2tpIeTgzvFut1T7A0icIKvu/KIkElcvV6yrYe64hgmnW6x8FfXP
/PeDfXWHevuOqMmO0EzzHRnNno1zsMbf1pEanM46FcOzuubAinWvO74eR37ls51O
WYrCi0tWHimaqb7DzR+Vq2JNCDgmjZ/f7cI9wjhL4Bf3YEPsXfUfwFSm4+89T38R
v/HUtt2PtRo4C+v2xT0QV9rq83/GFYvX7MuDDxPMU1yMxMf6VgfvLa3pMx+MxgQR
JVJXsfkZXG2NYZ2cvjdlZfaY3GbvPxiRdzU/JOc7q435z+g+1lKeCAJSIX5OQtxD
ugN2RXLK2ecor7M65NLA0mrqRH3r7IS5sE9h/gpoDGKp2daWA0bLjUfcUCUk+2Us
/PWIUUuPhaYySzPJlv9tnx7vb4GdWATYrkbhdbEVB6V/rOxfWL3DSnmNn++/l56I
kjNZFzG7WokzWHdFiVzWnWZrCIuisgJV8T+HZ9MQpp8U34w8HF/uc/F3Zm5kFNJp
H0XDq+QFdmTM9epHshY59k6tZpmN6UVFPMBcLxvSqx391sfOd/dOcu830W4g95SM
2JXzyr1Z+VXPos6Nf87KnPG9YAVC3bPRRKLYwbK3Mc5Uhct3zt7JfiEcvwOOvn1r
siT2j+o0m6pP0A9MBkuZNZULNjZIPaQ/Aom7Z3ySjo49wIj8HFO26jcDTYdvm6EE
xEnTN8umxHHzUVClIFY3OwFwm1Jugt4f/sLC80oAY8/Wvsuw8hrzbPMAuph/e5Mw
u8mfz7hHbaDjCA4d6dWsm8xq2xhqan3bTYhnYJpxOEJ8N/3rtdk+Q0fbXB3Q2lMV
gUeK4R0Og1TYkx8oqYTC3gx4tT3xLaaYy4YbrTzts7AyqKBkjxo49PN0Vbrlm/Al
pwPABaZqHUOqyfp4Gh7YgZvv5TL0NaEOfM6KLjKYONUr5n9E71qHPhciTy7Ez9/s
LJ7X+hkd75jRY/RCLtsNgGliqRG13sdZHhUgQt7rZL43rrC1BUYyI46gIgiIhLtD
p8/50TJ1sXgt0GFOe/QW/Q8OhGbYW4IcqFCA/bfRbfkFAjUOH6UX6ZnFRePWyQ6I
zJxd7/jC+KUoPP43XURLnpGe46z/WxjtgeGbLWK7Cb1clK0FxJuRRqTdsF/rvNxP
ADVmTlY4lRc1aLeSnJwJDNK3R6yEgvgjoBqWipJuSbnxq63JBSSImxCbCejYKegJ
dNf6FS33L4dNcuQ/QXCyDub0dBzxIoVGmb7hGbeuIaYmmXSesPZVO3UOwk97yhzv
cAFAhzJWJKebeX0/iQNPYJv22Km1w1R0eiN6XJRmnZNQNFRjoS6QwlEc3QBlegsP
H9l0119nXdiX0B8F5pC+zJjwPHgdG6sKkE1kBsHPAtWQm+be7HMxOVsnkOeKyL+Y
lnPCFSLYunhlFeenGN7q70rikE4a34tA7a3ya4otfLlOq7FuCcG1UlYsrR/ZPl3o
YIv1QF8R/V0TdTAY3BIpJbf4D9tVPOqcwc+mwkGrtSfDg79vc5shGWkQ8PBmdtZy
6yv2DQAJ2ZWmNnd6mALVXCoWiScKtZyMqsxUlmzkkdwjmDpGPF7r4TMg98VcFTVA
5sgw13d2ZbPCmf83cABeVSOO5M57nY9Y3AkNnxHtTjiBaImoVAeGhKIA5T+CjEvh
NzAkftWwBlKnJVrjAv37tP8QM4oYPnpkwc1XVuVRHYZa6BhcQvjWf8YBt5st7PHm
34yc/lnTrozibCj2sP6FJwonftyJqWgUUbpEmwM+cECZ6Jet3ywM53ya/jekqctg
kUgox5FiL/io7z2aUz4A53nH6Kc1ABGQ/uwqqBk30oRgdJVKyQvlRCYcqYd4d9pV
fRf+EpPrxTIk0dx5KmoOVEcEjpo8hw3vRhaR4IPHPQQmTzpnqU24w6apuDkMdYhx
YRWB3afJDzVdGNk2Buw2r6rU7FRV+H4poBt6PPJQyHPY7v9teKK78y/N4uQds65w
wEOBSglg1pp5SG82VMhyZ8YiS0n+UFylX21QGsSuu+iVk3iE0Jwm2cm4nqwufzAj
rwVRnM1O/j7b/MbC8L+tq23Gs2bD9gS1mvWTAGtce1/oh+lwRxB8at4h2rEv28qZ
yrMIas17mEE32o51o65VD7FIwUBbF9xU1mrt4+tAU7Eck0vBU0szl5VRHMSq4xIR
yjW1/rS7qR6VtQO4M4kaHV11AnL4vQU6ybFr84kMOefc/WoIJuizNiKrNCMV6cOF
cv1cadIrEnXkClPAAhnTWhVmFHblqUrjnCRQNgP7FJ2sX9LA/z0GbgQZYzOiq+v2
wYgTGrrE3VcJO4t+quO34SLIqmSG6s5yP5fnJhQgaburtRZHvZU3MaOxylmJHQFH
gn34tjtMyJLwpwdo7jEGav/TQXMucXRJeWVHj/iY2Fk2svENHOF6jQLYuptWWf7L
PX2pIUWcqdhmy2H4VW06GpfvGH/ibDQ9FXU5elfrjM/I/zdBMFiZgHHiLqhCiM1p
HIu6g2eHdnuLd14PEPTxdQmBa/4akMSetJLGvmaIWJAca2AgQDtyk1IQdejWVxCp
qmnOFK9NfReNOIp/ZI60QKqWuSZNNs+4Wl+HhxjsWNMTW8+/x15Xmj6sDf1SWMU9
oKQdlGZLBk8r1zc0X4Rbri++aSxmZPq14j3aP20x2/x4k/uXIuq/RSmGbQdQ/9O2
fGNqRWScRbJQdb62IY5sGmBgiTIjjnLbewpo9b+17ftojIriD9ZqPQkCrI8X+AXX
Di/ZxpyN59E87BNnNIvcJhQ7rUEn8JplCLS2Omagd9zdqSng1h7LL55W2PccTFC1
A38hm7JCBgnX2+79pPRbJ6L+2UgohoKRrGIligm/VPTZXjq9VbDsIlUg1/jECbUf
E8Vbo3HxHWjvgzLHm6xhJtAKhw6iE1c6cm/RQTuDvwlNXTKNoGh182sFS9sifmmR
Rn8rmBrJt/qTkmfMjdqhHcLIRmUDqlEdvyM/dX9ZNyNGn+SZnwNPouzaj5u+2jHM
6+2ZHsqpTIIgYRe/Ss+srIMUfbQMNlWJiQ9qFBM83+4BevzETqUz1u4ZVwIR88Eb
CyzF2nA1Iqp0SMRzd0/ogSIjRn4d9/dN6SkLy8AFJrlP9crE1Np5ZSMs23VnSAyR
dd9zDYaXbFeGzDNqu9JvBLf/PO2xVAGTmXF8UjkXF9w6h4N1REsso+Z4QeAw/duR
KvnlL6Soy+Fb6Jh54GDt/JCWMYQLjkeagMvy9Plwx58K6OwiSxUOV/hbjtBc+qWl
1/2GL7JGQfbgllGoBbvMsDhxVETttm/Ou7I+fkopcnIr4JCJrKfEZMPNWdgvGkuu
VT3Ro36sro2011Z0qqwG3gdv6HjKdGaO7QdSX+wHkz5i/RYgPZHinWOpEQEIm2Ga
2kZZW9J481zzcxwCt14ogQx361rrLd2YMmoEN2INgzAY7okzgyGBTthn0vHv7j4m
FD+G/EMYvCRKS+eiCnsuDzT9YvWyr+XYfdU4RLDjkTgKhgfMT29/y4uA8rK1rmxK
mOzT/tW50CW6HIMQy8QUCRwNWJNCdR2kU7g0BNcbHW0ixcSBN7qAWs2cm5NVjPk5
4GT51aCaxi8BcuqYEyNp2g/zWZtU21aaMaxZ79cRftExvHQj5JZlcCASoiouEJC2
o84Ichvw1Ja9QdacGn3BuRfIzVjm6PwrgmYgOIAfjoU0sOCk5Ks8oU5MyDs4wvmy
Mjbi4NGus10vqKrNutjsSKj+vjzWnqKF9xrO6og/rMGkqteqL8VFnrDC4a2kAID7
cClVE4X2M6cGGKY463BtMiqJHv5c5i713ZGm0UNJ2F6vNicPoeb5OcK5xD9lxBDj
J7q++iJ8akJ+51ZgU3tRf7doePdfO9Br3AMltMUfBebtaOMk8EJUaCu08K5xeVby
XrSBvklY/SGzBl+sZQyF3AEE1/4mzbsBmOifxXhrX51EetMfQ07oWJ/UEPeHU7Vv
I0em3Ev7YN1xK6v1q1lumCW5ZS+kaulj92S1jF8YUT/6pg8RwjI8Hh8NOt0nRf+F
vx11qUOwIkgZd9qIHkmiuNvnbCDHuaPezWh2AzgZgaVWlGMM5TUOzs7QvEuSHByw
T9lykdE+SWkOUySAWAn1OIQ2bP1GpNi1QNO60ZDewoCDdRUkKtN/0sIEzmAQlaM2
Q1pBKBGKexzmaXTo1i37gtCtzN/s77ssZjUheM7o2rH3PeyK9ZI5Htnty2w8QEt6
tbdECbcVI19kOmjEkSYalXqQhDc28Wq4TOB7JEUs3J0aSapCxgFPzZpM+SsDWgdr
sYjhPKBxXFD4TiwiUlU3PoYLLPcekAqcLJ0WuZiMjf/M5woPS81axo072ge0T83I
TnfxPaiIz+SFIImpTHUSXvAgME7//B49nBfqxQEtvXURnLjmTab8xXu2HbQgKQ5U
wHGmw1N/CoKy1L9SAGllwz6HAQcSeJ1i4hWNGeyczqbDU+5QlCOvj8DPmEnJI47u
eeKOGvGY5fhm3Sb/Y5IpinK90DVLmL3OuvaSCQqfSYlbGbFjIeWcvYO67S74+ZEE
cuqa2vhkH6DMzZCxAdSpZ7Tz7MF5R0k6dlhdwsnVWv1qKQAYdSYhSHS0qhw+lE1t
ttqZZZjqHPHS75/M7osrsq//lDkT0VuAI+7IhUTLi0+gCjuYamL8dSQommoNM18i
0GZVwE3r6PXhxVP3DVP4NaCjZdzXrQBIl5TN1uEey3ksqSL28l18MEjWdi7ZRN/j
8nnAS5KnWCVYJhQGczvucpUKJUBs0kj28+fNeAC+IdLsW5pL3HxqehIOmdXM5mAy
qFdCNpVezvcC8Mb7KsB6K7ISOGHHsFma0BhaZKcmebR0t6Ub3SNdZ21tmY0GTpxo
yS8873FlTjDYK/XAOWMeZcYEttIrBeamXF9ondNmY6vfJGaZECrzEK8xodxwNpHi
MIRwVKoXpEvoqxThdDkGquH3RyKZXSJjYf5TJpMUjlZbBoTcLtPNA6dOfg32OHYG
ewmW5JhRLzyCrKVVqQn4u6UqMLUES0wX91l06jtd0TkaNgW56Qc3tEFp+dkSCKrV
jYbQdC5vgAwD27FJlTnvocGAPjPdeRkWcEtUaqGYoaGnZawfgiluVdNXxgAYPSur
fBjOHyHtaG5ylY2jot+/2au/Vnzxb12jKvhZQLHoInvZYF/t6qp3/uEoiYKhizhC
LQNEl13ASzxoze4Fdh2U3suQ0oXWfhoRg/GBvNqJVoXN04rNOrAobi6FqwtQyM64
M2GAtahPX2g3Vvm8Y8s5E4lVHQcA7R16lhx5WUhVT9exRsQgETqdO+Xa3VBdGtTe
dzew7H9NXHb2iQW24JD2z+JdHdL54AOrPv0/vuWdIgiB7vz8NNH8Dsp9o0Js6WIi
b8g286o7w2+TCubUbkaYVZb1DWraep+cnZkcL3meiBDOuK3XUb+Pro9LspHS47ZB
FwgZady8ceTC+C/j+EO7VVB+ma2gZ2XFypAJt7tdd5N9ViOcp293eJHInnfveoWd
EEppF9GlMMPWRMClZKdsZFdpEWgXo7yNLW+kyRnrjN1QUh0KJLtDAZplTbMEucZK
T5x85XQnCe4juPagz2xnP4a3JICpJzpa+py8y97dVS6Kcq+FnjnZwQUb5zPAVEbs
7yJj6oh7vKMh8Agi34wup5vB0Dgxuz3Z9mC/bm2G7PWRbnqGP7O4bDLcS4baZq2a
7+U6gLHyFXFJ1Mdi2JIOuIT9g3JJC5R6i1rvhhakZ94XdvJBqz0XkqEYbcPjECQv
xhDZfe0hBFWwCoE8/CZluEswI+Ld97qnzQnX9vFcT3wU35W1h2Q0aGowcgsxy7vL
FH9i1tyCS6c6EWGZrFNsoZvMG0s7vsaK4BuZndizXiUfWVqj29AF7PgHP3+E/SKY
y7/KplkRwLlD93RW3z/hvnXDgsK2hjVb7AZTx5J//59XxpPotRBfTi8QLLLUsh+K
zHbGloLZgFy11/Q3b3eFn95fKPVSPDrWne/Iy9wvNFdb5Xo7ho+756kckjAJHwaw
4asUfLqAr4B55L2q8LEZMkjx/SdQ6cfz4EKEw4D5MtxnKUAc+kyXsaJ9WxI5z7fC
aAmo2wkrq4jyUeBWPnpt7z5PRebliB0J5XR4VJXpLUmEBOZZMFdlaHMBGlpJVmaz
j55iigX7clTk5SajE3yqE46HrujWcdajMExDP/fucdZHqZowLeg7ZISPn+oHxiN9
SG5VW3beRE/AUUbSwUpu4ia5Ub4WaX8z0+pUmmtKEkzC5cdPVH8MA0Xv+aOcObis
PhmLrD/otQGImfBv4Hs7AScyiJJrS3RMWO+SXsRltrmUj4l3sR6CNvf3yEWbV++s
d8KDqY9XlxHDep9iJKlnoyRcMy9Wcu25uAzniRPD7PGQh7p6BOIBlMJKEMSbjkX/
xx739wnFGeeJaATmkzg5khCeMPppSqe2elNLNlsMpNh9hMSoeGHgAd0khbI7bR9x
BRuOIfUxVO4IU0601vjwJYvyh2RgDKi62Llq9WiW2biyPL6nIqgmk2m+DzSbU+kI
0Q0Xo1EfgE+Sm3rEadkTNl0fLLQohjJEq8mtbikEDWXiQJaPEzCdf4A/me9jsWz1
zYh7miwbUFACfBJlHq9EUma1MydzxOy9Tdl5TX5EOuN6GUPQX5CHdt+2nQfzMScb
5e/fy0C0l/KPAS4iV/PdU+NnjzcwVYDQjg/NXvfxpKVVWMSxUs6TNr4NS1PEejF5
e5hxpZWwBXvfbadHgOicEgGmOqB7DZe9cM/Vbs5BnJzc5ERlPuq8juTNBmEMPXBQ
nRUv/HwXJ0hbPrDzc6KiF6EZss8bQsHUsmKwRsOxH95AHUW9PK/88hhly7zliI3S
Wspb59tVlyw8YLov3oQDn8fO5hIIVzIT7Z4T5r+CYjEBD6K9p+nFwY8viaOKGjEc
W2dMAxXKTUE13zbKhK53ovvNcXdJqvo6akj3C2/VO1FJnt1MPyJ5cO4+1LWCRpuq
x1qsU7Y/giS6hQJAG2MzZF6hhGu/RgewkS89JMLfqjmKz43Xb8W5+4BoPa5tLt0e
q2HtcYyH2ASfqXR2VL6BjTuqnXgbfl4ejx5HdxCCh5umzu2rUxtNODdJE4N7lLPf
N6wsnCCGmGDJiha8UhDd68iCTwNbw1CBwyhETSctunpArDFEaFQkCRoIaHLpr6Wm
KfNAKlpAbxImTXGdaVGX1LLxDzy+uHW5RJyy59B8MnT+BI5GA2bdc0xUza8l2BxQ
50E0rRqXZWCuqxjHMSSjXn/PseENYjj0ztyri7cvQA1JXraRuYuNFew+FKgxUkKx
eFcW0DMYMuW4oitTqUxwiCDWIXj/hZ72IBANgSJTmbARxnp/BAvI1k5zS4ccMNVq
6YqIkX8F/sbQfyOO05MkuIRYFMI824S3n4av3UUXLEs5XqwErjOhMan8449JpP/7
QkLXrXzhp9b9hoDYFhU439PoVpFn+jJuCRDmmG1n/D7I9zu/HwYbMRX+0PZZs6ez
qupq82hxIPlC8SQ0rmwm2Oa7rZWlwDinxY9nTtIwwk4XXpwiLrJBQUy5N21zHX2w
kLVzqmuJR98P9GlLDznjir5ekKFrAQeKEGvfij2INho9m8mODahxV9oFLfPoTn9r
3K0REn8cLeNuVulnOYAVNgxmITFxXaoYZsJkZ4Kkxx9ADGpQ0yjLsr+u/ffH8E04
M1CawRkRU/UTrVbBHHhEUgNihQQBJtg5MQki7wGB6HUafQ2zdYck/L2fH6uFigbG
OL39w0ABbCx8sTY9DfsAFnSMY2yHDg3rEba5kJDElKVpS6m77HKOK04W/0Y3BPR0
D/fkQNPj6N3D7FzR89hZd+Zl4PoggqjWBbWUOZDYoDOAJBxFzPwPF5IzJ/XPvBTl
rPqwCL52AB3GUNS1RxHawO6SdgeFFl9oL9+j3qXzbj1mHhn7pQGJpQEnwIRyH4ML
bdMZgbdYtsmg4WEoFbrViz7Nj2olJe4LCDCEskDwrlfpit879sxiiR7ceRzo6Svj
LQeTWdCxWd7cFo7BTTjMRsNbcA59FbV4k6LLjXqt60PnK/uvcqzVAqNSM/KTOOB7
0/Mrpt8DqP/n8tiGGZkOQcyMgcHjPVBZtzJLalmmGlQSM7HV42Q0LGiIfoNqOErK
Rul2ZOSqZNWnRENvIvGcNi4OyisNa0sIJPlr3ALNsAMklD9zY755FsVoHNn02F8T
unpo4I3Co7RMxwvC4V9uuB2o96Aq8/5aRrnjzar4e3TSsPvFtNr/HBx/lPWrXHsS
T4Np0A+ZvekovnbfhpxOdMAkFpC+FEvqIf7U2eoAZlq2+GcfhtT2vv6us0FUq6OR
Tz44HeUtAs9yykXXo8MtidpI72O5B8hSBGMgZqbkXtmCUrTGWJPb4cps5bqJU0/B
zjR9Da56rKcBRIAJp7r79Ia6ozFcLwZKN5o+1YhdgK8TK2MsUt+Y0jXJdw7H51DT
OjAXgSElYtnyFj9BvWJJliR2h+bjwZNYQ+A4LU1mdWNhItjzARC9QRoMpiWx9qY+
/RHuMg0FhUdOqvQ5ZUS8zoPXRlaMS5XEPo9QNxBRe5PfTNON9jmWy15y3wdMLIcM
j3b81Sx2laAiBotkcfOluEhpRVYs4cpMYy/1qtAptPOajnkhX+Ucy4USqBwFhX17
RI+wJviOD4M9PulOZA8VtmpF74IzK7ZfbcFa539qUOzR+bimbDxAH0OqVz0G4iRC
lNqoX5qHK0j7iYxfhoa0iSUc9+zQcUyp83rqEX7sAycLRY+xTPUdWpK2R042JoLc
dU6v4N4p18Ctlp/N1fHDy7YZ9ji5afZj108NblJrwSX6s2DPMoI/ywRpw7ewz6jd
n20Vhh20vU9AthnKqiiOEKBKN5Z+2/GUKjuwMNyV/CfqNtLVhwv4Y3CymWWjcBPY
R4OCMoejVkjn9kNlehvODPZwufwZxAkomAWmC/8GvOVYwgErzDbUZ4sC3yX9Dx1n
eVORs9wog21nksWEb5OMiitxxYHcX5qf7kc5CBuAv1bv/wpvbZSWiq1DtB88ixFX
dCbbhQGl/DEZ9wbLwlIOd5uwbwCRxvVqHEfq3TXo60fB/s+xy+3pjGtzegoivQXd
pnFWe2KCeuxwYTVgc2xWIJK4EjjJgxscZ9F3q/369+VePQxuIsiLxX956RYJTVfs
u1/S36QF/sJIuqGGP9pWgRa0j6sRhHpWBHjkN6IukcBWvFsoTCzqQPYtPVFnIhuC
sQJDI5lEzClt6WYmzTx/jb/QnuKR+ZOkc3tf5ARvDcrly0c9P6hA1H2tsTyxYRo+
2j4l/ozO9fw46HztV2SWCk3D+/pyxmYdKJaAjKGWszLWl+PRIXcj12k9CnKHTqOe
rktEE5wnUY1/+h1ayCRagddOLSDx4EMsssJeSETS/78SP00VBsQV/pB7+HPv7hrp
3kPQ1W8zXXwxDKAwWDZY9/A8afBNdfjLcNIIieRXZZE8O1nhouFdbEgAtP3If8X+
w+9UnFiSHCNIN/gRd/BZ6uUB72/h5Rc4GbpcAlFDMzOWOjahdbTGg5N+ajcgbizD
wva+683B12CDBYJl2XifRARO463dn/DkP4yx2H3QF+bOh4Az0htw4s1LNRKjQiEx
7cY/I+V4Am9L0U/VP0losxjmWN6+UypDLZqJjpHZNDbioLiTCfhrVvM7r1tQL8Fu
ZunRgoF5Km9kWx1h0ORzRhLh0beuKumSCki2Fzfk4yFEeVK/8glwPU8ClKgnrDIm
VqOr005K62pH5FRXTcV93jSCxdMNCUHs7nKlOm7w2HLV4dVgf0t88dqNkAKLq8G4
vzEWo20PrUeSUIqfnROQ5XxXfkPx3Bp2junTxEdKBwj8KBECDWo3olZT0asmgnno
Mf1PxXq6sZbv2arqQV5oQt+MIENYKgCScd39kNrpDOphjcgtKwRggZ7MGa+bCaom
ADZCs+km4kFtYGABofVI11fC5GYK0iLbgOP1YEaVZQCwO7+mcD/PcoQGbG6w1uWP
inx56HGF8mQ6VlxFaLWRi16tbk9nEIVU5aVWaH9mhjHkmreCHqdNpOA7pFzq+F0v
4x1lc9ST/0y5XzTzK6Y1CEibvdFvGifRgeJoof+44ICw9wsefIi/rRqlSWTgsq8i
anO2dwxIOfs3uQLope6VJrG36dt1pKLkEVzNkMjJbelJzs3QtSsA2bKm0O8LwLx+
D9p+6hdF/c9s0li8wcWDESfnING9pz2zf6anv2mzsKIAqoRmq3X27lDMECTQllZM
yybi7y5rmn2RjAXGzcUqol2+hpjG3M9Rf+8ORV1GrhdPOYzwhRNK0LXWMCIpdycf
dyvovM7lBK3xGyPcjdEgNhFmyKcwUuvb+WFsKp3IXi0hVtbqzjq5QBH6eNhO1Jc0
ZiacTXW7Uad9G2QdRv6jBNGoPjSnqBhK2dPiU3iYf/YV7FVsLdFf7QCQx5vf1Oqz
QPec106Ah4FY+kcmCsL1lw2ZKWEBYBBonfziLXMQCPIFZirH1mIm2aZI1wTEyqwm
N82qOdl5N9Ptk6huM9MwetWRvIJNktLJzTTRfrQXGGNO/AQDF+0o0D0FahjAYwgb
vvTqj7qFbsm0wJmzK9hEGEI4AtKhZQVIMvWwS3rc8v9kZdrmxd9dXPCR009RHK85
wVUdmz9TMsz+vHhV2WYL1lcL22N8ttsfU3uviTW32ex/c/iu+tK0eBl+lmWpmxBv
r8Sq+eF77+zwHj3b+NiUFKsH5ift7frE06MYvdI1S6F3OdmJBd9MnKr/SAEgaQHY
AM2IxcSnCaubOTFphCo2XnuyrWe2Chqkcv0q6hZp/D8YmytP9ExcsqWhA4IVFuJ8
ZLcZXoQL5Zjy7Nef0VmA5fJTXAW3sgD2VCr/pAgdb3WoXV1ihhNSmrPrGSbewcAD
lxiuhuCCX3aIOvQeLZ7a0bA35pujtumozF5XO3l/LUx5pUOoPSEYEacmnHmSbC5Q
a9DNAeb3mTFf2x8DDgmYL21Z2KZfxkrWzHmkd7HhF/PnCoJg6c9AY33gwdIAtbAH
glPOg+Tfj08Y3h+D6sjizRHg1Am/v2DKRZGUsruDIVYpjNtG+ql6bijlnVC7gD2g
gs6LUapoNHUZJA8FZucQkSPdMwds6yzHdGzw0gB2PeG7voXJqZ6/iuvX03Hl872J
apVHhwSLY+JlfDHaFrCMuiC7BfXO+/3J69lTVpjybn0yyufYs9iYRlpEgPrGncLa
jkEyhj8PGKf8b521VVAlbu5M+k45c+wFzfC2O1pKABNQxYpRLb6EBw4ugviFfR0P
tzuWzPH6UB28zpHVdAKBatBjLtHZGj2GlFItLY/Y1XmKuYUgRY6ydeMsInhAxPr6
wz1U4soU771tgr1LhYJtWMspQaYnggv4pKszG6tOC8aY4V4f+3xWJSlJBOozKeuD
KWVe6x9xOzj8t5iFbozmXxue1bl8i0DkRgIAZyxUo02+alwjAsxDYxrCzbW4NvgG
yFOCZVC1Kt4Y1I2HpFolNoR88ZP60QUZCLYSWACrwsrFXAC8RDeSjP964mXD2XuF
RL14y9mXhQzccQT1QUoomIMVe5Yi0J51Eyb7ec+H/a2IYW+fHjO22d1evV4OQB42
hd/5d2SkG4Rerd/v5G1Lj0uFFXAa+MipfZwBbs70L6f1e8PhtdUB6KBNtMMLLOZD
cHP5w7cc7p2PyWjdV9SovRq9pSeIkI7i09ovZZMe+egdnthnNCLIc4h6DoWZ2A9f
5Arj4tbdi/Hch1tJK1eoJ4LAAy+LohAYx6VZEUX+qzBKdxOX03gR/kZYc8wa8t6n
mGprDwe9+1TMy+4c3lNJ+wmRf2ItoHYjRqTJzg4YZxyoLS5ajZa9TAMCITq2WUfi
7ivATTA5inwgE1wFeBfoYGNp2wMt/k1BHJ3YLRvkQ9wJgi+WsJYxwVxPDQPMNsyM
kJkdYQZqRkIqm+NQ9UmJh55DO6UpaTDObmB3Uj5yQzsbwGDBf9vVwm9PfqbZqJtk
mT0aPmGCb7d623zTEzWJQFrKJ/ybNKDWOhBX0yZBMd8t+rCHQ3gD8T4hpgr1EI/5
Vvu+afkgoQ+yr2irnr2fzAwxDkh/ni71ZQ93ZMMwbUphx5wlpbscG1w+q9mC3DZu
YFYZeP2cxhA6RBZWPXyhlQrbkBO9p/VqtfmZloO0U8TOB9mlULwJqz+qxMnEXQe2
VGXQ5Zb2FGjjvoZPQ/OmpAt3C0qp5H9hYksqCVFPJnv4+whh151rnovjnZYeGGUw
vDibDfX+wuscClxvD0qp/tEn6RNYozljGrGJgELh+PFloXOGO1gvI25tr5Gyhdx0
fmwIqNY8HhjEea6zX6MweX2d0E5tJF/RQikVAUp402uB49YL/aHQxLRd5ASOFe+M
VICFBP9K4u8+8nw8m2SuED3IL9Uxn0W1/8tNJ1u9FvcX3XXFajUoUXtFZRD2SE8j
THPNaRdAuoDgZgB6+sxRjhv13EbOq5gM//J6ITA1AzblbBgM/06zkLYyLblokoOJ
Vo9UL5oeYvzghj/xrV4A5KVdBHjwxQa8oV6iZQPhdq2ZnAbZNqZ0Byu/geuHk3Lf
c9uA1SPEa+OXoUy1lN3d09u3F/Dci3+j/EN84CLwguw1fxOeDd3V7hai1YqpPNOX
STMT0266qlEz9c7yBlvcatfYXIh61Z56zAIZb1J0c44cM2vxPPhiSs4VA5ENHQLu
FynFBYvK00O9qkYjD7fpswUGAzUHflvixaJIC3EKt8P339AH+5rl6Aon5XxPwFTs
uWTBVmXkDbJ6tqbQiSFPemoEX7kZJO+e2oALluM63W8Q6ZJRb0usFsGiOnMS8qM/
4vCtll5VRLnP+mUJID1umxr6MT7BlH5EYud7+Z9UzU87Pn08bXA3HLg08eotn1Ze
IMGdq+E9WfoT4EeSM9kiAWA2niRmU8MT2wee9XXEVn7Btcb4+Ve/ee1bxKtWreYz
f2EOhtCeN0tDKV5RNk+SSBEyL5Xr/VSwmG8V5YnXKeJ1ZqvTCxCFRk1lyEqxBcFC
jK1pC8GmgrYx3rfgZRyfVR9OaW2rncLPXTlhvOEhGEKxinwbiV8penaEzkvG+q9E
JKSC7idinZylomwdt9y1kL4yFQjfylCuFbNRTY6GeeMEIumqf7sFuRTmgM1vhfMo
/CZdB/PLt9wTX3RHSx3aZB0Pjk2FzCYvvRUAN2bOXxSpB2KbTz9ad9yHivvwmJxO
j35kz48yeFVjMwxS/7Eda/Nzw9I8wCp+Z/kT0ongP3VVAq9E6Gwvo2Yv7xJW2XCz
6m0Ar9MjAY6n52vYa+0sDb3zhPlk75vvNyRb8mm5GxFmazmn4XkAYflJTL3v3Soh
rtjidNxgkmL6OceuuuuHpoTBvwMQHvS9QjoRH43VAjn4HYBGTwnSCE4EO7Le/xw6
54O21SP8baso3pwpjbBepTMR0c7s+6/3oOgg2ZyWtoL9LNGRzDPgDKiiJYjWj6nS
4NXDWmNsJMh9QbBP564AlThkzsplqtQPi8fhEN+BxIpj5RKc1JAMJQ4FryD7QKlh
hWmitWSMDDA8LK161LzHzz01x8V33A1hJR8g6TupE73S0BeLyMZhFXPNoYBgR974
6lK9nLzOwaHFk6EsbAraNPX4BKMLIqXOT/6dD69qfpCkBdMIVpx268+ljG6Y6gHN
Ir6r3EtqJEXwaNoW96beO3yD1y2soJYyeOwN9deKP64ahYVLYWkHSwvUoKUj6RoF
/+IX+8ll+ViG2hwhKgbj4mBfeJVcHHhFojnpOQ6hGSufzgoROe/qNiwAtpPTXY2i
qgZ8ZWPBVLGdHVBvS86RlRwHIHil2F+qQ3D1BGCW/po88M/Cfp7TRX99XEeyovim
Gcv9MjCZZ7fzCJrJUSDdYFysnPM+Sy2/LY5hQs4P11LUk1D/tTLfvhUSEPBfydAT
GO9w1iP9k/NiGO5HVq39KXeRVjzzsfMYnKIMzfoCT+eeOtGDKmPpdtaXY46LojxP
SYlhTBtVk9jDd4l+1d7vWn8VugI0jDLhURjRD4rdAuC2x0U7HYh/7YiKcfI5q9k/
MOLUEmeOwV5RJpi5/saGguI7KPTr00uw+g2jnIhBQLnSJd4U6BQR6ATlgw46Pm4K
A7As9cilgqFmrIp2kwqzHUgGRi5FtEBpdOpKLcIDsFP1m73k3vLrHIo6knl6FDIM
t9DTl+PbX1ZFlgYqAq5lA7SO+pBS+qnQGqLWBAtdVtci3rcV08K+gr/rPSR/Df3x
0UzfOqpCJjInKTemSkSW053xDSHlNU+24vp8bq/sFRLpUh4yKocHASMhAslyjwug
T9P6fIMiH64EOcriRi77ZIhI3indxZVDAPoQqcyjyxAz6F0gTCsBrn+mrPtxmT1K
G0xFJRirLRf5MT/UX4ncFfnCR7vKy474WqCLs/WGVq8FvWNKCAIfkbiHJI7cwyn5
AGe9Vsehkn8o3kDg+vynaGnCwn6VC1ERoJt/t1RYoFDhnrgwF0Zs5SHnCjbt+Xa0
aNBWZm7yjoJ2aHiLQsqZDkJuAsn7h35xwER2pe0WdoUsnv/16pbrTAv5AkJcB7/l
OCzPY6JAUShscy37njOAhSO9rRvr/R1dSP+UXdkrddrwmlcXCZIfzrdp5MIpsSvI
eurd3UA41uaAjReRvZZrvEtB0WLXzemTS1CD6zjPzrkzm+PSNZbnUZ/FUepZmGcG
12NHpkbNW3gA9iZ1+FrJu5TWyD4tkTSjb2IHEAKuV03qvxEMZVhfLBQlkzdlZVmA
1Eev3D9uonB1HtdenS/y8fTI6mWEnqneOHxxT0boYjBNHnMDoPkpVdXuPppTRfpK
ndx/c7CS1TEmbRe1sVYZaiDfsL7dBVu8FPhLmbeX0EnUpRMrEzze9ti6HXZOFNdN
TtxNnTw7dmdBNCJ+WtdZ8cJkx6eYCtWP+zkaGufAzTM4pfF+v+VBte3pZYHBh73W
R2Cb/3nDDDx+11dudAD1Eb4RYghFTqowO283ZuYm9mX+JNbnMStL58o2B82PMv7p
dvGwV8gzOzZcgubSXPPKc5NCvS5Szw3kXgXaEE5nYBHzBj363rKlVh/G/mjOSZr2
d5mdgG+L5hwAAGkWQncx1JQ+iM24+45/EWkKkeSKmAz7PKohL74IQSDHaEoL/ppB
e8y368zxhw+Uit02yA3AKeabhjoo9Ipt2Tw7HOg4VlKku1AbjBBiajmzkpil3nRO
eNsc2nqb1rqxTyQOpdAojNgs8hbVkAVdMnQPDuO7HFvX4CHMDxkxSCVvBGo6E/Ym
/8yxI6Gpd1XfgJ6uu7a+m4FzyUVziUUZ77UUVXADoqHSSY2ju2Y3GoABxaONj0Gh
8QncR1QAJBYs2sacnCBQs0Xy7xlfKB8Wkc7EqzxxXQztb4HTT53UkAapBI+8/fub
ddjfB08qd1XWscW6C+0AcOokU+JsShjViq+8vio68Z0QtKKFMr8EnixjPxHPqDpl
0FErz0yFozkqMmsQCUmd8sgvMAcXhvuP27ILSNrEEb+BLP+XP6Jp7kRdXpkxkLRd
f6pxsn0ISTkeZ02IfsSp94sqP+syHwiCw8ffqyy66hoMuqRmrYjtN+N85yQRoFR+
UfuTTZ1Gbg0CdMpEjkLIs8MqmXGpW/3hai6zXETJVYRQAahoxaTLFtL8G4h+P3WQ
zjp7DafcLgi8b659caXcBYHrMVj6Y7qVss90J/lqADDJpR2nTS+M2Sf51yhHXbKi
sQlDl9u9vk2Yqt60JUPDLVzuCim+aiviYevkMdIl9ftc9955BbU7W7ITvS9BRi0/
kUzVqGUkzWnIAlbm1i1u+w/50354hS5LSX7OAniKmfnvtUBkQnMZ0mnH4Zc+0Az/
LmGO1KumSPobXDAzrWuY6lkspt/xNqdQ06BBvO24x1kcEbv6R6VC2CKJ5XRLB4E9
uJblKUF85R1LPm6HjOOIaIelMfHyaslfoUBA4TRgc+YdLbz8gqDTR3YqNinhAoRb
MEqiglpnPiAW4pDFyTABmZj+klxtGmyQTJYtouYtzBpIuaHU89wS5WFJExYqohsW
txAzF18X4a3bfxmWpZjR4JyY0n790dfZY6BQltmEZG+z0FBjeUebJhxGRIW64wYO
f7k2OkaZc6wwLEj0cAFAHVnZuh1+ZB+SLHlB+/eSSkn5Fzn9em5O8Q5jmDuqRzLa
L+6O9zDJFyi+F9qpNg/6FZH1By/qkc9hZ03X89Cxa4urC6dxXXLzhVgQfEZc/dW+
uvLpa7WsKOq/hXaKivbvpdEwZm5CF5P8uEq5xKM2ja7/jUHLIYg19WD6zsTLwmlA
E9G8R74aFpNDNWaTrvVR9E8QXjoAmmwYbiXROSIfNgx7U0S9QQXdmrMm3PAiq6Tq
+HyMuJFyTVzUUtsQIEbTt456olIDj1rWiRBiTf9LUB0jirNanal0HUHwQ5agQm+p
g21EvnkbBaEOlQm2SS+l9Zhig5K4vfPhItpVe4htQT1QauE3rybib/XGDU9W+Xh8
k/uGQGbSXQ7pPwbFDzDVGuN6s/MN8BLcI0eCFUjX43bm20mdLD1PG/WDbouYNecu
a73pqu8siOQ+krOIKSFjlW8bm1wpNIqANWRGlWeOYIHC4d1FRSOdaThro4Qp/H0s
rw68xMztg2QZFAAjOh1RKZ9yMQJ03XJcra89B1zh/nRn4IKF8e6ggk55eUZ5r7ma
rF0sH0cfcmfGKqzbHOt5JlA9U2LeyWI3k/Ym6s6rvqrnkXYxpDGIVXRW4HBMTF/B
iTcy0HKFSQYMRj3i6hNlvFwHDpZk+42Aop9zqHh74OcggdbzexxMuEmDu7cxcPZp
eL/xobIaDFvCwvrJZRLpbOp7f765dVxbyFuEYIFmSz2DeID4jrTGyZjSsjSVCC9L
6e5b/MOV9884+sy+OMmRrMjgFIJQExN5Sb4n236fKhHdO1rhUfLc00xK3mtXTuG7
v0Zq7+3MA6zCgqLyaXTaJj57X6O0nv5UV7bnrZltjXXH5uxnvN1Rs49FbyKENVG9
diHGBHuEeSklQ481gZS79JahUglsshBmzNXNGA8X/BCnKI3h798XFbQ2dYR86+TX
9t68FossTNxCMQhus+I0X9b97S+DIuMBY5fZfxqD49W60nJJge3gVxPvUT6Yp/DF
Of0XfLXbzmSYnTHmQVJ2IdWiM0sAB6ONFhXSoFHwymsvec3hjyevqF08ivpT9XDv
nzYrV6PqF/DrO5foISZAg03Itl2P1bu9O6/sHpUxVHIz7nnBdJibQ+QFbHtrcPi5
SAfOKQJmUey6DQjOTk01AnoJ5yS9l0UiLsh2qnQZ0i3cGK+GQGHGT7wd/HQZBkmx
ha7b0qShx7LPBLWjwDh5Z5sDkttIQEWO++MBcUXjoHCM8srMLQnzcdopIlL9y5CJ
6AwLEc68WVFeWi4Y377wSeJm6d79ZnV/xWxmIyCLa/GMpYVpc1WDEAx7AV1PUAAW
eIOzhuE4Hec958Jj0EH9G+QLYwXiwUbk2b1cEoc+BQn88SiG/wh8cVXre4+y2pm1
OsWkEynLN/WBZvboGKK211hYlenV1yB6SMFeRl8P7gqNXatXj9NdAMUaxAoHN4id
pU1vZfHcx6QAeM9PFgSg3ojLP+/90lGo7IrPdQeMVM0Hf+iFbNnPfKd9i9FJoJAu
weUKc4+BXoubNUkBc8uA/UeFX/m9z55vsQ1vNweSzO4F/jEZEOYkz8jV2pINLaBv
T6N/RvVWLmzmDjSj3iqKvWx7PZvQApuihuZPyUAcbn05JgAwZMM+n7ptVy+E5qIi
cXyhzlltx6+cmFQp9o1TDDPUP2eFf+G3Tu5xoib+qN3lQ9UmVBi/ca222lF4EpsO
EklevP7o23JoOJBC4GdED2neTYUn2wu933R9ZMJt0/JwHF6iSAd50YyceXSscxWV
SyNc57wr37e6+L8DKskoWuHsl6r2lSfi9zaCVx+y/VCCJ6YBCi3681NEC76itQv2
hAoetMfTNvhwONkaLDd6nAbDipt0WQZNwQkGt1Mfpx2ocwdDmphKmGQAlJo3ra2W
5y74czJWYbPsOmSN2kPWkxatxfqQpOVqDNAq4izQz0n62Bk43RvozTe06ZS5dKWl
Wwx4EMwom8jmiriw4Qnca1u9hCdiO1fcR1odCvy3LPTeYQTI5J8H8PxWWHSTL7Dr
ekGxvG4zTznJm7K6uwnYKR9W+qKnds0nJuesHDe1y19RxPxYYq92Rkq+n3Sfd7/i
t4EBL2MgW7Ksui4Yo7AmYwHIUknjbfS11S0pyC3rHeDVbr38ZdAhgwAcbOSUZrrG
qSsAtBcmdg5EJTHeAIxVnXmmziUfyqpcHforEtLscgh4+NQP0meX4Ac4e/YQ/PHQ
Hd9Tteqo4++8Ax+/2uELNc60YdY5GWXLh6SqvcazXr+qjEvfz2+G2PLUWSM//kI9
/A0/DixmINu6gOMeK9voN5PgZLcB4IlVC2eAMNqPXIJcwYOimM7p34FrJWS01wLB
9ZdLf8FX1CvaVetYpuncSPGoAQx6/JoGMlhAoEmCAMzNTV5CPUFyzUSi3+ScyVjH
IHdvPSoPFhoR+g8heuZ2eLlI6FJL1yvlaZkU6sgAHmcET9u6Wl0vkul02GkWhi5x
bTDQYx5t26iiN8CE5poy3kwUfCqE2dyLE5f+/ANg3ncrFJseRo6DI8P6a0ZA5FNk
Cf3LTj/YV0uGSeFyxue2llFqtwo1PjEpAlBl0jpJRBqcZ8zKFYUIC9nMv6HpR9j7
5JquCGgIJXbW0DCx/PAzm7nqIigkSBfBlG1/e5lbTEdbr+gOIm1SsVNC6SD42gNh
9cj8Fe8rsZi594cx+Wj9hnEO6ngIuo+2nVt6Zo4AjHrvcG52o3qt3HBLIscUfVtG
m9fZ6pwLNLztqjuhdR7F1HJXG1GwLSH1QhAXE1kbV8LjeVxmZivEIo4A7VE4pSjy
RC+Kpb5r/9VmIDfd2mGwIAflZ1mPDnTBmXJnySt+mo9+45ybRCy32nnsLEM6w7V2
0kAfInsycflkS0MpzfmOT5CkIZbKX6BE9gPYmbZ202u5qa5lq6y3DpXLgfrl82/O
ZmLqoU83Qvh5V0hMDS0j1fVkSlr3++V1wVRhfRuLJ1wQ3SXQKvr+dZ6HWHyFFzEQ
BJ1Ji2j8uXhiDpIaabzNpOl9IKfFmPojRJE3zWrL1M21OEXVUuS8U7GWjOiGtN2e
l4O3HN5MFu6NtgSidQi+p4X4HicFI7q/nW5xV3/9j8z+e5hbjPO4DXR8AWESPvM8
RBlJH2u7NDmBl6FolOJVd3kgbXyTgGd/L1S1OksBmMh1VE7N8DZSGktym2InjJBR
McEUusgCVqu5rDqNUSmrK7kOiaAGYRpOJMtK5iu7z9YTQm9c8qi2diodyy6+ipPK
Ba+PAmfZ5C9uNmhGvTJDH8xC9IWegW8gLyDrBldQeziPPq+PvWpi76wPV4nj6NfI
Lmd2eOCrJfjeIr1S2DzqSCyfrKx8k6k4wcCED3s4oWe4dJh1G1bHSQ1b0i2fGyph
oRf9esOk0tIF7DsbezKjQGPs7hG8Mzt2Ziy7QCWuKcZIIHLsTmhAQyEyfQCjSagT
gojmaTNu8kufhL3ZKe2QBz5MeJravA5JjsMsE/DEmCr6UK9SkLueuF6qaFWmQYFk
kde4FtVuVFwX/uVff+0y//YKjxhdAuJ9hiaTrrCJr3dRYAZpYnwzPNxaorzOrYYZ
lpNbhOeRueomH4saZ+BJ/x3Y4cgF7njDMrKen4h2h15xsuV4K+T4M4Rs5YTuGu+I
wbBQYOuZenNgBVzghXds82NWii/16O0VsAfkssgKzB5nRsnTdizQryStiqTaQpVj
hCpsk7Il63SdXV/iXr/aYf5zbG1qyoX6aH2Kj8rtcfNFQFMPAKUI3VzZLcoxfycx
UD7M27cGFXNgEvSLoUs0lMYTqlC3SGzSCRaQb1R6ZzJXrGZPf6OmPqrALiz1htdH
UWEpUad3rC5ilSt65FjPXDIDQf3D06Zf6h8vX6Yu0Et8NZP75b6Rar1CXeqqayzw
DNeQR/bAIeFVbAGw5xAid5F65UZbCWGXVhZQFFiJSXfXgrl9PU55mDelJEKNaAJc
m9y+H1FwoxNdeNEX4rUCTruKponDgtsa2tKI2eQxrtIyhy9PuTwQ7eOrqdjGHBAV
BHZ7PA9t9iaFKU8tHuZ4ROwI1+XJ+FqYPGf13OYnusdH7FvzNRZZu4VbWtWe7Vgn
9YdB8ArshoTPyGEy/mcoAPtgwWiQL8v7rO6O5MyLe5zFvgYcKwcjMLe/L4QVhcv/
yAjbE0uIz6yno4iSsP2W4SrqGmj355JSzaGmO8SyBkOI3qU+xUhS+yJm9C0e0SX/
D1mfl3ofhIW8IbxO+PrhOkwGR1fbSvcpXmt4KEOoSKZLOm+8upoqztvXVhhJAJvo
OZX/xxR0AHSKLJL0+KDiaT8sK9cQuiNHU2OmjP0ZLZoeZVVNsFMkJZMXzlAxJFPL
90NSE6+HPy9MxUWqwe1ZB0IasR5O5LTnsJvGBQyRqLadRg+D/ginrFroGu0VmBmW
RNDZB9blICHxjyYAPM1jTRzrsDErSWnCK3pvRNrNK6TzJT2EL/0ixY9VsWTqf5YL
VgWAyW6qKnk2PjLD5NAtfka9tkYyzl10oTnL0Kke/eyVvUZZX0BGJ0LKVw16Uozq
MNvF0Xd18rfjT7/RbjKaS8bBb40GfZ1wi/Kgtu1XshNoBGJh85xzm82vigbvE9uL
h5Q49vuT1hI79TNIt8I/s0Eh26bEt+6oUGCGS0wnkQ5zOr+UaHBEmzNzMB8WYVEx
4itpp2lFF6y+GugNe3OVjnEMi7FW0qkZH4Gx8ahqctmQtgDujl+q23J0nY/FQ9IS
b51zfykOUDrpwmnBZbLwLyu2s07KWdCWg9dTq+OvAhqNK4Dvc9DMtNV9LJ8zDVEp
icaItvG0/XEhPEA5100gziHftWjBMHdi8+8Ls+5dFFsgS/20PN4jO1dxNIMZipkB
UKk2l//C71Px7TzlK5q4odAQ+PVpXx91Igxk5zQZ85gq09psOdjip8Ycbvv1bTw8
ZUOXipXzXL/OJ8CTRgJPT00QLTzXq2hzImntksyPFSq+6XfNyIRkPSxGmknPrlqx
RUC2cLthb+tsIiTVXqrfu9wtixqCFO07a716G0N7pqSTJhOPoGHRjkvuma8G3xun
5U8l9X2FF9ZTAebjJASrHHeCdQ8VPMXuT/wGITjynZDtW7RawfIsdqKZITkdCwp5
vnqivuKiUQ4uajVBRWY8pE8zNB2QYoRyy/blT8dMVV3nQdeX7qJTUHl0XexpXdRn
xyl9wSDOtIeejWPtJnB7bvfbCxTK+DyobgI+XyfWvynLNJqf51vujz0ZBUPPzPz2
MyozLfMmXpbwYvnZfbhv48nUEXm1DV39wVT7xXDx1x+6e166w+mFtHHIzeBCaPVS
pBmuOsLXAq8FjfyVxpNlLj+MfSRddStrwc4q3ycUN46q6ZMbyqP9G+rTE3Wf/vhi
LSIZ2mahJKd7zV1C+nLJsBLbA8+EsQ0nBCGsBvV3xkYzdUypfAoQrpveYgkwUdux
ewb4WS3P3+Q5M/6D/nPk9tEq1HhCGSvJ4vp0z9NXOwDO46hB//Mqh7YcNdf0zw9G
YsLaFaMeesRgPBaxkGie2J8z2+jUKjepB+WwuJ588rOHQib2miVmMHvo6jec/Je4
gAbyL1CE7nReqP54pM+ajeXPtCjIHKXuSoE9mhi9cbDOqTtoLC2/izpxIk6XtxhZ
VLXdYVEm+hITOP4sqDgYuBYUTKbB6h2oX1HHOMM5U+TA4dKI6/uR4LBj1jOdk0hB
TW9ZNIMlnUuutaRMXoEuLUOs8Ps4WiF8PC7SAss1AiIBMNSt0WiRA+heH2DkCXdO
lzpzzIS2uuduAgSKLqmSzN5wfXWahorGCLZ+JS+q66BluQ7aco1hZfmBkLiqNd0w
dXn4PC2meVnli66VOKJ/TrUme4W/le3SxbuA2By2uuQ7yiJRo+CJIoIBK/RiNpDT
2UcChK5jlm15GAQL+yeMVpPE7NyRjRCt+727M/HeEhS/AerQFQ1NSwM6gV0MlzPc
L/GreOGO1Qx5v4MImzLXoKKO98mIA/rOW5hCXk9aC+fiYFRSfj9rQiHreNTFJeiB
czqRp7P0HsKBtXLVlJuKRc2QyGWtTU4VSq55XqMYjnKgCV5ju1/ST44BhbR2ihyi
bZOm75+0VYADke7D7Rn9GDlpyKdtGiN1uy1wHH7poe0KABq6H6JkuwURrhlClX3g
Zqo9LW7Nx6RZyEXDLb/mSxH8+IQ8nX3pNRvDz3krWp3q73rUBgFzMj9I2e0x/tbp
c3qc+ALHYlPeD5YlOzNA4sZGH3FsI73vI9/O0KpvzOqm9OjxiA6N592FIHFkthX7
o0weJRAGruF2efnyYdIyfEYYhRxDbnTR+HV1jJRHavL4qjtS4nWYPslPEG1e7EUz
KY19tVmYvlZzdcZfuCdZyjNqZLkb2uJtfQhjp+qwj6YY616rpDQZM0z+xek2jtBt
fSs3gPjopXlU/AF+bYGL/W99zLGYqEnfqRbMd5HbuXxd5oyLm1vg7lf9JGQiWmTg
IRsxi9L6x8gTCFB1+QQNeSAfllc4r09CCQNigyOMUeXF/9ji3LGYzAF0lplaqqmS
LZLp5eIn90TWutsgYzNNzSvUwgtt0j2Yy81KA5GLkyfaZJzxHnCvvRduOwIzepE9
6FHfBEz8UBZfoZQaytRFgpZgpUX8noQIq2fnWFtvBSGpsw412ItNKfWDpxWdDRY2
dy/F/XDym1bo2d7BB5r/aQyKkQ7wTS3r0tEpI8c6B5CrtDHdLTTtaiL74UvoHMWU
u4utTTliGeSds8xyasL/xy8gcNE8DUGmNfGIDdlCYI3QnzCCotsgWmsnEQuGkav/
pjc6UKf6WoKdvSRAxeRbnKoWEuwFGMyVvpXPnMoMVKf99nT0PPgrG0/zA/KsOgmQ
0UtuNCtVhmkFRAYDceUuH1Ks4y2SPd0nFcjtI2dlS9I62g02femC0305mRvoYAwR
DvcF33jBE6/gYGySBVa1+/8d0NXq/nDOzRP235/7CYt/ZHEa99byDQskYUyO1UzS
uQxBpnMA94dGdnKSHHw9mILsRMPUvkjqToYvw2sG2hd19q1iWqtKHPQ/L/i7Ki4a
5VZTELf8SYBKthSG0aL5M+oxPGi4YEt9MC7MF/yMqoYB2Ub7lpR1L9Q2+3qgFJsN
SoQRItN9niSMQWi5V3Tat8x6jpuDiw1hbuNuVQo8tkE6I9GDObjDqk4ldQXVkuox
hmL3nKy/nKZxgEX+yhTN1a+LkxzTSL66rybMzQHnTZcoYmM23/+QbbgjmWXBP+q8
8PXcyElsyBHd/Tnza9iBucLCvUIYcKuy0zmakAbC5eauiEpzdyXdohZ8OD53W2xO
ZVURLXof23yppyualu0S00t6DXRo/CFHV6UTDNasydlBt/wop2bo2zvPAv10ikhx
hX2TwgKLQ15MGf1j0g/HFgAjNpl78SbwjO1NKMNk9o4/KRDTGCaykvGo3x05job6
IxB4pfagvsupNOtFbW8ypIrvFmflZ9Wc3sDQAkxKEX5IyCsIpASzPOJN4/WeiQBo
y88yd6jeG0pc4yWp938koe5bX5Yp5Ir7ZkD4/vyYkwksBQCimo4itiFRjLhlu23z
SQV4KAl+Zo95ync+d/zIhtsMUJBe5mwps72jKk7An5H3rOyUcA2CqdT5MFDrWX8Z
kl1KA0qMosfqtRp4yY6pUjckThfXD7AKk0JFXa+BdzTLceVLxCNqRTd2s6uvG40u
piC7w6jc/LkABiRYKv7I8/CZsLWJXNe0ASxqVmCuuU2oRb3jAgA/ICSyroXg344C
+XTv9JftCamXFl5Daar2RaV/NVH211QKYVNexs72ub9TGpIQCdrGCY0dqK+GY2NY
ShqpEs99KaPf6wk+oxtUEglewamkuty6UQUCzY8eRMdsIyrvg/IdKyz2NZCH3SZ1
pdRtnbR8V2Zwe/wgr0ZxQoJc7tSQHYdKRnKAkhIZu45Cwqf5lLTqvY+20zO9FhJl
x0LnIABPHYwAqI1jg7eN0D0hQJQBo+cL1Q3nmwQ1vjZ21WvgxT0iipWNfOgO+vCh
lY28PWGAKwa0MQehD7CLQfB1KAal2SoonNeJ5l2mYCfHtKmgIzvxpiEzj6gECQF/
seMU1D7StfPdJ4VA3Dyl+buKUhXvJ8rCd4nDYQnRBI/fexNcZ3J0E15a703LLf5x
pjkZ4BC7kZoag5QVI080oOiAGSwSkKTna8YNRfRmRC8i5Dps9hZY4dMOXKIBNa8d
LN7dqkAzr8iBViXfsfgj3dEaRqG2tpVBe50rjpEjtgL5OxnVi9/JuY0Nm853dopL
3VaGV5QocPbHNs4PEN6c2Q0e+WKk5sRlZ2Ng5VFdqqcbLWVtzrrD0wROtSaEtQu8
9VFKXgiVdS3HVAvUt30Ung8KM08Gr0bA7sn5AizPafc96fpNdJHT2guG0GsJepfw
rHrRo2yV88zIEsZRa5X1+Iixtl+QYgQQ5vRTcQsiH2xnIQfDcOkh+0ri6HlNzCFt
geqAydN6xPUBoppyOgn62lpp0Xy3uO96TP413l+mvA/siJoAeT8qUBlYxuXiJ7HJ
JTolfEAVjKL4J9vHvtadfCvjyMeR2UctW9HC2gIuc6kRFkNpwmDTxbRHoOu8v+5I
P0Jh4AzJX1/LzBWm0uUIwW0S8gEBvw2Pev436Thl+PJanvKEZ3fIJqW0q6BIiz2g
Rw9CCw52IETrAZP0s5ykf5YPvBcxGtNYo1XV5pgWhjVfguuJYGjTO8fmc0lW6s60
ecg38LJ+VTcs2vXnOnOt9zqnHhePeA+k7VgwWWXdNr/pXc6s/GfPq3izQDIy4HBm
jip9AqGS3VbwFw/R9P51jRcTgVDHbxBQ4w1bUdqnQXwdb3ggS4pXiZgvzO4yyH6O
ddZB0H4EwpQBJYsu7ZHbdXQes9EL/XgGlhhf2Qae/Gj0e2Rp60xPlI9Ie5b3j96+
C6sSZBEHLtcrD/y/uOS+XJZDfXOvl5wfr0xZsdyy3SIqm2ryB7gfG7K57a+4Mnpj
sXKSjEVDYNs6eM4xyukqecES4PQzSP11P3TiewmQUqO3DZaj6cQZvV5ImtfA9Dzu
7+dsn4HP3HNtLiVjpPdgra0qsP/tF5vdt5YjfUw8UlDvZemNAKpO+p6F0FecSPti
amoZam0/dYbMHrGiS3EEIjnA1dmYYXQ/MZXwh4zmWgl5uAiIi2q7Zz/7acc8MGlZ
prxYZyGAKKtwACduxbWGEvJ3BXVj2OsThK2J8uRlTlAIt7x0RYmMIaT9vgvEc+w7
wWnJwLUN++4EQJLhjkEBlsZTT+uabYMiFiWeUIPtxH8kjPfQBUMW5BOyl171iy2K
NuADvOysXHdaBfo/4rBTsTE7L+bdWuhTeyIkyUgXKxgM/ilakOPc1HxpMlRFm/Rn
YXKsxeWcVeJ1PDe0Lss2JQqzbibmM5tsHTkKixcE/RM6/vGbWj6o+fTDjiHW2oWt
CPe3enx0fX6rw8YdPCz3DFrLEk3FxlgDsQ3wXTAOOpjfhmiIcTZorRXdDzyF3bc+
a3hWp21A01Z/+nFHH0EXmP+XFRhdTcUdP7Cvq0T2mCo172TAM+5DdDeyIUasb5r7
cCtb0Er5po2kQkEPIlOZopDzKbZnxf3kYNmjxoSYGZ06d2wSiN209PXlYKTj4St3
UwDWULGKn6qRdbnFymUXi/+hnPVyt8O8aOhzaTZlbCUl4iBuDCAdZ/xpfwudAz34
IE0gX6GsACWCztLqm7Dg5zYIAnwtws+WeRsRX332vAitbZwU9HH5PuX41Tk7yIjG
ADodYAPQFK7ItUljCaK+6HfX3aFVfvGTFV93dvmvllN+f4TWHmXht8lHMKOecLlC
k9fFRFfi/Uy1T66LyxUbCmk0HGW8HEZyVrUk0zkRyMV9AsVaWwDo5fKPwSQHmBlr
6paPgXluI647OYxSelHzYvtqueWrj5+udp3t+c4BXIXrbYf64+IW+cG/uc1UyjbG
YBHSBfj8lECNC2nSt4Jx8RQ/QSDoUJDrDK7UXgjvuMhpugBarXipRJcdxW7LQXFc
8M88vVhyTbnmmxZ5B/x7DyujW4Nk7WNFLq+whlP8G6HlcEPzh0sYoZMIxUw0Zr/Q
YkDv7n6HpFQC96XAjlPRVZ7dgnA51To/uI0Y2aRoiDYvx/xmiKGF24ml/ncKG3YD
sibMwFfYXThxm28jYhTYbAXUJVsl7Us86m/y/EE12FV4sAoLQBjFT5zcw/Sxf3GT
1xv4yY+lxfSdGQmLEEPS53wx6fv6rzZ+yFkfaw+aNqDUf0SuOW7by4/H4ZNm2RmM
wCbvdWz78xUtl8kdVxQfNFmEb2UBCKwAuPcDidzoTVOW/4/f13lS+S+9sapYeSte
PFt5On40Uuzb+48LtQAiv9SYSf1WS29gM78x8tJ1aqh+4ZvfdjKcGgKXw5e32Mul
ORSfvP0wFM+86nYitC7Y3WjxzAuZhyg9MLcsiLaLT1LSlJPTAMZvfWLJe/HO5itq
zATSF5UhxK14jbs2DzEI8wpdbA2SLeVGFithua9MXeiuQhWXGGpTLsmMT1svenoK
SvJ3rKAYLzaxLzJqClgQKOcGSUKM+kGSg3TTYzLL/H6nKrmhUZ9vo2PDr+rL+Imh
vHthym49xQZ5jYGtWMQoDeFdIuhQGAVtL/U843mw++JTmyYI/loi8Z+aoJe5oc21
KLizaDbc+Ux3F1p717JkQ6wcc4b2R8a/AzwZcve5HGowsOG0DW+B3hL3FB+uA6yA
p4qoMLW7BotRECUr4EsGdhB8k1RSITon+qgt5ohXdIf8NoFbx1YjoRZBfHnqbGwa
DpSdqW5L1TNWHaIrkJ4oier0tbIuODkiSUlRLCwuIne6I26qLmREoyYe2Lt/T2iE
K7n4FcPOLegwOoG+RKRRQIlXO3y7NZsZpfIQkvxUneFkCEm7K0C+cKu1EIvMPZLc
eqerX1snCLXsu+byYojeAknPGZO8jL6RqLXfNngiag7/QXOydJq8UU86P4EmoRvo
GG5Oq9RN5XrwDWDfgdU9q2REfEAAYv1igJ93OWIr3soA5ZNjn5vTta4/LfOl/WQu
uE8ClvulHJrEEWd5d1H3M57B6Bzys33Pn1iBiaexjLK9qjzrRdfNCOtVDn3/L3kR
krli3qPsFiVSPh4ivhJoSqO0CgixOeny8dSa0N5xHH5JKvtJIcBR6RyS/A9ECCzZ
ROBMoZCXPfFyWdX8ves0mp1cCleoVsgLp0YCI56umD2fXWdWGuu+XEiKHTIT6rDQ
s9uQPjBaqWc2VzLtb6ECjqLQ+k+ZCeY9dQRMyghLyG4iSOtfawP0y0/R+Am+G7e8
eCCL6NcPB9Gbf4xqI0jPNdoIDNS0G0unlREWNyMgryAfBnt3Q23lmhqS8A4GC2vJ
oKWSShiyOftA9QKNDWUHAsopfEmgZj9g13yy0fpfud7KTTJ2ueeb5nUdbdb5VgVX
95aTusr2ojJafPWw0BytoKZ1uVJexSDn2OIRr537+CS+Eudpm4WbhFTW4wEZymo4
r8diurKIQYnHck3rFlo0fGuYXoSSp3Uz+5Usq7Qv2oBc5EU+XGaUthT8fFzwYbHa
TOYum6a9HvGcsvzYVWbfAVq3wkbmL5hPVRwHksrXVDip99UWqzuSTbDpDK3cTH48
ux108LP/8IPFjTRUS6IkvRy4kgqJ1bPy+gXODgL04KqWaqQE47O/FAhFlQDmW5Mc
t8wCLLAd4VhGNtNBFahB18EITQBSc+sAYvgC3Js3cvjM9j3yXVZf1rmPTWwtGDpu
EmUVAjrZVlROxjofSTyri+LNyYfCssU9mMJ8Ej32cJxj4bRJbKKdrMPjRFCMzYR3
pNXcJZbAauBGiGK9JY47Mh1cE0RM6BXEm2bqxYwIEDz80Z4cJNZ3DtCmgfPJNyr1
7TJ28eWxS6yKgCjDZ8R0nwLr09Sw+TgkWYXrd7QDt4smEMMxeV01g3KoZg5P7daf
jsel3oAp+ivDSwx0dTdajt4LteEuLTwStA459TalKLM1ZuoMPeOZtbgK5sZxhpOT
eWkQkHYGVS3ypgI+x7ErxMdtSi+1YJcokZbgvTHls58Bcdlb+FG3LMqlE2cjeXIf
2eWDaMnw+KlbnOEH1d4LikJpoovXUmSoUA7c5d0PrL4K/x+vPwhX0BRryteuhmAo
DvY+Pb2ayG1OUnifESD5sqVlJSYsIjLqgebtcJwKyTxUgmg92s6kEpWiSBm3SHY5
QDxaofrz/3+GahIeYIUneK1FmLA/UpKQH38t/pqEbKPsAGMOQWl8D00Q0OMTuFlb
eRReRnBn/OQzlgsFyUsSKxqNBwIchnAluCP6aupUoS/9VA5pDe5M/KgKqJ7kSZpI
AT23i+2hVFS3Nv9/4MabC9ky65rijtpWa6PyHWAgiO/LUJQyjUvw1P0bdN+FJMtH
4q9D+Wp8B91ilZoYYsdfE9Pouc6ALaBA4JVZBQ/xGScJ57z4Di8WIYUX42aY6PPV
5bj/qaebnrOlw506cc+vPTp06FJl613Enm1b/npdfaXoa3j6c+IWuqrL42fHXHb5
rzjtfAKVd51ZuYDHIM6UxJu4vTfbFuezcvsiVzT9k7TaSMMe5lBx++HzSYLBedLs
Mbd0CUhO/1PHTUvMUAOUNY+Kp33lM48yPnY1hnwoKoYrKqcQGG6LyRq/zRW/eKtC
q1EtBulYU9fu6DiYyV/gA354WVxyJmw7/DyoVe8wHcyApmI2SFpARy9JjkW6IlOO
biEX1YbA2KbEXocwIcg8Npmi+FfcFNCXy749552j+PG+EOB4PPBvYTFqvIosN2ry
Ou7eMKhf9ojPrg6r4cJNocrnSyF6mpUCsbOyAP+6fAONXU0eFkb77oQ1mtEuvdgj
tc0+WHDMPhnLDsS5Vkdgh8dMlXYKeqD5T6QsHpE0PfqhFK27k2SDJ6GkIbXkW1fw
AI8yq5epRWrlfnZA6WUZUfx7Ptlzmzyoz7oTNp5FiPtaHTmb0Tln5XmGz9/rKI4N
APgBNOneWaYuvvY+OYp+YyUFVvKUgYCGt43vXQL6peSBmBSGA9NOhM1qTwION0Sm
VWBn5ePIEaa3+BGJOEj9EjQeoDR7AvLT/ewEDureNrKmMt7hZ6D4v0slTtl8s0ZX
lirGwKSTkuZ90icJoLKjcPVmSWRDPwS/pZYHxM8y9zGCdgE2bkjR5++QBtpQ1Oh8
b3eZyjkewBDO3sL62GCPyrXj+mzgiQZzObqhn48rKwqIEZb14UTpwhLlmlCRe8Sa
15ep92mvOkddOP3YeuW6nBdC89OnNEXjcAjqlQmlBFDJWdiHwslixaOHBMX2fQuZ
jRMsGTitbO0cHODGUrZSvou7Bv5PrCcHhPKXwYIWIJtwYdce8sqLpAB2UxBTMPzj
LQj3OX44Yuh6x9dqMb8XZO2/vdpvIfLPKobpreIv2leT8abEwX5K3+fdOAZTKUg3
boQGkuvuBpXmFeDBpB/INnHM+kBPFkubQLQDHPVROJtJC7UhxJDV6jxoN4D2aIJy
/sZ6WpfsPSVqZS+sdpyIj2ZlZ/Cvm5vd+j2lxyPoDrCmsJoPS92HPlSxGRAA/xTQ
Z9LzL7PFClzfnAAlwMg3sJkkkViPRo9pWVpsYIFo2fRmEjRbrpdZ/zZzR12CePtz
97aCIL6OiVvN/Y30kUr79qbZC8Z/HHnbijzoZewo1F29ykqv03+HOeDkNJSAaHXl
H4T+PAzoQq4yznfV6eoyTkZskIxPD8QbXy14IFlCLV/V+BJuy90wXi3PyH64pKYW
qIGNyPkBuqT4F/jj/jQqX+LzDyGfZE4uXh8vTBYcdXuSOs3OdIsBpHoSGargfxZQ
mhviov+FjbHpda3vHlZoaBIOCQNx74MN6g09sCvf/KgtHZe3aYXPzfnqIZuxIilx
NusV9+WdpSm6x8ZlHcQ3gDTHKjE1hgsQHouiJkNDP+xjLrvyy3CxV6yYLPMoltSy
LckzDy7TXtYvQ6nG9B+aguY2u38Y/ajXv5SZC7V5xI8yLlvaKonGwIfzQNilRKrc
LkaOFQDepFrBc35/fx6LuusUIEy5I3H7d7HZEjhdXEN5TsYdS5+ivRr0J504Vvne
EgSaaJNduzJSreHieb+Ebb4Qeh84tGm+/TgbzDOHvYPrS/aV0cV2qWqwMgT+OvjH
7ZZsgo8s7EJ/0XNxyVe0SQ1EJIPe28KBNEhQ4W1ZxRjDLkIyRv4TDFEAEhPHRiZn
utu3oDeiggcebF0ID/zd+eIhfv3jL/3sVoKroAUjBZUTZTsAWKkteMyLTwAJxkYo
l8AQ09UFQuNa1S6eejVW88HEBw4uKjDlDmUYx2qmJOW2NgHURpFh2C+hKvpsdAi+
hOuV9iprq1PEdMQGtYcYxNIRVq05Lsw5y6dQklFviO1d7mAMnCWEkIlRtqL9W5Q1
YHQwN682WdqQQI3G68q+g72zsRsHC5mWSr3wUR+mPa9zhA5gBfdemevCu9zkssVU
IU+9O2EimH1F+UfIKFOk5ZflK3KoDhur0Mi1z6K6aGlPaqV+cVFe5TcTxkqUka1L
WsIi++BgxfhtDaxkg/QlUTBboQrfmZb5dcWbDzzez6T7N7GuabZRCrHliRzs8kxV
x+srjcC6UbE7nTk9uE0xhAUj13J0ikPw6j96n3/2oNLnw9AWUiDcXtxkqNKltKTF
qvDF2ZS8fgIbkXxKp8binZStbKAhrB3SSXJyvOpTGPZO6doXKBraGrL/aHdACu5s
K5+0PeH++xchmkJD+eGUxSa10Ep50+PWPNGlnRs6pP88J65S3F9blEnfMUtbNRCk
GAZGwjx8gJBZzYkq/psKa2g0lYi9y1EYeY4fxnl9UbOEgG5zytTcDHIC3dwGqAz+
L1ZzgmhyCjErFIZRz+QlQ+c3uvjRL91wC2XZc6R4qjsNlTGquwXFjbQc8LCVlM4B
Si60m4CNp6Uualeq2z24Sfk9aJyK8po3uKEKQi3RWezYoUHV5VAEUJYxFAJk7m9I
B67SmLCJB115MTgJTltcQWTsO9CW4MgfXKWK/aJocgtbedJW+QnSR42cRtTO8NAF
8ROFbsiPz3OUQFAAW3XqxSR/hMyPYKmGnqKbjgZMSWTVs9ZSWmcN8jZkyqrsFO3G
fhNzf6/Y3B90lJql+H3c4r7fBkb0wJUDbe/jpwQAtboiTOsHJGdde6HwJ2zE9pta
Xz6oWd5plz5zL7NqxZSlybgdXrEDVyRiGtjO4Xb/cU1U6TwSxby6TZGEMxxkJGth
xU9WoznPUC0GX6F/fNfgEMbzvHMn1pTbRO65ZcZILvC/12Ob7MlghIoChpca+pv5
kRuVdBFguqJ3Y6V7wT3PUw/iSFd4Cx21uBHk0jCO85OGDHJWbQi0fJsEj5cal8Lc
2i2s8D5vcbFI/LFveRpz8/LEEA3OM8l+dd5ZO3HZrTTGvZRkeDRsPouHk/VGRuyM
jv+jhzdYeC3wnqtKn9MZvNi7pbnHK3og+OlvQPW+pxJBNtE/HHY1dot8NjMtSzKD
SFdlDnuStls0pMXk1af7Ql5bDjSBCC9WgOK/2eh6gEkl1T0rqscwTapviFw1ID9y
auy7/K5PzQYW2f8IbuthB4FwZAMirU3KQeqfG/hao9S/bVNVyu1sgT4d+4pX/sMc
lgOge226zvdn4NY7y6/9JVUfsM6dEyJQnwOmkcFmat7hvwx2UkcobAlfPhZQ/TW/
dFcdXhFiDphEL9rmYd+R1pBWXg8but5IJWvrY6PRU4UdaMXwm4+TXBGDBg9WjYNx
DN7nFmTpNffJjcMU+3SQlhgmS0kivBYv9Lp6ZKq2SafgA923Y8ohHHjGIR2iv3vN
wQQgMQegz/lIgOrL8PnMQEOsw91ZSe9WAwpRO/3BZ/xSYdWjxRS5xAZwekZK9EvL
5/fDO6kHmtUNzSQAgiJdVEOE5JUh9GujN/v1yHmBBD/qINr9TXwRfF9W2C1dc+EI
hvDBwHfKBaktsnVEuTEpQGOe8hwiNucAdCK87jnKvxoG5szHeJ5QHciZ38QgCvUq
klZSLJt/P8mXg639dsUrVgaStkfXy7u+BXImxzeDnWy4tMm7YVV7L2JOJ8zl2XlY
B3FTn7ifhjXlUIY0C7nq4jRnS/6QG9lF09GmQKc9gGOsVKRMXYQzrCz9uQB4ksPP
NPKXIzZikBHD05F+6uuGJnQq97KDG4WSw9t2MEXSTtOpKg+hxhDi90xXE0VBE99h
V2d425f8kWo0vf24ct5ngbtksJOosI+bnJSc2HbevbZW85+vvs5iTJSOQSzYx02a
vL0RaX7uJUuWwm/6PaaUZZlqdpw+uYScSBNEJfJklVCoiBRQ0hCtcAWMvHdzlU76
JlthqXLH9XsaVCAUq5Cw50BmMTtmIa7m6+wjetSygyuSMj7CtGg2m82jkInlk4n1
P4erh2PqBehJ1jUgWl1WEO2WwGqN0BaNtvm4Hg61VESTuFZGkeJnsHWH3tnLnrtZ
hecoIXVyaaCBBw40+hA/ia623qMwivKrAn6i5CBWt4Pp0y7EhZdz5nVS0qCNbbDu
F+0tkv715G2X28jv1bFu4cskaaEg3+6g7A55gDBkeQfOHlmL5lcTL2B8YYZLGoqy
7x1cjlfWSLHInqMTpDAUnUA8CyFiHOX9X03EpGK0hKFmN+sv3c4rdx7mSXe3qudh
RxwIdgPiVRM8PtOMjMBlPP4aAio2tK7yNACbFx4mJi9ODenktVpF51xlTGCmgWK9
ZIC7GA+m4UphhTkbv+OfC/EpUZEv546XWoVi2UYkLWgWNzUhgwcecHNx5KiXVWKi
88boubGTqSDvaHrg3JdVfGWY4tTXRBCQFSeoICYiAmzv5Z+kYgvkFct1DwMlnUif
XdwkqTTeJQKLosSE0ZybchqT7AtMFbT3QUF+Xcn9gwp5XX/AiYQsLzd5NLd5K2W8
uf82o05DbBRpg3f2PjowFq0U0LI7fr7Xr0nZ7UwWfPADVoUAamm15gKouEwReHqL
SZTmjgtp8pnZkA1FcPNAPxh6VW04G2t9zB8gmaZ9ziaASb/FQsMkSktNdYtKI7cW
vIgdROwxTgQGl+j+UgT3Rr+ds6KfxSyEnQ2iVNT4nyr72y7eu34JZ4gBSJRyrvk9
ihiJhf/4E6frM6cYz8FTyxYtP5TdUNzNDDRVGX9Bh3seTu1sgWqBerpVZ4TAWMth
RRN8+n6QAW/gqmwMk7J+FUpudVdfIs9pJfdFfV92N035GBB+A2THnIAKbPNSWMzz
cdWJnWB2W6MFoULwafPHKmEEsTw5fvN6BR8sn9p44olTGyNIxWeXERXif6o3VEEi
KXoLzDiaxMlGqj4RoGe+yg7C3Ai2J11a8QaXXftXrbbI8GXvZRkLm6InQUa1jVyc
bCaHkOObgxVmmJt81mof801lZvSJLJUbVRx5qyxX34Ta0IS2nVXguCeW4Z80nFyB
exwNQw+fcfvnfpaqmD3xmUFVlAK9rsQTNRgXN8KagCjTQPdVTAyz446+s42P01z2
70ixyG9Esz9AfMkn2QHBh4VKvc082COS+yv1SJoRBKi/v+d3gnT5s4kHZfM8N16f
VNtLmpsAmtaAkLiz/y7G1VREUuCvQN38TKbMvpJbiLAadWT+a2rvJntEqfKuqW4a
niSktfQ+dswkThH+u7HSzSln4uUvo7UXVkQn8w9gxdiz7jvSZwCuqfZzbBiLE4gY
tSttXV91RyCHJz2IQiuizbG0hK0PO7z2iFxvqceec0NmDFqccu4cINfR9rVcY4gS
5WzAbZB+HtwS5GwN1UG9A5+NlT+zhw1eIeh0dICIVjDYbH/6dyJHvokgHEXoTK23
4rh7DsILMKNgcBBCwkDjcsGNT2+siwvWrw4oqSGBGrMzjROCAyIrBO15KRiNjR5u
1tEQ19U2DWIEPP5HMyvQWBhzrjykolj8nAFxghI87w3mrf6wXapYK4QxqajaBDbZ
Ya2GkaN3PqbFt1a0uY+ZF7eGbAFKvtAeRgV8fvv0juwPfW6DqI0wLvUPDCMlDIPz
H32nIT132l6e9viqzxY//E0EPPcXiUbfpxo+ORz60Ym3hNGKh8nS2Z3sesuAOW1c
xqE97YF71rodj5mncioF8a5UfPrFoszaWwOAu4elm780SznDY3sGYRdd281/ydxa
dVvzoaVsIZJyuMReTdrLdHZjITMq9WczkHhNw1hRaJ2r0dUNAlKdU3fNoTVzWh3+
RZC+abx3lNZZPsiOEw/bb4GlTPPlZY4xAAr5fp3SIWt8QPEjVszeB7A59FOuaIX4
8Wu1TA1rioJL6dVOiai++GNZY1T2DmhVGJm23zAtDCFbgYk7pI5MmK5vbwWHGn1n
6M4nD7GOzL2mlC3oOB4bG126pZyp79yakQMu9bZ8vGEu8uqMGKi+VVmFqyNmqB/t
3lCKZxkIx4LE+ibEtXnR3VaEP/PPdIlzJxVDltuNmgktbeXBXnx8ojI+TyN9P7s0
RMUA/sqUmRJwmeg9DabMKsfKVCow3xEEJBDA6dYIMKI7jwBo02zO2RP/dJVsgaS3
vhgEO5JVpem1vWhtNhzB8F4Qs6AqXfAgj4RLt9su42LomPx3nNgpMMt4gi2/0A1s
JtjiKhHK50Dg4cGuIglN4B32/+6mhWWXkQ/tzFNeDePG0Y1Hv1fe3yX0ETZsRNnD
KhhBrxPlbqSoiEWbOUUnbKPd9i0Q7jVUZmsIyMQb9rYMbFRh13Ud9lA5XD14Bfke
pKGV+INORBiSYCb67/LwGL/Mpj11Zc6bc96zkvZITCR0y4HJwdy/MwN6v3rmWMa7
+67tmwWU6RlPQqXAPYYVZe0lQ/3fxlU+tLCSsZTH/NRll4/g5cQ+USHmXdWz/b/f
BC94uqLY121pLKHfALCL1O/onQqTkkvr8GFgE3DVUrYGAfgopdbEA320lEPX+0Im
spgD3OLolahMXTqaeyLWsmY5sUelLMmQOX6C7okR36OCu+5YMI+CI5OfaJ1Rk40r
MuQwPd34UCChhbeTqdNjcpgeGZIUeIsxj1pfzYagMSyJYw+AjNc7vl+MdQr0Q9Ey
7sgJQyryN5FpBAU7CtuBopUNgbJf4bgLHo6eypU80w4QHfvBoVgcrxM8k/isOp7D
V3MkWczfXoQr5MBVmPC0ReYilPH3wcXUa+0+LfSZay+kjvZRH3uLsjaNbaxkgyYp
Q4L6krHWFIIxT4mDfK3+NsKHfU10lks4OsUp3+q1prL5B8+/pIa0G8f2xJW8LWxQ
af6tXEsKxIM/Lm9c9MB1oynWegrYh0lMjf1jx59dwAGonga3fasz2s4mumV6ftPU
o8W32zgcEZbeXNwK8ZJhcKg8JhynJWK1mPr7AgRwaiFT+Wyu5xw/k1d1s/bYqzTe
fyKCxeqDo4rq8FzSSznmuxQ1DJ7otp9YqGGiRTlL+wyprrxeMgXQl00QQRCBjqVQ
WWrZhTqWpu1Qq28I9VA4goYf3y2qIBXX2AkK6jszUGbpsKLYmQfaCOo7V/EsZdwv
xu2kPSFiL6zMczJ3Soa6+/dtQo+LMr4T7XO0Ou9in6iPIq1OM2oocFKkaVh5tljq
T+DxBgRs6S1M5EW/nIBaouTc264vkGksV7V6wKPtVQdXx+BOG4uXmUaTkA6Wgvw2
jFv1nrtlVbijpbK7azY/bHxDw6nyv0vMuFl2rfH9o+Xz4gFvYMHsCx6+0VMKEf7Y
1BletL+BMwCZRcCVjkQ9+/tz7RprpIAOaoe5fp7SKwFbDbHBrIhi7P7cchBWhmni
DGVNVVVIovO6/ubjxr6GsBK2Il0HziDRY2q3zqTDn7NDhbU2NuvQT40TwMNor2qN
JdQ82GeCwe1kvucaGAU/VcoUpcW1eK8qFTi0YARxkgdPhdPEjxTFTFUYj9pu8Xxk
2BoXVutTxj/zkZN9Uccfkky4hmsaqQ2dkodvKy0kDTIRHVHejM9E5ck5tfDV/P7U
o1xievAFLD+W9Nkbu54gJfo0S+72Ew/4T3fXlDjEqC+rC+JjPpM0hCuyvEglp7OP
lUVRjIBwZztvdBwI3uk6zrPRSSGygqrMXBvOz2iZywNO2761slfmAfj3TUB2tn3A
8TBn+Ys4AVZlxdVO0c/NyvcvK3lvp//UkHvySAj6+Y8iGaw7zAplZWMfb/nkEQjw
+fpL3NUk3pWKKP2lzQPJw88VqAZ37zuLMgApuIQAUxY69EeZn+5s1lBES81voXdP
3PNXTN1Lq+X2y2HfGqy12yfGB9bekICbgLguQWGvzEt56mZBOeFro7gAyMGoi4hk
pPAcCwg1SVnDbIga6lZTtXyoMnelExohVfOpdswuhCRjjxhTI7Y+B86BlVvQaRXZ
XilWPKu2YBJ7JVyxq074AVEFxWhxTcvxzlq8r0fV7O4whngpVW+RsOWKCuwq5Gb/
7LsrhsfsIDeaSczLuimjOsJlq8lnWLSpXRrUqRvFRN7udHT/6mtalcCi59uRbS7O
pwu+8okK5pWknIQriIUwIeoH34/hoZrex9y+ngaU9WbYI1ZvIznSSzBKc+aNdN0k
C7R6h2SPAaih7Z828+QkUX8A5t/PsLzONWyj0F3ytkDWqtp3bHo+s0ILkAbsyFk6
96o+CkjtDoS2BC312S695RdQ2x52zs7iYzD4G5kZY+XhdEXnc0Gc+iglGjTQsGW+
qmtQI6mJBeJ1PC04N62POzS3HP89/Aw7UTx3M7HZrotTuXVb2EJOgvT/vJlJq4VF
VAtZuaw36Z8CF5R2OYF6k/zDkvojUI/PsdSZUZKhsAiYk+L0pVe8JAOn/Rdnp2R3
UQGtg+iCYQ39dqGXxIt9/m8OzaMLCngJGHXEfWNNzjfH/aXvr5Sv35ziFdPMPunZ
3wONkUkI4IoZBuvjk3Jla2b0QMIKRFTdIH5qVoZFPKtyYTl+AaRUvLaie0fT7wzU
42clEbpXYUL9uTvSBrZQmlys314wlt8xQYRfdz9SISIHigL3fUWmABK8aJrRwGXS
kQIqfeYB5jouPoz5v3hDIc7ievS4pffbKJDTT9t7a28yVnL+TtPJBas+/l7xjEGF
f/63j1zcA9oQbI9/DvNnM2YPj9v0SMCmTL/XmO//4IZvqiuWMZwQ2kGU76iNmLgo
WEcGmPKiG5b8YWU+IGq4TdTv4sNee2Ht+JdJyEJlTpanSSxYwOdUr4pBV50pefVV
frEJEzhQe13+P/P92zITDxQGgFJYX8ddI3lXqmHnbbLucBMNR976QLhSKM/8uts3
gQRMpX9/0vh+YTrz+bHK3wZRgnRp7oq4Loiom79feuH6i35WCcWIRmR++3m/1v/x
JmzYzlqfhx9xtZyWarraLydj0Tuv39aMtu2nERGrKvfuN4z2SgppTJxQwRDyX3gO
vC/Ay8MIInJTq88zbB/O3c9LKA3cQ+j7t7J6FsxbJ8bBK49mUaOd+wLHAWJMrbk8
cFDvko7W1drx740Bj7g1xq+eAg6A3xN0WeJcSpn6IT3o7Hr9/W4cboYEgwsqDScp
dCw82z9jCB8BGVz7BSqEuUG2e3rdW8nt2wxWpaR4Sr5DjStS+YGwf1HLJVFUjI7z
PcGGlKMndzILzLNrDdVd7ofZu0d8EECiWAKoCblfUOwZCr0ffKUV7+0inFPFPNMk
11F4+pvQ/6u4KEwkMLTtAPaOVaf+Pi/Olc125+HTeIqU12yD6/nQK5rr7TRiNpbl
dU90Q9Ho8LyKHjhNAWRIz2tZpG6hp1bZfvt9eAJoRYP80KyJLlxf3E5ZeIT7GZUk
uYbsWLqYRcmS12kjDrNlvoOwO0lIUmYn4GJQznWlbdVc4VtQdUIy/SNAZtb62lW/
q0sYt+PYS675WNlD220wnskyYsad9gXYLjaaYomsaDURHPrVzIzGUNlWb9XrK2J5
A+hQXQKYUDyVKHQiYGUcu0/8959MnF0cvr9djtdheVkxVULJf4D2NMsH5nfCsMqK
4Utl36QvOLz0u7KBwG+9ZFiVKK8m5PXYwgXl9SQzYU37R5hPy07APcgXVwk++yjq
8PTkG9Uywwo4p9o9UyYiSy9x3lA6rjsFGhK6M6bNCxpawWfrxH8f+g5dce/Lq8BE
IhojKQzVryrl2J+e9HVDgrCVsPJNO/hSoNGAsUUeOIvnNN5fsPRRc+Dw4v+2Nd27
9RNOB1QasbLiPainuFTnC+EXnxGWWqNznIMUQv1coaggJxkQ8LG4QksC3aMF7rKg
E1XkaZFdvEpXyh/d5wPAvtdQASxjoBeGJfsttKgTRiXNdEG+a0k1SqyWZrNpBaLG
JUdkJ7SHkBJTBtuA6TrgQEbjro+wcK3LHmbLTW0AAU+zBvM2hxlGkMdn9/FzTfcN
d4w5vNKB71pQVKpUQfAwz67nqS5bivhedy90dtrCQ9mrXi4E5iKPTNUxMeQo5SsH
WfDen58NpzcxGjxHrgwfnWDqV7Gwx/pt4GKoyk9V9Qyx32S29bfL3vMG7E8ZoRbZ
vlrrH2iUGjTTxAHwc9khGrnigK45el2uVhdl23SWdRuFdrdsRvJWuuho6B2ABoKM
Zq0awYfMQZDLrXqjSzCn7XcJHhedvaBBGUWe0WOWg8KoMtuAeFIin6Ni5PJ3A6cL
ElrPqFbSldhR/NSPJ8FpnpGML9FxdmWCPt2xzVnG7EpAoL7p5/E9efoCPHsKUgZ5
hYNK+Beu+f+aGkKRa5NUIt9R/A2xCuNd3eYY3bopvSTL2opzq2BfL1sDFWK/ZF0J
yNZerlEVAOKR9BiXQuhmTnS1HM7vQY8/Ys5lsD7EM3x1c79jS51ddIaTYnVZ6y0Z
8IaQySjITIiKqO5/IfvNeeuwRg+y+7mUq8xEF8M2dmnolREIx5hjdSsABQDPS6nu
3X98RUtKYSomgxSPdfc/1HAe2EbA42iG+LvW3+YY7dfCnYZ4XgHYdx2jq8WlFGDZ
BpqBitNizQfxmSmjsg95jBygGeAfmDW56CapuqnsAWjapLN9aZx4R3Z6iv61wRYY
RwFzQEOq5mnKHJTnhfkOkx2mgv2lXLFrKwzblTKkXgbw1uuT4pb1rx+MUumLGE4O
J7sDfNsGv/TE+wXz97vbpkL8UqoaWW4Ez6Cy7RaM/qPv3vs5UpxyXF0vesMmXtcS
8ELFI2axRJap6da9Yd8OjdPSNSPSm3QDH3UdspFII+iqYGZR7lqX8/kmIINuQgk2
d1P8Nh6ZfgdBSNEmESCaa9U+LdZQU1G9FtDqOu0+MPVZJWyc47tbWJ8Mdy8Le4SO
2XSFPZTGHbRZAjAmZtGbIYlFY5pqo4BN8cfGHBcGmdwUinikVS5c4LUx5EXNkCJy
6OUFen1R0EiAX5MNpPlYKLkaUDb0tpZNIPWQJN9BCt0r/sN7gHhlepbScrUzcNEl
/QUL1ldrzaRxaXV8QSVp/p22fLta09YLqmJEFplof7w8ZurixYguUFvsey0IyMBe
aF5ox9mWzqvkcRDxVpJ8A2u9WeZbmp5zFPh6SSs/A8Ie6J+hlgzdtMCeRmX0gsIG
IHPfOKHCwfenXj08iK/2Pz1eDqOmCUMtsITswbRU2nQaSb9b3UL1D45hmKgpNffv
/u4mIUGViJLuNgDufsvh4N1fr+uCEA+kNuYhz6SP86DPjIvSjDgCUDNHBqU411ib
OZGl8AicI+qSZMerVvHEfCh2KxeIScy0tNggPEbk90IJulY6CFBuQb7oG8ygn26Q
GdYrnHCFm32B3KrIiVU59idnVVC7MH7gThvMdwamlkaD8vkXndf87cARgSLGpg/Q
ZFHEmcRQI/ikkHDk6pZ8TwGw37NKxavWBK++I9zdSrO3TPpXmnWm18b08u7ovR4c
3OorORFaqXNSnchwX2Lf/SIszg80Mj/5J/CgbCy5Zg1a/KPVmdG36qJ534nexr6P
woJ18C7Ogv6tnmnZQGbp8qqCr3xMeQwtp61+9wIJw7cl971GkaJgAGJ2WozqM2uW
nfIPMIQxhagQT6NjV7DOBDDOjCJcd2PQmvEK/+K0PWrl8culPaJsQyiHH4galKeb
NROKDUDOvVxn2Nk/Je+/puOdtJcLN/3+zF/BlWuVPnJdsrkICyOYkiRi47GltKOj
sRSpXayiQahUXe/+HY/HiynhuNdc9oVeGXIvxvmI/G//Pqa/fMvVZzjXeST4AhxW
4FIxZDr51z1yOL6Cw4EYGfKwvvgL67MMp/Y8fN5MYAP2mzP2Z9pJOPAiF1TYHQdZ
WpOALTDxEK6lYTI+59ruqOTzkreimNH1NXfQUz2jsxHJo/Ot6yStCg5IBX0lIze1
jVvAjV5xe4BZJKyuy6M/x8g1baacORK6owNMBZ9waKq0/ypFeqfSHMKX36hXKkyf
3d4WorvOuH3F2V53a/TUTs5Z5Xjw+xTmML2GGmwxCSGpVyEuVBJfe9dDzvSb20K+
CYAwAd51ZQkZaAn1EM1io6XQ1Bq5C8K6rfxGmcEPd2MXBCZyoINIWpHihHtrammt
Hfq/XU1YffeV0jqBqxg53h23z71Rf8vB/56+t8YrftnKsP3JJB0p1PzNVZ9rs/Rf
sERQtNHOwMjb8Aafk2dBXCmuJcKsWv0V4+Q74MT6qKyfA0cP+k8N35INXvcyS6Ki
KvyJx8VuEtWBlZc49ou0CHAWnR7QaCTYQ98MTgW8bTk1/WU9Q8QkdPCMoR50vPR1
2Iv0dHDKSgfmECtIO4wDATMuKYx9TFAcQeuKMJMRjOk4O4sZzsY0+8/AIg/mxx+O
Kw6S8QDkUt0vCkSVvWNdPrv4o2zGx0h4ZkYS1VoO5DVcgbwLWEUM7oStPa+X7Scx
NrdNM8uH84UWOgY743aAzj/ePkHmXZM5k8qfkMMu/t3c3Fub3kKTS3qEN2Rl23Lr
C5naOXMqteAFLf2FJBiMuKoqjfPX1SKFaZ97WKlbb5eFq5oqrhoDS5FULxcsb0C3
+kxmPgxb4u6VIL2p1T12BNNAPQUN2Nin+PIxo5kvVbIU/JvFwlUpQUOVfTIY+NhF
7Lg+DlnHR0AYYoaCCZZSl0CVX+kACHJZS+YQbX26gbhQXs8Wd/1m+Qg0KQtx8huY
2BcXaFyHDqLPkWaU/aYMXc6DaRyNakysLDhwOEV/HPp/rT7eEElrEcOX9E9a8aTo
gITcGL9B+Y2zrkxqS8xH8WZAcZNImdkyQ9eu4fNki9w6exNtCvw9gv1lNr68Arga
9WXKuY65Rg7twn8OXMi6pVu4HZzpg/MGn9VGxGwUeR3syJjTCUtSC4G5ZSaJ1BWe
x/A984+bblIhOONwY6Sf8vFI4BdhdPbbQLGjJwdS8PQ/Jw/8E3+jh1dTAyDZnGpD
THmCeCaMCfUOeZqOzzfp2B/dup2swr3Fv9aEQMl0qrECY0oT2NQ/Al4CZihivckn
1+S/XS5qMbSTDIwYfC1E/LLgbVmDj0zlB2EM6LXv3voeb2mQjsIQKcDuk5UOImqB
U8fUqZk1xHDklG+DVFgJ0STOmo9mwqFA/1FiXFUBy8R8xkACYTHKwHh5dHlQ2CEH
tqVfLIu68Ppg2872SUNbML15ja4uE1LCaPWwlkQZLy6vIHSVZgdKi3pF9Q+CnhBq
HVbpRUsllHz6TEDIga2sT87xW0ArqTvEFtx7OPiXq5vbrVKoqLRN1Xbrlw5UMrdd
MJ2EzC3TExow3scYmo/UuCD8H5jls409KqBKKDD5AM10rYKtxIOaOvZepNI+fe5P
inIBdJcwi/Qp0v3JT7hoJEGlKqECmqaklJ+L86nIWxGNrAtSz7E5cryKn/Fth7Bq
E/HMUr+08GkuJAnAdQOVpZVRuFdspNXhT9sdp91Kjzlyatbv1cEMy9ELewcCr6z6
ivRlORugFtuYM+Lkmd3RDJ6SI1ssJn3sDfofHOFUSOBiUwfjjtOR56oOvoLsS59q
i8cEf2v3VFNOiQds3+rkfZTWBpAexLELvPsjjMb19/X6MV1nv1jAOzfCVYIXgEgY
uXYfWiS1/raWdf4TBOd03HZahl+d8/b4zCzmzLZcMeVHubJBrkTeFARcZrV4hght
Bye9XTyA3fM+FPIYz8AQ16oVbmZKcfwdyYwHoATPSPUh6QRGv9YywJ5EMorx6u7s
6iC3DAzkgY7VyRi8bu7kLT8UvTlnVvB1p/g1TkGWC5TMos1q1dgybM6+ZHoi9oEX
nCggL0VyAhhX2Xby0w+Nb7oOjY6r8UMtNDQd8dryf0oHWeMu5bLV0ciTQb4rSsHG
6KRXxsGWIIudqTxYtJlU01F+paIv9/dY1fvQc4NRVadjXAg9sleXDmBL6KUoPEd+
fycUucmmcMFPIt0WeEFLee/o3XZyoihegR9VhnLsTjIqSt2sqSzsYFbdz8BFk5qR
sQzDkZ68o6b4KcMFbyVEDw88nK8EyBDYaPC/+L6tuE/09LqNudk7971rnd0khJ5B
BVxC0cL6nacE8ECJZYCsyfHIA3/JBOFWb5kF4ppc0dU2O+d5LBhBVFkrGHnCZck8
1Ba6ELtMQNMyjReftMam+VOMbDCF6XiMiaS77tszr+n/HZURtSFk8wHsDYMiMlMj
9Xhgor+LTLSXkHADi2jaC6xdXyIA72Q31Yb6EYsee/zDrRCLIbP1kjGeq8HTEcPw
UfP+nFnvE55Oqe0xdmwgjF0UecL4rpPeLM6UHPEzDJsWmPPlWrDHx1bHeQstr4iy
vfF9t9Rp6O551IeyfH/M33BNFlFISkgzRXDC3mycD8K3ari8Anjh9I/wliniPbpG
qz6H8yweXl6rGhcJPpW644U8EMelHPiAf7ZTQVN2ztTMCVqswWhmJTlQP97gos/W
lNMvBfo6YrY+ZsDiEuc3RHvRjyw5rCe2bxEWVIZJZ4hU4FlD9wUqW51SSs0S/aRB
NcnSYMmNHQ98eKPuCG8grYh+yCt3vXQ+3Q+NRonVEPP5EFZTsyZoAkp8Ikqq5Kxq
fFS5sd+JzKhLBCxhUnf4c9hJ5CrSiHMmNU3eMoJ34R4F83NV6cJvM6WWY/Nck+Ch
NwhGy2u28S8+KbYe7QMjFJnuJe7snKdSArse9Kt7ZRnOgJbf2hEh/gNdfX6jHB68
UTPb50ggKLR2WSBctV9onPpoHiLlpK7uVX7e/6HrWdFYHmgcD9PJsiefTBmOvNQP
Jxs/xEoJznMFHhOItvZNAfX+fEag3oLU5I1M3AI7o2KNFAKxbsQbU3ECSRRyUyt3
GoLyTXtR6HeXWlV7zsducNIN/qd5WnadRvJAq5OORm35mpRgreAXdZwQ+bwe/ODe
oYZQ/D72gb5MQajkcXw/FlcazKePuw6K9ssHBRqJsR1xvp95sZzTRbKkgVuEniYi
8UJcXSHaaBBphE9VY6+qh9ckZSUUxVC1CKkU5tGbYV8B++6YDNNWzTdKmez0DHdJ
eaYU9gkTbUslF4PtFRD5UHPmr825HVeODWl4o4lgW7htq5iLb5Mr865RrZJgvcfs
5xBxdsQrTjxKElRxhODdo/6K61rgruaDBwDjqWt8QrO4JwTfTDLsK9MayI6x6uiP
vpkaL+sTxt+IO/AUycgNCFPVoMJaZM1IwRKu1o9xAKWWRDgI6qzJxSfDR8fhdkCK
+cIgpiNU1G0zBSSKZykjmNHP3+dGSuy5Ny9zdvJVPFMDYaaLs1aioUpOnUzE14/6
HRCSQZAG1Z/WrrdcQF1HJeT3FGYGH9S8+YFu1xMAc9PUjukBn2fsJjcEQFKOphOj
3sXWreoVdNw6EYe3rp7/A7rPd2SFGwRN6YJog4uYYDvicOVihVRvv8I2NvhK9sQY
aeE414tp/RP3AFMgKfHtt5VSENlBycu3WqAJ6Ap25cGZ5js1QA0l0aDA8N6MIJSQ
6Xch2NseQFh6FihvqC1Hyf/XfXrWa3KLHEwGZ1+f6M2T/JMoaHE7aQzWVCToZryt
VpCtONhiMxOD+grXwrRR4FO+cKlzGq+pMxAivK5hv36TnjCG3/jUX7PE1TxyF23k
LCXRUHj7QyV+YOSRPh1R3wCsxtrO5w0ey3sMhlkTluoQYwvCNebCxBj6Gl8/MjOA
vxwqF9ocAUWn5TgqS78UPr5YZKhDpH7snXTY7v9vNodLf3qVXD0gFEorDF6hX1eX
HgtKk3otielFAVJtaU9UqQkP/HTKdUKoLA76WnV/6DtZ/TFsaktOhigYIyjR+TY8
Tsqpy9f5jZ9EaTLe9D6tCKJIILb9LJbjQjd0tmH+21VaRynMwIJ+fB5M2iPEp4AN
FYUXmc87taJO0MSZTRzvBYVRHFhwrAX8FCdMF5+kLwVuLcx/JXwQv6SXQTTOxqV8
hoAOY16oDKOLwkSx5TSTSCYsanzD+meda/61C7PsX1mwqiCRX9IfjDxQvN/EcL2F
mQRJusMfEKKAIl+EYhnOIsiVjRX70TRD3Xggm1mp/+IhmXsO3l0Lkra7fdq1d7sJ
8Sbeha2TsQeYnL1uJLFS9a5ZAXiwdnwBTLVWFd7voTR7kxoO6Lhe3NhyRZPlKg7z
T0Dq5WErCXdwR/nskXLXWsThYJLxDOocyOO9j3WPS+bWejJWhQiL8uS9uwQiPJ0G
sa8Amb8/o/HPaZhwg5XwJ6Q7sbjHlzqSOX2ghc/0qm++aeFs20LEDPnqNwc95I4O
uAfYwRzoHDjkmu6BH9qpgq9lH06b4w7GmkDstVURwFQDmZxnA8vG4ip64JoRZNYQ
u7ltqaVdEqYhu6Px1JrpKj4uiU+I9+pnxQ9r5rIdfKQLIAxFZN6wTThgzr1hLlLs
fLh3Y2JFXh7CzXW1opGTh3hpEA4nteU5y26WX6NB90ULnA2228K5KhUqPQn7wxmz
Ihl7kJt4GpT9od+YEaWun00oR2Tx+Iro1swunnTLWP7qMjeQ1XJORV7gEWfQK5QC
Qe/3iGBFu68UigRxt4WTeYF3gxkdSwpf4ayk7ci77VXLTS2EQI6ILgTGnodQ5FXE
+SC3BqOQ8PBETtyFoOBxsYTAlZj3EiTS3IFMTcsDDgs8yDyBrziYbNVpnC78oLzX
vKF00xe9wT0RkB3FIjdhUkK6OQQKz3gTcpK/bQ2+l68QzASWk8jUAiUMx5sc+4Uj
+geSaZqs9GInpU7UIMXyJPELUayuXQe1ctR2jmA0Iaekl6eYhfb3rfNJXjxC5WPa
a5yqXiguHkvfLZCguWvTsC7AReO8/Meo6Ukbenab+t6N9ZSx/nQJK8tuAsnYIOad
MZiH9ZcVISLmlgbaPqeqxlH965Uubhw6ylM0+2G7J7Aqz1G4xq9/K4cihIOw2cf9
h3BzasuX71NOKrIzuzAnEg0DMGVLuQtkBPIL2jt/368FhMLiQENe1xlN6Kqz06wB
xCNt5g5fzJ97n+nA6ZdyQLJ25mDeoobQPzkxrpnoQW4tnU/3JEzmUOqUUjJ97gak
yUoLJPjoTgmtbBDdH3I8JbTbKndr98QRSo81MsdMbbHkQXdDJH2vzrkVQioU8DJI
6NKoUpGGwTizsdYCqY7DNgcN2OvwysEJo9tdyHdv7YDN5S+AllKS5+RoEKsMXSBe
hANN7g+MPdj1FUVO8ZwaH1KqpaayEyryWt/yxDoonJhJRFtW+lgjXMC96Q/4m0Uh
t1fo8KZQOrMqTSG3vWPuJ+CEdU+Uq2XIfGA9AHShGDCQNBRsHpDqkRnBtsyCY82b
GC5j5SNa5gpeLZbOvGRkyscz/ausQ2mgu42MZf/40FxewiUwhXVBOihQRT71RUkv
pq0eLtsty73t9uiNCs0FUB39CzXuSOv1n+PhnKXqaFVORwRrse5A4QJzebET25r0
ycrM/DXZjb7uXgXC+/GNgceUgdbNAZls4PAReelYk3h1yiOGPum5x/YPiTlljaNs
v7smGSarWU3Owlrh2EWNRx6WAaPdkZlvSPu8Pkt7GG6288F5Wrhog1GsvbiGdwGl
UvJepxJAkxXUSsSkmy10fW/1ZcZFkPAPXZNQy7IxL6e/h1dT0/5sVeNOdlV8/YcZ
6aRh2E2OmH/5FTotXHpDAjEVuwTtLM2CYrZBcJm15Nubq4M0Es6uGGFSnQqO7prU
6gQ5t8DQHeSRyIGQZMc4ztjhWIJsafA41yx728w8GpMRqM0FmUmm0Aq9DZtU6BxH
4axZ9g+tHg0+nigx6jtY6dgwq8HTjTUyE1nY/0scuRbIilrjtGUJeIAYslnn/vEU
28Nc4JY1j6kjS8qj4trjVFKasV2Agx7pKJJqssnGtduV3az5/VvjRSSOm0dtPphK
Gysq44qBnZ6gO8xJm+bg2AM2Lpqtfk6t7dBuYIKPhSERazlcdcuZECb5tt+Rrqp7
If/kw2Q6HVgCw6FVMBcihrwh6y1XeowhNgCY5FTCMKotNiw6u+AZ4zgLSbQMy5Sa
2odn2NL/r9dwTQ0V0OxUQ9nPZeDGVLHXoJYQdppJ3Ga1K2ZlEjw0piNrCQLwOmFr
92c6L/FWIR+hH5AKA1NsXkJVej/9m2qiLE0ONE7FCqR/5fXRXLaM1Iwon3wcatKx
HryjFYNEpXzzMkALG8MD1IbE/E+WN2qxhanxmA5sNmY8KjWuZC/LPOEO7YYAin4L
/tR3QBdgMRa/9jhOoLvbAB3CdIEBzkk6ihTzGS6jvqIqsgmtBX2pf2PyeXULlLH+
s7qthz7fxiFxWRb7fJljGf+4dtDmlmgNOhBxlVdPSnbPd0p5fyoRatk6UjDJdc46
xstR2guWp+iMNNXa7DebPT4vrXoN4Xh81wW7rHLNBeGo0354ezmb2g41biADa3rB
7DyUH2XronGRVuEJ88663FUM6DjU9SbuhFoPtjEiE+ZqZQQFvbUrdnEkD7fhjVQ4
wDQDrfOxnpSIQyNHKDvxC9HI1cFMa/T97JM4DWPeS7CNw2AEZETpIQta5cgMAQRP
vlROGSgFwb4H+32XeZm7RvJe7tk4Q9K3IgaSLgcawRiCO+dmYV8SYDxJY/9pbhan
q/kR71QjzsE82l7t5B0J6uE/I8QAiUaZn/OgF/e9nx0yepyFOMy5TjASLdTcLXJ9
7tOYSkjJ6FvTMWwAeHf1xCVz9tvEj3SogT6l+rbWyPgVU2+XROxxKDhd7yfnSIIP
aT3ZEcDdKQu/pLIks7yx2R6n4Lpzzg0nO7S9MCUAWwFdBYhpdypuIls+7VszI6Iu
CkGn3BRQsiMQumfSuDcS9JQDciwWeQMUB8cejTC5Xv5Pj/e3QmS33cznFR6MYnKE
PsVPZpndEiOuZMnZIsS2T7gVm/eCCNkjYLx6qHGzXtrHLHN17wWPnQSiIYakZg8r
LY+2BSr6NEdQ5GjP4BJlaSkV4fuaUNWT9D6TnVT3xrvqwDVni1Wj7R4zsHDw84EI
qyro2YqCrGf/wtCOGAOfBivKiiKrFfaBhOvlE2L4qEHRj42+VICrZlKoLmU+SjB0
si7aPpCpGi4fjZB682WTNZDwjsg7mQhQRq7LrwJ0BbcAWSHRP3Vg7ejOaTb0/sQL
Ge8tZkWZVVWgUjAjviyiKEldR6A7v6CzL8iqBK4Z1/DaehiLMB+i3u2gB34eVr7t
iYsVJp/CHnD7rk6vW+tCOkvQXf7oUBCqAyEr1b5g8K2u3VDq5e5F8iDFsgc72v9r
Guh/Y5ea/xVNslgcd7kJh88zcF2YCPBBip1oeIb3ihDwnTj5v17k26Zp7V7W0RZP
tbEvvah9BYaN03BxFNC2XCqB6C4v6KRNhT728b+pSF78+QhY7XtpstHlWeRGXUd2
8lF6mjdhroTkKfuK/BWhbxj+oqC2YlZFxT0+04Kq/zb1VdvPdhOaxkEP3ucE+PBm
FDFzaihDe7+iO4mXclcWqiNZVRplBwK6WdpcgmCfG9g0/zALlir2i+ENQzlWH7l2
6mlRUHqZWQFUF14xdoNlJP754EVu393HkK08LHVBEPoN4JxO2rliVQ65LksKThyA
/zxyjAGpEqBQleVvWFHEtfzaq+kkYFOp/KiMiuxhp8+xdUy2ayUZgdLhbFKti0/y
MtZH8gq+QejXnaVdrQ8nviqnCFX3Nl9nyDKrOrx5vGyKmLO/tRha/R7gpXZzQSSo
d7hHa2Upcj9e0+Tn0hRWVwCp/88Ibagg/8dIR1tbzdOm6YwcMOvssO2HZPy3oMZY
a/iRtwTLLMXu+13z+gM3HjAv9x4dVt61f9ynmay8wFn8bJI3O3tzzvmO2r679+wL
xGAwwJokYOJHV6j9zHM3rivb5+KqjAUI6wdj/6M7SO+YYnDcRp8F8I+BketrUwtO
yLos0TrcLGVvSv90mv9pAt0J/ZubMKoM9dkcG2eNFfZ0o2Oq11oCfnw42D8y0dRf
mrbwFzURUBUyfhMqkkqtBPZCi30LEq9YIFWUgfBCFTLqmIfHuJ387K/sx+TA2toQ
8OKTHBbrdO554OlqdbqGm3yqWlvwD3udR9FgVqK6Cjdu1JtEDS4zvhnyLq6Ln/OV
yfy057oEOk660oMzA55AYZ5+GUxT/CiLOO/IVNc6rLsZNO9vJ3qyQAPCi5UYHV9F
dY9lFZIyGrnnIjTMYCdGPi3ehQq44NxKZGVOV2/GXRHVnpuMULKitszgYJet+2Ip
pemJ8Qd2YL7GvLwytHCuekej9A/PYJ6pF1w4MtsiSZN2FuQYImKP11I94k3Ob21h
A2U8L9CukLmm9FEQLdkdrholvDdflaYPRPkkyWtw86mdpiDIq5TCykx3TDtA0N8T
bMS66U3a9AZRhUdKIhPhoO6YFeNks4Mno34tE7E1eqaSatQiRVtmJ6uMHqsqMNJl
IWAc7RdzPfdDaso4LiV4mZKh7/2ISpmNfF36uaHqprpV56mm2U0aTcjmRR0no4s1
BXzX7iQPPuhehwUirGh2X4GmW//OeJsY9pZ1WCZCXtLFhc3oyhHsY2guD+wVl6Jh
Y8cvFb/AQeN2zKVTc6mZuEMPbIJRGqt1bILzKSmQEWTCf5cT0lz88vTw2inFtcWD
7iOrawU69yAext1J5ZWGBzI1lYv+fyHMQTcADHeYhiQXWziD9/e9hkF4ifBCPsYb
AncNikHBgcOcArEG5UISbiy+uA3R9xJ+L0lXIMe7eTy5LWbif8R9QFkqW2DvalK6
X+LMr8kGQe0XGd454VPCjbcavsr1EA8p45/CK8jefZVRwepzOd36KAHyPQOoWdrb
fs33E88vWswoZUd490OhrNtI6fsHNop3QpdE81WM9ppfgLASfJdlfA7uq1Sf26z3
EnRr3PeyKRthQAq6LbCrFzzPhf1eTgP282zM7J/UmNor6TlhGpEt49j5UD1seM16
ou0A/UhqQwRIiA5DByLWZ57qgq6R2XfugdY+Pree+hm1mKxmpGwVHZ6weHo9ERTZ
viY/oztGp3AMmACeRrCnAylMRNLyPlyBqAC4N9nDctEPXjtQez+Ljr6ENaJvn4zO
3oJacQWK43qjiuuPBdAmsd2VjZSuaDz7CTEKESWvYpNBRYz+Imw1ndAD0BuPmx2U
qTo7NKCJW7o+ndF++pSOa2HXuCWqsFWqxXjgJH1Hmv4rlQ2NP1sh2kRe5Y/f3Jq1
Yb2OXDhbvw5cOPlyq4ssw5TeooOabKB84N0z2ggj5YPGOSO6nwylq5rJdv2W9E24
ZOui3BEUSkR2DPECIYom+XlRRX0HHm7Yqdk8pFsBcVNP+jgQohWxOhTImSkzxMYp
tEV9CfK2BJIdH9dZIhegXba5Iu6E1bFaGtFeflMJJaPAkyXk+77mCeEJN0Gsr+y2
joPhHfJXcfw9mG3eDhofgR04ob4y26Nryvj33lGpu1LWEPqvgyp9eqRhUR0vp/m8
dEOlk8hReNeIZY1/ahYEKLKc/3mYs32yBzG+dJeX3LV7+fK93IWRHGTUL5o9e20n
gQ+0oacjwoXHB2YDSaXJmMuMMFXhfxqIfZOjGYBXw7qn7XZPlvVDwJA7MiNuJv/p
ly4eNL9yeLQ7oYeP6wP2zhTuyV2oQhZOcIMwQf4iPpsDgWwcEbwRbGIEXRQH1DMq
EAFvvl6OQJm3lTSOtOSMhjmGdOZ+ku4e/0WCblCDypwGyopn3B1VXR6KAaRJTFtR
PDDj6ANIK8WIBoueUsFcTc2rcqhDgKRLvVBsN5zbOOU5bQBGHIB8cfJwHU68dCT0
Gomt1UuWKn6dpkhjAdzkKl5+rcuTGqwsRT/ErgncFOG7zw/DQjAA4BftcwDIyBup
sSvRJj9f8Ov5mqs5Gjzl2t0vqdCi8FW3BqgOq7NWt93Rc7a1EonlXRMMrZLF0XCM
AQXGJfW+w4JzZ8rhkcI+iEmrt5GPuWjD3lVjZyXBBOkDHAvjCOvfXjptZUf5P8ar
/pbK4FPyhr/axJeiC1JFuDM7S+lAAFzGu06GsO/Wq2n+T/zFn8P0X6yjPQ6bJ/r8
hsb3laa2mbJ4izUoUhPFqlSXSvqNrXm3HWJUAPkQFbB76/pRW9ZK36gJwqb2fyeL
Too+lVYrXjo2SVCFQ84UWzDDwcqBKjsRM6DNVteHXlqA36jEJM658Fxm4ZdDC9T4
/v1ya8AdruedSXla6mzocsVAHgzA/+OU7/nvLwM4cLinQevVFwnRgQaVHzYfbNyi
R9R5Syen8c6ZwugOmiqNuP3L+tx21Rmiv1awpie254ZCDiYeaAxQxxxuq7A/W9+6
3yPrGkdBSS80OMjr4xn2kItBDqXVTsg7d5s4DNb9GtvP+M2sxmtHCv48/n8mBtgF
gSvvL1h5ZHPlj0bfPZf/q2WCSdd78RlApFFOHuWw4LD/bMyOsoI2kaL40ya7NDSK
eFKuBNaXUJkSWOdoizq4u29d6aWGGr7Vzil7kP/nSkNsamOpqmcxpBJnV7I9lQrR
vHYhSc1SNgesb5MgaV1a0y/Y+PuTmjDFmelOlvQeHsyn/hCN0paxzAA4qiCFBu94
JPqp/UI19Dy4kghSpkEnpbV8tzLKB3Eya4zO4HeJKQDGqPKxfy8tQdPwxZstt9na
IEBX7OynK6BO0/nrBI2DHUyGk0S8TAtHWjOyYo83KN2Wo2el3ALYWuIewx3AsjkK
lNosyQbffLuDpKSD/s2qYiLWizWjLLvo1uzcA9sGWPhNqZh7c4b9iTjvRddjEGkd
9NKpCPXMHAAt4/boOGABEpw+9cGYLeSu1qPvIr88qhOnS6nq4CBJJf5Im0X6mZ38
7CsCzZBVLCfTApbiTWXT9JPxW6csYFFkSxxFw9C5+iQ4tlT8RYrWTNvGPtjIq23+
ylb2M/9O0/kKHkTbvYBvortFyMpUFVL2azneZpSmmFlSQBnG1CiSxP3zD43ZsIub
mGLxdsOv/AW4VU1usc/v8b1izuQH6Ed4oGVckNKCR/T7XiSHOLkwsoq+PwXlhwmz
E2OLQGQZq5MaTEdVY+JXC2eukADYAz9+knFEUXx0pVmX5DwoGYaJayD29M2AgEv6
P1W4dxicFcfIOgcjTow2aGa/uPvs0cgGOSWZvIGyrHjSjHHe0ylHEj9vlL9QusUu
568iWlF8LtS3ltxWK1Dw4yelL4KdldW8yhiH+I9ky1NzZYu/ws6VAUS3n0185evj
VecrIvkK3HWjyzkPAG0sqnRLDkm1RuK1GyNtU9GrU4VVm8aaEUNQBWRBBA+YmAgJ
+PxBfZ0qL8hE8lrim86Bne+KvjNrRfrLMf4qJXykuO8LSrwj4BB5fgh5OTICvdg9
rK8gz5z3rERsuY4ukyzfbycdUzW+wHuph9uBqkdFG5/ewWWN5z9NmQifaSv48wGa
xSWMCum2YDkxeJoxGBtJQujbwFc/DhYvEWJq0/lXGzNMOeERR/wI2XZ6BA9ECPPO
E62zwmW9xDC0lAp+XPHaz63U/lxd56B5/0GBxK+nYE6LwbrCpLIn56u498d76b3l
bX3dS8D7MvQF8NrotKwbe3LTsYa9syYbS2ZPfr7OFuqKJsy85HNiNOSaU8nru9XS
vk1f/X5Q4zViTkJx2NlhjntxSAmobJ5YMGSvPOFSdbxUxgEttz2mEDgSkKnr3gUL
KlkMaMGpOpb4YZ+pzn0qqg41LtBSz6Bk25n+WR5885wOXeu/k7Zt/B8bAGgrJamv
W0ZmJ7kmTjbQPaDOs2z5pckq3zsmVAInk3+YBGDSNmcYQ/90m64YiDUNg3ocoOy7
X1MuARJgnSyZOQdjBTg8MUes9nuRo35nCgBYxPhEYVtan68a/+NkRP52PFVvwkN+
OeGMeSX84pqfc8DBol5ZN/qmqOjp4V0y1JWmJ3afiwTH5Bd3D9aNa5hhRPzZ6/j2
KyRArk8pAmHNQhFfRAnhjjOviQ1pFclR/1GNH6+xejkquT0w8Hu0axDNlfPExaMJ
MEvrhCcgRS1r7suhdpWCnlZGcdyOGao6m7h1I8GUMkWALvLZHhgpp5gyn3XMBIn/
Q/HZGH9gsdyAFOc6oe9ct8vcSntx9nZBpMiVCQ9aLUgBWDQP8er/IbMG4lPxbeKm
Lpd2jHIo/NWi6AE/vza+wjSQNOCagovnuveMkjSwYOOOggYCHOs3n1oNIS81dOoc
3l+t/z9xRwxCh9+svK0pzse7WheeKtoCcgzMuyLm8rS+QMosXR9mqR+FNe8K+9E0
w/QjcqzQJnEWH4RjH+IvOhkxmxt8CuZXAPHib8s1vWW0dAfPKtKTjjIvCM8ue3JH
5Uqv6yarM7pBS1lT7kUOen/a13Wyoz2Oh19Tsuv6Tl+cAcf3VVLyad7XE1jBRn2u
KFYePEgjhaP9Oemqg2xmtsM9LGQZlRhtx2aSdGBxJe3br5XH+hmrPWjJ3oXGKB+8
0wqxcfSOlUB3nRnR8HqDbpJwQZ123BvuyiooTXbacbrNEU7Yr22+eXPlRgIAuvq2
MGGgUkK2zE5uLA/KCPK1Unqh5wZB+29be/KIWKq0G4T9eCyDA/e7ZRK4gNeXJddb
TYv/XZYRNxJZlR46/DFnSWXE4whzey4F4FS4+YmmAL30h+aGnN/mCW071VR7TgbN
cPRHafDt3aFZKjsB5h5I1D5ql1z8ytsaSi7e+2ymK4uVlMuyd39uyUnPxfDdyIQ5
s6jzBsfbCZK4kIXIaQP5nFdGedIJurjMrxjO82s/8NTIHC3mNVRLq6htsK8W73bc
XKw9G1Kz5mBwsu4bYK/ctoVdWQk872Ry0j1WgDdHWMw3ETgm/AWKaizr9XqAg7e3
edDWQgnq9yfDWt21B+mEIV4tGAAb8PETWTt/sIj4FHIMU8vGTFGYUmAob/N2t05+
NYh7nn9eVkgmk9xlJ071wh5ksh7xV4SA+Q7f9/mZp+UzeSChZu+er3VzXmjyefl3
Wn2nmlSbHUa4gJ+Cjg70YhObln2+lso+lzSiCd337KmfOon4pLWGoLYOFAbBwUeb
uxzC++SzDu2doKXmCLQ3nRmEMV/iNf/0Wz63vTT2/e+g+tdUtoxEiCv2ncLoYA1C
9xUpkukOS2nGF+TcIjySZGaBamMxM6qR63T3AQD8wG0Ot/RjZD1Vm7pWsP+qeoUn
+zCULP5eieeLg6a4MBEgpHmaUYTRUilifnr+ZnMHualGyXYXoPTcyGcpl1IKwuLG
bdZDk2AEGRxXEul41wDsHDIc5nnNSQbMBYqOlNIFmJaBvU1Qd3xCCEPcaK/FdUEG
+/ZMLp5aAthyRiwMwzDGUHTu6yVaecBRr4tPSi1HR/t0GXWwwKlZloPO1l75r/eG
u46w7Wmc02WsF8yzxV35t3j9Sb0Y+aMoTto0gY1E8FPiTa2BZhd1QYMJJKV3FKXn
e0hOm/e4v1JIvATdbiuP2lzO68eLAzd+iDdUlmS6YJmsjqRvr65EtwKzMNGisTsn
+cQ1qF+3W5ftpGQpMoVwYYgX8eAjMIGab/dYQESiA4Jw5YDs5Mz8TWmqaKLUVR3E
TlwP3d6yKrS3Q2Wq4CstpPJfQEWqKYx+l5nzQ4PEkjdYRPeF3clt2RX/5Rwnta0i
cJB2WwbSIjhTInBALOkXR69GzmRZ0ClULg3giFbdnSwMZOFxYr6BAfQ957UFtVrC
2bXKT8b2hOIWBOQvcJetdAN9286gvZlX6NnBkA3tcJDZYwvsbpvDz6W/fZkozTO5
PY0wavHSSwfqQF49geuwW5EVJy8cYYOKLXwnwFy5nzU7pfVa7pVZ8uRXRkC51ExN
3RlQrKr54OM5RCpeIKFeTJ+RUFk2gtvcFBT7Kq5Lmqs7KcH/9Mgv4njrfURZNuwu
w6euZLnI+brEYqaHHqh3ZzLMwMcnWxTR85KW6o0zqx8OksFYnqgOvWqeQjDXE1uK
XpsIdxeNtS39ZQ3ZMu68sTWVldDT8I84yrD0aTTUyG3cYuRIXVwiqcZgaTPN5aeA
MUsjdmu3quTuDdp8sICRoqGk2/ONS85VHYkpkiJRZFIQvzdv2o3qtKgsRiKjPfa2
wGw3FzjITbUARdYQWpi41eO8trUMWSpxaG40gHOEsxj9LhwCOk553JST+UdxqEcv
tI8nqRbRrBU+Co8+Q68kS4p0zrRwjr7mcY8J0ttHdww8bM8KVntQACpbZtmRQiaS
zL2gKnAJL6+Zpc1DRVlYnf/E7to0vwDVIko2yIFkQiYuOMMRhm1JJyjTHUf9SHDB
C+PCVBiCeIwO50WzwGixamh33bq9JndMDW5SaaIlfWVp/k4Cg/84XtXjNsi8cuuE
Px6dxzs7mnxgNHXWspuvkXLquXcAWzZp9GqAr91XWYi8SRZizwBgBsCTEcUN87o3
ULx4UM9eOYkoY50pFihWIRHYu5C33sbGUzAsmNvLouLMCF1AxWGJZ7T9v3XL0VHZ
wArniPLUDo7aPYk/Do4DGVJFHwG/0MyPFJAAXc46Q45rlmyXDyi+mXlRYSacuEBy
PmTJsac5AE3COB6UHst54G3UOM5pz+RP8wJl44Ga0Fm1MqcmcbT4wj6ubdVzqSff
tgWJDLIELTbW//S0Kn1/TS7riFp7r30P6KjCTs3hYTv730gtUSs0bRza58qPr+IV
aoEVKp0aTuKhUZLSKvb0ne6ZbzIPN7CCav2iY/8QUAL1g+yTd7q100pPwsRfyQ57
jTkAk086KaBwrpr9Vs8Ds+SgihHX/mw6NY6WGDhYgaX3WNpnNRetbQGqBWNNzVk7
2nx8syMR0w6gCMLAJ2u7ocOhctHT0RHq0CehsmcPs3UsOVsNDmAetZ1KJNxqvh+u
PIztVivVMlsSZKNDY3sZOHGxVDyZduhJWzoyWDfDwbhjXQsTR3rtoggBBpBNH0Cz
r3xvPenFJ1hM7gwKTOiGUpJhDSDw+zRlNIqcIb3aHwwe7P/OM0bMZ3rkKem1dDnb
7d4afklLFK9/MfFUh9gHZvyGlaSRQ0OPW/a+xqMX/fuVebbEGDxjOjlO2t1xKPg1
Mcqg2r3absdj0EAEf2ECZ1tlyohnUrmgykIM9M5sWoMX1yRGH6BNIWSR40YEijnh
iheAphjWflVFedlgcW++zBh5qbqjebJ791dPbaJmr51Hx+azK4USdeKGa1m6xC1m
Lm1Btp4agTthPcUa4dT09bquH7rt2lh875QMeXHwCzoj/WBTIa1/KEgJUJ8n4O+v
+UCrhSiTa55RK2d0DD4eDBcnt+JuoZ0ZqCHZ/1cfH6PQocq33xFgvpFnxYjaoT0q
iFsZt+asZDN+bH5RES2zBmgoQBuRuIvOqYeTD9y84fihlOsKn7xUGgl7pSnvQSHV
DTxweuXc1+60t3+ytkleaffhX0Owei7LB/yB4a3ZPhuzOYS2ndQxpNAvsMAOcbDQ
eirHRJGwCvx7cT3FfoQ0mPK+Rt40exNfnyy61pkdRKNEo/mFPSTkbDO2G7Q2UIFt
1+UZWGOi4QA+698so5HGgJDm14TkIfrJznSeRVAKExDU+dHtijaPw9wGRWITJ5fP
IIv+fFz7UbhkGm2Bz1rrfMCtreRI5QHRgYXGyYC2r9GbrDb85BxyJGu6epSxhKbU
BOn8jL0NHLipQhDaFM7CIcytoltsOPi68f3DcduT0XLHKgRoC7RREOtPnoFYaxTI
Mo18n0A2xi/JwZq+BVUiU+w4/UaUpSSMN6z5+6JHozx0CgNjoV8A+MXMDw2bFVy3
DCqc83ALwnkBKw7LcEYt6QpRd40R/ZqCAMSSxxc2X7SWF3ItHM51CYW7bPm8kREn
4Ys09G9EGKnejNF0wb9TSWW0p6fRsiIzApNhs+5MhWmNZt5a+0EHDmqFa5RAbZCS
2leMoHMjvV8U+/TNurtPCU11600hQqlBNDRB9faSU2lhyd71FufxBdrwY3FRTGJ9
cavfPVh9E4i7SHx5d7eL6Ek8JoMKmZJjabxWwJQxPqR0F5D/g9E6jJxsOsVqKGkh
2KUw1dR/qf3eL9680UljLT73VCFG3BzpI3rBF9rFxpTbg/23Y820Gh1eHMWxS+3o
rUYCpm6cwPFzC6RBLbN522RH7zXSgVKrKA7GAayOIrhFww8XyjDSQqyMWzJRzRlL
bGcz71hj9Eg496/2L66PzryF0X6u4jY8nhT/ItDhy5iV5TCpMRofQqpwxV99oSeb
ajNlezXsN/QapYSB6rbBgdTEq8cXF0x3pwH8jJXOIdDHW4omsu+5Dq3jEyYQMYpc
7MarOWJhS7isL9rfhpUju3VJQXEmYjwVtvr8rVLPvMLNxnPFAYQbnWvjjFG3T+Bi
cRxN2Bbw7YlPuCQRj0TTGFmJWq8xdYeBEyM/zBZuhpue5sDFOF1q30o7e/gEWHPH
xOT3/arwvwJhwPMMtF0Z55IvLm/Uqal6OScG/OIZ9/j3VEF9mlFraiuzGP8uYVKb
II63Q8byK+pTuhWmcNO+5HjHRHcoe04ecGqPhBbL+x/ZTbUgzTdsdJn/P3fttMd6
hfPLwVZj2edeyiCEADIYj9Tm7D/Ztf11e6Ujz7lQSRHPAq6GTB6zTzm98A0/IazO
0zBSLuD84I5/EX9nknw3DLYMuKwqC9b03lNcFANMzXhabbUK1SKjHp2ZhDyd0oGI
Wwr9Bb1IBnPKtpvlWxCrVxgadLPDBDhcO7ECGu0McdrIJwW/HRjiLaE1/qyGaRXm
vyPD69qLePPQgctE6D96vzGfMH++azb61AxQ/oKnqOoGegO6l43prKEAsXr+dYYj
NIEXdOAWecb9R9y80fi2JUJ8sa+qGyE0WEts8t7aa54khVVVbszrS98cJMIgeFIM
1j71l4Rm/zVznw6sMbmQaDSJKzQqcIMBBPc+RJIcXEAfypU5VO/j/YhYWY00uAIn
f+H12GtfbvADpVgcBNRwBNxaRQkqvL3kQrszVYyOh9oMKVzEJkjk4K5hpb2oOlTX
e2sLoZgOVXAnyDX/WwlmfZQnkZnXah0iMtthusUP3IspknHhzUc5FDGtVrA8kuZv
pfzcCNcOglFfe9BK3gSZ4oKLYmsEDBQNWOfxCYpjoF2lrwbLUWLW1n+hM4JnP28k
P9yHzt3m1GJJ5NpiJBLlfCiS27Xqhaw9cQIMWFloOZvrrdrf1SC3fILFTnDRQ4ZZ
83TEGWFA4JKwa3wkNxbt9dddo0k+9vuxMvCvRjWTrpDQvTt8bYtS+DnFqeqrpmhD
RGF8yqOVoYxntcdaCBXP7+xUAZBDe1+NMNh8l1LDcgGQtvkxCUKxekwst5fSY7V9
V0JRrIiOZSEnij0CLIE4D6Hwl7vnRy1jQGalN/fjcARGs5JRwAC/R9FSXnRcdwid
67SQGt5+YWY1GwfK+wRTJ7bDpvXcndo/WHxVCpmD6jv1aX3/kr7i8pKe0W++l5sl
ClsRnnxCl8Kl1SZ+tzCdO1Is7p3x6uKe34z8hGQuZC3uIrzEqDux1K758bTXKjNQ
+w7zGODWpXpfOQ2k6bEKwpis0W71PaK9t8NngIAboJveaVyjM8O4ip0kjHPydwlm
Yy+tzcVtL5XwJ26dMeTkSRAHiO2CpCMcMkCg7Mz5Akr95/NsW5VavJVP6q8M8yWL
a5gFuCY5+720s5wSkT6DgdN8dpqLT3zyZpL1+sgaJ35MEmIlOoPcVAja0JC6iunl
M6e79u8e06umwNievJaPAiKK0FmS7/8uozCcO2ZmH2cSliy13VIy71clWgvfRy6d
xH3hSNWFmsqQv1ZoSyuiAPBM4gfUt5JQyL37THgzx2wqnfGglVGvfldHWwN3D0de
fYcHV1CK7Ac+YuyMchLrNti7ICN3ajm0vR0cLh0ksoiQ0O9K5Lt2qDfyvIY7PqKV
fpggNwe6cDBuee1TCJ/EdasVw4I7I01QMobvGVhsRiULS6MzMTlLi2e3Prfgg607
jIOM1Ncp/X2OcljiGrgd/C9/rS7TyFw02bKohusdt0YNRiBZIRQXCKZhTZeHVaKo
JZoCNsQDXgcUr2MgGRWYx632t1HIBBaO9nTpEi8lb+aYuGXNiYKtKyOlNd4nnRxS
bWXba+XtacY3wFxeg0d4olqBmH1xdlpHJAwbu5m/r16RJc3ZJi5Cno7fcYVBMBwT
Tna96hSvLCGWOwM89V6S1z+zY1eRCQBhv+dLqlxl0GHibTGrE16Ob9/Zs8Ozuk4x
BZ1swy2Y0UDyEka2otJwof+8RFLmp5ANaXwXY14DytQOnuGDL6b0v19IjlSsvQOO
qWcjlT3d5k264GE3KfTCYtUVoOoEY9fHYSVhUhtX4TrYS+BfnQloYxB8ewYAanBp
uKDF5C3PnVr4waTwI5KyM6zrqtPMC1WZo8Dr6ME5fWHJg8tn6IgcvXG2R30obnVb
ECi7SO+c1zM5QgEt8kxGLrL9YY2AUKtVjOsbxYNYdDy7X/wdufEjsz69HEuQYWhr
WjyoS5/qsZbeBXYwgZKaVh5fWLn0s7perIMjwAd7SStORLH3X7yxDAWoOH+xmep1
nRmrI+000xu/IBvXuOpBLwahZ0gHKVvdb09XsCw8vV+h60hd4Tr5/8SWy0+AfMdW
g18/op65V6WxdfXO1iAxsjHBB/nmqTjQMdT4Y5n1D0f2fZ/E7lQhPfieDeWUp4Qx
wPUFVw6EmSnQfnbB2JqvVmMuHLabyQtuF5os7Q8lRzUWVC6ToCOZfNnE4Hv+SA1c
EjcF9jFpseqB20mFZaMP8aSiSIZBFj8BLOIQWB3YUvp6oio9NLXNy7EMpBgIOog3
dv9FZNwKbJQHqAzsVH79//F+02GsWFFZ4yQ4H125dq9a/592WWCT6l2uR+eDO5c4
aC4OwCf+W76qtbAyiSQp544YrB0bx7PMpt96uGwT82JXI/7ISFlv3wxz55FDKz25
woAgAOVj/VAcELxIIeJKrYqAXSCCEtm6c19GCca2Uen82LI995xF6LwsQleJmrWX
vyh0c0bbpMhem/mZUwj1oOFrh7B1G1cptNuBBKT2lrnXNFY601BeXYe9cuGWs00j
VfvHcUXy+cjgDMkHA0xPaZzw2sdhtEfxe6YuLMa2wKgfQ4digK8nlp3p6OiHPBD9
cyGPSlAzWw/thCjz/F0rX30dMq5Y6iCPE+rXAuyvUL0tPJlMPqjusT3hDKbrOg/+
HcJbC3ZRL4FaW1gOlLOl1WYscxmneLKwOgA9LwLchXdr3X8jRayChqfJ7xy6e5yK
5rMj86ZCEKe6+53IkTa4z9SNEvcfgWEQ5D0PAuYVE4iDdokTXK22DQh3HEnw0Ig+
0c+hr7WCWUPd6KMDewx6V0VKdNsCqA14TeLc/mCR4kYs0qNPzv+KRlba2P4TMC74
EEOD5RZAs3kwdvRYG50C7FiRjaTpCQ9mLkb/aBd4D4Olwz6luKwpjWDP+o6BfADJ
TOxYjJkMbWIeIIsw3BwZaYDlisDMWV1TV2gq59mqO2X2sX1o+oIZvREjFC3X9Ez6
/W3V65ryCPsQAM6XCnxJ+SLyU6ApseGNO8qHbdXF4pQoZpXTQl3hKuRngXbw/ok9
6uu3Ai5LVPFL4Uylni5ZueQVmNr5YQLQEHg4nLNsgYYyo8t/nCe4kWHJlOXBCALt
aQ4DU9EpG7e4bUbeYVRHrJ0MNKuK4iU4lWolBTX8MabYnXNH03C4B97GVDJ4z+c/
UaZDz37zYXbKdqb2OSLjiOd8cGX4/ds3YpVc+Ycpq12hxpOsRG3QLNMIIg0X/64i
gQhdtr2QBuReK2i1QHLI7+tZ1pHACdXsqI/YTAA/nYtcpgxiFaPWfxFxAH18QwIX
mUv2ZdHoHvxv+q5wnWQHx6D+OyaES+6C65Wqpixhe3HBYEMezlA+O+rNAEnc8ppP
kVkpSWBARj/gGc+6rA5AQl8Tdp7dV7TfSw+spJUcL/4Xby0BHVTQr20kwzVBvSfI
xoo7fcJnigILmhwq8QT1AYRvkRXSFxQRq8EW0HzkbOcH+SIQLnirrCY10lcVzVvC
BE1sKV2Ws2krfN0N9lO93pEZbg00UgfY0CEXIbLKb1/Ql0Uknv+tNZZuoCG6MbzF
mktAjt34PNb1jEVg5OFU58EtPV5mDqkULOSuHcsPqjWynDToWPVwSgqWWZNQ5rzA
xhd9sOCUt2OqJKgOBGoSLZC51LfSjykXdPHrp+ch6UnUg28gvLefiX+S7yGMa4i7
P4PlIV747mlkzbrFVxsegSt2cluiQMbwiaOrBjWAnbcLJtbPjtk4xmBvtVyLvfCu
m4jjgKtkLNY02RliaBO0BMXc7r1n8GATEbYh5MTZ3vgvK75IoSgn/PIyl9FLHa2r
qin+NeOfr6sJTCoyPPKR2NJbAn7lnWnSkCKkYDdUxKG2L7hN9o3V8mosEqoy9pLf
amES30FNBZ1DUuow47HRi9zpIbj/KkQoaPjo79o4b1h2MHF+ggLC72MjaFvoNvYw
i4xIsojTxRMdoXuEAmROgT2jN19kSuYrW79+beJubPZcmol+54lsQyWIwMxNjIpo
MYYwIqK+PlobBPBSCWn9dfv9T9WJdbEqoyp42j1RWUqonA2nFAjc9UU3eECNra2b
rlYkMHsxJ+69q1/NGab6g+PC7H7POgghS/JFSROAqwybmZNvwOvJt1A4OFM48mfN
O3qZK6etQroc3W41kerNCufwBA0bxkLxlh2IZwm+gfJ//OKyK8kb3glgKZoV7cQq
UOnhEtFxql+52XN44bHFiNPf8QFC0QEwgA6XPURSEqlKLK78BY4ldXV2lwf9xMVP
4io2LqJZi1Bp/kfJXQ34fxno9ODFxXKFmcYNOswWa4cF4/n4vol6wql5VGrYwqVb
yGGvI2ozgvB0LTqfDy7T9RTo5yqnvPWFztoRHrGfUKEuGGtMe8KKMlKuAXmpyyav
P5lwE4Kwp6zGS5G/BrmMvtB7iPsBJINNlx6DW6+ElM/KpyVWoPdY1lxvQDWkedWm
4cdAKS6NFok5XAbOKpX3A/9e4Jta2oFX+FgJZIWIpsYMiI3AxontWhOVD7jIV1z0
omDMpxBd5l7QTIhkxzEMzBy9fqYnbl47VXdciT3BTTBbPVk6+3w1UUkf0VorYgvq
GBLhMWJl5e9aOPRTu5iQbtzruIk5qNiF4HaZobXynwvvfidnjlR4gvOXxgRAIh4V
JH1ubUWPpTwy/TaPPs5I4A6AO3f0QNKPdsGizrBEMirLdC+DRek8PnINMeJYKgmu
gm9DCwqeq9NsQ/Ckvm72id9iUUFM4uIGv8Hx9SISOx9zrgUs9iQJrZ07WFqDkJYC
xJNOd7j2XtorRA3UhRx5t7t+Kxy0XNFWYFDx/YhXmzX5HGStxxh7k9GR/pryby9n
EARhz3Cx2sZh7gJQxQy8BVnppJQTobVY8zI9TDdWx9h5AbPFzThbFhMU2ShWXsUn
t/uOlCWa426GY1panlgEpZvBSj57lgGFEOsI+Kr+0BGa168LhkPCfy0YRuxfZQIj
iA1Zxl3bYPrPl+MuL0RbFA5dQKlmvP1Y+e2QhR21S/ERPDsWSNL6+Upd6uiPQfYt
HhaGrLkVMEbThZh7Lz1g3MMyzBV5qL4Okm+fak/X0ORAZBHOq8r6DG2iBHfwMD1P
CdfaA6Haa4kCVFJ8SqCTHKpKbBlZc1ZH1lV5cHlQGviA8zFVaAFqenQXedRALWiY
xKE7yApxWnH+G3+Bk22/pItuq0MHRarUp7Hx3Aa8ZylsSYt7XpK39FTCEkz86Q4q
20jF7M40P+KcxKoqzeOWy1Bv+pdfTqEaZM0ghopXXaOG0MNE4EgABDVwiGJWq3dr
ZMWl0xSuzjvFF6eCp/a6ucFiM0vUGqUQXOc6KtY6+YyL/7jYOIaZnMUU3sP9krkh
WRcDbEUpgFbKf+eQHVJspudHs4qovPGnsCAe1GAiH18vVFjbNXJRWKR/+ZgZgPwD
OU6mc+e6XIr6Q3mrymjGHSg92Zm0gM7FzkyyM3cBfINzheViDXBkG2g3e3uLDhGM
xej8gVSRmbZVhpe4hgzmgGSh2UOQq85r+acA7uESSBa9TYdXmULj/z843Y66PrnQ
G8N9K9+bHZfpPFWoOGjupiG05gn9Es3lIYjyBXSq+btiRvgMjAByKSC0S5NMBYjj
XXlv8f+UxLBllFrd0/YxmRuoTuVAzNXN8G1pYKob+30Rui9sr6Xtl+aAm3+0NcT9
0EQEp1Wh88+QC2qgqiqBQ1Ljn8WgbZv605jB0kIKWUVGqWQhJWpi+jrDM73SahtJ
Ojk9/XpJ4Ydea53/fnzHckJulVs4LWNsOD64+DRadWZL3aav3JBWYhZ75dIWG+Qu
NWAodOuF6HlW2aB5nFw8zG1Blye3dzdsxTUZRX3BJr17mwvlBZd6gFDLrbC2gfMt
1h/DmZj5nsd6gQ3NZVltiWF3oG0fFb5rTJREAKFeHiqFnNPDw5T16oCktSPbdUdB
hX2ziIbtMdr04nXDqlUF8Pt0fFXi9sX+4Jk5eMcehF/Ulu7UPRT0Erwuf5xUfFrl
3fU541+pY9GsSb9yJdEyQqq/mQoeQJIV4xQn0B3Sv4hRlb7BSKChiqY6id+eSjk9
zEgyX057Pp1iKHtJi4BjkV4X8TqDq+PKwSz23Gr+3/0jusvgqr5QDQmI3V4/PdYy
oh4rDaf87xplmAksPfYSATumVE6T4q7JUOXvO3NtOUXzHnFJB+jQll/1UcBuuX53
bTv3F9lWNyRnJ9VvyoYiWqotdNgoi3bXKoHKfLyfGRXejoOq7aDtbLvYzfYaV/Cp
5jnx32rbPg/YiwcmV0FtOMvcWlUu6jfMBT33ydC6PgK6ZKrMpIwvPXaDkeHw1gwI
OhTPWiYRBiO98xsgBzQ0sF/MhN5JfkZhGsNPEGlCtCFsfwA0zBvDnwNclKDU17v1
+ZMeJJPdN+EbogL7oU4KuoE+LH4Q/dCpTE4N511g+BNKPkWa2r41xiM5nCD39qsa
UR0rdf80+k/i7XEITF4tFV+Ht3+95mDaWu9orPTicZDSZeIDNbjt1GSOFf3wf+Bh
31JcjhfkxfNmnALGVR6UyGaifF5eug7UNbeI3+Hw/M9UTwKcfwR8+lIdd0KbynlS
vDkoRrtDmcQNuG4vKyq0a1raGO3uNuT6AWhdWPuamLcmxKGxOovccCEcbKPRftpM
umWSewpPk5dieXUxrdC7dC0PClSsvvRqGggYei2co0+YLSWv0VjVehw0WNLCy9C2
JyaIv2wRFEReT5wwo31Y97IgEFZGZ3no+jt3y3IjmIGZT0qtTJim4wIVnAhGer6/
v5rY0m/tLnvC39Ow++NqEJILYdm8ulQjY+kCEea01JR8bZk7aNT+iPhRFxNlA33r
FqEZNHh6YRUlDf0bP7conTDGTf9r+KksOpGyFAncM3Md7X+07mcWLRjMuJpxfaUp
4g8Bo7gI2DOtOA+NlGx6lJdAFgEBbkpTo7z2bCR30z3z9S4AZHq8Uv/h48mMVGAK
piPCtsFd57uvitUn1UqVDTey62ciTG0CbbpgIoS1pwDOa1dmCFvafCodKf5Q5LYu
qCgKeL8TvjJBDsVYEADqsYz6yc1uSI8RGUch+FPlIYNw6jUI9dogI2jkrWCYv7xc
cfeLIj0jHYoPk//63vVEEsp/QpeKsO6QjdPsUS9kGen6siz31cRQju5w6HVrZq10
Q2V3NZ78XhgKSGYFBZLdG6CKJXrmA4sLStPIuHN1a7NHvSrq5gOZAiJpV8jKbCzX
AMGTzCyiGGGvyyxWueO6mM0D/4WjTTRsAwJXxActyMTkBukNbx2AseJKTZvi7vyH
3kVA6R382LFfMp8ZVgZtNKNSKN8PwWuvPIJQSWWMMCNcfnati9WXkyjTkzZ2VgK6
l5lXQjkgmWFu5OL6dwSocjoQH33nVd8smd4Derqrepegi5F1EVhgVWzRd8Bj1MuQ
QlyiUqhgyJnGv3HQBjtiBXxUkV6VpESAWah0IboCj4sCIgqlWEPpJjxVB86J0HUV
h7km/lDtt/6/R6EIwzv7u/kK4GlRZqJqgfFv0bCXHTx3NfmFhU3u9TKuz2yCl+CD
/x5bvBj7V0j3qcbZO3t4CSiHNlhylS3sS59ItTzWCDf78zMmeGCRYR0HI0OyjeBX
/EuZYE/6cOpCYOOjn859hAQB7+kZV8xAknIXqRYFwlmqPAeCMOpZbs2mQQHfrrE4
M+cg9vEzH6PbQT1rN04oyakh3i0Z3RAQ1C5SYktM4wgBjLIsX9B7m82jn8p8RVhZ
jBX/jinMAuP+He2NGTC2oKw+9m7txCrXAEMiAvC3D8VAx3sGsmJmH0dv7UegY50A
xWYv2VXOfr4TBOlQp1tRJovNY8REMiax+78BzQ1dA+qO36O1o4Kqqds1tc8hrKHP
2ZLAYsFl/0OKaJ0FZo7HwsRWZRfeujz9a2fjgN0Rw3CGOdw4fbzVIV/kF0BH1/tC
7Ops2HK4tRKb7pqTwUS45FPq7uOVJVgVC2JAA5Pbbi+NoTRpdOYvJDlyH3cW9vck
B+DUqZLjAKBHdCC0E35UCElbQZ3bkxyZP0RKElr8viHfqOLtK1YmegIV0Hl01tY0
7ScaaiT8SI9KEcAQyEjBIJbJTPCrwocIuf9N8P2fUyu5vLk8+UfmJdT3mgvecczz
VQWiRRVV2xQ46/KcIn1HgGQ3n5sIsiM4YDLPgnd6ydq4uFwJl0sU8xcDGSkNJ7qL
AP7cZQM/b43dJZJRhBUwbH/fXFa7+XgU3bO7SNsv4QUuff+0zTEex4r65IWXmKeA
j6DMna6ErdXMPhZNFmyWROZFwrZ9OTyhLfDSpEaq9yf5aHUTlGdQqwgXyvfAwCsO
JGB+iMHZxnS3LVDYP5rKarG4W2cQir6kQKD5bmsuj0wdjdtFCzoeJAgCB7UGAhAv
HqeV8ZDR4wdqaYf/EK84r6cLokOo6mww6JGoboVlNOLZhxDmGlNTcALvZCA691BN
EM41WUBs+W4Pb56Gn1kvvo+RtPLW/Fut+8bK7d5m8KGx8l1qtCggqg8/4QbnsYmx
WIyLlTXxalgob51zNAvVihueojzpq/5oBwNw3UAhQKupUv1NKtRZy+4FTmFgRbzY
MPASdwS8T6l6EWvZy2kvrC5bTEjpkxQ3Aqj4MflxgxhoDyKutN5OHbPdBXQgQrNX
GV+lHH6CyMcoLCcktIY4wzlWgD0dxhqrEF19Lm/Ma4K9Zjpfw0wmaaLkcyavIOpB
nPZ1avM+DwXUit69Hk500wcZgUMPQXciM1HDPVbH/dRh+fufAdfkZawZ8K9q0JZz
1brey4Rgs4133pkmJAFkHLL0klQ0XEWswIufWloPJpJO8Z9VK6lroX51Rxv6R906
yEB7ruLgnbb0MJDyqLnjvLJg45q1ZaYZiR9QhQ/1sZtKqvDNUk/JlOQZ33M6B/rU
ygcs43y9DpBJa3EWh208dqSyVh12eEDTDQvnC/mMFqSR2T+UzFaX7CRYfQxJGyIA
gHzskQRdWLGHckWKzSfbo+PkmvGhlJiphb2yXS+qfYYtBogimUJJNeRKVhuKoQml
MJElNVVO09D+0Pf5pIflYNbYp90encAmGITF0Nk+MfJBzF9ZzXKZ8VHTkuEYU9RN
Hb744/uLAVLpqFPE6o5VizOHj5ZphShrF2PNYmx71e7NwKYO8edDThLRAB127wU9
QQDnWJIZ//FjvW5UgfkgSA+l+BLa6/YB/nUiREodfDXLAR6ua+kk2QdVI9fd5pR1
R5YTCxzBBAigtLKuQaDXV/TTDb43RlsK/hWqLzG/svWe3xVXrrJqTYeqMv03UGLS
2pF4/4QxFcagfw+mEQKD2IfwmlO34xRcZbPlrspLEcKopHA51kAfh4/1wEqtX2yi
KWSgP2v79o6KArBEXsf2QJW6rxlVw2XcCzOjKqa1I8vWEJEF4BGDS11yJ86U0xC/
oSgLIc2v/+DaN66B7vgVd4bMxC4AAcUzICtqu5EuDJDTJSBRIZPrvXTi3/rm1xpP
PsQCXjP/hGHufNxmWtgNKCJ0O4LMUAtJ3rzx/1kMoCYoHxKSyskU3Xc1xosHrbYi
mwsyC5wd5Zy6KD5Q0QwFUhz0z8LEr0si8GeTpJ+/cVSV1vsKmPn3YEoUsI+Ey/a6
EngjjwtaKs8wULde/TQaIYs6c5FQds45rwGo03Huz/jEYbPyz+de/+n4yGEszSju
UWrZ4T6YaY4g1qNyBm3nTq7AzpKICQi8/0zl2XxrK4TsA1sKWWZXw6Fg6S7azLcm
PeThsA2L3CAZmO/ND6m+yfmYRPs9IpCuaa8SJrXQ6Wzp/F4qExJOptW3He6PtZqS
ITXWrWAFKAh1L9is32c+Nl8sfI09nitxCVGIaxOLz2dU00htECazU6q8j70ANSUa
cMTiGJ7DJQIKNCQPiQQRRm/pZMSB3WbuUiPZ0KhkDbBwORPoNzSWQEVC7ZvwFR0q
aPcq72euL2hSqgvTS6WI77bBi0l7LFOV4HLiNs0KnRtPwYkCWu2y2HL4iTnd1CRC
MsdqRuQKjSIHsyRmBZDHtyklkyOTUgI+lRxXEtAAdgVkINvVugiGq3nGH8g+Xk7g
rcSZRmcoB3SSrLxW9/gRaNoxhaR7h8QQmDD7Ou2kDTTupjFnEhkjB7UL2ZfGWWDQ
gArRnREb9kpQkWvSxjTnwjBsvRlnR078V8ENbyoq/XfPEnTyLXnIr8dRNd6MJYJn
ju1mFk0CUE+IbvhY75NlZ4sdYEuUle8BImXXErhzhzT9T8A8nsNybzQj7gDiiYEW
YEAFTqaV7pKNrKwe96YOoSUi0elprOUy+CF98fNa1KM2DYXwAtf7Y0gSXms12uMG
z3YxNmN8851jGW8rVLQ5e7PhASVPLbcnswrpCMlMhz7B1PWmiS4ik74XWXfpp3d+
MvSeO5xmJ2W9NTRVVHFeZWd2BUvZzfysS8tZPzHSvsyQFWn4oZBlDiJW9YPot39N
UeGRI9imNlvkXK6mEmnP//FLALdG5/Qknp4KCHqalcbLAh33cxQdi9ks6FAAFX0u
uO/+GWtMh0q1ts9gwCgzWuDir/wwC9BetznR1NQXaENZ4ayprGeJFLIjJKbi9PuT
erwI2gPMqpymr9S09UllA4499BR69X0B3OYztK02WMX9KxDXsJQkixhsw/QWUUy8
Ghy2yxfoXpFBKyzRFhxpLhrOcc0IekpOqoKEqTADRSu8X5neNX7rW8x1v3IAGXd5
pRy5XCmKeR08WhKjvj++Y07wppuFinb4HmLGY4O79SgBlSI1IUh3uPcwYnZ1STSn
IiB/fWk7tlwMS+X9MJoBBOJCjwlHS2Fz2aYByMPEqVxFVpX4H2OvGfHLMAaCgBt2
SwBPQsf/ucl7HCUetwO4gs5qs7fMS3yNeVWnV6F8+4ACo2zdBmvNLJju9xGAw+xj
NJJ+ufObpp25OdozekuGl0zKkQWQrGZ/BGcz+rDT5kxyk22uM7uHv19qGQM7kUR7
jsJLxXrnvuAeq4Guju9ZtdTI8ke9YhwLp4mfaWb1kCGo3nT2zQn154Tl/v8hbqtt
z0Ykt8gDJYK/DNC1eJDpjJeoU8gRqCNa5/oNmkf9IQV6i31he7rMrdCY+cQTfzLc
x/NVoc2ly+qhlxYN5GZIYd8rVOKzknHnKRYv4vwFtDOCjlt/wxz93Xno3dYPbfZH
Kc+O3687DZIqEtSZ5UyKwxXBbyV5G1UcnCX8/jOj+rsWy/sQfWAVVSrv/TqAUhVx
/N6U+uJuaI0J+zrwRStg/E44upvmhkc42wo3QI0SOHnt89Y8Ydl73SvgXUK6ABnM
dFC2rcjA5W6yHQR3ozxZwM+snNM+HhFPmrDIZHJetrYPwlIY+GDUXudQhlViKNjA
es0q4mX6MzUHac7n63+yHZch0yDyXyFFrgniFg5PG//q5y/t9Rf5oX3G2i7vPKBG
EW4zhPMu7QvwR8hxiPyCWt5jW2IgTNn7SsDYD1bQy7fGobRmbTWNGMPdfBQv/b1m
dIv/wQiHHUgnnymVXVcYtNddMfZr26SDipKcvupTZaHqUaXY34ESOU+FvwSoVxsE
SbA1LJQ5QYuR6wuXSC8DRVXZHQ0gBIlnY0lZPfFQj8pi57cXnPxfQTpoFoghpGtD
s0rQ6hKtP3CSaSLhDHwRF7FWVqncQ4QFXEo5+MwFqfrNW2Pq6xNJ9FFKgVESS/03
QJXRK7RwYSQZMD5Gh3KSqge2Atijt8PzcfLkKuQSmvGuc0n7K95RHL2D2btgtxBQ
+tqggzPbjEEG/1tfABlG1+qv4t4zX6frAYC0It1d4JJza03jw3LN0ovr7QN6w3KQ
rfUpx0t01pFW9OX7LXaJilM9LIuSBuo1q9Y/nnz67KD6cychGvWevdkYFXF7AFrl
t07VtiLH209+5n/fUJn2/omKZyQaJyG6eeZ/0GgLwi6eATdpTZkPuSg7eXi83gQ8
LrzSEJlOtTJVomLndrlFocLMNgwJSDVsI/C2sJPkt+Lt9efPp2pa2HhA2mOiDV6P
8wBOwFdqkSUKn1zNRgB7gz8F8jue3Vmf+H7I7DPR8mgcsOaJprGp/e5vDY9N63up
Z3v59gKIDsvOMedpz6XAlFgShgIbwliM/Ocg5DR+mLH1cTe/jkiAha4zDMemWSE7
8A38VEJB93sN7KJf2c2nKos9y4OgCa+msNT8Ctv6UTSp/y1MXJAq39uz1/u732hB
RX5ytsm9YDSFqxmwmgj8Vl1TyrM2zZ4UxiXWVeX+AWhX5SW5BRWDdgAOO67Cehrp
Dj2DhnxHGmJWJYsfjWerTXszV1/C3yKLheMUDlNVtrqDlD5uUtiw4WrmE1t2o47K
Em1Z6bOFzCQEhFc9bBzzNE/yzZSnWgMMoZ5bFLLCilGK4deW5rBQkMsnFqZS6bqf
ZxHYDeO8DFn6JJDWpqNHUhTnAS8LVs85Aimz3ofBL54CWVe6qX87W3HWar6myAeg
BzgFpZQouUihz2An1pLYWU697KM+QSnIcqhhY1bAXOFGTStH3duk/PVZ0JR/OEgN
XZO2nhobEEZ6ElGIREqbqK0tX7Jo6lxpcrGmiEKFRNLpJ90N4Hko7DdTOyEPEyhJ
tht+mASCwVcTPIsAnikO9n7Ln0ZyA0EoWpqB9/2omI/NWBi/e6b73SrbzxzTB/7k
1JeJWn6Ik9yaREIbIa2F3hKGjkQ4hkYdVUMj2gXLLhDJXkWpDpCI21BL5XXR9imk
VMIuJCmc7gHZzZI0W8yZ/n4WAkSIKySqwyuisgXEzx5g8s9BfJgbnTn9P4slQrhB
XYcBPK4zyGKzMURwra+RCggJ/xO8HGJGVDOoIQXJdQclM+OT+c5W02KHYVNDd8JV
YGCpY0z0UKKJ7pLD4WWHQ6ytbjkDB6W0tsGhLYcJHmXm2FTdyMwngCGMZ2cOVOE6
TqjRNf5hUCq58HxsWQJ2vKkQdAcudGBYuECZW4b0dPwr2kZBCAf3cxxWIbj54p8S
2Ag3BQ2l2RFBpfk8hr5yyYENiH2IIB07EDWlx7/5wGUaxGVFH41Y77dFdJMVfHtY
rlN4O7WvX7DMH4cyWabYEtTvEipYFf8Vi2erbGBs6AbMd+OO3mvkb2qCtFZc0mRS
BTzL8uHuBfflmzr37mt+fz/ejCkdPsW6nwdUDmA1ZlYABsX7Ld8iBFUUD4xj7ilT
NSAoLveEtmW2uRDcCHmfQiYUuK2mqPVb3yNNv1aB7tmYPnBQXS2kwOtQUpqjIGSB
a+5fne/gsOZ/6WSxPKkli9BaYSUip0LYTQdw/J4xRvYO+mn3pDLxmWzUXAbFJ0dX
9g4Km3f3DiZFugycKaAgtd7pgBzG7Vgy5ibOG0gBcfWdzEMMBCHUo9TPRPQUkzZs
Jdxt0UjFpwVgkXSLm7E+T5fX08dRxEeUy5g8q7rEiEWwTgHE1dGjEKeUZzMy2yDC
3U+b0F6WIPlDQKGBFnLYzUOFSYjV7pgOPGTOwl2ZmCOl5/dUl+79Qo7/5BXDAILN
qcI48DTimkIDZ6D/YlyZhr2+d5u4Rogp6+gD3w8gU9BdwFwXwd8vLHXySMxOAS+M
k/Ok2xJomWOPCrJUSC1iE/THTjOui5jrQ6UKdHf0r+GJPHVxACXESd5j2sazUd3F
AF8BKBwrUGRs6/dR2ojg8cIlLJvCNxJ2JjioZBPlgb9xa4PoLZPvCRhtnoeeMvgk
2czGUN8VYfJ67y5vfzVYCJ2wqloGplV5HyN7ezDrvmTJkqajnbUTAEvzZc0xUx2J
rJI/BQkWtNzkiKd9tfjCSimbBjbpXGJ/h5jw2esIiocGzWwtY1nMPbSXCWxfokee
EQea+nkBZnaycOIbOyKT+YTkb7moiIKyT+1KNVSby8ombFSU+jBC6D3f4lqygE0c
4BIX90AkMKSnbfVKlyFRB0LSDm4CZkw4Iq63XFYF6mbFSD8bkbr57hWaW4FS3NX9
WFBdN6E2rb0aYp1ylWzr4sfXmWK8NwTUXYxK5PmKhvo19fsFtVxDl5QRhAcR8Smr
O3DHxbx+EVhICdCejQh1lN2owO9nFtPkQjpZwroxPw9x4kCpuavVLLex7en1nqyo
uiP1uY3fstgW0pEWe3twLJqPQjVy0hSvHh75tZouJjRL4QZGLcZj8ObAM/1ytHET
eEBtzwrGUl9NU96OgTbwA06E7zLE0e0VH7vOMCqcJoeABOMA7Ldwt/TCwVbH3MzE
m+pEOBs/W06SyW3TEudZphzfrgXWSQa9VH5I6HNd1Hk2hggg+z71pBiwiRpv2pEn
xn+mCKctf7o/WNSC9Ocrevz2+5hmxqv6hWFiWUJVaZUdTGXztiipmwP7s7NUl6D6
AwisG36cnozw6qUbEBPVGm+JkjKa7+jIny3U90nFpDpybHqB73+SUM5M9ry98nee
l0nVOw5LQAiZAsZK1IQJw+9cOAxs9L5zonkqT3DkHcDWmrMmE33Fe4/Lyqd6fdNZ
kt0OvUULgMv+r5Ui3lZ4PEMRjs2CLh40etLdUgpYsyRez9uwM1L1J4hbQMmtzkX8
Tom3m5ZCDRNPsH+w9qvgnIi19cFP4cbOzHpeYrpx5LnwZjj9+AFMDZWnQpLwfCv3
+HSg6eKRVz4DcFGjjmVIqshW88RGdcz6A+RkWhfG1AZsivwYeHY5lxixpPdmHs9d
jj1lyKg7zDk5jrFcfYshjHCFQUH0aYXpGxuLdc16dXzSRZG0ps6tWuw56KEJYP+A
fIpuy4i/nbWricXGuaXZZ+2TVqRCGxLfPseFsoauR+FNb4Nxd6p6ng+VhA3mweOu
kub38/rYQKRHgmXDEHTgf19XVPLDjhya+yjM/y823N85asMwALddmLmyZ5GAHWz4
EHqrjvE7fld/2d5c8lTEiWfY6d1HycWmybSngguxkhTKw2vOJsnDPsAA8QgMMqfJ
0h9b1q55TvU2yV0lZ6mda/p5mgcexIduNklK/oH6UZSFt3kf/KsYtkn8IzOlRhSz
k+iSdIxBr3ga2J1CC4WN+7PHhn1FO1+S9iJWYaeZQeXbYbW+O5mnhP/Kt7bwHVqP
qpi7lkV8ujCqKEBPnUyWkw62/OWBx5YCDEARXl+ajjZAwdrEcu36u01o94by9/d6
zYVcCnRd+6oHMl5Kigw0ogkH+PItqVWdzwcwZuxEGdXULHS1BiXq0N5T2P73Ivvk
PWnOxgT8sZ5zdBJQ3P+mQkZPgta6+vo55qc5eyUKU53ZGH4ql+hOn+LAYFGu+QGS
OIeiAdlPfPBkZYnt78U5mBrxL9AgD75+InoNXVsv9JebxJFxe0h+nLtyv/lBpfGv
zb05/VEVNuk5kOJg0BD4rIx30YZo1YziOgH2V5Xn2fnGpd3Lk409AL8Emp0ZOTtM
sXxJisq0lN2EC8SfRCHmlMCFB0LeHN902jomRiMZ66CtdtINA+1TphiEHE9PTOmp
PtTE4r9DNw0YognKeADMuBpzirOTH5GD4Ab5WMptJx0A4JVPrLphnIMUYfdbNIzn
aeaRMypimQOJKWMO3Xd+fD3qVFq6roMWxJQsTwrNJZxLOQEA7KqORrAGFtByvrCz
s2yD1OYM+TWl33eeSaF9OTWKvp20AY8JrRHSwcge1fR9n7pD9dCvFA621qPK4/eY
pibs3lxVrnT7uVwFZEUmqIYfCSNpKEYAmuLM1AbSEOezJ3uiDxloEu2Z+FlT4LRf
NNKV13X5TkAjOo2bCewR/YN+WgID/aYL8Dc9MU1Bf7/f35fRr86TDFeD5jWbh37D
8QaFBPivlZVNXSxdUOG4r1vR+Sj/D70fzcjIu2OhYugnOd58EhgGj1bjHjmCAx0b
GJsMw2HTqovX1YgcN3bmpDzo3CaaVha5eGvMU/f7jd+RJVFTk5sDbWLkB9enc3Ti
sWof4FwHoTwbdmqsDTrWBgigJ7CWBxaJopmamSzT+e0ajUVaHnph7RTd8deRAGAB
T6W6OeyRD9hmOuTCPJqEOvSyWuQh59uDvORk6XMWFa3zlFnNJnxi/oy9FR9N+dIe
fhBtWJicm9Q8PHCMJ3gIwg8p/1FCdj/S3TpejyYX9jVZvI5jY4EHwh9/y1I0yWNA
XGuYWxDMKF+29JHvHv8B1UkZOnW+81wEQNqP7VytEfyaAPXc5OUWuhUUiAl5zhWl
MEMifntc1qgCUOUCQHaH17zOciyVyslRB9aF46iOcxNx22uzYj8ZXvvQzOanrSyV
PocXTiMXZcw1SjENHhVe6e/kFphLaF/MSP97Kr+1J1RftL3A//c+uBoxNjt9svyf
GzY+UiOetYtKFB78dX3j3u3nQlTRnjnevIfHOk/DRsafNC+xwfbT8gbBbtCmC+WI
QGuhwaW/+/f93n7zJA4I5v4zFGMK0+Z6T1p+4ajkUw+rWdHDGXkwevBpbb2+9ePn
lqOrydznLpUHXvgyZ6C+XKJnc/FECAjhWx/Eu7DjlRfuwDvGJMgeG+VNR8qQg7d9
6XjtvjaaJtNkXcIH30WsjuRNo5qF+pE/raxYJSwloxkPD/hb9Dppve1tBHTwb8Ts
RsKkT5woA+4DejmG1viFdaLerkC6uUE4JfWRaCMKQY7s6hWblJKYl4tozGubxi39
dIA1GxyRZXP6LP0OFpkmJbiTFDVVSWvtYPhjYK5KCdnAgGg9ATfj2p03XtFFXc+b
v0lDdEbTR0XwixT4IIKfwwjRW4UiqahXLS2POrm5t1ORcgdA5jFzcsytvuPL92X2
CPZ5BTBfHYZrLqV8czaYs1ovlAQhyVX8lqxkKUdbl3IlnAB5rlM52nPk11yQlF+2
rNF54k8/IY4tOmlFUd4JgpDoVCXr2uG6odMxNsfKJL5o746IHFjNV/Otymjrf7lZ
85hg4VoZooHpiPMfVw7Q6bWBE9qjPHqkmo5bkMYcFTSYHV2tL/ZBP3QKDZNnqsyf
q+qSFVieuQ2pky2mrTKB66I5Fy+sOnUyLLbvcej7v7IT7ZTgKsEMii5mEdtr7ewA
+kGno0e421aV5CLIrbS0zhL3DDUalhZcGQG7vOFVmkw4XAdwqFkfVGyRZLyp3pHc
uNJnDtEC5Cf7YfbzbFV1rarXdFXjBQSrPzZMK9vUMsfL/Vv+D7DrT2SNt/KXC/p6
KU337iwONJu69Rr3f3Udpxi17fhlYQ0AhniCApKi0FDFkrqodVcTHZj6Si7yJoCR
AY5aI+TeHOLboeAA5lbdYhnXZHPuQ4u8SX8gc+RPQ67CG6HyndL4FMsXc+96o4DR
1MR0YUfAbYUtN5PBJH6aGtm9pum83YaYt0ojCf5LsWRfGQGunipRt1qBXGurRVsX
w7ok7+ZXtRwWxMNGc6rcFiPalU51/ZXLdGIZbRWYWdN101FNsBcmkNbxLcTje27/
bG+PhPq75x8xGa6aY09M/QlyElB49NdMSS3rP8aO5lSche5027xzOu/hJ4IZT83z
Otme9+k+V6F15XIpnZcjPtxfG4/YDPw1lv/asSGwR59784orCVmMw/8CG/LnpphT
V41Hn5otzcOTi5nbg9X2IUmr/6YIpcet+60487pNX4XyLN+PLRAS1W3PwLE5KA+h
SUU0NS6FTwXARHN7mi31ds2LoVZtCKvoCxKr42zyppZA7VSfybtqFhLIAprMDOSu
5v6yvWXtN2gEA8+Ti0FdU/4IRJrm6umtyO1R74ZhZWvbm7yxEtCmmlDEo1juw2jg
zRH9UnzDxexQVlzYpmF/euEs3KVU2M5eay2557wx6XlT15xduFIlyGQ32g6iXs52
9QccFkGqyNnTYkupgGciyqXp8An+huyjdBu6RdimWlKVpOKoTfIvj1qP1yYXGyrb
pBhnwuXlbpBmvwG8mEb/rFimE1TpkgvoGUWR6Bvwsmiqg37fvDt8VKtXDXZwMz1e
RWZQ+P6cF8C7ZwD6zyPs76JHm5eKvzbHLydhPvo+LRS6hi/8eBpK3tiaxotqMkIt
+lp97x8cDSDtPmq+9N2BtVsYPP+5wYnz9eMs/b2ojy+r3A1zf+KrDx7VvLuM6sPi
RlBGtURsO83QLKgS84yl+2amVSeNRDqbJE7tiTTKNVTfXFcXitRSQzrOA2IcXhfA
yItdi23XyKY/2AIN/isEyT+0aIXSo3IUXoKRErtAFIN/dE5uvmaazM10Z0dHO0Zm
yf116rj6WLw/0Ckwel5ChEi3Vpsq6fIarb61D56uzOR9PIwKIiDwq1rYuW7dTV2o
iUwXtoW3a4ylgZswdnpQNwjhN7NYwv4uusKoQaSYhOKoY8oGFhWN/n3f0V0Tj5Vx
6nmjymzJTiqVZFKU+HDsy04lAFYWBOmwawUirpUV+AJZkLxX9qxgYijpbUq64Ftw
qasY4N1RJ7/4QqfZ2j5LZXTR5HBq+aiOl6bBepYUNhZInvvx1RVKUzxTemrlzuE8
BiD0IdpwfmCzG7TbIJhpTUqcr07J/lCYKCTmKy5m1RFXYJyfj+hYvxMyMhJb7EDd
C0Rqw9HwPHCqKDaDpwA3F3dwIU0/67cTVJzcI4vIP4SOZgM8K72XBvF1yEc2cAHS
qm387X/ArB0xFNUr9yQwU1cjHXC7U2B8rQbrMprQb0BFveUpsQ2lJe34lEkleLdd
t3ApyF9WgOha8lr0hTUy4sx33Yi8OEFEbAkQiCJvQ0JWbUcEj7PNGSq/owvcS/bK
5tlC2ofiZHJxJe4+ykZT3IAB00jJAQoMg+1660vYyu/dBvbS8Rnhe3Ru+3+N9ien
/2BtSlA3QXe0Jv6Hhzak/WU3XIKUTpCeulE+enwgRPkaKKO/NjJ3cDlGyzaOI8/p
i2NiN7XcCb7xkpMr2maD3ZmSPQqmlgYxkhU1auFdh4oHx6WYu3009WPxxJJeEGXg
tWGGGCQ3oBxyrC8UFHXYB0oXZG2MLEfnj24waG5NiA6mUFPiZ0JsmFubJ8gwbu/a
w9+GoMslZt888E+id/ezvpkZiUsUOgNF9h7BBo0YGbxJ1Xdt0ALy8NSLeQzjremT
GZZnsAjQgb42yG/og876RJBb5zb8fsKe4ewDb/AAOZbjP6rY9/Hog9GN8GCBAplh
79lFQVzu1lpsztTJjrtRViO7i/nD7DRN48Mc8HRuTPmtrkL5Nxx557eQf2KZDbNB
CwnULzX3iXjIjE8ZamE4Z0BqTTK9sbLM+HgS+UnKp5UI+nEO0ddNfoitVm0hgtxm
vPJYW7Jh7rpfxBeShVLXZjCos5iVRZZyh4JxHz/6VD5ZT/6Nh3cfJ0YanoVx27I8
sWIMXUe01stMIpCyom60aZhXVN3YR2SKbODVfHww4UAuaqJlzWBpWMtpst4ZQemb
pKo2ZaMY5K426JhoXU594gHsOrxazpo1Q7vx3B6Dgs1hMj9EGuNYsn+nk19snbmZ
Jlm6ZobUAB14Th1Zd+jEq+2BaAfwPN0TAOOZVjYJr4wJrCq/2x3EhoQp+y0BFz5S
EU5KICyvb2OXMDYmpptQZyxrxacXey+Tz6qbI9mVzV+aP9sBs64/ViYnk0e2BYui
EpDPvj9AOHgQWYVPj8uIa8+PxqlhnFgVFk2gILfeJ17bGSEq50ydDggflVDVOeIf
gy74rFisZtAGcyOiCWNblb25AzBu6KGr+7mYt/lI1vRZ37BMptGaPoHL7ggqA6EE
pKHJ6AQ4yohr7ik+TSNW/RMOVtErJvihVtX3opJjdHzUyyMBptKOCTXt/HZ3vTsr
eaJmO6QXjPPyGVmcmuDo7P8kkmaCG9nElNPvxlQdPdaCzzccfsd8iyyAZOR35XBU
sXV39V+gYu3H8qjkNjo6W7VEaXuXB03uxHwWcVP0KkM4GR5XXIABB1/sDGf8ziJv
LwTolnk3o7kb0Ssred6zdKJ3rD3Ad9aL8JfPKam/jr663GhKLGbLFtl3Rch0jq5o
Xem8oCuhtrv/M0K8N5cQpVHRzB0u5CTLpP0/kWoSaRU4SvBlmulcyDL0XVqm2xpw
iqX3LB5zABs6txes1XlvjxM+6QiM9nr2nKBzF2a2IRiIw2SUIpr43VVl1dYcsG2d
KhXOZxqFmGR9INUeSxp0inou0EMTKjCIbkt2iFqkJGVDYhFSqUG9GEw5FYhdfBfJ
o79SkBcs6Eo/i46CMWCokr5fGUzTgJnQkV865w1V/Vdkw+YoYLc41DGFvavyQz3G
vbj9GeBwYTgtAPpwbUmE5y9E0HMLTHvs0VNwK9TA4B7xUFuw5O0wwP1L3sIVgEAM
7cr05fdqWpY0crrX2OntkbwoK5u/G/Bd2uasBWav+P46sc+X5T5ZOxaZMK/74FCD
e9kS8342RyyvmoK6/TotfF3ZKQ0bL+QSK1dEZK7CxgM5Cv1FXRgfXEV+/YWPAfVX
q2muXYuDsntdLNQp3GwSjOKO5cWnFxk95VZnM8Z45Xjji8yK+pr1v8PZ7uqaQwYR
JxWrtgwhNG5t7AF2Air5nnX+d4grK9IX0tE44aXBiSGV80diVg/p2/Ul5t5XE2vq
HoqKzhLnixJvcvYw52BVjKTfrMqJx1g5OWUdz4/UHEQ6i3CZVNWyV6z5gfl+oCgv
kwCIOgs1Djn6QDPxYAZc1pAmgExO1rYn2quiAKTlJHVjiJxxCkeaE3c2EgWPkihp
F59M+XooanZ9e+nJFFnrMdUki2UNK3M7fwljJSPrlNsDF3sNyw8lQXuc828YQb2Y
KLbfWXDtNUT7sI1DbXbl2DzaQojM048FYlR7w9ki2yKSiWHMcqBErmjXkk/Sz1WI
zYEtTXUPmvC7iCZinjcnL31/PmWD12N6kXhgWC75zisux95/mAc7jGKBzJ9tQvZT
Uh4GnveMnj1/6la7uk8xySOflwNV0qyQPvMSvLxOU19Fs5f6/ZHGBgzBCmCuVxhp
B7doXiW6kAzvLju9dVpS4elB6S5QFMz8OrHDJT1uzat+Xl0o+mh1MW/iN+tCZs7m
sThw0SEd0k9x9NS4SiU27V5PgapDaW+x9bSBsbpPIUGaZAeonYTc3yU54EQyQZ9K
/uFhLUpKd27spE7JQhq+cjbU57WBZv0lOmRlt2HU0kNaSak3sxux+XWWNZgK3R/3
GkUcqi4cyGwK0Dol0Kwbea88MErdPmhTyZoY8tzgj4r10nHvkeuRWfGwJrJuzVxc
UZ/fDdcvw31y/Jk5hBi3QeJrNZ/6R2sug/ZeDY0PNlRUcceS3/Dmwpd9TT3V6xGc
I7nZXsTOfiNpbY1MLrbuJ9w7GC5J/blkSuTgj4Ofr6npky4Otf+1kVFWg+fry0kg
g9/9pMJlBrdo3EoADCoPQrXx3SlYcS+lr2ScHV/RnKFDOxCE0AQlXaXHZPtUHfgv
CyeWFOOPHHroGUowp5uRwQn9uwuu6zl4khlIV9i9PmQaHZ5GljmC+TPtDBi9rRsT
xx7wdGbFadbCWLq24oFCMwCIHcQx0ze6ZZGbRe+yrDff5iJAdZikGC69IZSWeI55
y+HZBBzmqVRAzaXeg206XSuZShEk1kA36IpkDkoNIB3rURN4vYlA1AtaGNsQa2ik
bPpFFN5F+4wsAEr28DyWyCCb2vgG7K5WEIGFR5NaTAkD+FwIziGTgK4pQNUQGCJ/
cLuJ60wbxB4Lfe1fcflwQq+V/cgBvn0jORWQrCsVkrtKNL4hlwzDQeNYXOM7z+iO
S9Lqh262WthigSwUUsEc94dGuYfpuWFDRI5ntQhkHh3rb+IyiWzbXBwaoX9kCFFq
lSMw+DYPNvSSM/+nFaGxCfCiRfHaOTj2FS2U15N7AQoUtfquDFhoN1+H0WINHRcx
3Il9ram+peeLDGqlAzrDuua1oHUgYz8MS48/yMdEvNTDtIByd1SIdlHUuGXyfuae
dyyEBljlb80WW6prMg8W8+g9hJdz0Jl3XAdb/DA0USqPblbZkBmGF/j0t52LD9hV
1E+2J6QSbp0Dgk8PtrupO+/2Mx/rApORPZS0cEapN5suKw14MVB14GPeUuaDmSkq
EU4siC94pWyqSqrE8Q1vEK9UJUPGkQ+EuUOgGyBzfppPJ44TszBs6K8jnPz6eEOk
apw29SSxSmpgA3J5BmHKJjO/D2Iz/99vRxU/65WBQ7Fq/GzCo6p0VDqmlfcBh4RL
ruz7YxyX6gBo9H8Ys7ac8soMGCAPHu9F803e7QxH9gAiuRkjleykxJmR9mDx/CsM
xXdhYiZlVyq7CKdqQh/ut3EcCEvyZbTICmGnJWz3G11p0opK+iV2l2JMuIsNscmf
7W3j/Rw6XdsQOYxb9uls9PF9JRJrGbqkgyviFCwkPDWpQ9G/XfbIaGOmL9wqqLky
x5LUBAcUmyl2xfQQQue5RIrseNH43utA4WWpOxbpOHWBOCM5HOkjgs8ldkWyxvSg
+/4QH5Sce5cOHHqs+dHBaVK4fHL9ee112c30vam45QovqXNi0BTfGf3WFMkXYIeL
bMydNQsLNX7OxRXdqs2DGlAiw/LQYD/u+FBU51v6qEEYlqYuQH2r7v7yDO27J3xQ
BKGvnXXpJZrd9ctu27XhNLuyJB6m7ShMxJSJ7AMTpbVTn9O/vAq5grhJZEtQYC4T
yyFeStNDgbMJ68OC+QvJubXiODMSsrG+wwoo2fDY/KRM/tIcOV+b9c7hKAOlzwjS
k3XH9buHGBgPPX38yB0tkHiy2fNfHvxmN7m2qKidWiP1vhjKyNSCB869g/PQPpEq
SVIhBWkfGA7y9fICNwDJCFfwZe56KfVBYLHLGmKLurm8gkZRAW3mzpxMW7X9hrjw
Vp3NiqIx1ieNjLIwA7bK56QotjvnZWXifjNdbLoh0vvjPQeMgqPRMMi+mETSwBWZ
qOz0yBgnDQZNlsBy1cvLUOXUrlhg14OExNsUSwPwuL8tHol4QVtRL48yV3pq/mov
P7bkrOvoK5mZ35FS0uZ7H6GGvNltL8rH3bsv1nulY+4o3hhgX/yA5iwD0EbdJVH8
6rde9jEfl4lPnofyqnxWSNafpSEKLYF52fWVFVKLyFBvrskCnPodcPG41zwaFMzf
Un+qbsbk4RzSNa/dmvWBtukqZr2oaGnCjt08dr6MUqi/BJ74qn4mkGQGXrdtxnFK
BLC8ecPZ7MMQNDHsJQ3P8VwkdQjJzHLLAm3Y4J+ycxnRvCInlSfGtoPEk/cRlSH2
XTKIpRg2ary9ES6bFmZE2ssVsloqz/tnV36gzJayAGY7aJazmHgiKWUEy1OOmvzZ
K5EtxXMQagb/0HASnhYEniu+exSVwtMQGXTFLXS13mfMcI04z2xbNj8sEA8ImHp+
XcOD/u/tJ1SW6j7YAL1yOp9nQBTIFobAutmsCatASBnC0b24cNa+aSFMb0Ekbm5g
l+GbzU5iVICkFc9woFMcogSYtkvA+n6Bit6CXx3HSEZoDuHbsSVqORY5T/IMxf4a
Aadb28CYGandvpK44ROZdyrRjRwphx/098TsUq+1wQgH52xpAY4wB51fXstJj7Kg
m+mzNr6qzCi7IQVU9MzVMcqmb/Q4K4lEitXvgZqg9kOHm9lEad30035LPDpIsaDu
zCzcEhyOpk5qeS9OB1+A3U6ADdtX81sNxTfe/fOFoIaNAL0xTgBy2qNNQSq+vPTW
IB/Dk8khG4ee6FoUaqQ06DfhgeeEXcjr0BUWPX/g4IkC5eUzNGgDMu98KgZh8jzX
5NnQnbpRtA9EQZV1Q5kc6BqYJ8CHHI2nlD1s+A1zxoqgJNtI5k2VyIKAVvmJMdOu
AegryQDtiXsEU7bWOuJFXMp3UIMfGzE4c3faZXZD5a43tmwk3ShpKeCfHzaxZeTV
O8b4m1IRVQNMdwcQJ658XD2bswdZr85IvkfEUOh7BmQ9rIzsa0VwDE75fn+cxWZ2
HfZuQqgnkMr/O3f7QroVhybracm/90WuCWKf1GA9Ebyl+q05xaX0Io3bitiUJrbX
N3Y1NKMDCz8gSHIH4g/yD9dCmmTNMRDFPjX3NkOazYVnJFoxSHenUT9oQFEu0XZV
1ErCIx93WnGCWZWGPawvaN98pZOSQ2A8UYzmtkBSIZwCvL6C6CAAJSyeO9sAGeR2
MwOWTD8z27+TffhzQQBHCezgwGhdCi9hBwbkXJHc5N0KWRyTG0obEad4FuNN9ipX
RwH2xF0zDhn9iz2leA8BZVxUIcLEdbFboqIEr0cjKlld08Ed7ZfbMB5+nyvGkSdt
rAHYpWm2lsZQRso58JY1bw7lsc3nUJWx9cQZAj8a29de/JPpfJHh5vi4UCft5ihU
l95rEf2svb7Y+qv/06BPKOhzBjLdvQb95bUDJRN7cwpVARZtfMH3hJaG6O/J9ywW
IVVSVr0gZzz+ffwjwWCJRFQlnDIAlvDfnkBtj7lPINYjukgniw0Z4lPnV9S3SKSK
MZemEUT9EnwHiR21WAsQHohf4T+64PPmmZwyTzxyPpxJ0nsQIduM0wSVfBMEgowh
u3YTAwaejGt1F3rKgSV1hsKOShDDRg8YVeI+LCPe1FmPOTfILa3rg3CiXW3+p+BD
mwsbWmasKu3qhatlFtpniVzuu4sory+3xnWd7mm4nLOiDnwK0csyFKVnPLFvX/5t
UlF4icOS12GL0jVbT97+AWXvLSAI46xftXnupy7/tf8M8xWfX1lbEoGXYNyH910f
kF0kY2eirIY0KmdhrZ2ke8wMptPMsLIq/xe6TKZeogpQD138U6pREJ400x/U/vPv
eGbR36OgN/XcWqhIalRQB0etnMUsYbFPYoYIXwqMyDHTzP5dcpAtOBLQ+Ow1cdht
Cbwq4Zdg2kyWy54/ylHAk9kYdUkvbretc8QRapczBYNaho+T4FuW7W6sOuta1ctB
QxiUmxchc2lOamP4C8aqHqk4SFEkE835n4DEX6OXUgY/lWfnTcJA0xniCaZnunJ7
nE4JvPMhNQMc66a2QkXn4a5k6kLnNdNzLbUbu6ZfJME+1L/Zen7zpk7kUxw4Zp/X
UIXF0Pbp+o0CBDnmHFBIzW/hv9uWb7+jA0XJ72Lkqjk/zrNN+1r8ubmWZEQ1OvNI
Yw2OVulIWJ3j35CQHEv7/mCMF8IxYn4Vfs9v+Wwum4ixVbu8ZpJ4doIZfAWEwH0S
926bfnljKGZLGZ2pxdPqRY4XOMMXlnGqSRwB2ZmcPl4GGNRbfP+6xqMYvgBfv2eC
4ZWNQtXEWI1FvxSz2qbaYS0SocBolZnEJpRtC8FKO90dqWKBcqErlAF6SPvD5WSh
oeYve/sSqSFvh1t7GHALptplJa0i4T40Ds7GzqGzjTrjcSP7x/Mkkik8NTCkinb7
y1ecJWrwozHrJfSk6hdZEJ7pRmHlbA5SwI/LsIjzlIx6ff7c4JNbRbpqUpEaV1Ir
r6094wt5tH+Z75UK0v9lgIXAoM0ygfQXzjnjS0IuM1cRhIq00Iuchoq384/njN2K
rPfyaFyVQcWKR5GvRyJlAjoIeqDdd2+7GOFOOiAgcuLTUyrki+ZLW+QOOeLboZLy
HLvJA3TEaIWMVqSFGXHRcSbt+k4N54kEQDUvZZ7q8Xo8xyHy2PrCLySwoolpKIjX
ecHWcbhUumlGsGHHFhoOMnrKfC7yDWf8HzWDZqEqWRzFKqGYSCqyYUPfEQIf6Ab0
LI3niino6vvkAsYBtk5Jz4stKqwXOQq9FeFZ35CqRew9m/JfaXfJNPzqqr0OEZ+s
53MoyV7GVJynUdcHBMyiJwYoYD1XVPS9QLp7B3fuLFlqXGoQC/Yl78toGj8rBi+X
8XckfhKpdQByLWcngflOYdPb9NdJjtzelHSPFRF1YnvIMiqrXtpyOXbDleRbrKOp
1y5osajBEklczwgyBE7admVO2Wqv5RgFY73lsqUvd0Nh/1RNRz3xAnNoHN583dnM
zSgb37AsfoOGl0wPZ+x4L5BnyyOHCwdvPi/xClr/ZxZGhfJSrf1NHIfmqLz5M3SH
MDGl71MYnuaUKpUrAIYsOOhqxQ+dNfOuBhSjC1FtTsr5fZT8CUJ4JynL9fm5xT9Q
lmbO+rfBGJqUPgtLky2kxT8TFS1Pv11ZYmp531Hc1jH8/1oMJTCu6mLl7cRdkTrI
f5kdrgUPMZokhXSkogg6rqz/6GVnsfXROuUlrQavymt2+diJWiRHP8Jcq4L3QGEG
hnR2Bz13j43knhHe6S7+YoqNyETNBNXvKzLew+ea7RyC6H3YsdUCmRA7euTqoAGn
DIA5Ag0CmX4CBF81Y/Kst+So1DzSbe8rYCxMqr/szfgLy2S718KX5kNlB6ru7JGr
en2sw7tbL1Q5Rit34YAf6Pnf0OzXJHU1atFoy/m6d2No22CACDfIyA3XdKPtXPlw
l+ZMqDM3D3vhXmtUA/W80Q98dtiTjlOjOWKbE7adPJbfkxl+0QfnKxwARVTX08C8
ZbBl9AK0pvnSYyM6mCwD3AjaLj3vN5k1PENfWyDQcKErueGa/SKyKxTHptaIx827
8CvY27F1dqevlbXyaro3Jx6pG/COUPnPcklpL3WET5BsgxsQu97yiIXKLOZCBtIa
FjhsVmIEO/nb6+nz6RjfWPGJ7tRRaY6+p/NJhejfWXxh8oYXgemLg42Ox1uC//ae
OTFajDw4ZVsfl9kede1cCJWxZRd/CZqw7MAXuWPiVqldDRHAEHdedufnUsZ043gY
XZhmvXnyVLPUyEpqQ/qYoP4M9qM+RNO6OtvGriXQCSNUX0zWDvKEarpeaULdM6mn
AK3dhsCEYqOKRkxOqA4TCDOhrUQim4nlT0ScjYd3quVsHTVJ7H0f1JqNHUXt+23D
ffRfyhnoMHFfeo12dIpLh8a66O+0Hec6HPVivmW2l29TIG0SnuzZ7G7fVdobftzd
7nRLPxVPEFG2rsMaozfA0B+ewoN9rCny2LlOAgV07cGJuLm673357KpklsmyAm5N
98UDUvmY7aRk5LxgSJ2JiO/D5RZbN/nu4zRkAZ19RamXxvqDaf5IK4Gck4/rHhRP
1+OtgCUAjC9iVXz/Qf67D9QqmYXGWqd/cSCKK3DQV3g824oW2DNIPZwZxb1eRGSb
PgFvlF2H4hhj1Ohtd/lAlWeo+dNDCuT3RB+2fDbukDrngl4FcpsGzio3E2znkRkn
p6N8SMdbMw+VOtw7zXjKuTsqJhHJfeXJjEYTmCG17n8YFzu0HJ6HHZKLAbPxRFc0
PqLNlSvEEdJBoGqU5v6X212H8gIvasnBYm1+RjiAfQicjgPsVFcOLUuv5SwX0Q4Z
vpeSEsZbR8kK2z9wtKoggimWH9CEtpiqHu5oFGDjVRFNG7F1z/mod/zqYTcG0ROE
Xk/evyCZWbfAdRCDY4XT9updqxaEgvB8LAV0Pq71vdujX0xWntjQj1aN7tH3K8VG
Ijy6YeJh7YsYsc4s5EvooeTzw37sNFu4cQeMMnhMgkyJr4xCuvccxXRSGybEDgQA
8L+FY7z9WWhTfNgw3ezS+LJp6iuh7IIlVJRoZ82K4qy95FdkHoiyRopEMlI32Ji+
YiyOywcEg6+vpX6yNV4bh3XSOyDgK75DbmvL2Oy9Z7g2ExbEqvUcpj7z192Mt4yx
VRcGbS8PQMGZ56quX3V32anFZ8141dwJod5FNWBKZJ1CxpEO0OSdms/RVJPu7vog
Juj1NnnkUiHcmLtv085/LoenRJ4KNcmftMEscG633/RIKtX2L3PbWvKMZ4avbO0t
UwuuqbA4jvVciVhKsbokMKntjKdXRUexoRwq5fF32zT4LKcHr+UFKqx60OHh6cP+
bvm5LtvDt/cW28XJaByrAxV2NKUXRFSgb8NcmzslS+8JMktCkCx9uTBV/39gKhwZ
5WyUEAx+hsTQ8TXL43yi6nMy7oVg1nQ2yGcm6xnW623TJzLbZ2Bfr5BLrfxV45DY
kId2Td9S4rN/aU3CiRRb1zlbfwjKErzb9XruNK9ZMyGf0x+3y1jUqZK6Sk828O+r
yxxKZw8Tt8QeWLvgPEgzEiqr15Ep2GcT/2Y+4Baam07zdLmr2eAhUq7x6ygQumbl
HiaqlPt2DV0Lfe9Ojjf7vISndb8jVf8o7qOCGP9OdVdhV0FU+Rg4IfX1/9+InKkx
XKT7CTKXDvdFJWDYUwhKw91ODvpAs7KBa7nMIIu6u2aTUT5cBMWBubPspQG8s0aN
erwaLrAZHMqJr+z4vNZX7XK6/eB10m7ti5gzNcTmOcBeoiWfHt2jt9H8hWCnYjRo
8+TQJU2aXyXI6g9ZNpkZPLiSUuiuN650Szp2OyZEdFpqu7sF4SFbRlUJMAgTcxie
pG/KkP+aRq1+gA5PBf2bTvzNFl6teFl0chgVhAbypuP5dUcU0SdbXaADw95s4kEf
o/n8wcKJYqFtRpibEfb9sLE7kd6HabtqGqCc/+fCcDYzpZQfQncqLe0/CuS6ftn9
JZieN4EIh3cg9Gflpmc/XCKxiQoyLKsY6soRBmBGJQ+bGzOorSz6I0Mjh/gN9/kq
cMwl+9ZdcoLqJwVHS2ggUpZZOfEbz4o/KGoYrlJ6jHRjw+iWFUTlOR8rzglP7Nah
XI4iRq+3SGm8tkc82pFgSKZA9wSze2mPdXlzoPzKdrj6bXec/MWGibtnEKIkaJDU
fi1Gpj2p750KzN7xAlVcnx6vML/rFqv8Kg1DrR8iwaD9Qdbf/09KGO6ZccB0Txur
SUk3PjozHNHBrh83i5K48F7deT1lRVAKcMKPsCWCoLckkCTqgwBsbhEVZamsieOI
V3Y+65NokHp9Lyqc6fLJhRuiWpRnrSTNzSJvLqWJm46afQj40fCRPn4EPmc6PFcu
jYGhzhc2g8BL+k9xy2lUayD0w4eMBmGDBKc77tvrXjsVXEYtddDtLlIRfPxhQblx
jJsIohIn0jVGE70KOHs4eAhyCC2Lg4fgeawXC+rrxiwyHGnu5u+7CNWk9AVQXplN
rdRf7rdR9nNAzqwZbCpxq5svUOOEDGXuv4IL6HeCqjAV5ivOHH02Z1KeIFhWcEma
kIVjY5iR/q0j06c7tKHfOAgiijmjim+uqnelsTSv3cA7jNxc814BDl5BRGI6C41j
x2n3CevymcrJIf2HMo83xK/n8+pMWNEr354UCl6Xes87/AwqMs7L/BFow0T3d+XP
TLrU4Ny00IIb79OxNqweicE4CajBAbEOj8nXLC+QArLvN8It+Y9aRjq3fDtUsh/X
zZPMTlX0hDgnLi06GoQDflLfTUxZAwDCbIRP11vA3mYhwfCUPpEHDofWQgb6ObZg
tKzPkMZepPnqXs/5gralrPIWEd45tj2cibJiOuRv5uR8QQ1SJ9oTGCx4L13sJtqz
ARFYQIoCIr4F9rKeZRsBkVI/el9WzITPzWVSnBfl92eEMae7JkBr8uKiuN/nY+6S
qmInRTSPDOTamCizV/yI/9JDFc5GUiVMQhrgnFcEuVDpBQ9dPly0yEyh/oxJ+y7C
zi17TdDF6kQYqwog6CZccLtjWRNHjhDQi0O4ESsASm+I3MU4y/O2HT8yn3S0Z4+W
STJVultZu8Wqlywya6LdHJSC63KKnonlR+jskSi+95hjjbIVc9zV8fIR7Oz3ttpj
AP6eWTTt/1T6S9S3NYMYJDxouPvZgTSSHOJaBCK/3/I3ARTaEOcdjlTYDMoV+m2g
bQmVxT8+QnOvFAlU3eoxjsF9gEuR28AeGEe9m7SC3Zg1Ea0ADH9MiP3RrMBL8bTY
kLDwnT2wGwpj8WLeP3931sQvizvkACNT9KikEi1dvB6VW8/YZ/kiTrw/zeHPRosN
cbO1jp44lJntaY06JsTP83M/oGhELXBz3DPiKIYDHypF5iKc7OnPt4JLoA1LrSYw
6+dp/WsfEzUqsHsVwBuCxgKU9fdLJa5TdO1Mkmy+BAR2d8dqIMBqAUCrsNXD/BBg
q+oqvAI/ohBcEZV25eVFn6E5mDCpTVlaSOm1a9egzZKyoe5sCU4ccB9hh5k5WXIS
dJk5nn3aox1igQoJzukch1jRS8WqjhWcg7KsxAeYcoN62kqSC/OjnFMdomSW4iKW
9+l5Vwzow5zdGGoXd7VJNo+Z5PBK2l5ClPSntEu3Yh/gfbsJs+8J8/QF6SDx5n8t
/SVgvZbVi9ZkMuWmBaTDVllxqg113hKbeE5ArHGH7ycZpRSnr8QWjU8EpDySYfqi
C1QE49xUAsbquNnMBr4q+al/eMLAKjJp/0dS8QD9k5S9BvT4dAO1DAnVwbGAv6eh
KisF/mfgTaY+TzF8TUpEz+0WfNZuS1TIlAz41Vt0teLLAG2u85h1y9YnxnSgVjDl
7u4JxaX45Tdt4xZF/pPmD16IJf3/cq3uIGlcXVMLp8bV3BrLGogFtdONvQHECzTj
a7wiaXcZrr2qEEPCKLNPu2EdhtGxyLH+mcd9R8+MSvH4YkaRBlwVxShLX4SJe+US
A/VFRgP5uaEJz7E7VXUx1lAoklw/H1e1C0Qxd9eV5CLezyCBHCRRXeJdd1ROFUqt
AL4BjwxHayD4Q1yIXtTP8HOL4j738J161gjmeuk3srn4dZTVX8lpO5mJsYrV3Klo
Xqittos21eRyazp1bfDWZwc9682Y+VHLqC4QomO5H9KBllAcN7hyCcV+ycydo+tV
uJopv+1rUkhBCCEUAS88ZtNNNNxOyimVCIk4OIjFqWGk/uatOfB+2LCqekZ6lfOI
SgjMq9a5AyVO0aAiwAsiOVHioetSeZTWkTC7MxRRJuGdfQK0yz0nT53rOQu8xlUG
7MANIz+EPJKBrfUlMdXk7xWMTNKMryIjzn0WhAF7W6GOEKtkZ7loTh9wIr8beRLn
bvdQ++UGdvUH4xTYzBBDSZNIEwUN1qx/syIcPpkn9jyaxzR9nCNV6IDrwqXSezV5
oihcIOSArHlLC2RD6n273MqqS5ZX2z59aLvMT7AScIAqa/VeVsDUvuG+KXi8wkLj
H9bSZ0ZIkaG2Gbk/7vPalIroe9/cA1TP9ECVnVYUuH0bc2w2JVsCjBww/pLHFAaL
t9X8mPErVW0bbbDPQYn3fuUYRaGXl2EM1s68qeuyt/PDgNXQVi2H9Bcsg/j2Wk/k
m4RCwUTwGz0Md7cYnVdpWAkelt3DK1pP2WNgGuM702/qMpJGYhgSBG/H6ZOdqhEx
rKHJG/drXwmnk5paC6wFpZxuqLf1LYCihdDMgpLzu+HYoZQUXUAToYAl14f2P0Od
lqmSzYEwzh8v3jiFHZgjzxSBccvbuOAPBZUm4G1oEU9aTMsdFha6utiFsuqEVLVM
ZAntRZir4fMil3BbQj0gaG0BpbRtJAb+JDE3+KDRc8famcUiV1H2zPJbIlJhgfyH
Jfm7qxCHm1KDa0wGLlRnriCs2XIGnZmj/LcYd/qKIpVOrw+uNJKLf5mWAmd+sZ70
qeGe5jhCI3HsE9VqD9s/q7cHjEdZCOel3VV9ZWdEphLX6CY9EieQJxKPJ8vy9sEx
KvzggiegaOekS+Zc4gStYRm0AAtqf69BkImybHXNIpc7RAkjrmcTZUsxs3iO+pH9
ur2/gBgJJmwRj07fFIulc9S74ET/xl7GZlUyhf7nfLnC65hq9O8+o9RQEfuORJL+
cc8FhlNbn/GOi0kGXWSA7i1nk3stL3v1O2BuAoby7XfaC13Z+s/KIbW3BN8XWuqz
3gNL7klnI6IzsNMOVxDzYjwaTOehJbhk0P0gFo48K+5K6lhenu2F06EwyhfwEOIs
fTVUfKivcpB8xxzzgjJgj9sEcj6J1HaD6GTkiEVzAmYGxxeBDQ7gZSYqUoEQhvyE
C1grmWeQQvpisyEIVMn5UGLTi3k6fMprVGHqS/LNt7hicteSpbQRoVWIJ0AvUSWS
KM36qmVkMV6BHpsinU/30asIHsiJu5k7a6sRNjuFv+/AoagfbyR9Lr9vxlJn4WSh
4IUmWJC/UaQHsepqtbJlDLYomr75Pib5Lc/3fUpbPelvlafuxfVptMeD8N7E1PTP
3eOJGvkwCX2E+TaxydDWdgZSpN6aJalgzC2ZxuLOZiRf1PmhwOUpqbfZj6h2nUqc
PFCYQiaKjK9EL9m6jGVf+R0fRDqNlV6/OJRlRgblR5MwA+EGZX885e5LOxNTaLFQ
tZlbs/CVQ70rFiDQnB4SFi6XXO3avV824CWjzegcu5WD2abkDOr++hUXfFmpNt9I
QHH7JOPVk3RXm8qKZ1yYypHwcDqC+lVRSUNn4ZEKGIpJcpgi7C6HSBSediQww9l8
t9y50CW5MbtTJIV7dURTso7O/PXfOuJ1r5YVCZU2gIZJJBJLgUHx5JvhVTtGgIbl
Y47nRkhVwVNnkTdqouSsMcYRbU2gPQomxs6S+JmjOCQ43oGhwjw0+BQttf42WdBR
jzvFmaoB4aGIotwUm6QQy2bZ0gNetmiyRDDnZlc67fFmDgCJSd2qWgfZQtIwK4O0
CBLfFy5+ydyXBJflSfd8MiiJSqvzfw58DSmQKIHpIFlbCZuXUun7IfECOpoKpmV2
jRWqVUSxe6nSUHm6bUPaOBjcQHLwhZt9mVl5k2OJfJ3PZwSTWf/feY2eyYtYJZGf
jpGKjLlidF2OGrxJNPuDPqp7aKPJGgi4DVGNkRpKjhsCJNA4iTCKU+ScSomEx9jU
XhO4dSNe2OCyhJxrwEY1fiRi/d2hXsm2nkKdoNmKZeCZptflM4dgU7NVwk7W6LzZ
OyGPmIGo69uLS0cBflz+q3oNliUQKtEhjxyuJ2So+lCWu3jPntG3QgrXEjbasDgz
Ke6WO+DHX2s7wNSENCcsGjgWD9ipOEWewQ2bXsU6cVk85yj4d7jaCOIBOYHwl6b1
awUBCXXwxR11TI0G6go9ThbmsKS6ojT51ytdxoZs4fx3+/Ibvovb1zGzOTT/FW56
bdw2uZ4RWDd/6fxMMN8ki6GC3WGXPCzDCQ0I643npGjvEncUqzCb3d2UvdLhYPK+
oDW92vrj003sq6I068BzdhA19BalizMKGJ9rZdleBIpeIIZRD5hRGEzqHE8rlTyZ
k5ZC3C9gK9xd2ekMdhklKMmLpT7VFR873r3jfDp3XR5NJQKeGAGbfcKv/ocAAlvg
GS3q0CCUPQdxiDteZhWV/I/jQ4w4W88UyHbgFmPTrC205o/wzIhaMVEnVpsE3Lk6
JinoROKeGc29bvmROc6aU7tCTDeEEvd61HyndKewHdu5NjBu9nBnDmfh3MwzX/Op
Lo63JBeCaIWrv6fGWJRfdjMtdlPlNUCehSbXNY1rM8bK2mVHEAHKaRPiHgkJxtAS
t7UGC4XA+IsoWqSGzDtv6/Ub3ESRLTaZoJ3uf48cgdt6YBNjpgKgGuElKZ3fB/dw
tKjy/1eBxCTlksXVhXBQgC7SIxRFCgS02a5fm9l0FXBT5RhZPQSsPD48ZjXsHx55
zX53sjzDtZu0mV9v7/OHRKAdt7ThlwbAALBO79WTI96thFd4u43X9sYOy+ljdJ8H
wJJHavqqL24Hz0DDOUiIgXoXI+vlmEJ6s2I2WsNmGWrRc4cExHzHWgGFdP6y2cBp
HXkl8L47rqsHI6AND2YxjYBKCvNBD7Nw5k/zV7Y1uhuFgm5XVmoXbnViL2z4PjGx
iiKsAcpPiWAw4/ohv2Hs7ypIQwTqrNEo7t6pOOa3z+yHhnoKWL5Sz4eHXqt5l80Z
u2m6hpfaJJ02oM7w4svPkodGLAzKy6l9qDKz+jEZZMjJSfZDyqFtG7aNI8oeFJaR
HIHF1PIp2QCjTV2Jk73gAYOvtJcbr3EkKeTf9VIaBVOSOJTnbNcGrzFhkBVpA36V
g9BsTqoR1SEgA3tCRoA6NbzD5KyTMlJcMOkdJN33OPi4+JLNQJWJ6TBeWH/BLPxP
D/cONNXlQGppBd0RU426auSgqo5S2qbyRsKRPF2EhP0XSoW6l+/8hGVzV+DTQyor
se03iRz4e7HeXp31Q1re0pGZ8P0koRIA5RUTyUmkimeFB5W/cBmVOi6OFuj9kzuj
hkH9ypLJd+AEamwz8iXwGAjVGK0B7z84HovfaxvjruA9ydEUb6qc5cqgdVEEdsi8
ZvwezIxk9ERKXKb82ZiG/ZCzYKaJbwcTxislbvFA2W1UiyYH3u5kbkudAIL3PnSQ
9juem/N92kz6IdYqUIavCbhE5azTJ3F01z/Nl1Kmn3wA6boLGa4uuZHXTKIn7eIn
FLKxqEBCkG3cFNfMpEbm3VcInpUzgKzbfpwlcn8MEykztBkqQwn+UmZMbHckWseF
2eRv0kXZLeEuHhKzmGE0GGpf4dPA3pqGtHpp7IS92NfL7ZNKQB8miLv0TkpxuLxJ
FnQHmGxBfpw251S9RZLGDHWk/CEDbZZL77pDupHU2RjpyxGbrPeM6fIX8H+2fCJe
kzWAgoA4cyUVcZF+9ceemU+M1Tyj+adzUV8cojPu2P8ZT2EX0fvhI10S49Z/W0s6
4S0obmVT+io06J+pBnAeAa7vTkOdAx+jB+Vyfhl1DbnA1I47md8sd0jABqyC5qye
Ph5w3GeN1+S1l6LMx/IgHWEydMFA7e8nZ2ScAfh13nbhaHoR9MixXUml7XMgKhSs
rHXw7kcyuUtNNGlft35f0rjU8zkLpQGqSjPdwY/uwoqhHsyV2r4jV7hAZ/YZj6/f
iDkRQBG1C3m4iSuAFLto6WPZgHdtnZ1FSSD8C4y3WASOUws2bD1Bgw8+iTqqzr5M
zxh5Kpm4U6JBKaFNM562y7bjaclr1m0jEwki9oehqWPDXZxSZkrwnjIYDFsn9eo+
hcvQWSilIKJudiD79saOJX172dwQO7p8KHtSHQurZGPU1+vDt/MQyc7QGoGpZyY/
kiKUfzxT/YQTtzILZg266hkebjTa17uOFhxEE05mE0286FpjJb7ojpD10ZKeEiij
h6JToC905J0yLkaSEQaeVwIx3bg0AMAUbiT6Uw6DjBFxWXIalIUkwWbhWCLNqPSN
CPEM8IpTZOi1N1nASBwm2TrTYqCCPmsDLl0N4CcO+sbr/id1WZkyRiPiVM58nbtp
P5UWhBX1Htw6H1bMpMHo27oAONrhvLGOJu+ylhOXqZKNEeyJrjAGFgeAle3dwESo
k6sTeMAp8ewYgClMRIQAgQ6bAk+55knQbvBPuJ43I7ZSYetCbv+OfJOv8OCH96fa
m+0GsXvauRwEBfPt6IPKHYf8lQ83cVEUCVmp4XrYmsIJcdutLVy6vqKiE/7hA7/G
Q59odDWVp5c7jF6dBMJZ9+4I6KnlGzogoBSqRI+g6TTQt8Kr8YormHYaPtWUYAsv
2ithPXO3CXmZpLLUM3cJGbZUf3AgK8aO4jbWnw1poUUjz1Ms5jgYd2Rl13HeteEm
DD3CnlqxAT1EBtCjQB95nGuEPh5p9BAKefOqmyIHehf2ru61WTIxWzYp5p30XQY1
lwuYphoMNWSQduocJsitYA6VSDL85hT/iklkE7fH5RJ3OCd2UBWE+DZXAHlpMHPt
yAkxAEWdKzkgb1FnPn7/H1JnAK4dt8FumQL1ORGCV8mowQQ2Xa0AMUMrqQtuwkK5
wvsrxiHub+TSPskN+M0nlP1hS/eKsDFQkhOZutHkuvyOEZg9FzCm9U/9hl43+8PS
x45M2h7uJ9C+oYfZN4OFFSX92bzA/jG3dIb+t8LqV+HFiwGdiWA7xJ0Gi9q/+ADo
H842gT5cL7jyZCdL9IlvVXIqGldSZWSQgbeDa1kW7SIMtA01VPlpfpRiiBvI9rPm
wMiVqYOE8QTTfE7uEOMrwfsGTe5eMX+kaajLL4XGSn9kw5vnntHSOudccd0AT5w6
RxVDxyl0M6uAWtuvNOFVhzJf5Pjl+n6w5iTFMBtEG89JAQWZN7WTBXJOE4O5z3ij
kOqKqwkcskclZMDDYFFohjjHp1hzUAFiRsALL5fvurvlHgp73y16IKYN7IdTSZkP
6BsWl6SAxsom0LD+uOqsfGHjCZgwxQIj3zK5UOrGwhH3kShZ+IXDzzeEOQrU1+iJ
0lplqG9SHfVmcvdu+egQXhC2fypvC7tvnFoxwmkzib9akwNSXC2hYwkUY8rm28Qo
RQ8jIop9sUGNELyOsxJ+9bPrrqqBluDhb+8pH5E8Xe9TfEbuLdOvZX/DPSHeUiPk
a+y7W4e4j5B4BtPLZD6op2a4eInQ5QJnc47q7GTRmO4mlbTuymU8qUTLQP+I/RA9
e3MGRWW72jJUO6+ktUFzpEYMdL4P4MKF9+aliBNxfCEqFeZGncBfF3CpXWw8s6qw
TyLinKT4L5DXRIYE708OiggYIfcBC3wgTTEpXry8lox6yg9fHqwWI904cqG1obp2
USlzymcovpxf8kF+ueQZvJ2cTIlyfj+5x0Efk267UV9idZ6u7dXniHEda8pSCBS6
qEZLzfs+YaDYMYP5yRi+rieidXa6BxQgyjmS1wZyuMEgZ0NgcktXvHdvxO7KnIZY
z7DrKG/1lttzpW8EHXl0zi9Z3/vJ9BrvGDpGQojl2RabKP5vPUML8Po+mTCZUp1t
hVIIz73J++R/5SBeT6moHQsqz7GARXhzutD0aq+DBtAykLRkD/J7PXQ8a3lKT5O5
kwcC0oOxYKh/rhcbEbXPUeupFsKpv4qdECIXZuxe5UlhnY6M08ZOqWlk4Iv6mfrd
oYx7dIWNBIZ3wpFSdhiQooKf5FcNHKMI3DFUUWg5hXsCr0lP07S7vLPBhMsjI5eZ
wbeh2+gApfRYC9rZvjArbnPq1CK+v9N/RagDmb/7eq9eD3VXrtpepKnZGhwiEE6l
d6C9xGlOKsexroxKj27yGEg1etbWFYYrDQGsSGAhrIzYnFO4Pbsq/cV9dkc3EOyv
aL5dSOceoIHydTFt8qy2qLr2jlDZBix5REzddN8TU4J6j919yUKh4W3GJYPJoo1m
2a955L6WkpQNf+7hJE1ARMoySOPpAwygjOgcxCqltoJ0+gq6QUuvFZX/LDR8tdOR
12NrNW3xH/0kz0Z2F3nIGwK2NQahoLYG5Qh5iZdEYPs1NhHukaGjdhFrfcGnvNc9
mTyXJxAyKwXEfkedzeACdR/R1FAA+x1R4B9FXEY+mORiom9y+/KZTh9Rx0bSHyu7
oHZJIJkPgLfoH2mEEd+N1VgtQc89sl3baZRIb7WKdVbG9dl8JAtA+BvVO9umAFP2
2NBPw9RtI064MLIXV39TUTWtKLfeoZZJd2l/IDQpvY+FBHV9zSYl/RmdjRCT0WIO
NUWJrpHlGq4k6AcVrFM9oeBZxVFVP8piZI3jGELRdZMFw5dyvIvh2Y+A14UJTcWO
ING43LetPhlnTkAr7hvqFw3FU3kKX9vuPBqaQIMWPqGP3PUmn8m2fcCbabLhlGHf
RExOxpw5Odba+zoDH075ty8cMCg+k6BvF5q5rM9T/6vW0bfWwTR7/BhFJPK8RiCT
gSqkXSbhzL+oQ4uA0IGyTHTf6Ss04CjilJTzShc/PKbZbGiI5h0u49H8tqZ1H3ih
DhFKgtTtiJvjIlmX4Tkb5BkAdw8UCu1bYGVjz+YqJKWs0A0QiSnfFuatmFH0VbQu
9zuDivnR7C8Juq1wPCWyg9vtPYmnAFBfj2vfClikSvSpTqfna8c2cC279n0kLbcL
IeXChLEe5/nmhhe522ChPZ8IH2lsC/V7FYGEs1vR9WT7rUCNxYgPN/2Gfz/GpnCq
Wy3pLBGA1EEf35DpH/EV8Gwkxn6kGpJDssP0xeosPyHhV3Th6LD4JRzQHZ9DJX1o
NCG92NRJYQo9WNXvYkp5YzSBObyj70vNOb23AcKxFSWhd4bEb/VWIg2BK3u1b9fb
KbAuYoeIqarv4o53uNg/ALrcXTCFxplRWuEG7V90uUeZYZo7AFiJkUlty29tn9WV
TOy0cNBw97uS67YBt42ctP2X4dcZThDKdDz8s3FbCySv76JC/ejBp983Bo/S1aUb
JsLX617bIb8yTUGeKwN1LnDh6u5qGuGfYH+ihVH9SearjEeOmAgIQhp0wKxEXQYy
huElcqRpGw9nvX0DZ0s2ZwIVFdMvm3LoL2L6P9v+cSbxFpto/qImS6OocJhg4KLu
g/Bw4qeweNOP0W1O0OuNVMennWt0Y9kc+y7/FwR8qjpoUa9mNTGmzvQOUGR5DQgK
5i+8Nh2N1yUSi4Sn6FXhZP0v46SIG+cD0spmy0haWkkWpOEBRxsm1nlzQ7lJ250j
jUhRyZEqoyvB/UTo3X3XiO+yIiJRQQZ9YfZsREKyZtLQVtSQW1D7pN/6i+rdFSqM
dN8H0sRC5kfVAiEe7O20pmBmN6Q2MwQcuZmBRbKpI3j9X2repnWDtfak0HSbzRW1
sgYX8XGvEAA4mtivX/zE+5xnk53KJ3Bsh0iRjg9VlmLw25L4aU6TFCXTDhB0KmSw
n4Q2B2ifKRZs+x3yW6AZOHjjnhAPTgeYxl2Ek27qtxPcYohzaOaJXwcrEnhdjMUb
K9BZo7L9G6Hf3yiS4V+IZYdC1bs87dhFwxB83TQrXPiTWL6AXg/ZXvRC+b75IRho
VHhYwLlwByM/d008XcSyXucwitQqYoNvR7FPqI9429KzdQrb4yh15V4KWpOcoJ6o
ICkFzpvct3x5F/38Us7btUCe9r+jQnAB56F7hJSgLW2lRBMn6b3dFxZkaEphLeTn
inuhaD+jg4sIeSXo4Ht6PHHy0UiGNM+YQjpT/U/8QHFWALgVI8ngsnWHG2HuUhdh
PNXLi5m2+60V8RCXfkWUGo4r/1eTT2XCb7D3RoBGiRueGx4NoCH1Bgz8XJSe+QU7
2Lq6KI+9kwZCzYX6/MnYeOdnfq1Vr6bEDVvvgY2EHH+l9oqfSEu6nLoFgxNEzzpC
C4HeQmstyP7mjBr7px6yGsYXluXGarFQwhsD0N8MjwYv/BTbpXFrCTRWdSVhmI0e
Ij73MCWMUB1OWsU0ae36b4VYy3Z+GR2ufDjNBFhgNrZvKZnfHl1tWYZ9JOxz1XJl
QHbfQAwos3fjzI/Cbqc92fX8EEHQNB0xxqQgejRZWht7a3jBQ33/9Q/O/CFG9imS
rx3wxjbSuSoAhsqmYOeFk/bwWXsMs0zTpJAwfeO8lq2tD45l8tSLVV9iC98TB3NC
WSyn5xJizi59vLXG0LmhgXHIGxGRwWfg0C2C/JoKYKsWT7cR/CgfgBBl5ZplK3yY
stUNqb4+0j+yf4KM8FQmuinrNLvqN550d1Fe1IdDdJ0N9UzpdZvNNP/Zmebbf/Xj
9kVqbkOrfk0GKZRWlBAFINg5L6Y121m1rUAeZ1z2juV/9IFBR40YbLKHg4t79mAq
Bxw1SFhXHMecKZLzCGR4WMcRRmEmOfJ1KgSkTaMfqDNvQizZweOR2pMUQEoOJtm6
7nRb/syQ6b1onBNg6uPICcxW+5Hic55yw53ntrHPk14Fo5zRlUbk9x9D4IBHRWk+
Wh0rpug+gy6hCLW3yQk8rIC4/IYJrfU0WbhJ7h3wP5FikYgrEoCDHqybJ6E7TWOH
MZr2UDG9sBKQHsNoK/pvHgy3Iqz2hjVU0lQ8FVq6jrTku5SbVUyWcwJKiSOO3gjv
ZYHGGyQSOmrjzYsMswm3GFXQXOb4xZTec/dfCo13zg/8ZnQ3Rz0m8Sd34J1gvIwn
rOvAJSn+ld2sAE48dv/LF9rdBeaYiqruxKU49z+FbXEIWFxFA9LOPuDyVu9xmP6C
Zm1Y7YTec1ERei7MAz1InW0ye4kbLya6/YSvWNQBvhhCrg+ubwm8LHtKh5WsS35T
/+QSrG7KiVVR+uCiJ7h+Z6p7qDL0+CS0kdrqOeq/b4Vy03v2P68ESsrVLfTd18Gp
t46sxRuatq908xAnj2gDPhbDcaqjUD32ZwODCHXVOsykM7cqjU3q8NVF/xJx5c+t
49JU1k6xd08TpYwmk66kvL9VX+FGk+V+qELzlbmtsJ3iRAL7jMzkl5tqbh9IVeO2
SzQPHA4bxtyql2VCoQZVXSYfsHtEoSHuUqp8kAeNDTATZx0zlhNy7lRDF6MY/7nt
0e55836+KFzXI6XgsOBIwm8/sovi9FgvU0RYYQYpi7uc/w6JWOaE1K76fZRdCehN
E41LIyEobkYHPOS+gIFTwh8o4uzsSOSRgAojECT7D/r1vSC/FUAtiezC/XpcuWub
sXltkvBg9jKAJ5MB4kzvtccXXeSXw3N9RbFw7EhM+43xIXFK2WMr80ZK1BiaNfy+
jmxqHTDFOkvG30OEig2Cf27HcKjeq5DBgewA0zNxe/kTJrbrTpOhwCgIEPXOW2Xj
XryQOdiL2TrcFf9G7Ve5pR8xkYIyI+r8bpKaysE3Zoov6e7HPBVL6xI53PhYAzRx
w03ZmUmO5iIRD2JOixkOIfsZCEEpkDXuSpHlr622aiirwJ8UKI9cK4lF6QfdvrAJ
ghWEvU5+f00RrK7ecXZa4p7vVLWPBX9IVrblhgUEjmAijcWkKYuswejUtohlXVsk
KLMQHLOp09vEPE5N+gDJX9YSG6mJJwCY5JqI0Duc4E12JnlMP7kkHUsizDl0p7l6
veuQ3Af9ltJEHmzFVlVV2/rwMKruBvB7FUknk7MMpylPxDnn3F+clnkdK7XumaWY
FXv0Hglm1S0KdQzDVf1GbxSPcgsms1duC0p2s/dNnOkSqvG18VzPY315kalO8BbG
m4l7txzNEbTGh/9/1x4FwJLVO4oCxsCZ/YufEBnAZv/oGV/6+mX0pl7V0VQN0xsZ
yR/3SZfNwno5VZ3SUR4asgNE56c+/8OeaIX4FElXXh1dk4sE5bqFv3xAaylsWViI
97HEIgCA095kucybmpxQBeQa6q1O/le1iOtS6Ofv0ydaMSOwTI7tEnowKpYx7YNm
KJaJgLEDV3SUrKwlCFXh1ZdM15mPRbHzUR81XKxa+O/opyfgCYYhcHIPqpUghWVf
uhWSyPrsDrx2qTvbfUJ1DjJLhT3nzfIZ9H7+Cs3AzrckWssjt4qjpnDn6klP0IEf
tNaYNYkbtK3QART0IvTigptrSYjpp9STBl8MIFut4AGMFOKYwHbxyFqsaq8+B+N5
XUDsV1Q4ov09d4vc8zmvkEQI9QuhwTqdrvSgR8eBH4R0UXp2FiKrh+lkk6bAKaQo
6mJUzcDiSOoM9V2KKxOeFXxWmsMRNU7PqTdlgN+M7XuFJNlkh3GvNo4iO5ayNOQy
xMkJXC/xShNlZrHZdcqaz9Ezdx4YxX7Q5wGADzvolPPcd0KeGovG0n6eEIbt6ZZ9
9XACOcC+CPqg5t37yJiPiGZQpFX3Q7GcHSHJX6C7JNT1tCUQKxT/UO9hCjo8rMY5
B0uVacI67/h6rSOGf6nfo8C9+4O2NTPZDKZ1m/YYOePjPz9sUpl+SZuUkDFYZJp+
pLGDvHBvkp5o21VEsW+2pTZiyokk7wi9Zcw4m4vqRk3ApEUiySqtXZTlBTgxxSmr
58xhYoZHMSHozpZBTS42A03XVqsW6M9D+HxYnUtafoHl9unCSQcFCDWkNDdAFrNl
1hNSj/xKe9BoRqvNJsH4F6mxGdTqNfxxQ5ZsBuggSJV6dP2bJId579SzDw8azO6K
ibs2ze+zrwLMsoGL3b685UW9VjQTUw9WW7D3uye4+tmcBXScMBey3X2kspFoOsw8
Hzsco2bd7aMait8zHE4jlEMpNxNztqFpxYrVbQ3vO+zX13Td7F5LzvQ0+Cmsm1RR
4pubV+v/CfAtumfevrzp3QWSLoGfhgNH37WjkKskYIcZ0v/6WNAv7dpY5WGsQ94K
JLcp77zPFNHIvsZW57tUMqF60xSRqN/sc9r4OGqCDYab4HE5rAnKdz/ocWMt0jwj
1KMxTJCoF+nYF1jUjvl8k22IvRlQiHZfSdn8hUzDNnBM01E530AoJhs9ChdRwAjI
vm3gWbFGfS2ghSRwdg7UHSCOuYO3lObxe1dGTFGWsd22KpjcdwAxHHpRsXuomHtU
ZXWzXtvG+ohZF4YsO+oSQFANP1S1AWYVo4LOgtWsHyrvvMMHmk4Zx/mzfVg+nW0M
b2WbrS8f5XFNFULIhzB7W9K8Gb4C+gJDKovjn+sGzdBc81VWeNQKu4PN4c4+pZzs
n3/9oiEMeDxXncCmnCrlfqPFeMUX0eyTfczZSZhyf00kQpaV/F5qQZLF9/Oc6gyO
T0+MfgCqf/g6R8xrW3uMu7yuMmKoUM2ZypiXmaDVxJE6r3p4ExRXpRloZr9fKoQ0
e1uaKTOsRAOUZqUCA1YINSZfb+cWqbOv/SpxpyUQmTrtJts2sz/s4EnDg5l5aLru
iSu0HfHMQ1Ayd+VPGY6cYpC41iVakgstsCBMbeWIuDYbJddkMMEY7G2gnPaHMU3k
Scx/WSMsS6wVXpLskkWII1fWaZeTFZkmMyIiWVE5aNT0Ez/FPp6AHMRLEH0wRQz+
6/9jRLQMJW2ij96ggGti9o6jgwOpCU2DqdbhGFh5/cwIB92lyPekSdOEulT7H13K
IZyRv5eH/DuJQrLe2Mxbrt40Nu7scbkRowjL8SMNdrDmF8Tv48PqJSBerH6KkAls
p3QHHHeDVeuwAEQ36gJrFAh8sDuck9se0dBZsq5lgQLh64zchDomU/SosiA1EIf6
Bt2zf3yBNek8Gvh+WtokNBZx0Ng/yIW3o2t+EJls4kjtwTZtcZVgi7Zc11FnqFPA
u0eW7aQYX/6kg+jLCsyJrZirM9rInouFTvNNZHWDGlRyuZ73J2sRLpzihlaM4A4q
isBWjPriuEfaV1qgVb+FmpkH2rdf0sBCmg5njrMrA312mT/jFE3aRd8LEmNJcr1C
gbI+nqCO3FSBP+EcvO34SUsbNdMPkA4aHxyasoZAlpbEFMUtFSoHHrZ6BCS8DrhK
tr6bPBn0XBirDbwrF+D3NpP28BQDRnJJ+rZrD7orVlkrAs5qcXdNp+zvNMpeDCqp
Dl6AnWNd8AMcyYoOiOlOpyR15pRGbOySB2upP4jKCzTn073WrNyaa6S7ruIBjTBC
0p8ND41/imf07T7Jq+X2snUD23WPZwDph6oQVwSFUbLKvUY0eYhD9OG58F/qCWWo
OSWHtcYZNlZ/f7SYkugDZilPvCbRa1Ln+r4BaEiZ9Q90lYmzrFfnKOTAIjSIdi2d
o/V5LAMQH3w00FfzB0EK3aRzyKeeN3yYlJ9/TFagKGRSI+UUj5X1Nc0ioiSWK3MD
oSGN8vRcWN1GDsDHJ6z4YBgt2UpO18cRP6diY9UfrOtZ0PDDoPRrweAUP2oSQoq1
+UHj9IY4mbmSaXEwdFX/W52WVRsBtxr4zxilRxX7jYQOFTHP3ScXNpyHtxZztIpt
Db163uETKNpF6e7iXHSLooQWVW9YyGePlK9yz4IqS/gZ0Kc0hJNTfoIfU66QBfl4
wbzxAFZZ2388Esyuil/L4ZkA4iRS9XoqAJh0itrLpxVsu3rTsOr3ZzuvZg6x0LkX
FwyTLc3KLEyGi34PA8comACSz+Qf6E1QooH+pemsHb8LgOEDkh1YSc45uT7yNA0Q
XjIi/0KO9vaVjE8aDWWXkSizdDm/Jf+fmtzAAs36Y0KFqqV1+AReQk8OjHnl4qTe
P5Jo9MmQX9K6mhyvO2a1GpqmOGQ/fBV4PcyaLiPc0Icvs8hb1Iasu2kqGv+qbYMO
eZdbaxUvu+4/hi8aQuytatJtzoWyi0flEtx7grZdk0vtLrT8WBApk3+yTKU9hk4r
dA1y4Wh4ZlRKgwlfxSLXtE9haqxVVpY3UOqkk9XeY5hpO/sB3ggtWTb43I5hFDqQ
rcoT0ViV+aVZR/1u4XgR9gJSCpYwwpa2A2jNwsGQt16c33IpyXkKLqeB9aWzRoH2
MzXRrSbd9VaboPy38XqXCMBgPB7DkaZgYqRYylhgedDJA62XfNrD+cHTS1UhW9cI
b3dUXd0t15EpDxXsanEt+3bCofZpNUcmPyd0nFjYQbQJg6bMHvZTTr66WNnKea9u
O0D3cVFUMyOHfv3aFHyqa3kf5nwIjX7iXTR/rt1+u0+8+rEmLjqKVqphFq37R4+g
g6OkXLnxKJPluM5h1VcSwGt+Rpc2lajg6Dkwoft5IIH/n7934APVI7RGqzSvZ2ie
Z+tyDqCtsdSHaWgiQFaj2zAgRvBIjEfxeuD1svGJqjbuphdPsZ+0/63hdLaJ8YwK
RNtCh22/qABXxrXt1dunMgET83G3Oe5cmBOR7sChd2jrRLf3v+bg3ptwPJgr3xUA
eY8hhBQRnbtrPHgfrS+d44uHtW6od7t3ZopNsS0RvkkW5PxOy1XONXHpHdQfmyUH
TzpLv2kt1wF84hrzyANjL8TLnxBav35CnecNqA4bAp9tKc6r1sJGjdcsvOIjJawc
9GGjw9mosWfluAxsEJCvZPN3QkdOAch6UoYEmU+9HABlMgB9360pGLXDUGXYaWaj
nmg1ENyQxCjoCu3wJ+uXLZeDLn1H6SRr4C/9JL4vD+JrknI2rdPC3MjQJ4tLpxeA
KlB3HGo0z4Q089NggZgqhGOOfuaL231vX11EYbMryRzTybNYh68BVfLxyfT0/co2
aHGnWWP3dmDKrP1NEatt71q3BpmWWcweFib496eq462RuC04nyIU2ETv0AhxSFsx
WsNdhnygeWszw8RGUow1RkVYeY759KVJkBPC7xnz4trIUudG9vhpMwyGIJKrxCK4
oyvQEZQ+vc1Vu6kXRogQ1ph/7WPbX7xWBqrC0VCvS05eYBOSdnLPA2Xfoe/mnR6v
d0wlys3+/PqUwNvh0D0jYxsjyRdgBRaZAPxZTGBfLC0oRCmVnBrvJYsNAmA1Xlj4
PC7jlZ09P1nDmYqcHNC9wOqReRCIbl09VDA5+NqMJsExcQrgUb88ozIGS1ijPZaQ
4h+VwZWXWGXXQzMdBi5dN0UaP9sJ5mHXrPpiVQVFHFKxVZD8xPMou8eDhcgaMxjg
qsUyH0iAD6QpLfR0r/XW4YKZKRpa4Wj9Ds3OrGgHHytPcWjPFNdz7ejwwAVw3mpk
JEvJ2jMPlSzbnEXfPSPbXVcq2Wl5Q1IsFkuVaDBM62OKacOmDK4OeLZ/M6Ai9rR2
S5JHZgte9oBDBj59O8+vAKlupCw6QPI+3Z/Ie3VKtuChlbPbj7gUc847HUMn/vMc
/tD9rRVY2MNYzVZBUSp7udVlNt+SDFvkPrsm6zhcqm0gmQwNfSemtqS5IzoKTnXn
q5+SBV3LsXikiPwNLShJMbpG1n9Q/koPYEz8Yym4jNtT+tdKlGTFART7r+FNdnW+
fJpCf0h+Qbd0iqh41DEV6hJ9irkGKsylzTDjgO+fXQtdCOE29qBvk+p6Y96EnIP+
1D+fKyrST2KMAVY0eFFonzSOVYeY1x5TzqobkhQlG2z/tNdVARLP50yvlymA/sIu
rKmeH7gGnQHdvdzPt4KNCU7DzxxCNqss18skTSDx+hCVHz4W5R4UNkF36JcXdPnl
GGTrUzjLHA7u+3gapa24aGouH8FwZvb2kcKo0klZe7IPBtxocH1OBimaII3fK1/g
UrIf5CEkX67bphMWHkaB90fQK4bwtEjj2SJY/ffmucbcT0STJt2xy3S5h8luFZLl
UMukW86rBtnZvygwzVlF5hg+BMZ7fSppezbXPJC8ySjD2GEO92XFGfbdrhFsl+UP
CRJrDpat1/6cljRE0rlsfoCv8j7hVxAe8pPDV1wD5S9rqbX4PqN/mrXf0Zex5BdX
aDpCIdiPElZn0RbsPU0DfQSZ1QinLEY2a6tc1pqVTv/zJx0t/mizydS0FNBBznEN
eEOAsBHIB8jnFI9xjxJkOANwPcX116YKl0omdcd44zSMh5RBy/kJ/1eB6E89+KdP
d4pyhjfmvrX6k+RcHx5RxPq+jWvaQLdORuu31OG5/fI0Y9hiMUo9hdjagWkUhgcW
CcTCAx6/Q+04UW8ikEUI6MQJMudhnshPokBqvXLTOJvC32KFv77Ye4HT2Fno+0dx
JHJ3rZe5zhnWuR3lSzxyTndk0l3YnRkkP1Kq2d4t9bZOkHZakmofRU+ePHCsitMz
ox6zue/mKNGpgfi546YtDUMM/QnZuB8HNOK2V5pKCfnvknmUm5eJ204NyGprbl6g
wbcHrqC2jsA/Dwb0AAM5kKYIUeYAnugpX7aKUDmPRsmfZlQ/HgpaeffkMMqnGJdA
sltQ/1etEi1pKa5sOeqSbc+AzmJCdFI6WBw0YxVPz7F7qKeWE90gZvUBYd1hrt+D
zRPXXmb1ugtY7W6iRVa8PJcmJT8rhme6zkE9yUAzyn3VJ9kX/iJC7s2L0Wh0yALI
xQJ+IYDpadsky/QPTsYfH2UHZ+3Mlgg+puGbH4CAJMM1BqJAbgMcmsxpCengwhIX
Z/lC8TrnWjFx2NWGapI5ukVk/VWHJMLCUVwZXNXAkn6TQHJZRG4qCLjVgveO2C+6
OjY9u0Arl9i9jzrOSgmVbPEGMaGula+Plbr5q2D8zh1NPXekZae+3HG8QNvAD/Zy
XNO0qObXoVOpatK1Adt3oMFj7wIn1XkllWZTTd16CC4dgkeR361dMazaW4lMHG4A
ftvmP6PM4Ir4Q3j1UfmnzcDGLrOChYzx3+1ULyMqRT8mKFwF2NsO8GhCgpy7GrIp
epZVYqHJ5VkpCTwzMROaJqzHmnMCiUcil2j6DHDXRcuhqty3JTcLYNxBDcnYB8jK
vOGoyULRQhVA8IdjNjAJ1oEXN266lm/MEyZODXsdFg0fyPywpydWfzr8xVjSq7hE
Sa1+ArRmrDMDcxYfyzhrNl9aEC8+XHn0AefPhuKNeseFdrMnZ2Ct0WSt983UmyU7
ooygYeqhKgnYnrqpGbiALO8MbNXTXkzACiWMO2T23btOYDvGRzrUVEVGuZleAMPB
wvSC3Oeh2g+Xt8ZSJJCSSsKvs5ueI7tCl0AYrNR0uvF8tQKKVKNIKAttOujJlS1z
xAakk0FcoacW4X9e/GuvHr4Rg9o3jbInFkAmULoMDZ4+YqlgIKvsVbL6j0xv1k6p
EvYaKhpZQ2mGZRDWSAHEfiz7ucJ/WozknMIM2X3i4QEhUwceSAIAu5c8C2PHDzAs
4oPRQnhf6SuslRzYqPqTD1lqvD6qMhokkx6Mypb4r9KjnsS1228hD4Cq+R6K6JMT
iHNDa9ygDD81w1FT/2mOToxvsiEDpc3dpHZcB5TiWAQ3Fp4YZk7XFwtmaP3Ch/7/
K9FP78irPMlUw1bJ9bf5oCrk8npajsJSEegDtKuYrc1vkhGp8KJrluzsywHs/4j1
2vXIHutMlSSsd0OjJw1ipPd/xy7DMmJ2Fz6CQwY5maLLoa2jGiTXL+1Zy/ulD7BU
2FU0FE9VrJ5NEPDKNCPj7UAnrIBu2unvqIhk/yYmoUGneF3GaU0OXyhkNoRCUZ1h
+dPwUufwBOF7MUY8jMxqEbYZEUyAXcWWHLugpyrAy6C+Vp4EcLOqeTL1/Qod8qWA
OjLdTfhnrAE2TwJdobR6OlyiIVZtL2JSL0aNQjHlcDb9MdZrikwP9KzKg5qFKBB8
D2tr1/fVCj6S9AYKCWpYzd40WY9SF7bsVgkcndVbv1xeGpVxeI880TNF8ch6M+L0
EXG5CrnfudD5usJid0wloGNP3POHq2GIZ1JKc95fJCewienZRawITiuj/jO2WtBk
jhoHJAdcENUzqZy3tZ3YE4iCcSH8GSkAcMglp9rSbe+MxKDIkhQRj2tGa5lhtWNu
3wWcDEQ9nThZlwPzMfJhWMsiQ8zDOkcUCL2+Xqa7ijQCVJQYtlRR5ou0McG/zj6e
y30bOC9nvfdn3oWPMhvMeqkHgZIqWosUOSGU3gorQRV8xiW6hzNhwDRF7HC/JFu0
EtRAE4tF35wD+MhASwqDEJFGe7uYn01AvRv1sUTlsPhFH7mo2AJaU9Iu2O5Oq4kX
47dnpJKOpzvaE+1oP05ybPsf/g+eziWPVhFGbtKXsQ1dyMEcQChwwMBUnsbvJr4A
0e/aRfdA2t0bbpnUOfZ+/vuERlIAr6RC7pRrlSGZMl+Ccv4I8A4L8ksGC7mUhZh1
vjFXI5JiYleEKToZ37RpnNYLS+pN5FHHYa2K+auyhqj2bdHyzDpRdVCHZg08xULp
BYZumQROD52CD6SzptuhpemhliHTEUVtXuQDqugB7w2rCMESq5A50BpvLSIKryPT
LAJWNzKrqpjjwxqyTtArfxjzCxOz8tRl15qp0AZstotmQSathH/zxQEQljZCozZn
doI8/rtMp21VJS34cqNP6t3BKBHBEChWLCE5blrAzuy21sNV+iTAgyKZC248i0U4
rQfxTpV1RftmRRrPjAz2tRE+hYMR3inldnn51wlizNJpRtmi2xh/o2AE4OF9Lwrq
g3iU+GoZmr1MNyIRy6dNjg8oHa3/2yOwQYVarUQhnIwXKjpiCfb3mea9mT/04mWe
SqNVCFxZjVtzmTWWAq7dvKm1Ks2phqRpp4ln4aVKckgbCuY3OW2SFndwcXvC3iS7
d8FT+m//54lUyEegHvB/+0aUAYbKM9GzhUobK6m1DPhb5/BPmZ6rsftrhsJcvg4o
1yG7CVsHzIIURmcKdz+1uj/O9ikicK/H2h86tzH6W7fT8cTa/bWN1246GfQNZrgv
U8sdLoVzs9ybmoeYmdjC6jE1y3GIPa4kdSWkYtJ9qWME65/bI2HDaXBQxtFCBN6g
heYs/XHXHz4InuWCh7gC8rmMsntahH4PbASlDk9j12m0mLelLzChSAiRGDzc/LJF
e7rB/iTBBnCP0rPF2W6Nquqjd/xLF47Oxi7wlbNH58lZXqxb3AdSwqX3+fekNy8x
bFtxgsIWlC6y7i/XjnHXsQ4bA5i4AOsTV1t9m0aDMZKffOoWhANWIiOsWxXAXili
lHbk5UudVMN1/ZfigBykzRrgUggq4dwsx8PI0aa0z5mhTaQQ6Vt1gzvbxXbc/Y2y
PUzYHZa2izhTTOfK5y47qMxzom3Jk3aNKi1WqMlQnohZEkuJMeLpkQWBqXw+ZzJ7
Z4UwiIz2eujA9mk1Eb7V78DIHensdZ6+PW4ReOn5Fkq7Kh2IXq9Y3w1biu/FOqlW
mU48VaOSId9FNYG+IIpBRVKdatjc6N1wwnkzvQ47wge/mx7JsGc46sRvU6vT3cnf
XW+i8TguGDOCTlvpsmqF8gipyGZvkePNrCDtZJ2I87B6KwJnv8JIoddpye8PFeVA
d1bd+euEB8U0Uaf+Lx32DXGVPF3NLaby0Kjq9MMu+R6/g4FN1X6kqmrzNghVeQc4
JLsr9JTkeU7LVdh4akEdhtcW2YdObi9hTPqyPHh0PkOHTDvKRbtwbTWvSXNI3Oo1
tMizESZJdBc0Us2M6UiOct+Jt/oka2XXDxbV400IQyrxs+HV2wU0nzfkBuz3dRsJ
clYS/Gu2B5hWeaSMy0bmzNZBAbaXL3j3lwSVru1Kx/Wola9XtOf4nk2O6OHXSoY+
tvOj7wzd1titwBeP8s3dNQZL0PlRy+att6SD1JNAfk65HwEfuxVtYQNKPQJVGT+Y
x1qr4lbeTlpXweHG6z2LB2RflDhGbve2JeLvX+2A8mGzavXmTeIMqYlfMUoPo0zs
3zoeAqo3Qir40eipSOSSKBfUFd0b4QrgyzXTUAqT/ITn5G4RmVNRKAwt3IqCQuu5
8Ye5klQehOtRC3k6Tv0M31zeo0Z40H9+gLot53WeLJMZNc5M3tiN82dBUU6DCK/p
Me/A2zH4ugQWQ8DvnjKHcaQ8nxufc9PICsQenkAV6PVs3MxwMgDXvxqKFaSvRkhR
lok4xg7By5/StSBhWWo/vrPVk/xnVdp3waVU9En1QAIYFWjK2If9ZQ3tTzWHWaSY
xHQz2HdVOJ+6QwMAJ0aEA6fks5uFqBGF1MUGDpJjkwE0cIautRMVSS5agJ5/TUjS
GGsQQCbx9bBBRHbLxYgHO4giF4qInjQ4HuHdYokxl0JHz+qIPMTvu76MZAYy9hAB
4nWWOR6NS4otNDUagbEUONnAlGjrVntJssJ3n3cGMkF925n3dJEh4LWtC45wj1oS
YsitSUcvmkZ3+ZazkbTTerQBJIxnqR3DbZTLoda+myoFsaEUr+LslM/rQedy32iF
wgOwMBTqqLiKUjoWDw2FNFUUStRRPzTrYY5iAmDcJIytyeRYcTVM2caMtKkjOdO5
wkGSeXXd+rruth4rUjATe2B42xTJFq+vWWNMdDeXMY1v2WPnEYFCAJlsBU34JOMT
ttm9q5r99QMYerWsHGMzs3fWniv6k+6OqAYBFJ6zn5N2PPDR1oYMzcPnR39apwcn
DNTWpRKEnPHrev/wGImbrwyDMm0Oh0affZgAgMn0Vyqc/04zhviy8wTxeEzCicCT
Lf+zfzVzPQebvXDeZQrsSgqFvUgbEjWiWDdK8DPJsXzA1saMBDOmF7s+OmQI1k0C
IbZGe0i66o/oEs4YdX6CRhOPLfs9qV3MKWrLezPejYX//23vbskxc3V4yR/KeQE/
Eq4b8s9br6g42LJ/ZyC9Lo4f+3Tqa1Y9gcXv+cfdwGswuBRI0ELFjPOooN/TLchn
hQzA+1hwTBcXIby0W+NgR/kLT5blkwt+MS+g9/b7vU6L0JJHvi+wtiIAGlx+C7V8
jr6XH+pFmLBr+Ww60Gw2gILU7jGLV0+WQeYEcNu4kFowl6cWp8n6qZGD4L0n9XVL
HniSK68SoM5+2ot+sG79rcTShSUkkZs3M0seqUUtVA2GnrfmFQ9tdiYzslyV+Fha
nQVEZwzFtVtVnW3RnEi9fvUwLj4hvA+57pAmLonQJgH0TY7RFgrGZWy+3jqfJfW6
mXqdUNmY9F5xJPBBc+DSwMjg4ZQ3xhOi6ukWO3UX8vMl0M6V1UYTM4iOlHIoUiEV
z6P3U6S9Ty3x2kprq/87cYNz5Q3BcnKIdEcLs0066S5Hm4s3u4bIlRRg1xXYQYsI
s4U3BjpIdiwuez04j3A5DwYgMPwBtHizazkuVBljsyQ8RA5+oIWfyhrl60vMXDgT
vsRzuIgGNFF8NiC+CdAuiJGkv1zdzk+0X0wLJWP2VVrgT6lEMMLOSW2iv4DBJ+cT
RjplcRYfYlT9VvZl2echUQol4ccUYS8fKa9NWmef4cJFRb3cgpjO+p8g0iukLZ7k
v1gxN0qcYjMy9aSmSkMQJ1kQh1lwfPJjcVgdbsLlc8vg6UsluE0HsoQjIKIuDuxD
Th0O6yhW6eKCb/H3JH+OwU3aZTbvOcD4Ixrq6AQn4Tr4IVU3rPZi/Cq/SEBUu9dx
WFzYeFpyj4xVEWR48yowf0LggM2Jig9iJarmWUWXU1ogQ1ZSaneUDYEDlZt2LSB9
xVYxug7fRysvI4XhcP8wk53ysWnJkCK5vn0UzViG3AiZ8ws6ziCCaTG21NdL/mrF
Jv6Srm4mwBd4zb+B1WugkfmzGHKAGUxWhKo2soVgm1P2cWTuQDZxoNk77CUASgkR
LPPOb21LRtvnJL4iXAo9BItL83ByJBMiBUgaZ/UNUZW2wv2tWPZztHQxxWeW/9jQ
7JbCSUxUaFGC+dZZlZzfROX7Qy9BcfHIjZ3mZKafTZk5UQA7uBisB8aUMwVqrNBr
LSo4LYaf0+TO3XtvCuBXvu+KC9j/0ziM29foPCG4mEGQzSf81noDNzADZj2lt//8
VeiPCmgRjqUZiptbP2x341JVijL4+jc0n0FyZZLYFn71wDgKNp1toOVCbwX29Gk2
0vCVD5tEwE7m2NDjiQimlR9OLzgyiQAdo/LAI6bzCFG6TEbe5s+JyIfYhE7p4Oaa
dw2GR0X+oqos1lShxoXMLxi/1mvQEqOypWoNsNac17qo3hPzota2C4/Etu90jGmk
qVIE0XIQLjjST3LBCgsSIJgaedDGqz8nu1mvTP32pvIB2ag95VzEcqRgmZJut5Yg
xgMp+PTDGyc8mXG2SqgehduMz3ZmzrWOcglLXNo7DbLX2LixyW+bm+RHGbSQTgcO
7UCZ6X4UtoOT5+WJCTigvIfOFz+vBIfobp9Ft1DGJUwoa9/NRVD97sKOOCN14Xtd
j8+zua46Izj7bEju1ICh1Hc8kZlfWUbn/cwBQbQ81DEesuXqxF5n0nJE8gISXyqq
UwqN3udVfPoAtU7dnHhMiq31K0eH26URJPHJcgUY8LWMbTAifvxfh57Rd3z/v5Bc
cZLky4tPXmRZbMDZMurO/98zhO432PuWrdDCLfSqkj3xpI03fKmjy582Rg/XmQvF
odzTiOA61islODIbL454r1TSGePZ9IfuPuF/Wsv6gyvfk6c73T7cQPnaiCKdyHfl
NQeelTnecWfGG1JcU/OwXQEghTM+58tbWWKdouMsbGuL09+8MYEo6YxshsAGojaQ
30rLQ7XAH7BQ4yK8rBVpxliYnKNDNDpkpkwByIRz5f8ZLOEOXOssdGzzWB3OOJ0R
2yHGlkqduUHW0KusRfeJ0256m8uV10REz8/Co7g/k5EGZta5mdFQrtZ+xVoEU8iL
L+MpO3PjTx7WsZJBP5nDyBFPaqTtHZvKsiWHz/bEye2LXeyUXmMET7XWobiLUbG+
5Dvb0p8r3U6F0QBLiAq0Tenop3BFVCFQ4bkQdAQupmlqN/1WLKJys84GaemOF+15
gZq8jXB85UDrV1GfJew9S12usyk7NnvnwVJ9ZE0bLipGs+0T5e9rQRnDQNnbTx8y
iFZV/3xyTkUpOS+9T5m1KcpJkYMBRPv8iAxi6NropvpFArNY1qfzjHPnDa41ebZd
ng82Q30/7kQ1fS08PRG1QTpN9RYHTB5cS/It+im7d4FOTWqa4OVDKlY3XGz1Xrzu
14VXtygrKl+N1R+GPAKkSxb80AZk6DZAoyQ5a7dOhJbBnYays+SCxIwJ+KZI2FsP
fna3gzcYuWoOW3WOONa5zEyWJAyp2C7NN1pnefVH1Deu7dfSHrM3IG8FGdLz4H8z
teWQEBVWSWRorF4V2iZht6p0I3KLAogbV8m05oMrWk3SZ74C6hShXGt5AliJ6OpS
8ww97+egJfviksv8BMx/XQlTQjzM17P53zcbisFeD03jusi3booWmEEIE2i7p8HW
FvXOXRsZXsSOKKuOGEFC4x/hlS/IS7HcoKjtJB2sxK95+TXPT4VHjmL8Tu+efAb7
l5AQ9Sv16pbAtwOngJIFLh0q3ObEAbGIYQSp0MR0ieQT8ZnPCA9X5uRAGLjq1TjV
LDgBnKrOmJpGnasFHXV8ybPdTPqCHC6+mN0UJzKqN+HsnzwaR41KLoQdoGsZavV8
w+cEcP5dYyVKd+80SQi/dj2KNTRCinMvA8XAzv62XwIQAUW+xNczh8LxotCxseCm
FPpg55yAT39x1u8CEW7y31K9n3vmFqFqzItG8PLOcwDpwTklKq2kMeeg6+orOvcW
FRr9Tx7gbspm/sTDrKSJthHWxhrYHgS5A/kCHmnsvAU4PSHTW4SQzN/1EPC0/hP/
SXLV3iBnQlOQUHxnKPM55IjMxYv/Ekp+vlI/f8Vyz9dM19ImVFZd+OM/IJw+34KE
zz3jAl0bNSBm17ltqbA+1PcnucSDaW3i0WipDli8zOLfjav+hQKml1ryn5jPqDan
phX2sueEgwmsBUi9d9e0XgQDzAPxK7qNs85FZtcGFmDNFdKm8tNVpU9J8drSuRl3
962fE9DWT/OsaJKQ1AZ+zfUr/XfEeoV0RG1+wBXC/i4Oh+pJSsXh5SRJHSuymgSc
eISCgxAh9MiWkuUJUQZtGrpPiwcUXq8XIURRGMCHWHy0Ibg4CBs3UkBytJiDYoZK
mKWZSFJwR4zTCM3lKLavAcs79RiyUFeEjMD6kFom5Re5017ekB1seD105kcwn+vB
H04t1sfaZkQ5EXGcEGzMXemwYz07mtkFhdTax+3mIcy6d0ubGlsd0c2zmUoLEKb9
/4WMkHv1JTaIcwKysUohCbaOquvwIJrvsQSaITVLeYOOs/IAQ9/+nYC2WPdRGA9g
+XBaRH/OEvW1L93aiKdgGRptL8/als9PVbDfe3XyEwMnpI7mqKIuh2wKv3Pn+2EJ
uaaXwH/Cui8ZT5pbhnhFhwf/5phJfHmyXxIqv+vqm9hf31CgekXmlKTakCQ6Pq9h
iMmXAwHpMNpfYfmXbYtDj214WZe+EIk5A1j8jhY5xnlqa3TRISmD7hN6fy5CBj91
Dgq7t0WzPOzkIpUvXmABIuirGwkuWIomsIFclOHO1/5c7wzfdTilOpcA/beSRsKr
aj/Q7SbOn/KV4a1v0UBAFDHdcwxs4GOud8PLvWKpdPnijAfsY3NTc0FWLTb8nsMz
fP0QRhs1p0X2IpWmuU92MUZq20ktizMayozVj6M935CTU0mjdyHAxNqGRsMCm9rR
eeVYR1L6Y/yd6mkbpiJ4pQFj54w2jhTEt7CZIrPVO6VfIK9v+UPdlrxCUEdDF4X1
rBLkMU8ICvuMGkISWFEcJAra3HXh0zTMpuBfp3s+FlgUk9y1WA9tqYycszDF/Eq5
Z8+nkQxBrHUmjDX6chvAtXlUY8xBCSOchbwM2mh1esYWhNLHnL23NIQ6uuLVpEV8
+tnoiEy/WOJ1HR/ok6MByVd+4kNh+xV9DtgjJc3Yfqehohcf3jDpVf7r2qbC2k35
CUkYfpITZuhPWebGp27leC0WNJe8b6tE0y/flKpZ1ClR+2zUWx+ZX8poaNXhn6f1
s0iUwzqEJI5L2vnqvr74w6c98iqalg48KNUoD7Kj26N8+nSjfcP+LJc2jnVLeT01
heu+e/H+GE7piXukBcnX4KndCiYB4ewXgQldOoXJ8Nk2U8KiUnL9EjjuulN1Q4Fr
A3BThrA9R1WPMe8Hk1zMeagWsly8TdIWGNukPsNVnbvtgF1i/1HIZAfxm7MxoW68
fg73veyQTw18nBpqUYzVhGt04qGnsay1bmbSS2wAHhViyU4g134Vjw0R2MbrNH72
ZpbRPG3Td9ldnxwMcsxokMDi5PfOWA4isYVqT0ePIFkymVPEsC9ST+GZbleq+OT2
Jubt+hGQr0FCENN0pYm5YgBFbPUdEp/qAfT1XrdJUC/aCCkrgzMguHoC4k5dxY6L
wfKXvD6y0MCqR/Ob7rgjqvWrrcmF0zCIPSQ2sgA0U8xoXvmDBf4kb11AsF+tK1kV
XQWfwf4SX41DVGHLDyCVQaVxDGg1Z0GElo5ka8qVnJmuVgFKeJ99hlhseGi0zBJE
7SquAG90l5BVJZHLneUC4FvPwiW1nTdzxiQhBwh7R2eHbJuvJ1e1tOHwGU7gzWEO
pDHjVFlaIUwmeTOVGpwPppDhtPNpeqKgbMaPsfFu/0OH18u/66E7oDRBsYMVDKy3
A0WUsJUW6JNAzqFKbgeY0qQ0xdmNH4+jIMYzlQcDCZd6zmWc1OS1clfcN/iv9kui
yi7gXbxO/ovEVQg0Fe3YsajWhL995F/xLOGd96EWrL6cahewBQdi+X2u8a4V7GQ4
folJ7VgAk+h7PRnzd0K1s3ixslkxG/zATV79yJtcswY5/pC6543KN0UhD9qz7WqA
udgyEsF74DYiwE4OWhMkfIwzKJ8UHGBAqU0jdZmXhYQ1kaF0GTv1VjcboItaRgmY
hWzePUeURzNXes+WvYDvAp8TJmi4pRnrG5lTtxM6JZmjdoP2imBeuNWXGmlFMyrk
pAWiCN7jgnZM1bSIveGT6Tjvb/5JUYjqmWJYPoh8tfWe8hocHcCyC+mJ2S6khKD3
MtMFAYhhBFJRC+AAeVflXtwIBvKDn6jUzHsCQf+vYzjxA5DMN0cacQXLZ7eY+YPu
o4f6TixIuMP+vCpvhNCR47ZflP5csSSIhpCJLcNzOeqSYo9SouRLBBb8pUlMgl2k
m0MBXylx/s+Tt+vnJwK/5eA2BYzX0Y8V8+wlUW587iNPCQKhObPow268oeKSz8Ak
NiGJ7sQe+1Zp0+h5eybhHHL9GhEy+vi/ektGyMb5XIKsFUl+Uj47pw0rCaUNAOCc
F26rYX69kyOLq30686mC9UfsRlNFMRuXTGWciZxtiT8tGpvf7eQJQPrYNbYzdkdp
V+njBSi+TZZcjDrdl94/LTmReAI7QRymHNRuiGtpZ2WjvPRBHF8XraU8TtJg9Luu
oBdN7dhk6NQz6Ubvl2v1z/KHhIhW+32aSCK6jn/QEOhEl9wX1CwXaurv/dIVq3j7
e+3CMUe1B1hIp/KMfIbFFo9yiBFdUtEhs+BRHiPhi8eJ85+LWUGPb0/REESsLlCF
anrR3g2lYBfX2NwP7rSDivHxHB8KxPYShQWeUO1cFGSmG0uwRXKevjfQenZGQMP9
eWzCbLwItbjO1e07f0MQHpiR1Qd8uFkPDZywZ607brE/yHht34vtVhxur3GMomgu
IX63Oj/JUEB9aF6wnmOi9rW30QZDn1lkYIMNrANC9tu/7HEUoUOV+qHZEFPu2ZUE
xYsCq9c6kZBv86v+bWez2Ev+/MuQg7utNNp/5WV/oIyY6X+jwZ62gOG6skwmEzZ4
TXh3HOLL2muRXd4fbsku7ZIZ5AyhucAMpOokFdVDoFBokYNC+NSB9oi3peONH2F2
jUHuFFXbaRVWTSG8tRCYmWVkz7X38+dw57RTCMtYg3sg+9MdEdeCkQ4AR1A+RIip
OYfC8FkOZAYHhmRUrfGPl/OZf3yeUu3m8qLYyL3kPX9GTvNZNrmgOos05wjjOyzw
2cMVWZVzJ4GyRGWwCUpSwLWaLod0errlmknGxBKKiind/seL05cYKnqaix/Rmv5w
JIT0NoJLi9d/dUYntz5OqLkHB+SLQZSkpDxmotL5VK56GOLj+ON3UcrD/E4UIa8N
bOJFGuSDZzOuEa//NRD7jpL+1G0V6z2utRE0kayXCOcAqNLlz4KY6r3W8EWUdM8D
smCY0RYxXZyvY131zb3iaPUkfQKiSCBXTzgv3r5VhgoeOKxSf4pCFDReQT+CMGnc
qD/On9qG2QwLkzlKq5OEHShHnh1wA3oeTyUNBYdwhL+dAfBcQuYC5+F6mFNGEk6s
5pQC0G50dvuKOCizZ5/6H3PWmHu6AexcRJg/uDGpac/3Iiux1wrrndAMGto3vBUu
fRHIgixIyHeJ8Thp0Te1hDv4Trpf71ktZcHCQlSaTjbkYuMCXqhgIeDBQ9TVP/2p
qoROOnXHKsWmsu7Fu0xo8vFR9g3Jaykved6HPmqp4ijUzEnc2XzvWCNtX4P4yUiN
y74sOG/IsKMhmX5aWI7dMAipMhdb+SJOzBv0QHEg0JFLyPPwMaUwtGExjntD/nVE
X49wBAMRxYbcvh2P+IiSQD1S89sCR1YC9pwgFPts5QJ/ahgbJCyuZbqMGjqhVrTX
pvNWlu31TcmbTKGct+EP9Y6HiO+lUuBd+uGLEjvi8c/C7UmTuTT2Ps+f65xVTZ8e
Ry3JhQ2xIlIj7ubwT0kmQKl8ikWe+G40jbP2IlbXDylKOeYiadCsG8CDgQsMya0k
84mno/Epg5HNj9hpEQLFS1B3UgoU8TiMW728aM3CjuLY85Cw5s/o1GOx7JlpzBqh
icqFdmLiZ4ptQ3GoYNH0s4GQyk2eJzD6MFyo1M0+ezfAo1fJYMX3IOrmzDQzM0b9
te40PixksQXPiGHcNMzeEbTc2YyZbfxzjWAv0ypejDPJzXZiIoCim/RDOL8h9Ab8
JfLNGxmEHTp2mScTo6yHkBp8hx0jEtmXdol764rxlH1qDJYr9kml2//+KjP0KQic
NaXSfdg/yzOj76ERE8x+yrVC2I3N6wnbzf79SgtDYrHCq2UVDLoxhMC7W0UkknnG
y8dvhAqI7YGO0edpEAG4Azh7TGhchru3Asa+IkgK+d7Uoeir/s/ZdAJfQCpQftmE
0riRTAXDs68UHmeiamNBfTT5Dc1+Y24p/cEq9sTDTtmdcCeKiV8QSBWib9wrYc+S
8d+L7w8Ov1MXjfvUXAWWpl05QFG2dDDcesbDjJYDBhKqOBJaimN62yma7sfUCRZt
6iucWNxgnOSXUPSvG7koKL/k7GfdfRczFLJG2Q1DghkEUZCViw04TmR5afegHLT7
gSfwh6ZQDMeaMu/MJ3T2xruyRc8LKFmyYOJbyavrSTX5yJnVPjnlx1wd0YQaKjzD
pe25zvqQVrwoxXSWwF4pdVdUeP1ahXahpzEDJGpR+NuK+05vTpz2zl1UA2t7mBaQ
UkovrvM9U0Db+f3/bSEhshA0E+Ds9M+JKCT5fpEGZOI15VNEzyop6vXCxBcTNccT
DgF6tEaIV1J5wPAVK0031/ppEvt/ZP/qoJqYKE1Lb5N1Ey6R3uAsGjadExz+iLZ7
tBbniWcImfut/KRdIzNcGoVVpydpWfiLRHvIcnfECpQmR0ramAlc2e1BFzRpM7h1
YClhhsvPucUhRUP//3S2SVmCuJuusi/aaTOUm3TXOVkjZLYk6i/7lbis7n0ifFEK
EOkaHv7Rvgto+bc5c72UIBXHP7gOa6zdKwzP8jzH/T4gBVoQol72iTtYdy4m5k/e
bWEtYz61rHlD35i2W4u5FDVWnx/ZCNfAKOQNNCy5rZYFJEqSedmq6F00EdzosQ2f
NHtDuLBk4hu8U8QOEWn3tgmVXPZU+jIYwoGQ6LxH+hquj1UztPi5qHqeJBI9sSLV
B3vanmTN49tVw+HxFwXh+UDiLJTrtHrc2Upbb7RKGxsg6P2fUBD1TWAKlbUCDfgH
4MhiFFkm6wi3M0V0Cfh/ilXQMmJOJGNhxm/FupjD7HQbTXb3ezjvMfPKcZFrBstF
5ITks6J5xZDhvWuBXCznN3Qfyo/WAwOcewwm9hzN5r5NreKgyVPzHp2/M0aIymqj
VNw3BqsHaesYnG2nfI5Z0cO7GpxlZ0w+N1hd9AvFs6y+q8GHBO0D2yOs1JZ7y9dE
EUJbbCbN7JK/zBTnfNJQaE9s3RqZfben26c+Ij0EeQlh9fkik9fkQyCrTYXzVyoC
KoaNqB/gK4xTW/l2XvKPJBJFaEQsLrY2s5E+7ZzZ0J+AJb6v8WAZpL5393JPZAin
taN/Mbvhg5miQBs6sG/Ag+RxkschCiu0Llc1fBWMIUMEqSOwVCFVuj+w/PPNBCQy
LTOwXl4AiFryzhTaFA2UGv7uOp+iVPjTvbRipyeKu461391Zg00PbL4nPf862Irx
tzAFVLHgfYrHbzonQj6/Gp/Yxub/HzO15rRS3vS5OhUkk/+fQGbJJj4H0EUSSPgR
VJ+LBUHmJ6iSI9NcumN8r2noEKKRUHY2rPmYeNtPukVA7xmdgKwPCxa+TdWFfcGI
8fSKpXIc8N/FzaqlR5Vzr36w8ILKPCwgFH+7QRRbhc7JVNcLTPIOGm5blIyRpa8m
mhijX10tqnS/J0pyu8Vy7+lxLHklOi2yNHvmC7ckfs/FJGsUtUAUDUi3f5TgPMh/
WhG1kBADzVsnMs7Gs+P51BZdT8UVjezn+TnkzkL4qrFKZzzC0GzHFMEq8P+7ZjBF
JfJHYWcqeGuaYK5NPAaSsEyCz85O9sMAHCr+877QONgrDTHB4DI3FfTFwz9VvOen
8N7fcQFJA+7Y+bOnkq7/W0X0oDLDZvbh0l10EV6pfKNGpa1UR1Ya2E4RC0wBs4VH
vTWBS0rpJJQ91cked0dCqbLNmfinY5zSQDHpBx838MNM9A6be8AnZcoLkmE24haj
8rv1yraGoIZHhdGheMEq/OtIHwdyAqmqw96pA7sP8ILtxula93vlAoJjGrLv5jJ3
IfAvnJahsdTeE6h5oMgWqob7U0eiuw9ZO0Ramm7tXAbZjSDYkLf4VPJlDpA3iG8j
w410tVeSIzdAwfH4bPff2IaEKOo5oFbb04kerEQZTmbSvW5HJryy5fNOdr86/86A
CNK20jOZDwpXjptOvV5AB5YHdHCq6x7JZrikDu6hrCP4LW3/F42qvEHqZksiUYWV
+DvmKIGzfmk5/7r+tQZol44TwKbEDJdfwymWACZEDLgFOTJeH/i6jsjq4XRjWVYY
YTXPfCxYw+wlXydiCmpPbTXaKXJquYE0AoiKE/mf7WdNNcXVvcVsCPrPSDlnn3aT
nqojbb++Z26mT4Cv2inwQ1NL4Og7cbznR/mcXUpZTchRyJVXtjb/O+79jzVXQQLI
zA20f60YOq14lGj3wQeeE2g0bvgUenwExYdjtC3VZuBpTAbmEYyrVcV15ry0taOr
E+fV65tIdYGg58vewkCE+ANJi+w8N014qH7zWqDHwA6gsTSqMyf8sM6snsw2Ring
VE/tg/713twQeQBBtTQqb/OfekqjNrUQZ/rZRxbVg33S1qu7s2DekUXh6FLKbW3H
1Ku42wRVG0AP0kSda1hdF9blaqwnIdHdqd6Uug6ARbQND8kdW8ktVB2jWTZP3XN9
2xp3xv5Vz7jIOSdv5ct9K/qln4FN7NqmBX3wg3jDd9VdqvX781G1CZJMrsjBdClh
i806Orb73SVMKDkgC7JtQFyRhQZKZaLREYkHvBPOGsvcd6l8c7igIEEwxGBLfKvr
wHHOeMtCgOFDi5MTQIVLOgYvXB50mgzYVnR38wTCLV44IQ3IUV67MVH4tun7F+xv
oQuuvKSQVTox7E2JlzuilYmz3K0S/+I9s/jEYPhbif6lJqkfuKDQGTePtGs7wPP+
9POxRE6TF9S8YvUgNTvsi1pQb5xV+x5TX2Cd6Cren+DHmMQpGUtf2N1lIDDlf+je
3QK01vBari2SUVTUv+Y4GL1oI94rrJg9GLkRGE5oPLXm8Ot/oskOz2i2KU657045
czm10TPyw/7U0rxY8B9NrvK73Mdlkc2VpUKBHRq6F8GEF1Vy2yLyWDuxNZZG5Odf
+hlR2XaB7TxP2OdmmNpFQq424zQX5cULI+zFOzwViRkVVtjuVyQL5Y1ekhoCjLE0
bHcbZm539QD8QZEmkCaPGOyblNkuc0/959/rnNbUwIe+H/lNKP4Uh4lBCKfN2h6M
aWejz+NSWq9a3vC4zA0WqQTPbMutJlIxOjkyHRL40tLvS2JY2PqdZHrnCH/y8RF8
gpBDxV1kKL2ilUaOxKjC5Yav2/Nl0mNRh/+v79uqLoRT6hSENJzsxI9/o5IWXhsj
kkd95qtx9u+K1Fr3JmhTCJcNTMsAJI2gL/TSD2aU0kLJN0Ayc0/F9LeHVpXJwGa9
NrCLBBytofZ7r8kVaOHk5YhULL4NskMFZXMhFwHDRsXA2OInsrSSxrzzumKgp9mt
vt+hJEpt+LXbQMJQ1ObFJ9qXn+Zc9YVTY+Om8+KEiHjaM6atJRKzgt373T5FnE3z
KurB9ojYabW76I/bXfM9tAe6dnylCRzwM+Nb/uH4+0uVGOvqkQ04Q0tbniwCOk6z
1kuYX3HGR2d3fcT44mHJNhTGFaB3u9o3kP0/Zo7KjXD5g9CQlJJr9bOrW/5BA1hu
sUX/pTDMbXK2NIrdjbKb2+Z9PNz+MMPsJ5lvyOLlTC9H1PTZPhfIvDznhrXvvY+3
wnz0UZgkTnlLAdvuLH4KVWNoGDHoB7P/gFS8hqiKTJVWRfUF21cBbDX1FVrvkqx9
nGN6G5tIkU0nl9SDIlp8llyIL83eOj9on9kSsi/xv1ezZVY4YYTMBib1MvD5jFm1
alRg2ohXtO9dBSURvjOKeSwGv4ibWMynrkNvrBaCWniM2es/PYYzEDu6Xsubazpw
fgNltP8KGkGajlHEIPh96QKdYG7aPpMWADCI23XPswXWLV3CByGMRTLEVcvwVJCQ
ySVtSmE9BLMMmNjbm3QFkAE2tFeWgKcHF/omHAgL1qe0afGNjCkFxZQKeDlILq8a
ipu5C9ggdoYLhQoRdcBpFNRKTx3QVvleZUeSiKzhYnGWd362VoqoEKLiNfFV0swn
zfRyrDGCNYDYFbQgnw1/FWijkjdfgtIv8K5/v86ONB8OMiuNKfUQgG/xd6/Vzqc4
8tfN7yeMKu9IvmrM83YMhHt6hEkoym4ib83LpXTc9VNnjii7VOi4HZ+G6I1xMuER
0OJYtYD2j5JS75PXUCNv73gHBb4rcuAgV/mfvQGycpVMwY6Z5W0l+OpUNwjkVeun
56sGwqcuxFdNHdz3txZoh8jGrTF1nCGdlMWOfZ6kLOEaqbzDEIVU+lphGDmz2QSs
XLPS6o2qUQr92EbN2bsTaxQvYZ0MYvrU8lvHJ6BGxBVyzEiPXDj1Gi4370zSSNiQ
Fi+gIRPDpRlQQ/D2nlqUyoo+K6a2sDilbbJeACP8tlugwmm8hjCwNxrker7h8jXr
6JV/nILSAGK9X3IPljFBkI/7OtaPH2UVGJ8T2WZ4CNaQWEJ31HL6DqhDlsGx/V5v
zwqvN/l4gWBuCHKMWbAVdv12r2VDf2QodzrseHYfjEoE1DvBHnAavhySvMuat2x6
9cN9j8Uq3Whr4Z8HjpOujg7TLVKMl2FoKEaURxCzhCjzyGM85PXRPFB2XnKXUnsY
3OV3iW94JOBJtPjQuwWWq+FUiO2e7AXWtFHodXMNLbuJSAX+t5y5QJnVPiYbw3XG
XhVO/u7oDOydZejF4mYm7muJHdaOq2u4V3cyOG9eerEOnyj4+ynQ8sMeAt1NPZh+
VeDfX/j6WMOGla0owv6uQWIdPBA+6GUv8eC5A4pCtmbChc+EndkAAN88YEDw3Mns
1S4gVgy7K1OxsMA1NW1AL7vN49H0/JJIbp6mATmfxiQn67tUS+S/IeSx+YvnNkVK
K57LPlY2VQ3SDyVqOhp2g6IT6B8K7UrZvokGFl2fA02lbuRZnbf9MDmIcE2RKmiA
yBqcGYh6gWLkKsPC5HDR0cZes0IBbO6o73IiLVCfv2QzYUyqSc41VR06oYJgPDEy
MTGQqfJQ01JSnmTZzzqrQOxGfxRNV7qaEEc2T2cWZ3Ao9B4mbBTk6HNNsz8K48GR
GpQt2wAtpamE3v/DFH4HgHtDJqz0Zf0gGGtHwPAOMRyNci+VbpIU+iunMFOaEINm
sa24XUgEwn/aQexKPaRW/sN5NBQt5h+BOIs3sKlwjp5HEb6ig/MD0yfLezxWquOL
c3BAV9t8jObqGjKlSt+RHyowx2DSNbPz9Pney2DlM0P/8PW+z9oltpySFJuJzG6S
2FymcZpE+Gt1/VJbHjsJ0aj02i/WvdLeVvDcg0cSVWm8SLHJ6dNDwGqmB/NXBOKA
2aVScMIrXcUMLILVQgUOSprS9y+O8JVX+t5NxYTpvVCeYgOaA6xHyWrV2iBz5gY2
KqkIhBWN0+r1/MtSBHUIScIxSyDBambmEZOL3ErlSUZ0Vku6Pyc3oh4dYTXczOZq
IIgoVS6/J4MZVGPstNM71Y5YAImTy5RPPMexJpTTigAJuLPkjL6tpwy2iz+cUWAn
qc30x3HxbfeDFNa29jDVMdECd+GP7yFbSiiZ7Mqr2Vo+QRlYk31O2oK8iCvEhNBr
sq/G/lTZV9N2G8nZapFUA95H/4MrrMMLYsOrwGqNxJXhTE8SYWm+RBt4IZQ9YdQA
qMs2PSq+vevTC4aCiReSHuVHQyRAH9Qa9+YB4rZFTTn7r8QwhFi11T98tByrU5kG
9uY7lEwwMd7QGqt8FrmrZoJV4Z6aAJAYyHSuiIdn9j/LcFL0vRR2A7GxIHYTgFRw
tuJUxSxUC3HiG1hEjPXY6srIIjAxhfYJSb5FXkrA3oC5LfXiILDd/pf7aVfMQ6KU
zOf5vzsJqOafjJzDV7o4At5J/NhBxEGKA+IA0LEi7C4LkF91NtnVc/teOZSA063c
GGEtHQJyoR07oDbxrftgyoSfM1WFQ82OtPdMFnNvUGVMSwbPGZVK9Zdlfd/9Pnj6
8acjxgbR6shUDmPHP6l31xIza6/pvyVRhRqAKCwim/rVi+YjLgw1nCqIcrCYBd29
+hZPhsPwzmmTdNan5/5ldi1gs57/nx/Tl/bVbyjXEKlFP/+DhTKjhTKbPDqRzueA
3bkbGKnLqClQzbxLY8b2VZgGZwLCy8DjPGfoQcZYCwx+UaPCdP0177RPItvR0CS6
+NZbSmMw0BJpZ+pgd0nwxuEA0QVzb2CQyJQ5hUfMCsN9hvan0DZgxX0cd7Iwqxiv
jbfZ/UUv+9WK0rWN0YItdzDTJ7GEC+9gVGdpTa6X9FVWgV/HY/Hn1S69up9PlRa9
DFkV0s9OQU23SxkmHDN1vngt6922FuxaCil8sMg5keivM6iL4Nz5vqocyvY4Adp1
2QauZRZ+1HffBEGv5BZ5DdMc5UulNMmtuW9q9mvG4jMOEhYsERpdlQ++CLs4x4j6
VYX5P2eOoxAzCSV9c9yuA+RqbD+dy26dzZ7sGtxmMnr0qlNAnjk2MNGfRBGWqEF7
o79TFNSF7XqjOntypXSReOfxU1aV+rgIQp3r0fBuuWPBg37JhOgOZLxXrCa8ml/W
UwDUF2vRnIWRMCJJjcYUzsW2qM+djSBEOHOSFwP+u8G3QKXK6JF7G77ZGuyn1+tS
mdS29h2OcSfm61MxQbT2vhFLxc0UvMxZBbsW6TrXG+M9Kilq89TyuJWx0pEqc8ik
9oE9aDPoo7BGGOouUzwqObr15gQl2krbdHdN9j6ATibXFWBWYiRdK3BxZYobIvR8
WhFG/mTD6RtXYxa1g07/iUkZU4Pcv+JrG/man+pBchR+kcB7JV5LrpAFYfAuddal
OkhPNpk4kDUVmSWWsGF8ANICdq5wBe2sJSfMgVO0qQ2Cjv6K4sqfXtYD5RjU4i4f
BmSvcvkrUuEizPOjlEvZnChojKXosusTjAU6reap5NmteeyWgkh2sg6NtLYJnyUH
YsJCUsnm9kj4Xy21YoMspyqN8e/YuxFRMMBX5aTiw/YeL/GhL8YCNGeRtDfJiXAX
QZr+2wYS+hEgkOcDUnHi9xgJvdj9og5bRyE5CNLQ4PZtTyDfRrSMfYJtxdjqyYMH
/iB8pd/Te23HoHP5Or/Yl+NSuN4jG42pRVAZR9unHssH1q+JGxcJ0Izgti/usvbK
Aq95qGnWsSb1jdEEMeJSUL1th2C3kQBdcK99pZhnW5Yl0hFIQfEgg29Q1C0ovczW
OwGNMdo9aqOVelqh2XJbkHNXENZlO+CAEr0XlO//WaWRNJDMxF+VcqZ19MCKv8Sf
2xldpGnVPPzaYXOMQXK4jY+6veeDIvenUvjaQVW5kwrG4yQDlzFA/46+Z0Cv1E8R
X63AQJxOqLXYWJbHWXzpM1Vd7lOe37CBdP6AHPLLKlCtH63b37lvQQWSCRwllYtE
LYAJD4Z4bwrJsnwavJxAUbXmCGFbxa5W9kb3tvzDpxS06xK5ie7ZxwZ+l5Kp+mkB
SbS+e7Y+UCn7fbCD4mSBXWrU2PU9VCGScaYo2CoDGnuO9mwtkeQTUVQ0u1T8pJ5r
0N0yECzN4mKQ/RvQlZPIrgBBG6NI94Qt1jc95ljGkIkM3V7UXGIMkC+Q86csaBv+
OxsyO8fVtx2zSfo7NOW0IRFsrH1xtP9is7jvLG8MwnxaUxlwjjF1j/F9S75dU98W
Xwo7n5+Q/kUS/BBQDgLC1bozVrWCS7slQMCWTRl9Ro7hX9Cgk2gopU7nwauPoEOs
gx757XO4fLYTcivQ4qNadKFOU5vO0u0kM3BDNs9Tyu4fO9F0hgXgwspOPJTz5iM0
YsGWl8IrbUzmgY0SBdohQiVq8Zyp3zArtfUyBnW8jLOwe7HKF6ImcW24i2c8jcGU
OJY7C21qAsUdwI3hwhFeVRjFhsIEGrczDuTUkdx4TCJL4CPVi651gjWwp5vVj/0c
fksvgXKu8WWsMEGDfchqUv6sRKafNygcqeikcO3FtEXgkX+1wBp+HqSd0Ygx2kd3
kvECm6I3ruLTEo3+YdBK0qV9Ci7VPkbFy7DjZoz/joBdJZ3U0XCLOW4HKpN9KQSk
NOKrX+4VPsq27T9BDSfeJWxxuCvecY9ear515TYLBtbqF3wiXErNdFdX2J9SQoXO
UvW74oxJWSWaMvje46+JrjKVO7UYDU3N7qarNFySAiKXD6kvWgOND89r29dQeTsR
8JJk2OscJhQwuMBpqvgBHi5/ddVkf7kwHqQeGytOoY0JnJAytG5p2UlmNlbloBNG
cOkBqANkdboy6K4jc4FoQh5rZhWoZkG3O3Vcu2PXYP3PE4cXABP0pwHq3XF+Pwkw
c7giQhWNuxxQFDsylueA4zK7Beg0I0K7DbHH9XqlcW+W2uNml+CPjXBCHsc7ngjN
/LpSMmymy/z3M5IJkBAzVBthkXdaPj9qCG4kkw6XEWDlsR9P0FBlSZ+A+kb5dmx7
41AwPNM/o12C3iTwvqkJ+mNyH5NZSdedFrlycnDH0go2eBXLL15W7F8vP9AvQUxA
8s5TDuAWmIWxOhAi4jn5FwTGEhrbUYhlqfWGZf6INvQLd4u+3eTX/6fZHQqmQT2N
3aVTr6QFdwmiUN14tniT3a7l0MJ/WZaJyigJfZfw8zXCL9g2m5mc+uff2N/5exIm
LTFmxtYm7XfLl7FAIPhmc4GTaKPF3lzQFD1cfX1jSXU3s7u+CeKCx99ByAvOUdWv
IVlB6pLDItJZ6+ToGhHM+gr0/4Cpt0tCFhMrUpDT9eaB1yR8zSRFwTURojzeAMtW
2T5igey/41L2n8j5+Gh+5TEafc7jLfxea3/YSPpic2zvaBP8S56B5Lt+ypcJ0neo
GyNSoEC7GaJOYM+OC9dPE3uZL7D6X4wjW3OlQ4V0Q/MhTU0/+0rQwqH4DiB210+b
UHStOJzm281KyBniSna2bc+wsr+i22Mh2Iq1V0+/2opL76IrZcUnfv55E5VuhgWD
aJ8fwexlnamkbkJEmB+16ItEYMPVmSUugxAKYyw6/b9zHNyMEnxWK46SgzZMCkNz
yS9BubZ/mnbq3qZGWYt0Ud/m8VU0e7HMipp3MXd8sm3oGTzOsWR1Tp7jU6AUyGZn
vd65yZJLUHiJS0w3esmTAJWigaTgK7Ofk7jJLv5SVBJvpAP+mft6vy2AwSZj3j8m
e4XRgbwCsQCaW6nWs7g5b4q8XmEYhe9o4GOQV0ml4MaJukdoB3W5mh3Q481L5ZXZ
twdpt4ditheVGh0hhT6VO1BD+iZHLm1eA3rKKPhox5fqyew9gWlg6pz3OuVT6p0p
fUQYzM+ucBHJDRfyHAFbNUVwfKvBoGzGw/5E/xIIcZnsk8cIBKRHh46dPJpQ8Jrh
0BFMiWARqdJMxMbLPV1tXlEjWzvQ3pnClrtRE3LeF019vDB5WAbsLzUDgqAaD7JZ
qQv4QdLZ7AB6L8bY4OyAQaEKpwXPSa6u69xERTjcInjJjkGhYz+lJogZC+XSi+Lu
dJAi6J41JfTZbIyi7XZyb4x28XQcAHcadzk0+8Qye1zYgQaYZlr8RDSD0Q3iDAaP
VRJmMq5O5qzWWs7wYErQ50UngL9FS4Mru+P/m6jC6WaYXAjySyqeTaStLAR+RTtb
is0LRtY0TAAsIQPGvHRlm97uHsnSfNslUVNsJUal6UX/SZSPEiKBJQGP93Dlexdo
XNAI19rbjTAww9s5zycbZvazzwZF4j4MagUvFR2zDVPTp+/grzaV2xrwGfyYyjON
XAjJtBn/iCm1AQQx850TTJeictxVPnurU1rOH/UPUZSGqb+qAhZnETbxqIFeL7WC
CFHAGwVr8BUH7XeHDN7cyeGndqQ9mjG3Uu/LySz4ouIbo3+kkHDsWg/1cW8wocyj
M8CQb15TyjgWnVd0JXI2Dlc/TCFDhN0T2XSgUccaHXWBhGRCkeb0iqybz+oWPUIi
gatYU4ipt+2u8uJB8HXHQnV5u9ffXK6omOclSQVIzm9tqa9nCEj7CSrDpcXm9Zs8
4ssBQY75WfoIgZ3zl5UK4JUD9rLu3ABcZ9kaoSzLqBoKIwMfKnqIzLmOKzK0KhCy
vXHeLjDjtiJAP9+i37XqkfDnc1KW5LDksiaeCG9KNFuXaJoecDG2azE8K3ZakzDD
daeFu6I31b+jaeMakmR6DDCZfCTHXuHi3cgg1x5SsZda44ns5/tOk+/bUI3ycFw7
eCJ8EfrC/XwAaejbk+fSYLhHdDH9oDLKAVFsianzASqKDs6RHua6rFctujDImZHM
JmFQgoJiZy4DShUPaO4+gZPjGS45ZFUb4xGwUvL+uvzMNu5HO+lRSIg16NrzZ2gE
08md5tW6wwluRFhXLCw6WGvdkCdZPqafrERa1U7T90lHnzQmShH8Lf4pWjG6w5lw
l/G8iFzuyDIk0urAP7HpbpkPaxFI6bVlmRR9vVfRScl8BNuj06UrwtRGIhIMsGrI
wsSPyyfFlIj7GBbN/XLUH5tPmMqTpAh36D/ERMKnsikZqAjcuLpTlw4wJRQR+FDo
z52xSkgyvK9raa0KRnUsLSdQnQ2nG8KXfR8ttzK12qO1NDri33FfFkId89WQIRaF
3AM7pHc7EXFGdpok23INUuN5JdKeiOQwWo4AMtmzhtgwGod5L2TtZtkPDzW7ABZ/
AKndS3QiaTwHyBRiyag2ZVXV3BUSwaa5GTtZcZeBjKYVuZ5T4eBeZHbMqyp6NZmW
CLxIU8zfxo+b1kJm7e0Up5GSIM2KM49tLTRsh/+6dQ1lBS8NKHVu/TSF8lmK/JVV
xBCaPdY36+UAVs+OKuEZ11ur9qldHfGufELtV8v162R+jyPvWUqQ7PGIxu5YxSg3
umbc+ZvIir83n3MoRB5QPgkU1ahs+mjt3aCGErDdH+HXIbufBmPCQJgd5JeHtZjp
CeEpsu7tspRNd6tCvQ9KK5op/vMANvxflVvMmaOXp4s1ht56WUrLuZ/aZ0mIL05K
EKDhGkUUNT7rBrPdHsEmWsl5afR7pbQVEn09a7PMHBImEFAvep6/RtmMpxPcaZpl
JXGR6+gd3cwoQe5ExjRF4rB/ZhTkpJrFNJInUnHzmJSbBSCE3MKd2U0Zv6Ip+jS4
Ox7L/i/2DRMlTHhat0oEQIxrkLdp863aD4Jr1VtvzWUkWZfyotEtR+9BX6jrf7Id
uKjHI+XjmcZxpoXIPgbLT9dUF+cfko8OmNE++PHMhe+T1XzPv3eIN/IFG5m92yop
/TOXgUFARxpnb3lDpB1UdCe2lwivdRv4TFmtr76b3OZCzoAloWduqhxnnZQn2UZ/
D3D8CeSCaRJLuX3PH7est9N3zAMLqS9rBCojeiQB9m7GKVVsIPYOWHVInXwLyHYP
Ie29KqnqpWW/CmmOYnWhXk9oadKovAJ4DGnASZKlncGlePS8wNP334Uds+8+OSwz
PF/8cTRcYhYQsELzNqBqT4QuqaWSxdwFE0f3xEFdJ/3lI5qJu7YpmlSbp/jRQxQ+
Hy1fsAPoQ58gQdK/aHeJQIq0fXPy5SRiCvxft5wwX6Us+QisE2c1VbBnJhwzUpRL
bVmMZ8Gx0LgFCnINFiPk1BErXh6pXwk6/PCr83tDktZss4S9gAbLa6odsVdi5fQL
wdJA7b3e+4pyjRBuPWnnZfrbEyQfKBHYNm+TlYa9Oxft29rjGoeNTD5stSJXXaC2
ppGY5DHP54leI8O44ietwZJT0/OKLN1jnCH+mPAmPBWKUx1QAp4EW5xI8ngkCV37
0sEmhg+4K2SjYnbCrUEio4cx7rWPH2vGFJoZtfz+Masl/zxFhwkbIAiyicmm4DOn
J2DCQ685jv/wcyx5pG8z+3R12cnI/4Ok/Xw7iTS7KMGavoW7bnnmnQMPEuiAitWw
JkcuhQdBExnWH+jq/1hkQK6NmLEgY5KZCl/SGpurEmL3gY5se8hk2N78yqRR8dFw
lrCq35m6xphZiYw/QSTTXJMVEFDeWk7ntELupglbTrlPgQuk4+g8NGdBN7UsX4MW
4xD4wtpLwgON69KgI4X4ZQYJTgWlR7jqXy4xkFl88jXW51MKt5ZyvXRdlo2GxkJo
RdwpL10fcOJ1bfnmMHuKdAr/woymY01T+G1UZ2yhRMNmGKVjzcC810OE4mejVzxB
JoJwgKr35ICMo6+IK5gSYRZqqdFFgjNJ4nUXQX/hdswQWwm/3XFY36OHIkAlOVfx
ugjm/hbF8Llm8nerfOxAfCyw9KPJ8pwjXH9R46KLf94xUsMe1MDy8AY+c4IXGOU+
csMDo0bExzFUvgG0w7+NbsBRslaCdDcf8/+Y1Z5idX4IUyicvrc29BqPqyjFMCMW
j9cfV43spad9RSma+f0ixZxWDDWxqIAVsde/zORxQNrazlbEOqq/SUI0c+G4Ihw0
fD9U4f3VZyYw9N8NTYGNwIJivXuHZaR/NewEMFtGotFdq5OXGvm2yxzaq+naoeut
6OZAWiYjvrctqvsZlggwbJCzdf4eAoK1L7Yrp3I2e3f/ipjmf+W6krGPWEalqYph
/oWPzsPrOmroF467sz1FQNhFIlftNbPA8i00t/ZsoGWZDbYWkH9wZSlDHkcrEciu
dExvJiv+32B/sJtzswYviwhBkxpu5HthGfRZi3DTN0/ZqF8d2WQNEkp75aYHdhGD
lLwQ9z1tF3XZC6dzsLxphBT6Uv5aStafHNr1q3b8NBvqXmLw/yyhlpPRczWhEVLj
UtmhoJtST+6LxHIt3ydD9FoOPUoEkROiNQuJEP5LQLR8tmq8g5guvlU+46/GonLZ
FgJhP21AJKQKfVTNJY7V/B8NdIk8soVDnCIKa1yjauZNOk7g9uS3VwaNZIVkkB+J
pM6X5PtM1crnCfqEvFeQZujkHaIgPz0x9Oedy0/3fub2x0+H85wCxw4lCTPVi3bq
HAA4xaU/34mqcBxSyJdDrF6nksBUk7HEmQEEHMW0LkXxr0l1qHetxZyBfiIlKGAU
y+b6hymStqEFoHP2Ro4H2zrhz1srkSZoC2zKNjHr82Tb/HG4L4J/eXQNec1M93ld
HXMW2KuFC/RmixkBVv/USjX21KyvvxadE+IDidOil4NcnEI+QJM5ecHZ+Ul7ozhh
OXsKYjiYXzIES6/81322/Q5l/bxP5jZunFYp9nY0MWByJ7+Qp5PqXbwtvFB9+Tmy
nPrjOSEOf7Ed13r/hZra07Y79oliZFLju1BgGOtNqNA48EKqK5HjiD7KF06/IBpq
pXhkAHPFYyUcL1u2B79aKhin4fARfHUDzLsWvd09r86rCf494QKPFc+w+oED1xdN
bHgcyZfgPo0KFphYVZdD/0+YwfJfIoxXfAdAn/n+UEC4Fdo8OED7+nwvyKQd8MOl
hH8bLzygCHlcNvFrNeQHSqaH7XYaP3Hr1xJxydvWjvznHzGMR7zTNnworQ6GltJc
5Yrrt0TjC2xYvcRzX7VG5CikuHNIZ+8HiUC4LnM5ioCjIIVE2s59c/rqkaYKmYka
017JP4LoUYtJ29PA7EE0YtlqjsMGJ7smogySR/qLm54pHo55teKVMRd9aTPdj32K
f/wPMZXbSsuDo2PKfO3BTZf8491IkPG3jSt45KVZABriiIOV/1H3lvZ8qKuyXCIk
u90uWAmpEhtLk/Hth3LPcQDm/4ZolG8EXLdoJ9MIRbMx/o6lA3PfXVSOQLZRayhY
awy6pXDMkEOlns8O9rbCPwH80z2dz+7J5v2r/UyCEvEU8QrHnB4xLxrwoL8SxHGP
UAihg4+tlFN8kmSZSa3iebI8nAafPrDGimw1UAEcLOx2H4H502LI2kIKXjYnkGt6
bDYDHyu8oMkSikDrM0RzLoxP9kHRdXJOCP0nGlDj3MLamMLXsc2w0/bfFtlYLBX7
yy5Eq8mlTMAGIlnZP8CGV9b840AIcjPq2K8nv28w44NSjNQMhN772DesuQhCF2UD
ePSRp2005LOh4YednB4HfzrXEsauLoB6wMecEb5zlhHBSdbTE4+oj1f55A1OYXul
vaoubmekUN+7dMACqjhp9JFgg46dIese9M3T2plowL5OnpQtJqn1gpy5TScq3EIp
5bz81iO7PRaSW1Btnyo3FFfee8/kVhstMBPv9OWZ8scRR5AsOw97Ku1ViYfBszT9
raYsTnJ1TcfCcaRwDiyOg5wJkl5MmmbplFbEBGMHb1IuA75bRPeb9PMX0Qe7yI07
iILso7pbvfvb/YrWVXJvrr1Xjlhv/OiyF8KLukqDH5fGVHwV/Qnd6hSDsFag8odM
Xea2ZhEj2Abf00E1ul/UZVcXCtig2wzUqhPilkLRF2qbOefTWd0CDepSgkkVIN0f
2duFPaQRVizqVfoHXnk9rAbewcyAEQN+gpzyt1LiHzsWoYZEmH/PZW+e51WCQATN
eZKluaGHYfzWq4NeJBjBD0ItbeUPaCKXkEDUqqWMCbgr7Sk2t+D+ZOxveOThglaH
e9ZxAEDow+Jh74B17YoUNh7IQmF6pvgEZYhZCQVzWO6fHNEFhGrOb1kKeMSghTkP
Kc+ZRwZbicrlUwBA8H9qsDJta/9FkOK3xXCY5rHvasMa/r7rWMfS9vnL1+ve+EY3
fNY9K44roAu85w7iId8Qqo2PAT1ZGwGKboBt32I1wl1ePNR3oalBtKoD6FHZcYVG
WvBdkiKk7xl9IPNhEShj/Q/1J5kI4asV8p9nGMkWN/ucndQhSsIusObDjtq7FdcJ
DYF09fyEpVB/1P3pCkYhTyuHQ005XMgRbOb1i7UsFzPKb6/nPI/NQKksGtA0JKsn
kVTs3VIGrAMZzMnc/ko5FCDx1ErhqJ+SsgnWc1bsLrZ8gCSg5TaLTAfYAQEcdsHq
6iIAAfqtjtWMc5oiO2UDCNyw4LnEO+uqv5XrIijfG3vFuR8WroKiiyyffSx83yLO
b22NYdCIPD6Oft+5b3WlCI7IgU0jLiaZhUEKtvxnVzJ1Sh7W/F5Tah9S5siWfeTz
8mYY3I+9j4K6mhWL6ZD8kYwZe3HNjwD8cp99SLv4sN4K+Ibf89q8CIXyv4IwJCKF
S7Lvjq4ZVop+6precBFcjkBw/fOM7MQmowsJAGb833PwSkslIK+CLWz1pBylJBtQ
vbykQdYc9QjqP23kPq+etC/xGhC7oQbFf1tQwOl9V4qxtrWIO0+qHL7p6L2xEenO
sCkCmqUcPcGu+NsczAadUA/BOQmA5ds/uvk2wraGB5ZpzWoFBpd9dQd+w+w3aneC
y/U0j+3e8D4IWo8TiPBmcb0LPf3hzqXNg0HK6AIeNAWGrnWdm4QyfKbPSvGwzZyY
rFQxkp2Cx+YJvvPng9jqjnBUsQjaNrHtYqWBuVvwzzy8qe3CYG+nZ2ovALVN4ZPX
YPfbyXPwfGKbvaTi6zI2mR0/+tpfzVSpytLR0SGTw5D33AztuCJ5lA/H7lvJBYf1
zY7EPohd3draSopKddVIdIo1hXZ3QWL/r7GhGJMycbwTSwlRUjOlMF6QwDZtVfJj
5Lmw0l5kyDS1o0Q+KK6J2cJeaYw/7Hks+5rBiVUkihJqWUEY/USnsj2WXpGQkbCb
DXuRtW5bS6Ngvq37T3VsmgBNZy8lk9miUZiKDYhpkRQZ/6VlsXpIbbOpjIkU1VwD
LxAWXCrW3A+ZMOH44T7Eg6edkHI/j0g/0psmAFH6XOWSJppoSvbpawmSfK8a7eC2
/lACHRsWkyG0vUqKnnfAYTHYtZmhVGT3hOosFUoact0zoosvo804/tliBgopNEda
gJ6icW8xg1ZEje3ZcLQVMrKVb3sxubzPaUT3/kSvvtaFbvUegHeEJ7kTAZx/rPYM
wT66HWW5w59NLZCT8+9JxtAO8mn3w47mNgDGN67GS5iRN0vP+LfEsOqzedUHNmjP
Z38ZAqCWhqKWVgMjshca7VnYpn6kRVDWd2xiquHp49QSl8pj+DmiftxI3rt9Gwvt
xJcA9H9inmU0A3Lvu8O0LPeWCoiNTY6KuP4oVtA03bD0BBD+1aGSvb1/GH8n1ZNt
/hMkQZjXZ++D100LIN8eTBQNxhD4Oj5lCIWQawEn8ASzbyTl8O0j9y8cMQHfPHvx
npdqi+2xauXBDoYfmlq3RPCttC3+BeNYMSbKnv9fKHBTqrakiNc3ya7S4iRZKeyY
DiB3CMXo5nZRudv1QyiYzIZgOgG8Vp5BJ/ljEuWMS4cxZhDumORjVX0SSdKdULmI
YALmjQWVigi9YEgJM0dCmLFLQ4u/D7ugrWO/CA+uMUYOty779+KlPG3fXD2MNbgU
PXEqY8duPZFosVpZArjWc2hvFqbO9EOA0Z+UnTTeVibiCrE2UUeOmfjxOmLO+C/H
OfNiCHsZv/Tp4d0mVZ5KeSEpD6OlAqFiIav9pHzS6/1u3J9wxOoF/b5VKuxznfRE
qEk3bhvYnyOF3vtmRrjeEFjQsF18XEj4LmVclNWYfd1wsuM27VGa0l/paRrWa+4t
nqorYeJnRlEEadocH7AduC+deXDf02H18PIRfIFnCtiuV6dNpkX3tL66vGGxG+uf
Gj9RgE/3YIoBgGeHYm/ZgMFAw6XM0QiVY/xBoQ9KTHhlSCHzLlBxhPYo1Ru9LkkR
jIb1enD7qAMN+uIE094JXje7SuZpvVxdDTINzwkqZqD1iGO5KadTS9iqs9ZpCF6K
anqSzviaw6/afOgOVUMn02jrBOsaqItrJjz2Fzed19NuvyIJMwP9Yjy4mjZrdklO
1sRQder1NPbhU938IxUtufzi0Dt4qaqSXmFC9wo7+hE4CW17LqXWGnHjqZIbBdKM
qchLQ/2YfDj1Naa+x7RuZxbEnYjCpzeW7VjzXotsI1nmK4HMpJ3qv3BWhPYLqFjw
LSrntF/Dv7f0GQT4gACio5Y3HJO3h6ApjI+xM0IOj1O1InhJ7qNM9sBB8up4pQqL
ZjdYRwGc/AsR9UaZtMVt7H4+GCNkDbvJyLOlsvMnuH0XCdrWCOaIA5FEu6OzHnu0
Dp/UbyWeSY2BD6fLhww7k48XQlV9rBwKOjGDWjePV2fWYMGVZAirdwbnYlGJyluX
t0H6zrx85Dw46EjgNiRSYadXiorXX4ssvqBvFLckJsXwQhy5gp7g+w5gKYvdriS+
RWFPx4vW3ks32tCHIb4/6tVqVwGwg0NuRXFLE/1YPoPg77FmK6+mS8ygUyqvR3cz
hQBlfstqOf9g36Aj4y/rEWBWUBt3CEgJxtkDqH04hhnC4mg5goHR7r+m3jDwr4wr
l9u0H1yK7mVRA4nRp1KdK/7c+3AF8rq1c9Iy/TUg3JMRU3YVcHYo8LgO4sX4VJyj
Ghm7LLy8zEBBZPCh0zuTFDa+ahjrK5piuQIdPYyMaAK930xZp5vh8aWpnHmdQzxr
sKNzff2JG/tBHv+AH5Qrhlux/A8ZnejRzYUjcstWBQsUrVOtFchOWg00PObYVILb
4YyOP5QAOiXxTLAXUkLf641i1c3rQvgGJPyFeJqNM1KWRNPyXBI3b18jKg3N6pLf
W9Xz2GIsPK+4f4QIqrQFQLdpmKkWC47eR/bUlUjkZ3e5hFN+LsmebUqE2EYXcRzA
5ypDAtMzvE0Z8nGDT3+C6m4qarCHqn2OCkpDTaE0NLozD8VsJfRE/EZRaL3WFKcm
IkpIK6IrVGeNqAzFGnz3zaxtUfPj+WUCTj0WFY7FBzyQmq8JqA79PEiIZfmk80jk
x7he6+6qexpB4hJyGpiDtjamETleQslZJoSzJS20hvfjSkdK+4CS6D6X5LfM6RFf
w99OfPY876BmgpL3gDRi7aOBa6hZHDliyTCdDdexYdlpyOD5btZtRFZ/VnnoRb6b
/pJls6Ml1bdLpJEmx6Cj+Vl7572TwRqQ2w90kVONdFarxSSDgR6hNnltrRwuLbNp
pR8IcenZjPiV57LmerF/BnaYCY3C3lE/cEhOxXeE1nTdDRnSDPbRq6enS8K4xYiY
xyELnUtvJD6loepLiO3RFtHcpS/TOd0f8I76lFmGEsREBF+bLkmI1ZrS52ulJdOp
zyio8mi7wswYzg+SjHPDksGjDlPF3ZLhfJCn0liunIj+cq0+CB9Q8GOtyA3gWH1b
o37o5JTl1zkfaToVgg9VXyOJGmB94DX/k2S6gWtdi9YTNCi5oT23N9zZQTygy+gC
reRo3/+Wjqbnu6/gCcz6cM+oo4nFlbdkH9rH/KqzNhyKbrip7f+6pOBvSEUgd+Z7
Vb/82jPJdc4VgrgTh2Lb0IyL2rXRbxnAq6hYsggkNij7/lB8lXazOX8LmSaqEwSl
arVt4lCWZ4Wa7rCh+aL2p3laEwP/aG4AIYueM5vT+KNm6X3a7LpCFeqoINIV2Htn
4h3bEwe2L1Q4PzIFhIEXdsyZ/pN2IbWS/HQJ00uXrz84fPCBDTsLDS9nKVCrNd1R
8I80brhVHsvptsXBdwe8fitkv7Lc6WSb+sG3aaUnHmofHn8Z2GpUPclOlSRGMX6z
CYxDpj5HqL8oWtO0SEC0xa9ZuxrzB4i5xKGPYsMjVYI3xlwWQ/OLG6MnljbhnghY
inijxtaTFlkIuZacihp1CS4pMu4eoh+NAJ57pQiMiCQeTjGYqKTr6pck2Wx2Z5mU
9opPb2kA36faAGqv3Bia9ML5sH+rKu3/CX6X/WPxKwpZqV/K8CjXR5owmfY+VTcl
9rK+NJa3GKmBOulvYQntRe5NcPN2v5I8xW3pEwmoERRVgfP2XEMwbOeanas5KKL8
EaTwm35Ju9WARrNcVZIZ3QM+6cftle6g8MzS6fjKqekdVHwhL/DptQFRF0I0+MXm
75Tz4TfPwOb0ZB99xyVtAN5xh2zy15uAzH8DynJkWy047IEm5Az1+0i18jENu3gW
NRuH9S8vY93QJlnmM8B3u4nsHGUrkD7FzSEZQnqOIHOGvwZJVoOpc8vnQxbcdfSA
OyIKy+SUAs2fojHqmf5KsjPfWGKetfzkVA4xZHXm6M2pti+brcPvp+eZ2QCQQ3Es
eeDB/pxuCr1bpozQGEX9rn56kViCwmyjnsOg0zNgOxnJenLPnyqUEVoK+5dstvYH
B3PLDujvnXVseF4OzXygUmzwixepWqekKkfRqfOxB6DLYo/67nx5u24IF0SJXWUY
xX8dQsoGKdM/NmKyfU5UpVubWIdYxDMbPe5DEfUWEd0BqziUhNaYdyQ80PSALJYs
Up1RDqN97xnyMJPerFz/+smsiBBVcJjrVhHOa15Cxl8qQB4pcI0N/mwt7ZsmHBxt
eXxkJxaDxAYAGaEy9Iiz7tiz5lk9qmzznkVkcdBLPRDrJDifMz2NVfQY995lS4LH
v83KklBZBHTM8H1mReiE34RqJKbFcxsc5UILn/mV6foT4wLxvorvOlBlJgbU5xhn
jlWi3MAeWan7xXTncYV+KRbe9xKF+PK96zJM3GSBen09VzXWaujYbUeFS5W457Fk
9JeDl5zJFr2IRvuHH7pKJ1s5pFyDBnvvzdNZQk1li06DJUTX5G1Gc5KruzRwJtB4
5nNeyNISYtIZ6K+RByBPlPOAvbxQP+uZj7nH6eMlWLGTDnoyonZbZKuaBgTDz0hz
6SPRBpOnJwLlVRtcslmXk/hCA2vRqelDWT0yxRziJgeEtrd0zoLF7A4FjymBTu0F
oz6XgzsGYUMZP26q7C4UbFkxpZn1LUHPSXgcK0+lbGqkTUuHL1V29extiyC/NUHb
anUqA6m1w1Xmi0HMSMITQmb+PypDqQxgQ7kAxuUEGkGJ0K0kg2Ey4mndNtgCJw9S
3W2drZwdqz/wfZ64q6hUfJv39KtadvlWBAXlUNpgaHP43N6kWkMefVk+8g4Z7O0I
KcASW09iTvu+lpjSbSzvnKuwwJGoEmZ8bIZ4SCGx8VONcap6TOHMZs70pQ0PPz6Q
bEq0IfkJaCbfqYtjeSbQsMHBnagSYnefxUU5ksr8mUE0TNQePaLTgxKDTmZc16PZ
006Y3YMqCp4vko/m44j8qXTLPjhNXxp/sN0VCb6dZkcP93GOaQFw55H3Zlp/yMem
UmTqFCAZqd2UrLTpFSk3J8/p73WY3EUpMMl1y5j78pnOCSe/nIHVwF9nSJ9n02cL
odZwOcU2Rv3NHXMmupvRUUC2yUq2doaigTK7dHlbjTAHg/TJUG1NsQvfmp8s8foZ
apVbDEtfPckFO7IcDizt4D6sPeXeq9/T6pMjGzp5BfGM6/CuPpYjF7y0tGw4VeSo
euYUjDEb9h+lGjaHARuUgH/n0KCxUhGcT9ckHPW99rO14ZUFUyDapcfQ8ipRFNlF
nVZpXXrEQIZw2subXmsSp1GciiLjNpZYm60VYM8p1q3oobRGcwmU4QrLC4DzV5L7
s9pHqfDas4KCyjK9b325EhamfJPHUI22n+XGID4vOB3zGMYZASYCSNS2N2vh2ivl
2+s4axBzFL7lECG7Sd2UKnls58deWG3LDx5eKNTYD7VEi0wq9hIplNx1OtmHPgwK
mJcgucdg8FeEOG52/bMzsxs6jQeOaTvRsu184v0BjmUs0L25drYxaQAadJ3NwsPW
rl7ACJUwRaLFoO1vckbyVu/nL8a6nx6a0NfvDmDgXgoJ99eDtZhtDtTMvFNxkvwf
4+mVBI1g5Co1VgHjhuriI56G9m9o5MNJRyV8YJIs94yeir3pvLH28aSeqlNwN7vy
mUznQmyhM5Ob9Sr7TK+wIj7DlbfQS/AjY0aX7M3FpMYc+kMF1d9Dq5VlUBL0RDrw
uj02cq6tvEUckfm9T3EIBWAx/dwmM9ai01nnC9OMO+ENPg5SlmEaomY8yGh8p6TA
g9F6TivK+8K+2fDNvYTUiWrapExWKWvoEIe2qPDiE+V0I+pBQfYfm6p2tx9fVn+J
4O9gt51ZQGXLz1TUvcXMAbYxzizpZJWavCjxL3aZVQRcoYjju/TbpsYMLmZK/CFy
XJLsNb4rC4fMZHVru7EfUFmd2HBoee2xq5RvpOEXiGKAUJCpBwmNQFrh5gY6yBr2
WNy/BexMaZ9UyABJl708an5dUlTQ0mg/A8qMZJoH0MP4+9HAduLHnlSquV9SvfSK
iMp739LuVqLcaQq8FOHoRRWkkdmzl31SVyfEKVUx/4zxiBWZavZM98P4vIP7IqI2
vH/gLY8tGwGvhwfNPNPdS7J8zRoZ6C/jwbpKC78l37fprmBdSq1LeFkhca/Uh+gj
sUQL1hAZvMrFo6opBulmbBoyCGvua4/qvBaQjxDC5VddXou62MjPGGUlCAyz24U3
K4/haInvhHH9k9z1inATc6Wm5XpfMobYgcV7nDf/8WTmUks+AQyEO2MXDB08ew5S
asyH5DyqYSneH3vHVTbr8Hdncx7X5aD/u5ZJ4/fTEylW7xilINGoHSiznWeJdjMQ
+juzU2H3FbEi8F2meM51bPvI0gBmJUwpiCmLIHXpYqc/0SGkJhCgV6jU+QFqzy9t
NrqJtKsBn1sjt/ZJZUMGgqNqqLP3698rb/uKecN/sonQpypDafh9/t38fVPny7uI
dDjoPQtr+9czbzrEqi8kMKIE+RN30Ipp/nkeqHcogiHdxYg2GhpgDSIKTwEyHxIW
zWdurOyCjO7D8cPb4+xbTMJdZVwbev9Mw3/L1ofl7Uj9KF+VtM7xgnVWYCxjMrTr
IfO6r0pPlFELItnbpyB+ej0YX3F1sb0JSVuSBa5dAxNPIPx1KFNsoSitJpS3DhIt
Hc82HQIUkXyDhjW077OGV8jaPPOu3imgxbu0ZfB3Uhn2tK1LtjJvd3+i//DQYwX0
//Pn9iub1WpiqA2VHJ02SwRcFWGxV8/erUeLHeFGOjwbe8I0dNUzzA41eeylLIkm
BZgQC936dOQEQq1D+i/x+PsN5iid/66f4vTyyqN8TOuiK9t9zohiEJwU7u/EcPwt
AqWaITPeVkvQ3dOnfhukypnpSzq2XIpkczqJuUDvsz4nlTHZ9qXLu1Dze3mAHsQX
NKttki1VKeEjz0+OTf/2QdLNMGNIXpZ56zF2C5qCDug7zOjNlIGN0BAYJ0XUnv6A
aZMehUMqDEW6fFt2MlHmmptkjMVqMGkmdrVQhvZkZsIUHyxk8Yym5ZwdNdqC+KOs
X+jH0o3SBbTZvNu8ML9shcnouZ+JBULsZZBz0ppiim/sJdBlpKLovdj2SsNaWO45
xQPnfSUiw7KCWD9CFvEvT9sTWOXPQs4v6ciZYQ+s9kkzd5o+CpqAJwSyNh4+fPiA
WyPKbe4Or+Ou2e6Z40b8g3MB7HPuW244OOm93x2fKz8LWSY47beXe8l8Fxff0L61
IboHkl8+Irbz79ww6PcUi2fcdcpUnVig3oFmkNj1FY+0q3Ee/fEXrYUpZVZFxLcH
oOI/YFNkHceLxpbfYqM6FAVVFDFWc7LxZ/DAtGOlkftSGx1jO+5rWY8bDr5ZlzM7
TcTnk3dUhDXPRmlWtLSSvGKTVWWt8Uj6MEq7FUDRXDG+Fzv+dcN/A0tNP0exCNXM
SYELI2lcAMBpbIvR/eo0JGN39JyRSHp79DsSjCzzbzLXX3pHdRKNaxclupa+4ww3
YA2N7/evp0fZo3DxLEcuE272/SnBnlfrFk/b2LppuK7uKVd0/V3WIuyiNCIyJiAM
W80AHBodViB40BaUHIwvIyYy7AZihZ4wCoZNqmlrTk90H4MNmCCncfidkvAGjk+l
h1A0AqI8FYTyqVh+30TY4OfxRuQjcTjgqbXEV6Q0mdYAhvfz/RDpGPcrifa0vxne
D79trH19nPJXn6OBfzBoqyNljEpnSIDS3/03s4Mpi+H7ZY1PGjCs+RWd6vBqJyFj
IG29cwu61eRsczt5nrH7cFXV4SU/bTMrAqFy5tPM4lvhZnepcnIyr44ZH6J8iw23
bYYOT+3r5Gr0gLHpVkfR6V6cQ5lVQbImyBf1moGypFWtAVD44sTSXveW1mur8IOk
P6/dHsPDdlpxdQI8OGuPed4uN6VsrYkZyVPC8eImyOA50eaxTUuYBFabtVwoyqh0
UBCZ30SMW2tr5bwe1zHOtSVGfjgzTI7SuziPgRy8wcXUADpqmsBpwOjlxdEfaZq6
3p85mPIBDMMGmllkE2rS5G+ycogb2KevI4jNOcWlXbdcBf7o55uL/+d0ohoWYQh4
fHl5A+9OyiQkZwcTuOsUmAjxMYgOaOT5eKTwRsEhSlvebSPci1ZaiZQKfk+jSm0j
6pKQ7IiXRS1hyEbgy3DBgsTT8PewHQA6so6IJjOPPntt6eJ7sWe81GFk+rZ3iC2X
Gmgw1NoAnqi+aCGATLYFFpgoiZcYNH/mLNEsnF22wKcD9hZBr8YOZ3ywi+PuQuil
LKLIxBELdmAnBabY4DOrT94uPBENDqV7aX2++V9uGrez2vkPEzZhOyb7clAI8sQj
wqEnBoQIMYCy87nTIAaJFDOQQHKk6fU0BrfmJqPaATjvDV84k/vmIE0+z6OR5kVY
cwlJ1MpRwEptLhDECPVBYbX7syRhsW8qC6qkQLerI2+HKZw6rttTRf3LULK0wOSq
LUx3KQoE+sxGMQ4WPGy24+nNIZauACHPd8lWzwoQSLGXAIVEhqBPj3sHZRtnCW+j
RMwGlsnVF91Xc6qnY1L/n7A7a5NUChJySuD3NT4LqgN7/65oVD0+IQivAwdDeJ4a
ZGPY8Deorcq3VxtSmWE+F52H7cgYnmqYp4XtS/AS6SQhGrwVHv5K1ynTvfNW0fd2
sypT17/+eaM9sY55QZy6/dMsMLA47w9kMWLSevOvFOpe6GqplWhlDnNwfC/P3yTZ
xLAWD0UYuffb687J5L03Yi4drcw8QXDsgu7vUyj9AFkIGvDyJozfCo7tgmRBxJ3p
V7CZvJtH8KarP/9giwfLuWn0X/UDnP+kfdenxDvBb4HbHWLen5JN9cltfLeRC1T+
aKi+DktSKFMrf7PhNfYZXaPmaQPdgAaKrl/xsg792z1xp2ukxTHYvAgf8uUNmCb0
6aIrFkAy40ZQTCUL26W972uqO9/Dyl2s2m4S3Te7CUWMKWlUBgtlvjYVwMWM0K9q
8jFq4i6fs9goy9I37UVlvGlHY7qkHVfZlmAQQLUu5dtZE1RDAoewTPVwk1xZnJbL
BIPQc8CclrbIOLRqACFg+uQuc5QUc/bfQKBZ94lnwA5GNBL295nTOqhwU0eu+2vt
hNzq5YpBSRy30pA1YF1CS4emyfZUgXbtUXuEDIp6cW32uIEHRTtli7oNMnw+RQTs
gdbTbVbm6tEY9ZpMJ4LCu69+rPIPCF3N1EPqLPDtDANB+mbAtK3cJsuApFroigsH
q/Fzto5Qp+glrQfj6OG90vtInhqU8y1Wb3fjHm2pSfgg/ZTMgz20hDmcldMxMOgG
CPFDNTdaAATtTnVenxNuFVwq6HRXy5HeN1HNfzkIPS0ZLAVUYpeP5eDP2Ummrgur
kiTKugaZ2NCIBl01GHpC7CMB4RrECaUUNKsWxvyM8g8Cc+FRfrn77g9iNrzXo3vu
2vCw3ToYLcBcpoyqJ1niUENquDCzt7bjPWrzjIZ+8MNA3sHScpTi+nLc/1OX2wIf
197w5wKLrecBE0kvp8g4Hz+WPcNGiWQnGEM2zir6pFVQqpKybhSiOUfANZjmw/QW
EzKupjvWLsXcbecuFdWyKzGo0vWH2ot3dnp3XWI7Iz8dCS8oZnSCoBa3uwrl1WeP
kPHtAAoUNf1y05vxOh2LZMU1fcXAILOjzh8eoJmDg8ES1N0nwkGl6rr6A2gRWtbm
1Z+IsltQYxE7oSRhc/yvfYET1q1TBDJC6/4RJ5yEJVKLzB9Sp7QfOBjq4rJuX5hv
b/bFBSqLyNt8E191AnvJN/x1CTScIQuPN53qnzRYH0S9btX5LAJ4ix+JRbYrK/qf
9wAP+HatnIJ4VpzQbE4LlHIalqlsF0Db1Ej55a6RpcURsVwh040Li0vtH+376HfI
5cD1E2z3bDBtLw4UOhCrV5Auvej/8ZxjK2+zp42qxIjq1AgaNkJvUgEuPW3BfrYD
vqfyLICT/gVEqlykV/7QPLrysoZKZnTA+29FWp3ITcKx2Wxh1xUIopePCjW6NQyt
AGCwghNNe+BDLUC/RDFn5UB0EB1S4UTD0yoHBPhHK3nblP+W9pTPo3+mUdXSUi7P
/MD/4R1x7Jz0R79n1MCQA8rqHYrD+Wq19uZ5zq1crY7NC9V2AHXCoT6I3cZTixbq
U4PPVwxTqv7fZik3GY5V15uXMfcGz94IpmuSwlpPYHlLRIYcVtlbrD66LV4xeeR6
dENjJu7xsYxatro7kQAqH7vj17HI7sD8xF+W+s6X4NPv9P5z4OPSk0Hn4HwNfBw1
J0yq5Bv1YanM0HxzT1OV2WZ9dQvK3nhUYErCc4cAaV8ghwDHoRPghf91Ijo+U+3d
vyP/s5yX6BS77PB1ITn0/ZLd5qW99aiPlU05pII6j25unXhDldgJYPbiw33iHsGE
pjFKR3pnoG2biwuGBmC77g5AoqKEzBTv8JsJNfKmCdYGeKsxF7n9anCGaY+jSpHC
pneuPVkncoqYtAMQZOs8w15NYe3Qgz/vSlD0kA8u/rrN4E+VUmTIglvgiMnDLP1k
0XcNuBPHYUQyTAPJgsmgbzsk4P0dugF0xtIn7B+K83utXL4hapWD4AgqQ9einx6u
dp2kOPzn6pVtgL+zLBfa65k4XTRPKpFL4rbHTyj+nb0+bQCdeYJE3qnMiJgPrFJa
lIN3GchacH7NIVi8jL0xM9/PUj5zdpI+rkqiWuFEddcKy3zUXArOi40r78scRASK
SBl/r8CYzkbZz8IjiLpavEAsN2hj5yavSG3mV60kDf2bEBJb7CippkQPurOp0Oxq
2woXOPNRblyudGvx2YOZsbu20f+aiHUYhMK6oZSNUv5OpWSd7xJlW4cd4Q6w5KMf
hCfk8WOSXssuLndi+NGPEJnvaaBzGKLeKtmUV2/QO0tcpyuaiGny2TT72Ml4rK9Y
SuifIx0zwGlZfRR2U962ft7nHutsq+xTjWRlzxXtNLM1ecShtocN3NiHU0P4GazD
PkKCeIqIxYA9akakJKpPpNQLs6+KBEPAK+Kf/66kCdxfNUPK9H/+vnTTuQGg7MBA
+6X9i5Bv/WQVZ3HoCEIvM7qXanvMZ2sRP/+7mMYzJtTykmokxSYE+uhR/EuLd047
AKf12FF+UhDpIcQI46rS5h4V/bj3XR4mSZbTN8hJzFhE0dIQOmCaOju2fF/mFnMN
Kvip6FYUPpOCE05R9Yu0oDR52lwAGsq0RAr84K6G+Dgrg+vnL7pCjbWNiy/FzA84
3Y9Mt7X4RpFKFhZzMXe+87+mxxXwIaczY4V4FwRv5ZXlwyXqtUPixgtZcWXXYZZj
tRv8u6kb0dusgQX3xVrRzf77Q/aaC2AKA8UavsC/Hs5nG2wGsU8dIg52zQ1dz44Y
Gc7vMMSZ2ycpoGo5Jos1hvvPHBjPJDwT9apPrkMEZC5RkMgk2QneC5dsSzjnK5ra
2ivw8lq8pWq3/aIFWHVgSlDMT0lPdil49pCV4+XvqtP5h80wiqO0KnAiaRG3pRXG
w+/48yXzTZnE6lMcKDhtb4IpwHk17cqLaAgPStGB636RRh/2DsbEjN6SqSyYFwR4
8rULPVbeGmTscOn2oOExGF5P7u358xJxPdbBJdPUmdeMj6TxRamCl/9C9rsGPdnm
8fyHnPQNOlXJDCl9c9eJhBabIoZYAIurO7FPFnfb5mKXX2PUak2qNGxuhSQTTEuW
JN2WE8Fseqe0C2KtEvvECIbbsR0n392+pdFSfUWFPkQrHtI3dSQoxA1lo4aU2lK+
kfkaMAYnIdN6NbmTOIZti8VAMrWYQFrUsq5hlhBtQCtcD+4XtiWjcftEnHBe1OQW
NVN7xDBonTa4VGUTKOQx23I1S9A4YO2niTHpTcflXc4fIWTSpmzYKlooEpEotoAa
8SRICjNVmnAlJ4bMc1Pbrgks56MYUxS0l2THFh7zTTaAi7fKHkoU1Co5L09zCIfU
faw8V0b8gQI5/R2mHD9PsAl4xUE6G4E4s4daV6PaWpXWDoHQcRK+g75QmUopLPDI
Lk76rHyTP3U5L4DSWfLUb+SVhenH+Ayiv5MPiq9zLs17GnsfLbiQ0wyBaiFOwNIz
PQHRqjypnfA6KNFs5dQf+LhYGOoX4nGpQFOYm/rx6TUyryJtmsRKBRahT14JafG3
OEZz+//pg1QVvZY1+CFczNfXzaY2gDr6wgoQwaHP9f+DZZX8Ol6u1s8u/PhW6BL5
atZxiciMBkIa4kcERgX+yvQyoz5MxdyaLAJ9qmp6AWO+5X4fFfcDJXptpIwz9AKD
PQkj3/I0VML9e245eaGyNR8Gmd3OXJIVaGiWH3NiSVVsxQhCkAOQR94sn45BrF3K
nq+Tl6vy71H4FqsyF7KD2BcnZjHBBAzB77GBx9cBy8+Hnm9oiH9YlXsHpvN83BZi
DkW8Z/a4a7FfOvG+fDY9LaynMMoPP/Jj9L1aJ4Bp50xFdJ2IeBZiAKx738b15OPQ
0kuO2IaJzUOByAIHP1QtHNMKXYod/VT52VII8zzSfGZlWWquiMdgLObvXMJXEKvT
uiRuGX7OEN93oD7mNSeZTRFMljhgtQzzXjwabiKu0iwZf6FDZ2Hq164V7FpIiXYU
raUMZql6j5n1RNzS9YxlgfsdpL05K48hFlp8KmesYD1wK1Ig7bDyV668M2SVntEu
F1y1cHe/Sj7Zlkf48wEXUCJQiTDBFHypas4Zv///wxkhEXUxqUGAbuFxmmuKTX5J
sm9uR/dG8CRS/FmXxAj/XUhryo0bKjIAdGUFzA5c3r1l/BK7GwlD6IPfRgZVx7Gm
HHqMpb9mC7hx0drdbSnyJH+EaJHepUGq4jXyQvl1h5+iMmrW1BR1EyxP5nrH1Li+
5YHK7Xy9iO4edKVxUFtVZ1QVAt57my6N3hOo2NxODm1mcX9LWve1x+408gVIQtcQ
QCRrWzOTgV/87ghcl35FPx/Ul6s4sKCY320/ZqWAZgq+LTc5PYQIIdsPXya1veqq
kmXZN9nqyOvjhjl7ww/pSQYHffr1ZIrKy3UgN8HzRhM4MaWcieIFctUbYJ5kDuJN
f+qHGpPsecZDqIoZxOXHML4CX07aA3bXMp/pEBfuSBgrLwPaG6cOUvoaOgS8upx9
lGi2JUrOGd1BXuAUdi3MwkacX6ezIB/RAOpMznQ0jcxHRtuWDtY9eMri2kFH+Zju
y20TxEqcJ6LXHgyReHM0XrNftJ4QDGEDRDRs3RyAlsf8EAYtZa3RTS6GqiTMc4CZ
imyIxdou5+VJTDjcSNZ18Fh8k/EqV013VyDtqoDDFvU2Lj47so+CT5nPf/40XeC2
46CoCssyhe27za1VLb/xw4BPGg/qQ364ZH4GXejtFDiborbBqrAA/pQg2K3M0OL0
CxdfpkcZbv832m/W6bLZTZJPdmAiBAM/952S+FsU9zehw1iHFHjNB0WvGGJhvIsK
kp3FgbZfzoxr8r6O/aFwrRqN0H4MVPX/rTiTHVCgwCsNGxK/A8HeRAeIkOrMTuQv
f6LN0bu3Z5aO3cOKgU80A3W3qEUvcc94bTT/eEW8vKji7nP8O/owxufwg+lf9/tF
sNIAzWUB4aC1KSabAdwhHS9MsIzz+kqRB+VfKZ1K3o8iu890vxJVkTu6FAxepPAq
ZDkREeRMVvV/FKiUo/BTkk0tISjHzvAT4dIaUgDiMETe07l2wKXWueQL2SOQ0ezq
6GGJesUvIb/b7zAEDqXiZxsOb2v3+zBoo6Ru58h+yVuVrdupWqwDZxkIisMzdRc8
furCqv6BXUozouqO3zcpAkvJh/C/sI8iQDl7MXOjWNmxTGjn0suh5gARNCYqkI5h
hW+Kyxvv+jyZDfzPDo1YmHZCaNnj13fRh/jE0WvbJ10I4mcJpHBl3M3bF1Y3LrIR
fPkJHEtcb6pfBwz051oe92KqJBe9CrjaQylGgQcgXCw0pn95wJG5DvoALLltvVoc
T3wqLLsXShmwW4GJ96PMbd4BxC/w2gA0zP6FeGPXFYI0OHlgURJ5eFTnZJlXmAvk
buPsl/S8Ot6URZtnf7rwa0MsxvhqvGdHTBWCS2+FiHiO65gztzOlQEJqtxbVAvJ1
gLQ6ubqsx6G5kQs/Rk22Y5TSX2eubatK9I4YDuw/fzq/A98H/u6nlFYdD+B5Sz6L
OewQ0HRKP2uKM+sGuV6auCXhxNOBRB5+DBpBydikVhKrfn9p3m0fvndoZBhcyZGx
Pep6osV9ZyIEwOF9deIexrq545kYqeRtgXs0e5GvUI+8QAqAZIW5xCsdA4TPcA4R
8tAk8CwBDdEXg0QmjKXLiXzsUXvzb7LVb3jNFDfv6VB+dwU0ZC8/nG49HpDVHMmy
tZ8KRRaZ2IlWno1dx9HTF9AvMeeD8WRl880pmaWHUnM8kFp1ePMZUdlwYrSeH0rF
IMK5/Hu/3wPkM6Zjx5ho/DmKJMpBhXN6Qkva9xV3dWHjqmmvfedPVoLvTabTa0q0
BPb/VBVDEx/3mKVFtFm0o3Sj2jssVycEz+vi3M2aZ2EF7BJzdX6BYYBKgKq6WnDu
TR9YD6WckPIpTYocZSHsjv8jy16FKQOFBlBIbQjWm3UqFRLjbZRq8wJVli37XIc5
2KKtyQuBKJXz9mi6/sst2Me9Tzq6eI+APQRnjHj77cSj7J2QSnXUCslQwMfts8OL
P2qfUA4px8pGUmFTBm+nyGExzZAhNekA31ULObn0kWAYCBoQmj7uQ8UeVfpos7FT
aruxzSDV2vgcROtgDrpHDeXsXejh1ypSRHOMNMsBuA0zU3Ql9YX6kMGwZVbmQ5ed
KWhqCxq/Z6ub5E3BEk2wfHCdhU3ce/eF+/uAZwzbqzB+a8uX6RHvhx2RqO5bWc9f
pvmdnSZ5JA2g1CspnKjgKicpyn/KlkMkv0TAdvfIWciX9ayXNQQ+gUgauNbnqj8o
1n5AlUPW5X5Id3OMNfBRheKp9cHbJP0/Zt3PuVCbkxBY5uRfAD7uQCOxLtH0+uAt
0yTeRo6blQSpo8fyPgTNPpDkCxoE5ZII+JZZlSGxnqeZ2v25eK6xLPoWgudH1PVN
CvkXj/yPzYRT2e+guaS265HcmNVBRM6Oe+AzZD48tLHNPvcOWUouY87KUT04UP5V
2bbATKJFVdwVGln+sAs4G9kzEChlJu2LyL1Ol1VYyd7wdwlOgy29M2bZp2iR43qx
p7g2amnAWpSEf8/IXhC0/3K0uS4LqTaePSsX84iXS/nwrBxgXj7AJfk9g3qnjcXv
R4aLQCfEUj4j7MADtjs361TcIFvRkCa/vJRu178XBOmOdIedje8DSITkT4Q3If0s
XEu6HvrxEX2ieMitdEanBNCxHqa9oBYx1mHmoDC086Vqv0AL56IXhikgMUWzMTU9
ne3aOD2wxR1eL7BoYLO/ovYX5IXv//gmc46pjjTxpDphVcPA/ns+O+i/3ETGDKOH
hsxiTAOcmox37TXdcupCsuYkfAj2L+2uuri7DD7eArCnaqF8pnclXeVLSXo5scxx
mEdyANWoeC0AbtuDcWjio669oll+qiZxVnXk8OcXSSYbjAvH20vpRSxkX6+TD0K6
z8/sUgUtBvcYok7uL7VD+mVDrwJX/mzn9If5l46+7/DRsP+fNMf8SyV6Bm83MqwN
PmduESRCRHcD8BmkLhp+iQjFIMR3fE82W6EMHeW9VyPevgCGWMbP/zeYaNdIbh1X
fzCR7IaiskJARahR5DKJqNyXCN5guUa9AzsvEydG5d2S6bEai/QW6uKFUenIJv4U
xpcDfyhYpTX3zJXDW4LqmQUFueenb2X5czO9WM9xyPwsyqxP/ObyAe90P3oPOOgf
cY0IPNWaSKYmsuDkQ2xXTfDeDCxRawiDcFonYjZBITpRRFyHFKzRle04t/h73dfp
Mz/9gq4PO9tcG8ameLjzQoI/kmR9pJ2xg8HKSfDWUe7pne9Lt6BisztcvnWE+zj3
vOM7Df25dzpfocdVbrIkMwmcTy7Xq0nZ+2MyNmfl5xwIVb4xlRt0YdboTJfWwB1v
qgHbgeQukMo+GgjATesEGNaGIlZEsp5dyD9OBshV8+8ts1y+MqkQAeQASOt4bjxR
SgEiRQcCtTzqnG+8CjACN03oYrb7lBYsj1H+RfMTLaxIYw18Ln0A+BUxbp10QHON
3WT9RklBmtgCSa9m7WjUvLut8NaDqnfemtB6opwf/mG9qGCG783f0hUQ9UhGxBf8
L1ncPYhYkx/thkZ6BAEPRpGob0/QVWFRNkwRk1aMDP9AofjzCwjnoD7o0BJ7iLat
6QaIrMt1HIqP46+ULNXTJxmnImGopEYDB4AAo+dZsJptXO5NUXahZaCws822kDzl
oEDogok6Ut/io6VMcA6ahWwKmvH2VG6960Z8DV/2mb17+98ATlKfFOaykFGYoM3d
gTlC8XSTnBAmaqZfp7pDULIS1TC9CyHLV6X6dWH1C/BwurHzUZc3K7D7wsJuAtG4
anz06WIPPGqev77qjHbTAuE0/va5RgLqsaBidq8f4t6HOYQPXWMlU3sRRY37nsTR
LPlFwCDVPuyR3gy7N+pXe6DBL6EPaCTS4MA6AnUhCponV2Fv+qZd8v+0TTfffoS1
Sk9KswoF+IPm76ZI0u6ZHVoFgk0Ac1iKIiIACuMqnmti4eazHM5ZSptwU3dD9dfj
idAPvgr6eo7IKaVokyviGSFb50V5pM95IJRK3XwiDxYfGcpl+KqlmHWD9zvlTIAZ
wSl3GKH/xiy/w1ZruW3bV0cHL0FtrsDJ06I2I4Va2uO9+xHvw8dmJ1BZBg9NGO5l
SBML+P578wxPNbn2Xv4Mc3b0rRbamFOcFPQDmpL+YpQi6YHF5aB6phfR5jjlYQ6Z
vSXy6xn8NAiz/d8WlO3hrO9tNtjH/RsbWIeq5/DZeqAmUosXscEq+zXmX/aHtjgl
id+cdzHzLWXn7huekXAa/y21mCkowLXqbyqEA+rEzPPxidqi2xl++SJEpq9kCwTn
prnOaUR6dNz/ILDI98LoPTt52LsTzYcZtXA53/iOX8JUhTx4ZR52OtGvyoMw73QX
arJkmDTr5MyGfWkwI1VyHse7aftzU8FKkmIqZ1hha+tpaiO/3f7gwzGswLRo7wPC
FOrr+o1EZ/MvsM2XcQWn3KY8XTCh0RW8Hvy7LeZn5wubFGyf5aJRclKTa0rGGT+d
C+9P/Qab0qUrh+xzxe5c6DH0J/fM/6StzKroWmIvqak59z8OM1mJ2STSjBNzmjkE
eWUSK5CMMuTXPaAEtr4uaKLMRVA0PvbhkqEgzUXMfozRUM5HB9j8VFX4Od6LciCA
/LkT5ZrqlMtuO9LfKaGHiAqH1HbIhEjHF5Bfk94ZEoIKBe8l7vO+puW2meXNZqq3
pnYeT52vr4Ljk6RMsvaYbUMuf47vJ7kbTNmoOCE+mLy0be+yD8c8WKegBGZTmuLH
0ShR9s7T6bk/xR21dFL99nekWavuGfvVPV+mY4qN/NKCguc93WVlrdluXYQ8YLYF
JKhaBHfJGoJmfglEIT8AeXsWDdZHG6tduBGMyChPHE3wTRWiFRpk+2Eqs9KV5Gl9
9kd510pIwZ6VG7EuUKvTMSNClKD60REEHlRos5E09hcRtJNcT+xRSDkN7dgt01j3
uirNV+DRX3VAge9xNkOlJ0EutD5l52EpwYTTW2X9TqUNQpHhNoAYKCXsFPNBFLgI
ql0u1Bi66PaoEDdnhsMSh1PI1JR0TLGdUZutXqUyJSfHYveQBCaKWPK742u8ZoEB
ndxx3Pt9ln/sdH+fdajk+dCXc6fOiY8QUn5FWlbH3PGoPEwdQS6aFqHqePf5tZ15
lS457tSmuQKg6HJCqxW5Mq1HBB9GAY6LiMsBNPzxB1AH+WwcLjOK5nmmvTS27feI
8dTldTH67WOeZXJT3h+hNv6yA1nvRE+wB0QHg16drZGKhSNFwYQqrlpfezGNX1HA
rTBhR6vaS3vT8sGQUW7nYOcqQ2neJCNW2Bj824TozxRheJIN/7vZ/YSrAmSOX8YH
kPfmq30GuXwQL6Xxtbjf9AzoWr65opsTTrPtGWxfMu6rVQrzNIFzli0w3mFg8l2b
b939YxZHhrULA31+XRoGwpizrOEQ3i24esHU7LBAR397S6997hlswz7OcWoCdsVX
0gHZo+ReK+3K7NJe9Gzs27P+TpSuGiIdkt7YCg1WbwoS1Z2PSsPlI/MCzibX21Lg
1wALgeMphem7TVuJqLWIJmjppRJ8IBMuQOx8mEZCrwiJAGJLY2In2jFHSesJ+1Fv
mkNjxDviTS/giD7AFwf1qsaWzie2/+d/SeL4ncjC+m5+gPqv4jXu2JXlTYKC4g8Y
EQ4ndhq5yzQY3HoLmxB3KKu3OBASqzL0qAVYaFcU+1ZwuUAp5bht2i4FAK6OJ+6z
JtV29ysTIry9aq9BhehiDfMiew433yls72s/5sO7L7Nse6Uks95FZtNAVohruTXi
BrclLpKQV8yrtN8QDA15aQCgA/zQSm6v5P6dXHxxlkDVouulrj3y8ATib64utR+S
qozWoWEnQayeIPAgr460vn9Dx4BrDkHSmDRV4l67wt1MtrcfCfZNFrqUhXtC7X7L
ArBgr0GWJnVoKLzZtXCJHvO1fNIx2g5oLVRCqNB98sPL3D7IVbTsQg+azvpwabYp
1asxYt9y6clmMB2NRtl5z9qweU8DcdRVgYPMZxOvnKXYGQ/vC/eABR7T4NK2OdYh
2vvbt8F9kVlNwAiZVVbM6IaWsV2+m5GzkLo7tCdgmBieX8gugL4GGkRxd740FA6r
NpfWFUnOWDpzUsKW+IdV/9iefATKRCqokA4JUcNd7cW4gzRtuKTrIiH0l88VsVKK
bps8ICkZL0TLPEJtNep+SITys61TbDsnBcznCUk1h+9NWZakKFVFfzrhpVYtcXLA
ja9yzeQFQidlnEA0Q64ItjOniGFHItQe90VHLwemBExpkfYPu9RKYDg3Jv/2J/Et
ZmR5RSEe1mC35P14edPwrFnjkQEQY3VcFdn28YdbmsVz5eeBduDTRHpkWGStG+eo
MQLQnOwAV2dQAatcvQBAuesqunL33xbOQ0bMKnbf4FsJWPgB0WSp5ZKS7AOlaSDa
NkdZEsfK/bzaE0olpz/ZEp7OYnBqjQmmJp+BNQycusIGtEyOkNKrML2JbCCvYHEr
XQDZBixhuiUOh3krrNUBRd0nsD8Y6vTZWB9aFqlc9RgsVVSMHcuK2MfrjyNyLaTm
6NZihMk4CLr99IV7LJxhK5oyL+jR6Dl7T2T+Wm3/qTQzzqjxxJ6qxiWxkpKzHG+F
EN5lq4s6QYRJDyz9VpIVQXv6FztNAOK6rzoBH2CS/QS1Re66ZK6qoV+2cn/hsVKm
0XpTk9p+ezz5sWzioB6BYY84nG5J/a3oqJB2qzCufLrtMd2ppo31xwtIlEJ53+XL
JpMIOGCEcf8r+/Xio6seyKPb/phUbfeHdXIFpsEosIvHjeRn1+N1uRnTHBK4OoqQ
afGufocb1oyh9Z/Y6wZxJj/YxR3bAG74boWnqw20wNEvN5C86ZbUcJY44hpn5qLg
AuY7LbCUIOcvmhrX81OO6AM/ywLGl9LRpUWMVY2liLv8+hqKy9LHAdEMgmqNBr8k
H7Iuc0fwCXhCbaG2YCy/+VzN1nx0a2gbbRDMwEJeRSQ4ledov+nsbN4v+UJW5C5N
RX0KFuZadTU+l42q+dUMZ0A8DhAoGxxvuHK2U0K5waNSF3isr+mVc5EdBpSl4qFp
Sh1VxCZcaik+XjhI/MGr49Zdu4REZ/cPUk5jmYJgjIr3eeIB0257k4Rq3W0XihDS
Ij86uDssF/+DYJqxCHKCi8G5dBGd27g1RXA/kGMCQpoR+IA/9F2roazPPxmfnQpX
Xv2Ptzll1RsUzd2nKC6aPU6p7Tew6u5fMsRBu5KOzkBjqlvYrpk2aTyzElNgneQE
5EFmiqe7ZRQLpzTH4nBnbvJpxa/3J4v+sO0PlmouUQ2+31Azj97Lb6ou6JRO6xhK
Bug4ItUwjTA/2TwPKGnka1Ij+4kyXWSgccDXun2veMLVBtnsNwXKWJrN6pQXMNyb
sOFlRqEkY3Vp/hvY1Rw+QV3ppyj5UgKpq08beZG21cagTw6+je045uwyMN8k/ALt
0vad5McXqN4WtsXipWbKakDa9YLzYmiNa1mxAnYf6Hr1ioB3GebFAX77Ot+rHLFy
NNx6FcAMAEzHU1ckfSd0ONjBGWUJgQZrlCxNa2q00wqvoCsdj80XQuWD/Lb6CXp9
KLKlQy5g8zcAWKuiMBMaTfQAdS1rADSel3myUoyaVEGRbNGqKa8yNaUZsa94+yKX
q0qlGL3ASxh1DMI3+m9gwuwXRrzZvrzoHhO9GxKOrCiU9itVjqR+/13Y8BCF2Ds5
KFv1lcyFxT6Kw0x1AhRCiFvosb5dXNt91teJO/29EGixWEzOQV6b30o/XZLiRS2r
72+nA+Q62ySb4Eb6hPLxPfma9VLH0erVWVhim7UxzsC5d0e5JByyc3A+YmNOaVSW
n27xqVRFLy/JAEVZq0nMpledEZ8cm3zppYcY0lV8IGpCGrCeDS/sGYATaM+CaSLw
E1C40acSW6dovCxZLrscu2R3vanCoxb/vt78jTKNdv2S8Cfcf0xgBAibV6xCUXZG
4FCC0oKnbgSVOTwd+C2VSk3hHrs3f6VMzkl7bTMEMZhnIteGj9iOhzd9KbAI2+OR
iK4jDWNEawEsRVNkg0r9hSFTID6LyroZ4Nor2B3dxWVsn3cQ8JdDOSiEK4jrS+qR
VMO4D4siCvD0SPU9KpKAKGRz4Ct2vMvwJLvOz9TC8MXtTMqwQnAHb5U6xS2Yt2c3
OeuutICRvCLSqktrr1ZpjQQeKZ2e741sLGnXP1bQLtMuPvxFLgTsgJcUmkKex6GY
Ev1uHurWeVFOWV1m4WKRN0gfXs4oE7aXRV8eN39E45nnMYApTvbmD7nFR+0rebsJ
P1n4WTNegI/0eiA56RDNZ0/etdcJLAx1+KxXxPIWgTnbE5yiRijLN6XohnhhZKO2
rJgA9egqXfo4OG2UM5YE2sjhS6ckTJv2hRKjb8EfINmCmZUnFIaxXXC9w9Xlg54r
idoirnz9VARSzZtTJQctuDdiLRFvVP+ILLeuHLNlEhsLloy6bdEUwsI2UuSmYwUu
WaH4dws6OJAEqQbFM7VGngPHRdcutpm+suaVGhem55PDhw8exq0ddaqLOk1KGwBf
vBJNhC0tbH2sW16VG48A4xN0v5RS113ddS/cq5mb6+I+MMv7mHIfCDjZ/0MmHug7
l5qbrHXEcZB+O2EsWNew25Z79aDz0upvJtc0U5uZ0v1ujQ8jCYmFzUyEZeV/X508
FDww2LZ3vo3iTJOMp0Lsb97wbkY/wMON4WgiuLn21IIQdrpuPEmoZXvpCfPJUAoi
XboRIzmhcUYt0LMO2D/Bl27WNQksqVCvs7likJspQ8J35M4iuAnklOzhct5NmiKI
gPumsJPfVKM9ADbFdx7a1lBrGyXJqBE3KaSZKJi8ck421PE4xamdTorNPsqjCv8V
9kKjpnPlRV1wheX4Kkt3M8K/OP46uSfAGPkPlKS7WvIrhiJ/mAM3LiwlDj46l5B2
Vl1MesxJEIdeXxpt36Fpem/pKdxN8RR1EXU2nqxHcMSlBu7CWQzUfXHJ+HifVFPC
uSheN8oY4U1DusK6P5orka3oeaq0t5pv4/exXEvblKEzhGRE3kaETgHPu+DflBfq
eXEiGj5HR5Jm8D5MMqHAKmERWxx3HIIzWymAAaOispTCF0DMIWptRITNAJBXpUuu
B1pUqL8cRvoBuLZNPlYUus5ivU3hmrbipDrLP+B6HromDyxCGTs57XQdRsTfpGSD
1vpVtAxkuSbqWunJoBWQK8Dsvug58oNdYU3EW+lImDsMaGY/1xupwV2sgcU5UsJc
jx/8Sr3Aq933Oa/6dJYvfvrMraN0dxLQJxWZHkywpbTNqeM2yThqlqggPkJ7mKzx
LLWGGBMe/TQO0G5S1UILahur27tcFkM+JgiOy+y/k9vrojpE2UtYZ4BtbjPw2czg
rwRiUYGhcp3TjyPbWzbU/B6EBHf+IYrXM8/GWFnaJ4oJP5enYW7D1Vq1UH+zLlu7
rZy6aHMlHVc9XqttwZJXSdOSXCLuopCmp/mOxjgujsTcFWRQPncSwYBUIoPKRnEq
V4F38slEfUFx+CarwbosU0wfeAvZnTG5GlOmDXgFMYKeNzgIGLTD1cfqEaY3GEte
BabfWwulfBeW0OUo/oGamtZMmE/o0Cn/NySXT/eGUqbsrLIii295huKEfcyRrs7T
JdS/SW0n6CDrJ52WZREj/aUqxNP2ue5QERbJanANG+IIc+gH7Lc5gklGrqISBPJM
vnIEIlB2k8PDWNVDKD6Fl0TgRbnCkfXz+kNH4QgwTbJwGGNchsYDNXI/lFQ8KuGb
TRfKth5yqzHQ71oD5CdL1rtvxYqaQYANIqykGBFSp3INeSq0x964c8LyyrSB1iVM
2MSAbCY0p5dXk9c94OvK+1lJoUf0s1ml29CcV6c4lBWGhH9Z6WJ4ZEzZk7kQRuOR
++L7bs1Th/7UUKwhws53r/pfeSxJoKZVBPkaZpOl7EDbLVsKmMbCSbLQ1il6lmzR
KqjURnGpZpN1+lABzTJ9n8HMiYGtGAIx9yinUicCCihkuvELMXuZw8gBtvpBY0il
i8Z4OC9xJMura9PWbTNGEQc+CfAoEHeF9/Qqbe0Xc4bHyJGNV0KF19kCvGBo6nG8
oPdRtnFPBoFBCOPkIR0auyTLiBFmpW25UNeDUSyGTnzbv8mqDAUhEFD6ghC0QpIC
h12UHFmNl+mThUUKGBOF31078hDqSzCPi4T0T3e/YUjkGrrtbOkm3TBXA8ZDwq0d
YJhHveSvWf9CKV+AeRyHyPibC56d866l4lVcHaCKbmibw/CvQrJfwTExsMMdD9TA
qgHNe5ELnEd5km0F+TiyV8l9hVbtpvHa3prxiIk6kcZ9E80YkjGt7w2Ou0EfpWzk
FIoFaiaz4HyC9upCJU9k7vISKRGEZUPw67wnMM3RlcNO60Cwjo7b4d9uCfkPFzIp
xq1G7YhTzhN+ollKHC2obZ7fm261VPbPMrZreha+5p+gyvEYRoe63gEUFCOT1Bsv
cQMxXyk+Y3XMHQZEV/+MGaZ72A826oysm5RY4pCtupp/1AzE340+EMjzVUCjOAdk
LUfsh0Zvj38wi5VZD3zdhlMPj1jMu6qNQ6Wh2gplmfNMv1NV9xfJ/O6CLpHXkDGP
rP8whT6wZn+6zV65iGuo2KL5CKCWGk3VzNl+GznaTbKVcdBNMBhR0GorSHN7AAG9
ja9332/mWwbt6Gx3ySCqUXyOPx1OiIrW5t+eQfgJpGzNl4EbNn5LBSmZofkV0ADi
QSA2ijRIXds1rrWLZAIydcJAkRwGrdm9WFXDH4y+Y6DqASqpSRX2zKNUM3gzK0UC
9e7cx7yqC1LqOskoq344rRHHHKZU05j5qCTtuldOd8S+N4lavxMD7KyEfGh1+eMp
ZSXoriEIt7PirR+vusI+fBrtJPBrgif9Kja+wP+wjf6Q8SE7jpd5Bg31+jfyWKJU
+HYqAT71dBbcUfDz/NgXpi31hAdr6q7E29ehdDPFkpb0GXCUd+MYxKDxGLTgxgp0
0gJBw81c1l9HdRlsQyQOLIshMGOWtT5qd6lcbS5uUwNK4ZAjo/V6R5DOm8JetzA0
avc3DObqXTg5Ebo1lSSGCUPsL+WXgi07BhJuuGgsE4Tij3L1fV4rv/USE7PL7jSj
XqNaWGrc+aAIsb/uv6AGD8TrFvJBEg9ZZIVLPfAkym1C5OmubYFosVHrHS7ZYpZj
nfNjMJy5poBuKN5CRLyn5VGlQHQV8Fxn4LWv43X1I62joNLYN6I83vRgXR430ZqW
KvW0ZEJPyjXA3pQRHA2HamRGJcMx3S/LWUczMNtVPtY7QmnOBlmKw+hFRyVkEelL
aO9Z9kqn9H9P+gB0xW2sJOVn2mwYUXK9VKGWL6faJbXhPYpdU68aQk2HxI516GWz
HBxHIQVy0ryCqcj2xuFeGOJ5khi5RbR/DO/1G2iSdKXRVFmEmlRcfwfiR0zR5PZP
O7XSYxvuzuj1kgeB89bPRZdILxdiqvPfesp4I/kmBakbY/cM/aqbTXavmrzsfYSD
KUYh+jk83DG7wbyB7u8Q1gRc46KHC/CYRIVW2jhCwAUJKc3P9wrgL8/EgeBO9pMY
nmJEJDF4f/5xDd8jEk4Su7yFgBbN5KT7xfJ3eDxwuBDEbOELhDNerUvVst0i97zH
jVSAw9miuJ48M3AyBezcuxLaXvh4AtWtd0GV4oHWt5qI2mMgjSU/F6pilpyaZ1Zb
nI340rb0Hlq/UVEJ3arf/PkqXQvkS3qudaDYSJQKXvZL/6421PY3rZKZrZ3KAK4Y
L1B6dGouKqAXfbn6Xbh9eGXLMQjtDEDA4D4063vFBS97oNwKbKMR23AMpqRdSwQ5
mQt1tPaLixbE8tMwtAPtYMY1/tsJd3Kz+eIWEAAndq3lpQTQwyIZa4BLrjoSd74G
o+65OidYnjHhxSczPCn2UI1aUXNGfB9BtRwMtWLwVu4sIMG2Ejp7ti/t9ey3+yMU
9L9hoXIF1+rSgtwLv1iwZywHhjguCeFFyglOOOZ+cLVOYUODOg/mOh4+QpxV0b6q
7W7Z0SEfQaavern5Lk3XtoK1+nM1i4zMGqctgy8YRdi5ojgs8SVo4UGWdXDQ5FQB
xU2fRA65RBpGq0hQuDy/r3L7qzKMTsrylfjGQHypkhANyAx1uV48Zsi9nHFHD5dX
xHG1xuDFw0H49nhprBaoyZ8Y0tD56+NueZurwnysEqhfUKYm4buZFvsfcl/E15S6
rmN6by2WnLqua64Rb1m+BC5fwBh2lEoAPNAU9D0u7LJ4hVORcoCIslmByTf6d1tx
ZJ83pLJpd5SFe/3jDdUlXOuNgH0M+q1oZ+z6jb3k7Bw48rwMhGhzaLhTgatcm4zC
QSmnquHZJVOzqOTOV5YankUNl+WUB7pOnQWMy75VzpBbY6zw6VuFFNO9ClbiBLWY
FpBUpxPjZtFpBR0zbys8nrjW9ZfC7uukoxoaxHXKyAHPL4sju85iM6ZQsrHS6Bcu
pMhgBznuwFXpJ6IYY/liacq6yM+JehOC3//wgRLlSqbVA9qNqY+ovm3XAMiHOLS6
i2WD+sEcYCh9AmZCLbR/oxaF71MLW4nesJCaGZY3twdMAgnTWIR6GGsigGQ+9O5b
5UY2jTIqlNs/ooZywqEQvCrmF1jZnFVcVqaaFfkEToj9ZY6ShQ9l5Ij4q+HCA4EH
QA+bcN+o67G3SIV0u1rvvbKRX+j+qT6RFwLp08Fmh1Ivt9vwvNz9kGKKQa5pE9px
E0NQJ59ZdnGFXB3OkZi9jK4k+/W76i+d49ALHj7AQG6/4Hl8KSrHMCK6Vchc05/r
d5RAN3V5pxwIg2FabtPahB1t+RW+Dj71gZV/dWqkxQ4yd5Cw3RJgsDOzkaU54f8F
GJmx7+muX/np1kv00A/k5aSj61o4QofL5/6JINOLcyO01IUL5moBvicurB/uAzvn
65s/svd4IrcRYHJyihfhJ2DHRQfG7QdFYNcdXZZ9rA58Gy6kasmCoai/53fQCCPm
TDpCUu1N41wNpgYZg1sy19UHcpIujgJK0lCOCqKhYNphLNT4WOVj3MgPb30RgrNG
YZSAqAReXO83ncRhF2nHEoNrT7UWvI4UzTyiaTe3mU1v6gop8M34C16ttxq6a4OS
3TSqgfeVms8LHUTyfqTUK0ZsKaQkaORHB7IMv7NzP1bMW7Se4fwkeHD1HYBdLThK
mircXWmQs0xOMOMlHisExJvsIbcRFseOateZJjPnyVyZTXeF2K6xu2tJB1tg60CO
BoAdjDR+B024iH2aaeM+goN4dW2wKlwexyVoiRQaz6V55tdZj0BnttjHKnlaCYqC
Cc/CWG5fPXsToeYaB3EBXJepU881ss7s2J8bTet/Th92+rk82BKeen8j8gjlSfjO
z+Qd3ifyZQ1X7JOMrWNnh6SBL3rTRXc8iA+xQunc4bcsa5gDWbYA4g/QanDm2woy
8v4c8LqGNb2+j0VYEmNdQcspkbIvq/f32TKrgtyBiBesaVUqBRI7B7+Ix1NglOAM
UK0PJHWTszEwD/LJyTETXpV3yXN0Xy9EUgizuNQYVUF5a2rlQluVOArykM/5uhC0
nJPEba7aI0/XtBBWhYmfyP0A0MbnbPz1ttziAUiC9N9aZHB3lghIamnUyv+cSnuf
YNB4hSdjopmZVXOTcQSo5Stb2KdYva+jlNSI58H5SHnlYHAKaiZbzSiVYqi8neTS
1fANJRV0pU2LTBBcQGtcd+u4X1l1XWh1foont2awhggFHIjgz/Xq8Hcj8JEesZY7
ycxW/ZCOrS4M7T9PjX/Yk56M6z0fOq67Rix2UPzCX2zVN0vN+2xCF6P9aOiyuq/i
m/c/37jZaeVcSasn2r/5PSAJ5utJZCNCs6yM878q6O9iMaL4bAIChuGzOcAlx53A
BlQpsYRNu97ZeK95AezJz2jGW6a6QB4fsR7e4BBmpq3rU0A0sG15AVnybkiDPnAK
wmhYYN5PIwxuCIKKBlV/wS8coxig2p0qskFaA9Ss2Cg2KCvyotQ9kwdE5nqrkq52
fG1F6xX4/RDhf7dbc+4wUS/O2fA3/VNXcrdq6uPG7cS+ehWDDwpTpG1tTbDbvtjj
JMrITE9gzCleXeNt7Hr6Kq5+ADAGBPHPQjw+dJVexFTAY1+zapH5hvrm47on07UZ
XHK4EWfu/tDs77K8q7xgx+ND59hVIZ6DhSarPo3I9eGdaWA2jJjqexyowQ7QHNTF
17HH7UIzA040M5Lm7rqL5ssL0zz330Pl1TCzAHgtxxUsSVLqRLr/kMDGL1yyk0uy
XnSKZxdXuey10M8RKK/4cJ5s+2AHUgPmJEq91vaDJHdhRZbkW33Zb/4a5FJ3ikiA
OlZj73IHImRohuaRwMnUsLfAgO72q7GtDDGdLfhWSizAQdZhuDOTiA1n2de+lKUY
o7k0dHddnc+eYo8h/XZng8U15OAmb0GUfhUBNUykIEBPWNXF6NMk4Wqjbjkcb3AC
dTeIpTH+DPhR4Q8NZBtTVhhFGiKcOFbtB39VY08sZfItoq1PkT/n7+eb48/QsslF
JcqQ9Ayedqbxc0y6Fpt0Zj7HHq/qV1H9goj+YqjrNsMKCD6R7JdxCPQ7ACC8TEC6
79LcyeTi3gkMF4flHAtzWmcri9t/Iit9F96hWNyD0sBp1m9KZ9DSd7FcbKwMtoHu
XLOb/+CT5GW+LqH3AYUGlmNJrXYafS7d7Jccr7/NB6jYOdpFKRfQJwD+jc0qCOom
CPKXAVe1qn1fpkvsmzQI0/oyBV/3eACX2FA/+I4PxSE68WPZsPgPa2BCwpiH16F/
+eqtCh2W/aMgYf+QRsVfM+mA/GP9cNzk+fOBSmZmyHJd+MVi4IEDyXGAv/Zy2MJX
oOr1B85fYUSk5D2YT8/cUfzIknk+03AD3uWvmPf6bJX6dYM38j5KHZPcEcwir5xA
gOvp2pFteLEhnScZxt56YnFaxVtC2r74TROdGQK4MSMJcLJxuJtpmbFXzbUHSJkd
pS4pxqYAcXvgjWhaQdmCzECTuT5PUoC2vVL1LWtalCbsw+/KKJRoP3UXJes3LQpt
EpOsp+Sroi9B6liSQqBHwKH5zwLlbNjsGtHOxjthJKROdXxLwsPodERCubBzzRn6
LfC1Mrh/H7tPC4Se7LSiKCCos5246/cyVxdRZSjkns71kDiUwH5ChDj6UH1wR/en
r9p/fUsk1r6HYgy+UyJOUWG2bk3cSTBtBMQ2rCsAwAzHGyrfjh2x0dbsn11EWFPi
yMzLpd/irvFMsUkvVSORHCMrJaa/eErC5wi+SUgs4owfbuxg4xYO+VyfpwYiOI52
J06FivQGCr+JUkgCR6jtA+/w+SM7a3vJdVVY402u3wuOcZOMiCXTX5FKD8DKyUZi
d4rdCj4aJ/bEpw1Xhnu2Yepl1CL4/zgt8rtEPcdDniwybYN9tNUMDbaDHlMEGhh0
q05G0F14IqVKojcHofmsK1eVvOfc04fdUKnOzaNB09pdV8TSmptr0leUvPKF4jW5
PVPChjl5YyWxUyNWGvEsqevHa8rkDU9GHB5svO8RD2g1RhDa8yKb700kcFrR9PfB
OWXBzup50Taw9Pkj5pVDFFHyDD5zu9rzzYE4ekcsnG4oCzl0JxK9/P04vl0Tq/WN
4IJtyKkU017ILhoBMNYLn8oSJ+NoAyb0HJzcU8GyWc9lpetn/+gAEl1H3/UMMC9d
OEbw5Or2iK0x9Uedmh8ES6nmn7JB6oebzAAfAx+DKNYVf6rt5zbuWxiLbfa5EhgD
BgfjPJA31UesPlqjm1UrpueS21yGgHuw54r1hbryVKUNHrC4HrEBRgKt0cF03J+y
uINGx8X02DNoQSCRbXW1jgX2/ko2UAulvPzgU2iv5sSnzJfUc0Xs4/DA3DwuL4go
hgm044fv72YVBnHhwPHKQGBuXipan1ma/CrIFl0Ma4lUjT9UWqD1t3iX3ppkey4K
2qrdRZrY/1kd5dQ/lHTiw+ENItcAeK/tSuIKc/QbtuXt8exnrY8oYQw+mQpkMqye
cYO4ryHk16O6NEr1lUKzkVDLom9NjTQUE1KBwemqhLllGXXRQbB5uJxDEjJjXtjW
b/AIYs+ZsJ7vhcOnsrNDzqDFFuIyLCR5zpLV8koEg0iPydkadY9mCPmSadedDll1
U3EfavpgHfAk7ewMJO1IRY3w/Z2Kh44ojxbA3aCIaXY29+EpIXFPPoj4n2qBMu4n
1Iu7QHwi7hMjGgyEb3l99OfYhtdhkXfhRTavgJQr82GSbfkr96p3xYcV4wTgYifs
KJT2mmxDsO2L954OWteQk+m4TupSqbaSGk8QPUDC3OYyalm/R9Rabv0LaAlh5V9s
mYH79jMTzME5IFgzT5KgFuvYtvOUkaMUC0xUWPmGHSO4cFnPYOK38uln5n8q6gij
R3uf9J854azrA0bXlXUBealYuRg7ba4H49DVtWHhpBNL4eybkHHlEBJ8lz0kVdGp
Z3foiozGMeBfcEOWgrc0uywz6zCfa44l4wbu7N9tD9sN+DznrGU/WalSZrR2R1ls
UbIl9NS08kauvjmMSicfqT5qyGl8WzDhFMKFUNT+2UK8/YO3bTT8d0XLvah0BiQR
o2WC0p4skLFbTL3MbXLKaOfrOs6OIUo/PTXVOeaE2zvbR/W1i8PiwHXAYllxQpQS
YpIp6IewStEy+9WBb2CUm+NErHL00ZwGt6BGHbWYivjvpZcCOuLYJ2VVhlNuRFCt
wljY2qwbFlzqXpX8oYJTvW5FTOssILaYFjNbI8RMxY+RUfrtEuSkQHt0tXU1wlu9
/z9Z98voisnOKNh0yZStRiDTW6VHend+5G22Ab/DUUausID64ILc0m1gvX6SmQr+
gemIUIVJKoJWv8ZMl+V8wwHlB0nTXLDKPwXdQft9lZJRbZGfH/pt16fMFDHBcpBM
+nC7cLBJ5yf0pIk81uIdx88BGCQOyuKypka2/nfaB4cj/O6KJ1J4K3Y/kEkkYFe1
I/nlRRwIxY5254IFI+nwnUDO3Dhhf/ltIuIOeyw2/bsv4U/M2ckrBdoAoU62eVb9
QOHOVlD1ycOsVzdGxtPkTjn1zK/qCO3zBxhR0jlg+WJX1Q0+LabbJHuow9qyo6lx
xZseLVCTRDIyDtX4XfbjqYF4IELIg8v8ctmu3P8PU21hKuW/x+teQDAT+pCwaJS/
EVeIuGccaRZGCdt1ikmy9oZb6sEz6E9VcQh3aE2/XY0dv/NPsPth9IOMEx33v6qs
Fve2dLwcPaQ7yAttYzMuPcV+LqgbV1YpPIsi5+vLPv9iIJtd7Vuwd0OXAfTygK0f
FU8KyWjMXffud1UpK59EfRXiX+j6LsrmSxqzpDzWY3Hooc4/nBNnsG9v6TaIavX1
8/UMPAQsaTRjh/KDHQDArO34fjvdpNz1WthUITZh+e+twf9153Xi0Y4//IiiKASk
MVBg0xiP/ycxKb6jmjKVTPyShCrEcMAfjfBu5xYrEJrPIWddQxKss0SJkisIAAH+
b83DaYw9/PahbMdAv5BE4M307QJBFaqpHf4bnk6Pb/wyrJo0bOV+m+9tL5r+ul8v
aYJiwKqB30Fe8x61zlawxTvAL++/hHhLJ9TnAAV8pExMZo7t7pJhzbZ5NtpmgxGe
G/T9xB27WOI/x5PlcBi9m1uwFQABNW5NbpZtkJcnEZitCOy0pzOcnnRtom2nps8u
XXBm9JtqiKT1q1DsCP/WbdS6cDRdwEnXLlmlJmcLve/XoSnXBMMarz9UAXtvh77j
cIy+VBs7ZvH5jYTgvPwEnxBl9tRai/rG66K0gz233rj9WzTDoHvti1bEKWtzqCC7
oQ7+XGOSzjgoAiX8FxsuKuUOIiY/0a3CIeegHrgs6G+QEB5CmahrjOjzcrfqm7/q
F//N9BHATUtdmU1lwQyi83Yu5zy+bMjLP7Ia0Oz1vZzO0rH9J0u12aXc7lB182Ms
vOcXBBOYT86+leT+x5dHk5AsXUF6cYLV6ROt7i0GpmrhUHa/qFEBIQZz8H+CqXsH
dOXYHuCXwrWap0DxkJewKTZ/PpkGtCHxq1wP9cY2MWrvU26DwVuuPD5jjNr7xLwJ
2hXk42CZR63kMHrjVqOhnFFjtOTgCLdHG+K5d7i2htU9KyLjjH2Vhp2ZGsteqrSr
whgZX6WvoXu3EJUj/UYgCBQ+ZLR8HfC/p34HJ9FpCQsaUchXGuQXLtAy45mPnoSt
3kiL6iDfxT3/hNQXffCgKSUatnCYIAJARNRw3u4iDhdgTa9254jkXVuuE0AvmJeZ
3bl2LP783GMGUyvC1yPJIBkgmwTnQe/sAIzeMdtvyeGMpKGB4xh6ap7pz7gcx/su
mNKJMoJ1tG6RxHJikiOpF3OaJfAKtrpOZdumoFJ32rZAJCYngp+NYt2D/foEdWHu
nBqehdEnZcxb9UgIHlDN6V6L4QYdrykGV9Klcn1BrjHL/Zk2skfd40XEZPnWeUcy
LsSJIjzoG6tKQGajhItnOeAh4twSEDgkXz9cYrjBzHEW1ROoma4RdIOC2o1Yoxa0
XCYDPF2RFlv7rvg0O3MlvUpU0EBWpOSj0jYyK64c+d4Xrtps3oh37JGxW5AI5SOu
MeT6/lu1cT7UVwFFqy7/hd5B/urg0kQsrPqJmiBy0WB3u2cMSo7wm6XpUbUAGJgP
uXS6uyX6UkAPZ25rnEx0OVCMkOegBbaZ4irF34PjscenNo/4dzSc296/RP5RQ1kX
1PsSR60cHaW7nMu/Yo4+fvEfpeONPmr4FKjqWHXAwrgzV+22vlW5h9AsesUmQFo8
BZNHK+oQJ+DsMffFWx9Z7CROXiRKXYpmLv/LYxhDY4CDHE3AXZW6eXqrx8BZ2TvV
M6TSmWgfd6/+mXsAE3jMwmcKr8+UB7wbiteE/iB09N21/CYU80D9X73E47HMNwu3
q8bC6HQBAGSBQVK3DXfUxN63rxdMGUWBex9nzWX8ZSlVBpmpk7m0d7Lkk1pfe0EY
kJ7GervAaKByamXjjEXPDg9urYo2jBzQego8skbpOOi6EcF85FwO/3TxJyhyx946
zcchxrqy/RQKbin6yWusfKecehSNUriKkAAsnkKP0mliOxNtc0P6J5rxQd166Ild
GV03SAkKhFI1yg50EN1jPi2AeZOd6i2QvUxItzE8/JgB3VOwOt/iz1xJwCmyuDod
c4trJoLfH3R1L1AabS1fma4CpZ6ciw+RY5mWapBo9Gjn5rBiFUcC7ebys9BgZF5j
4Sed8tlt1V9Iu4uT1lW4P+eZzptkXGvVnHeYj7WukEzf3iGFKtG1ZVCb+9uDth2A
5BBGy4TojE3oxMGEV34SPYp2br2M/B0wTzNp4u51rGj6r8wHuq7OWCDYO0ILGxGz
3fTRSabJnY4zLx/3z9zz2lxVsG6ugzEy+hrnu1il1dRmO9dnbacsOOR6+lAPSF4S
ZjFPovTGXexgT88GsN1RuvS+VlFZha/1YVD997LmwnCkky90+XahKRPay+AubGRd
U3juS4JbVUsqtYsxPep6nHjVgbgv4ACf2K/SxFDxzUG8mHgILFtCuoUil2kru4Gx
I1LQomFTEUmppVWK3kVM78cfEiwiGiTgJZAWnB6V6ronpmLv0ALiaSdHzZ9gpOmj
BhS+LnPoeagayxoDyv3e8QvzrokxA/57Tw9BSYcWkmAOY4Z2/joWo05VWCC44j/w
MrDQ8fAjs9Askd9IugOF+6AAqIvZNVw8VvKoNFu48njd6DywWLvL4UPbxCm3sISU
z5hLfhs4ahQ8Y2E99N2STiKnDspb7xlUftDGqgQNlo0CPIMNDqj4RmubKfB7J9se
STVzUAKd/UfKDaF7PkntaMmLi3q0boVyK3SZBn8neBzt5NMeCroRs/4j3RiK3zyN
wVmkMv6HDyqA0tM5TPQtWFgfuw9DdbC5LuTjw+hbOXqn70/mWSFEybbynroK/uIK
Dbt9HnXm94NfE3l4DyVZ4Zp8hVWmW7IITdQa14GyGK3EJtJHnOlZG09wa/HQRr1F
EWwT97XiMzPkpgdCESjDtiG5fxfWR3QBnHoXdv0e4eMldw9OS2Fp2Qs8OxiDBDjH
IKCb20IV2vezAqIkxtLha0HQfcFT9oqYFbox4WDi/jflEF5pXUjyA2/OjrI2BzuD
cdAkH7sOM4XpnIwpLM3WG03E0DTlBH8QMA191xLtY+8nU/ti1qSFZZmvHItDpQF5
D05OTHFaWST+eAgKBHc76HQJ8ZRpGzhWPjq/1oLk2ylkuwLleSGM4mR/orvw9OAo
pK2kfiLIgkfvu3dCAhM+lYPQg8WZCwm/RN1pqQhola3bZju3dgF7545JHddEyuUJ
/OeGRX73M54VVevaxNJr/dAk06Bkux+48ogkEoILo/fabBAJcayfR7N81DkxQo2h
oXkqpC1HIcVNU1NkfwRbA7JGFDDteaqxA8xvYH6/+57fIgdxpkQLi+WSHFmNBItu
zOsCiRdaBtbxZJyVJKsIgf0ZKdlneiY28m5SKnuGBRvTNLzwQ/GqP6k8Rlr1sJca
wPPJm/ysitCYbvecER4idGyhcCIbuoR1pIEcL30as0bmTJoXeMFNFhxy2oegSCGs
fb2o4It/8w8EVzVWBGMdpRwH+XgBbMvWSQL8jppBu1WEnGiJRbeF1JfLrib1BwRb
MmVWurFwqWT5MNZ4sgoAr+BcEjQsnP3LjOdQD9t28n70u4JP8hCgQQPXTLq4O8uZ
ZIooqQrPU5UPcRf4PKJl5HphgIoEwV0PoVQACajUJdSF8CXcEJQGWBrxt8Abj6/k
zIvbs3PAzpyb+6ZMfU1XY/OoyY5a9R33sSKNB46anWoPZQS28JfIiwHMQw0fpoQH
vB/VzsJWd1cJ39Y9HposO8PFHOHmN7xPveRtrK7gELgbUtA8g0u7hPgC8QPM3SdE
6XnKsyqs3VVQspdj0m/cCcQkVAELnF/d2jHLmZX0kAokX1RxJt+kO+vdxqE9XOqA
cKj2y2l8cpXCMBnghwrGT+rOI+nKKskRF+u2bGZHdOkhFcDcoghGHiAtnvJGjTpb
NUVoornBUZcT1XzGkwh60tpDX9Km/F+F+JHMvbhMg/tNoYaZKRuHBCrcS+NI17oT
9a9vjp/1t6Ez/+o7635sE9tevAgWpRB2q1/JywdpVc05j/69/oubhbOmwEry8wCT
5WHVXpvWFpTWL0cfrzrQ6/mHGDL6sM7aYZKCqNzx+2VCvAx5q/krxUJMqe8xqmUy
m+LHVXrdeK3d7UXjH2ZL1cuBEAF8l47DqPD5RF3+k+oIok3KGOMtTdixjacgJutp
bilbt+VSbR+G0yZSJVRpFcjkrZgX6GEJ1mazP6dzrqFonZovgMTkfPLfEfHcXdTw
jNkSwSa9WfDqKiDW1aOyJxBM7ovfVyL6n4n937hUu7xhfIMbTs993gnfCk1f3UPw
C8IFReSGzm977zrfCVhjFny1yhKTBybE+EbJPs5zzQVgJ0sbaN9A5R72z7U1Fh/A
6+NwsxmgVvVLBrLoV5dDTQk9x3cHETjYsxZCxF0YCF3KkM8T8JwiQKUQRSJwFkXl
JJ8PT2OdfPlOrzUKtSP3xbL+Ja8ULr2dL1j+JJEJ3j1XQqBCXjhq6kD4WXpZgaNo
aJnqwjOOfcHKc28Ag7ZfaT3UQGURuIDDSTYAm/jKiSwuiEmPyfDQl0XsNQR5XC1B
MuvWI03IbRmEoSP7Rad+V9lgnst5zZQ7zuCl0Wwi3GhhuNofowgFP3pe++25vAq9
nJ+fo+EfVNxBjMORxK3upeTeJQ6fCWNMUMYbqI1IyV+vMqAB5ldVYq6KO87C+6Ye
/4v9ss/3K681zJKY/tsHoSAvVoP4BvzvYClrJKtv3pJxBC0ULIDJad2F+3Psnv+e
c6NwmTQfI0L8ip48RbtkOfGDnpVoS4zOaJHyTnv9m8PtbJuZkG1LXOa4ur2JYLAO
nCMDGHYMBhLijZethdr75/+R9P9yYRYwjQI/nqvORqC+QnsQPFs9qxT3ln92z5jw
u+ia2VT0/8Cq64dEuAFPcaYXshEIVm41o7wegYQSqYusOnjFrqzwQ5mzFMe+B9qo
9autLRqjmCC6wHvnPO9EBmUL81Lz5GTYITreO1lXTv/AqHSMnJjMejcuvkgSl9pY
BfTQ7BO9uLkI0ovTSYA7J/ikIcmt2+d83PZMFUIIZBe8tGcW/rRQGNfYUISNcEa3
+zOMM8RWe9UFRPgCsulPJaKwanvkYZ4314OwB/OWdtEBjnpg9ZdPZXPh5qNaeENz
CQr0/0eAOtKtEN8+eudKyYy1wzN+TOvox03sgxeGI3hLS6hzeTGzbtTPOD43wFaE
iBBHvQq2xFQDXcx41pIDmMagSEwvN5mNhERoquEywefXdxnWEdfqLAd3vMgozkmJ
GiWRsDewDMNrHm/cuFmK5FRcWUVImMaCO28NqZVOB2FL+97amctEFRERQDmQ9yUI
FIOa3eJoQINjbBwkOdtLAnhJaq1ZUUD503X3mYCbvGwqtCPlray6ryVPGuetLiDu
NuwZ+e5ABXwoMV4QVtvoB6il48usMq+IegDX43KxHQSeqiG4vdN0PSKfBGH0YqLb
adWLjijiwAceN6S18LWLeDugKO4n92ubAxvl//YXphfbJ+JsWbNAtvK3xK2h9i6w
Ww+7ZzdVNjlLj1iWHBk2IY+Y4uDAZkRw62oV0zYsSQ8cPYPfCryRYXI/wcwZ8Jcj
GPHRnKLygpdH91GIlX2Sopy5GtBpuEke2IJ8xnN8J3PSx/xK/RDGSPIXUVuvjGVi
SJB2BtpsfwRWzUEvAijS3lHYujXs2uDRwF1HKH5SOWR2Z1M4UrkyNTSaGk0FbwVp
a1EXu70w4MK0TGCZrZgZPz1IaUx7cHe42XoY+WD7ucy5lKksuRV4Qt/UOC3thLxv
hYpiR/rlfp2fHQRTWd23fXvRBpU+oV2Upgc9eVFTSIEyfFbw6rhQujDDDkC87imH
6Xt+f4HYD+PI3hXfamtlm/uc6WISHPLESHhd8rftQF7qZYmyVXay+i59q3ndm8dD
6/tYM80M9JC2SW6/FzikzZiEAHE9V5w+rpLHxvzgjAtIuxng+hRafS2bzGhWf33b
WKs7uqE4r7OktX4vSSaH/ry3LxfJDk8ru7kdAPrFOqJW2yv0QeI13pRd8UmCNUq2
LB5cMles+FtUNYu2ItYYxaiqHsl9u3zmOrvEipqneUbszvCgxqO02s8b3LVdexNG
Y4b/eJfQ0uo0qbC+QVlOhX2T1vi246stTbDC774O9WIx+SMiTICAYIxIpYnxyRwD
8ugIJhuzhqYdlYcPfTPTP11zScH03dhXFxQj3rkJeVqmFCv5sXRWS2sozdxGvyye
5FY5cvqnHk7lbjof9g0cM2lZus97G8n7agHZIjACOAS1BNojXb/6DkbujX9sPuyN
7prU9Fi+lwqzhHW4Q3lTVxQz2Rm2U0EPEwQ1hmEoFKly30IPOWXGfCvXVH7ZnhNr
wPeAfiX/KS3C+2Qvlp2OH3aXX2dQxpm6KtIwnKOLJtYhoUj2s25u5U1uwBXiGdNt
KOk4r/lPSERLV3bqLTPUckk9BTB/wS6sQ8P6/m9TPcP0WC1n/yhisOyFDWvEAt/6
HBk5UtA7GXco/bHgM7ZXdfe50tF1aIM4BGZ+fShKkAb6nNHpD6ABVI98zZKBZPWW
gHwt2gEmFx+BPAXFRzhI5RXvk7zowr+XkZc1Pr8H24IW8nbjiSJ6oC9efxf3hjjv
JFtai70zL4BumR74HK7GE9T2fFyV9V8hj2EzMKoJZkfy4obdDslaKlmOYyQtqWX5
DoxlQG6667sF9BZcijYUzVOheBwsj2oIE4HWMQn0fYZrrIPoQp1BarsTMoIdH8dR
gczfhQ1kulBXVv/n5ddHZUHIyyc9Lm2OCO4kYoIIygF+Ybs6y/vJgc/6mpihEUtC
WmVxMrbP2Jxo+vZSQKnwmhLq/O5U/7LEWG9dfOyK4xlGbLTTII1Su2Bss30hXEPs
FbxP6a7zx3D7e1x4wnasfKtKAJJRqu3oWE4PRHD+cNnuxDqmu4kJI2oL+Kzol5fD
NNPyqgWnpX9Si9VtDjskKPjlNhHOEXPZ3uptDjsmwKvm2xaj7yHLPCSRA9fs7YN6
gIQ9CmzQd6KvDBUWW6J6ZV3E1S90K4trrDQg7YmT5Urt8XusNXPL8oY7md1YJdjC
twRgMd1X48tcpePAExkjo4kLmeurq0w2KhTcbF6nJGDqGB7VVy9edtBzu9dlJEbG
WILWX3OKJg27f2+jvf/hm/9Mj3nw4no07+Ta+7xIRK80E92jCxWY+jTAHtAsRDTk
zb124mKbAk7kB0QQOET5zpEOf49E2+O3H6hsZfik5gn4qTfchz4YdtPfbxdzWMDB
tjONIBORK+HfJ3a4x4PgzBHdt7ZPqcwmyHYX7cZnlJU6AEKIXlP+0TbOtIFJQr/l
oZNqxl8iAwW1o0hSRGYBGpHTjMewTuz7UJeG/tmwVcqDw3kfsqCwRIHIqAFXccJO
rISaso8B+I32CTfRvBHaf/S/WepYqzu48nYCo9K8v0lA+fzeQqQXISayTYp7Uaed
CVT6yBt/1s/SUsti9GbOWCrGyiAqgOdwVw2Lv4EKunXao41GomLqWvRPA7bkxmIp
CFnkq0hxgG59Fx4kSkzAI3NvxrWXnVzmgYPu8CsAM0qJgObpWHmWcN75TSIHTqMp
MJ9G+prQOWBqpVCBG47igZTwtlNyOyhkTk2/qMYIJlRuKGm4g4QHScZtE1rjCrF/
M1ZT80cmeUWzpmXJtMdTTj01O/CUHIjbV+5gQePMWNTAVOM7EFbLTSZYBZVLjpvJ
33SRExcaKoKsTZzL/FWL6WmWhHuGv7XIvHFEYNcLg2VaqAAnoMxp3e5f8dy+VB3z
n1g9xARO8GpjEer28FHyxuo/OAsYeq7CXsU4+IeaCL2sMpR7LzNcW/uFH61oyId/
t3GZy0+/Z/B19Vj5LIA/oD6eei0hfS9RlHPOhe1LQIZQMdShOqqck54Yg38fwQv5
sMqS9OUt2tct7x2uobtovlhOAv8KFrd0O+nbOrABwbPeN00OzRmsQDUJk+PjyriY
4aY+aI1R/iJ5CkZTWwPDUe2U0/8f4gV8UJT4kUwzbdoV0qm2/nYiZEWl7D7QQqsA
ttZI1KXbgOuPozdRWWDVQwo9993GipwT4xoBWw8pzbiCpH+tC1kF6ACjiqQ6z+Ft
BZptvdjdU6ZoIO9Tl7LIKObL96iCufROzel+JBTDCu520FZW3TwcUjXsz9CVViS9
QCcDvazG/Zne1d/Sdxf0IzIdzEM9G7Qo8Vqxd6WSNhWpshsIkF6gq+6a9XdZisH7
DHckiSPirf86Sbzv1P73MbIlfs3IjJrvCclYAVP8IqHi1STQFd+9dnmTRG6h8V+7
cKz0Y6iWGGk0vyyh/F4+D1NqjbzvhtgfObIr+KrNm7ngS3ujeVZEhvaGpnzngYsX
TV+pI3k+jQiHiFEfRbRHdJjcGncQe7BScZmEB9yva48vNawdu7v3EL1jNZy1v+/A
/V3Agwm5CvpHoc6t48yMXtCBswlLNOy9x3qXJHdYg0La6LhhgU1paYR/QiCaD9zB
pp8B/ONG/209ySx6+nnd5Lyaqo9aO3xd6ImUpnfiXNHO6oFNFVqEtczjcu1Gms+6
yYs2gdxGWR2LDdDA5s6o5O3DWkwsZ+bugqagsPGmJtbg8RIg7usHuPKUAHSQ6UXs
TPC5vdyklxoC8d1n+gKQ+VtIJbkMdVGxg5KoC+AKOK+mEHrG0I9Q6X+cukJXrLzY
98N2Yi3DtvTTmSvRCz9VywHLGueaCOZXO+pHjIrSzMJ6i+Y1SpUr94uSdhPJWEhP
UTTlWq4ugOcNzWiogquprM2V8BrCtziXPKtuIaYHv0TQJgvvM64eyOg+Z/Wy3lkK
E2h15xAOw8I1WL+UVQhS294kd6n8CwTC35T9v+xMqAcUR6jGpYHwp/d1AQKyJTOK
KH8TGWI2QsOS1+rbLucUmsWqCSwNIQZMZ9ilECvfNtHfALONsKmcyLB78sHgrkPt
sJjoUJ2iLkQf0dOokH3BLBvmJzuNOwtWdJcZU515Bwc/k3d+jqCpotBMk7Q8FMc2
gh02TokUwhaU5J4OgABvpwWwKpZvBfAqA0inBCTCI5sg6xE/7pj1Vy2Y6+3WXY40
Z4MBA+G2OeC6KpZXmaXjJepK/I91vvNxxOI9vHZrEf71dojcf22wrm6rrUPqFk82
mf9jG/y8aMo8iw+mfXP3OKLpfEtyApVs1c3hIXYIWSh/hcftqknR91yQWhjLZjZL
3MMjx38xCoBiCa8S+QIe9KpgpQJFe2rok4l37aRLkUhyVZFVl7sSV+fNghLvIiom
AcPrWUA0YQUA4MRS+7fh+wUAj5JF8gMjxgQ21kU9i18N/bnu7g0q7YDYAW5x33yi
NuCe2p8+7gmRC161lsBDNIgva6x6PIA0fzFqSjW7G3ZSrvDjc4uwkUqOo7a5sXX9
tpBgtalbjBVCvRnQ7qW24bn+p0Nlrj6cx5oMRpqvqEtT1bTFQKB4fvg75yFYtUTp
+G+ouNQ7kx+62eWiQLUqIRm7gDYCjGAvu6ru7qlDNgqJlIZH69E3BVgpqHhmaoMM
MZtx6I7GngQMuSJ9nGScttZ5No2xoR0ZXkEtV1R5gQd/yM1Ep913IwM9oZXNWFZh
dG2PBvPNVRA853W+49TvDALeLejMQrsgpH0laYDQ+r2LtlZtqId3hqUHBbir3GMx
4VyXOznCwcdXfYhMzL5OJC0jwRrAfTzThIwYFvl3/BJ9XScmo4AhhNku8fWjO3lm
6mQHHKGiQJ+UOeLIpGzsTpG/QR+wDLfOAq++BtU/fiOzI25ae6lvJtYG+NYlulYY
K4Ncd42vhiLQ8cGLWOQ0AOndkz35wugQspn9WrDig/K5z2jQKiGozDmnSmVntuu7
PBGresOXLSUkXYFv2kpbmdK3VrHP4LDZR8XGZ5ZtddebU8dmZDkIxv3Tr3xMJ4y9
s+ZWcXpsxkKtU3Uo5epxcuvOh7+5ujbwxHVOhI+nIxEVJ1xNcO0ffWeH3930Ntzi
yuQB72mwju42EofeAYUMCo57yYXzi44p3ZPBG21THGvMb7KFW3k8M3IJ9+cF8VJE
uFKXXNI4rMX5c1kJnrqAquMAYWXZuGBY7PnEcED0odEF+eEa6VuzTAg6hQZseo0y
VYwhQ3VlbLsFMXtSvnL7pYVE6Zuq/dAktKOHPDubn6Ak58VnggLoySGWXznd4/ZF
3GiGB+Gu0p29RYA2Wonn67oabbyh6mYW1xmmg2nru1F6HE1qdEoOkd3gQjyuU43v
eif+RDZPtMV+0+VVepzDXl5rC9Vmf6wDkQRiNE/E8xrFOqPsT96p8NFpgKC8aJ9i
6J8PquqLh5jrWkRbqErqF4yMywl1iFQuRYxwOujATuY59PTnF0aX1uXNFrJddAbv
/NkZM4z7ElQ/pHXQ0u7wPcB7ZW4FHwXIg3nI57vaysxV8il67jrPPfI/BmK8WjRe
FjS4gY2OAGphr4KHEtQUnucq3utTkTJgST7mSvYbccSFSWNd3YnoZZ6sDaduJsMr
+xGEk7rcPG2/Y58RFtjVGJ70AAn/a2ElR6Kwaf1mqLB7Jdh6fIwv/yHGTgBBZuyG
SlYPGoR+Z0skkiRFNhIPI7+0mCbT5am9RlxawGx/ZZws5a+2tRAsvFv5C6wZbn/G
dX/tupgJRe0nqrrFq9dN1zMKEB38cnXYDqlE5E57px1RnQtKLWrZQIIqNy4z1uMH
vkDlAPPXbeHvMy0iJPoHlJj0qVHF1NhBu4fp0F6X/n5qPVnWsQ7XHOWxT1qQsdUi
VH8kS4WmEBosF3MvbMLQe00E9jAIphPgpPOmo0yDpYJdt1tf70o3m6Nbbrmwo3+E
Yi8KNuWzVo2ObsavCTjPthpjqeDDuuBAM+xxYAEbE4x/LV8HKtWxG0dBSjdFlFoS
xdVARAFrCbmYoNI9BLC1v+DJORQYHxkKFuoticcjyRfpEUCxTzinLnRFpTNMDqaN
/pXZPZ78F6MSju6cBHcoSL0UXJDEyUIsmW66wYqSq74T9hkRIt7Kr1Bf4Om9VyGx
zWkKYwHWrmkyb8EX0VW61Mf8NGRTfQDZglQYJnidWmqMmczwvs91NuL8t8+Ah+f/
fZGuP7NQGz1QaKm5lK90qmMur/qLvCW3Vv3snL/aqVuygZDZoOr/kh5yuD0DNjgi
vpdibyZYJYBuONU5PXaRJbjMTTmV4Q3UTGnnxgXEELmVohTZavHgagGeRSEN7RTn
TPqiXgJ1eCuGi3YZJhIQpn1x67tIiXKvL3xiHaoV5sA/Yorzz+hcMR9zu9wQdPzV
/kxXdQ3Qx+QsEkHOCU+PLRRCb4q1qqBbumEADKefJkDXuvBAZkebBTCbyK/3moaD
5KFfYvbnlgG2SBvcHrjzq3ea+TSeytydcqCvwEucb21l8pg5j7hIqPKwiG4AeK99
8f0n6B6mBkLybga/X9EIiSsCdU2fbWrYpcMf6ulffryoI/ldASwhDKUXKkLeGnEN
4AkCitF4H5JoizhAVpRJtbCSGK981t4pYoxdh1ABXFQwO5SEOhFOV9amvp3Srxq7
XKdv+IA0wuwOG/aXCdyvzQc0ZoQJlhLpzQ78X8qRzd3BTOdkjAsxj+crkWb3F+UF
I25l+OOmBvGVhVO1ARc7injIfWaaO5AKSX4cgR8J+XqwM9+r3BUr/miKb5DTPN7H
96oAtmjj1X7zvcepLSbfjtmJgziMf6exT2wXviw/hQz05H6lR4+0a8XQkwvUnaLA
pwS0m5jTCR+ovsDk8AXMX9e1bU2TmQgiyk3O5aK1ugg890mPUro1ESCG5gntuoOk
V9KFB0ihvS3fhsoT1eVhv7GcZiEmziUmkD6TKZtdU7mZYE8wEZaUwYkUOPDlPXDZ
/BLVxgXzfOZ3Xntoabpp3tQXmuAHb/aD+NRzxjSNK4xtxmMnbSUH1+krHhWKoBlS
wttL7fW/m1cLvCyyouARwC3mAyLc18RQP6tASoR7d29oULTTkP35BGQFMXnk6ZdC
KW1vBQW3ZP0Ia5E7qnhgwwtIAN79UNNtQddQ+AeTn4szKaJ1FbpnrpdXzNhTebPk
bypGISMVJF4+S0tv6ILmeQ+BiLtFCbhqFT/bHkgPFU4AyFfNVhenKCTvbPtBuH9n
6a1p3RscswlgCiItGMeyBCy2jhHipcmluiEh8X1+bu6etcoF186ctEtcBoSb9qL2
ZIoI/18bTqPXszd867riNBlblKk11rLfdY+ou6JnoyMCgHc94bwzpne9OHOtcPUO
LozILteqxQxyAfH4GBVv/QB8wdb8Yk1/TktdvfNKJ+RmWAWscabFQLJUjkSDwnE9
H3cgEpAQqhL5Nu+olDsJ8m4ZWof2HHW0G+G398IhjTeTyin9WvC6qIkIp0jOVMCQ
ySNC7w47RerIjmdklS4OWdudLFKLrEE0XYO9YL9u5Jw7dGL5zVyPjjmMEOy38bvh
5AHcO+lzZLd+L4SFGbfo0As0aouowvBZ5N1zB7NlgF0yhVx3jJ1p9fXQhRdXVojh
8M3jkPsC6jXmlAeY+hrc/i8cuA22YSu420KPDl9RRruhbHf5hgcTX8vG7RQYxlWF
cb6lsaybA7lQMp6Si+OuJNxG+XfBKOCzxdQp19lTf4coLYeydsFYONimV7ZweOUZ
64bDRt0zvadI0AyKpz2DTdZrZiQId9Yl9ff3HhZOh4v+BSqbNxXp7bl9BpmGgi3V
seBzk9Le2Jrfv6eN/23wiUknQSyTyUQ1xggdQhmRXt11//A2qwkxsKvyB/1QO9Jx
W1zK6w/bY/XFD+vRChWSVd/GMzMcufPzDJ26jT2MWL77qV9amlnIA6JIoFRmSpVh
MCuJ/TFpcOvIAOvHyHFSlpkJs3COpf2x13wP3n6qMod5WxlSDpUPRDEnpjR22aDp
Fve6HLJVij69yWXF4ETSGbNYK6PYU1NfC1xcO58Nqt6GXGa/rbWAmOvGanBPEOpE
0RQoon1ExPm4JdVwufpX44uIizRbxtLlFvvHmodnzEBkCdHIlMiGDSPCSY4Q+WIC
XiffWZID0HEIuXUioMYwjeJxFMSd+8t7YXBQAn8Sm5fsQ2WXzxAMPUb96IqkVAG+
2+L6aaEYMzj+NgxhNRg8L0Xra9kyYHjTqbNExyg4sGeX5IppBjXGonAj7opVOpDC
PZPQQk69MSjG9dsNOTB+lHAkZkgIzGjnHVTO1FXSw7jJuVU986Jl+L0RV+nE6Hu2
x0OTQy6ZQm9dwDLZVGrF3LQWge3cG5w1NDMN4uqoP7RrxhnNs9GiOj8pgIeIyKVe
wyq/jP8FE5Ie8Sfd5zN5jja8yeAV39SNuDeB3cZbXZYhf25SXYr2gUWqGi8Eh2E6
k++6dU/AHvBpeuwg0BE86Xd0857sL+hW0DgxyzUYnxteihD/lRMcjgaS3OzRN084
J1cpmAoApBO+i/VOsdb483vTDbwFtZ0Z3JJ/3ThJjo9v8A5f00BZfmRpmf5P5zko
CQxHTrgmEdrJc94YGZ79M7F4x4qJ/Y9Hx6Kl/3WAcr5tlIDPmJVfm29C14sd04hN
aB3QPje7GHuQBgbuZGa8o1zyvwEUgJGuFgqff3To4xCWajSVi2opU45Th0SoIuFS
6iHRyyHSpABIsqARCI0LLbevyy97uLuAQ33yWkGeuIyUy1Yg1fYKZI8juLWFtSsG
Rhly8wtPQbLPw4mlySyyKdImjoDfPY3WrE7EzwbfbGKxkG4OwOcFcRFVJQtm/ElL
2hVJBNsQeDjd17KiMWRO3UE0C4hqCSGSVxp0eNr9aw1mIVoAUKjvFiB2lwlVvg48
pdyJVpmcf9o0PlAFz2FHGiE9zeB2lwe4RoSGxvC7mka/QtJ1GrZvGhkJSdQbVAln
B/YczErlYZwLasknhjU5wHEdANKWPSLeX8v6ZPg/MRCaabcc1HTf1SpDyV7ejjGY
OOVdaf7gzYL0vJMZ0Puv7CkKaMkMFYDx0H6Xa9JCoDmKYJcVwKt8TVubC72mq3cf
g/wQFAJi8bRzRpYTXhOooXEMMGmlkvzhvpbDIrIeR16/8zBBnnEh/oanR6CS7yR7
iK8GDV5NQFshqR5Qr8jvWZudYwrVqCVqH99YeHhZI+NasYXMLbfgIYhbaBwgI8q1
FSHuJ+hfNC+XiPuvYYH7+RIjYGxrlJWW8xbtsvny/4MG1n3DlgUD/f1ch2Gp1FwQ
YXKfmNXi+xs+u+KPVk2hiLrq044C7maKpLQa1NMRYxP43vMjPUFOwdvIXyAe8ds1
6FScEThcXb1erYMuF2GzGTegLrCxc9EWALjhxkiE53FaW69uvApfzdJUDSfJoumd
KY4G62hj7bwKhNc+QwiBADrmOjtOyUrPD+93iGO7fsZBjEZTTdIuvm7wIh2uB499
SmO9P6LY0AIfBBz3zeAiKEV7wDutiiYko0aTEGm4yTC3CEtDUzLTCuGW1jwSoLNg
cUEdAi/PAGAHOV/rOhiHuDdR7T8YtoNQI98mHhZxBbFJjsAAD7n53V7xw0E8nF6t
XO9f9EpGHZKA3N/t5CTIixdR03V3/3musA5IHhp4rQuml70pEcY2dbHXFDBMtd3Z
BOeL1/iwYMPTH5I7q8sD9XAVseClp9ohNhKZZ01toVoaxQw8gv78HBGSnQcEnnah
9K9YJKzwPCznzciJYaS4jUOUNY5M0C8YuSEEzakYYLjw1wiqLQ4tozhDk2s7okGx
iMVEq4LnatMl8mzz9VmFokW//NhpoRSdi1pxnxA86Piqgpw++MeRwqi18YGP38QM
7IhBCHdb5Gmng7eyPo2jWmxZqskB+PSX4mgk2UeohxaSNJ/YXE4xFWE4oVBV8aR5
5NN6LZF8y0omNXrIOK+Axx5DNEJDz4e99P+nMd31a7nbRnWP4bsTrGc4vU3gMFUN
wGRi5rMQ4U53Nw+u9FRzUs3YW5OeedHRh5rRnR+kuRkjBKf0QfM3KlI+3/rXwz/L
ITUAq/kY+YsAuXVQkNOOqebBXPrKHqdU5U3nOHuz6MZK+8ABVOeVnH+9QRlEEFjm
/bPGTvK3+J5JGzDCWq15hhgwypQMtfKbCyVHN7Rg6gZ17WkzhBjiTi/g4hQRN7QX
76GqWjNAKly0Kz6CVaicuKK6b9aM6ueBXgvIUBZI0rjVGoNGiL/tVmJKhofdjOcq
roxKtqb3nG74ardSOgtWvAHr4eI4wmvZZ8o6Oz+LMpSmlKxJhx3byfBya5UaXazh
1TEH3l6yGij1OpmFjvChVV5dEWQquW05584WaDGPd+WX7AvT3QwZ1cVzNKFoGp/V
o5zYe4R4ICIzSR99wmuGzUk93arqComCLklnorADy3DTUBO4ID5ic5V1dNBhu60u
dp2m6eFiNUutDEVxP8kk2qpkBAisBqSnZy0eG1IW0dslkK5QMWc7Xzkvet5iNBJK
P8ca7a53MdeicoqpSuxoMfbCcxbshWDxTw6TX89ECxLdiEw6TCtmKTri6FKWaaCX
xp2aPu+jTJAJCilhedGZtm0OCscFIdib2oiDEvy2S4A31Im3Yf9XrOTf6ofjPjTv
trL1JOWX0HDjAe7GKGTIZJ/bNZ+OzIYYRuSWfS3EEdmfuGLM/ifoqcpeSHP4UT7S
bInVzo/hBeC/jFEQVdVt8CrnyvjA/MMcDYK7sz1EGLqcxg0920y9zxO5K+AkLPJ4
b2LIDXv+46ay0mD8Z5ysY39fgUoS3ODcD1v+xmLaMR8bV7gCElqudzFWxwI+j/zy
A+MKxUm5Bcp8TCY051TBb5NRe03ugOXSoWDKICAuNwDcMhpmIeK8dQZxngfWXrtB
xefYu55UmFKtrlXWAY6dNWgvY9sIEQpTvQ++M9gj94B96nUc9sv8QTbWAxOlt7A7
xgNMf5imBt6+BQ8VvoHgBzqHBW/U/CK1pHczRn1ekkc3v8aXi7g7fgOvvMGpa+xX
1PmqocAlS0HtwEV1EAJw6iP7ujMLKwK9w8PBaE94MQnHnjXSwukn/zsnQ6OD/n7s
4wVSNiefQMI2+peMepeZOvX77GY+6Ztkdmxp7/EOBz+hzT9kcs2ainGN8Om8rujV
MpiWBGcNCnkK0ares8YfMkC5eYrtl5tz0b85YlZrBAka4MleyJJPj+UqTTqHVGZu
xKua4jfg8jnULsUJRi716QbCoDYwZXCFdKqXuiPRXjBs0qdDWkoWED8fHg7wzuKY
/eSkQo4Jo9/82i4ARRGk8P53JV2m8W1rz7V7T/wp2EKpWi4FnVqTf04WjJfoactp
GTE2uT1vdiz+QZM+IDGz/03xQK2XTNW+fkaHj3u+4IUEDHE39xiaxfxWWrkfuMfQ
HpzgD+E06LinDKI4zJbw22P0knenlooJrPaZiPyGbFlKLhHZUp6/qBySyy70UOyF
wk9EKdpw4KFE7DbUF95HKIx/nI2qbklMU1/4FYypboLJMq5eWjxegtjutgcZbofC
GG/l5PsZPIrqM7ObyQKJXa6gaGBAp9yiNZ1wb4JYMd0X2hPcy66la6sJ7BH3uiPG
FXBFP7RkEo8Gvezmu/dfaIe74VsLpSn7ZFKD1XDHiSmo22LUDGr+RJt0GprbpwUF
Cpt1UKs38hpspJhLe4cw5vDjBbHQyByF6qzr3+Wsx/BR+yaqAbhRz9lhoPlFknVX
RvjQLyXt89BPXiArzz6CyWjcE33nKKC4fEKeP78WsiqdEnKUpA10nL5FISDwlwUO
ELMUafNslZeC5wNIPxM+jd1xrDiS2XJ+bHjfyC7fN9caX3AQbLa8Lhd5Ou3wRroe
MgVCKo4Bb15IniA7CAV2ztsqbssrav/pMXoog471kGD9zEBn8T8+4q2+7nnsMFUo
EXw6VsfkUVT819zrQAuSGWhS9osYu6EazkOrScrcM8sqQupTK03zsgk1I/bx0XJN
Sv9evtljKQ207w5k3z9DwdsiU0EwDA31OqCc7HNdSG/YDEbl0xgx6e02mSo3ZN16
etfURIZmrMxqG8PkkZThnzP2/O5puevqVHW7EEqKRSCRcYPlZTMIs3G1gcXJdfBL
ID3+RNtah7mfaii6Eqt1tpQTb4BCleZG3KRAhGQ8rcjooJMj4rnGW9QcMAQOgSv8
PpPZGu645c/r04sUWwoa3Bsu2WjlLJ+HN87kZ68Pc067SRvKL7/a0ZwxvFkuu1Kl
sUiPHR5m2oIKTj2nhFEBSFIxVelUTbWelrqWu4QDU6JAZ0DVNMyh4+FQEuwOhgUU
W8BtCyLjQQmmHRxGh/0TiGlTo0RS5A8dvpuC43yCAKzXTfKB7VNznFvVDFPdtvdN
Xrha3ML0VETGdDlVtxNm/Nvpy/8f4oc9Aag6fVuUr4h3l3OFHPfRs6sQ9ErR/sLV
hyyY5o04cXXv2l+CypOoxQwq1vbNzycFcN+B1vozgs1YX5JndcOe6gFkN2EWiF7P
Cuso3KB3jMgK+Twe9+Nw5s6+HKHOYSr4fAvBY6I0vEY14z9bcB+nrmutErCZXir4
6b4v69z8qxxWdjOMYsdJHP4ZIKFz6OOb0+t7hmKHpC8R6p35dwJi21oBVCpQFC37
M4+RhLLDyYjjgP4vvCSM5PB3SteY7lRAktn3ipP5qcrp0GZ8pHC/00k/C77jWIin
ew7x8zDnzeFJZrBH8T5L7Sfajbe+hhtCIWe2j4fAd7I4G3l9X5dG4Rn01AiSzIpY
0jLcaSzdx2K9W4+Vj5YW7BrufyffRHmOKeBUr5YrUTEpSZgcYebsBj2LPspAAU/H
bOg76xJMzlaEFus8QZhogy9be88/COG7TXiZH6X/a2Jof4sc/NyKfGcLD/S69mdS
Pyz9jYaJ9/QT+vopTvNvDRww+WgEJiBG/VY2TxT1Tyj4hfEBVVHsCQNovKFf57pg
TGocxOsMdgCVmdGv6Kg3Rh7s6FGIikWtBPwq1FAk1D0OB76lthTs/HF5WT1As/td
3mmQre4zx45MCUE+ss67q5+OS3s8L+w9+h2UIPpMec/J0Q7NSE9PAHvK6T9jDVob
pduxcyJkeyYcgGNn6MTz+IyUUgXC93Bj8xbz2GNv1+plMB8wf9acnU5H+908lAO+
eP3iaCwGO0d+LkPe4mJOVl2PvOdT89BbYb8DsPXsdIkfDiVDoXKYs8adqc+TpXfU
adDEWJitgQtUEV5s5bqxzZvTs+qrwo3jxDK3cZHFe/aWwyqv6ZRtM2tAZm+gMLM+
IlMkx4+FH+VRn4KdloZkov88Idi6iBYYFFSD1527gJd2TxU67MdcMKlS2U+sYKgq
2Kehr37i0M+vEvU/xXSpezk6Zr67XjSO+kVpykkUh1gFZCsVjcMSJcz6B/1skxuu
2FesPeD1Q3UrvBjHVu8e4/pZ+j1IKcL1UT99RNsCLinNlDL8KJOYJ4v5EEJubWkP
t8p/Wd5Tal80s4IZ6EDI566psRAr5D0168YyuG+tTUh0SmZNX4uFecy4f+JT4xWw
HSrgVHVEbEjJZ4K7Qm1xhtfMTZspmbO9F13WDCW4xNWUiERZopENAUGAhvltjeY7
GI9We17ONLHqRdXgFhRy3AL4Hmz/505xpFMkS8grQ5E9DJFY3QASDNQrjC6IakPD
HIVkYlNCMa8mgrZRufIeZkJKq+DlkOxyDaBm59PQ/Pzf3CnhxbeVCSiQKQgeMWTO
efR/BAG7UoBaDzb2TjO4poCxX5DjijMWGHU+7yT3eqdRCmuhVWCJRb3LjlN5/+RB
61CichMF7rZgD8Y4gGeBuYtsfl9MmBUIol0/P3/ZoYeDKRClHh7WJVP40AxaYSBa
7zcnsPxYVmIiM1HTTRPy2UTcAsyEFt7Bo7O6EOaAnrW/JjIUwvooeMDAOVOzBLU7
vtpdbX5hWfRbe1zWj/eH1cPBtlNUEs1qkgAjqLQoU+UpJBfPeFNWAV+bFdDt4XRE
0c0cUcblnzBvdw809ujzFrPcfCzH3olTSA4owu8WJRrPlkMSYNDOPtACYPQ53KJu
FQa4C1mKKDNpfoP+94fKvqR0vw/6u86vKp5KO5CTN9HU7G1spoijKzXkAmOJSsjX
41TJy1jAgtA5QZVx8GIXcmqQ77ccotqbel2d+W4geq8nLnMdF6I3ejWpFIpdRQuD
sVWoiHvpQzz6K4iEbrNrkg8KpjoIiFrYYB6QWLj046ZxS2Fl/xph5sY4EjqazHBK
lxPu+lJt36twUIx3paYYJ+2hLEk5ZuHqBXs34ReT+5yDkRDzCUUrkI0u7VVaDjCf
5nYcaGG3O6WtXySgOBJGcTgnfH/V2eVJFgzSztCByyRzRLQoXsgS7RM1+tCmK7PS
EzYfhGIk8477HP+0tCiAXxenTNzR41E40MS2k5WJ6c9ZBVN9Y0RZ1gxOLUlKNyi9
L8O2g6NyLllS9U7VHWy77p+4VXQBbMxAXK5pbUVl88MYDUl2dTvz3NaYx9KcD+tT
BEElthky1NLqmlQzdQZsRxUdtWMpiwKUynZqKxNX4O6kjh3+uOJbdylC++8lr8lB
uXQiIjAtn7oi4tz2eF5PcO0YMLVRrpWf+k9XoTDWoDF7+mY7vlbK0DDIGG9PvtsZ
SzIG1Bb1M6rupZNRxvnHulkC4eDM2rgAjsBS4LEtv4tRkh947Ppf7+GyfguETMyu
aEUdcHsKQ4YFOCLaeSgwKcV4PY//38JXVZ7DtNhwThA7UXTGIENG+I1r2hb0x/S5
TVpvosSApPKYF4APEU6sOkA0GQJc6f8G5HMJVjJ3gy8pwye/JzlF/9W9YIhWpqKk
CHHMX4dn0+O+sEUxtauohj294IQJOLp+cvFSjtfXm7yUbnXLxEdsnbgf7YfLjEXC
0IuowdciBwf6eZVEk58+4gDJqw7FnXDqeUr4XBpH1w42Ju5vBOV9IPt9sO3yXNX3
lQLX/Bz9suIxNdTx0RC1kYFiJRSkbysj0RArtW6E389o3C5YCQNEUoKseQ4mW9pI
yAIhnpn43Y6J2r1GRfDUgtk4WuaFcHRI/WhB5+fqdgeRnYEmp64xFgMMYkF0c4ey
+Yu1UigIv0Iw4MJIdwY1HMT7z0fneLAy+9z+uIWHle6meMdNV5ODBJPty/zoS/u/
iA1SYtjJedq2ZzDWSYKd0zGVVTq1FlwLEPphCfH2F1WG2FlH/C7WOeaz4BiPoAbv
z0X4iFFyw6vanlcBNw+YYRnwLFl00tBjCIIFl0uomEDhBN1vPz2u2wKV0bzcyFdz
V6tM4+XH2edUG9kIIMOtDsHYtjziUbxfasHZ8/C9PVffG/23h9Yd1Jgn+nDPXQur
dNbzm/Ct47A3KCxst85wa87JblFSI2W5AU6xf9qxLBxZntmxvXhH9ytIQdsnebpz
98lRUiOhSwJnWTnFXNXDyBJMNSULqpb9p70kGwvMWYBt6AsMhqdICqk6qvQ8OqqU
3mn7w7h4L2SyVZyq8K8qL2APpzkOMxzXE5HEf5ZCuIljrwI+lGPlGj9OvZX2jNfr
mt+v5b7mWDceFItg79Q72oidPeGMBixBvcY2z8imnlbTpyPgT40eiKN8PxOAGlP1
fv8C1eFzij1RMwWT80+yjO3TBRjOOIq5IZF7/jUJLqGKZOudQlLFDby+3oIs+aCL
dYx/n73Egz73JN8YeyifrV8yCs35dhVS3AQzE8L/N7xA1/Alz8Rr8HlgejzhI8cF
1lo6t4BglAuORNfHd/3vgmrnACpmeDR30JZ75/gskHLo9UpBk2A+h/Ygg10/kA3Y
uzRyHhi5OdXwzKRv7xnD2Brt7LSjcvFDvfpQc6ibabUzAofR2fubV7ZcQ3dKsW9+
KJi8ji9w4fiOpE9+FWNgEmaAE4ieaGOs+kyhvlLD3+/KGGwKTpgXiwxmoM7c6Fot
KZb7VJp+LjzqW4Sbwbh2BKf+Cg0AG3f93QX9fYZbdlA7WCKfT3nicVPOGwfn2wL9
O571nUGOPwU/5kMvZEIM5onSztlqG9yK+IC+otlJKE3zYWjz1x59FRprpcZNB7/6
6mMjBlJ392l0xXlu1K+anBUtwrYTInSbiqHIdm8a4ECoa6Zd7gcns7RMbxjLhqh+
Rg0/D0VcL+zLFrSJwxlzBSz3KYiZAp8ROhJtV8k4iBzr6gi0EDfnml5Da6kRTuOD
I6k1IbruS4kbcaBfDdVTUkkyldYIL6Wu/zquSTUImQBPjSxfjAQa4dkHbu9klI81
V87rWe3bFO1Srao+OREubtcWTHtgsL0/cladW6HG4RMs7rLnVqqWvsAa7nutigON
VLjIe4wQXai9ZjPW4zsdlxLgy0DpZTDcF2bMkpUXup5dUrUKo5ToOw29G3RvIK76
1SiA16qpJBrBCBKIr8cdPcxgGd1jwy+d3gH0jreU4MdY/x0WyE8NWSH5rIQiJWnB
W4JCvl/jdGp8JBrwU1oq+Uu9m/0jJLMbmFJLJQyWY9cxZ4bq/I8XGw69lGs5puZx
PlkoFD/wjqmN5F+UCzHUr66NiNV4aSI0J3vCDnGbFxC2ekl/BgVfXwtBl5YwFCIl
HGQs+9SHbUbyDr7HwoaqJK9QSg1Uw0ZTKiq1gxEIar3DlySTweQNLzHWYwCgFvGl
w+XMilOQwEmQSQP439DTkRoxUzQaVKds8g7jGI2EgL5S2OPgMMVXqkqQ5q9ofoBA
WcOtO1qBrGCO2xLhRyw28PG/Bn4sLCZqCI1RM0t8PFdFvfidFBwYc5xXagVS1UTl
TlW8xkIZpsUHIScPXRnjm/x2WBec7lCg6quH0R7Q6Fghnm6B+UlAE8EeYloGpC3Y
EhFhrOM/5sHhIpf8IKpHKG7Klr+f+jN/939rTrm/2q3OwQ6hf0nnQqISJBHLLC5O
lAPCq5jAHQpVx8dAU1he1Rf3tCN/TjoZ1W2iWQZFIXhNAzQQyo2ZcU5G6B2oGLPB
qHuIjqi31GYByWGWRSKFBrnsG2ENRCo9rnUYu83SQOpfUQApJplwXYufxc+tidgt
7tg/Qigj04IAR5dPeYb/en+s0A9Gfz+k8BnpLjHahYeDMwdO5y0qjJ2BF5HN6G82
5nfAWHBywGg3EqYfaPExob3k0jLhfOH3TMEHxQOEdDEpPsk2OwG3Dw9oK2hUGRdf
O/pVUO0C37pRy1ZnSKh5euQuT3ZDuWYWrWdWngFL6IJhRA8fIguE5jtIMN6h5Ns6
FpsTNTOG+mrezr5w9ABjcgtoyRiPLpYQg7RpHLsdK12rnRIPREyb0cJbioXn0u4+
kHdLFqkpR0XtY8flE6vllMjKv8XW6ZHi2oMwebPOiXZFgrOLYMoA/THYanqvAPpP
g+R/xnbXncTLAW8FynNLniK1RNMHsAo6nuPl51rcF/Bf5rtKt6wygO/EcXx9wR9P
ZUj0jSmKxkcADdsFWMfP9NZW/H+4qsJd04tpNqBFwjyuDcrldA40RbJe2m7pARO+
M3eQgFPtu3PKTBafELU4EqxttqbuIE6b6HYygYZ0zM5TXxhcJFOsw+pBeHUrtXIk
5zxeURbbZnE0pRwt6V9sXqYdZA5sGBIr9gBr34W7tjXGGZ9Cw+PB7dUqGK5kxVfF
cwySHwzwmwqQ95qOBDfLwDt1M3CSP4IBBKHUsWlMBRugEWO983D4L6gIUOg+gyHi
g9s3ZEKB+f/SUW6/zlrsOdbaA+QmdvyGj4am7D/KqRvpI/ojv5JO7TqNz58ZM3m3
1wEK605SqsKL80je+lm7coDc8H+6t9Mzf2Wy4c9I2z7YJetADRNR3is2kbte4cz5
4jEBWpS9hxPVmKkxUL2s7DjhDmQOmMsF7VtoumPL4uKHv3ymvxjL0a4sXcZfSgX8
GXvFJ0Eb/pzSzANv9L3Necvc8ESnwJ1Rv+V8gKfSedBTOO7DpbDcadoqUDfSxZ4Q
G4D3/CSdFjVwZAAYa8lnE28eZ+8N3WUM7WRNUu9bvd89RfOSrGSCk4knWg1sAb3J
ApqAijBE/s7NJZOVrdCvKez5dCEc90atTlM95jkV9WpiK0CoH5J3BrhtFBO4F14p
U6rNQpCHpUeLUf3lLvYZ9USv2SoQa6Wd5S/8+wyCN7UG/P3yH26B9S3FL/X0YlxY
8EndF35xgBRHGSwucQb++lQMuLIVU17U/6owUCoQ87pfoo3GkZVWWPT/CSWbtTkF
kAL4wDXoL/Ke1ZRsw3emmARAw3P6zIcIaiZktJhgfGcNwFGmhNdF/QY9pUhvpVw6
wkHA30GxLeYvBqJE0OCaMI9nOh/deeXhGsJ3Y7wkujZwQjFZU7BuhjDiqk0IkuUz
z37qFNnWK0UWZj8z9A+11slOfjyDEn0rcZuuanzHgjL2AWrgzjiRnbwh8SQqmnYk
Tdd61xAs49kP5ipSF9YYWnAMK0nXur0lCUxynnuWXlqVmTfY1r3WY/OxpjhldS7u
lB7NJBQhBLsgCBw5LxuEKeZWe3/1gGIMzYkFcglCnb0P9hfeR4qWea2NTdi9T1o5
4qMvzRYa/f/QiQGVybGYUYWXFnLVBNdQC8emFhySGGMKohNvWGX106Qls/jzqZc6
FjpFbpQpkkClfJ8DxlzqN90ms3MPmGf24sbBP3jGBqcREY7o+MT0DA8hx6BztR0e
gzg4IrV0kNsLjqVVQPyPrCzSMPu7NtKlRcf2g5YJyuRmqLFwKLBCV8fwGRvuzCo6
fQ23bQSRmKN1DZacXhHFANwmU6kW2W1+vn1lx6tESQLkvN1kthERAkvuont+pd62
/AoRT+UbJ8By3nVcB5ECzl4yZxW6zb1gTPAIFMMgDUoXuaITDdtjt6x0oQjoKnZ6
N0sfhE42oc01AzHjLpTzaOYslfEPD7dvm/aw5TQNgi087Vec0ihlwX4a7GMqmjfB
yfbygUoD0M8G+zJgJZNzaP0lgjNQh9dG5BwQ1wOGBYXLYMUuQ7jRkh7AkJmGkmo/
U6UpeMH8mCwmN4piPqsvjjQF0jTWpQB7L273TJioT3qT9bsVHM6pFU6U+d5FtOcL
VNPbkBcJ6oO7+MOXKyZTCfDMMmbL07JRPerYAkfNa2ZsJ1N2NGgP+RakumASaJhe
TGzPNsB+xHdMCP+j9ycz8Gto9on0CXwzCCi4vd7SIUbqDQ+iu+0mLwzXfwPHwi6H
4n5i2FYGiHq0DNeV8VqPWh6EJ7Zq0IggQYnwY1u15lYwmm9ShbNIAyVo3Z4lZkLW
duwVmfVzf6V9hb05syuRxrk5Ima6gsk/Bby/ufCSz+0aZVeegQHdOtwLK118oV6I
cxZ065t4MyJV9HR9x7BGVEGlZoax3hIcz//wnB25RF0mCsE1M4DMjMHY3ZuWHxQP
cP5ByaGcmmZXT41CmiCYrfW8FVpqPFTjNm/si5RBGQbl/AIT94ReQxo3mCMtPv64
9GifsSs2UEE2SG9u7DU8vT8goBg6lJpcPBzZeqUcF0hSB/utMmpwMFbB7rbV9krl
LAU5pxde/fN6uL2sij5tuVbJVmOmjNzvbp2eCe49v1hYVZYHjm9j2flDE1gdRsBw
lXpM9T4oeSRlVVohaHdXkzGyBQaOaDTbHIF9TvBLoXpu5KFznyhAKjfbG4/h7JFC
VZxwYtVado26tmyaxi1bFdCVFefCW3vXB3Hmt73MTo1CQa/PrkXjt45MTbRWw1Zj
z8N4XwiqVpz/69Br9BJK0sMijE7DBogYcXISO8pWZNSI+9TBxCuE94xs22UlMHrS
sauBMo/0BG05FWOVlpQE7JcqnQWK3cfrfq70l4CFoYEmgYAeTmdmoZ7RDprUV1y/
MQYE+47HFM2lr4I3uPXCkTnxhFCHRhBofR5izpG4CBTH48pCRzrvG+IkT9hSAVMV
qEJU7+bkqmOVBkghgvVcuxWQecj+AxqmvvYcxxcDyzmsxEMuoiPv7h2CZRZQAaBf
C4snmMQalJkHP0AwDgWbKqdaYvmbdJtViqmExpfMYQBTlIB+3yZ6FwB2KW9lP9Ru
GgwMsnc6809awJY/8EJPKpy+qO+H7AlkcVZOgmPijTg7cRdWecjs2Jlgt9QSa78b
IgplAhBTIu+ZCScPXN5R0HMgAo5qq891rIutU6tWngFaLEBAV0Lcarhg3eGzeP5Q
uPukN+LbYUmItwN6zh7++D9kFuu9K8Qo1YCbNetusllBlnfwZlAXzA8cIeh6/Bpc
1A/FKOp1qv2+By8A/m793MsEuFg3voj489nVw1ExRChsUV2zF++CcYkwGL2Y/VNa
HVpWvMSsRpwoblwhG287RA1/HraX1lPcQ1NQrahuxTioTpD0WFsj2wdhUPHpFFCF
d8GTAgmHKxTHSk4crxp7VzOl66OYntmTGu7xF/lhYOpvMtNrgd8hlJfBjx3a7a9W
nfYAICTisj1chL7fmqqvCyq+puE0wIH+UtHV+1rC4xvrW/GBNxbBV0D8fr9d2Oh6
OB3Yro9VU+Y3JRVSH0I1by8IUT/W2DwogObbefiw45tN5TJWdeCnd6Y2CGAPqSSc
bQxUNxTdO7mV4xEC2KJ6Kve+SRHbd9E1bsHKYXlSGfKlTSdc2JNq5vO6iDtJVx+z
XzgjaZY/Zfo75IM0scLS6oA1N4TxKBqVaD5tmYVSoysVG72bauFXGGuUVUjdccS0
hnF/YRRI7KZj2kiGMDD3AF9+5JvQMn2Onz5d1UJSo3r5Bb8DevSj66F2512tVuh9
khBiFbKwAI58nh7SKhpiEiFC+9dfRSJwXxEkHmLi9tYqj+iBvLKm/CbPqwNIRRoU
CUiHMdl0SyG9/KAdlP95YaNR84oxeI7siOo0TYv1Lnc3HvOUsV2wiRAMSAqCOT6N
KQ4EX5m/YrliqnBGHjHed/W1X/k2Bn1Yb+lMF/LF9O/vh5RJPSWQ3Of2oo0Q3uW+
PnwvusyC/o9LK80lbg+sCEM9W/tPVGAeJJVGRQ1t/e5P1NF7t+4z1uzihRjrvbtf
BFXWd7pqi44VQ4dsFy/Y2HR6WvZKec9x8dtcuhf3Jhom0m9FbKmdwyFHSahTp6Ur
IYyhTforeBXL4vxzdFjFtM77cPn3NoOyuklKstM4MIZoCT/60JWGivFOMJQb57uj
q40awfFc6z4fhIfMAp84lhyjGKYd0or7YvXgbRwJDuffXJ0myaVQLW0ZCz1xnf5B
TfIfm1x/OUttjpd7aRQ1USR7llxlUDCy1laWfGvAXbLMHpoN5680nAH3CHIzZ3I0
9Z4mgiRh2G8m6imGfrYH+QWmOdBK5+UkBYKZXHEcUjxF576x5231z2UFA4S31+ak
E1Oom/xPHueHgVU4y8N97CQUm0c5JNkTP/TJ5fgZVueDXvRGRsjTEBuqJ6e+FBPJ
s1038IzGRmaBckvuOlaUUKGXKeALz9XgLQPOJX+MxdE6UIzPbE+vx1HbEoCrEXRC
sed5uRoysTitbngEhyMxSTcFTjsbvKTB7Y0V/TeqOBeG4sdPaJD2N5SEx+bGodEg
u8mg2TdhPYSOljUVjLZHAonPR03pA1rDDdM3qo3/NMhjFYzndcr685gL5d+Iw/iX
xddPBvXl7dEdSiS8T8l+1GdHIVqKfzngUQd6OKJ1/4UpwzLiTfKyAph8BpsRWXmq
CQq7pADRMjvMdgce9ifwM9DDkX/83kFtIJfTZfzUoA7PXoRuDyYDsx0Uz9RbHJsx
h0j1C7HQUane6JZ1vTtkt9NV82JmYeL7mjQXmnVt0mt2qZUruTO4Pzx2Zv/qaJJQ
SoruIt6r06uLSqbaSilvZVUfWykN37W+B5BlMYRY8rDauAU2Gi07gLa/h9s2beVk
oxYacICV2R2z2CeBSfg+dblyntDh6xguOhGXSlynvNh6aQaafO48TzYbITw7TwZ2
CLo2bwaKDT7t6igFTA1BXaiZDqU9xEmsjxkT5LMSCu+Zk/k72O+pACZ0gPn7+ZaV
GZlgiRtFzdXxqQBo/4TvTz7gnjQd4WgTsrSkFvZcjW6iHckyUE7TGW4ob0iAC1uG
gv8bEAnKaudhq5qv9h2MeRrvOtGHMVY6nOwCxYBl/jvXxmVz1TKhy9XafU3Zqr5x
wLZEWizvqZ1uBNhMyPuZuuz0KfzQza/DNLg5QboiCM95bjV9JqhTljKZydcpU05l
ELBxDK/s2anCKEeSA66QbydRcDNx9IEB1B8DRGM5QpYbl4T5ggEVtHd+5Msp+A/r
Rmf6KqqucBIysDmdHqcHkTdkpuYmeYlRMy981RMg4cs9Kph5Je6tzToTzFenUKjE
81FgFPoIyYO+t+nLF2VCLGgBVgW/b4mADVnT21+hBve5PX+RLuN1IHGtDSY+7QI0
KXL6toVI+Tk1HVPQ7m6P1AR2rWpdkQMCuYvnSeGzwM3AS17lydY00FfQdf3nTyXZ
72oo/9gVPyODcuiGagH+nuWZYH7jLLPeopAuUkKj8b1lAvoHqc9PC6UVVc6Ii+x6
0RfJ/Wn7B5aZxXUjSDeZEfNoPQ9lwA6+6CYUj4OBM11RXkTJyzp+qR3e1T3rlzBK
8/ydbMohvTD6/7kJKQ1miHhKM6wBiqs+IUEPknYW4dSLIZsSqh8h/W4fb79DrK/5
EPOuFvXxWwdW+APBCLG2BTE/Dth3TgVlvSqi5QwvYASAkCBI7xVWwRSVJLAoYOlF
9TBnQifg7eFdW14+57+fLaWteCTiMKFNfc4bN3az5lH5zs/TqzLH8PrUZfjMRXPX
4e1VS20UbJHF7wpywBixMs0X104yF3PkO1VDwK0MSmoXwkhrBPsXmd6iynh+kza4
XKnqRF/6NVMrO+0R/HoRgZC/MfeYAcYFVy1KE2cjLB7LaLJht0Gih77jIAMAKuDM
dCyzOSOsWaZaHuFmnXJbk2BboT6Cu93qO4cksFhL+qFeyT4Qh6EYB/t+6lJ+qMTI
ZATKi3tBzDPovGkexUzb8b3ec7W0hdo8JIg0HYqAhkk35PHsE1Lt3yLP94QfrGwm
wF2IUfCxesgxksmYnin9A6zAwkCPsXDiyyVw3Hi2nloRfbjN5p0VntQj6IPgPbMf
byjV8t7DQNRkBRykPTKWZ/XLK2iq5Mgo6TiC2BXUZ3YxIebk96j35PiC0imhF58Y
WCEZVgOC35YAYbbx06A7qPLR7LHVTOtKCfaDqmK4cOgMlmHjfN0ojMaSgJRDxmMt
5y37FwWCW5xf50TGezQlqL7y9CLF6MxwvliWV4VWqGeJ2KXRGU6g/Jmw6I3WRIvZ
2+53iDEFlAvC26hsu7+RRE7j2SyOKd0BN8PkwYrKrP49iu1idr8XVFT7UEkNKV6r
+Y5aYkmb1TmrfPCVOyjwSSyiQkREekY8eAu3DIoE2iFFcmE+EkBvAimqe1Cjp2f4
tIFsaVWu9KoJElmBBX/ejkNcXlKO2XJl8sVE7WXhpk38Lu+8lMa/TDK08hXPvaxo
CzC4jxfdYFLOWeytKSYl1xwg6VjzDWnTQJQo7OAOYyhafw+XVUtos4Ny5qjP1f+v
i5/70jiT4Hd8k2Dn4CbpRW7oVH2OjGlUpEqU9AB3jMnPUz+2tzsVqmO+w7pqAWTx
9h93ZyEf/VwzxAfDYfH4Trr2o7RU77gc5YbaAEnRAYJtHcw1hFQomUoZJc3Q318N
CNIvLQGfhKqHGGR22FJsY+hUjKiqOve8CeRknlcyCIH2PUXDy/QFx5WNhBLXtVkf
aAKpWWAzegTC42c9jZ6nlZ2JD7Y6I2WpYHM9g0cuqfrVfL9xX4goFKWbhq3Gybtf
c/29FD/B7xPMgx3w924Xyq7/fDWOfjaww1MpkFFGks7IDg+bR5awrY4aSW2SVRE2
MWdU1Dqnz1Nm3od8urKAix7qglR2XE9PfNJsdyFGw6RnvIsQdmhXpkdAgC5k0Ui+
ieeCJIx5RhhV/2W7H3juUHJ8opYyqWKVt+XmMCxcC7HBiOD/xFOnR+ioH8XRKLo6
kxN0Dre2zcbSDjG3JWZvKWxKZWpTM9wbVOjJBh1qLl71xBKnxdm/VdoJqZILJEoB
wHYRHXx4x0rnU1V64Xf5vaih3jV5UC3qoxwosqjK+V7ruSw/NBL4DV31ziny3gMC
HoPrrQhCjpapSPlHdXubj0gwxZy9IrLWQ1W51E+gnirB92XZRjUgjQVNrZMyCh0L
8DEk/RuLFB8QIY64I9zHtb5BLU/Hyi/QLMkF06YXtr60157MUx4v7f095drqSfHB
nEH/3LUk25ei9Mp7qFtLLrfApGev+4XW679A/RnmVXVlpNa1lZfGk4JUHDWMmfLd
42fCcQPHsW6yjQ1N/9DI0OZ3bUbmEvQjXcz2AvRMGTj7iowGiquE2uhl2BSVx8qT
4XE90r84R6cQnGx45sDrrsVV+xFT4CK6tDShASw8CDGRHtxGSIYBNyOoQu3xhvjd
SHhRic2NVpbUzwviYA5kSXQmhCH/0MGUY1ikm0sOCQMONhmAEUHbkdJUcvY+3pa4
ECC06NKIkYJUnwPXEgvXbF8LsombyGVxM+dnUJ+i57UAjgC4rqWIkQk1g0+0obJv
1J4kzcHNUqz9G70STmkXICx4DWMEQ5KEYsiSVj/NWAUrQjXQfGexTJWgKXWG7ZMU
zrrPJJKcbZmvQcnbKjs9OUfXP5pbEWLMenvDgT8oQL4N0IyNWXhGq7c2rwD1hMbc
4Q8Qe6QwgwSBI+hPSyek/XJVste37UqeJ7x3apDaqhGvHaEv220QiNzU6L0bHf3o
GWh8ht6ZGm76ppoNSq7nDweY+irNiGvtUU2GfD0HWUonbKU7g5q6tykI1bumY62O
45KP4Zaeu0JfaMKk7xj3tq5n6YFjtmAZ85beE4RkuqfHI5jQywi1Wu+xQcZ5fTVv
eLgejg321JGxG2/DUeuw9SYhwT/2PGf69drUywaG/Q18idRSulqPYXUTZUp0tJ9r
BBg2B4JxtiwjRgmRhQIvRTwu8asE/PazzDS6Nm5mgvboZy4opo2Vytc9BGtakgM7
ZZtSokVoAGQpjxKxbtBuKuJP2qGXX+m4riHgoMm2wnk4T6RQPfV2LmvIhv9PkEgD
tsCGem30gBXQZIB/szKCgtIxIA+gPAs3FFULX0DUCkPVNNeSZf44tpGUFa8CiwWQ
DaSw1RACcNUzaWTyG7x4RBAK9ewiGO5Kl3NJDQpT//zcv9MVNzg0ZhKFLO3AwC1u
jSv12hpAxX1+lMrpN0lfWGoQ4THtvkV7ci+tmFvG61WGsDV1emAK+DlqwbbK7WVl
2z2yiKdyAJ4letlbwQOck+EU2s+BLiaCkoqu1TYrSTsf8Pdpz4/J0nZnrnVpaOuR
jfRteK7sbT4KBSdUKue7xAJQi6+UZQvQ3WlNVguQXHwlpkxmUSBRpOWO1RiFYrjb
hQ7D8pRywIyoOlBauSc0P8v4pCQsVZ1a7LPBXqK/hhLVujyiZ2/3WffVqm8iQ0Fx
3u0974o7kN1TtLqHygFwQgcVmsJ4k6GJKTID12HEDEmr9/DvSQOvI7NFhwuP1RCv
jj7Gquu7eK33iS1RfhuP8lpoOtaQZkiNUkq2j0kG4MY+RsBJej8KM9TmbH0WYo4K
WYYv6tehfc2tDb9QIstGMq6WULAQ6ZIdZXpYob4hB8dsF4cjSbMIj7v+uM4HBKs9
IZn8Q23prRUZ53RmbgxXTjQlRm/AdMvNQr+HjuTglhtWBttQ+DlfiUqpdIA6HH8C
ZymuW4ochCUx9lYhsQ4pZHcz6LFma6H5AX24jVrIc4D92LmhWzkYnldnl0WcqYfq
KqwZoJjzU6KasSOHf3J+Pd6TmZACIxZm1WiMFVPabmqWxwcIP1EYBej3R6LlpPHi
t4WrRW8ewSlJWzEzUIWHTTZFYYalxvBzzezucyAeFjWNHu2tiRqwYdiKrVtomdmK
hzNsTQKVJiBCwSJ/7L2JJ404/qndE7b/03zsmQJASEL8xvNnrQWMRGc8LiPDh3LK
w1Digqw07P/tnVDrYkRI7TSbremt8RZQOMCd+aP+wHE43zl8TVhVRO2HaQ4GV/D4
sAAsQdoZVVqIM206kYKHgCj3iChHZtcMS6BHa+63GktDILizZhJx1DxZkNSBv4ht
6Txp0g09go9u13YQOj9bE5fE6NxGOR+P7tWGqaqccUJjnN1JbRj2vF6gByk0kFOh
EEvY53QlFcj05HPO0Na09+EsRM4PIvUA+AYQkKefr35I3vKRDJOxoNciIdB5oCkc
en6TMVw08T4DUxIB3VVj7RvNasm37k5Ucxu6reWoV1pkaA3rtLqY+E4rApUicjb/
6dLrTptGOYrpY6VpAOuwdUq4VzFPDefiqVnKMTiRpO/WtubR+n5NHmmLPuaAitkN
ljpYof0hKTG4OmSQkwaoquSG4kWFOvnOujTCkMqgJX4xMTdMMhKdNc7G+fXYpt/U
XkDAN9ygQdI8nHUOgOIXOsPH4Qwd6td6IgcFP3ZA+VIZC35ovkVL4EPBoI/vSi5D
oKQLBqqCN+nV081lwIze1GB82X57eUqfjX0f9cDqRWg/qmiBaK7Ed0G3LUcl1v2k
DIIgJcTo2U0NbjAEYewCqwTAWfRtXn/geoQgHYQmEWfu9udNJW9QXOI9Qrzs5jXf
GLDzUm+vn/Uh2du3jRtBig6bNSbm0HGHWSQcq232NI/bJ0Rc8N9emlW/RkyLORvv
8i1n+L03aY7IsQLdarFXyHv8lrEatMX2WIGpUL+g5Cwx5ohXxt5VLOTPXeUMlKo2
sWPgFQ3/KbVRv0xVPfgJ9fOY1wnMj9/2nm3nzoPxfJ/p38azP7GWETjVLetw4MyH
Y64lsPBozgE3MQeDWNWAWQL5WcTNi+6B/5MwZaiFpOjYn4xZb4BVZWoErnPXAbc3
RJQQalLDEIMv4NfJkF4YPfOOezuy7dLhyuw7QyPU9t1eUg5gXhHhfVTyR++34sH8
HUHjRbwNkBCKw0Sa8kv9wS7ywN9j0r+rwW4usLJ4KIq0h+PAqmcZ8W6vLVhbp1sa
WG8wjB0uBZ1wZ/6pBM17H70+Z2lEmU57Ff1ndufHw83zc9j0i99k9qcAXXmhnWZ+
wQd262e1m3sQbHHZefHHRL67fTaGa3Pia/BfYRTwxF3b37Ak3swyqolOHVU0hmjI
08g5+wVEMPI7NYHSQyCaVxpCHJbKO7+t9bKg9xeFu/qbyX+Yp/6MCVNaC8oUHnFR
g+KvdulFo/OZvxWQw/pITgvxetTLquejAJyYa4+lNGdy2v85HTjRGG0x1s629lJi
HGvCmE1i9XRc3YHTw2u0oO3wr+QT25V0BBTWGgZeDBayluZImgqn3p7i3OOPrC5X
ID8DH7IATdttZNjFXZv60Y+aJdJ0E36wD7qSnkS8jCwyHSVxdXrc9ydCI6zBsOqD
h4i7e4Hbh+LkN2jySDFdtFAT/iVphbKZjkrmllngnJ8e5oErNcZhgR9tVeCUy7Ub
PpGR+SOb8YI7VvYKER3nneCNy8MFqUA80RAAss1vNp26bWCGtUCf0ZgO3n62oG5V
TKadjY6kjSwiT5mNbsN66wDtEGo/jbNU/ZwogBmK8a8mHVboeFBzegXnnh8uyjOc
96/vY1Jax4OkVae1PhQlDIQ2eIJOliuLOOjFXtZyVaKiyErdUphJXnGySU0pLcLK
VO1od/PSvVaiHXMfmqAZWzQyvV9C85HGcRIrngjtR24oRgf4gtCnCmm96GO64Pn2
pjlLz/5tmpmBRQ4VXV1dLrYS7kQGwvhQcYADdDFmLLz2YRznMaz7p2FuDccKmdIf
Cl/dUsWcogUfkHaYKjJT/lZzc4Y5kwHFHP3C+4rahAE+DcNrfU8dtuIFLjj9fiqE
rR/XXJoV1QwA3eaO9ykPzNrgmG7NEnzorspFTS3lCiNUJtZvyZdQ9R0Rdkvr9Pep
DUUO5l1sl/zrYOZasFEMRQcwcFNF/fdV3PbL46SWo7OCPX9u41fxkTA7T7t/v9iS
quduUPGI0x5K9qLJCs3AReTwcpIPRKEmbCre9Ttd77jetp1yaz9bLgq9IUpjTA04
T1FUIxSwOV2OX4b5+qx5p6BQwIMjEBR6564EOYkXbu0yPzXSBNQqd5YMmcv+44Ks
6BHWGYUkRCdPPi6pTS4TXeWXbQLySajA15CFb/PWKvirg6RLh8OxMTWSHsPGMRpD
Ugy6xGCDS1VpXYhJL8GDCU24hwVHUR8WA4JSQ19esxSvRMhKGuO/CqvWKHCMsrlH
oIuSAqCUvKGW4wz82QfKDiavAlWNiNDFM4DNUZgO7rzHBmQj8zF5ORCD6cdu0tFh
vP5WEnwcr6itOL9Za7iDElOTg4wdHTH6TXickSOa0HNvHS9nnBHu28Goip7pMCj4
5nESUQHuBlLcJcE/6N9Oydm3v1MISH7sEPVwcTdrhx1XtF6fTf8pQmZR1HuGGck/
DmEKOe9NhYfqakxIjZ2Jf2cq8Q8GXdJNfsfnMJMd7W9Ojcj4EQx2r6+vBxxT9FHS
e8qYctkTkNsFApx7PpTQDNWaMupORz6zY1oHhA2LINxIYzD0MR9pvxNeAmBtjHo9
atFZVTuKcIMTnRhC3f6XYiWtv+XVCr2CLd1cAG7VwnaoSYuECBPf8S7Oy9+nAyvD
Ojw/UxWYM5QzTP+3IkRShNoe8tK5JE5scYCveKhT+8rcJsphZteAxa8EOXvsE8+W
Ary91NH3Y0WiwA5ZZsuwcPWx+P7sOOM1tLAF/jCKDKHfgQtGPSA0bxpc7pmNegEq
gyobXUlI9uv+cfUWrpNPm84W6wTks7D3PQ8Lc8bDWi2y6ADQKMiclr04tF/cau8O
dm2Bhuly+KnJy4/q66frrpBamK0Uz39v3g2aGOSmzSZaMuwQjcdrDa5ubkF1btfT
VhuPChbyOG/K0YsU407W6d8oW/lNCqJPSbn8axnQHBQjgKE6ZIBt0BSoEW+sTDyh
vw2fL1JWCY4a/8zwNn2FizP4nMelbYcRkf8zj8gXm8uNnuFJWSV3GsWm8gNW3sEX
0xGUz8NtG5wL36FEEpo2c1tTPXF0GO5taujlmCo99HeONqeG3xFMmukukTb2NKCH
83efpkB7VzbR8pYwE2twvwzNe06XQ7F4w02rtvYWftI7ElE7i8oUD4F9x9IDl4mv
D0B13W9HtT838phLQfHSIEH2pg957Xvz/Cx0wqTPBFjgM+WqFXwQCUJagO5ECUI1
MUO8zc8pYgmBCk57gjuSfhV9Tqp5ipVmVK4fJSM1b8ZMKIlN2xJuIHLjnwINSCMP
Eu75zV8XZGQZKHiCVeG1CncDC8ryPb0tryHuXSp/0Az2g2Dq3i9gRxxHE7AVSpNB
Fc0Ynnt7Xardi5uvd9yEloOxhuFdV/kkXemSB2BkmoBA2FSMp0YEMCIyBaScis7s
5ip2JAVPA11CRuzZO/UeOzF5C61joiKm3VnRUH4viJkUaYzJEYqM1WXg0XFFbSHU
fM+D/pwiaVawlnBsBXEle6vPfqcQbbk0BwUNNYeJMQ8wNOfMthJE4TkvLYRR6Dxo
p+k+Oh1+W9pAAKQdsjlkKyMQbBXC2jW+08udB8OejUgFZS+Job7F6JMMJRZ0T8GI
RywAULOcgJKwvZ/ckIkFqF+iz4Zd7QwfRyvx0b3kt+kYnP+RL9GXlu3ijmMdkZXr
/SMFQU5g5JHFlJ4fV5Uw38U6CPS3+FOe2g2t0doYo2HvBCt+YFRWAe9sxWpBR3vI
ZrcWo9aFMaDykl7gpw+k1JEeeT9JJH0XCR/J2fKrK8aNdg98oDD1vaHEhiBvfhM+
XfAj6ALzjD9KSKiBvoxvZ9woO74LXzaQR52vQ/IiwbemNBZJ85fSE9PSYkD5LOwo
7aHKpoE0Ve1QtL7DAshS6bleJl/vC1ooyZ4AKSAduG1s8SzlNRDbKAmVgmU0l0Bm
NjqYY0bS83VeAAshA3pSRURDj0epWkVXkv3miP3SEFs7EGqmkfkAPHrNBFQmJC6G
+zXhmU3iPhatfsm/K4TdU8wwJgLRwtZgjrETdMiyNRIW73A4DYGZ7qfgvNm33Yqv
hOxEupM9Egw//b1ky+PWie8jJHKdHWQn3vAClu26K3msl1k0/Io+O8SBhHbHqWUD
Hl7J8upOquTzc8F1nQ/YxO1fnL/SGEg710nYN/K1PQhwlwE9VhQGOy4H7SIKL9R9
JqBYZovbgurwyEQWda0g5ZcBUxxfENpHXYfwG9BfJpl0YHDW5M/4BAig4/2VyCTl
cy/E325OCQF14kFBn4x/xO1W8bousXKTQus2QK2+olfSvdVb+6xaZZphgmkwLSFW
xPut8vGw78WY8h2ImSjUwdmDflklWtocQ1I583cUO8GiFoyYIZwtmUzFxf/3EPST
N9ORmgAlOPHVqzYQeHiqLKBf+bhoxh+nqqKH+5aCJv3r1VW4szTfRYMY6C09esvf
wNZ759UXG1ODmGseggV9bw49CI9DVx313Kc3cS3C4CUgbO4H/kUwR7Q/hG2KV/QO
ttecbFXpBg2O/v79IPIuP8AdJNGSTE85WqHDiGndYmDoWXddc7sx9TJPxOmvqkpX
pXWkttGdpSUFw8MZ3vmHthdoGXhbZ4GMZAPB6ugMsznizNhWWyMpaqeoyGJU4Lgl
ZaeBohm3a76hxC35yD/94JjitaVMcqf3qmJxg2lVCUSF1UAbuJs9kc7JtuFsOSDj
Rn46xY8eBdtGorxZBiXMpbMBourq1LNdFnsNjq+Yc4OzSTCkRoDwgX+a99Z8vrdA
3kswZ6MhLGQC8DlBVwol38lnJGY/RUxApxn3phE1jClL6bozLZ/cQRIGZt3lYFJy
wq5hCeERu+ld3AlNcUPJzUb7KKJnMBw+RPIHaRRNU980R8u9E0JpbhqxPlEk9bX8
w6iD1AaejIfLh0spieqQ2G2b8wn8jyo1brZXmzjXKhLXtwzGDUzkJHXfZjfTS41i
knEsc7PgIhKUHjr+rYjy/ZXSKnefb9PDiiRCbOXUeApnK2gWElHcDy9Wm1n2ev1R
7SjxyUjkiTpPB8/2/+XHwsVc2StdHH9nkPw/DMzeYrUenDTFZ8YAQrNvuydwH00A
hGHCDXdph/MnKQ5tE6OqDlsj5DFQJe2dBVJJ3eoMlwceBLxx1iPOUnwFZPQI3Qwl
4yJHWm+B4QoKkZmTwdqaG44s9rL+5S7H+Fq9k3va9wuw4Kzz7wwF1myA2IVmPx3+
/uwx3HFINZBIMaKFPiaFNkNyvy4+QRAoY3aizyD2aSQtxPmrDCpxJ1rxj3BTCFBw
qftnZ4f8sWxrJugw/abYJCMR7N6CsOXgtYc33emqIOQESq4OnwHFu186fh5NTxuQ
JYitUJKAibwdGx3fSGWnyBfQK5LQNfOvuRMG83220F8KkjSQK22xVLOFr6OQ4ezQ
yCQzOYdBsxiHHq1tHWu/swjZBddUzD2bLEtmPQChNrBXoM1zRbP5fFu3ysby42j0
s1or6UVjwwJpdNL7Yu3wlasajUlz43PWxsK24dIXF59V2z5hIIuCkOUjV8vypUpM
128plGMGQRNLaqhzqe3ZOXN77pwTo5whPKvnb5lYj939iiL4Y1vVvck2ysgRCCBh
1svKqLHRro7MWPIWqnKlRmsdjtslmDv3avKMzMKSv4WjJFq0NwDfs6pBrLecp0yC
j6oU40UAD7W1rVdDQ+TXtcNxf6bzWBozI0R3SpVVfdE+7cZyHqPawidA+VEIhE7r
6CiX/DkKN1LPaSntoTKuadH3kveMbSx2G+aGRyNUxAhXmik2LxgkzvJRdnkXMxpx
ZBEF2SCLz+C+ql5bwKpzAzoB9iTebMv4W8BNJEGH3DZN7gSN/Yl6i0DEjZA+pLzK
xYNACw9te0ofAh/fkpPp2oAIFmldhIswycuxvmGO3FnZc8tSL1011361ZyYxIJsB
zPdPdZVIlJyTf1DgfymLhyIqy1VPYytB6fl25EGaSqZv3Yq0+NqZRU1dju7677zS
VUW7XDsyEkQSfizpsHa4Nw4L9blcfSGWKtGlHKCcMKZnZ+nZ/0r9L9/v+8Gntp8D
cVI7XtllFe2GgD8gfLXZ8f8D57Cn2T3iQmr0akOXXNvMR4OHqcqQ9muBuOy85G2X
utaCVrvUgdnq1ddBAuio/IsM+uInEJJ2Ln31Z6InWnbXXZpXJCX+mkzpkE9SxdUX
kvIrLyCGr6jBiYZIvk5qg6XtHdvP0D5W4GZSnCcR+WSKhytRm0w+bsCRARhXoV+c
y71iRcuWIFDkaQcNwvPdWBsqwD9/JdZYbrzK6toylMpm3iXIphizcUa0Hlic4Upx
gAweeoijA7uR6Hatl84vg6wn6MMmtwSTFGbH0hbZGm9vclUxql8yOoScIcIK7aZA
l0wNaMew5JTaGN1gnaZTmKV7NKMKDtrP41DoX7nCtw/1Cb7hUZpk8fIeOJ5js7mt
ScmlG1mB7fMMgwAKeVAoGqJna2oNAtTb3nQzAVNRPwFczA3xFzs2ftwtKjIaW3vl
zfA0ubfPARIVK3gBxS+qCIyAjRzZxd0cj/nb0n4kYqFQ/KBECW48k4AgoD2FB7et
4nydSWoXtw2ZliZJ16QZ4yrntWwLECx4ZC6HAk5EBtXuqXzGAMcuVf/Z9BaqlnSq
6u0+oHSXFjENnqhPKNuE4YHolGWrqMsysGUDih08i8NgBW023wh5XQYr5UFr+/9I
QE0z6ALaECzSDJt1oxT9Bs1NPN78COl2dgCDqCfVIdEqsYFSijaXSX06UU2eN3V5
FnyigLk0w7IRbRIZG7lvZds17bH4dUr05sphtrhGXPojForPZMPKsTZDJiw76YON
NJ3bZL+GwHl017EN6B5+diGN4z3R0b8ZWMLCQuGdXxgTzmhCmt7HqBCtE/7Cah8H
gyCvQ78uzfpzak77KwmX8PD04q6fTLoUsS+t042sAlDeKM6os8HQwhSs/A0SxKIk
+Yji1TW88mogjY4PLchZpiP/17g5qlsKDyVm6J8hMscn5TsgO1fT06lKTrEXWDyz
3WxD5LyoBbyn0aCP7R0pULN4NEU+F5oMnNczxV2VCInF9hhs+9CMAIFrGQhiMgk6
3w3282suEQS30lVLFbu0TYemkkNT2PMO0D2GxAifujF6MxldV+K7q54Sl6uflcfY
LxL6MwOQ/aD3JXy6M3l/yDDqUp9E45T5dtqJ9WO2pPV7MjjX4LOk5WpZfDNb7iCS
34hZ956jA0UGHUO7MNkr+vAXk97f6JxV7yhSx0lfIWUQZdIcOF9uB9VdPXxHEnZO
b8+ruGxFg84r+2YbmcKWbQyc3u+u7gtFRapQXZ93SHqQc2fbfLlQAWEeaJRyCrwa
G5L8AtD9G3+gqjUhdzuzbZv7y9DLkgD1lmoEKpNKPIH/D3Y+pOulONLfdxqJRvAz
RiQIq2DYnbj7jwjKNSOlIWuijSe2UJnGxgOxkJwCnzmLuLmmLnRzBhBrnVVEAqJl
opGZlWboMUfVXhQeSuEIspKYAO0VOX5/fb1gPb6YwZ4x5+8k/S3IpAs7hxKO2jcL
lGqCIhwf0momDKz5+NPh8rwk4jJxFV4vON2xjft1yOl3Pfw+Uczq3paDF3E1ksUE
ENfKvhGo7MNEYYWGqDBvGRV1dxA/Ib1J2ru68ZzGfW6TM83kAnptgjyHaRZCFb6o
b795WEaAyPAX6yevv15/yvxaP1UVVhWJQQ8dS9/pb0H7TqOzPpuGc7yMD52/zyNH
Lh2hJ+7J27vX7Ebg4n0ykDdVXfH9mA0NBGhG+SlErbzP91ZN9UJLOQQrl2A+dWXh
dd/I17mvz9x5IgPhELpkFesYhvR1JUpZZrm+e2fChWg3nfqULjVrPmGg4Pr82oYg
VBpCbQkDVJK/z/xkSHmvICr//gwfro4iqDSN9ClQx3upBx0GFL1Q7tk6B06xP+Av
wMk7zMxp4CyKF46yvih9vwh2aLeRrS3+GAX46Qfkhh7ZK/254Je9CQFfZKzlw5ay
Ib8fTdRK7aXxjDxGdIHYIDPG9A9yRUOW0vJ+rIcc9D4LUFlDg/YNB4QmuGAoTLw6
jkOLEC6ia4ko1JY2bnqd14VPlE6ok00zFMwTTVwsRywl6umNzgjphsGyQkSxCNV+
Iw/k8BUsxrdKWnCCrsAI7NwbpUicNFTZvcDVDGW0chf2dn1nG8PGsaPFBvISHXJU
SkoDAvg2mcQQFP3j+TV7VtzhSVPSSRqF5y8Oe61l4pdx7aJ/uZTB3KnUejvU5E2j
KzmcCy5crTxDiJqKrbYjkku/AXwYpTusXtgd8oa6AZdjhGqPrpQ8dujoMp5qgLD7
zgBGn7XtQKuNn7uQ1SbwW6rlHYGbt+a9QEE+sHKFk34cqLSV99IX4fpgdZoTg//e
EcdIEbdJGEeeg8EXXQ1HEFM8CveA+LKeDx6RVNvKyV+EcF6lVRDJd9Epy+MKoNLa
YObaNvLoaAmRZbqO8+la8hsJqnm+/bfmB7HoI7stmrp0j4IXkM1nYjuY1TrSU2bw
dPb+M5F0GpzyohjwLpGsP/dzot6gwWMvJcF0CiSUGAABvRhBj4A5naxby5xZuO6u
A3KdkLTS54Is7q//aG0qZq/CA+9MxLvRdpUriRkYfaTCGr0ZhddCcDwHhPQbsA9a
0PEwhG95HitXmf6D7EhJ/e1fsIcK6n47esh+SCfKUQDJSAS9q1P4tPq/v8YwcrRE
i0m/97oFY9xP3rZLE9/RdbvXZ2nTYHszsFyp8cIqgIB5w265MlOJ1qtp40mZuoXr
6BthRByA85jq5u0R6jmkZrucwvTHM14Z97yw5wi2nvzyWWqbrXuTAXqMKGRuB5KU
hz2g0HcZ26MofFnTxL4TztqpVmHMpAIWDyRfPL6efB9RdK/lZ8mI3Qr8fXU/l/q6
WCqOmNfRYkrkDAKoP60mLns+rjbSo258UwydKnxrMkkOUFqkdCGDly4vmRYfWKbG
xOK0fqqvmuuIz/ljgKJ2x7CT9V0FHM8FNB9oa628BVNiEAfLuMwujoaeuqKlYb+D
8qUk0xDJftlO9uYfjGJmr0Vq7M5U1lEc6odns8hx7vsF+ntwCaP15DFWai1GDbeV
/1BektjOkkRByIxkqwZGHbQNzmg9S6b4E7/lL+uf9Z1qG0dL36B8mzpg9+n1XOmd
ohS7tC4vMzpsV1dloGDtfJs92rd8ijV3O17wR1vUnF5wL98vxTzTvWPbeb7bEMkn
ONkyT/tAntyauQ9RXQX1RgLAi7Ca7FZk9HkalJCpAjBHEHz/VtRq69KAUAN1HQPp
GO+1gb/1VBPXMPPBgV4ZQh1+b8ZKrC95wfNhLf7CtGOAxxiOWoXbjQp/0Yff00jB
DvJZMidFGyKEVUJKWHHZ9VEQ8bt7/fZopj3KcjFZqdPg1caQjv+YQ/e6nNJK98VU
a8UreqU17lppUHDlXF6WKvRNHVV3E36GABDmax1xDdL/6jkfECXlNIFS+T5yGcIT
vocUvtNBO1/ZMxycs6/KOlOZ4wyiKVMM0TFtey+urihbcPl5UERMpQZ3ZMroT72l
0WCzK+jThdgHYqltZYTDZ2JFeQWDR8DdKtCrsj7LJ7eAqLykDJlT5sFsWCtsGek1
W8WNMOncYJn3WMrN5nTAtUG1D6oEVF3Xg9stw91j0TXSCU4Yvd7hvl0qKWmDwT2h
kFqqarPQ4ezpu3oNRvah81zdLF9cjuDNR6w0R8YavN4CUHFh/tfUibYKvvomQtXG
MXwWp7mW4H8PDlhkFUoJphalElRoGw27ebXDrnNwTInr8fnepaPkIDGxuz/3uBIE
zEtAzhxp0hCCNwAifOmBuhEst6h1auMzFiUnUPquD7hEvpobmtcC6jEjhvQgPtTZ
tazBJn56Rp9HHNAusc0zOoXqT3WmvYlu2j/ISEVL3XlN/KbE0SB8Ytkwh1z9HAc4
RnFZ3y4vjyu8iai+tUWX/FEytfKvcGa7CkhW1IyyyG75CA2LeAsPLAOjCJY0TyDt
5B2kIT7VQNciDlQIPAKVjfjvLWqvAwFlCXQKT4YglxnnFZ2/qkuwdegG+6RIeY2+
GWJsKRAVRfvZnT+waK1XHDwrv+ZcmIf95FfsFCdQyX/nsfLR8Gs1UR4Eg1G7Ikhq
gHBZV+ziASO21RoMlruP2VPvJ2vya0c9Aw+AC1livhQhWTNF6TmMhRcoQhO2QvRN
9bo97OBqLhn5GtrZW8eRDk7MlqrYXwCjWTfxUr1CqS3qwf5faKs4Ac37wSx2W3Vi
IuSwCqu1d44T0pJQzQY/yVvA23pa0Rg8XxFwqfltpwP26tyLu0hqocE8bTozgdbo
BdWFMutSl9i/tMmoohpUXvSVOWBAZc4xQX1o+VjmNWP7C89m6jjKsbTryeJGqZN8
7hv8M2zzpOVbSzbpDuFcieNWaWXtpBQPancE/tIwwOPZi1UyDp0j5Q1I36ubIk6Z
xe56yOgjKBjf507swcAIYJkll/TMx/MhukcpUOTtBSCzlzkI6suQNRvp7f533EHe
oEj/dR17LGVzf0RIy2Stv1T89aoKDXCC5a0dPcS7lsR+jiL3AxY/P0glZ+jSno8N
BrxqRfqR4dsez+IGyae5SaptIJuW1mV/XiCh4AOlq4DH0PBV2/rXpmjChqphrAlj
F9YyPeqb8itUZ+oVMeyidG7ipqhW4kwyRiZXKjlw55FAygTLsVZj61xKMVOIsaPk
1y1vKR//6ChmKZH1EahDcrooycdN5e6sUeTo90a4EU8E8wMKT7O4MdUUN9EaavGN
KEh+X/aONCZdHblaBdqLJ5c6httnQ48eEI+L5l/5Kii7RqzuSafbmwFvoOPGp9x2
Hwa9eUX70wDeQiG+ZBncp4CxRAgSE5JMr5or1UC/+h4eRwwLtsGUOzHw4JcBdUyW
eMlGhQvfEkwoNn/TF7Intl36wS9USLdmCikSkhdiK8Z9sprQDZm4XkHMhrm905u0
dPIyYEvNAAkvnklyZmIP62emcePmiQdnSN1Ymz3+z+GOwaWViGeSqGO0iDM187bS
ARv2ZbaZxppFRH2ofV3ryTsaLyWUHX2Q73RKphpIVE8O+vMsJpF5zC+PhJW+3oz1
9LhE4W8Tcb1n6jfpyokFnyjgXUQd1dgT1LgqMrU/n+3OpbE0Z5FCWcBLxIufVwPD
vY3ZJTv8WjIIawxUl/kVFSfBUbBzdncNMTLWmGG3YqdxcdZFweiw7pH7uJ4BZzPA
yaKkIOLEiSvRXQQVIqfJHdkaMEGp9Ld/2ffrD5VRgfSwYUAdnpBm+KsPF9PTb/LA
3ySVtf1Vk7mL0TEn0v+DgI3VC1+RaXrMF8+GbN3HJwV5Z1JSm1cfURMuXu+LThpf
1ErXishZLKNBVoyASKe69SmPn167zHLj/D5m79542AJt9cfwGoFKFZTFfX3YL1LQ
+i1gR7JWBnyOkTqFV7U+O9ik6BAKqPZoKz0MOc0487Mjz376BZczUlLBYu4L9YGz
IjyV5PqGP6Gyfv+dPB0gxq2q5k6buJpBdRqXm6806Jjcl77dhZECKt21i5tejwNr
Uv+hCdgddVxOqnbtzRgtiGoQJyI7nzUui54Pqq0WV/z/JPilnNtSxO5Ep48nxGgo
tPLzzTdmorxtk+ExRkNbbZE6CX5yqLZD/xt/lAV7MZ6gHOFT8ec91g/AD75fS8rA
sviuR3QJsMtQv1KwDWS8zEFyr+hP/HOnOvj4DzxiUDsAXYsEsOaf5iWUoBMOJuiO
7D4R4ebZFUoLDTlOYEitOCRr72t9q4eY/hKFQ82ShJOmm3HuOjVbmUwK97fanQnF
pRR/SP6Khty8DOJcrDX8njYsY0MKlTo+bcS5XlV4r5gdNwKmdoEfPRT3ghDCPGWn
DJjtPRkvM00Wqy2W7TKTuGeHUkm1tsUhN2ZWxowA7nocDKJz5vY4Ga0lOu1z7p1m
7fLr2T1qIYfwZVMj4DCFSu0TPSm9brc4ap4pScuJ1vkHECiR+K2a9Mjf5LuJl277
oDULQnGxJopkFFtRu3XwiJmwqLfG4CFT4IXjlLLKk7pxx5oWNQmhN8lOmttT4611
XBPTtK4mp/RavfBvEFDfGzuY+utYJ/1MRf4a1cUhFZG73CX1XSNHxlyfQlHvM4FP
fB1uhfRf9ccPjnPCv+FFsFelii+stafqf4KOck1Ap2pKYOV6/+99lfZxtM148GCR
3BlVN7S3JQ+WFaKMTP2meuCo9f85agrlzShdQ6yugClAaQbFEhcow/nI8CEYWGJv
5QrgzsHByNYQlRgTR7YOeTj1ePrjbg46QyYfvf033wFmRC82IgEwEE2QGKNh0cR4
6x2EKAV9DaAdiGiYu4XolE8m3aB5huTl8/Yic02/3iEmLogTJC3cC/yRoU6vxEnH
pV242cF9HZ+ileqq+O+zsPPmQbKc1dse3N7OPUHYWf1+QyDNfmiwKOFauC33yJj+
zHIRvWUIy3Csncqcse684z6s4BeVshqyNxNqCZArLxlJnj2GvSDDszwlDD5APhPJ
a89wU0Q4jvO06uwmKPUWb7yVp0mRCygTG8xvdgrRPqowWnUOoufd+D7xixhngbHS
iJvj1lLoV89dzxMQYSU9zwq3A8WFDGH+T670Z5LhuERyip/guFu+Cw5QsdxRmiwh
Smb+PI+abBAaAAUoZmy4X+12iZa4lgRmjJXLX2cnrGk6fYNiEU6e4LkrX2LIvBRm
jom0itCh0VCnRHCxCS9PhPUIix/NoCobu7xEZLhnldjFSF5DADxXGu1emoGTW6wR
R9d+PTqsyYVGIywgHsne/ZjvIba/Y60FFjnikAAwg7+Lu3qWqOUxwN/XyU/+evtK
USILPwH0Hs9IX4ReXti1JZYYk824rxRAhlu6hOoFI4X7iU0xhFRLU9Lx5SSbo/9l
n0fS9TymHoE2lnm2SIwFy1rix1sU49Gi3QRT2TrHJfVGMc+wy1UbOjIk+mk7XMxC
1JUvKPCf7zK3pGzlwKCTEjd1jEd5BBhekcgq1vDXVzb9lf117w6KBWWcTDSkKiHu
Ww3g7+8CH85Eh5wyzR00eVidt8Kt+Ju4I79lUFxMHBmC62ecrFSQlduXqri7DT6Z
A4o2a/PQekioTEQYKX0kJ8f4BjZ3vYnnboor03VN0LDuBbx3qE7NgVZxKcfH//np
MBhUdm8g3lAY+W5mxn6XbDlOxbyhUe/3bpkt+kwgVcP4mj51Csqw27RO2aL9X5Dv
lIm7NsCOu9hCJp4PzA+zbqkXZHdXKQoOx0kpE88tpvq3XbHyQXaZzEb/BElZCdjt
thN/BJN2PzDnqbreiuzq9H4YB9VMydjMUICuMrfUKsep2SJEwnN7W7uiXaLNInc3
G6yTIUuwbSbh50q5vr/CdCh6tBYjmcjBs3WCccZfOOkpzPv85Gvq9DjBuWTtq11/
KVkgwCcNZZLn15oPzc2yEIe8ocpH/13qsIuXLheyEmSclYav0qQLMEfLlTFd5Zq1
/V0w1hEhHRuxUOcQskhtM4mmZl1RaPP5ZIkb20FvONUF93G6VLwDQu+F/Me7YAoW
gx65MMgwnRqEDr2LiDNAulK/UEHTuBteukweuDA7KkaKWoC8qpxPCEkmQcij3YHl
CJK3ZAqjHvhaU9CJFb2px+psY99qhx2w7WhtN9NlVPDNe9GVVn/qbZvZ62BzHlD/
mSmuYTzHRM/FbUJyfF0+Mb9hAHr/OLOQaQxYbzoOgbDVgeMW9eMr4gUWOrFzru6E
oCFS2pj5wxo1z5Nez/jfyiAZt+VoFdM9MgTjADdKYAlIDPVFoTzuYUuNkHWwiFds
5JB3X1sW0CUZMGnFi0U8U9fZZp7ZFwgciEblv7Zg16MCtIyco8wrgP4suxhoZptT
472AXqTFoH66CydyQW38+gMMpCQ3MIuBW0O63QoTWD3GQpOuBmfIaAwFTPUcLAmD
EVpfVIK9HWfUjW+y4V5MV1Rl9k7FdWP0jKMkWk627BqrxlF4CQHd+VPvrmg/BmZ4
RhEAFHdKEE4anNoKxzaVq4wBAjGkbXkFRysbdkjWrfl6FI1Mln57aAGjBG9HEhKw
ch4qq3KKH0bvcYMVfXDMfBLb9bY/Oa+1gInzk3UZ0p0/gWXRPPddX055hsZg16Tt
SzS6HfUPuak8OOyJ9u14vfZeCEbO1eJ6pLAnNQqq3rL/qwrroQmIlf078lg6IyGw
95XDVFL69kbtiLgEcTUaX25+G1QbnMlOS1KNedTvlx7bbXKOxSxaFiT29F/njGcV
otu6T++gGjSCAaDLDBv/tHsMwCCtk7BDV5ijcNpkIYqWTh/OO6z9khu0E7DtpNW4
JcnRYK+lpvasgAioDlAV2f+IwEqk+zUyC2fkNO3KNQgtTjhFCRYeGTKGouqmZd6Q
0rRFW6jCJpU9pYeg/XWU+kT2h3hWWXZwu8QkTmqUWZeT9HluPea0JFlIBRPBcyK4
3xZeHqhizPGv21pqQoJbC63xV7xyDEUSf9KGjddUByDC2q9XAv0KHUErA4uUH+Gv
/ukmx+sQLyNJNQAaC//weYdwJLYWcQRppYX2CxLxpurTmbRQnW0tb9o7rLohHrHl
EPYMDVGURXUIZQ7Igcasrs6+E9USrBVb0rIW/cnqkt/ds/yAqJdo2XMefWrpX37j
zoD+p8UTZPTry36V8xs1qrbZCUpOmaXuENgaGDSq3CtYy7TeWidsG3Rf/+/L5rYV
R4JKt0erJOynU1fKd2Us3PmRQYNuXN6aU7y8uRNITvfYFTddHYSvWFiKX/epfIfG
O9p3B2mdVlDL3jYpecsrCyzQomEEI+ztvUjI4RItunELjcWbr5mDBVYAPl+XVjXQ
ylw5j4l97h3dXAVdsqiLEeKUjW3bO3C1fm+Ep0E2BW8weZxToAvGrem3a682LOL1
DT+6rnIn7R7deLcuNDTwdPWxeLr5n5G3GSMvzDWHw0QMTOwtz41+Wfwyh1UFtES+
Zb7U79Lv8jenvZdWt4fZGk1xMZH1uqZDwMG/Z2M3Yp4JkDLYFjlkyizdPW4NmHXL
1Tmo2TYJyGw/ZvtfeclqisxOrUsXlvs7wWBO+/ibvgQsyNiPDS6t80g66P3x55lK
4Iu7W1piKSw2MxfO7dIswIewZjJP6nIIxQPj3CGTnhdlvSg78RFTIlbVBh0nOt+/
hX0/UjJr63Lu2t7M6GKbERf5jzi+LV8Seg88k55bfB2SQo8OzzTZ44f8+BniCLVt
M+qwYWNjLtSWinX1zIJnVoQW1Th+0x7J4iCRZV7QvnZT1wMKykH/Q10umqmpUsjs
9Vc5zhOx8AjS5cY6ULacozd+lLD6iuD5K/lz5JSpoRwrkiqEyRO1X5DygEuacAUU
9iMCZeyTgMKOAvPQ9woe2UI/Y9x2JdtiQbO6oabuxvtFXTOJ7sO5NnwIQwT0obwn
N2Yil4QblY3+llIcVOfVGDN3oSlZnHybsNjCjqOOBMi7Iy+g1MFOdw0CAuMMl5o8
rGKnROBXFaEboD+H8J+BmKiDAYJ2UMQNcHZ7piIS0516eOOxijBaUCop8e5su0dy
KhSwGoU0rSvRxN/Xzzi1DgU7fNE7s/pB8nLe0uAqfCFZUSigHZwFBn7G0g35hFoS
tR0b5h+dGIPq5+9i++VODzDeD6e8/en8vMmZTdgzwU52fnRtmhgnjnG3o5P/j6nl
n7WhidIqUL8R+tXPaIFj0jblLkSCReNNmHrMvx7aTldfxP5QoISR2szXF3U5ENB6
SqLwF8sqU+ILWUtEl2P7ajnsntr18psiJAKNRj7DQ/Ugc+UEbeOuE3mrTCRMMY28
kO87lGSSHKOACR55ybav0LIr47s4RNxbSDteM8cCIn3v+MPX9kbH17Nlyx69zFl8
f+b9nDqp8lTEs2V/L4e2ZknTdo1JeyTG/KLzPygRnrzhmEmPBDTdypZDlnDkB/Cl
2VkjwD4u6FXXgk3LCI2Wf0GksSxVIFo5FSoMCs0kuyeZvetrW037XMzXbOtVBQ1r
fFAcNAUR9JcdVKW6IHs7dp5/vgyQ5BZD6D9rCygf9vdiStOnK+bttOJHqjq+5jG0
zquA1Kh0p1jzC6wcCuuhHChZOUDZTbKMLiNz70pKE8uth/b5at14bcVBBsOC2mP5
Y3pFYAF/qD4f5OtXcrhCBg1qRNeaKyzWzjrMqo/mbPI5959S+Y1lAXW3kv/XkA0s
x77jyccr3oXVeZBbSMSMGN4dyrcFHWtR05eDBYE682dId7EL+gC98BgGTasDsQfL
5BUhLk8/YGK2vGPsusYfnjH06dGv4ylGR7eBKFipaymLe2deOhg/w6Tx6q6SpRfB
60R1H8dfGymr3jIQSjpB6kSMRylCssBpR1c5Tuc9D+y0iFLYOe5WzTh3ojk7gq0h
AVrjlEvuNhQkEDrCQD4jZTLyYEp49r48Xgb+c5liAp0VoS7Cy84uw/Gt5ohH/Kih
g1lJrKTlSBZpG2+VfhX42U82VxT6L/3NGFOlm//Kptaz4ShOrSSL2n/2vuVaKowm
E5gBBQl/9AyYVJDzQEIPJbzCPx2JwEuY5MMpnbvuyrzPPi1RNxJ9KZVr00oGn6o3
Q2pAO/nF2bxIPg1djCaCfR1Rr28OPI81vwBnRei13Z4L1Xf/vzg2YQOZnxj8SJGp
hUtbFsCh1pwJvvT7OqG5HXcCDmXGOZc4B/NNqB3ZVTWpNGvABqwO3RxfpcV/Ixm5
3KTgCL5/ehN287ogkveifE8TzpXwlX5+S8AJaSW5/S3PJjRmNE1CZfAuDkhAPHDE
7Y2q+oEtVhJariSR5VqUQXNrX/lX5tr8EggZH95Sk79MuvAoU+q6MzDHhj6PSZmj
t1ZgX63ZgCKuxKuyBerYpMkvAeGQPSvb/Bp1pDLG96TmABWRJtuPcGz6kvgH1t8f
34frrHkY+GlgVLTCOXGKWmaLoeGufRjaXJlzYb3+ROGN4q2fkcGuNuTefnDCg8GW
BtqNNp0Ko7A3JkCkSHD1MPKFC2t0O+gOTBO7gwDraBODDzOAROHoTxGptz+sX8XE
r0yEeVTkVqgbaf65hZYgzzOZixHkH0kfuHD6kKMYYiJH8OPfi15Y27w5z+ejbuhr
pApk208x3N3YCjAuEa3s6MpcUkV0xwgvbET8TG3XTIu1nxILelhgGMlySkb/pJ4t
EqnrxMj66oW+6LuMMWtdwRwFzU51MfeiMuGMhT7eCIyqhiERc5KgAbyPD2ywmgA1
ntXHvbF50B+3qVC6pCqbVrF4RincJyMFnzVSzDmh4UCxt5g0K5nDmDfRw3UO0F8/
eCramqH3KxZh3XQNKaIvE538pYvHdInUz3OrdQcR0A9whvp6mPa0fzLAiXuDcqHs
kEJtdW+dArWcz51V5D7NG/Imh1Douf6HAoeiF5lPYeaHUH84wAU/ZYuIdat4S6oW
YijCdZAK7LhNNAcvZKqY6yvOOX4LPKyx4L/UcdXrXgcYiZWykHSGFp+bNgqUbiGh
P+Y1w8neVcjnbnaKoPyzJQ1KT9p/xtOZh0kKlQLGSEZ19udhGg1PMZhRIfVo37Tj
uJWX5uzuFq9hxqnWLTNXW+KRglU6U2nGXkhY2R8Z6TuR5ZJzsRy/uFuJIkSlaMnn
uDqAwskBCqfSmrl4bnUYAFxNgLW/b9cl7k3OPa1zRBLckpSXLQdoft+pft7t2JZ3
A9L6S+TL3wziiNtnV1+dgHOvdCDe1Qa4T/H8GSqLIUdoZ7FvKwpZjhBx1tiTR3J5
JTBcuiHnwd35val0VEmmShhvLzpoedp6kBeszhu8D/AD/QKAm84PFnu8WFlRYDdx
piQXv0N3rCtF/ZD4z9agyqeeRRHOj8eeOr33Cb+fe7JIrbZdNibbOs/CHOt8dNP2
4HTIR+aGi+ne3gjge0kTihGnSpJwq7g1ft202Ex85dljtbf25JrQAsf4lDlVSV5v
pMws5X629IKBc3aT26DTdOiOzKmU2njsLeeYkkcdunUdIbUdEw0TrMHxibJK44Mc
Cfk63Zdank8QcXEKs+f8gt1GlA2MxPTVTpXo/Iu2mJudUiDxyLCwp85DxZTvbLd4
pQYvqBqqbb3He4t8HumRZoU/3G61ECrJmTDA8YqZNlpDOdK6dEX9WtkdWsWIgVIS
kV3/+AZ7C0/B7oLZ6ZctnEJLNxRec4Mc4iqTnCp24NNJvXDGhYd2nOlZf9vIdAUW
ulck+wDn8xJADlJNL51rQi+ZCye+ov7LIF0s10N/lJUgCPR63ZHrjN/cjkLH7QaC
HuIZzbJMC8NpZe1SSPuOWskZ9wW7staK5dKBRHGvarKaWUNo6f4dreS+GYToStFw
osvglkULysjIBJqo4FirjV1/7JLdF2IxkJeMpsRTkCqzZE84uHo0RfL8L0E5Uyva
F1ghp5K0yDM2UmxtlJHcM53O0OakuPq9uqjy+1T/4+d6eF4wak+RGftd4ynVvVmR
K53TE+siIvsJv8avQSp4C8hMP5/MIrs3PbXsIEsAk90d0AkXZrIY8zx+SaRF6d84
10JEFnzqYciCEGZOwy4ldQ9KHDcQ+ySxapskxlz6MOvRBv/C5SUsHN/dIs5XPaGx
+nXpyfVKcgUMeq2xDlM947MvWqy0YJQ4nXWjirnWSTf/6ojwlGo3c1Z4nXZlAk5k
Mdx6Vg/2iNk0MEY3u6bXfJEqhoiFJH9Nf8WxJ1C9ozmjyb/T+5j+GZuv+m7VR29W
D67PIntkL8p5verK6A7LBevKsHrMCw9R1zd114LJUVyRik/L8gjrSaw9uBBVjI+A
bztM9v+sTa4fngc/WepVqo3Z2Bd4M0ZEoOTYuBxK9cLFD0BQaod23XedEcdPxUWv
89SGFMrJfnTegyfe+t54YwyTKfdujbpzFOt3vQA8KjNvpC/PGa8tJNbaDyfHCOGS
gEP03+2CWxaXo4gplIocZVOpIjwxvWeu6jFK0dPWtg1qCloAniDcUyposvLMS5u8
265Wd2cD6uZ4esaayYIS7WhjZhd5eU1w0dAYAe+QHgYbtHkO6b0agjQS9986x0Gu
+OkzcP7GZQeaKHpl3c3bc9h6eNCerLfeXHKhmyECb2U+5peFvBQJCCk/ntxZqkRy
RgvniYg+3ypzfAjTxDelN+NCQtltpZpZeAllvOpb686k6zOAiePtdtUF1H48nyT8
rE/+s3T0ymsD43HZxPgQeIXpDf/b44F+MOYEC7J19GivXBfg2sSMb90CgSuFdp3s
5f+SvVRC0bcvzuZa+mj279ry37A5vEk+3wmRH846Z1CpFhzCdEISf81ho5AFnZ/y
tbx1PBtBejsU81z1ZWJHKJtamSP0caHXq/8T3wFT3uUHMT6vgkDRaMY/ZoIajt72
Gi8nDmgsiTeX/Oq6/lmWKJNnHKzFmgvP7Ad+xIninFUZbAFLOZiJrkTpGZ1wvue/
wsmyFUzdsi9slwFu7TF4kJRktff+K9M492MqKZHTiidnie2zLlDOOk3LNLO6VHWb
Sfa+Mhjn3EY/GxxxaM8V85ferH9SJnySy3OL2hlW8f7UjEdBFsIwn7zm7AzLs8IZ
WyNQe6w0PSSeV8NO6rTHgmuHla/eumg6l1/l1zXEXvpazQloYtmM1h/+kM8DwYEq
gV49kw9Oc5JUM37cC+VDHF1rYYkRHwN5Ir9GtVXE3WXfwBpNq5fl3BkC174B5IfD
kf6MAWs3DCpJ43TWv2BNSatKcp3MDUcmOXvLSvlgaMoT5udcz/r4cyV+O/3j2x8+
S2VoazrXjkrxuDdHkRB/yMkDcRyDcsCnAOOZr2k9AK1GrkRiLK0rBgAmeS1JRoCj
On9WGBTyHBjq7IqQrQEFtmbNFOzrslYVvb+V2dVQd03S9cedA6oTZViP5SDwTUa4
r/O59C/CoxuUBjTFkVN7eSBy2qCVFGUq23vcclzr59oybm8saU+lAABrUncu5Acj
qumC4H3yPYO19ChObWVzeBDX5xmy+ncVVrrlCMA/LvKpMCvkj/llOPmWXeIprrXQ
oCHS2l5GWGWHeUV8jRsD2o600BLqetlY8YOVmUBw7/CAw9GnACpoVzDmBilpv3xs
dSB8o0LrZn6TythyVLQL94afUIRPJ5iyqwoE3WipKBjL+r0ik2w5GPtiEKbASAiZ
3rXwB/qvLWBtWBsrsQv2q0K+CHVhSpoKmMZK2e9k/kR51DXQACMx2zWI6kRu9VG5
MtfmkpZxMsmpI0cKEZ+24XOr8eTdD4YuKloszRyKvtJ0BTlsyPCqS+cEgYxfBbLw
H9JohEriLVVEFAhM4WSyT4mscEpHJhVmTCcrRJV/biFxJP1Cs1BnHo2ov7eGLVxH
ID2dML60JNhU3g7YiPYs6GVIRgKiLYnvksxPKE8W3XCb0RilUP5Ajh2+Vzghot/U
rBxPBkm06UD1uePOXhgl7ODwJuJMtW44YqE78nMvjlFcUJUa2zv/ZOSbfbMyYDdb
GE6Zq4agcfflYHuzzU/gEzY2MFAzTDVciR2a8EuwaFg1lOB/QRMPvXqCHvx/Ue8q
v3ItjOApZqyF6P01yHEo3oepJ+l4a4pjrvGM+QQdPI3wsjwwymlcrvfUWjjxaymR
+VFaVexwyqcl6rC4cthQ+FPDz0IVOMKvUCPzLR4lDKZzYrlA0/CiBdb4LSFM8zR8
fBxVt7buEO09sh2nJ1aSNCM9pa/wbsHQH8bHpBRL6OpDTn7s1HIpzDDaSJHcUhCo
iDnBsA3Sk9L2/UOHzm/TpjuZK2SyK6MzFQkx6tuzUhz6cJM8OF4lKbMafbNSlXO7
qdbbv2Vg9uu2owmTL3SExxImwqfzhlgp38PupGCDSCfyMk9bETtXtBIcYtKpAWoS
dWZ7Dxh/dlTzGUk4b+W31zKVnY4ikNYAx9yrbiHU55kuZh2Vyz9qFF98kYM3lWif
Jqh27XSYCxwG2A6lfC1thnRCELrVj7l2PMCcL4zf7r/UksExi5UNQEBcyNxE97tM
xl8FXchrn8Zu6Tko7GGRQ4eOTieUyGfrbEf3nMIQTutC2M4dH2+Bhyk6YDXgLz/7
5Xpiu9ayNFMh6vbKnowXeN4ZwMC+7ivCGW8BlipZB2lFw+JdnczbHVPSyGLqQTIR
eW7OWoRYQzKNLC7CbmMGzB+us/uqiZhKx/bT0ToJsJtP2vRKYnHbBHQvCl1BMjf5
zIhW9BCeEnipl7EFl0/IBI0AgluXSNFFpK/ZnVYaR7RC9Ao6sP8PmbpW96aDewhe
SlYHbvNFfYdb0hfqsYThvP6Ygej7qvOw1yLPPV9MQMYpn+8L72o4Q6GefC5/WZxl
YdY+74pqIrgNtr/Rz1HsqeiRHwT6mlS5Xz+jE3wv8OBEJJCZ+p8fctFIZ6gEdyLN
ehf9u7Mf9cjaRcCiYCVbWJgHc7kc7jF6a97UM30dXtR1AhobokIV0yM07vURhz8U
Vc3IFF9CeG0f7REIfyCyHYt5dDgGVut73B6C3Jv5Rn1vspL7ICW5z+MUnBFjLOkc
NXsDnCkum7z5/2ZwnvF4xVgSqpu2JWXbqu++pfEPDHanRSp3IDUFVKo0DJsPAf8r
PogqZkKR8CRFaB6euZExCPqVOKvav0ldUEpIGpRQqVOqHmSAZ/C7g+1eliVDhWcF
refzVasCJH1ypqZngaYvrAAQ8nE/a4XJSTPwiKMX27j8hn5jDXGAYp//ZclKPJnQ
9N7yFp2+AX55AqxfR6DtTgYNHT6xEPEAjjLElb37EvJKsBLJHIz9dfuIuZ4WoA2f
qzBqhKdKc4lYOZuMzaYnUpm6VQdUUEHJHoME1/Iq77OVg3e3+uTUZnDZA2A8Mnvs
VQTPWh2Q10CC/s92TeEodZ2FV7aH22SoxKJTYdDW2KI/8SRkeosHsBeV8PqOceqx
sH6whDrFF7bXbofu0ivxzha+SqZDLyoZ63HVhyVcsVmvvDX7ulom12x7ef/nBngr
i7SgTBuw/VMVzFB8oICXI9bUGOdJATWxHjUYhfoiD/VtBdAAuQUPoNbmuRNRlPOL
vxifF7uYWR3SjOnXbp2Aa8Swm8D50EFM0C44cJLDMzK4YuTZIXp/M9ygjLe4tBrP
dGgW0mPIsK4IpZ6mHf4xugSrkxPwx+ceL1R/fUCsh3mmumFQjqO3VvpJTDnZmpX1
kuFPTkpHPJSyIIRcWARzTe5Dk3ulgsjYeV6ibjCjCt6Nt7/CdX0HzuSIBoyaEhrH
vta3A5yccqsjJqvJqn3/AKBFP8MgBfSw4xt9oZoqv7YpaXjG7JrSflMNQLmRmeel
Sg2RuRIEt/5JTI3MzwqmR5XVhkky6LrtSKeSgtKFoJG9tHVCVGgo/omeC33xzRkp
44Nay7twIIJh5GNtnk9cuHbVBSq8GlYLihis4VBbCCssuW7wZ/LkHOgYlAVgZGEM
/m096Ydivlnr0uID26qhRw/pBpuR8dQROqDlhP6HnhjsRIuNwYtqGl1yI9bUzuPP
9NhZfzREs9ce3f3uNxZ5iXg7EmUIrXUic6826bC/QDt4/hO79dn2rwyIaNBoPVLZ
LYbW2XncARxIxtxV6T9eHM0zxomrm4Dm/dMtaN+pJ4vkD6b8W3DI8QtnZPhIzjP7
lbgUiYL3+bJceP+9tbdQRk65+uVRXCSkQf3gUw9RAqLoWzwVmfOiQXfEPGAJNWbx
CI/+WEpMO+uXK2XPsBcTAK5EMBS3zYXbAjIHTyWeJwHRLL9qf7pQD1U1r39xaCVs
ufiSuDGhh24gO1rsKJUfZcvG/Ly+3MqCgW/3FADmOxnvse7Glp7GoiOIKuLJcNrP
x/8S1kU5ePXm74V57zC6jL4kaTCd1yNer7HODSAJH7a82WKDMzpQ4iFck+FPTZnP
tenR9wW7Pq/Ev4Inx+PNx1CRW+fuNnP7baKiVFuoBNC6edJ/RHrcVrUaDjssmVjn
KXL89jZlkjjiZ5N3eAg24jJM7AdpHJvs44u+OabHN2T39MNv7uYLo0at6ksWPOBs
79LvoVurrTeLiPb3+Kn6RhYaOCDqTgJKxWxFyCQZ1LOiLz/sygO4e3775VcDFRYx
N59j8Z+kfeG1AiLLhDV5Bx4aM/6pQv2RA6Mlk2Q1F7nFdjGBzftN7qurSlAfEUB+
C7eMv3ieU64gjfILR5VdFzg7EHDjOwsFQUwDU5RpbVcd8bD0kIiDom5JgTeU4W/k
n5ahcu/8Dfa80ZAvbhA9+QZ2qs8DhvKSQZZQ5uJEXWU3Y1tsPM8keu+FVvCVrvke
/o2fC+1cEH2du8lE2xU9q9M3NZ0/hGrtiBJktsA1jRC47Z0HgmVIHwneY3rXopfT
mpnF1520KmFOeKzritSYOgViymN39zaidg20t781WcU8iHDXTzF/DxefPe4PC1r8
RbetXucMXPMLITdpySlKwT6xOomV8Veu204ffDDxD6nKltIXAosE2VBxZQBxYhxw
w4z6fQ+1QfE7jU2hujqdwrSEwFWu5vjYNnNIFOCrz/KyLoNQWRfQqrfM/bCUwjHb
qPDJ69N/GHYfndmy8G+9Pc8p0/31Cv2QP0NezrAO4EwHAjxZodRgrL+hxDoWSTPs
YrK3XEA2Lrca2EYQIZlfe3A9xxfNhMznkSvOwVbpv3wHT/dPAbEsiU8DSqtOjfbt
sPSJIRpl7wQxf5F5k6breJD6WwbNyndJ7m3R9Hbj7C/W5kHkvSpkseszOb2b5EfE
7cBpVALfdFODQvKOEaWXtwOG4QFFaidR+PtymeeIuX3mdWJCnjvPefGjYATBl4A6
bxUG9/G1JYsUSycJw/jE+t9FNDVyPAOE53vltIl1GHFRbfzNyTEZzpCu6yvmRLmC
AHXQUw01hA2JwVKNVFixNzceNce6GSPrJIGnATRC7XV0Uvw0eMyhlqje3Nz/nrqZ
H4aD34qb5qvzom7cpxCy2U+5WQFWxtxFmojQZxcaRmvNBK/v8wG4PI6+Wm5f4eXf
Z6xDaLYhVjmhcFxiUxeK/8njjZZwlx0Fd5UmhjNNE+GGgdczxw8eoNFRtbv/+1ih
2K0svoI4diKxrDIQFdipi8kSjcnsb/Znges/apXMYJpJ5vDTJFmC0iO6FEySYVjk
0UubXystGLxhdSNpp8VUVHyUF5zKh1WSNnmADzJdLPQL7bRrrkuc04ugLM0uevLU
OMKqa6DVdSe7EB81XMvfer7WrKxWCFWc5N4FzX5oZqFjxubenZBvvu7QkecZ524J
Sw/oq9YZro7rflIo6heWLbotTL8xFZEJOxFIHH1athN3vjh6mPn8NFZM9KfACpPK
0LP+13XAM5EoiaI7Orv4sJPBwqcuoSW2BxuZxp2aXBkqtP4J6GbHSb36lL5NPiFM
NYVaHC3pK/gmRzdU2UTH5xhFu6m1hOy7J5IhvMVjk3S6Sf6GUt08hoYjnE/qNVkQ
6wFozwSCUBNTLRGfhCC5i/J1v/w8zqkB5M69d4axXcOu4IZHLYCuL+0zpCPjEyab
uwGIEnZhgYZuWBBbQs3U/htaDc637jpJbL9iR2XUyO+L3M3CYP3QPyM0uwlgkBz7
jPa4mT/Asq163c0bxKq+CE1KNZe4uuQq/cr3jHGCsMlbaC0NSvNzP/OuOO3ugTZe
xOvUZ67UGdKwsMsKhCLsB4O2KQ+cSwueUSKy1uYC2Igj/HFMgHFmnoerubaoQcAx
+/kZVRUMrJrUOjo5wA/aVGCjr3nYZiykGmqHbhRJPbPL1csVXnR55f+hUs9vHInj
PmXijWG2LNZ0B19IJ3Hj3cpeeoiWM3GTBIBRBypsf4Uy2UfX7YvO96paT6RosTQi
mRWFhLrB+Uh49rVT6OUBTCVmOscBJiG7mNF+4TgxPdof0C38bw2lSWjR8c42LQBv
7xlAPmNNf5CIWdffrSwB/GCgu4QidYNXIRlCnIa0mqeEkzI06wOoSjRtr9yZ0AH2
BOAdAK4VKDcO3sBP1POvT+PGy+UixlMB91TgQqLKkDVUOTQu4rv0p5IE9Sh2GmoR
rlFGW+kqDtavjlfqRodmA0ui5rwLrENMXZlYj+HgGs6f4Wg077NhD1ZaGZ7n6DA/
LsdRaFVDIqao8oroXR0az4V+OMfvAfenkk7spFQ+1JrVIX4S0lxIpS0noRa5cztx
WvK54ztnHNbIyAbY7prRTe0mQk94tq9ikl9G7bpo6/GpZaMBh+cbZxZ0l8fST9zE
q5LUL9Bay7kk6wBYU5RasAdQCF+GcfbkbMYX9LctXznpuCrUZFSR6dAyeR5YqYVM
XVJCgK1pEEvUdcQOO82peRHF4+PyBtkm0Ug+8Gud2LDQMamoRIuOiu6wh5Lotj++
kGXg6T1ytJpIQMt6ZyeyiluvulC6sLp5k18t8c75jr1LqrE62iVaNajn/ubvCU4t
y0mR1W+YAZG4TgAI3jaeBYF8jR7ENFPDukHvvbS4v4HmT2tF1Y9rjxxtcn90ubEN
VTPKnWVhyyDpTn6Uu071wZhdearB4kR6fEd1UI/n5742yL/kJ3bxFor0/yXaJS/I
WFGa00B/woWSP0Ip0PyGsMU4X9S6+ZZkH3ag++CeLYlq5Tj8EJqtppZSUZnSJjvJ
KOLYFodjAF0RlXbBb0SAu2plMUW3B3bJM11tcOugT8/NJdGR8jqXHPPZJz9GUMEJ
LPcsvhuEfeogHr4w2aXmXySrW/nXGaaEsXvaHBZFEbAbnMRg9PPeXttLtp9ClXdS
urJDlSASS5quIhlx3vdeVVXY6lRREHrGw/5MWPcfd/EaomMK+p0v7uY+Tts2UeCF
tLKMBcoHOmXrP57ES9u5HW05lLnm+pibA8w5zdsAfnxZpBxWQsflLIbGQImqKBtu
vDWz1MJnY5GyqRbScfWQT7dWfwkpKl/dop42WdqYCWg14yQcrgJPeIs0WefaTryN
IpRVOUmgxIwgrL24swqtLek40wVjIFczIM3OOFkWrGHaQqE+ThQd0HmTo8OCOCQH
Gz8YjoPVHzI26ye/a8OeibaHIyRYo7+BUcRttXrjt4WeeuVZIz2xqu8Hx+nHQgl2
HZpN2eadKOtt1+EZYVM0Q0wsP7ApZ1RRdgMOuW5oK1lv77vzt9fv8gSwip6YgMSg
gia+XZ11tQWGtW0N3sd19GNdYE+WLIhqSkT4E45woYxtppA15gt43gTNXOwblXDq
EaX9t+7Dih4jwRu8OyPmDo4q8Nl39aLohgY+/b49dSWLTbSQ8qDEA/MhXDaxc0MW
mV78ajj/1zCQiltT/AsycTRMujZb2nTqpGwco4lZi5aRC0rJs8yUxhkt3tY9GpU1
Uw0DC4LpqvhtGUwydDNyRW/+BlpPnJcBENVGa85nnZeKBKjbzLU2G7r3ae9XVIir
Fbi0qoLqn6lBNAbW0r7RRoDOy75CrNzRmtdXoWpB3pl2M4707PoazTGa8Coguwg9
oE9f4856AdUpyQ8myjokyCczayQ3Nitf6s/88wptFKSdwwwuGCV/uu3kSW/+/qgB
2ZCWIsiJ/Ff69pHBOXxhDhjpNvTMq5EDjYrYOhL0i8Z7hcrHho5hJTO3m3V9+NJr
8jyap6V7SPibhmkkf0WOYBx8EirisAB2RD3ttM9p5L/A1SWIw/fN3IE4NRLmXAoQ
YhrI/NdKj6bxXf7EiTcuGZBWdqm7Jj0rxkG6wDRwd5mWEjzRr4LolgFPhK2oR2kp
jaTgIyqWQf6Y5XXvS4CzYS3jX54W9p6jjwcXKNFDFb+qOL2xfxjSaUg4EQkTgD6Z
Ks+O/0HF7v8y1Pn4d2lHvaHpeDJ2W+1t9EeQF/kbXNahhHwYoL/N+zij25lygNU3
BPuUe5bygoKmWgVyMbNgx9Xmsu0n829vu7iBhaZkEOzw98bYswtpy8fSZo9sCR74
38lNIuMRrQdm6vfGi4px9bGyhVqL6JsgWXzqsOo9ExAq0sqcc5S3JUPuZC39muJl
mp072+8VuUysX+s+78wCGCreenkpaqcK9h/nt3FkcCzPfPkcmzoO5hg2CbLebbVt
YPIr6ha/enIVA8F6UqdYA9tbNVM/ATQ4cz25Hbxz5WSdnIycwJC5IFmF4k91BOCz
jU8lR3KpG1h2a7/pN0Oy1c8LlQDZzA7UvZvcf/aNTBO3wS1cgUGu/fPjQm5/XKsJ
JKEras+HPFsvQ/wYJlPj0rD46UwPPIhiwzwS31EqabCRqkNSdJBXOEJbZYO8IOXE
EsOBNsv3Gb35EyIIpPrjKMzSy22s7SkEkjFYCCBZEIW/Utq+OVwKzsDZ/38Flb5b
0A5rSFlONvUkodWkMvfNDnL2GntQy8GnQMZjlLdpUHerKVPH62QuQ3YJIDRGlJN2
C1kvWCd1lVOfxVF8EpUmsqkznQcYtmOcn99+IJwSeRoPVbYN4COlDC/sgu9ru1DA
Ghiq4/lL2itl37gFL221jsfHVX/CE+a8RnP95qB8x411jzSL5CFdaiy73B45Gbvu
Z5X70KOiJv6JgYTIK3wbmKv0M50nLqNo5q/3cEa5T7RzyS7rOeeGVVcteJV1tYHl
G3oMnhFxpo4yYuSuAbO+hftx1Y8qyzACOuVtOgCpSdiKAuHXHl1ARTsQbG4pjb3S
dRW4UeQ3dH2xYiC1uMRgZea9+3fNy5emuIDeA8Xf9CURnBxklkjGjd8Xer70/24L
U4vTpEB0LJUMbEjBX2Ktch7of8N4jpAk1yB7ND8ACdUurg7+ksbL0e/9Wqvz6xFt
iGgaYRSpFAReHPpOxV7uUf2rmQU1nR+b3dMEoITK5UF3CR4QqlvccqmqDLcI3qS7
zhbhdHq6Zx0FXCH7Xh6i2KoNha9alPkUur7QHH/LkM4TH4zT56YlMR6di1PT9dey
yRxlzhPVKANBfZ/rNjhfHTHePpppkVDP/BOQMZXdiKhLy1dN6OK2Upp+3ojXaJgk
YkkcE3Aeb+3nZAxVtjS5HyJ7ApzKmtUnA1I3S6dBdSfYh2/XZL3IiO6XEv6y9lgK
8Lwvx1A2HiHzyRgJ2DvZZljLRx2gXLiF/PxAwIp+ZFilBhb2IXPj2ERPJGexZs4U
GMMXQW4IP4MdhEc3vr6425ffH5cEiy+5UFEVyvOE2w0JyyTT7U9bx53XgdUBeiz3
HqrU6chdDjPIeCE1NloJfvDsDj5sQpf6b+DpG92Z9D9wGBxbV9K4UjsylDM/Frxs
g6Cyrwb/nZJy8pJ/HxqNFv48L1XpgzcjanYjQWxdMxB1nV7293tm/Hp/oCKYTKZa
O89xMmGK4DtbH58yJWggZRszor5ijQdp3d0YlGZNIqimFExWwILIrkpWMU9DUEWM
bj2rCK582cNc7wF9p8yEvJiMPjX02DxfWobgJJJB3OnVBx0+4Uo0zAoIyqQmmsTc
Oa7scemkhke1AGyr0vBJQFEAtd7wfGMGYQsaT4yPavpJRhFJ4lB5C+nzfv88tJ62
7z9uEfzGPRLpmIHn2p8CELyENR9tklldejUd0JiFrPmiheIDpM241bxQqWb06CLl
zfSyAqsEnKuMZEs358Nv2Yx4/uUx5PYa3oZSuzQvRVi2QSmmweQgkJbj3O2GLmMd
dLGp6RplnRaA0jyBef0qj98YVDhMeSndzktzIzf4vc6BYu2t1LsyqBvzYnHOVNV0
VpCIILvsnxnZ/ZJ/K3VWj/qrpWIv9P8hvv6IlP4Bls/sYScUPFrabd/WKpzBv2Wy
iAlfKmnpP+rXExuuJjQIfTHXkWN2CtxF+QESRrLnlZt7qqjXW9WN7YH23SWRgdpe
YamZof6hMDaGytICMFy8h1hNziFPeas6/pavky0NruwQV8q5R7zw9r9gIFVSensu
um85tbpzQrA3P5V/EQtSY8JgFIbr0EPip5DCY9JBJVD7nAgg9ib4TRmL9uDKCIww
pNAEEDxQKuLB1g+KpdZ9Dkva8N6J4ZwaI/qL6PlVXdVzqOhBrLSE67jkn63DPj74
OOV8p2rmiTrweQgkyIfylPW1F9FOqGSR2TQKjXrKpZ3UxQxpt6TP5+h6MuErVIqO
s5CBLfRUv4Gfm2h6a8iOEsEqol6VeyftgtxkQjIdkamoZOc/VSGoCpZlDx1FhzdP
QlpuGMdygs0AxqPda9B5LOut4bQe8OifixQRFvUXmF7xUL7UJ2fhXneDAr/dfFz0
q/BzE0j5AY7zdfIKUoCv4BD9Oit+kRugcAJ8/KC5fYPc0hHlgYZ7pA2gV4SFFE5m
nGjk4nG1qTYPjHuY9Yg+nu9JexH09nw6wJNNNhhXb7Aq2rLmCnSS/QmCyJ4uxjyP
CJAorCXQy7WTKt09pOGvtbdIRKd8kWbhRScYsCZDerFyhaUMxLhnJfqlBRFtQgOd
BYSk/7Ux52ix6eJo7LSTKvuJrRZsGkaqmzZf3wbiYzkJOtimLY7TcJJy9Goqunoe
NdPDMtE/z49WGdBC7CqxkzarmndV/L1gfk1ww3Yn7qvJF+2v4cVJQvjt224vx50F
kxsrvWpIWY2rSbHN/GD+3flLjT6sT1/ZnFWyrotn+YaWxNBPsfcbF5WeEltbTN5z
eood8bivsEEXivU7qsYEb2eoDfJlod/GZ4kaQ+h8WnIlXNATAiwoUgFdaTjQkmow
9LpyJDOmBrAXHIjDsExO0zGXyv3A7k/e5wCvgFyZG2JChK1EcwNaLkRRgPxjHxlV
OmMBmDkLEyWuKNYhsKgCYkaj+Ym6cjiDJVXmJbYZMbcerHCeqeFnt0V43MRv8RP+
KmIX3Yc9FzbbO/sdIzZbXp+GQfoCRXTVMPa9ZwKdl/krfEDcEmEIcEfTxGDLwlZB
UTVlmZ3pQq7kxiJx5uKSUZSvSEghO8m668d0N+c60Y3GZMsZlDaUB5RtxAKH1RKN
J5NwkogISPSBD9gnw7ehA2TYP2W4eErehGZIFZpA7VaFXYF8Tez9zG+qkkgScz+l
LEyIxEOPE/CR/WhH7aeODvx36wW/6mJEGEX71+qx0nc/Q/rKBGA7VzUogKt528gO
kCXUjkO1pt+LPoiLewR9miMG92UPY6e2oeJWTZ5NB1irJTvQ0epo+fAc+2XYtJv3
KlWbJJDtcsQ9cuaqc8DrFFla4OjVxCifA0G15fcM9uwzh0qbBWuE4arJ+/2oyRHu
cEU7KuK7yLa8TUaDBo3WQZUz9NsWTWNveleN9USTe37k7hhn6tv0i2hUMGCQIZoo
nNEg2vSorapiuvg1LL0pAAYzzdlg3kqp+urxYlVwqt+pFzCjqBdYhMdyaLQh7Ubz
UrYgpXJyJhAyc8XVM+W7mLkLMmrFVM/XZe0gL/Z91pKR1It0i/A4QXReUafo1tAs
NXLWyJPagaTB/W1lmOKe8wAkEUXXaE8WFixaNGM3+oGDYuTBHgwMSYZQKqZVa/Y1
48By7r2ijO6veg5vFbhmq7EXF+cP3zYPpAmGMz74/RUDCBK6OevTV4318KZYY0xt
43smBql1MGoPL/XHRQCql6FTJNov9y5qW8qPK/mvWP+R4eFPSY6x/LPbce8djA10
yad8rUHgS6CM297tLmjfBwU3X2Mqdjuz2cStHkOMA9eZW6ahDXMpFdGYerybbvAp
qTMX6TVkUjDv7MjVd0C995drcmT1eByg358Hg7hlhKRPs3ENNe0USRDCvp0h32dO
BV8vLES6q95dPdFBfhjvvS3UQF1KWC4Zju0JMWL5qDCTl2cV3NBlwbZ19/enfLL2
kXY6u1hHaDEAG4NJ1D25Lsar8u98ne0xVD8VR+MPinMD0fnlXZzg1orvxfXcaLMd
O18TqEGfm3/PHR29kFTRk8jGnrSK4gshWwmz7Y4KReUJs1E2jvw12F975DO43tdp
uSrud7P7zSubooRmX7mV3KOKvSQ35rKHBHefZdRF+nCTJZRjVknYm+8UYVp5LaGh
Tx3KRKgvrattgj7pfm4VG0UW4U7xaguYyL++wDR3JJEraz042OZMoRThXQ8npv/3
/sOkjSnjgKHCYFGdvE+7TR7tN6v2TOnpZ+AJAuwqjJFhWNJaEjj5/aV2o1Eu8Ak+
cGXN4ptAcWn93K75OuAsw7JsqAdndWAu8B1Ks2KKcmiz7sAcYZ5A7HJXkl8/UjC8
ncJpopJJ9KChlJ5NRraoBERycjhYkP78ghxctZKct+/3sZFLKs4uV2OaULXlrVPm
bu5F6NDK75h1iTvrXvqyEGrktPPv8LxqV8KEGHsHeSmmnqPtcblPm9JnQ5Kve+cO
W4Grv8jl08aklWhNGEK32un6WhWSEbcqPrnN5CDDnjhDjpcLToMEHqjReYcvzc3J
hc5n9CueNBBtc1Zuq3baMV/IOUtPpjlaKVt4aaUEBJTDBYxKPZ7/hqWGM0b3RZLa
qOj77S4qbt1XyS6zhGEIjd8bMPwU5brZ5IHAm1tJJa+0OgkiIRA96z/IPBcO7hrt
b6UIL73R72pGasz1+21ibbCuBg3cZij0dG+PK3bzOj6bNMVD0AXqX5l/cf0QW9Ah
hidBdR6esu9AM9NhGPcE7tH8Pd7GkyVjzWZ+J9sZfdTHpPx5dNDXOIwNjqL0MEjf
GfKyWxwhaSN94+CedzRzKGXU7A9Acluv8OpGttdrnX0dI5LaMuyR/BsbV0P0wLBt
F/ioEZiObfusmo05tKpPEepQ8iYRHjZASEuMpufzPgg3HrIS5hHOutzflzx5fdk9
FUQNYGEKcZaunRYic4F7CnwpOWfQBVP9ZM7Plgj9qbUgv0qX0zQxes1HBOJ1UtpR
9wWd8KMn7FsmB7BhDpFW3/+4yr9kw427JsQ1rCTMYXBcgA4rNjpAwOnIMQSj/lyZ
u/IxWCVCNn5cv6MHQiEnMXftCQxBKYIzGfxoAPySFyM3N0eVBoBL2/lZoH7fcqdU
rFJHYYrgRfrVolh9SDrUwNEcBKEzEdktv8qZCt5Aifq3MKjgSwGNvbymSdAosaK/
aEqK3tlJ4W7z9LY2XBVjU2dPM75/OANRFKUnbIBhObeRYOrKuWuNvBNX6Qdg7hd/
jp8CRQo2M9Vr//RvK+pQ5vLAHbyH6f4DzRl8Ou73RNIWj8ix/gko0sjpC+lc/O8W
dUARocM4zXK+vaQq+nJePJV10KmCesP3bgaC4aggpcPFYxUdaCTYsBDbnFSTJ6jt
X8RPGBpfdrJ9k2wJ0CdPb5gVzvGbjqRGjDvaALWjqQZsH0dCpbyLg+jEPCzfqCEy
/bnE+xoZD8ElZmh0wW4ZCwSYL5kcGr//rUlZWwTo6KRGJbYJLX4DusC0w/TR6ohz
TmzbyalEkmnZ28Ie53OAuBFa0htEdyL55Xu2Vd1pdTHS9bpHJIeD6DrKy3DgqXAM
p6FMGXJHzcQewJmJ93g5wHuA6XxCFQcIk9QpU2V39MAlm+q/S8ZTF521ml4xo396
5krv4vEO4Yr4yKqM14KaTRuU/KBbG9orJ9NojOJt8JBiEO5wOjQkhbRE0kMHYYZr
3PakGRmHhhbxueehCJRTTTpaelnDU6Bv73b4VdH8S1Sm7bLfeMWpogsOh5o7BrM8
APEFKH7q5JljEgfMs2Ffltft37R/TpbDdxpBHgjvOmgjzfDycoYBBXVLDTk9i2fU
O8fM0xvtHeUFDeM/8/iA6D25+rcTBN61wjaUn8XP34XyBB5sLQW5VaLHog5ZkFr/
T9xe/K1+RgkvmIV4fxwrvA2fnDNfNhpdGLyCED2XEsp192Fu1VhvH2r5QFoK3/FK
+O9NOFGXCPj+tEoOCO7d+xvzGJwVXwhCthPxB9NQN/Ko7crCcYOAIDlnM1/A9AyV
+4oEhToL+TY2m87j2hg2c7ej2R/ETYsWrlHNfk13s8/o4H+lAH5UBhFtHK0tIuWf
XoqZRhjXH/ympp1lhGA8ro0TFAay5rPv9eGjiOyPoBYJA1vS6hYCMVBIJsD4mBqd
EMIXL8OkkoHzRSZtsYSFDzDkBZP27mFAuDSHHN2pPLanLCYSil5FQU551aijKaA6
W1J9OH7F0b+yY4o46RaUJjw+JEPK5/qFRVjjxO/wJyl9wG4TmR6agXA+Fv2jiHcw
fMwE7+ivzvpf3g68p8f3KjzFcSJ5mywHKo8QUDMewdq54IbK9g6AoYCwmrqZ/xla
xe9iX025+NUdVcGZBxnAzzvdKD19a9NQpowSXgM+Xzy4b9PCqr7k04gQoKAyJ6cg
lJd8fG0d4iagh+3h1T5zEOvuJZnO9hEy0KH+J4UJkAJF7jhvRvmEsTOfhPCtf75k
XdbyPdiMNfdb+1fB0cypof9FDphfvzo0AJPC90G0i1/d6EI5M1rA6EKfz3AMT1+N
gYlQx65+BPeE+Ac5hZGO8Vg02cz+2WQqJFbVXxT8nFDB0uq67gxlYBlTBOSMaKB1
444/XQUkQ8kxw2y8rzElbHv8wtaxtU0/jmG0gyYBMtW4cDmSViOHU+JMm6VxNRQv
MKs8CVwujo0I3/foCNY8qU7gn3m/0dhVfxkIQxIJZ7WUsSiCsKrYj3FZvLVYDV+b
kBthqTUD/pWjaQap9pCuMOHZjLAHzzDcAMncP6iswmuLUVM8pNaQhFEcvLBJqVGR
cyrBjn6ukTmJ78gwLqprmsGy61dcWxoNi3JZ1qZVFN/K8tgpvsTyTK6jQO7nCfej
MoRPAKGgkPFm5id5v29b1KyumD+fUHjr5gOmY5mqYvFi5y3y9AnWFwqskXCghU0m
O5iDwsZEFTSaJvCNvEaHmLKSRh2ppeMY6U0VU3QN72HhOFkn2ovy/YnIJTRC59Ig
85UWwAWgU1xec466Z5Wntg7o9pq3ZF10+3kUMTB32K608sgq22NreMfPwCbqwTqb
fQVfEf4bPv9DSVeailelUktQg/9WMJF6sD23aVslDsnu7EoLmyp8kp2NZDQTQ2XG
LT+7gN1/EAySqwG4/YKPvhFHhZcIk9fVdQS7SZyFCv+BC/uxqRWhX/0qyJMND9CB
PBnnNZi89Rk4mMP8DkfsCBrSw9lyFJFEG1HUxi4IJJJRwIbLn2cx3VkPvQQXAEf7
Ym8+/ml5dxkUEbhD4QiVUvkTZEpBWAppzgk+vY3niVt82w1gi6syX/UT5lOExW13
liZPyKHc6ZhE1lEaONvWVuV7TYo461c2D3+tINQmYHJZ+dJ16V41gG695rEmEQ4D
QGf9G5YOtXXV+Eb6GU9mJnRPaEzkNJb48mQbcYR82O+aV7ynneBsj8G91tw3RuzQ
yUtyvBBrt/megdNy8NCICUeWI4Z/JXAbNogPwJ+pwn2mAuOWTAddj80mh/4zKJoV
FJG0HGnR9veuS5ueTC2I6rfiNdmdI3wQS6xfIPJwrI73Be35lpZBaY2VPCoLJ/7I
Sc8FMjgL6gWjFnVYBI+4eZSDZpld4nitVVMYQefiY9HBVDruD4jXsfBFYMKtHudJ
GdIohvd12z7TWaP2pUcrDtS0twP8HaUBpRqNQN49AlkCOY7GPUguAjgID4wAhUrr
RrN7fX2H6RN2yqFvlHq4qK1Wv7+tLFhry/xxClOSU3wpr4nv6rb49hswBXXNzXzy
JC2wbwZXvAMzyKQoh+6whF4k3Y0Zb9y9BZ4E6biEd6G4dbj3csU61Ns14oU3mr0D
2WJhvVd9xKr5JDhwqwIPuU0WFWhCQJ3PwC7bfYZdODd1vrp54Zg0qPapjNbLU4ME
mX7kOCobCgI/QgJ9f+Ecvt5ZZn5fzk+0paU+nCxAsbFg9IsmgXScSOvLN1IOCh4A
uu6FdN/7gYiOmah19scytI6vO7spv3exvtuzNIkctFRt9TZNBvG8cRwGvOMVumCf
IMw3IORKDMV75sySqpUbQZ+o7Hf9CfQ0vj88bIBUduozlL/tsau7rF0ZKw/qCtcU
9YUmaYloIK90xuNwcxP+YneEj7l0Mt7UY0jncOPuoso6d0O6hzsoPCtoOCrpG2Rr
G2Tr9auZSkpv01QQ2AMEKY1gCaqj0vnusldnlv6kLeg5a+Kvxw3weNZT7xKRvDhe
GbbtxNS5buPx6M9E2k1ihEzacqiqmsBYHLzd00kHJmOyNBKo+fvfvRE5zjn/VUxA
EnmLU3+4D4JwsRAVgilKhK30AdC+jKdsUuMoudh02GSZDJSa/6PanSmZm85cQ3jt
k40dlF37mapcSSdvi1LDG9Zm+9ttQXoCsEOMGj70AouHaQrlHNronaK4osQp3RLD
4Rz7AFG0HhntCGt2ZNPdJsfa1OGtEadBqob5KngxUJ9+D+WM62DT9aZad1apCaxx
4EUAWFJVrLzRvH4qTV54kJkKJTRu6/BaKOc2j1u/E3uVATnmaY/WT0VeKokZpq62
11vP5VEKQw6/8a0PbCD87Zj7Ailz7vbiLwOhicpZuPXDzZ0xUIP7QkZ03tLyEzE6
g1m7tAU+wYeacPn4onWj6aNRYpokTi0xnFqY1aXT91xDg8yG9woP16Nbnl/jcfgh
+4+KUMHqimvLMZdodGj+oRxYxMeW9Kw/SWz0bbZNL9Jx6JodgvAVU8+0RS6XVFZx
0p4nlvwbqcoTV/UdWAjc9NWOY5/zZOY74CnQCIE6XfkQrPHYjO3EndPdjysgxeu0
a+ERdZzvevbXmqFyM6F+HvlAM9L4z9+0df4bLN95ajhQvj8G5ue4LZFw4dRUybi9
sFXH+5ds5ubreWU8Uyit8LYx0pKimRp3vPpxdmIISzUJ/XxaqqIqk91VFTIY1N0Q
Gncv2wWjx6hdWor21VPuWmHewBD4kyI7Bbt//ReY4Z7OEpMt5mUyntLhGFVyPbe5
JUrinEN9fHq8RXu4MImy9kxlMVnYR/eS5ymKGVx0TUMeL3qq3EbTVydCX3PzorJQ
ysm3/W/oqS/ImDrRlmd7UiMPNcmCzvqykH2qIwvn18f6jJyPqZsaXNApPwmcxhtY
5SEJrrLP5NbzxWhOkiEF0ugYV52jA1eXwXYr5L5N8G1r8STcDc5XV4bOmEikdtu6
FwtVlEkMDmbJrWXg+ODcPUxQzsaPDPcyOlqYpHhgals7dYZAK9ggpBbOpIqarHqg
n4GirTJKgv8iNpLbUryLWzYpsE3EmkjDv/ZQ8Fy/YVNfAPR1pvZumlpVeJCzAvou
nOppRPeDB4BMKUW+qlHgMiNz4H8MZ186BF4wpTdUNVjcrStIuzRuiXjRyqTtt+0W
QbPQsJKfyv7ypCuQxUh+6iYmp9UFvWwtlee66DbZmVSf+dvUufCTO4V6/qIfHpKk
kf0LXSFsPH7T8UexVzOlrTepJx1rMTJmNQeaPlUHZH2yftPBHgFHXMUu957/MRaA
Mmh0hBiU0HBbPAJ3VZ6JZ49GZOHTzz2N6jLXZtnmMb2hKspSiFp8ky2XFd6+hkRq
ckygM/dab1qOL5v8BxUlYtfRQQ0OYzT1vABlA68z3fQeMePQhEq7T71x9+VvjyT+
0Kld9kAhBJc16ipudl/9K+JEls206m/MDCzwFeXFe2yKXvx21tA1CZ4SRtnKRlTv
nhf77b715+Bjb2OEGbdazhBiFRBuOn8oG4CZqqf4uFqy7ogSmxWqcL7qRn3J63ya
3+T0z4lqzEKFud0VV4GZcn4VmKgW+AUhGeYj3ZvEJemqgDqJLtPqEPNjYjjo/oQU
tiQsxE+ouUUfA3EmjAtl0VoFFq4itHO3ntXMHN9CQbP1A/TvSlUtPQLqbbQFHEPl
cVvMzFoiZSutujNyOb1hZbln/UK/BAlSXWU2COqa2NVDQ/A/9yOYvhYyPIHb7OaG
BX3PwpeCc/pYY+BbwfNEjHQ5aA6dFmqmo56MyNVrm12IiQYhreZEGYuZm2V9p4Z3
DlfMP4xENaGYi3SjOHcns2dv1DZdKgw9umDkUJNFW90WCgUU/fxWaUBqB/xxckgo
iMB1P0i1sLSIgpPdaEXZDykcz/TAetJrWPi5FODyjRbPIZGFMpUp9d2ZFlw+v1Uq
C7KW/7zOi/sDhLnO+rtvxxPhJfIGpQ0DfTwxwdJMR1DEr1bAfsjc9deouIqSWSTr
AiZb4EqEXqE+wDsF0/Dc6yPw0nOFp/QCyt0APP3knSWzP3TX9RZHFxA3XqSLL21q
4AQGQAnFaYnX4XsTQsJJo/HHvsDWyb1t5ThrMWI379Qu2EA7ASNY3Ln8Yex2VGQq
L2/DNFCLMn3x+H3BzXRgPCistmZviI3Zli5aD0IrAOQQ+s32+EML1T7eaqYP5MYF
JZTqYORh3Qog0g69QYTlaHXoz8AvL62ZLk/566Z/vOMPfXJ5dzGJnT4mkpn+dN1F
u0kWfJtmFiLxgasv3b/xvsXnfQHUMIpI2/aCF0z4TVCVvCjGgj9mTof7yAkoIAlU
ew0zfjG7WYptyA4eure+SLwuFeXAN0nJt/pE353seqyvFg+/rc9BF6yX8OUyCt7y
mh9fk+aBYErfHEzjyopYMu+Nn9PKFoke0vXG7JWnc0P9IWRswxFHNtpHa5zOAZDO
HV5UhBwA+3jiWKChKaqAed+hswLVWU/ieDGi9kAcp4XGZ6mYTsCRCJNPLoxaNk9n
+XB2vO0TmwHKQqzlIl5NQ6+eD5ntFxeF03qPCX9OPSnvjAX8XZECrzOvQgYgrm1J
erLMAfDcpFUyxYx19f5Kl5kbNqDneMGwMw8c60DYhqb1q2dsFHwNefdd8RMuuuH9
ckK9aRmVvuhmBOa5jog1LbMvTGVY5jozV7/qoXprv3gA1vBln/J74426hvlZXxlR
GDSqM7mlPdKASiuf6YjOdaqQ/WQ9EVs8b5mRA5Oh0qFLOB0QTA7c7LEvTUNWUh0j
6O8Ny9BhVnMCOuQS7AKuToTDAp1XFC4cGXw1xOZF/WG2KhxVMGHC4AOy6D5bk6+6
/um4UJXenxiYt//FMGuc3j9J42qgiSbTOCwv5rPIs1u9KRvRqvoMfFTA1+6PrkfP
TkC1ZDF/MmzUuNXq7+cr2gq5JAEf8dOmGQroLZK+pZsQwJbt8joj/p32htVweiu4
B/HHkgxjRlnGfsCzJGgHC34iEW+M083wzd9jKb60JaBZp5RQ92cY8v6tNGa4MshG
+eBKfoHxFRDAQHafk60esKubenbZinwTXrNBwwqW2qE24CTPk9wJdklM4SYeH0Qv
19UEI7+OUNFCDXezCAbspmzw6thVEjMZjUxCw76aVKEI+ZVWW2dN3gD+ezPJuX6P
WMLiWy+NyOOI/wMqZBzopFKKRd7tB7+kmfLXXIkF34QhSUUEhqCVT960t2BIy8uV
g5TViOL/xLWy6TZQfZqluLTuDnr1DPWZoTFPZA/GFcCzhBeSNmuIgxAEG/nENCQi
Qh1CmHn0XjR2tg5tnSoSmm38EGDswSkJsiQFh+EnD6hX1ovKFn5kfNb2wbdGsmN8
gpxTPTDObSARq/8fwPnaJEutxPw4gFN+3a0KsWVr0yg98ZUWrMJV3/8sYsVaaUvE
rH92KdxgV7n3DN8pZHY51eo+IxNyMv5sHy5rBb89xXfVdyH4akCx00n8t2MNlZzO
giFol1nITLvry5BD8f4Iduh3N/EcgH0H4LHkBZJ6EIyNap7w57ZcsyBfI1HcWRm0
zI5Lg0blbghxnc/gSyd0KNAR+PdGf8541KrSYUdpbIVebDae6iCvMPnAqw09pXnW
dpgjD1vGAoy3fE5WznaoaZJyJRoIS/xpCCS65tOEI21fpy56C+vyCwrSC67IChTp
EZANomCgrRZv1HNRlCoG2t0HVMwSdL530kirgURRj0mgC+4z9ogX8mr+5tRu3PXh
pxAKMyCoC7ZQxmhDIe0KK75D7WCdiruaZ3Qv9iICDOUUSCDVO33E9A6v6UKyaMbN
8q2hMghsaAumykA58V5SoOZp+GfRwZ1LYlcqQd4jzlmHLsRYqqRqyzaIo/WUicoP
VF8R7MXJKkWJZpjhHvLXh+0VSBfsynj/c/lreQl00jiZG8BFisIbuBfRdAqTV/s6
ju9JMg7otduEH4a6ju7AW0EzazuEb/OOzAQDyyfzoAPJm6MfIkSTww4f11+Im6Se
3Vv04gBwqn3EeoUvdtGhzCl//d4gCDhQT5fg38XuuhOXIhwhFoFBqklc1w1YI5j8
ytjXqF3zoeaQfQJyY/LToSy9hS74rbeL66zzW86V7hr8WlpREL6awp+9OnK5+ILF
9C+y49R33J+XVWgAg3ecejlzG1g7ml5e6BDnHH9LB2ljHfx+n/GFxG8ilI3qLYMj
Su/TUCNz93on2dB3GFPeEPXEtGDysh6HFLLrDgrHE+VAQ5Twl4KE02Hba1Krd4ky
aUME2BvFMvg7FB+7GmzAJz4AQptYh95Z8pOzgWVJuKMLoMlQYBmadttbEiIXAnpE
o5MU4HzcMQyesDAko1z7M/PL3iU6VFvQZ9l1wMEy2Uu+TofGQqzYOHvmYrZz7OqE
AK+svUkhLi3kzGYl9vC+KxfolMKX4Ax4IEbWPDVAB6hnHke4moqmV68kPfkP6SoN
1V5Vcfb+Egac+sHEPaaNrCCjY0AAf/KSaLew/Pp2OCLw/4ppm/t0jdZbRkENSGr9
besPQ60Nl6VY03vl8zEiCdjo8hMf3fTFuT6iNV31Scww6yroIMZo634Xxa6wWzUL
whhKyDRk3jLYqUsYfKKvLOzNE9y/Huebh1pJWHSuBsMCWiELhO6MbsZ836/6zAoA
mWwNNGegp8pNDEwukRF1Wxb6ta/QVVfK5I6bma+JcQCRCme7Xmq9CB0+YyfxE9zF
fOQML2qQIjM3NPoqMB5fsfh9QJ4PfjPjtqo04rgL4LeUam0mpJ6RJ341Un+wTWbr
HJttK1Dui5uGbCkix7d72zR0R0Vi9VHi59F+NeLodGL68tu9YV2mEbAGb089vidg
462IR0RIcO7htCjKZBmzwGLjvrdCddunWSi2B2/WKyq2iP9aS79r3QXTrpsyx03d
YsHQ4/HnshWYj6ZgJJQVb1w28vthEcX1uD45MwpLA9FwcREhDfzK4X37xQYUQEGI
qWFzZXv2LkGtNjj/GU/VDR/zkTwYmLsNPsVJSFAmeckoXB8133h6rvjiwtQAFFfO
6xV5IqToB/IoPksDwviMpqzLhcUI5lQMRf01/tOsJq9Dkq431OPrZymCUlqXB8hH
5ZHfl4Rjt7d1PhMKfOzTfbGbAX/UQ8HcdSa6Q5tyFY/nb1+3oJRtqLhaQhNjKzjJ
KW+pI+/60DJl7d+FcxgOqc191xQ8sp8bInIv/AnMdtFfvAAIVeEMwqTQ43ruxus1
dik/tGCBLLOpjtvDMVo0NH9/68WD8W/9mZaD1OJgi0CHeOHdjMNPKEpGeIiWQZSt
JW7QcSlZoXFyw6/UVyXSdpI0LllcLDqlbrmfcLS0kI2WX6yB2Z7lTXn5Y8xHyHfS
tjZ8raZze0uBsmNVrfcWEHuJ7NU1g9Cx1cOG1mi1nXMnFmrN+gM8bTjhK8JY82oV
c9ouoxS2hN0toqwL6ppfe3PfNUr5Tz+uIBPQj0azlMm+fjkwwW4hYvmd1rRvkEog
BwHR35pcpQBpr6dYkUXb1xtwiIx/FqT/2ZOOksHcFdUmksAQRNcHjIeNvMCaOFn4
KrPEmQTE9yEyGpb9fvKlSFWmtb+vIoxpquaB/nfdSiyGIsXaMsI8EN5yQ7XcLoBd
quIJ1Sxfwzbv1D58pMF4cvqLErnVYINPZXQ8uCuMOwB/gMglRNTdkT2ySzDCyvWP
YdYv1ZbxRp/rH0lbmqe1IxOHxgCN3BkADrMr6jidMaarZ4gUaSmByi3UCg97DnD+
qMywxzoElo6Nb+AATkmaOOGFtEFJYCSMQ5FOTbPpIaEGRf1fxInFIKS/qH9hKRha
jQikBFztESn4qy/tElVq/ZAtmQhfq/FNMib8IHr1Qql9jAUjNxfrpQAHzZgqMyHi
bEnoSwwnfdrgCj0JRHkruvhY5oBjTtwBwicX57uMaBZuxL8WjXiQ22k6xcUzlXvo
c4M4sdiy6Qf84LACr+XeN3g6g+W05N6SBFOY45mYz1XAIs2lQdR+9LVLzno3Urg+
we7BKxpIcvTYBjstqQuVML+f5d5iHxeG5/tNXl1e3kMPQIeSH1ssHZjiNEDycwNg
G4lm8SpfibSYMmzHYWZbITJqw7geAhcG4rh4fdJdMu4jRt3HmymJjnrWtzeeIVDf
mnY8bkkreI5/sBA0iPMPwxEtR8Csqm8eJcgeMOe8KEnwl1ApBvlVj5fmZy+KQlFt
Ph6oA+lCTcWAsiemfHZNCUs+2F1DWuGdCG3uF3b0McMnvhPOb7710wEDinw2FYy2
vfhOvgtEsHMwpXSZwmuypuv+jjoMJEP2lMLmyXe8IzEtn3PGeQL6z1A0YQfTA7xJ
B20rpwLPrKUu6gkCftO5Jurxg/H3Pj/2rfvKKIe9CyLh9//+JI8ivfNESQxc/ocC
U/otAURrhJLGZWM68WP/qY+800Yjq52E330T2VGR0I9m3WQv+ZrTsumWdWqZuBaJ
/l6p5OH97rIt924b19jmYs8JbHMHieaer+fhBii988t3xqHEGoObz3deDiY3S/UO
vJpzrHv0Qt8zbfKLwWtIs/5btPB1ZrTBKcUxE3xOzWTRgWsntMnOT9d9p5cHa+GV
9MzjBfHqoy45voOobPexXXR3fY9W0hghsAuU5r5LifKoGbeFJuQGpj9q+jz+cbuq
sih2eAq5SY+4cCHDFH1CdJxm0PwNmFUZHlGP5PZThsUiO+u6YWmy01I0PVOEAUqU
q9V2yH1o7PaRquW9QNBSfbp1HAE03FQTY4WM0XGHyrDAHVPk5gGN/9P47kIud4BY
MvuPFBB+VH88AvMU9Mwqyh8KCggvZd2Mv0e8NQmT1hpsodMybVqFEFjnDmxHknKQ
QCJwuWliqK+M6VtKAGssoOtDmbILU4m1sEQ3QkcFZI+6u0HxwS+TNL5VTN/XQaE+
Ev1yGx3VGm37sXHzR8IJOge9mfWDZKnn/97/xdXaGzZEc5900TKMK1ADgwXL6Oeq
fMYvhGyTCZcT9bSEHsqjfroWRCi3DNF6/0MhnDONFW9Cqd9m6RAVJrFfb57rqHFG
Hdo3QBaIPYkSG6Mmg30yWCWBGxzyRriaQbXddfcoc/8k7aKYGg1wnobVC1cJZ/CH
3qnNgo6NEYIfv4YZ1ePqgc0qlMkh37Bjjk7BzY60GKU/n89N8C43SmbLgX5nmkx7
xPUvqrZWOdHiIKnWA/eKF0KgYoG/NZBIIe7eFYiPJctTpNUe6FrQ62HBpopDxs1R
iy224zv777K+OtpFgJbE13Qhz/JtMj9fkbKLZzFzp7fmHKzocJFLlTNv8VI57fdA
gNxWVKVpeQfcUCg/AKf+KaGJu8X5lcW239/Or0W66zXkq2BowwBWniwRAK2U4iV0
zDZ/KppTUAGZMPPehePU7pz76acZFVtFRAi4bjp3tL7LQZBy/t5/N09sl4hZgoxl
r13vwoBtlnLfVn1zCstBp/RW/AK3me1yGhsDlCOr0cS3UIqD/ST7V7RmxMNSpRtM
sIlGAFpR2/cKy1PW2j6PrzdgQHpRbEfhzbRG40oYnXFg9g47RXZEnpFsQPE+mc/X
Kgrl+N3RufUTfZjcccQrrdYMuyTjyOzD5flDRIExvOueG0syCbIkwqkrYIEMfexb
SyGauxpbXJEu8Nn/NCK0Yw6auBj/hcu+v8UFA0RfaVrCRwImHwSMg0i3WwINpJ9m
W2VqB/n87kwagEXrCqN+X773jlwlLQkbWNx5r5Rh2mmkLkpcnIfVz8mFnqdkmEXV
B5xvgpvkb+Yb8K3rlKKSW1+vIdodTuMFj1xKVgPxN2RmRzAQF3Il7m41CpoTvX60
osOoR22FA/+kxwDhDL4LurRrTliVPWDaTciRoZmtKfnsNBlmQbl6bGuvpkg7i3z3
JndHyBA00Tn6dzJWx+ZJNFIoZvJ3+dw6Dyonkb2NdR65ynQ1msY5vhIykyPDSGQB
yzMvjAYCP7Km5Cug3YnWgRGyUILnn1HFfQs9BUWAMN51oIIwgSlrJ9t59M5OPfdC
70NgmUcUsUy+RiM4o/kDDiIPsVkhOyznHBe2TP8+Ds80YddncgT8vSIEkdcgA7NY
Q/+ETz6OfVrXYYIT2Q16RnoAizWwUUIiKKaspOZmGI50d/DgLA2rFBaaHmyfA40g
KSD7LdCvu34ud+m/QvszP8Mgw6saDbgQhyx9FC5I6lkyQE4DHGT6KSaFoP5Qzn+L
14hyacjv1irKJEpBQE1LTC5AJihRzb86cdecYy6RsBsqgtTucS3T6P/7zrx7gJQE
LPostXPPXdimbFEp9ePItxEYRzFlv98V6Rx1yZHcSO31UM8dYck94vFbOMUKITK8
w4Pmpe8gJT/keaYA6aI6ad9EXrBFSrtF13sMx58ynH+6TWVoIwvTz8nZEbpTJoKi
+hIwadflClEEo+wrISLkiLDpD1DEq0xvMAzuUvS7TaREmKbG5L28KjVIBqpsrpmE
hh9Frp/x0459Ou4RYLK0w8WXT8rCyyWfWVG6GdcynWMcvy5tJLZ8Wcz+CmvarXev
axSV+sAlT6TUrRp8BDDSteRUFKxQuYNeJpNzPWJkxwjpx96fhzFgn5P+bktcKpUQ
5gec9a9CVjfTG5c6DRQuuh/BHvS4nUE/XNuYXniQQUZMhnF+nsdwTpbOBWeTd39e
w2pNfP0Zv+O40TME2d+neO/CwDgqiub9H+8zumfUR1kGoXOm1dwnk/R+EXcIGF3X
ypTKG3OySJ10Fzvo3VU3S8VCIDTbzmWYQVq18WIiaIsGfhP8eT4Zy7ZeFpfCO5nA
aw4ua8MN2xbSOSZ96yOJf8rKneyEGFwWZagzX0FIkr50UZ5UCFYqspksl8J/1jmL
7AIP+LZBkf3SRR7gQX5ayj/2xMU0sz5eTaS1X920uQvPkh/846hkh9Re/uhfp2gv
n8mvXoja6R58ymze/gLDsWuvkJf+qdTSv/QnqzAPZfFcWInCx0dpK1XCYVeUxLCb
Vm4ssEsscVa24LnGOAuohrwSGLmk7jAbxDO3IDX6bOj92edBSvuLdtIZzYU8euqH
JYTUdHItihkuXrbHZnOe/dlj5y2e3ClMIaz9BJ2paxEw3qDGKVAWOXZ0lkJ86lLM
X72n81qOXNSyV7vZ+wssCBIhlipYXrH1MVLGDhWbhaPEZtx5AamnEkMXHmrrTH72
Tzo5smOWBMGp63YNEvOnmVaK5Qj7j/7WV/VHHFT8y/S8sT9LVgqb3Wcnc9J9dXPo
POrbPBLvSm+eBXaOmuYOeMFg0sI5PuAirzeV4VaP0Q0iQ6ZPE16Ic6WrktnfD+NF
cUbtyLFIBzl3fW/uH4+0gqIgnN9jBZIy9Y9E3cHoL1PbqAvA/csMMrkS4WMs3KJz
RQEM1LXhqfbq/Q65UAklnVL7Z9wVf8bknKsy4W/ASl9qs+BKMDZNtab/dDpHJsKG
Q5Gwp+Y059ACW1Dj3D6NwJNkzew0FDEaOgiJwKBMy2Bi5n6qCRngN2tmfIwBm+IE
h1VOw6fKhKcY0m5JNK1+yx9ZafU0kSBXsMFb96wfdIWL8EudrVy578pB1mQWDQ0o
ihWY9ce8SeIrSPC+1NE7PeXqruOjSnu/Xx35WLgBqtWULWgYQA8mKF44nAd/70x2
1VKZWSon9df4ddPphMZ2O8Iff8CeowxBqYWw9mGq6quEql9yIfVEdFof9px1NXqq
scgYU3HK7i88lfKqrNquIDue5uyZkSYUXviL7x6I5ZU2bhY5W57tyIVsYMpuzBK9
yykMMusxlDnygivaSKy8HBw0d4JXLehVVw+TGpxERpOo41uF0UcNIgZCdEKAgIA2
Hns6P+hWIEvmAo0ldqEirC95UOR+AMMy8DA11k3vGn+FVKsqQtdtzHGK3M21aGRz
M1POYTi2kKHmL1tWpV553dlmEQ5iyLYkRjlAnr8eB9AItNkDCEAYdOUfD3XhntrZ
SgqI0AoQeqmX927UkexGIqLMgrTqzrXu7iTw6P3SlemrzpQtHn5AVYQm5HODdhgk
shOF1bUpCybRrHwbV0uT7vABxvJZEp1CTWfDtuIEQT21eQEcTNLE5InpnP9X7eqx
gRDDz70HdRSwjQFvauKndEiBOGEd3VHsmllpObgQNo6pvUaRyUkFCOjjE32DnMWK
4XzBjoZZOKwP5GheJyTx1iEZxoxjWNlOwZb/f7JVtAQvBn0U+bIOEX1mRrOwRFQW
O7diQP64WM9Ns2/nTcEjK67Y5AjK1h8ZBjSoY1ul+0IYRK+yPhF6Xm9024UYhy5W
vI+NWY1zyQ++KyDwj4EP1Yq11rIRK+SfmtXEuL+Mfi7d0D+owXkF5WMeYZFRwNQQ
R47AMkSBkznfM9Eb3dfkp+OM6YN6dsh6V/MG7J6ZFXY6S8gkUVHJxSxKDj3aoswF
SLGctbH0MTG5+IJdYi92sUghMGcF12bXuqfWO1reu8C6YHDOCi03U3YEWBtCis1i
laqywOSV/dcTJREE+qMskXA4VZzuihVQSOViiQcr81iwrozwTeaHNuV9uy7MXuPG
Xwwz60dH/v7bgw7ek+WRPNOEMha2iMhqheyKiuc7YV1oGeVu9XK+zvp1Fle5XGDL
j4aW1GCnOub9inVqzSbdFjUNOlZZQaDvASfMn1YhjEOznAzwfrkm6kLIa4raSGy7
Ej3xgh2ekREOPKW2bBAUEcW36YH//yhfGQuyVkQbAife/IRisqOHtV0ZS1DUV2Ju
ZUwspsCXDccB9sNxalA3Se344Iv7z1ckAevW2s9PZkI8hPUG1qL85pzdkQt5QYIO
LHeitRIhOUphG/7h9DUXYSQ0hPD8Yx67vL2KeZ+aWSthuz7ZTj4PbUHty8zna4DH
ARxH9E5muCKTjWPG7p49AfuwMiFwiCZZy1Vcwfm0VFv11CbX6sX/EriO8xfi9TZ+
V1hTWwse6Fq5H48uakw+i6R0XnqcjPNsFHbuWLVdNwlirttoI/qCi3AWtenPRdlY
Zh79tZp181nhgA6j/tC+SNy/mvXmkOLsN1IRWkVkR+i1T4nuG5lAHNyU2wMXMaDd
9K/rzqLhKVd7Ki3jQIbiHTyja6KuI1b7Wg+INuqca/oWHE2ADsk6BM1gY3TZoEDA
LwFkZWSqE9/y0kGidg8HulwBgvyJ0e6PKF/P0jFhTxfmEss+aQw54Xg+18Nj+MLZ
dKGtaVWSQc6w54HFy0CxqYAgY75X3blqTf/Pwet3h/pLF+4PaIJZqaaCjICUbqvz
iGzmBqM34IxC1syeAhpWdxOkZy9MstVrKbP1/q/U2wMuCy8rk3rPeok1OhJT6d6V
mAIVOYRd4oYBMAG6091zeL2DhIhs3wlrF0KaA4CO9qDxHKwuTl+nc6V+t1IulhUD
lMFnBwflJkjC7pQLLl0TntHYpBYTERWNANTZmThugHxqM69Pu/J0fPQAxrD6CQSP
pPKLJMTgymLD+XBSov8UVjCdsk+nfYQwg7XCU8CctpOuSvXaNoSXx7hAbQxQuBAJ
wMs5xVhbbYjjwL60Gj0brIKmZA8qtzLDamzQ73PpA10In9gppHUu6JfJVJoPuJb/
ok1OdkH7fGPIRgJUlKuhjypMZl2pVJSkLDqkFIx6UMLtxeVEmElnkQOl4W0Za6Xz
pVqZ67IZA6Yh6TCmSNv83f9bGkt+ws53UD1YHY50jEiRS0DRNyvWzfX8xU+cEqSa
LrZbgV7XfXDrCHJxjsZa0UuObEhwW14PwCk186gBWF7M8SyPa+F9k0yadshNGulc
EMYlOsS08ziDZ2lb+cb/48ZEmFOng0KBn/70FQPiLkt29hXj3lB1Caxbss1RUIqr
xYwPvEVCnywAwEv5697y78koxC+wwANfvku1b2XUy0SyVaMvZbUPT+uEoRIRLVsj
Vy9AdC/q5zakoYu/wHinQKsWFLdDfLLQpxBP/nj4Hljiw21yKDjBWWApC1KzMbw1
1NdRShsAaWMiuQqLn1Pr4e8RSFUjK5uuLEr1qsOgWEOPJwowfLBevtbKr3MGgG4f
S97D9VWMDXlV88Kzx3YEuumgeyHrY9cidYlg2TGha55cqjKV7t9Tt8/N3ZeFMdnk
qYRnjhA5Xhxx01Qh2OfcFf5M03hOmDWF1bGglCBrgeskKWRZkeXYeuWQPDWcf6jh
Go0SlETJEHuOesxQLa2G0wym4GvE4H6mDDxATpUB53QYN2blSzpVwULomWXinCFb
hFNlsaEPxHAD3oldq4i7ZuthY+t/wpOD78pNZy/Wc8NJo4lqli/hYJtQ8xZyMEqh
qWzLXP49BLLbRcAP6UwnDkE3uMd02J4mRhC0dUpCkVS8LzuT84PKPfd8bIQ9NgJy
8OQI98KJ3LMHLdC6CJft5hURLZbeA8KxmRJLw6I6oPr4ORVMIJZWjIT8iYTLwxDs
gyGhVs6geuFo4gKBabxoukVOjVFz+0Wo361PeVrVeXKjuW7zJOs/pklTNyXRka8B
pektX6otFbFtwQ4Ce2yx6lMX0q+VwbNLwVfEhUr4FN4VC2jVOwqroH01k91YNRCA
0cTSvfUUdj2rmFFNclxogRlWK/PC5LuzkjwY1qPRMq9QEhT/J2vCvLhMmTahNg1D
mmE/MNTM7/VCmCAgC5o0R42SSIE5qoLhDDyYULMy0Z8pw+JXotfctvb1HWfZQP6r
JYu9IKMDmhtTK+v+v36trlfOiX3u1+uDcnmrbZxk6xPD+QACrLtsB4EhAMWM7YX9
G3M3h0Qcv4vFYN4zbXcbiANjPbpBoESUg9CvWK4V1jN91l2fh7SH87iW0NSkS3cf
W5I10PujN5ma61LbEZPW0OmloONUVCnBYQtKi0EBirF534hF/mQ+4UtDGQlzs1Zq
qt64Abj7MDVCk6HJEMHXxwew3NS+otPrUfiCV+3MkjmAKu8SGiGByygBzaj96uIm
HeiePIsveaYCIdxQP1DzDrZgfb6kNGJSdvb6e2pRct/pVYV9LqPWkpf4hTp4OsFF
s3qH57dadarbpl+WSGqRGNxsPpekVOdNWqg9w9/jYFbkdRfqLfPCg4E8DS9cpsMP
pGGALKoRhH0eNb2m8cGupezTFqbZm4lbpb55BD1I9IfZfgbXv5LQdPe4yNwZ0pTH
tF7LbHqIp/bh40P8X+P7QvhhJ8F6CFDCMSubxtHbn5bkWaYJBz6S4yIgx0pj2JDp
7zEZGLBXcF1Uk96Ez3OFBidkZ4cNL2xD74BxWlCCFMv2w2VvifjUAYrPkX056t1Z
lJxvOUKXT9UdK9hlsF9RdLI9NxiBmPsljTmSR5potXh3x/KRuH1IrK/VzH9y5yH0
e9i9exrntkaqb+v8v2oAIcYt0sWRt/v3p72DUqc1QPZ+UuuFscaGqHNmCzys59bd
cXC+nWAVobCs0zpJAMIwe4wOlFOuz4jvHOpby2Qh29v105+YcwgJ/daRgAuhcZXN
m0fR7B8NiUntkD143VJ0H/I6bn1BE2SL2Ei/rgpxICM4qoxHHpngBguIehQxuLUV
Y3V/Xwglu+i+Is7X1RCJvdnrS5JlaFABpgeNH8kLLdBIOG1198OBCAFPsMISuK0v
PIQ4PBXdvC5fE5cHulFqjGrbmkNedpkibjtXYf+uoijK+j12bMgK8qpfEDgddzZJ
Pxp9JHAf+DDNqBYzuPLjV8tDYGq1HEq1PcevSudGx83K+BSol0OhUOEo1dIDvvb7
20CzF1gQV5ZyKCk2OX98mWerZpsXgX18TY78HIGzPTwn6A0uMAW3AlnXGgEqmSJr
zJqZvd5hXYQuyBx9d7Oli1v3xvXP/YrecQcXj/XZq2yJNsBpTBGR3V062xFLJHxy
lLo5YCUqI1R4UZaLOatqoIrN6zU8fJrmxHVAvEOdayp8k0BIdYwxifxppAZ1Tl4H
Je03boJ5TzoY2ou52pIlYTGcAp7iz4rhmsRfGEuhCAd8u4rKFXNKh8vrWgLhF3N2
aZuwNMDE/Xk/yAZOD2UaezN8Bk+yB56+yRCrqXhQZymvUeZQFPOKf6qdkx1U9THr
9RtSQh3bY7XqyQXLHYMQEkYp0UsR/Gc2aa+85RrxDNMjMzsoELQn/fjoQ+wALmHT
31OYY9vNrXXr4QL0ziHLyQhRdXYbV2PXbuUeMRVm8ut5DG4fbHzoxybuSrzR8G47
tpl2VKPsbijZ2+NaLRLZF8HDSu1klyw03UGNCuwxR7eqTSK/fZYQ+uouYN2H0DEp
kk1cJDqzfqOAR/iDaTaL0Lrl7z4NjzOvZXROfiRcPrJpv+JOsEKgTILu0+rUTFOe
0xXXYG3bwubBjg78qQtkMGelwMsN7/+QW3CSCUoiwnvSwYwFgbbOL77Od5/ucz1g
ouSh0UpI8kxiPozMkSpjWnTRBPlqWMfzs1sCIWCvJORShm1KYXy1K4ZbcnO362W+
QHfsi6DDo3/6ZzcjFVFhD6EsQBkH3GB81ab24pPPGsOPQRhJPMeqHBvc18tRugG6
RGohwOZtzaM5MDd4nG+MAKVskXubT+r9EzG8NrdgIg8+PZCyH9gw/nJ803Ly86xn
i8mgOPZ7TQ8j4bpmvmPKswulBmEFeKDtENyU6UsY/3xgIWz3rWY+wBipg9AiS6R1
T5FYq4uK4pVKqtCRg/bl4S6AJkzvccgGNajFI0U7gfE5SBzgXHRabTYeQW+Ylu0T
RXpNTzFsNgv5sSaq3CXgnPztsIVns5MYImkhxD6girdO7lPKLjZLsvh11yWhK4Lu
6GiIq6TeThg/IIZCZ2Mn/HnhlQTFNFQndPbUquUAXKuruFbyZ8S7sBa1uaPGNhoO
7BLPaoWeMiUQBOahv1GY89Ha1PAin4tX5TBFcxRtxUQNXp1mUtOL2MGW8+kdg25t
KJwyLT3zJTN8kaeOVYWoS19txkkXNt8Ti4AbvXYRtlBeeMgDf6hYaFDILtne1o3m
1yPhHWh0KFNaLnaWN2ezOM0jvyy6z+KPDZDoJcSjNUghVPnKmz6duSKL+ccpIUUZ
bGLKWkVkzXGbizdXBvp4LjHdN5Ez7IWBx2LqYIXokojQ+4YeKzV/Y0Hrd3/e84Jx
jiqMBtBwAhC0bfk7hqyEmlOZs9+RcrNxGRVQkggNetGpv1kzeqnS4fIdlNQz8RWt
9B0kKX1nwb7Dtb5b23qd+OI/hMQkS1+y1XfLUEfsdB3fIGtumxzmGrupFwZAUKIm
UB6JFHZwCEG/bh0qsXhr1jtjiBt7Pd0qhYNL/so4iiwJpeOQU/k7fvC2vpnPnUph
l1/5sBs+XyImr8gp0hvT/gh/JPhqH/cUZG5l5Bl1GGm+hVyIdOtst3W6nngoEU0T
+xqHNUi28EXPF4aK1UahpCCVabiHy/V4FqOf/0BGeXR7BRwGyYBd33QMD+0/kAvh
IyZI8yCV/aWE/8zJVJ0Gwz9MWvz+0c+Zk8rAmbXyQFZJJg0Ft9LDE7eiWaRW4VMA
zlbd1jzzadNp4GilLgwDt7e5RyPm28UjiNR8h0z1UjCYjN2OrZ/zWoIPGe9HAsvL
Xjv2WNTv8fjcFVLwtYiKPfZDxuwV0ovcpO1hEoRWiL0xde6uk/KqZFWm3TRr9V1A
3j3StItLl7SNLWNXvObEMd3gYga1TprgnpNX+qS9YotSrl8yP7tQnsmiZPiytOJR
DEgx6XD1p3MHHZwsnxWsDUVgnr3gsgVh9LvSxfzWdox4SOih6JHAIJibj0JrBx6B
5va6w5WPjm9uUz3BnlBmBlUZZj+sIuHCoYeTGBWuE/kmn94lZtjAvR+nTvyAi4z7
H57gzLdwU/zZ2PwZsit8ZK+nSojJ1eCgABrPJ56jojV3P6tKyXNENU4b72sqVCSC
0vLEd7pKi5ttt9bTsXdThadaq8tvBTuEfHhqII0q2isaVBjlGDjZtfVt92u5KP51
4GxAd6no9Iu9LVl5AChabnSEGJ7bnUkRba3XbHwYJ2nlKEmPbuOu1CYgyiwrex2F
2XjERg2gV/B46IVcFJ6VfJNI2Z71/c7L2WHo7QeCdQQwXop8WsUcA/btN0qmY1c2
UeJirACCGBLVc8177sWjxgxiOgJpNZZZvl6rV0oUM/iUiPl0zLDa/6IYbQx7PQn9
6j1+q2XgkS+zO1aoYcc4OxuYSlqfTfLqkfTPVzpK5YoiQ3CBtBglHhDOT7Kq9JkG
SPluE9F4WZklzHu8tTuVkTd1EdWNClHPgg7Aa6a0sRAiogX58yFw5F3S+lguzy68
dVHk1YePkCQIYu+YyNDD8Oo8c947LRg3Gls0WkqUDB+Wa087VcS/vVbJn+MXEZkt
s3DyR1nMrSqQCKpzyVxqPVz9pgp5H6yn6iRTw26ixf+EbFrEEhDgUGG/WrOOuuh/
xFuLQFR/Osah6KY58N3FNGLDhHLiWRl6pENtNwyQ2unYnaVRyTQlja0HeFbKIEQb
ETq9+UsMiZUPlq34R4aZqs3i9llqawU3F1X1DQNLgBcbcz5oZNZ8sIfmoee+gzM6
+vGysy3qfvvumTCg4L7p6mOw2VTCiEUVS+s6I54v5B7MMQiSPord77KeobwY5mVV
JKs/0Mt/uj5L3Pbhn730vzVFd5I38ymRFRqMY6TqsuG5NijQ0FTp0KlWavbnJDJ/
QiucCit4o5sk11cZ9YUN4hkYiZj5Db/OhudUKK41hUIQOYuNdzmz7FUvGm+VerK1
TO5sYvZ2n5sZB+c4rZUKyIQNVmt12BI0DDaErKzva0HR892hfTu+zlKjtZtj+i5b
/8HMHX758UBHg1RrgB3Dtjqo8lANVYoMrfy4rni1eNSFt/fIammE+VtW3K8m1udM
gFXNrfgqWI5kjTMI1h+Sq8PqAZkLs4jNJXdkXBFmjp3v+s7YDR/yD4BbQ3tREHVE
VyfeyB0Z/dlD9n2vPtqwakbrBGCWndw53Ahl66cM2bR9bmXo5Rk4PXtz3s4QZJWo
1l/0n9C7YYfh9BZCrfVmS9rm1HXNzgwJY6MrBBdvlVtVxg5t+fNh3qGXjqJPFm3H
gGf9VipIl+rudxCnQtEXXymIecDqH7BVCIuXavZC2+zT6vf9aSIT0VUx3j66qEfv
LszoGi0E4VJQB4HibWjod4j7Qc0NSDCdIjRThy9Sda/cqpHLTw4cxMiy0OLxRHWI
DsawqPfjxBf2mCajPIhdSXE9C5lEQh5XtkREyau91O7xXbBwE/YnnkZ9RL2rOjsa
iGKZlPOq4sbNpY7NqcUjrS9k7123CWYQ+BBAHk2BrvfreVq+84ytcsWkePaodcW2
Wxack3gW0e7lVEG6N4v/c+n3WKju6RrfrHwiGHqkmsIph6uvLWzIhQxy9tOQ5+S3
C9cSMqqEU066WljGu9v+Rh4Hxviu9Jsc4g/Q0e6FUHvHRqHpSaVzkAyG7pYyaW/t
tlkSn3FoPMSCFSfJJj7fZz9djOBaTwqz1Kc+UzSmuOLgdzjV2ik2HeFTGDFhYbbd
1Qy+jat/PxiUPL18evNMP0L3U4VC/rO8Aqja6v9S731071PQioVeKrfKbnPMKygv
qUzWYUEiS3UPFJ+rds1MPRxUObVijRqFW0lYA2OUfs+bNFpGfRGg1AqAylJS9CdU
K5KlKoUz0+0rnnqv79HG083TdTWPIPnQxMQscsk60fOBtEY4uqP+PxPYEjelxHcs
pWRE27X+q5GFKaBCJqjU0ufY185aOpHYdSt6ilPVQzFdDaykpvAsH9zsn43S0Wuv
5az0r5uT0BptHhYJaJg5CDr3Cjy+yXLdUjGRuR1b9FNVbWJXeEW+jrG7vGn5qNmU
1l0AeMRjvAqs2d7qID701uPzfizSV3A9dj8AWoc8kjIRCkd+ILctFmdPs2xMGhTv
0M/IcmnzFxtdCbzAZN8+alyysDQP9wkELJsuDI0AyZBuxmL6amByiDc/PzCQmxIz
6lyASIq1VjRVPZSFDE9UVo00zs5waMcQe9dXsIZMcvav6jRFuE8MEMvVWe4w13xo
A/9M0MGrWJZFPB5l2tKR/IlrZ863pbLZutYw5s0tv0/dP2WNj38whruyx9Erw/hG
iswuRhqyEX3M36OXj3U6lUmX3yM92KmCcXrIS7DsCLMNrSt8P2natjNlECRKDegx
hjU1Nei6cdx/Tcq1XBztwSq7sNkzdCyJX9wkGD5dQ2KQaF5s0EXUxzqqJgsbADxJ
ybIljB7md6oscEpNZahcGR0L8CP3HPRp5S1lz3pDHu77Otr47/LpXBYyrUi/hA/Q
vDipWoMFtzhmEEbHJ1XCKd5Oucf+wSkSXRBjasvpXN+lfAA1aeyPhU8im8kGNtS7
OPgOyrvDeP/WaDQYnbb4p5pHIayGYHi1K1hEZ0GRDOCQqUNd4joeQVaNxhynVT0Y
Lnt3bitPv9svn/FkfoJ9TVdT29aVTGYWWPXP5bXDybdNydNos9sAGpqIbWQV1T3D
ziH+5mjA7kpi5j/J/qbqan+InAAsxhP1TOfCffuiNY8dmaw9mxli0UbC56nNNUjS
RDjDe0k4GMGYdunRNUKKjOSe898cU6R8ALy8XKGV2yxQvo1mwDG5zTWrRimz0QV2
8FbVI3qRn48mSlKG2lMQrc6GQ1EfUOPjPxZnM8Y8gPH5Gz5KODaUtKWERnCmp4HX
eG/RkMIXqgG4WjSf8gjTfjdTqt4KWJkrcZnc1GAvsXZDWED30r+FCuUdHj2F+9Mu
11v3GO/6vC4OOWHG4+yGS7numFlZlRqjVMstWhIedEyplMgBBAr54B/zVbX8814i
KoYT8/rMwf6uMqyVJ9bduJPJ4dHisE3z43/jsCu54/EFSIuUGUwJgsZHPS5vCvZ+
f6dlkLrPDutO9RoQ7WIYopQa9WhHkVOn42JMDwMG+qZP+Zfj+5rIq0p3mJKlyWs/
2u4JEYmn47ME01uxJiRNijszCE840lHq/eP+erLCydksl/1Zgam0odeV0P0DKZIK
wX+tawYgS+LyypR4yzoNmC3nI/srb/P0ktxwyuGH6R4usnpJovPIsOIkAFP2Oil9
VBJYBsXqfLxZ+QNr3KxYmzAOJpThX2gWDsddx6qO729cUMsA1t8KbXx5JmDwPT7W
I4cS2upFv1ua8qOBS3g33qpVC9Z6aVduvqmsYhVumq2yoHZU6kfa3LIvI4e1triK
2Zd/QG/nn1bJeB3W4SVUQWFbnlMQF8nPDkJgU0gbpfYvXeqNOL0d6kUu2JxF75eZ
WJdUjA9m22wIJ0pT7t+Rs/Z1qzL6i8hqQtGzYzXjN9NGNHqSS8+Y7QfZ3OKSumGH
NWqNGxUQ6vjTmwdZ+VEWBGQmAh8JfdNTk13tdDPc7qt/mjszInMjAePwOh+YMr/G
LRwDAh/eIQUcaH7OGJNIEGHQjqNobMoH78hRRFU0Bk7fycbYto5BqiXXtyBO7z2j
h/Jjzt/4cT6KbE/O0TmhCTD3FBFGWy6xkNq2iGBBk7xtDzkOBpqFA5iKScPBBNcx
tUrJdQhWV8xcMC8EF4Fnq8z8AHSI0YHMSILcl+vpvjsATEwczaUPlhsMop/0WW+N
Nz+pvZ4ADGsjFHcDkYxoUAFpV25WCsmqf7d3LXmwn9n2FvLNXfB1W8vz/TX25As0
4gyxOJs9AuZr7UL81yjGwfXOo8GDNrDjVXkDH6I9weYRpnP8do96+maPM4mmzcYG
Q5UVtb4iURqAh2zVk9kXZS1xqEbcqpc4ZR3JCJy3YAEfqc3IWLv1qH6AwwAfvOAI
zVahumiGn92LerTtDiR7lgDO26kroV+4cWatpeVj0hTkSyZp3cmEzV5GqxsQvSM/
jdYvBUTDXrYBJEXb78IqW46VXNeuilZHwMP3A++gdNw12oSWOb6WU3IYzwWag4lK
+fOQ/aaIsov5ajxP3anJq0FHoNHSYJwf71RZGV7JIOI7SFCuWd9XTJdLLjFLiImO
EKkuxY0C83KSj1kCDNYQKtpJiHKs0iMOVjQK1urFbQLJGQtL58UKEh3wE/BtG5vr
1e+MKw0JQcfTMkWY0PaDXQWXnasdi6+rv+LAGMfX/sMBfD3B+eVdnL1kXg6J+3oN
unpE2SQoYcoxR2jZzDpS0An2O33ecXsjMHVUwCqpccqwPgCOlc3Zi5rlKGsbZfGB
UdEPfu18OHHOQSNxG+9MIAA0imXRkK4KxGm1TwPUqRcmngg4Xi3T0SDyhhmRjbR1
aW8k5J+qys/aQSlZFOHDfoosWE7gOHUybJsM/oGzysaBfL+U2sh5bOEUkw0j3wlC
MAneg/xKsAdYwjctoyrBgtbHamKAwnevsSEgwLRzdSjOR8IF8cccQHG8iLUtgR3e
TVTnOY6faZsWz4R4WwJk8o0kDMW9resG4pmCjht/odC4v7yoaKLZJeR+v21hjXrX
uYOi6AEfeQsB1U7adhMLgHBytveejNp9lvWQN49UDqF7YfduMwCmiatfHRhgiryC
dWFxqo7Ilvq/DysehKP69SxYFNyk6m2KS2UdSgUHNIwI1/BFqtKERDs6iB2swZ+6
FYUDkoAxOifG9PZr4O+TEnSplQD1fwrfT94TJW//n3lMUp/K1yoEXMhOmqWQAJYE
F47H0nYqjZLStMXbmtKULFS1DzufA+XSGTJXJynMoBeesu3Pm49U55wyxcwCtHAV
P7c/t+PqY4vgMh1cEtjfQ0e0PUJbpPTPRTGTiiFEYnGNJyBLfOb/KaNMfFXSP4NS
JcVW4Vawe0LE8wO3du5sehEXclmyVpZoI+T4VfLrXz7qEfrtx2oCn+iuDNiEnXDP
nYErV6CUFdftgk2pZ0yFSr8kD4D2+eMm8JAy8wRDLOgRhKc6h604ltjR6iiJpzs9
hFmh0ZOuShHdc1xgkz1WkVZe6B4HuaTVB0NFzcZ/eTm4R4H3X+S6n1eZW6vz1yfH
iYng2JZe2GLmT7TgZCowYUTxAl/uoHUlLD5wgE+yw81M+QH3uxRnxg+gDH69YX+S
Zog03Evy4XxgkKLMPvcPqPGsqznh19h4WaOY/m92mSO/ZMcCeEEw79amjLjToYYa
foPXpFyGpi2Ck+DltwyncJE3EIIK8HN8fyq/EmLmX9wh8D59DJr19FGf3GGrx+1w
4BLwtWNx287U13Pvt+Qr9sD1NldekSjGnm1GvsZJEjbHhkgVvAGZOlqUoe9k7/MC
66l6AF9TUexq+VHi+RG1Nj6/9LhML+TZWpcLaqsjaGcqreLYy2gjdhcpEGiq+99L
37xVsx5y3Iopnm8wCILaV396wrcwyRUnaZV8nZnmhLivbWfZeR+vdC1Ku/8Yx/dl
esIh7VKeImZnKK6Ok60HHsiozMVsfVOqqzNk0+QbjF8eMlrFlvHHIMH6xJ/4BUkr
24971PENNOI9AClbnFXkBlJ+YzfsCEppTla/C6BlMKLzAtYRodbni6+GsGyYLv/9
My68kpiJj9F0iPSuj33gwswVKYrusG0EnKaBlJJ8U7IZzzx2105rZ792NqzqWehg
Cc+pXI4l7pRiB7qIQnP7JGsI4UJFBpL1ViBqfbu3VxnN5oTai+z0QnyiM2wLVYMg
+/fJXhHMLu4wpSuybf8QbRToS3IfDwBRf7R9rp2aRXybN8mhj6Ag8XZo4ZmiVcJ8
2zdGYfGe1zHeYZa6yZ/a1zn1CgmMLkcJMQKimP+B9oc8rDF6A9Qki6ZKl3V6LyPB
K6mNv2w5ZmxYWDDy18Wjtz1wzWf5Q23lePdRsZTFJH2XAZAvFb+ghYTVFQM737A1
fO9l7pqeFUqEEEsu4i0bJlJcnHcwyGOc+8chGbIHwvbZGa2Juaac1yqK1cVGhBcZ
+qaXAyUfI0HS9GwFX5Uj4tI3Zs/ajKWc5mWbjrMzT9+3Ugk7t2sYWyiOdEvhpzna
8q3TfSWsyaeAzfd39DAixxA1OngDpRf7Fl1fPtYLUFerPNPpg9B1VzflEzPq8ukT
9G42PYQ/6DXujG2/i0FPgDk/omNGvLCIcydnz0Ig07nTV6Z+EFYIoFlhsJo0BEUo
BUYJ2Lh+aPiCU8hPxi04Rrau08aShKat91DLr+bmqqrNlZAwY13GrWWjHnbRWTVC
a61vQd8AxKGHtgnWpqbcc50j/FWRE1dg/H9snr5VwImBo0J3AiA6zV7WQIb/Iyw1
/gtuzNDG2J0J8rnydtJHaGjfDMeGWTzVL7tcJnuG9yG2f8ImVp+u2YktxoCKRR1H
PsVhAqGWMQxHUUW6qNLPNRXHV9JPQQZ4wXTJ5iXFU0kiw37lSzvjPdxrE04jljUx
qilX4/7t+pJoa4xZZbOmiOotTKJMptby0TyUVyN+vvKK6EdUSDTK4Mcrbi2fwJjZ
ck8rqre4or3U7YmQGKWtl9U9mrZYW747jWxxmpfc2ezUW9EQQNSfLUvGnZKDyMbY
gEVJeKdGDeJMFxE/xod+eamOSs6Gji2BpqHeHEtfA0fsT+172vPO245pw8O49JbX
A3XipKKteNkmOq5xCVjBkGxMfqvmVAQH6k6rQ+PhCjKwgDNXyjde+rSmqiGKXxi/
FH/GV8KoXZBnXtSaVhoJImpbMRVvSr8+VLXMnzkiwv6AYSA2gSP4V88gA+Zt2Nzv
Lo2aO4bkt3vnSXgokVuYXgVE7zfkjsYVvzxVsX4zGo+rKs9AJJFQj4y/N3DTft0A
7cALEQC5gSRD6ZRq5B3i8Aw6zX8nf41WcmK9F85uk+8BRYD9vaFdj1x7VTqf57ha
qrpq0uw1mTdJWxCaZIRQReMJYlygJT9cjStv/NkclndVr49LHIXQZGoG32sH3ljl
UJ+84UFoZaoDI9OuFvs8y+p6xU0prB52MvcWX9ix3MbJJ/iDvVHPYCXToz5Y9vnW
9UirEmJ1txCPSXKvXcYa96GKzSUrjMFjtXcASZRtPrjjYvLggQ5CWlCMtlMjNBBT
FCIku08GbyHXnknFj836su6TFPZP2/QD2QGWa5JWbui5Yzh8AMdOQXFOgYywap5R
GcrrIbKPvC3PHDErrfLS9lMGG+79Y7fc4jKvRKBHazKeQhSeHMEl1Yh2aXjRg4DP
jt8w3xxIhp73eIYy5ac686OY7XmrZ27SCcFFwVNj3rZ4XI0kyXFSTLl4Eslj/byn
nhM6XDjGqFMId1V4KYsseRf56zvIOSDL6yEwjHVf+wNWA7CxHd9oJEXR+bIRjJsv
q8y31Iau5BDwzNbbB4mVSi8qrDtlTUDQWl2ALsqKselub/wqrhTmEUS5Dy079YQp
FG8amH/OuZONgqd1XLFNpaYDgKEoO5uBDBVCtlcC9bpUFyoqt1f2cWkLhOuQCm8M
JkKWQOpQKTxJ33TrRT/G5tK/xQIsy0JPuw2ZUJBQOHrZfqbYYjuBjwuruJ7CeUj6
jFFtCK6Zr3t3GYP7N6Q+7qeqf5vYEz44cGdyPDMCmLO3ssMx/ujsY9DTPLfo5fRj
y1Nj8D0GxTZUR6Ru1M7ONT8OtG0Xx3HZoI975I/iCtcZPuIAOYUbdUNwCDtczgBo
M6gtyFn/tWgUY/4oW1Sm8SX4PmqPh8/JSUpt8gMDn2eDiJGibBwbL+oml0pBvTMQ
CsVWRa4lfThz43Sdjq/wFrBfmllipYdaSmAnYXJH3fxWk9wzMUmL8xUPbqhEEEdv
3vSIOOAEIbJyK+/XOu61PG4d9Q/1LfpRI0vdECk4WHWkSZYbMJP0mmOMc0mVK1C3
otITSnyS/t9c6aDGTo5YoB0bkHIZI7huMHRbVw/7sSdC75CLSoCF92DbyD7pVJcr
/JgHquvrSapB9mJMCc99vlQI2bHq4wSsszCa1KF91Nlmfylke4wSJCoRR1E16PV2
HNaocRDPQevxbSOsFl2B3uPEJQrB8WpntZ/4YZmomsni8mbF7V56mQOXKKGTSC2d
RG63hekM2Jof1byRtG08CccIxSj5kdXWhC1ltzQ4qPliELKy5KYreca5dsSPeu6a
P0ukxam1du2qfiOChQTdKe42R1niqUbhiBBfnEDlJASHgPJUpyY3Cq3s4wHPoukt
9g5aASow2NboSQh6C6HPTk+LRi00H80gZTzF7HqkKTXg9D9CCYzWPogxn2HbvKZY
ux4bnk2pKM0xi5vjYyhsTkoyr5qkQyHrQSWyWJax/yBAJhJYDPj1K7MpMVqhk0k6
IOqGnFwY1YSf53uaEBtSMvI+8aWf+70Byj13Yledo269DvWeAeeSvoHI6E7iy02e
HFsmLQ6hFDTR187Wqr3JbrYHtOrDLCntnu9K0RVdK4E7t0/VH/BVnXhmImuTCo2G
HD2RB/y0LiKMDcYxz3pkn9CbpGG0SR9iueQ/S2dlNHlqZhlLws0qkhHZvE1br2uY
hFBGOQySrFLhrym/kNLHTkwYBBSLiWOMOGif4gpvlffxA1iOQxWCyBibZ8GeuLV3
Nnytq6YImx4qS2h9VonJ19f6fPHhDHpYKt9WWUrob5T/W7inlaw9aGFauX1LT0Bp
DAfmGVZCFAFFc94dXqkcHQuhB8GjnRq0uut59myyzta2u68ImRGCRE4DsIYMrvLf
zjvqkTIJt8a4DMTFGVwrf0iUkpVfwrUC6+ZnFwk95I9vTBxueQmvu+wPRrDE68SL
/kfugUmTfCg1DRHOlTgBFz7VhYdXO6qAWgPQUXJ4aC5ccS1LoBJKILcGpW10BCKX
6AGcP1ajwvPGp9opFtMcJhAajfGA5j0b1BaEga4OsMZKZmZnKYafVqk55+4rXifi
2YkUnRQQXUicZMPe5y9d9pq64tH6kKcgYcT87AN9VAqluXOSk2tRIPPezr20HiEr
fPgyw4apR1umkthXt431G87zfyoYGq44Ws/T/qOJ8AG8y6bw/FObE7UbPjCmqnF8
TYUwGRwRwYuXfpJfmH2/ZyQ9Kdwymj10m+yQL57rYakdZAUjdIr4T/+0O3Zu76Pl
en/+3uhldfWoHudtPfpiPTdXtfRQK1PTEPpcI9oWk6enrQoZk8WmE3n/3z1C+ECg
H27SukmtiMxjJL5u3kruNyHZNl3VlF4CVjDJv6xaJ8li3gC9dj4OSM/wpPS4pfqh
igjCukYxeE8T/sdnX5xHCPFp4BIa5RtkYDbkIlPRdACJBGPiuOCV1mEdjJ/QySrA
Ay7D0SY2EJO02hXiyLvVbeUY9zuQwHE6kTpgsnDy/npMBSQMclMaAxDzR4yPv9Gf
irkcMogDBAIt1MTGSrcLe1l2vfYoDosWUSW9sV7AzprmQBkPh9ioSburu+sBJND3
aeTqdQ3nNZrSIt2COiv25tboiOnuWxb3GHK4xzEVvbuoc4pNn4FxsGz4q0sCWLoI
kwInUWAm8kWuDDY2Dn/aI/XN83Ni5tdFR2BkrPHdXX6D2NqZkZIkks3GDwSLZQ5E
beXzIprwQ0FXA8h83HaQJnrq7zLTqHXoGt3NLQVwYB7sBL/yKTlbvGbW6Ieh/CMV
oSobmzOE6t3RHCPTtY/EFfA/0oduCOgUucAENe5Yu3T3Y5jTn7/vVj9WhqvTKIQ2
QwLR7UKK/n1NeK35nYKbQhS0VEfqLO4MDmwsyzzu6Zsol+c3H5Zi+qqfe8nG9lfK
WYkeXKGvXx37wvhNk4LQ4SnmPhp0E0NI6TtzKGBT1kGZ+i4U6E/52MVHmJuUfN9I
2aYLIIRY1Id2U4zj7wHqw7L1d2tJ+wxVGHz5cp+4BZ/9VNjk8FrFWCx8TvbkdNgj
zMAn47NHfTPZmtIcEBtGDLZlvRInM2M1pz7MXNcZeXC7xkzgQpH5U2S61ikNaVCa
22VsK2wESC9h4bxHEM5antp4/3c+xFdSyirZt8mG0aRNIwmKKR531o1YP80d48UJ
4KmLEZ+9Kpu2N/wgKQXoUwlXi1bdUAYv3G2h2BS7is+Kx3+/g3ChxjjVQGCuPoVo
ceHY363lZq7SJJqUh2POLYpZVjI80ttBS9AbNd7RM761uv9+JQHVDKdySAu2RwpI
sVrqnsSE9bHWq2g8aNvmoJuVZjssN8rDl/vI1sc1v5JEWiFL8tvqnn5MnnD5DGkK
wQV7fc0EDT7k5Y57Q9ks/lZ2HqLqO+bhnv5n97R55Y3UAPRzXsK1tL64iqkLgSZv
O5HqlQ4Ddt7OqfeXn1Jr2l2CwRx9+AcYkYXWxiX7jnkRIzuuyGPy1g1SVyT6aWWV
0e/R+H5wDISsD9ecDT5Cqy3SLuscU0JjUHdT0Ie/pUKT48leJJ1nkHq8ACKfImGq
q+elzvgHEq2EW5j+Erbt0talhK7WVaY/xorDfELs8CNy5YkZ8HckvAp1c8i0wc5l
rhn+KupjSwaP3UPGzhrlZ1CRlKeHn5v721ZNmdeOVk8zPShCVb9up+bKzwBrRXRK
L57HEIucb+0P3axi9cQbbRqmPsGiZ3xKeN0ZYfdxoBYnxEV/YiZ41WXDcPnQTScg
mPlg9MCjQIyUXthd3qvzBjg84HbjXOx4ZCWfl14dm94h5fsHz1eUewQdFVmtQToh
DQjEzklD54KUh4ePSy2e7+NBm3uuAv2ILvJtp7UCzUg96MwVueYjqNcF5/6hzngy
45no8ftAgX0AYjct51jBJmIIcMMlHFDAzRagTGBLy5rV25n5k1Geinmxc9814Lj4
XMvzA+2Zkyi4j34HiOcTbqGJjAUvk2O0RKaa4cfhoVNrmz09ChDCeOavnx+Kzk2b
/tW5m/G7d3ZQm7RHharNrIukfBpx4Kqc7NvIKuIMla7BCtGdpkQYFIio8AIsOcYt
TGxHKHj4QI4JmBVDkBMoNXahK79mfh8B+iW4DB5Z08FKQ/OmGHDVP5AV861q0Drr
1FSvqaxvIm3PPJm4UwNCryoaZLlaWViusbgnLqA3N3fUmVg2hBdqcHSf6tCHl9yk
t9zh779/A9e6rOPho0dRs9bmRC0A7I2uhD0kQ9zWVf1llJOshVNrkIsRGvArqD2R
x+L2LItmGbc4U/ek0DBjftKZIl3D8soFk5+zBsOq78v+C8/84LhPxTdTz/3KSScz
CnjGKi0viqPH9oqsKufDVJ1+AG6iRJL2rnxs9ixxFlVWItKEnzhrMjvaj7C1MYY0
eqnd3CUQ6mkFgC0EDGcOcWQuN83ikudO+C1kSx2Uhwoyk7QA994YRehYTKO8RasN
N9CE0XEzFVn+N/MB7YTvDoiuelGl7CejXkESvIc+K0DUmONYgsHkRvv8CuL37LTq
qtuFWCo5AutbX9thU+Y3NnZc3qfDBTiH/6e268HOyNza1P46udISsV+ZDOzNJXuu
b14rvUJWX5ocH9wIxvg3FI3jNQjoFULj5kdWtcRXNtXz9XISy+VcWCu3g4xCCDLR
TbwTTWzpAkGY6OnlFDLBoE7c+kUZe+7UkqHglFjOswVfasghCo+AcDtPuYpH9JRv
gqqYOJxPY0vyPw1OLa8BBA6AuBoHMSeUDSf+nXewQtTAhXH3n3hEEVWYQ5pw/SA4
j9cmyF7UVRyONT4B2DzczcCV+Gw10s40T0hKt2oP9EnpYVSDX9SkpuP9n7qSE4XH
e72mFJsTwR4LiY7Rmgc0tVyUrEdMxNgNsALU+kwEok+Wnh+e6MHmtZDoaY14yBXJ
tbHkF4MuAXCv4rqAt/PBQwQ16tPmiN0N9D+bb4/JYoRSGkURpBcbU+DN3ulSKcro
z8JhhmSNcC7b+UWyrRf4DdN879T4HVkbwooHauuJKX3NJtjcSr83XhyN0/7r2VVW
TWpNorQrhfXti3kJRx7j7xH7z97eROkAjZuMFNR+KZxHFsqf6AY+5ucmkwRlicGw
ZOACkn1AR7jOj7GCRzAu3qkOFtrIftdIVo/rhP9imUUbQcDsW3JLOcaGJz/5sVlx
msVQbtkE5+LSyZdltQwyaIHmw+WYus0owbuEab3zWB80PVHftqwbrDjq+pPqrpGm
gYnG/WtnOg5OveW54Q8R6EEsYHXJ63wWACgQgPSqyCw42S4lJBspT9QfNaIA5jiP
GSaM/Sdpjro5py+HL5sI6oloN8tR1SVvqz5sAU3DEFeCr1vcuMIiyTEQbtF/K7jj
CZtAJG09zFJmiZ2X7L1SYVfm+yj9mkou4sQpouo+mWfpeotDqgOXKo848qmH9AXF
YVa3MK4m1p6s6erfckv8L5QMJigd3+OxnQGdMQYmVBGST73cBfkrmD3FRfrjx2Pv
kIMvQR7ITOBz2gSglo6TAZ246eO0+mY0JgLcMfAOc99N15E647y/qmz0+0GQ/0NO
5Ftgd3ZYjkvdv/sVRMviB2LblJoeQckTOUgK9dUQhvV8KU0VeB6lqpS0hqJKROCc
tePQZTj0hPYtmDQDdjYI3My688dKRMvIyRPOuqiFvbv9YhC+gQZ2b9vy5MzL+Eya
FZJaMZ+sHLMAB8U395oBxe0acjTknjiId/zQ556xdEbTwOL3srCBYnmaL7inAVjP
Ewr+BEZbF7vRGqqeygT7TagyCO07ko3tTDqobVBmnxYv5cKGRiMUHFRc0x9r3VNj
BCJtd8DetWOWqzy6bfrGPM7r2YVcmJIc9n/w+QF2EKHgoEqRcwNx8TI9KBzQxErh
bK1PixyNpd6ETq1TbUcUbb/2NkLcj0kh3SqWQpDP6s8eZ1nIij1ohrOeyrFn2vZL
upv/bE0mK+YIWx7HmUR4NCYDkeYzDWJ/TBSaTmeKTqGlaRFVy/bd+K8+PdBl6jdG
l6QVATWF0t8GKxkdd0dJuW8DzPi7AghW6oPouUBW5WPdQi50Ek+xzsp2hPIOhZPe
LUz45DfsP+CwPsWbt/dImPTwqIAH/8pp0Thxa1oLgOPg64Red5aocD/Xm4NP8asx
KHsJzP3OGAu5m+EkPh8rIw23NV31WY09SzZ+kPL5kB/tMk3e+FnBdX++bGR7rEm6
TQMDb3PQbE/Opf12212VdCp9vSOdm7vA/QFGdFN3w+NYOCbzH7T6ICPE1gp2B8vT
HYkXDa4C7Oc7AH8rLlD3vyJ+nkLecgSCyNUdScX1uZEVnMxNiBsxC35kJwF/Sx3g
1qFEzDeRwVqPTDxBqT0z/pqh0Ppkh98BJ0KVnon5Eu0c+99ZOReL5jM9nzUNzRPT
7LqNU44Wx8jrzKYOAA5ogny7cqgML3FVuNM/Azz/nohefa7n4QgtAjtuEi5TJw4p
Ae1zEn211qoCsz/AzLoeIWGU3UrAbh/MPjO7g14OA4jm5L8EnYAJhJ3zoKzitnHP
03I8KdFOvdlA/qa5phFOElVWkIhsKyXvF2ypskRO6UbWcMjkNQzIVgQ8UbY/jDrV
UM84uXWWdMx/Hvi72OX6T8y7WnrCBJNnz/PIXuLdQKwj4bvOwtGi/7JeDPPUeEuA
kOcfNG8gqivu2XZGhk4jMEbMdElaAiKa3LIGwzOUsYfPoysw0c8Xf04//7gT6fkM
fjuO0TRn4oCPqvBkpDob1Gcxgib4F+lkfTOP9oxHlBYoRtVjY25pCEpsLLbTwg7m
kfbTwQzcjLj1E+BISRqgYWWNyqY7QrqVdYA/2/wW5801XC4QQz1kSdDWeWubFCde
sjl5W1thGhjxMcR6Gbseycy+5SC4V1VreTs+vud/uQ0tYByE3ROpuBT5oizsYh4a
6RQ9fLWkg3aBHWjZKZ3XGwpLjBRnnGzszaCBnPPDTao2BHwwF0rVLUI+vxhnekOo
s+7pOZjP69YDU6CS+8Hd7FzyGezgXXDkpAb2+AvEcfZk+HBTPaIYj0Mixdwl9kEG
bJZadFwkAwP9HRryQlogzeeiy9NyWpsqS1x7+1ix0YgSlalHQVVafRNzdFnktqro
wPYuPqB6rXZ3j3g9wlQH3nQjaLk6l7nlE1ra/V9No8zOGhNKdv4HVa/y29T+CA44
EeSNG//aTWJV6EYe+cEHbiriOJNutqddU6FSzeQN4NOB4ljAtvPqUHlkSS672w7A
cVzSmZ/Cf4wKVux1Z7Ym+3FoKE13YQHiZid+nmaM5ATcgbArnNubUMohzvHixKbv
N/BYzqM9PSlpfdJbYG5Ip3CQE+r8SlcjeoxvcuYpaVXSuyQJ2AvzVpwoWXY8SNWE
ewlR0rveDtGJp7e72iJvJkp7m6FvXk9/cBs6GopYkLsL1Rx+zT21PXttke4MjrEa
Dn6HpYYDnpShlBUTbsF7wAUUBnxmcvPHANDR2wKP5340fY1C019fJpr/hEpnbra1
jCd638PNY8/s3U/uhzbqQyuT0T92F2EAmR0XexPgsOPSx/7EyjV7z6fpeifv+JxI
mXBv2CkYv6ohctn7c5oposwrghVtX4XRm2uIByKpPO52BzXyVnQ3GDWB4m2B+SdJ
fcPvI+2ipBrG5m/tPsb/BvvD8hHhf6vKwOsOKE7+0XJS0TSkQfifmMUtkKdbMDjb
1/Pu1AbsuVVnjWHqFTJJTJC3M+sleWCz/YvvwOB1l26lh9+XAisXTGiPBV2v/BK2
AdeCgYjUm5uCy6Ydm2dgTih+mKdbdU8ZE+cfeUjlsZe0EWjXN0WD0MmYdaF95fzQ
+Bl3Q0tqnFrgtkyCW1EjsxTghSiFRd6XtKNQPxC0kTfyUXLh+Y2Eeg4Rvxqdm50J
LbFzLLEsesEu+n/tqO5EAY6g7V+Ed25DVSJqpsZGyInxkMbYc+GVW7nsPdGehwH+
Ogisrg6o6OPmbJH26g/loca+dUik43MItKBZTWMwpuILjKI103YnLJZIC3dSTRpp
6B2BDoPANs7vib9uOy2dvIssGOYXgZgYBnMC8kbbCStHn4dtZif7ZJZ5bP4E/bb7
ShfBfkxlOqLZ/Lo592MOS9ztV1BKE5syBWJEpx0A8vfYryWB5i+oOOcZxpqrbYdb
0AgSiPM1LZ76KHeWaG222bt+u48X3BsJhJQHXxgYUwkfLnhmATfU59htssvrjbDw
/ypXFxzbbwvv2L5We4lO+41e8/Dg7hUQFOxGt6RN4z14p7nA0Y6s1bXfp5QQi5sT
Es/LxIpkJDPUQ8DT9pmwYbbdhjDNix/SD7N8U8g6T3YkwubNulPmyoD+MhWRaq10
0UBVupCtj9YQ4dAcRHziLwIsJrq1aVxAHJxegfTWKG3erQQYJgb14AtmYvFVNlTW
1WjwLybHmqxzhx3FzkJhKujED2sE3xnZ2NPwGiaEEgo4VvA0+fJyQscGAH1R58cL
md+XpbHFNqQb5YpN53iqE0pcxynvWxS1zQz0hxV3c2ENjmKqgLkU8POTnezBnYDh
cAMC58caTYAua9xO6sX/ZzfISIFvRSCvj4RwnpJBiNnm0PJj5gIa7YZBjQ5J3ecR
XW9xVBKXNAdj1AoNxbTZJPdJlKMQYW2v9pqeX6OAQrjguNnNhtk1SyKsOyL40P50
Dfwwl30Rt3EIkcLSUDj+aEpLJoPIRAACWolqc3XXmzkp3ip0dkCb65jZUBQlSr7Q
kHmcZO/kEzgw4KOHbY1IGLMO3gR8uA1+61F+RSP8/DUAq9yqzao0kIqoE3yna4nx
v8GCGTXDOPBCrL52hkQt0UJAH/fBEDjJ2bWnLFch2jfpevajT9Z53lRM6yRml6GM
thLCV4aUjFH2uxfIkESGVKou+Y/uv/mG5Rx0cR9gzON1YIlZa5XgmLdQHGeKe8MS
zPnhUNKKEuoQRj2ZhMZkO4U1SYwCBXISodQU83e52skgwGpsGxXkd31nmZcxZwTU
6v9hvXzhpngtfU0KcQMiULUmWNJgT9MbEvhGYJqj+T+M1ZiJVdlnv90JBcKjXx4b
Z86r6lPKo4rnJFMLJdcyEaLwDQe3I/2h/++gW1kwY7JMQaeC/+PDuCh/R36g24ck
6/sEZpDV8gKDYhkGl6BtAZIcayGRvq6uJfggMYbhlroBBGDkCSx07PMM6wPwhYiG
zedtRQjLj6sOMSpa6MRcg1RC1TXVyZUHjy/27gs3FPzTiRNcQRBTF6UHXBIm5dvh
4b6Qa3IhuPq1omspreJSW1ZAjXjBMXG+SeNW6L+FEpSqN47IfAb9bk5Ir3p6XrDd
KE8AN//SaNm150otDn8xx14d+ayi7r9CIwLAks9kRVZbLtkk09AlK6yEMXq9Y50m
fjzrBSOE9VEZyCHPZc67oBIBzebB3Mugo6wqpg4qGUDIl57rI0jdQ1AMeYhlnN7T
YQilvFxJvq1eRIabgIxBis5Ar7W5wVz/zl5idULcN75Bbyjs/WSeA/EofU1X/fE/
m63ZF/zDZA4C7yEZFUVmaG+KYEtC7sFyeQuToP6Uw1UuLHgeTCDysuftj+gyCNqc
56ec+cgd9T/EArO2W0GKYSAly2PfC+lyvXh2YCx7iz6/PgKodldf4zeZZ5i7h7fD
7sekLQp6QS1fKcAhCsR5YVZ3DVH77v0TgEnjdkmve5pcc1y7L+a55Q6LaR5FcfZF
8Hb8OkfuyHXDvxJ26GmLAn5U8Fnixt2sv7SaJ9cMsMrbzrekk+62BCpChfb588os
Rn6eHpBRiU4rfNgJXv9uwAzU0uiFaWUa/i8tIkSIl/bWJJ9dNGucdcnsjes+FwUs
NJcOPP8O6XAkb67Gj8VFXxh1UN8iP5jLuES+V3QvyiJ669NaFLAmmUJIi8ta4mhA
CEreCnIiai9Za1W8421k0feobenicndK+toMDR8MRp3++1m+n+tuUcjccrX8ccnV
QW2ff5AHP029ovAyUJwVJBfHqaJMBJzFiYqmv7Vvc3SYBzfUnNgzHX9CA1MTWRem
nCkKKDjcz0sayUOob/x4/UQgD03FYbd8o7w1ZNFCsiQnWEgFrTQMTeSFbIh+R/SE
I8UJ0dUX4X8LgfVuzjXxWLQhvSHBp0JpEf/nNnzHMMCkqjmnnzWZCFPMJgi6kdsW
F+yQqn0hYSjpCFLU/zlhFfIq4C2Qn6Ztt5GCDTTurAFH/AgmboTHo7VRlmHSZIEZ
XnMUiBiiVk7FdWCJyRgQaxAj/kXroXQNYFnbs2NInUhZBGF8gnFLKyoMpfM628jR
Ag48viH5bN8pDqphVZUDCLTrB2FLkgI4f9wr2J7Zt6W/i5mBy/8FUlucAazzuVv+
rndX73jts97+uc/DXu8eRflrSELF3Zt0BRImVIBeQTo74uhJUXD8NmUGuouguD87
bEcVIN/J/+gewrvgYqiIQOTBRTcpihKYhITFKrCwwgufh54ZCpAuUq63d+sCck0B
LH5geUExGqhdMOKuvkIillbn8/z+MOCcx663CkS3/HwrsZnVZZegby2nL6/blmcT
ea65sOO1KsR0ZpFSNTlWIsUiQIR/s47C4xEylPe6gwm1TKquCj+rWr+/Tf1oZM/4
vB7FUGZNlk1trBCwCY2yHJyctCjguoXzvDZ48Ez5Ycj7kbRCeqKWMz6SI+8TDGBK
bTi5YW5xPPIPmMRorSEu6pikMKbCxPId5NEWaP3X45Md1uMn5rBBmM7jAsdHv7og
habzKLNlCuVg/e3FcjxwXbEbd+cECJAkh66QKsgUqWOC5O6EiDmutZ7WoMRFVgeF
/gwo7KYeg3YTWC1qzDTwjZwWXErQSOD8tFYDVDwHcIF1g3IIU+CB1tGuq++FDf+t
8k6bxJEWsYCE3S6XXIMQdbcejx0nMS1jPROPVTLwQkCfBtW/aE83fYnl1NA9JRIn
hZ2C459ntHKDyOpdapuqDy27zXJlf/rvcVex+Bq5MT/Nb/bpihCSkeA6Z11KIJZ9
pVUymeeo4cJ9qUIDiXpzdYiOMBRy6xoCdsgjmqNaSDLaQDi08QS6N2vITLDrRcRS
oaQTxcuYCLS4IWNDpos1KyArg3iiA7oBqc4VBepCDl/ck3qT/jd5MW54aOYHBFie
SuiSxDd7bXPXq0zYfIKZmlF7HXEveE6HSQB+sV7xkMIpVti3xMHSpUNW+Rzp/K2e
gb4W9doZkICtpm0OoIZ95Qq5wgPzHw1XmAbFTOBXIGJn4Ivi+TjqYLEFbzWFTWw0
7ckxuj9WqneCrEEfJeSvqQYCCcVsftQjgXdXNBvcfEXgzE6Akjpdj22DQnaGmvjr
n3Ds09uMhEZjBeG9l/PdiuxMdqlgrVP6/nPNVGAeCV92eR3Qchrt+4egcD68cS6C
h0CcPxtYXT8wR0AF9TxvTUr1o9IbcLivDgobkU2smsctnwBSulAUGTf7Bt5hX/go
7fTIVRMv5bK5eimCyKgTr7dAMri0um7k/hYELmBLt+sZOj02lDlAX1C+OGOa94DC
buNmMR+kfvH3jeZ2oMqHrmKmm970Rt4EHekSs9q2yfSzCwjcBnABccs9/x7tLqFb
xzDeNTdjvNKfcTqTYdIKIRyChi9xNUh0+A5sOxDyFe89juNB7mo4yyUVLscUbom9
QMWRQsHut9SgLYKs3zYXKzHPUTc5/lxen2lZvuBoRIeLkg0He4Tfe+dFn2ndQCEa
T/e62rQ8raBQaA5Xxgc8C/9bA/MJozBclVJEpFmRzfXC8x7PHIhy6pn8Js8R6ZgV
7AoszrOkNPDVm9bQT1O6vL715Y1jwuMQyP6JFIP2P+NrrJkigL5/HqqpuSWo9Mte
RAEtvLwed99FsNosy/uiGXVMWLN3eidRWydE4U0D5scDZfZY4JacwkPn4zrAtPd0
edfUNJKTE5LvwM3yXN7+WMLbXaFrLTxSyJAa6pR16zeL/zAI2l7Y2b0h1Lao4VtG
s/+Ki8jczGb8EfxuZmmo4vmHIWw/MQabx8Sjg6VpeMBEET/sQnLgvI8moS0L5taj
0UNdZKsu5yLti+ZXSaIqpErbpn/R/3Dc7upYsykTG32VooD0n05WgAtW28uzXCXa
tj3KEQVrmpg2FdBTpYC7gCISm2HM3qo6eEcxS6Rh8hxozTHmnP817OE8JXWe6wQL
AzRhjD3ETeKTDB/GTymxBtzMtydgFFATGL9Fwkz/peooqAA27IsYmtzjXR/DHNec
ekgOfIDBpbnYvTnbWMRHGw6pIu2NZ7ZGCbli/nGAfiZ3OaGeJJ3xCXZC423HGd8o
ePF6gJ/nJiO3Sdzv0t4OmrUVY5+OE5NOWEYaQa0a+fI443nXzR+Pqu1wynJbZqV7
2G9HLApXTUujpGxHjE/oGFxGqOZW1zuQJKjXUw0pdikBe7FQRClQem+XyxKzx0N8
WjhMwClQ50xcatdIfu9OGF8bdplnk4q4Oz1CQLCzgvBW17vHIfAp3ayyifm62YgE
BTR3c7L0wd7HvXeVIEfG8xty9NXfofbIJhqHO+mRQnb98gPaVUg0/Y5iDNOgibxK
J8hy55kq0JSvylJbxy8vkg2cfpJ278jxuKVv4wyzpuvS7VkH5eFBuiS3dArMc1/k
9WEtjkmm37njeT2H9K1VFP2wFtez1EGyBrdZCNxEVn3tdAya/uHw2GBVzy7OJ+o7
Elv4khzpYXLHEBLCtcHRpHbdObzdLMhNtfDMnrnC8s0LJSGCJDQuiTPp3SO/Qi9T
V0yj1Y5qAq1A5YSL09CtmGfbHCFkcxfkY94RcIEgAKj3+11Y1Fjv62iPdUReow/w
w4YXXEgUxVlwI3oFHPYLuU5OWzG0er0dR9T5wb8HHyWT9UnGeuM0rpyi2tWZpyq3
4wL0OcgMwuvrAysZelc7KqkvohzikAkn1qETbH6ra5rH9/C+9WUSMlGdN5JljULp
BU4awrT35lFXTR1y/s1/mHbLboG2km4Az4171PC4Y6DRJn2hSn9n+FipXbstmO0V
DdgCu0topPDTWki/b3QCgZm20IuUdtC6PJXpFLOQDkfWy1GX+bQJ4EM7Yn2B/UmL
7+GfI3RpaF4A/tBhlSHwXS8T8wDvAP7qjnCgMZtXgXEBZudZM/tU/AnUL59fCwR/
Nwsb4uM8khaYmNqojKqRpcQiIp8xHr16tM3GXZtRiUk1ndiRxAFPEPOKL0sVhUNo
9mL2Gu+oDmt1pANwWIFZlLS0i27HQdZOcdFUUhloazqccmS6rvte97ZXSP1gOSqD
w7SG1/FeDD1Ua0QmLszYvtBHUNgTD8Z6Z6SMT6zYmX5b4hX8OCaUmALfOZFcqOh7
LWTiQujH5NzUbaA2xnnNzfuOd3YdkqPTNu2vHqbr5znuOs9QDIumCRLiYAiHvmMm
Gyl8sJZTl/nSMdwXYtEDvAytxUWNGfWtxqqnv5nsjUaMEvNEV5TdILK4zr+7nign
OnwuiY9SSPaL+B3mpwqCdW1KxWPiVkHTj2iSsm0YnsyxFnEr0BYX9jpACD+5t+ct
V1a3WQV6qo0wlbntYv8Oum6aX0xPvCRqXRtXZmSgSS/DyNYBXtNJBR0QZG/aAyd2
fp+RHQQsvnwV1tFnN9gjznWfm599GS01KFsh3KITn53ifZ1ns+uN9Czf1Qx60jBB
3VBGFSA1hL1wsZI8rWnMvh5MfOXOzSH0tDePsfxJcyeBks6ROYVrM8NO5wBV75mz
IF7lzE0QH84wZdlgpmtJuQQtrfeag9LRrzWT744yRVGkGXr6+u782BUB8veaFesu
P52EXkVnzAvU2A1quD8eKQJvP7yPzgdAKRixBGzEvTJPq4qVYCnTmmunDpbS0WyH
JJfSDVQk74FhcnhWyRvScl+IqbRGWDdXZhoSxmUAur3Z/BRbCk96vug41RGRZ3Az
e9huj9lPVyEZ9/6iwsJAYoHfP0CPaEeB3VOV0C3KE9IdO0/ARLIxi4pg1Lh7C3Ir
ZfQFCQAcNd4gBTU+c89g2U8f3xTHPBjOuOkciOTJuh2FOukr+tp/xVObQOcvcys1
6mAZsPvo++FRvs53A5OKbR9ayufww1GnOf9laMV1rCdfTxgMp/eCO3UXmxdqAJNu
X+uR9mJ10Z2/H1Oz02j6CmJwC0W460EEhwaLfpvW/Hoxlc0VlSQUQfYh4VJ6dfn8
YUeUowpRVN5mIlrM72BOqeV7NQ0KKG1YVLasyorN6RroJNUgWT8zXdz0rEI6JdiM
WjaZowbKTVeggqRqoWLUTWvilHlJKQh6Go5SMP3yCpkkcxsmw26mpxSQmVUUXvop
B/SLE4IqjlM6piKcCc0qybG7tEEP/xni3HTtpEoANKPE/6z+ATF9B4QJ7CmthSEF
sMluNnd+ldAo/i+aIvMVcb5+XTsudwo/JhJTzFZdUrHYcZKtXLSCBZdoT0+S6noh
Zl98vPNxpfmbgG4U4sl+1vwbSt04mK2yIwqkjE+oT2CRkPrPp3tkpMzentphe88Q
Ysl5puO09+nf9lT8RgoF5bVXmPP9K4c5AlcxWQavgFH6+s6VOzAJu941QJ8oOWoF
VAtLM5bFE9LEQkAxSIxKCrxaxkYSXcGbNVgcspCSSxmoLHwlrysDVLS8d4MPagFa
t6O7dS7TZK3xHaB1VIfkw76GfHfSB5tu3lnMqKTBwkWKjuxaL9OEjh9aprdd3CNt
Bxiuash7L1hfIU7zb7URYzmKtZcFmEPQPcWUrYXO+PfL1yoU3NCURQupoO2VfEVj
CjeL/UPlSg8X+mINCYBuonaTKCJ9qXXg06Yd78Xem64kyP+a7abrApivIVlLUq43
B/Bytpm12PjJIiYEHrzodUgsU1LMAzaiEXzV4wBuFosEfGP5Y5FEvWprT6jYgBX3
BiiAs1nCYRJ0l+WtHdWVNULPElJC8G5dVMFnTTNGAIyvJyki7sTnCYPqcr6t7uPU
x+Yzh18ZVGi7WEaQ4ET1G80GG0AHhRCh5CN3YYajLts1WvSA3Xp99vAUiD2+jmXg
KH1UC+d9cr7l5iw9A3FdD0D87bLZyN8TN7va55GjWZDgshivXcWE2wLBSxSVq4j8
8eHfM83AJ+Zl44iIQkMCIXolbK60siYppJKhMUfEuuMd2/eYQEWmAAUTXRF7KxMh
QVp4IvMRiw/D/gQev9ldepw3wJPPcKnK7mkBKPTf8ZP5DzNLMv6G20j5r+9HHovP
i5TcJ3nFUJMXrI0po0HVh7h3oyFaF0pbhmHN6QY0x915J/uAKQDNItlkf6xUpUKN
mOCankKQswyLV0fy36eddTDYVNogZF+M/Ls0S98L5zGyHu8KZWkOWHPL3lJU0GF6
yygJdyOJpiVVFYBEIZK+hlwbhkSZ+6rX3dJ9nTsSulmojiZIF3mU+1BKRfl4K6qy
GmxXKvWuRH1o1gtKEityzETvgYjRt3v0HhLeJQFtiQkCfaWRkABbDmb13g6ifGLQ
Ujh3u5qmjiEwEDrpt+ARsqs3jxDJGV/+65/mZ1xNgE1zYNZrGk545G271VvVHxbH
mtcPEzWA1m1gYLGc+akdvP74m2BeDx7RvVI0SG/DkKs+fd78kzBAwOwBXsYaBIWN
4Uvkz6CPFtuWOJUD8aaiIqOfFEiJALvWNYRy1JWSdGPGgeJ8Vmk75tQsjKoABmqd
6uCaTSl8+LG0bIu7gcExq0JcivBt6OGadm29W9OQqV5APQcG8ON8pLuOvFr3qwgk
ov+hSNBgm3GcXkrO8xvkoTLi2mm70lMH31i1uCCpEn9ceW5T7edellZrqMoKRiLa
BMJ2cztCxp11WGW9JuYUJnydCpn5nwBZk9JhsrOFrRToHLTDpjhfgs82t5SJY+qI
U+a+Dcakq75OYJEcsUrF+HgdAzzTYIj9abdsSPm84ZYdJibtBtb0AvZvxaRLsdl0
qhaRAOlKt3lDpNdDz6wJlbFrUuNnomqZH/SKMJr+CB01A31GK8gzcQGHwPHxnlE2
Py/Hfo4M9TjKHA5TZqj7fyZiKJzkY6KSdNJWSoTadrfapjF9XpXhnPrvoHutzRJh
XpNuDpj0RSsjbh+c1HJ9ANH/utvRkfNf6X83WZoyLSYZmgfwoB8/HYfjYqoQ8qYn
9wwj/LWocok2AucAKcxQRIbNdN3AF4vXN8d0cNHOuJviOeHFUt8AfCitopCwUyGv
/Ltc0W4ztNFfJPiYNAbhJHI+EGMCwSkF8Dy47Wuzhi/G1pnfOEWc5NtEHeASdRpB
gK9HcBr96gsIBx6xvY3GK0EAtpEEuVwPsl09KmMJS8iRGT8h0wydCpkFN3C/OFB3
dM7ntURDnwuU/6CXDqa98D4Z0O8qrHhLd5I0yizgpzjG0Or8wTwmQVIUd6Q0M4rg
E151IMV+hIO/Okq1yA1LvVPRVEeS+5fYMTUHPQVzlifzg+6grFpkv1uTMtJAFlSI
AzpCQxtXEiVBeTvxg7f7HcLm3ZpAvID0wtPEbaF6Bv9tKphMVLy9M/2qwErXTU6K
g/rt1lHn0vidgGWrIfraQEC0N7s0PM44/6QsSSs9A3iHIGMw80bqZ1jBF5jRtfof
YySvDOpTGRfxVIUEHMixxNkVWy7KGIJBdRL0rSSolRNDGu1QlfrdFUNV/2v9CBHY
gU0zVpKOBMY7Gt31BbrDl3yJNMwH9kazsXcIO8k/3h5IyA7mxqULtDjnKP3jkHK+
jfm9Ma+Pz6sZ5mEmT7WNzsrz1OqJyt2rGA4sxTJeOeZ6B4oHofFlD1GxXGwegdb1
o0/gdf7GXo4W5EM/D6RREfmJB1ItTR1jI15bXQhKt+SSzXh+ObDTFVXbbkO0Lvow
3jO7mV+snCmKaq6yzSoXJy3SR9+hWL9TGGohrhfnRbWMYmVq0Ce+fTla8Ml/7Nry
wlBA0qJ04nsUiZC7ycMO1F2zRKg17vgKxIK9Zn7m1j/2VBSl03+Mx8oOScImmB+K
Ymk51Zm6d/cCZfGOq+Ich1RTrE7Xazc85k3OlZP11TP6Ktdnh64N9Xs7YZRzjZcS
qxuUH0adQyUB+QbqNjZm/Exzjg3IdbVHOuMyLMlqMJ3fP6kdRMcH5++Ce9lP2jF2
iVoGh33ZsO0eKMH3+2+vEOQjDG3Z+ISPi09lYjgmukSSfrH/D4LHi0OA6jm/IaVL
4u5KqgcJZynjJjLAAwmzKUM6xrSCsH0WVG5OGunIkSu9E4rsYC3JSURkuVHg2fxo
+5XF0Mq35/xoSmRL0fA6SRf1G2LNZsaU2rs+ecpQ1CQ1DzSwOy6/NnrQdSteOlTE
7iiBY2QJXwNPYetRjakCF3dXMUpETqTClAnoAJBpg3p2fFPeMoXNYpWVqlMCopGG
A/xse9Ov3Nr+IvHkXgzF1r13S4eVL5v8KrJ/QCQl3h1DRNVOQ8PbR4o5Ew8NMabQ
7uysOtygfOEMv/dW9Js6wuya6y0Y8LezirQ9bnJ6NsvEeZIM8+CfFEwHakVW+e6E
CVTo4JX0fmJAySu2OVJypRMcS6GNGNh2mx92Ut4rVTOBvUS74ZDTg/tWOu14yR/I
EZHHuplPX8Mlj5GlpRhSZ3IY6gMfpP87P8Y2pI57s7V9Z2rtXJhDAMNEHxZs1FoC
d8rfV8AphGe9zZAN+SKh4VulhhBlqtXndXCW8wwOxQvUnCm8In4D0SKe2LjNClXe
69at707YH6RElErTmxPeJy8nbcheKRcXagW6cwfV+MBS4BBkw0fUdu+WRM4GoENL
adBUyHS8TXIRvO/mgHZXQMhKIpdcZSGW8MkKApYZwYkXGSHzgd7vSla5ELS7GHIW
id33zTWBLMisREjvPlatvjvCpRcHRDTwUABmjNtA+HLYEgEHggx0i+t/92rrrnAe
dWHAif8mPpg4CQuzjkX15UwJyBkxHA2CBTnygIALClpOYZFxLGdpeXvQXbrUsLHS
tdN5zR6FiJLa9e1Y6jse029xb15jGRhj9cLlXo0pjb9sWreGJQJfow5Nxa5qD9w7
P1Ya8iPQi/Br+me44LtlmzaB5v5Pqd0kK12nRwLnLRXncD+Q4zuF188DvnHdi0Za
3blVDnYCzIdYQfXqvtYwt4BYguPrjckU8geKIypM5OYkxeLQLq656NSOuG8GwJ5/
cU0NRhm1MC/8NhBSG03n5tv83NqDiicJ4+TJ0nsHC/tMPh4eaEwMi9RXGAwxETiN
Eeno8yxDT7CJ0d3zzXAMxxWzqyDEK1Sm0YMIxiuv63u3KcZMQli66D0+FH2pgZ+P
+8hGhb10kdJ+36k/9bHa92ucK5tReXRIgVWY1/4vi4/+x8mKo1L3g5zDUCV4ZXVd
Ec10frW2iLPa9lsGxOY0UlxODm/Nje1O5epDdpYAgQgS4nAO/WkK42zWdVY5LJWj
AQ5SAWKABfavnGDgcJjd1Ek2QOvYm0fNchUOatTMRJXcCkhGKYuyFpfj05/MATg1
VicG/6Z/2270Qq5uLDfLUVOQcjPp+9M/dTlj8EbnLLle4Ik/TpIlqBEMmYRY7odc
qIQ/leXyS/02nJLfOG5ug33C33QT1CwAek1ZP1/6SGxWotiHJV+CbvHRqlQfoJ4x
ZuEyS/zb0HcHSc+1CDMwvB0ukjwh2/MzG3RSCI6X4xybETylU8oCsTgiEtmQMyBY
OPHcbNBhBOlTwYWvSCmEEBuxSehXzh79Bk8z6G0eWVePaMN2hPzAN+vIRm5moYGo
0hGUbUVX+5Tz0EMrQQs2aIkMNYZKlYg5GnD1uRsIiW5X7DqgFM3FL90x/mmG2S0Y
Zv4b8oVxSGQUfGdHozgwCQ1/nt5JOXvEF2wNr5ZG2l/fjHUEbD5nto4+pYCCwnoV
Ly67CTv08oCRMRyO/gIj9zLVXKIjrbQGhHL8VOU/dhwQ0uFBBwPQga4yLzeOjqEA
XTtycb4stv3bW1la6qsAiZGaJ575lAnTiQavKdTgRYtLAZ0Tv5cWeiMl1AUwxmtB
lufO+kDWtYXoO9hcOPmH3aS1I2xf9m46a7BLmb3khkMlGNZKFe4eFvyhTpPtBGtr
Y4FxuYVZp/PfzYpbOSaxGk+SwvziTuY7Sp0H1YIS33x6tQWLrIRK5+eHFu9U4KGL
A+KDhkNeklLUzHMUovHRrSY2JF1i+fi6uUIVA5NM0veKuMFmBVZSlYVBDAiPfDhu
qwdyGCClBfRdw4/Bf95wHjCb4tqv4znDFLP/tJvqgV9jRRK2fGd7rGXpjqkQInhq
WuJ5ji4RWBVpzmScXV0PKioE6tte6Q/2WjepYCM70UPxGrmNrpSgPpsbkqf/NI+G
rxXbxB5lbGWHdJVUS4xsX+vi37m9l9w5SNYKgKSAMgK/t5qEBw+lxiqMVEdBdv5j
wbPqr0IO1/Ohm2TKFtnfXpV4cJjWoXbkcjEb3UivybzhvNnkJ4sezqXi/S1VE+eb
V/Z/cuD3z3tEMiUiQBErawRhti93DRKo6ox1q8d+NC7S+oyzS2+vwX4Uzi5AoWTJ
K+OyrU0VHvz/XGZgRU55aJ0cKIqppwFfHd4SWrw8C42pexsNogAcmV369jW9NRIK
25nqqzThqErB5FP+206lvQ6qDImjfZqAwRVTa0R7whQxkY2UQxPBcaD2DPRgrD1o
aLMKOoqjY69jRwaXh47/9gayphRPch2VXx+lWXuhi6WZMIQUXmEoOjJ/bGRAx0Zk
kSoXqGk5JppqURcomagQYFKpH+YKSR+IIzTDhHW6xe1Y5d185cIlmflvqodnYx4j
caYB169MePF4wExbmo2fbQzjropy3ONw212cJ/OhJ54ZEIHUgtBf35YvIMrcdDpi
3Hh+7NhM17qjRbF5nki7TUc67dYsbe8zIWpjz/2e4+CltNJIxWv+8ulODKkfI443
0N/KzIS970cCvmaDfUDqWIBp4EZ1IT2YBOMujq9xOVDSw857EkfhOTlVDF/Guuks
GQsX/gT0gLeQ4njcZSUAczfMSmLafRyC5quevbmpyEIfEHmUeqQnMcH0QoLLZ2j2
jgFWAbQRyRKttASseQY/SXczl4ZScgFhJZ4xqG2BvQRQBUbJU7p5yDBBpEm/N889
qqjsHLyxTdOZRHrpe9vbRZoNnvKzpwpMYkVdozGeuuVAgun88zLoL/RjEvzwffWt
zALv2SjQe6fILPqHOuxXO4YaoGp4YdQrLESSaWR6QBdc9JBxFBTIn2ypOW+f1uul
HSyRTPyt5yFp/f9nrFCRd1bUlwzBmFZt1/qdY0hGiHF3VkxtSOZdV87x80tTy9tU
55SIjfeL18d3Af5seXpieuPmACWp3rl0+xn1wS9YRYMubt8NY06F1GgLH6OT1h9t
Tj4h4MKKMwC62WeC27zSwyOwkzMUwRr2Nm4pKOY5uxloigUFztlAYSjtbTLsxn7D
HppfSNZPaoAnPDYaB32T2IAs3IHq65/SAbb0DurhBIZp+lC7vd0KhXxrtLAsuPqE
DFfT80taMoAc+icasVelaCtZj4jgU/2VGnUo/yz6uRiKa/9ut5tNYY9QpiGOGgQl
26WCZINZ7Zz43LwgtnamnaXMGslGqeKhjLm3/MkZBfS4bjh63qNYd5QxGNUBQkev
V/3Q6qhQ31roxihKwF9JhRqyrbeHe0vYjhpfn3l1nvjY2vVHJGVQpy6Jh4i7bbjK
MfbPRon/Hw8WUncKNvR0EVZ9f7LufoFQl34MXOThqaferIfAQd0wio1kJg7OPpy6
ydMZCI+cUt8bnD1Ifg63WzeC+QVUoE6VUUFRYs9R2J/m3YLtvDs0VeBUOyBuBmna
d6Fu9OekaEMHbQF1ktdx2fjyCllFvQbhzG50kFCIAuf72rsYkHRi/l1Tc9tldYBM
AJWEzEi2qsBWNfHdsJWJZcVOkPoIbbhM1kCWayOjnvrGCeMScD6rFB/8o3yCy7Fl
A0mfjktLtsYJ9lXV3d8YYWxEyBBKMtBebd0R2MJwQT4S6ZaiF0yFwl/ANnsQkaej
idIspLgvYJeE76IkrBDaIkBorCCp2/LwFgFT00jEXP0rW0c6DUwWu+xAmyiNWpDw
PbDMBEOryiiI+AZ+Fbeo0UIaXq5eaiaRshDlG/SeLH4A15Nx0Kf26cQ8zAhWWMd3
Jdcwu/iZkODt13sYezFAHDQKvS3p4UkypKGSrzcXcnpqcYu2IVbnZRD2AIqBpM1x
DhwZLGEF6SbjxWt3nNCNHC6ZVjpQPcjTMZjrjJp3glxgaadfj62CooB8iDkJhAz1
mrlRHhHjgmTSIs5w8yUDZExhDgrYMwt4tCY7QRSGG4vovnZ8HWlznAxUsojLxhGS
1PCW4jOf6kUY4EDUWg5JtSSUfiwCIDp2gdi5YCuDo04uOuFYEOv4CeJlI9QKdBGV
MTK2le0YXetQAKYHh07qP388XYYE4ttY7V4HpRY54gq/J10kvJcrOzwuABWELhVC
XstVR4fpIs2UztMqEwn8UuorBRMCe03aKTZylZcZwKcXFy6tBWT1Vfxv3sKWFzrW
gLfm2w3WbHKgsdrmApu14hVyV466lnY4DOmpF2DwEklXm0sOMPm+o0ifULWvxS9P
09kMAy1ymxVdrXoAkoYUflhM6+uUAkIDvi4TtxV2arAEAsTXXRNucp4xCsmM5U0i
+yI8mgBqs68WATBts9MP751uBoov7rNR1/HGgQ/UvlnNGr0y7PxXjoE5lUqjdFUJ
Pg1e2sZ4tvvs+qFVnPzHDDPNO0iisseztlebnjs3xz81rCn92tWYRo9TsijoaOGW
utfnTog9eQClxfcMMsLj1q9HbVxF65uG6Cc8u/4lkMKuWB/qMveIXBvZQvwKhBOY
FzpL3c7zhQ3HBdneeqfOVo+SvXBomTMf+H1hbaWUhj4dDZT/l4EQnP8R58xWMTWk
S/w6yMz9/SRy4xDGdvqD0zpVvfu+XFB1CJabazEAZ8kfKX1mIKAk74OaewCIl0o4
6kcI7boLUgcghJMjreLCp3DknOnWKUphaAAhyeatbrVqg5gy/3ENTBSBXD8OheD3
sA+VUW6KXUcU6j63GBn+g/8bqyd1juk9qZIz7WYZHF7ZVGfB2LiBfiVaE8h4l7Ym
efsFBPoHWpavHaJrYWCRu5NUxH93FgrahF60ow2WwQwUTYlqCuV1814QlIh/tZqA
FwcpcV+hCgNTWS0mrcGMQOQd+/gn/iac7fC8b3dw4KLiAjoEdIEb8TVEAoXU4fRW
nLiL9NGt91t1+wia/h+CaY/gwrvNpTBZiog/iXB/DCf5Nf2A34iWo+CZUEMiyJ9E
ISBhAvXUzXhSG8n+imcefVgTELKNfwTSmY31oS+X5VuVt3HIJdEk9cxbEU459Kvs
mn/Kfwgw9MxjoTtjl+qwxDHSQl4e4D/ibQir/7mv25BBPKZOA7se2yIgsbFtHINI
QsSvodGui6ObuXUTc7UJ35L6z4cwBIy7ndO5Pzj75EtoTW35QZvxtzrI7UsUJ5qv
czRuxfyfZyHO4fW8nSHehi5w20BI6rK1YhWeaH5hVQ4RY1d2tOvEf8dO/XS5cVm6
J3pKi/dZDOnniPcBCIiomKDxZsFJbKHL081iQRbRTn99WRMokHL/29wntrSuAVON
1OtPyEKwfAP+dK5yYDStHuQ/UI8KfZv8PZeCOzV2B+imQHPzHlIOM76tlgdUHgY2
T6Ymm6QEkAlaGiQYDErpUjyxRLT3tGztxJGyRydQH9gafhig6haGl9mMQsA6cZ3h
lXtqaaA2GneDw7oTGFldVaJj3TnwqiwdaE5Q6m3FQvevSwkVsMrYWoLJCgAyhakx
XIUJp+tbG9JAlhMj6wClC0LgFaLGtlOpRt6/cYug4JBaZ+mU+d9uFuCm2Q1Hcz1D
vRkMBm/S4bnwWh15/hxoLyy7NsQXz6CKFGtE+voqbb84pdicg2xfpRaJpK0trbrh
n/YcnQbMm5OUihafbUKG4eKLopf6HFjNmwjuT7BNVPxrMfK5H+sm6bQXG/RFWzjv
cic8b39P9i24rVBzGo7ZUuyirRdGk3xvt6hMJJIBWXOwixcW+1/GD3eE+shxkAsc
EgMFmIHtXr81jFXKQOvlk4RFM+b+OSSaeqyFV5IlAjd3T0zZZrukWz/DRxojxjnl
gdTCshAW6ZNMTWVCrVrXKLdinfD4Pgkeyogw3XgHJjpPlnNGf9H7UxGQLxPKOz1a
Gh8SPr1WWjNKRgD6j79LwSJt4CWl8RaraxRWB2pVgVn9vDH78v4LcXcJA7r1oGFs
I5fn2hVYt7b1pGQcOz1Q0kTlGQdUFx1Wy4FAVl8TQzOaOifeFo6ulduN5lvrNTmv
Ro4C37+uab5+X9aRXTYWQmXSZ2EzO7lFd4N45VS51IporTQOdP+crKZihaqf4ASW
zsZdVXdetfz+Tf/STA03MBidfE10PjB/XBthYAx0dtIB9RIv//VrwK+pGflTeO7Y
/5yO3NfdWY2LhuFqtvyAfvRkXYQb0bxjgUnBzSv3mFOrbK6buQp+9/zKbSBHlHuc
5eGnhe7XwJsgs70hAyUeYCiyePMvbhC5lx4CGN6x8UeFa7EJwE52PC9LbYH3gUoR
q4ZCmjWZDJdaqkBH4F+jlg4oT+14wftqDvGxVj+BlIJUgjbo9KTo8deVpJLkWBbW
/OLtlN2HyHLRxKrm+u1IQXfZsmzXEN0dE065De0WE88wGlYLpGosy9Rht2tkEkZn
4h/DiF6AsmPgl0pNNN04FrOfUN1HSPuUtX4X0VQkA2ZjJ5dSJsxDVkQIt7o2Qvpj
1KdGP1XXVcirlDZQZZ/l+3iROwzeA2G/iTbbyse44cmoHaZH8VN+odv0yvRQQ9xp
s2FY1KC5mO1FxxZ4JsppdZKoO++dM7YOCZ+g6C+0Z1GUqZTxNJ0Antu4jZ1k3EdB
q/HgNqHIp3BJZ/AZ4V84z7+T7kPmd5hhD/5TwvkObvPbCsbVKJxVN2L9YWSWM43F
+PzbAe+ww+sKun66Y/OzN2azY0dxMbGsdkLc1NZXNSoM5YDVyGJvMg4GWflVxfNN
OD9AuFiyhybruNhum0RMCwbp1jtxFQERLAd7743lO+qoMXd0+tKXrpWmI7w7DRrD
V3xrx3GOr7xaBX8qXfYJM7zJvl+t6+l2MqbFbALUwYSY11uqZZTNShNKWKQwVc86
0/wPYOWm4OUhyx3HB2s57C4AL76KcB0t+lLmVd8/0vE8zVtzk+9ZBryhlfzhmb+V
hvTpsb8ju/UMoFOaGPnw/3BWfsUk5xfaYRCyjNl1ada7FfF4i//zRTyxJsd171kD
Rqu24ijFgzx8YFeXm+oCDJ4psA74Bojj/jmjI30zY/jVtYoKpW4lzt7yoqFUggSI
aR2M+TUgiy07NyfpxxW+OCBlYdvkiM150anMkEMcICKJrjWmRL0JJrOFWC0f3qy1
9jHtP96h+ymbsX/MFwF6uaMlYmb2QV96dcIXn/xJNk7kwvf0OFso55zoHDPq4pLz
CjtSaQDvtmTiKvmeesok6MYPcjkedqDDfbXs7Kk/SMRdT29e6tZkrDAlcxXly6lS
2DbtUKNmUgjQNJKHAuNQl6YaI5qAK3F+xlU3LbB/ZNTui1De5DOqBQ8LguDL7HTl
tj5C0WLLUEk/I3JggixD6zxWhf5PIauGHponYK+QVky5EKc4Mb666I8iKJYT9Pr3
Y9XvCx2X1TI26JbqOGq4VXXJLYZJcBRYkZjS/PLur9hnE4c4R1WChxDGGMGwPSGk
okkBgLy8B0H8xUVnPwNxpljVkCU1zoMN+ATMP3+ns0abZ8hOH3IRRusWOjv/G1sJ
o2UoX9lwkLo0ayGbRHcc0vaH1iMHdZj5oPAr3MEHUjWyfzne1uz027RVrzXz5mkW
1giS5LfyOkzVZI8hup6S4++jOXlnkp+1mJhy0DJ4iZouzDyGeLXmJInuKZgq84ah
ftzJNPhklWLd60h89EPOiaI4PQsww+YaJCfhn+Fq8ZmY+9PldmN4KfiVMToCsvMQ
sr/YAy3OaF+krZLtkAxtrQS9TRd6NVpeRbRaAzQyEjE/bII0YRni5yl6VRPVt0kK
Z+ZdC0MtPOLvgR2QtTVAA2wBQ4ma2qvbtwVt8VnskHFL/+K+UJCfYAf+lWc+sVW2
atHOK6H2p43vhU4CXJCXEtBGLXEKgQ6Xt+umXy6CjgL0rkWccB9jIVTV2ddG7CDB
bQ/K5d2FvegWkquAQTjsMjpr/OvSw3RE+Gj5sAU2UnBKvDwd8L18blSz5oGcuyxD
dXMY9esESrHVAomPVbVG++184fmC7RzsAms5A0SFKijs33g56CFFaXV+LARyKYQW
GagPaUyYvMrnaxRsqTmKKMSkt4izX0XvK7OC6KOCpXnzqpIz6lgE1e7BEtUaTNm+
IqyBjetvMNQnAiG4VyOAwkxtD5IQkakWh3m9hg/MqdaTIWcVBJHPfpr8K611DNub
Qp48/DxQPoOIlgH5TqFF/rUXlHvar1pvslq0+DaFzsP9uHWCgDsi7RCXS0kJs626
Dipt+0yxlIZpYuK1pW6Sh01B6iHBq5mx4PXScFNTTf26e5K0S/oaLfNFxqgRJhE9
5R06mz9P4Yi2HyLLJPYqBe4wgCUUYX+SmJRcWJ9mImMV5PdnJ97neVEphdUoSqkb
YGjFK5Rv8PJ3P+VEokbm+qeIMt3jAAi/+CGdcDhx8TJLIETzyf7rfgFSNzxHLGDV
i9AIwwIeZEbl+7al9AjemrTYcmmgtmKpSC35r9NXg3JK9H1FnnkUIH8Y2VAonwsq
+J41J431ZDRE+oSWyW5jjGAq5CX+vW4QM+3J/IR6ov57nBTq9JsflCkxgobfB+2b
+EIdJ/7VNL/jSaB/h4DZSnXf32uU6CW6MiXfYBQLae3krrMQFmJm2YfJspMdpA+w
pfe8xNFNZAO1M/Tfovnq102dtSCpyis96KN3mNG7r26o93Oc/JvlerM6LGKReoWL
k17qJ5gWZxBHVcTZPA+Jh1XHILUwN2zdZ8X6PcZuo2FOsiWavlRrppGJRK4NXXjk
8MG8pv2qNO0SS70h2J93z8hPtB8hUVvcuH8xHEisa31rtwrmS6HXIkA1rTlB13Ew
xMVga0xDOL1gLixzVop0iVj3+ABiuApJhudJY+Vk65Swl+X6X3RR3o5gsR+qUbV1
9Hfa7zCYCw5taafWCjVE1u+d6QGBnCUzFzBPHSBLHhdrp6FXn6Tk66PzvHgeJPTL
tT25IEeYslV5y6ynAjyaYbDX9G5blIx3ulX/r9DJOoPvQzH0Gl6o23h4F3eYkF3Q
FVlGvY/qwSce5gr+09r6kAfU38oeYy2wu7uDrtufX/VovjmVSXEZTTU1kn/3mnz8
iIBpILuNaLWrjQEqnN3N3hBovwG+HHk0GKOQC1YoWpNtLJViixUcmzYzNI01fM5A
ECxAhKZ0YXjpbSZi67Ha1eZmrZu6tsihcrn7VS4/RGRyENlHfZDKuRMy9ecm979Z
qvWkY/7ZAfYNASDCW6kR78wiZvMHIJ/cNrF2QEsJj+PcIZia7XfU69oq8FkQ4WPD
yXnz8E5yttE6K6eKzmyKmnnlFMa5+BltZ1FgD81IoT/pmXPRWTyEfsVN9vk/EGXP
XD4b2tXdCbeJS2LiyyjazGG/Tr+PW9B1hmR9FOWwiJLYEKmU4abTQvHzQzL7JK0f
EZsCkwI/6OmXfGaWP9hgFc7fdRrnmUz05nEDms59jSNfCFJWfVGdGrHWFHNll+Av
1BAZO0Ld3aD4ukZ5zWlbtUqRTHtV1TdSfIPBUIgMdAxXw34ZDjd1THJ0+KwAoGOL
na2SaByBJVyI12uhp5viZPbTYXRoDbfxcV+QcOwefyxYGr+ROiaIE3brCdDb6mP3
kU2Z89VBQz/IXsNuFmgxELh5mmW/xm6hsI5F4M2giQ3gRzbmrUiQd4vnLdpYSQVE
/3O1j9NfJr5L/TuoTdPWoyDEp92EbCmFFJNSmQ7s+swVeUIpLQl1fMMu3QRTXGyL
tVWArkWdwX8OGcG05ba7ddFk+EWAOnok5aeYGGxDTb2eb7eVicRo4SQCEB67mBOH
//4+1rmidZjxJJKTxLt3Z/T02vic6Wcw3oiu/5fHosKvwvvJj83qLxe8jkQkTnqx
W4uh+1NrMEGO1oKiIIforZytI4GxA/RdJnT4EbR0mfQCYU50FDoq0rytrZVAiM3M
ZmOUUOhf493zrCQb9LCf+VbvImomqldoZIVeRl8umH+UtiyzwzLra5dowM+Zb9Ar
5RXflJKGTEbOuDVaYbo1GfJvszP+oKVB7nUf1rTALzNbVT6Y01B3H8BIcdi1qZFw
LBXyK2Wx8ONCLorDbwxcwX1Ul/lVjfJFLXXMLwsRqXrANf5ix6dcISxlg4gRfwVa
PuhSnoRevsQ2Cnc9Br88hsqPg4w/u4vauHruah6YwhlpOPhjYkVlHvN4t9f5Ftt2
GWubB1h8aki3kxDpdB1JYmvZG48PI0S0TXZQMF38nkJgoANQ5Ui4KlbbaookjP00
EVmwXDBwFx+WJJ9vNIkQMQVI7Yt5w44rLJKnHVAxy4gYoIeLj4mmseToYZ9NpcQ7
nS7C9sQ0EWivciJfm4TMLS3q9A0yTI9rV8eQ0LwYlby6F9VO8ZbUegqEyXT56Uki
g8BuuTAyoqcufL9sD2CuFvSwAkH1AMZ3d87w4k6x4RsTvM01NiZSlO63qYWUo+x1
uaJoyFV9CDRA6Qqn93BaKz9nBqYZUUeCJ1dmbH4+SGLp8Byph1BRW4eugZFhJ+6p
f+DcRAjIhK4zSUPpfIlnbJ5fxQf+zvYw9o/5NGQkcRbgVGr9LtvrG0OgLelW3VDa
KI468VHZuuXutOgk+gM8bVyg2CmkUZxw8Q4Vf/iJ8Ty2z080lzvDiGo4c3mjcKrv
SsDO3mqC+ianxel2gJLvYhuAppGJ65RE/njyZokjcj3B0IhMaJVqLpQuecHvtss1
DlBg05paEOQ3ZGDlVKUpSxSvoyuR1ApsCO91o0IzzmwIARyuE4QgcPjZdD1JUfck
uyTLuyW+02q45GJ0rcvAA3cJndKjlkfCLS9Qc2fAm5Op16kXSa4XyLkDoAYyEBAX
EQ1icZlOiyy9d9uey6YFHl5Y7J3usKmSWvEu+vjNsTxTCeq/qaS1k9i1uyzCK0R+
l+wPGM0AoPgg0850wkqBTpa3V9/4i+IBZ1BpR4f6fbuHq6EIgdH+Q2l6vY3secXX
3ly3jC9FtlrB/QFEZPbeHKY/KxYGWZWfX0gi7M3bvaE5jfuitI85IHKCIcOq0Qol
YXiXCfzJ/Emdhvi5X+1t+GKbSiUYw5RWOKdxhva8hatQVvmQLvqzybhCEk5lKoOE
m/kiN/YAXXyU9irk+az8I41cWo23x8soqUyh7etYrpveOIyUIJHJB0C/LyO2s7XW
Ymyutks0Eo5z1PQ8SskmKbC6Y8LkjfqugkA2BAzUvocS/Ootf/Rl3QUDOh+Fw5+L
dShqyOlkVLZOg+wLr6/VX7FvpGscRcoOEYkmiFC00LJ9/dxCsMGZm0bvQ34m+voK
xAQKdeilgN8hhoA7c4K74p98mrW1Qx8DNPMUyX8xI4RFQlRR88C7u6HapxU34gB6
5tkmLfGn52EvxNpDBF7kGrPiT13y7owNLfy0JK9s7gdrjyfubbT/4aMIQptWlrhs
LlBwVE3iOJHxtMQ291gSHJZfcucX9vHy2pM4qbZ983RtPPJ9HSe3JeHtbcn9tblU
vCDusnZNzOkIAt49oynTzEGB3cEbzYFxvDJArOFtqiAwUD4RzOTkcqIjTstVIDKF
NLs94GFaDAB4WAqt2M9vTMHCYf9uJSEXnRczymlinAid0nKqWN96zS4Rk/nzB/bs
vSaMfvQJ1sZbvJW2S1A/yEVWlE1cscA0T/EhPd8SffadZP6kIvEAUXqB2gnE4PPn
uaBUyb6L8FIoUlwGuQmyfWab2AaUj3YwSLxQBPRB+VT/dBTEv03cchJqmTF3K/Sv
onkeauzocSudfhnHz7XE10/s4gMcOURI511cKtJQlRKx6XleNDWiqV5V1xFDJ/Jh
mC7hylKG2nf6CVh9+evXZla4thVmq6yDUu9Ybmd9CsXBsnRKbDLENG3HpPdDk4SW
nnAuRV/6pZtT49uaOlbsklBpZxgxEicTg44SYb+0O7BIBLwSYjhj6bjhBjzegksf
oEQQau8AIyDYanLTbPn/ZP/n4Xqs/rb6vMPXp76zhjGbQqBXGcv8GpNtDEXXsdB4
paejeBwiWesxSak1HjG7mZ8Xcp6s9WLqxtqvXGNIbcmdlzY7K/ko6e5Igq1t7bYx
zg6M4NKjeDEJ/7c/3fduUPpOSxwj5WL2mJCWUb7iJ50emGO2Or15UdACrHK4y0Gx
Vf73d7TqsIqRJmX0seZQApuQYHPglBbdy/P693q681HgXqHD6JljWhgbSAPiRFOX
/pxNCfszKUhhdjv0u2YNiXDcU47A3d6Cj52nXwxWyht8aar/CgWJXLi8mvTZkD2a
/XOavGi6ad+zgMyKNPGGYAOlQX2fX4RfS4EXxQA0nHnDn5s10rbkP9YxykCUZAez
fuT7Sa65b6nI7Q6iuGci+K07YkUGe5voMnraFUeh+jVumUeW1wdAZA3ZCJH8xYSj
8yy8YWrEW6+NQvK9K8XmpU8cswNs1tpzdA259YDM5lvLHD+JOXqNT5123rZjezj+
8njIGWfMvIeyPZ3WSp1Q3ogjCnQn1iKhk68jx0lN7SEikPTEjtZY1y6ngGyMSWWL
tT2farjf8rD8y8AzGhZRBwzJGOhcHYFuq/I9BLaL96y/6TDV3+Cnv1aVOPXxkI4W
9mk6pK1+Sp84aUIUJH5SoIu/bmGeUgtbKTOQ34NhHoiaiob3mhqP1zydnJ+IRdSe
871g1jPkIIj2KYabQeKyVuvnwXigse6cXBpoQP9jVlgtEoc4DqA82JCSV278fDOL
d9aLcweX4D8GQQX1wTsfFbzHIRVj17+/xUdg0dJr+DKf//qmYZwRvkd83wIlBZO9
cAM6R8+wVqVV6iEr2154ix6KBRLuPtM0gTVeq3YSZfjN1LxSx2zhtoVzhf+zirEV
0LUkbJTlLZS/EzqDy2ZGyUtjfEzYpsJl29Cw1WDceUo5Boh3rPKVxCPJaZjrUqx8
5/TN3tJD4iHHf8tJKBLsVZh0E3MQ3bawA2Uf1wStdJO5Z268XVfdlCKykVGD5fmE
tZpFJkfhSGoDNDTCN06oi2WgRfpjwmDNQ6Gz8KY8aQsty8hVu1ZQNRgK8x58onEB
sW+GQzgVtZDYw2ojn59iU60tql7Fbu7HbI1c3S5SVsmO3ZdcDB3XSwlWV8n7QWiW
9Po9rjD9o9ByHAuYJDgb83j9J6iIkVWEyqB8OMCKLvKrlxwUQVfiUZYv54qcAvVz
BqSUzrT0CVaCoiytoug7pC4i+vMc6h4BaeRZGN8EmzU5oakWetF3hS5LIK+cDKCQ
TCST8QijmTO04x9KLdfX2c4oa58ZNFLkxIJNO6H9yyJegpczysBxKXOG0pZtkB8l
iAaUY1QbFRZDDg3CsxAfXSrde+uWPM1jG44WEWFza2Lahq/Mj+HgMsDVfu4201Lw
uzcM4QiJtmAeEo9YJke484aJYiUROsJklGq37yQ72aGOjc4NGTEvfdDddtRx/NrL
Sg+qoK5V0Y4hyg8R8L/XeZJ6WUCebbJTyNE5TPQ/2grFCH76Pp7Dvcnp3kZ1EDry
SFSu17Y0RLy0ibJrfoddWkUWiVMYx3yi7xNH7ZIVyP9QYoNc6wMeZI02dkPXvFeR
2SkpoVlBknP9iBnZH1KgMZXqMALJrd5B1ct/WpKSCJtlkvAalPVuyg+w+oTuWkCs
T68HAbUXsKkNG+QXyvf/3NSJNl42lsR5lVPCMcsPSyWShTImRjlYxb/QDtU5kDPr
4ZsPaLw+K+NXoheU+UlRtmFsK5vSOIGIW9ESt3HE18TwIW6duC6lwDhXAInYPQP/
7hCJcconhS5Ha8ied+SaSRXT27WF0s4QRzu3BEtGtyLDddawrsmvKoYwmaHzsMGg
ieamHsWae/4B/A5SZj81wqNalGEAZwuwxVwk4i/aK0qgr3EEf0TkJkXe3OUwqP9j
IyGKQ5frtTpkpWM9w5SUPf9LzAuAwynCTHekRnJxIuVqAghpqvxESFyuk1tMuIpd
ChKHc/W1LF+oag0gZWi3GGzNxmMZsUC2Im/5ixE6vEDAS2Ik1Mb0DYIHZR1w2VOb
tS25+PdZzd2hoaAA34DOZmaq9ZG32gNB5nbqqAf2eRjhOI6olwu6p9T2vGNE0Xx0
w13oggflaYIgetL/5gymqwH8/N+Ee97F513+y4Sol1fLTCXLHL9EAXQaq/mMrEOu
Dx8RWeIeUETWk2zq9AcCJM5PrTOGpyeT4BDRCbpTp22Mx+VPPcQtVCb9lN4PTiKp
a/RZy05eCU+AXV5BL68zgyWypKh7uRRH0K5nPJHc2IPAXLzufi+WFszwF6DlBYIg
jdtSbrJDCQlt/8qM3OygHpW1KPWCSQuFNG/t1oyvpGbQH3S1RH8SFgc8omxgTEe6
UwHEbN15IPCBtUp1OjwojNqE3mOoQGeQpwAufQoz7k4wfakU54vpF9h5xEVpTc8a
5XMfC74fXNVgFJ/u5/xv1BFmt+QgnsFQxrXAirQ0gVPorPkOz23DgM8U7yLY2XYo
S/QcKpNrH4WX+jlknQRTVMtq3/81P2VYldTbWdzIr1wVE81CDjD+mpDFUE5E4Lcv
l5bnLpmsmnjEphLXmpxf44iI0qhvHrVnbrTD6tPPz9tFsZtfQBeW0E7ZyfisaJWe
TB8w/6dLhqtMl4tQqxNYMgDtLD78b3p4pl3//DiOFrTQmImQOtZ0CuNPJbVVoHcA
G+jvBLvsnlQ6E4EfznY8kAI4M6NbyE3kqTGWLlsIZMohuHI7+D+9pmFnlcuYzopl
N2bec5W+S0QyoOYesiL7SFqVUczpqYnq0ou6FgS3B4C7Kyko0hmEWsT3kwdyO5PJ
01dFuEt9ErRRsS1a5gOqQWNmcQWuHBga5fr1UTHoKXqvzpPTPzBC/irEuP49ubZn
IA5fc9NZiu2WPxPS0ZalPOQEmOlVds3v8SJI5uTPwXSzrPUoQ6nfByO3H6UaIlq9
j/PPlaY/5X+Zb9/deeszy25x3eomIiVQXz175OnuaNyumMRZWo/OeM8c8h6Fv7nr
7xEFjZnR3wPNJh/p96fbHOekgA0gM7GFhq3F1NN8KXpZi5XV7z1Lqx4+ejxKnogi
CRjvqOs3wn4E9uAoX9fGs99gK54ejBKX/2aCMH+y8tsLsA9DYnYixcghSN1ma06w
uJPGThwmDGHSeErFMs6J3bCPALR12+cKsXfdThLBJl5faBqm047dz6Uyan7m2yQD
XvYW1MBEgy4SDfvw09YWeWOss+hfGQf3HjC0oZiaHxWeQTJ2a0yzH5hAXgJsR8G5
JN+8yH81QHtECa5a/I01jSSEGNAMxXSm0tZmdCHgIP2/fOZtKpc4RVXjU+wPiLs/
Crl+f1K1brRxu9/PsSKMVpGWx5p4Ga5/IvkJvLlTylaogGLMHe4sidQd1rpMX7/E
41CfskMaACep/eSR+Xmm/PwJiP/ZN1PAwsmo+NblsN//0rGZLIrsg/YmF+7pcxS/
Q1WMp6PXlZJEVCr9b6qNmzbIgYwhKMTCW2UneBVSfozYQK/BXWxeDZYfN6T1gA0F
IABcZVzJx7+KOZJNiDMciXjrZAa+qSQeEChPe2PvesYjditVc90dcDE3SfMrlz/7
hifx+ntZ8Z3L3z1SApgtDeXWNDOWSwu9bL5R9mrpX4X2/2V5D8Eo2cKhLrLLxi6z
161OrFEdbQcsqmgg4l/g8W7LMZt7YsTUgmisqs4/r5r7rTfLkOGKT9qUzkKC+u0l
V7EBcHs1dNf6NPxxtuwdtUXtv+uvw5xGOCnIIr4Gh7P1XCo3NpMRMp2FfQS+jBZX
YDx8/P7MhOEaplmdtZI5Z7tRq5VIkBCQs3bF/PFweycdJrTxBpEzdayT5eycrn5t
PqP0Tcgr+ChefLQdjF+C53eBiRc5cRbWiI8dt3HVNaths99f3lk8Foye7lmmXZ4f
lSX0MmwWKul87ojioeO/9clknGBPBe5q8s4OHT18B1DxWZxo/G1ZVXvOZAxfhQ+E
Tt6X+ZLA+cGI63Ow7w0hv0o50PGajq1yQ8bx0RnTFw5AeYNZEk/RXN/HboMuiiDi
Oppra4YojvM4IcXMZPvay27wvyGEvaZLL/e6rYtdb+IXkfB+C3v8o1jhcxa1x5pa
XRFhH1Nz2ZxYhMCixuPPhDtE6n0Q2X7Rr7c7fVCc8rVWY5sxisSZyN4NOqCruWOm
Ul2c2qweIpHADV9gXNpLzl3kApvYjKEJGPmAaHniafoQPzBmr72ZCd9Y1L7kumBZ
Jbt419lPTcDL24NUB2cRA8sc+qSqO8nztARWdFk3DbEn5hcZeTjDPe7mljVZALMj
jHCDGAcTW0pjLXe4medZRgekWREWPYv1T0OQP+8t7a2yZwPgw+p2sSvCcm9cKFwr
56zoGcyFnSydPY74kAk5Rn+9L0y7OsU73qvUggCTzBPHFWvvvda3v0ANOqUDANoo
frtV4lgpb0v4RSI7litCmZIWTWF0xf8QuzwI+xyPv/PIZwPN04GUAcZmKXBizmXo
9TV08hno7i83ukVEYiC3L5brPK9SFkQvRrpqXGo2L2aV7DO5KvJJkUus3DCaXLwT
Jg1Sd35dvHbDTYVRv6hcT9kwqVsd22xwnu3hHHw/YMcbZ8KfOTp8bGpc9+mQXazI
Olw3xYYxNh30//f7EAmMO6GWZsVcyjmoq44OQh0YraSLsyiJekkQVvNb/UNRNZ8c
JflDPOjRGAc2QIe9iutewLCeo8ZA1ikGAHmwl9M/bhfj2wWfvw5ySJYXeld8ugIn
ymlcFeK7FHYY3VWorh4kX5+T1/VpTp6N4eixTM4etSmshKi5muNV2OUtchoH/r8/
MoWndVuncLj+17p0873J0Idy2IhFaD9qwdZqlzWY0xGppJmY3jfQBk9I4odjd7P8
PDshhwgEdSfxZWHsos/mA4UTRSaLrdR4Nq5OpD8VHlY93v3sduKSZSC4+tB1g9YW
/IX/7PaGVpO0O136+bGv/r/u7KgUeGZ2b0TH9RK7jqbVDEdytgHknUI9Xsdm1VsS
xD0+kuACGVrJo2LFToRKhV28hoLOjgEWn5s3J3MmE1ZVCVuHJZ6lXNfHacVEEXSX
uULBH6HoNdvZzfX1Junir8z74oLuJSymdFlXBqOAcIrVvTqHhkwFoI7Irr/tmt2g
gu1D52k17PMRTqdhII7BUFpOjyPRQ+Ojc4DnblvDonHJg2GuMPSfd1bZhEFZmUFb
KFqK3v7RIdKmXruL+eCuivyb2vaH/ZlUWISYtn/5CtjxDJ/1eKgGsEwuihFv4wco
KwMFcWFZ/uMXVbz0GThisdTw8/4eD6ec5+AhleGUzJQO7DleDN/y1GDCSykTj5Lx
u28FTeq5pQeNKcVLq8u++xlrPndbvFuV7MIrpQ44Fd85kzHsWVoTmCJemUrguACA
UNRnmUR50x4l0D/UUUgqQAdGMXD5UrT2qBOGcx4wT3L/bEMXKpZEN98shajrinyg
7pecslpIGeOjddXYLdhW+SWVVEpcXCXILy8Iau1KfAW5dsxPmBT09aKaLUFRVe4A
w5ngLTP/ai6wRaSRhx+140XRMmO1SGFW18svmxaK2AnZGcd7wcoyD/UbhIcJwh8H
q41DDk0mL4HzTE/gqwbYW0BWyQKl0Xk3PEIP+qIpXmwoP9kJrz+FiOkhAZ+JH1BO
B5blevH2MKSXySLAT4bAu4ez9U75eu3BkEkvCjzkM5vq3qr1zYpnOL/YwEwwWxdZ
EWSyDVxuophJzXguUYLxjgl8Z6o4VyoGj6Waq9MZ3j4sisLQ0/DL1Vt/QzAzPEi1
5GeqlnvT3yXRTELS7tw6iPfezsQeC/YgoHJ+2soxNhOfOl8g7q4qvigtUbRGRZp4
ZJsbxdVGal1XETj5wRNDREtnLantqCtC3fFDxzXrjRRAb1HAdnzYsgop3K9a281+
efWcvleHDvVbcn3l+NxvEI9TTJrHLjzd9v4MrYntwm8roFEMWpuCM3zJ6IbcWQMy
k6tpFfOmXMyQTwgthbZc5VcK4BiWuybLvwadsoMey5EY5vHea6yebFVaIFj17AYC
qbMurPuFEYYTT5u/E+EzPTaia6PTiPTVBcM7Ky905KMaQoFoUGm+lIxCNeld8JF/
ANA0sFFVURAMresKUiGgK4nIPMqLjHYwxE7814ktxakc789/XVioUGMbdArJJhhn
Z7IYuhn+JEfWqxC1YnirBfEPmkWAy5F6BLGB5gCy3tNALAhAayRzG1gI0YS5B1KS
6cBQQseOSVjZb8DEJwUK6/qTIxGHytiD52lpLyy+Xmb0vaQENmPEa/d75fjquiBb
yWS+z0u5gzvy9zAWNcWYixTV5KYoiJobbw20NHCYPqB02lwmoIDJvUEF2Nqntyne
nXoOQ2qyzEDu+nagSIxnGNv8LRogAU43lDNlF++tKadz9ieYTZDLESWncxyv0QyG
S1AYiKe3ZV0CJdZzFVx3LnuqFymL2wfjmWlfTTaIcXzeFk0ze9MD9nmvwqFJgipd
jEdDeNaW9XCzSBs9Tv71kT8icUJYW/N5HdjIP1isnh4imPbley6VfUeL3vmtoQrc
/xCioZwwAJaU0Ielyz0ztipJgr6CibLGklEEjqcIhNRxo7g/miw2KwCFYZUogtWU
yGs7aAX+UIJh6LLrTzVzGKXoZus6UvLzWJbPdztVcULwOjH82JtodjO0JlCK7T8R
RENakAczc6xhskJ1hJ2HKnBsCJeIFlxTQZ+zATvqSEluAbg3uC3Hfv9oJOG01FKH
Jmq6dpAMYuP9JtZWesmo7ua3+H+wkq1jAKMwWSSzuydusVZPVQWw0m0gXzgksJTN
+mKjoTvzgb4nzFhhyNqw5UoUjCp9POC9u+stwg6hPTwpdpSj2uLSiKW9Pxyy1Iik
RvYsWN6+lB7Mcb3CvNqC2JtXbCavIjPTH5oa7WhNKnJEB9sknIE7G+pWE4n1y/IO
kJOvKmWrI9c6VvMniWUiDNkvvHm0JbPvnD+AbFmbP2Guu7Bs5JmdgMNFFM+dcBOl
fQ2Texd828l8KX5BRcKHBkfTGYgkhqFi6X7b6l+KDrNU3AbNNlM7d2u+1L599wXy
rztjg6xDWB4PE4FuRcI+HHshF2WdT/C/1Okhq4aKwPBKBAo+ImeMY1TVb8nz77Kx
1TM8ITLup+rpegkPbZfBgGwGlVG44rOxM3ugorgDWNMsRzJhfI7LFh1uvCSfp97D
XJhn4FySdc2jKLIS0k7qjfCN/BKSU1sbUaajFCEJosbynW5CYLNQkDojS05aV3HL
pW5rsWYbajKzQkMV3dzBjSflgmNr6xkwcMWqlKXEwz93Vey6UpNLVAlAdncZE+94
hnvR3LcvaUbWnbEa2IG/ugwSaKDTqmwx1OSapybNWBRF4vPLOceULJ92SzaLjrVv
k7Kcy29xM73BzO4miiH4UUn4XzXZg5LQ+66dbZ+7XxjD7ukYSxnOEU1Cz1/GFgqW
qmQFUCP+AChz0lOG2XKYc2BzFZGY5nDtnwUCw7TKnH4Yqk0DRyzzticNOuS3eqCG
rd2YhNSl0+vBeIUsIpQA6gZeMNOpj0Pus6ls1VULjxJPtgoAtly+R/35jdUx/ks7
uE3L+VcoUlqNDVQffs4D3I+8+Qavrd3LetrSOiKkbiX/NtlcKMc1dwYqm1EUqffS
GU/lMAnoZuXhawSs6uyx3ivxFZ7ksH1zYBXwLCmnIKGOsiwoj5HgWcxVA7Id9rSJ
tT8nBo3NW+3mUSkdtXg1EgCKdEuCscsw8274i793Qh68bjWCG1Z17UmCJ/ZrqNHm
cKAniRFdRldLsH16gLLDTJEkpZu6xomV89AI9eh5BRauUuuO4yTM16Qm7yC6/yIP
BCvkSmIgNu5J2oIiBtSaM9yopYQ1HxmY+Ma+CFSVMhRAKRwrh4PlAoqsPGc3f1zu
9pVP454vcdqx0w5/HQ9ktwMZq9eTSYoMWuknH/FztLOomn40bs1JMSy9l2BC97yO
pcGazvTNZ+QY3X6Gk5UtuRYYautCtSiLVFPbHzG8utdtxHSrwbpFAS+0TcXGhqsm
nobnHSeoXppFAmiw1RMZ3hXUAqVtzkz7QC9FCH1QL12ECKF2YvU6mJeQEspXc+eH
bq1RvRBH431UuHEM9QRSoxSN1zKlZr75aufSfLvad0iMSXA+80Mc16hae+h4cutr
6T8H3nGRAqrSc3ImLM8CFLj6qBSieo+KFvPK2TJePkVNkGHCAu9uKfR52zTjDrua
9xSOF2nZUbKUmyFD/ih2S5qrB1z5683rkmfPOqUFhxsh6aZOkteyhn3oBMyYIThA
UM/zoJ+WCjGJD8GeM5m+dnP4PWqA3ZOIRTr3no0wUnxUVQ3ppYauToPRoM57ADpZ
Ct0dbhbDrq9/MujBNhnwARtCQPnAXYjLJC/hUOX93xmwiFHNHZXa3KtMLf9bQ6dN
LwnshOrTr3+Twt57c4d/n87QfGzK7DUn0UJdwDwlZaKay0CmopQFEJ08LtWAIiL3
l6ZtbC8qNgQ8EhauZBxhMgRakHTs9556LzGa4zualAX1Gf7XeIIaZfO36Uizon42
iJm33lSQZMwx+7pgR7bfjvV1rt0tws1m6bSYZFNZDG6KGeVssA7mAKVWyJFEPMfd
5et7EcJrAb01Rxrxz6L/fVJUckBuCbn/psTvFFtkUMnNRLYKndvcDx/XeJZrYgFO
BluPh83VWvVSskY3TSVHaa8r1jWYZVreNit9O6ottiZe4okvhUI5Xm2UjBHBpE5Q
oPkXSMezAxVxW3rPrb1T5+DEFbX5wWPDJNC5mwCd+4WkO50lEyzQoD/mhkiBxhot
mbsYe1oW7yF0DZsrew5ep4QfsORCyU/68hCHs7kJZmCJDZEqheBhulU0IGRkc5H2
rz/hVY5I2CECFVTw2tGbysrGa8KMeLVcQYCnbuNRyxfuSo2FZ1mKK/q4k7qzzMWY
M7Z1kvXUXat7yQ3bCxysRMShDNfognoaXs98tZnUhd5hOjV74xPGZLEXExDBSsPk
vf/Rjz7VY9oa2XRMhkqzdqTuqKc6U0yVwfVhW1dQICR49rd76Aj34IrFm+m/fk/R
wrvCLewsMXgVX8u+E8oBFstuA+OxJuWavdYJAb5DWWHS9/5nA4E8hu/9PXBXXWdO
xJpIx8KKE6CFPtl5jw7NNja/+XOebPRqmNmyCEYSjphzOEMfkhcsODiM1zKxQwrm
6Bqb3eZ7Qh9yk5R6byDZTQm7PL6dqZdUuQzTby5oUA3SV1Pl8fsz+1j0emOL5P3P
7DzeQytZlMZ+KDOIsZp7gGHWJsHJ3NgaF6fa+nff/w5UPJuMui1zDRovk+pBAz1X
Usr7Ol2+VmAHa95BTqVx5bqeqVIX8npM+T54lo3OX/c6jqwDURb8TG6fN1tJthHF
O9q6cXpyfWHJXt6zI5JVGuwMc+oGfUYYeYdl6lqo3ivpATu02leiT83q6w4Bpz38
Rt6Yntmd1r0pIGtyL9vnRF5zS5myhxaXzYQxXU5PaLMz1jWXlX208kbOl8cyddes
dnF5g3WX43hj1R4FG0DYpYsnCABa10F2QVJjTwxSARkEQ4U7FXvUcKMSdQW75Rrn
MVbNPMLsGniUIn2b3q+evMFF89vNZ8czR5PKrcqWMlQEYpXAlK3U5JW4LUM9QCtp
3sF8+4XZrCNEaCGvr0RfHD4PSt+sMBeQroMxdXflwa+hkNzeUw0zaPq/Vd8+bIK3
MuV6hWROllJz7v8tu8dpUjwk7d4AQjRSZ5J1M4hVEg4eQ2xz27FmEChgb/nvfSjN
1f/0aJsYMrJ/X6WxNLWiVgGHPElcBExsuREs8BXtZqqFFi9ox/R/ouMk6+AH7+Hf
OYsDIMoOYF5AhmAnHKeSrSb1+AAOW2BP57eooVHIVVuHwIQnCpBxpTQ/hlWAiDAD
U9C43kGuKDdJtL1Qv3I669Z6OR7bbl0EEooWYEXXd3cnXuDfJAjDnUB9m3tFQWXl
oawnA2ahoxcNNxsLYgD8Xro++SSeO56o/MUpOq9ltaKd/YgQrVe0FNGdhRaNoeVA
0TuGC7y1ndmEI3uMgzC5QkUAFziPfZMQDI/qRLP+qZVHseyctuStkExc5i+0p3tT
/sCAmIITFrWrQwf/P2vBdXCHjXBeLaBbuHkrAv+aiUdh4XbiCzBQwqrGlpAsQC+T
1TiFy4UYE4kXHKE1bx1ATYpszhCcR9X075UP9dvVMk3nbQOjLZg+0fFppXQtC+dd
OZsGUghtu7IPBz4lwnzKSRf6rN3XNWibYRPhcR88Ldql1Vyiq+MyOPB3rpEY7+NM
Y5qEvl2NAuHV7gQgMWrlFZHkyf84jxYNOO54pkjnB3dyokAX0lKToV2/CJAN459h
9w7V3Onrmo7TskpPrhZZSlBVOk6CxUgC6KrCwGn5937YWKx4vpiR+8o+HVO1ojpO
eBqvvbVa5+0e5loZO6CaEwjwTk+dNcIgiesg4Kz+xXA3bHhoFLA1Rnh+uMV4kFXV
1nNqNdFrUZY3i/xL3LsTjGtxhK5k/ulm8cpW8rcbrL1px6wLLVDRxy5squija+xA
6884XhcsFsLHRMSENjA7UEWUzm7fHy+AJSuMVurFTo4Uo1dh4v9VeDRGXe8FsOPH
ZVMWAA3YWkDbI7c+2jm6HRlSUAXhp7kEAGBBVPxu2/7MWdpXqny4nt8pmTcTm3lf
XFEOcpVULWOmhGiUs25PlAHstsJda3/I2+/9ZPPNXoo/uuhPgQ8zVpCAx+DXHUkv
3J/Kc+3DNINJu+WE2M4RSAYhabmFM6K0wdogstURDdnJNrT5ITL4f/cdVHmAA9aI
df2Ckphrumu0UGGop+m75fIi7v1MZl+EB9rYN5Sg97svuq1fN/0YMrzBa3wk7b+6
/3yH9+oeyFt7jgFbnGdtl+KQ1yIS8oLSN1U35gXouHucoY8I3WaHEuV+ARkKaaOm
ieYXhPdL4QMx09VdifmeoTpYA9K4t1ERcdJegkwYhEgqxvgbcMKgVMgs25wVAHZC
fInkWTyajp4Vq7gknrn43J7Woke7m8H+C+qlpxZw+DVnYsgzgZpUzdeOK0+kdSyw
zG2UfCKUM8znix4oKkxfQvbQxtAblRpwXrGK/FGh+xDXFcVIE5PUMzZv8BMxmtQB
OrQeSuPoDzJvjaCx6REmUQGRNVHRKyfx5Myy4mmAAcWPIPzBdVQb1sgS1Lq2QZ5V
XVB8uH8HStnoOk0w8IL2H6HUP2ASqF7QMxIUwzU0ky8f1zo9xNbr2yyeNnX2LVNf
o13lzF79zQbyzdhaD63soSgv+el8vPMNPWiDexgyoDbw2RzVvS2v7JYb7uF825ZL
1UE1d4yDgDdfNa/S//ZiGvCQ58jMMdRa9LqXRyREuRjrmoxhIDaDHBKf6/L+1+kB
y2EETj1p3psS0gl3mn2oMwQY7y+IrPfDlCmMq52ZFp+9uFKBowrEPpqw0m6nKMyu
7EuNn4Y7jGeqP82pBrpUycNpYEVAfHuTgTgCXB1fozg2Coiofqy/Kk/cOzvI36hB
bmPwa0zLZGyMBOcQLnXbmHQBP7FIERlBJmo6bJNYMWd7e5ENaKQK9eGmYpUzqqbi
2N+SIxp71tF7E31i6mirU88+oBT9oSrHuYpFY0Oxliz465YTcqHHfRdqfrlh6bfA
MlbNR27EbQaFQ9QvZjBedBU7CXiZ4lb6KZC7ctF9/eL3vVFSRkPn8u9uxY8PbABG
mKE6RCP0NRDLJ7QiwDyZJ8pGbLNOGvwwBM9oJR88U/W7IigkwFFcmtaz9r6ZIVgi
jc0MDajbwcHXgX8QmirMuv9Y4JBtR+HepyodSPyTGWK9zJ6A6EPB8hgu1YGMb0G3
SWsAYaaUh+vyadmJG/cNGvPfQ6huLCmrLdejPnyDDTLP0FT51+s+iDPXWuuwkR0e
FiUv1Gi43QNHQN0X8nrKpAzoLOgob/OI5rYuejvegPcFtRlcILQAbI+IRTlIxklj
wVs7X5X9489kw7OS701ElpaEIZSlLxDpnmEpwVkLbtzrwgqo/QJdtXrMA5M/mgmE
3PEuJVelW8inXEc2w2+z+McY/HdcaoPqnWoWbts3sShP19g6kLcgCpKBgifjQSQ4
JojgUO2p0Te5az0M573ZoeyTVT6e6hs/e4z4YjzqJzsUc39zAR+rpuFI/5Vtg8YF
5W5OtWCXBD+QlfQ1oAsSmoH0BpFSGvnmXF4la13t9fyG7ELlppmaDGY59+k7njV3
He+veVR5UXO8nEktYyt46RwSceM7NHP8hJdlWobfbjQcV+TWRp6L+Va+v7u42e64
HjnUA1XWCajAv/yXf3C8o/exzX5giIeXIxYy/6pPyPKSvywreCk0Pjj/Z9cKuOX9
LrSHfjNIQy/Co6rreWliIQGzuu8Ij7G1r1H4BgE+ekpKtRBRiIZNF7i6hgBZvEG5
hLjOe+EHzyVt+CWVo/pNnhTsbT0fHr9PHC++LNeG0v1q4hbasp96ZlEiVxh2DWtB
oSypdXqk4VeDHhcj7PanP7uC2Q/cfzalWRyWywCyAlgKIoLcvtUJZQ8lTtMgfJ7O
yew50q1Lap7Mo1dvFtjf9nYvBSKL8YacFT0B09hRtAsVyfRdzxeiRJPbRd/J1XVD
t/5ct0ceWWHoj7N2VY8Ev44O8Rvz3oND+iX63P9QdaTvnrhKViFhiF7z23gTDTuK
rXfGP3yZ/EUF83rLFMCVGXxwVadbx5AJ0kcioysI1N+ZBQmi8t+QO4YRbM2EIZB9
4VHg7SmBBaMZDIDTDwcIr7YqBhPNsqFCHGa5sVZbOtCvi0HqKmBkSdSOS3W7XGJI
+QmJw9advbkbcnnktI1IurkraJYabukNnZTFtLgYjEJQc5lYI69L+LMiP17G7B8f
hgASIUpIyeyGpVm2KN27+JUNBzNDotP59nMdJSrn6MN33o0dbVD7p0PnfS/22tbD
BLZvika99k8+xpVItgKwkt3SG6NYJNEM6fhXd7IfAbNajDCmqOyExAPihJwYhAVn
flhUjLdz2maugVTyWn9Ujiz3ARyux/kGX5Fm6pwDZaBcUmEQnBIBDVBIlOrowKd9
PmzD2QMVJXFbCeNawqqBrbuWGxPwmU+T9xiykxfNnBTbj8GTd6pWg1Doo7jnBCm/
xnyABGewGGNoKMUkIwO4WT/Fv36mGSUWOYrJyD95nJdTBdTta5RKHI8aMxqRVWpS
fcvFfiqj7l/w3EY+Pe3TS3fPH6nT5uKBtptpFu1+NDd7EGmI4eNOG7PrUGZedd3D
uVoTPP49IfxLYKu9F1zfi2Kgn+LBKKBpKf7n6ItTZU6WZVCP6pXpXeFFJbmdQXav
tjFu6wJy9yGBZ3uZuOu3PC7pDgBBbI2NK13PtSzQAgQcD0w6YA9LilxTgZeCV51k
IxY7tiQlggOF33gzRza02/VjWgZ+Y1cc5PQGvotu+s2ptJBszn2CsyO2T947GEMx
v6BAOUOMSKtQnWxskmIC945I+UqThdqLnaPSqo2rKDQMpdUfuWlCJRnVET7EY23P
IMqhlkJEHsQJUfY245LPR5Vcrk2pyYzEWRbouRb3GAbCHy7I876z0UXCmKfx/Yq2
feVp6eDC63YPtouy5jN4dxAmVILOVcm8bT1WFxSjpgnhvju1y0RexSbzZoImegUY
skpnIpHK8f7ya5+vPldJwcGVfTQ+PCCX/35Fgl/jm/BKNJRfaRXb/HVEIvCEIOeN
8a1xKybD8b2dztWgYE2sMD7HsypjEiz1MZWbLjStUv5VMkgMn88cVb5ByvCDJnE/
e8LZ+XgvtCpbqsHywwAkFnOp+/tN+TnnZm0NH/TYs5Hdm6nWDeKEtOr8Pfl0SPEx
oS3mNZKoWMBNDizajg/gFoFD3dUkA0tRW6wczycElzUL+QrZ1Wz/RtziVXBdWRuC
1n4nOavHsdHPpYI34P+9kbL/1zVFcd2HWjP7waoUlaAsZx0Rf02e8yQazLSqiNPS
BfypfrURryzusTKr/ZOl7QsKYGQY+J9kCRW8pPOS4+/71ujX6y8wvYo7F2n1TymA
LzT4XxwBCBM4eJDtc5ntjCPLZAQrcWl/Bm/VBxs8qgdu4RpU5AtivKQoGlls305Q
G41lGtK7DOaPfY8INQi9XjoWgri3X1N6tqFSFC5vHCrxirkmA7N2cYtZ5w9EfQ/G
UZk/Mlx5cRy+5p+dsOsmUw5JCR7YGUSa4w0Czp1rJX345SzDkR/mzzlxdgGb/ZtQ
DBLUqmT6peEmF9x1eKH8kYJ5C/kwyEdHi//BStM1xzik09xBzioRjzE55zqjvUWL
55Q+j3l6TJJ571/Uk4MynbCv1mfnBiszP34pX8yEj76fxQnQLoApoaKeip4JXSzz
/inkz2hQvFdm0J2yMgkqQXbYeU2bzZUXD5E/agfkA95eGQZMbJCaipVFTexsDJ2R
VwLZbDBJca/xR3gBgGBKV8nsYIuLJbGtkkYKwoyQZNUqjMhBCA2k8OApIpmUFU9F
D8nMX+bd5448Nxxm37URtiAgJ5yWtfU6iJXxzwy1qYxcaXmnMDrByEnJe6EQnc5T
Do0Mi7Sh7e0JkMczoNgRWl3wJUM5HpK6DKVfN01CB0F4Ikeoj6m1JgLI6/IaQVxw
nhHO4TPBurczURHDfL4NcGWIuKHbQA3aTD8M5oDkXWAyT9Evx+nVSeoaDfhBRi2q
/TnIXw0iZIvUCAE9Eb1UY7ckS72PhaLLQc+VkZgM5QyvkZ08omJpFJj6bQcaUoHn
q3cQu9lxFc/rRTLv+rkOLbOgs+VFERovdpNg9GzX4XCwwYmKsyXVb/hrUZRVyTVD
du6gm4M9XVLYyqlpSqt2+ijzGvMOf+kxV7DjZBbgjLynoTBOLc6ZQQBtYzAEj5Bu
bhTvGBn+DYL/igQdszjcE7Vo6eqC1gcKGwwRlReoS7UVuKiJ5bwWzknsXEhxCGKU
BOnCo7uVw3KHv0xQuTAlIXpqlQ0OTU6FQvUgEP336VHKZOm3yqzFU8maFIhdg8YN
xbJg9rXbX9+/kNd3vwE2jfOxgLeBxxPwkk/QyPbTTAXEeYPvgBhRhMN/n617eNmz
e1S5rJf6SSSLOwRoSKUDi3CRfaC8BW94ZLAokBVjGZnnmfug6U5DtRXFyzwmX3Lg
VUIIx7Tl1C2RtXTvpm2HwBPmk+m5v2x26PggP5CdBX00lCxmt+zUa6MdCkXQ4U4M
VnFjJCRB0Bl/kpiELJ6C6EAIALg0r/r361q+PzQbv9ZQX9ehIctirKe35pQX+hlf
4Lwma5+MK7Udpuw+/Mk3UkUt31AA3VGa/BBgof9u+wqLrrdAKkxc7+3kbi2viocf
Qf+3SvGsFk1PGqLVJ2Lu2SpoNpU6+lt6Q72INi0V/tWp4CGUW8d6sDF85e07Q49t
WEazJeNEl4hVPGxbW2bA0XAaMQNhaDFLdQeOxBAV9NvgSL5ifTDlyVb02xR36mxr
/eW6FzYeYv0QtGQ8nJfmUL61CaSVQ8aUX7tqmrX+5fafHBsAz1g9czdUGWAiHAcI
W0LNit7DPGxYigs27p2pOTwhFSL1rifp8vX2qj+3U4Ieci6IEA35CQE3j78DyQu3
PAaEy+JMk7RP6c2QSAtZy3b61/Vr5tDBVwc+SJP8Ls1I8bxYwdmPc4gJeHgUV6Vh
aK062Ec9y6umWYc+Q5Gd9Sy3yfhZ4XTK1/HTALR+NgWMWvzh77OUL3nIGZ85f+rs
KDwPjG7OdgRn8NzERO++rxxpPCmmFU2pdoZaG1iE2JAfylIgpKtdBDdJQwdkXk+8
9MFsKWCRDVC9dvRJ+kZJPxx2iNFq28brO0bfMbRRER3+XN2Z2H7vCDS3wCmk31p0
YKyqQDiYPCRNhnrEcSsaedB7Mc0DhImRB2LvSDwmrnAgQ7LsDa1Tgp9ZcN5vfxX6
DblkDpcHwGrRS5tOABIwYdhp4yAyzS/fmCkq7Oz/wZrHtSso02XJDlKIGg14AImG
QnUnhVARmyRCDZg4rP1J/8G6KlwJPbHrtvLlFrU3CaiIT/gahmZkZZ/q2TviC/xg
xqbC2GmMNBLfZUZB0HhWy6upGblr/fbkJWMB+aA3OcgNLW43an4pLPmHsLcvyKuw
4XcSphMMennJFtGGmjNMB9bx/J3/jkKmxaBg3IgBT36eakiFmr9AHfn+vP1ED4C5
nnnP2PIv+oEF3uI7XuyAG1am5NIApg7/Vbauq0Ro0Gn+dkIek7PhA1WBLrt+UA7Z
dRix4IrV8nEFUhFeJ1TwcUQxo+IchfCs+VhmNjiGaJD9+25lyrdkl8gKQ3HJypBh
OThHsZ5dKN6ElD4DhAR3gFIveRsGvQDY+afq636PHkgLJjQfHoOmPr98lsw/BKX1
AE/J0uGfdt07jZ9lmMW0qSFFUOhUoLopUr1rIQ0yIavsWe8LbSKDUwqZaj6cQ1tZ
kZXr4Sx2eFqd8E3B8DESQTi1VF2LH0JUw3g14vt2cJEtXlsNb++tcE3/0IE1eQW7
aQLz9cF0RxagpBJ4MmCMuHa17T/Kvtefq5latDwR944JTXL8nspiZIitZ1efx9bt
KgbSB1JIOXWpYjD6SQZZFlTH+Ya5m4yh9SlgBwgpwS2caK7lJTDvrphbgPJ0yk52
kzr1rRaW7yCRfbji+VQGQb1TUFoVVP9iJ6RF4nvwmpzNuK4570RR5fcjEBQnQC68
75wyuIl6pAY3iLdh2ky+ldWOaJo5d3KrUhUMv5s0EWWs9xymO58noI8r8NsEYgOJ
0vst8RSUDxG5X0NfyV2r5nwNMSJ4WsbHUWKAxihJW6gVp5lXNr8/xEc4+LaEaiDp
irvRRmPKIOO12hMHUXzt/QSWxzmRk1rUsjx/we0qW2aTpjCKI0MQOBQykEKvr/0d
169TBJjatw8+pU6L7/z+MfjRnOYzF1IuYHtBqMMiDDlrYmFUbW+F/Zg03/FkpiIo
+C5Bj0y9NSlplE6yxq89G9MGWk4ss0FLliux4YbBZTrTM3oXMvFDJIiZmuLwkOLt
BSEg8vtPYIuiVmz0HPWY+9K6YQSRzuTw15txmslEZHC/No6JbdhNB/App4EifgSq
v7iLITHaHJ8SgMnC6VSKx5AJ2lIMx8WmnTTFIA9hDzIe9fPV/yoWB0O9gcR0Mnsx
KGpKLQ+L7g6ssl+690YQt54Deod6wJOPPLDSXsDEGulCGE/2W9wNrEVsEflC8bEz
UJkHlX8R9iXs672goc0hzuAGmbS0bbpFXwBfpoHARJRQJGf3C51cDzbOIozLsbGp
3352aHOC738ho84ZThdoU3nvFq68y0PYU+D22S0Vl+zF1pJRo03DWcaqzKb9E1lp
jNvgijqxWV/EVcqinsCQVVPoX6mMKGirT/uvt0kVg3HXJS45QEmcQYOfQqTXmYdB
ZzscAO5saUuG2b2Q59UeafY1nt5hxATk9AgRRBZI9XcWiHw32E+bGEernp75uC7n
Z3tCn9jDsMTDB3O+IIKIecyjszneD7Pu33u2ZeHi0foqCfT+ix/EHovbXEEkOhD9
1I4eKaA6sHIUGFEoafKxVbWA1tPYcgBMWTDZn+WDz34q50EbLVP9rxsqzax0vMWw
QNUAhiS/VK3Pvtzt8LR82OivJqiv0MbMhmx59yfd+5aXwd/8GuiRFdgDBFkbPqIH
j9HOVai6Zaxp65zwBzXTAk5kEbQP7vgIeVqX8dlZ/AxT53gbyuqHuudlR3OQdERJ
RJiH7tYGryajAZO2vOMXHgHoShAuW4erRIduE6hGDG0CKwCt09dmRnL83Ik2deVN
rwbuVmetcLcbp66mogfxtlvW5oRyZzTh4oMLqd83hfbGpMawkrBkNpVsIyXZzAkv
Ai2j7gKzBi1FKYJiNUyRgzZvgwdykH1E5zUYVlMMVwcvENGe8CedD7L5a5BfODyw
zrBvgS+KwZWkNVE5tIMSX2AQaRRxY7PJflMNqSGGDU+1FomK+GHerzVkCTTo8S/h
ILlPg7bXgp458XUpS6koVQeZdzEr1I7TrCwAjMwMz6VQ8Kf13H44Oe+OgbCXfkPt
lUxQ05BM5QCvIc+6vfbNrShybCgA6u3EMZVRe96mucvrc4wqy4pOAWjxIeOIu+Uu
0hWLObb0SyJxS5Fjijsu2eWtsJ5VkL2Zgn5ww8eeo/uSmD8SYx4yFIogAVC79tBq
4KuCYNE3IoICIKs3VhlelB1k5ioRMIUbkbsGkQWfyn1JQ8p+WTF0z/ZBtXmPAb67
aFAB4CkAFm79hZu4rYvZEXVpJHmH7+mFgD9UekzdxyqDvmWX6qUZDxLMUckbfRQI
z0TUa1MYuMNYAbT9lG3o7Rw20oiTvFFgBgxSGG/2yiL3mgf4pfusqqOqVM9dLmdJ
x1YNQG2puidZ1jYOHQTb60iJXwyfK9Da2H5Oxo7WfrNoPhUwaZp5XpGFaNnrXCIf
dj9rjA1R9UmXnEIOQpZ7xO062BUoo5DsWF+i0yA0fLcupSVhAPxE9e48Ie8C27vf
h8tD5ME0L/npiTlghofnqZzqkNsI/SpLOX8k+pK+xo3rU/07vC3hGOqsbaMuhQun
bU0FtBMxKppRsvEwioYdodF93VuFImahC6laBRe0uxvd7B0ysuobEfa7S+hnCdzV
MiOGtTcvbOZFYTtPYTQ6pWYjRadIQVEkumegwr82FcNd/VmYjgkzk9/wRz1KTJzN
muJs3jcqPtGB3w+Jgphu1B3JHKtM8SxiuDP48ylHfSelc6UUkqdF10UEnqLrx0C2
uUDbatMKFfo10bYG8grr5vAgyEz2e4CVwjhzdtyw8hCs77XbuU3JsGTpYNPoKoe1
Uhep5f/Rem7u6eq/PnjttQnnby+XkWeCDgr/aK2DvcFVMTI7wYxmcAnsVD//wOHW
oD5mDuPrMrDMHTyhjk5ncOSxCsDBnyEW9YJrHCvf4SLHB+sdhocf37tQ+rzgj+Ga
KX4qiOmTHSeD6E/A6ymEFB2caOqE0oNFhSd228TDUXubF872vjTjusX/lmngWOvJ
IQlaicrrm1Cwj1DpEf5T3eq4Xz1nPEvwUSdW2kFI4SPnTDi1e01cQ4GBuvFdiphn
BswI8PIWF2Ur6srAKB/7ei801IWsyeIoWS25JhdJa97pIamR6hAP8xNltwdMvJKR
lgDgQFOoqgEFiViPy/St7CWA1OAHHyv2FCvaNdRm8Cbe9rlfI2jLzkoeJaKEAAqE
gMirnwtmirQJ/bZ1rgPV+hvl8ALtTTWW/Ktph69lP1S/kJGH2weq8Up0txWTz15F
M2RDyvgPcCbnNwHoY/KkzZkf8/9DMrLiHFYZs3MDRWDqJb0+2pFWVHERU0EoZR9s
SN39ntsDHsi4Zgc+Fc88VSf5Q933x7dSUn6nzdV7uwjWAaqgjVb86Y9EuN283/xI
oUnAeOkXK8rigHb4EXtaiDfMJVgaH1sYfPCXoEl0abbNKhKyq3KMoevkPs8i+RN2
i9Hpz1odQs50442ljuRIJHyqfNqEENj7yIE3vdvSxeSc5l7MA5rbQs8TgBj6id+h
cffdUOi0SCtAdWBKNHvo/+T8lG8/VnUSDywJnbKLbjB4zEyIixV9qxbQ3yGdFI6x
IW9ksJfJrr07rhvoDaId8xck9AJ2XXRV4q0XMfDnEmPVWrzXi1oTv20h0zpADPcU
ES5cR3EF/pc4Uwu8/3mh8SuKQXSHPvVS6OwhKY+HFr+j5wqq03CwBz1RfA0oA/J1
WOTs2tp8vXFhE9nHXWQJH4jgggRRd0pqgaGELmMa6hLh/+rD68uVg8M4e9a0RPvr
L51FjTIbFX0w/to3Afm0ajhU3J6Y6OhC3/ooUBF8P1hZY48lCuA734oDjyDXyAHb
QWv28af7lOUI3eo38CEN56W4Vx4yon4sbC/st7XACwFg67KRkGDmbb/2IuQyugm5
P0QZAvtF2QmKq9cYygt93ed4eICWuQED5zxfVAKRLCI93UPwNe1NR69OdeCv8MqO
MUZSMXuGS/5G1UnT+uEH3AedX5iVWW401Nu2GfTR8P1Uex2WMl66+QMasoP356Qr
5SG+myzIusT9pg/snfn6C6IiXt5sXUbBKuQGfdVQC1xbdJCe6an5OnmPIjheTMhY
HBMN2MZ8c48Vztscqbjby29zarh/Rud2LuBVLeVA8WPA20nq6Q2sg28g811pU45v
NTGTO2dW7aihW2tm0AJGLMk0mSaZRom2S37x1ocbxtAjVZkOlSk6EzYieEdPG5Vh
y5jyr8P7dx9wi8urqelo6Y7ZEN49tvuanx/ClmBQ1DmP/WSBZ4WRaB3UbnTMwupY
dsp3bxNlb+oTsBIpU8s5eQ8b8GD1J73LfkH7TU4zvypeo0KKjbKyXRKF4u8DLvz7
J8Qb2w/ww2KGixWf8jFwoGziPZ8oKRqoCw76xnHKELNyi5l6msS1K8HrfqNAIkZa
n6mr+8+9YFSVcoywz6JS0cOA02o5Bpz7KAfJkuAg491WzUb8suYXpWzJUKbEOt4j
2HZ07Wc6TIu8uZlhB6uP9QTio22PsAYvcBCOlRM5SD8lHnbi/Tm4xs8Nd5TgtYiS
tkSme7rM85ZI10D9mCJxcSSnRffhKUIA+J8fIoXs2+FaPSwANsxKE8qwmgowdk2s
xQWlQZV701nnjC93n9c6mp/xg54P7o7d3A70wYJrfFpN3Yxl6rs6PyM5IKUFrsqe
lKZrRdKU2zR72VPuDC5W4iWEXYPJf2ujomc2kE3pIDqRI4UYorDkJLdR3Go7uvdB
fYd8QL+/OoCNTnlMupiL0+RTuO+WxCa/gMnj2rYg+Sd9+RiEeQbzHA0PtQzChAJ/
UdJipq5Fh9WWcs6lJH7Vb1136gy9m7bKk/mIiIHx8AXDNmMmEIpGTRvcAm9g+0wv
gu3+ixNjTWZYaXI3DijXlaPzyC6t1wnG0qmbgpvlUfPWLqxZbpIAPIzUBAPaBCz9
1r22rgv3ACVMb4ir3w0diSH2ReRpicTAK9hZ1o0p+qLjaYnOsskuXfbqp02JyPIz
zaBijvhrKlZsPNFQAh5qxP35b+DNJ4CimHCV26roh81yEVNJFvmyBSYCKAyVKroK
7zEnW8YZNUvoIbp4eX1rNxDRAzhhf4J7U2ipMJ3WbO+II79ApSbA7wiTZvFaeDUV
OdeKtI9QAFGroq5Qjje8KOTHyKB0Tp0YxA/iEZ5lbVwVlUIqw0NMTC+wHZ+xLmel
OwfTWV1Jk/Pg5OA5v7IjdTjGhjrY8BcTaiVujsOUf08yw9KSMDtSDwSfxo2ONJuz
QhTmAq4bMO9XTQWCPZAzhlV1sD2dz8WGzNzUmg2hb0aru6E6g4fmi3vRiYoEjNpM
tISJieMLBmv3jUtAU1685X6ZFc9FdW1NjHExkxCzcAIKSaGtWDqgAuoA7cr3th31
YiiuVDzu0enhOmtQZNX4HchM3/PGp+GLfv0LL6sVGdYR9Mp6gzz7/Zao3JR0Et7O
6tXwrH+cHOmfe9joM/QKBaOrN3+6V9y6kJb+olqZ+FjAJwOa4SkdEji4Urh/svx2
G1V6T3UUMkPsm1T6n/NHICMtCTPzuDYpYqBLG9GioquGLei5TcI54kcHlMXOnngO
nHXuSEB/wl7UDGxTub09nKEsReVCOJft5X6q9iORWvYrFevJ/R5j+rP+7OsKYBFH
dii/aZXHJFJ/eEQ/WBnxx11qN6lSENYo8jvee+rxxUTBbOliTW+0fj80X/mMIzGp
RJT4uJ0n0TTn2Gtf4kZ+5V2PkPWlanMrAP6T9chI4eZeJU4tSjbC5Frv7g5NflK3
LGmksPZwOah9s9ihtFodo9N6BEgQrKsBqgX0YqBJv6QQHWvWfsWjRKB4C1V2E/ek
+NSl0IY5hrIdZLOdwqp3alAibUQ8REnrM119mfeYxJSQ5NzNv46NEMicUWaMLdrX
QIJ/N9lK/BK7QmrVasok2He/2KyC6+1wlCZr+NXiLfGsOGQktLgAr3Cz9v+sxhMQ
t3LsRrL1+OOGcX5Q9ABdeacmsYjKoTS2DtHf55nscV8pdnmEbSBoKh9ZtH0mTki8
rKNmgnsjzDKwANTll1sGdcZiQ161EAbaxOU93d/nijqb/Y2QnmYOGDPVPYJ44LQi
Y3UWOT6ogyvs+DyHgbnw3NhMFziF3kSulrxiKEjbQP1mhlI0o8EtYRLmpzNS3JOC
XTNaEvCar/oQRBa0LANBg85L1e7W5U3l+hKvL3eeHkBjUmlZwxZP3dd+ntJR9NCo
tDXBg7EB8EsJwt7jGu7m+dm35Xg0vx2KHOUsMHYP0nU+ZedY9xORuXMRVItpKqJQ
7i2WG4AxESrdeOpVJBOkotbWKzcBcxWPfKif7fXkrpqeAPgZPKULekBuaQZ8Rbmg
NMP6yg8Cy7Wfu3cdyN6Zr0dP9rDes10exLFFkPM2VCT4eJkx8aJ1nJmrvZP52cVU
Xmr9Bor3JnzuC+fvJkIuYxgxokAltOnbK9Ej+X3OK+1VpSO297CorKmG8FRRgccw
GnXa51nE/Rhc1LdSly3nrLGZeU4WG77bqJxry+3Iwh1TltBfoJFowW+kYagLexQr
MX8ruVvEfM8cE5s7idwE3NvlaWlx2uPhXeGtAEwVG5EbYVwmpXcLfF2B31xd//ZQ
WY8YBB6ZHkqWsah/gKY+dgP861/7VsZ5B1FcpGAJAVMnQbw3f5RtXBwBlIElNkSl
Jsu9hHqn8RBRMP1rqt+AoFLyN/Uh0HbkqgT6Oppp3PKnBq+1PM34b7+g5g/UOQdu
ssV736wokpVegl68rRFVEk38o1HqB+H1k+ExpBt7hpH1ZRwdbnRg/h/I37Hkh6YI
xpJ30h2fTXq8MRAtQTYBw6V/91MejGgcNCc4FR2Oe/a8+TtyvTcMcIa8i3gSWya7
Fo7oCKX7eAgGMIScabaJRZfft/cnUvXg+n3mQE81GunlB4bDrN8wgtjyJ9MhctWE
YUBpSKM4xs4j693An+E9aF725ggq+hA2+3bAsOQUpmYYtWa6y47nqV6RtRUthawg
S5yay5q0GoeMxGGlh8Sry3U8JRhGMpPWTgi83lYTGBZMIkV0C/BKxaieqZgbjH/Q
F5ci5kV1jjxU49Q5WntHLJaoQE/uksdR0w+D/5jge4dlzAsWQptFlOTLr2D5S3/y
nqqZifqBPt/Xjft/k8HfwC3L7mFroRaWhDNk80R5ao0Ki3tCQm7AuwTKlRukeeih
gB/+/H8iz2dzCJU9nwl4nNZ8lhM+e8W/pSYEsUUTvbPSj0HMCxEvGXYY+iyBzaK2
vD4IAdzICj2ZQiJdqjmZi0HfnIt0M1wfc0FGwoZw2abxfTSrzVHs8GRfzQRXvyRo
jUdBoBlwF9FCmQ0SrNXiTPPRG9HgCD6+Pd7jaC+JpuYDBx+l9DqWi2SRLwiVmgaL
LkKnowFk/Wq4S8aLKbyIjOCbU0KkSxU6yNbO7NlrtHkQdBs4GH1pZEzaRf7q2iyj
wvJ1YF7CmN0zySNtm1lK0iKtHZpfgnosIr+YJkWT/V8X4vf0Edcd4B+QSnuZXAnB
HXo8vjABRS2FRyCmxU9M4QU3lyXgDh4akLn9XVKfQOzIa+xZ8Fikwt8HCDArLuhE
n4KswNdN2P49dpVweZ5Fdbvxj0LB2Lx+SEvNvTxP5v3vqD2tSlaNWNfChvZQkv0P
nvX+KGjt/3b5rQnvdy9wDmkzuPRUZPaYn9I2nBFsWFrsXuoTnn/8v8Ri5/ZX2iNH
f4Auvb+/+7jLV6SQwYGksuPl2iSCiVC3QuUiDR/h+XGvit+EEoVSSxk9oyixeTrN
VnvGNQGmL3EIeSgUXJ2JMfSdfNc6LQMN2vMpAmcumA4L+1Fv4mJf/gTjXqTbGBji
y3QLq2ZjDWCBrcrZXcJ3GFMAptKVipsLnZVsHKAnAsZ0nKIvkfEkgQQDpsUH50A4
/F7DP2ku/bUnxxbGqqjpHW+Xxexm8R8lo4h2fYkOaCjs7VRF202IT3poiSgVIm58
4FrmrezT2B6D3D0m8RrR5f23OYNGbqjkqhS158WtIFi+f2nIG6sXudpe69/LCMWG
E/jAowyvzYLJN1rED+PbyNeJZ85WDyNcV/6l9eOjecPmS38Wj52PAp3X/ngohQfO
dujDCTOaqCRXM7quMeGFoAdFLVJqfxwP8t40cENC72hoSSzxF9SttTHOb6XMbbem
Fr8i83ve1b+LGCYpc7cQeg3RgtIYrXKwUM/MTf2H0VjmajSWCc4viNI80BNbcIKa
SDKUPnvIFQz1r97JdiSy+HsZayGycLBRimcaz5jZtWb7V3sbf/EkoiV/BTkLfbod
rE/kaPrERr+kPML3CgbYjd3vJzJiNMI3W+klV9EZ3mtQIjZJlcpUym0RfphcEE3E
18kcJ5tEPeOgIES9rfowsq5azfhx7sdBv73kNQq0PYt4LboipjDGduT8TT771aoe
4YFg5nuTSK7n92wkKMNSMM5ThrbmO64H/ExZ2zmA1eVtBzWqRTrNgaXIcjqKY1Sl
Urkoj9KOvmpCY4no5o62cxR+Hisxq3t9KEn3d5fxlQ6UhePv6xXG+s/1qq2rvo9E
l2Rnl6++EjiuGKKwaQHxRZYEd+pESwatK6D4QuEjTuOH9yhF0foff4KlzsjPjgJo
iCll/k4wXPNEMqMubCLxihSVmMGF6fe1LsDEVqpauIT9P3WGyQmo1zIDZJTEm927
j9lEGghf0ftl9B4E0ERpnMYzjVuKDvEalQVx7yiOEyfTfWM5O+ZR4mvOszwiDF/P
yg0g9WbkrUyUlhrJ9XDcHVRV158+TqVZ/WAGn1hS7UY9s0kziwUyASshVQ6kQXKq
xLo4pMCyvwQRIWjdo279XiVQrj5zoLrga5glIUxGSoJ033d5q8Rk2SKh4lry6Zo2
hMaeSE7KiHbWneKs4qZBS40kssmof9Rzwg0obWvA7AUoS9R7IfZ2paSCYkPYZQTb
xSoqJDn9qliaNIxut0sgY5YFGAMvYRVj9lsXR5nN23Vl5uQ65NNkOsDPyU7M9QKB
yyrqgEjhKAkFnWqpE1RxPw/wqtBEdU4DHtJaVpDnvhBpwGw3JDWB6/G6LHUpYj72
xuQ3h72lCHfXgPZepFgxo/d/FEwadHt3GpR6vG/E5IilAVImBM+l3pt7i3LHOBHw
7cMVc2q6WnHeDbh4sji581UuZit4hM0i21Jt1YxhihoDd/CTCZHBL1ELsXLsffsk
ggZtOV2tc7ac9VrO3xMv4LoO5oy/fJXWtyiPwWJGrEg8brPAmRYoFdm2ujJ6lt/h
yDEvbGJq1obokvL97UjzUNeRerb8+fIZnqn72dgudztggzxxBZ9HJWFQnQ970uku
/ptfKGjmJ+H4bOzWKi3g2dhAqrXqte82pmOFn8fR+MsPUA6OBTSwmLydysNsF+sL
pUQy6XTm6AFluwk4yJb+GvQEoRc/QwKhVR8pC3jnLowQU1ev4Vd+Keo3hYWKJmAD
aYUOZE+m4TydYSb+T2pN3xrM9CJ5q9mVbQdQi3U9FVXBB1XagS7SjIllIEsW8ADR
XJpr59RWoEq3j+ps3/GB/xYykmUoQi3PeIKJgzHPrX704taDfpQqwED4zwM7/zgk
vgNJKmj0zrK1iD5L9PC9d9A44NwcJ28hGtx7nqvmSkgaFL7B/4Nz56B7TIKXeQIa
DddcPMn0TEhsmObUaAp4CgBtuRwSwkOG5E6LRPchnFEYfuFsMyC4NUApOp9F4OV3
AXu8Bz+pDGBYbINqxOznkaNSuJuGau3BhF2XaMIMcOKYKXAqc60mgRV+Zi3EGqw1
GfpA+bZOP0EIYRflEMSmU7DYYJSomLjh0M5fxICKRtfe4gIfho2fle1cxl9knjSs
uGgCrVLmu5qBdjGqIzTlj5L5+C+n7vkF53hNp/NqIZFef09muHaYvCpk3J7aKK5g
wfDmzjZKjIk/Oq8Uf/3UN/4cBS+1nAD+h108rEMkFfSs8hu4DrnXBtnv2w4ymlq5
DTqIZHNiYVjL9xUqrSP0IjlYPO0lvaSfbXok+T4z5KsUzDxi79bfojZ3cU/im91E
KHexnGxWLRTWUplxHN+6iDyZP2IpFxdq0Uu9ArDCm0zLc93tLLmQewqItF7Kjv2Q
zPcDspiICNvhzCkyOLuem9XEkXI8dNyDU5JcZu/WkONmoGKCAVm5dI9LMg8froBc
Xs9fEIzbxWh2nuDqmHP7wjFpLOVzrDvV9Ue2MZg80DDCdxuSqVmzcjYvjQSvPgT6
2Rlhc5khra0OJsvrrn9YNnLf8Reb8Zm9PMGda9/jCA9G/z/WmwtoT2iYpTG4rNji
f6IXwgQ/5xzpCBZgBAmL02jm04Er70XlRxrFd175/6gG3ymxXzeGL6mO4319nIDL
fGUjU+L8Xjk93CLoRUOHdtYtOriu6RV2lVW0T2h+3kZTFztlJbA9UREnuq7ejxKB
7QZPYgU4DB6e1PWyVGE9lOnBKdAYEHEjc5jd/WhS7FeYsWuu/ZK0TfjTDeuf0mW0
c7iZVPl9rtNc+F229U9O8ykQF7nk2bNdY4LgSzVpr/9oAK9GbPMluUWKXeoRG7GF
/kW+ffxlqFC7nM+NWXZM4+uQ0zDGqkdciw+qS+4oXIdBXj7e2Edu+1oxaG1uW6Gi
A0wxw12jPl0WOMGZw5IBX9VnJjXmx1yNQsW5IQcOPM3CHJI1vEAEQ7Y4lCHOF5G9
gUxN0OP9ih2LDGXXhoKqe8iToLDojD3vnQqW+ghOBJs07/NAeQ6kcolmGPRqGcnQ
R44sgu0Tl89L9CQ094VRmK7yNpF3t3t+QM3gZj08n5/ilFQ3gZGPbscSV1maPBCb
BtZwWu7ZmgIa/xRBiiRVkOhgf4rnCGOdkNX6lCHixi+JBYoaUnS1WtHY0aAX5RXz
t2uOqjQueLAZu4K7JjoCeTXDK3ItNTvEVV6lis1V0OfHCDHVUN4GlNOSH7ZLHKro
TRT4jgxiFHpLdqfDgeZDjgN9AMqnAJqQWs7NwyQ+9Dn+XW3KFpUBqpyOyjNeR3vE
UYR5nKGBtTW+dZXEVgbfNOGfYRCgq7CWNruQprsf4pH4ky7+/VAfWjPzuEbRv6Tg
HNS4y128Iuon6nIOGmi/MqQ7MtiAGawL6jmhJQCMPS+b0GlkykQA/zpcQV5eQsMr
/xP7gQAbb1vqUJh6W17wOP51KLoMX504//3fk2v7/Lm4WNUkJi4hlrEXXABHLFfv
vM3QyVnG+T3OIKJHmHAQ16M3TCaITDtUTP0U639yEobCwWIDbiSqE7/uD/5KRsCA
89NklpnDwy17vjllApjDSyNNW9AmPB3m8kN8kE9kCZ9sPCGMVH0QsuUuqmpMihX/
asqB1i51ZgJWBJ0fSbtWJb7Jx6YYnRZjUGU/EBPoNHb2+tjyaXGIlumAYIunpXfM
bcWlmW4jh33RcUoYtbs8NOlHajfr+V34l9FMUAn8Y3mVJRrWwGVsFB3tRbe0P+3P
I++vGjRb4FGwctx1mH77YKDXjNC4TOz4HFtkA1fp76NyOhhC5TWMKGjmVd4KBTfH
Rw+pnh8xSA47+Mi9nAqPdBkjLW+1fNHdWjroLDoCHfExKTlC+xvr1t74Ajdns2o9
73J/3qIq1rw/Th0Q0T4hBPpRzd/c/1Ds2AzuMIhDkRuPU144mhBZrgck+DiYDYy1
OWE2X8kgN9pWiD3NKnlMMl6wkJG5vbrB3T1AXRJ9FRtOK+fsUxB1cn7tW9g56EZ4
2KzOVa7rMKkHPYvJBvPSpd2KVrcZiKkmHhJnYQuId9iZ1eSM6Xy/fviGMc593npu
z94ndzHbyapgmU0ZE3j79s6Afqr5H4Y8yH74XPzhxqFYXR49M68nibhRk7IBKJvm
18pAGasXVQdRNLU9R9PiDaw8ilTQuUN+KMh1icOfysoWvfC4YO198JyonFgYEwJ2
AAxAgxBnByk9JCPqiHActPHam8YvoQ7jIUH3F+77OIa4WahtgRKlwzaRBsJXbTIC
YCVokCGuh/xZdZcGtWMdHWL5ziE/xHF1F1TpCm4EQ/RsvWKo9DAfv1se1TadwChl
1gtkr9yH/0ht0FUBYCWYuofpLo8lrBB9u4VDc54GpyXOqUPpPY3w9xfiLZbJgWaQ
ADJaEnXoNLKy40g25spi/5MxP02ouEBZ157Itxe3biPokutIbeIqM2Ye/gFrYYZL
yTqbQ4rPoYr4eRhk6lEfslFFmpi+DpTsCE0c+7MAaqXjWLT0iZ2R2DcHi8gvXZzI
dYLuTtxBCi0mxyzlBGoa1oE9tlnSCrcan5EgjDb6ve1hT1X3AoP9iEuEO3/kevP9
LirqNzCYEYPahHxDbh046jV53tJSWsioXDmJF8T0sGH2QuXCx1QG9KPViQjIWFgA
kgaqTRY2GaIg235L6vdX7NqJ8cw8fF9dlbSc8HqEpn3IuGk5US8BVaMELcohhUI2
qw13TnztLLzaGcxDGF42noA1007SRGJZVfZ9qEd3zAT7jaCotgxwbmjXjgEIHJCU
EGMUkimpxEZzrKOG40iUdC7/RIiwNUrkV35ukE4n7k3nUPDm/RgliJKlPfYGRuvZ
Rhkn+52k8TSKdtIQDMp3jpTK7zpebXTR+L3IIZRUuKQluy3oKPY2bXVhiWmSusIr
q0MDW8AAYnrS20TPaa1J9NrFn/Ek5oYAczEJBeWaHd40hXFuXp3tLAfTSdmM3nGQ
tVkvvX9BJP++OkxZOMwUrBe/bLeQodpszZEY+3mD37cfJZhWMNTZudGtHtnqrYml
gGiLRV/weR99otnJ3RMDlFWTHCaQLylG1xjvyIzg0j3m4QOjo3ulZrrBRnntzd+S
ZoJel8iA26ah1OxacCYb3c+2/Ts7RfVo3y/uchxlMeTtzpQaGxczZrDYtHcs0svY
+Va8AMe/Q+zX+Q1dfnCXbguUyctQkUSgSRnU0z3P1rbb0jLSkLBiqBJdC+iqmE/u
r7/WRzQxp16krbeb48jSY9ZnuiqlT/8TTLd3pI8r6RYkefP61Ax8foVQ2WtK8AEf
ydHN6GgIztynBSYIegK9vn54ViZpzhK+Hz2b+Is83mKuf9GcQ6MOm9eb8eYkYPNS
ghb2D8PXU9uSbjzRzqqBjWfAgKAuTtgt/0tqDgFpBb7YqzGCjbjUwzlI6ushCw7v
p8feJQlMNDpWB14xEg7yx/a0V73osdwJ9POipJHw9+0C3rHKDksB8PKwEr8a/PmA
ChEyyGquBfZkl6kFP43N8IkHzr8BxQ2jE8m8P8KErKFEoV0SLJGjYFbZmJB4VmSt
5dSlW5CfmYaMGCTKK5w2rRsNpgLsOPjMH68bNGoW9CLj0kFIpN0NQrjdvu4g9auv
uuRLgykul9LSTu/yKV7KF9b9jdIlznYzTWjm69O7UMBshHCrk2PQyikRGI3um729
tryWWU1qGz3h1TUTAQ3ubLF9dILRCeILR82zk4O/idsx2W0qz0I3nj8yoFalB0NZ
6Cmu6TTsAhPombNaDNBOufOQuhw/2uskg2p4njfRGz0g46LXRYcTYGAKc8Hj/rCR
O/6A1CUiAmlWQ1pN+zp5EpLM11dwxEa8vu381weAzTh1OkggB26HfULM9lnNhbPm
7z1mzKJ8/nd5pG9VcHvm+5SC4RrBbmmLP8EqGjMrMB+UiNdn4p6cv4B71hb5BaU3
Gvp8ucQBkQgnnV1orPYi7MqEjMay0PhO6/C+LSbXJHoMR336YozESDpI9HtOscCs
rXgkCctNhPYPdRXt6c/cp4pvLZVneR94MC9yWpKgNM8uxaLKyUAf3HwX2k5X8nsw
llifYyZ/HlF0R7emj/nyM+UNVAu4+YoIs9O1Fz+a+FQJHG9x5hGRlkiQdSGpOho+
RNIzpzVifyrbU0w1SQcUFr1h2EpzT2gKIYppxg4ZrIfQyBW6K40oKqFD/6LOVcoP
/h5BEr24muy2Zp5iYrKAikSHbQ18Rm6KuFMZ/Nw+OEuCFCfdpqZ/v5d+C70xPVJo
dGw67AIsOBKNfUhBAcTsF0lORRE61NBSRanavCex56FmqwdTTjXcSveVPbnPfBxD
DRmf2L8YSSB2YuwyBwM/rU57xqEFDxgsAq8K3PPGNqf9IVWBQwbCzJpQPQzCp4PM
uU5rGh3Ul8P2qmNg6Yf9N1Dy7gFjaBg+zBhQpYkh6PdgCIfjKFGluQBNdzaKkWkH
Lm3/LB+tQ0SdWCQtYfbsUPXDQuuKvyUZGUqMq287ERNTJXcj4BMC9qjdabrWcVlr
/bVxughPsCdZrU69yWvXIymJVdIDpsxmSJBGP6iFdxz13Q2+cATKo1UU4JNaa6oC
6jN04jrtZ8hu7rPhUJ02klhMLY2Nv4BvGE663q1gx3OSduNdc+YYlIh9rju9OA9j
ymWhsMOI7TvKGeDPc9yyJ3rg6ouGzsnWkVeTgmm3W+9Y2EKVxO8rPmQjDiu32+yd
skbJFpC11f4QYUvol4VpsWUySKbfEBNHvfLn7RUCV93vL8VPdEAdro8EL449UgyO
M2FXINom5kW5vS4NjHIVcCxCZ+9GSMPuIEkfx+iBqzc4fmVANTi9Rn9pMBUTYjdK
iCHc8JLwF0bs5mV7lC3O0EG71sgYhlRKva11Ny2SAyRDunDL6zWdk665JuXlrLBD
Qc+fewqE9NWNOTRmn3YV6rtpM2MjLIVc1RAxT5vsn0zdm5eBVyXhUjkoAL/4q3E/
KBCWp4bgRbl1An7u8Hm+mvRk1n1Ku+vSsT7cuK63Ah0KpOXJ7kqQVyE0YE4VVhYj
U4uXdniQIpGzihY/TlnxeWlmAylXc9d69qLNPsj1UBqp+6eeQpkMzzIWjskSaB75
DmWrdw3zKSB6VyxTVA9JiAoNZ/NI0TDAGSOksUMXjQh1zP8WsCqG9W3juFUv0vnX
LM98tPD0LcZI1HjRZQnQiDGXP+i7nQcNgWdSANwBDgfUf/PdsoxQ3D4gYNhL+Wuu
AKmUlkG1qC8D+Jwj0/xEkSJ7I5orGScpf0WVb7GEOnbt32QXVw7AeKPlwP2cFbAX
MUXI21fdaO/SLKwl2/hDCMnzkElU8Qs96rEqiY6j5B0a1Gp4GlxM4OwMv0+81OKP
lrqcmh7cLd8ftOKYeIL2+7sZW1MP9JDqX0nB9j4pd0qre6U9vrKO+NgiAGT6c4lz
RNasKctFwsUF2Y2/WUaqOdwiirVyzKsGvKgRLGaEpnqL18Kr1n/6pQdYrh7LpX3/
j8uRawznnQGrb3v/spggdziO73G1EgzrApZZLnaZgUUp+P0ceivLhVEyftacOrfp
NzYkyIrA5cFDiS4XAuQHdSGk7hKDfyJBSRJCngA0n9Qtmy+IjDwxE8Ky4kVP8noX
Lsci773Foxjm6CTDM6/59RGA/TePRDA+hqOYFVg2V/nUgAA7FrdfQSfhmhiVPLH0
DohRy8hYYRN837CdrGI6oRQBS/qSGP4wVutiR/JMII59pH/8BXRT1zUIp2ZP6Uja
mzDxwcBj1HsxhyYJV7Lp4E3qAoU5i9hij2LVt/fQZBw637/hiVgX5aE40XQ80rAH
enduCqJjkwyHOAbPBr2lFh7nrLURM9ncHnPmY/W1U54vNaeg4ti3nW0dtW/gl82Z
LycVOPdgGbvn3+tHmIjM8wWUG9TojKAfSGzgktoLxySQKTS85GnHJtKUANLLi+5I
Lo6H3uD5D7alAIZachv0K9WHiuvc+eyfXaLhI/WndyE8GNFELI8jao4KkaECgkOR
MyCYDBfuDQ6u4ZF/kgYxhZHUjLKIyc89xzp2KFeOIhQ3ScuD0NIyt8J0NAWU313f
PDXSyL73nlmtIT05Qb6d/oZarbmUxsPkgdwVXrF1biK9fi8ZsP5PfiJMK1QQx3FS
s+60V8O9eV5HfjMLW/pzlUXxjmveAPZr4S4dKx5FfMamHP3StvCqJUHXrXNkzRrn
uJ0Ptt7aMiO9nMa5NDp/tSruL+kFumYN1w0iMo5Hk2ykjrWaDT2XFHfTePq4BIkt
AHFtx9tdjFeXsGQVvI1LfghUw+ljILwehYSF1j/amaR9SjvzQIVaEcO3RZDjS7gC
psAaUXqbTRzGfoBlNgBI1O/GrhUvNiRD2nGuZczN9ljkMaV11VyyFCXYnaT3QV8k
KeRw1cIp0DOleygMhasNjozPi1iaPkObe6lQi5MwY0yQs4uOEXK50I5WXeA8O2Ao
+BqufL1SmJ6NN8B+45zqNLWwHf2oNT9dpZs+b4WJkSbaK9yWu8MldbhW3TqusmIC
fnipMtJPURExm/EzO1iqhOmDd4EgqGlBumudgVzprFUMqBwCugVHLiMd5XTNCy7n
ZeHYtzp8dibHQ0z/0MnRYrriEx1WFR1LNfqnpTz3ooL/keXZxV7OxBKeiszYFf2s
l3u9m83jYT/wRQPOyA4SN4LhK/2s2vzUQN4ovh/FtXfkCMM+844rcRTOq7ngZfPf
09mFgNvCU3HcaJHvFVNWhPazHrkifFjC0QALit8TF7jWQHnAhDL3IqMo1XWtQ4DW
lPU4aKAsN1/vYhESWE/zuB+Q26r3OUzVfFxy89LIFU3tkWQKHYTQhx/um9Rc30kR
2nSuHIfP0CArHK/pAqo84pNnqXo/tjEqdEQe8pIuF/ixb/YnM++t+ePil5nYq85Z
F20FOcJG7sz8RvarlH/FvslVO7pN96Eh0iOmxqreUQS1GpB4LQkK8XTAfgpFJvO2
jygYI5QA/yuQvL8hF63b4oTyoCu7EZLXXoTvfn3iuf7bGAIeOo1lrRZtAhUxIb3S
NAdKPWzShWsb6UruqFJ+rS7GqWaRW4Q4v3r8YsD/ENagXVaPiY1XnSwqs8Ky62LD
pizxAGk10fv/Y7K2xQcPPEJl/jd3yQSu4ZSA/2oT2hiAQcYjnC+4cyDCFSt7tEXz
SNECPYJUEgWlaWlA8dQfwCgEoJLANJm8rwR1VUT2BTHPMQqIbfBRKohIP1iH1qmy
xYABdq3U3k+dGxePC6DEtTuRsi8oVIs4EoxcL3NutYpLzo/vmOFQuq3fpg9sF26F
uo5KVhZonKodmLVMNI7AZCI6HWgIHlaJRT4DkbbtS9g+qkvbpHkY8O16J5Jc8u0T
gMTglvfL84mV4QXp61AXcgQy8y6eoMfbRYBZh3yi2XFlXiGnOwVMI68x0BobIXK4
N20JSdUm3PttRl+L8fhL6vUa0IrWTUoNzd9BcWmYr2ek9zjp36rXEs/C3SrFL9PX
RATzJc3cQo63SCEeNDi6kqVCBGOvGxZUpCCZHZm/qwbu/xnTCR7zmQ1FrzH2NMh1
PnoYNzRytZSXakbq3FwFcBb76s3oh+MnQrWJYyV86VbfaJJbsiNZLIB401CpsCuQ
IDtyblCzonVPk4DK1cYdd9oHZ1HND2cr/FGtMdXlikwIMGXCIb4CSouSYISxqlZa
ip3XOrkHgeAbunGtGBTq6hHTE4iuUeBLyGEo/Ygsp+LubnjH11SXSr0nxm7nXicp
L0Kbik2NDVBuxwcWdxqMYSSvKH3DBws1awcQmRB0tH4ucdUabGqLYdTZ/k4NzsVf
XqNBw532LTVWrzf35iTntfxSEuo7TuNQmlefgYs5Iw69nLlH+DdFItzYJ3VLblGd
a2DD0NIH/8u7r431AQN2VXFI2hF03zZmvUb9trPrvGkb50v50YAhbB7zVEYEKDOW
1pBfkj14KP7up/9BDl6b2AV6zTs6Ci4E6X7jzYdprIXn332La3Si7TktcrqvBz/O
s6IhabHgZtekNfqgCZTSqAi4Zi5UO4IDTnL94fYdOILOvopUwcZTt8aDS77W+t28
OdXogo2mWghfwzeyGKcYnU0WMtxME3iMoIU0KK+JnJ6WU9UQtH6fIohPF2OnETn0
ahUPUuakpbkD0GxS13KWdfOWj0d4uSUSjoqSDmmomSnDDvMJS9GR27xsMVhxPR8J
OQA60YxLgzUZ29ukLFNNCXf9+SSiYr8FLJbHvfEegvSuKfikuYdXwKx3t1heVVhX
ywDPs3sncKV7g5Km+4CWcR8VsMSnxwV6QSR+VdRooCacFnqcN4x5+8XDyepXQC7v
nkPjAZ+TZ7c1FW9rIH+1JUEVtkk4A5s7HQ/Y6EHkraFFXHM2btbR+fl+XOTa2szq
RvAIKYlcsNfkJyk7942yF0xFNOUOcZ8JCJgIuZMVE4Nq1pEOlM4O8Gl85W3Q9l5m
Wtt/fhoW9USgAAFpCA6ePXGMpaDaBLW9r1w4m1YOxgbmzPCqRvaTPCDN8pKv/rNl
7zXMQ3mi6ZaSrvzOvXF4gkmHfSBEdF3ta73h/nBXmplXs/r5XqYQw4P47Qi2qUVP
4fJMfGptm808UEE4nf1aVjkmzYvZBv08usKNALrNqpmvoNYevTR4iusUbl4uTqrn
9BE6sdBkjrkzhu2m6pY6ohTJ5CtcvGp6yn8K6zi1jZaOlsYvLMEds+AsxZTbHdNA
+GvITdHmQtjEZJnCjK2nE/NBgHhW2VIR7d/i6WMFHsnJyNLQYQ1A4r7CmHmXuW0Q
HDlC5BLsMQRalxchoDkbLL/6W7rqJcbnEBYOqNQMSfdfqyugqXFw9sbdIxI0IXGh
zQ2r8m/qxHToshghdn0Q5+lM05J/YMN1/AsOlbkulwGyXm3YvUiDVzxWMeQsOeoC
46rpg7EEq/yfov6w1V/qJz2xiDeEZ5aPOWIPhxVFlWcyLtAY/6XNek9rGLzYdUrj
F2T9RcbI6r0/ZxrdQapuS4O34VtlV2cSV/ESnroSEaDD7JCZDJUUBvDUWyFdot9s
GXeElULvzDdkGFMwM3eLBqCq0LCSLTyflwhUvjIAw5lLmGocFkwOQTOreq53NvJK
uoF4/9l4i8xz61Qa3bZncvP4fazGH0dKUtsAjEF4ks7I6IcQsSaKKAHmwSFsfVN1
5Pww3FrFS6qDeHvkLT9gTKy+JSgJjtfazMxXkcw6wD/MYsmlv5PusqtUEpI2INM+
Uy045B+8Kky4KvXfFqcMwpMoekwiPcA5f+qTXSuH+VmDd3Pkx37gS6vNZpAixrIE
dW7uUmLGhkUEZRFM+i5C/+DOVFmWgbY7LFYu4bT4/eYRphLBbfQhSaK4XySR7XPg
kmjumfYoQcr32ALa62CNVyQ0kP5429QhfV5rokYKeEqIfTpAtyvmNsxLu/b5UEbT
ltoTw+DPtUcwPCxVGktvUDMoBKt3h43tvJJ92R7sgfdhCsnDLA+O5dtqCNdOjNHd
0lUNav468TnMGtK6B2QsdRQzp66Rx9Fo9i4bcw3L6h9UxPhJ3UXi9h2K6KMHbEh2
SEAXCBW8xY3tpyRafE1UZCDWBxMeRcO1FD8MKDR6ur5zH7BD+U629J64t7tn7Lxr
XMTcwz1uwERL8sWLRkgQPIoaUWlY9P2l731VI0vsunuB69E31haNXgG7VPTYktou
XlPeEZCeJMjgLjC+1JwSascU7NjeaTSMulNc81J/cCpM30IV2syxWViJJKvShvFP
P0p/20GLsbM6DGXv5uKGUDpK/5ByVx+3CGGtM9H1FDfhFUhOQo9uzCjePxyNPFYV
fYotE5ZDjXc7xVi7+utvjG4ErFd69xwI/+NSHOAX3sCGtTt3KhJwzAJf4CrhAjPK
XwzaegI07sWBZyrnZAneQUMc56glLRBAkw3/Dxbn2oE/N9XjAQqBTk6f/1aN2k79
C/C1/F6O6waZUnR9xmaLBKRNwEL1G/I5YO+wX+RmnplQ2zRz8nAQ1AZgWvFdAp5i
YGNgEBhEdSMgFWrB6UgTEDifM8f6HlxTuDh0+qSvNc6Ge9xwVT+qPSTAhqmN5/eT
veQk3rzShEIrin+9Fuhi3oGoXjsCqH+IkjAWBKG2Q+emjT74M3wkl329VTZv9Oa2
lQEOSKYEBpvC5ySBPOfGGQ2+vf4QQwT8bkTz2vXsQpZGOTefiDmKEE3mb5LQOmkK
coyBypkzlJNswMFDgQ5eUrew1lE05XBlGPkRspPgxvs6c7FqXMLf0gnDdPxCiQQn
kN4S7UL6hlEzbDeQKWlsv0ejxaI2/iH93MkKli4pnxYjZ6/ftPEJnv2uuQ5C2Csn
7jqr63LUye3fENalv2TTbwIeolpjVZwfaMq2YE2YwVHhz1/SdQ43zBpo2XSwEkT8
93WN913f9uMM9y5/gQK0z0DQciUwiV9pCgDFcaPW7U+6euuzLv4JY0C74ieCT29Z
k8Fg96IVDhg0IZ7vBX5xX+oqfs/ayeQh+fu8EY6JtPFdbkirj+BGBOXRrdx01lHE
3kYplHcJTVFyuJT1VSeT3ZykuK49mKv/zhJ/cVzI4jenb+UNAKRKB2euWh24NQF+
bj5YVtmXVzrnX7jVjy+4ItNt5h9jqVTmFu6jd7i6Bf+eRMoyTgYJzKLWAcFndLfB
o6SfwDKSLCsiVM5N1GbafveZOv+ebKsvXo1rv/hQq7q+0UXZX8SEWrot57oM0utk
0qzSoH9/wuIVHZxUbbD8MojwLYSuqq1UjVQ2+nTJkAwH29j+hDHU4kPld9mtIHhH
NfYJG+u4ErgvurDG8CmAN//XeDDMYOxHDPtlwQ5mBojv2E+yF098EezU7tIvGlhS
saaLkcwXf4Kt820eeuOlirRxq8teThSzMp+2LNLaaxTBcHinR99I+QSt6OasWipP
NAuPsGvsVuJxwh9mAAJFCEA5JJLWfbnDEUAt5ld+Mgmh43zz7d1mOxXnMqp7ZNic
xGrLV3Gi9DkAo4XgsGKJI9ST2O6N1zJdi3lVS84OZlbn3yMQpdczaUnC9vZH2huH
Oca9z00dZ/fbWEuyaxsQlLN2CouPGn3YU5p3njQLtzwkFvpgXikJxqUfTfc/1a7b
hOng1xWcENRXhgS9wgTuIDP+rP9wqeV02QJ/Uby1FOTh8o6AtHnXHw7gkmyC8Lyd
X0rmGAGTH9+hWUpoFXXbdAaShEEa5afAPPuY/dZrydP4Cux4Q9VPnPSKCy3TJdm9
EvPFkEo1/bss6sm16Mz0X3MJMUfefVou49eLVHcaZv9DJxH41FMkeJm+ru18BMP7
FVRtbA0mbnnQ67anJYvsXXhO9wiKWEo8xlq3Mf6XOa8+6Swm6W3te0l+p6jEodGZ
qtmvrHx3AbYOMhUSnHhKFid+Ee0cGzsx7qpr/42m+2FXqmESoRLTnNz8QDN3m+pg
GUzlOYx75c4q+7Os7lYxVTJRFtHwJCRolUm08A4b3ziM9ZthBlmTdxftDXF5et2a
LmnOtBxqyp7dLDHg14wrHR5pRHLQWFS+X2xclKVJwK1aP+jxBvBNucA7OcuEDfUd
Q6he1T1mgFLheae5HSXFk4Tsnymz6nnqYktMl3uPYDQAyB5KmXP6AF3qGTZIADsm
NZ7mBTB4e78mGlvLodWIB26tcoDXlfMgKvHUIMJOabsjleoBMNTtd7lAnwtEI3Us
EK7Fxuk5pXhU04lkXzQqFfwynLAjBYxhkvLNu6Oo7+nZLbF7GlKbciNvA9nv5hQ0
MFCdk4kkgOheU/YS3b04WxIG+4Yx9IjDfQuhBQ+y97vhqoku2LNCgxjYoIDF4/N9
G5+sTZThLA78prBI1FDgdLLgQR9L4h8sZ7/H6SNWBJ8sOQi0pYiko6jaXtreujdi
4mxO9ed2i+qeIXNl79nBi4zqhVdK6XYaKZaiGxc1vJFeSqJocAEINcXq0cG4QGVU
y1aW3LWVgSm73F8utBccBKoWySnIGAvBW+68D1kx2ENmcfW/gPcXvaptOmxh+jFG
WlOKmJjaiv7PVWzMuPlqZPOGj6xGbr/lejuXBLRQb0eJ/t7nPiJ+ctqWl4w3b2jl
4UsY3pR00Jjxx+4BSHaPDshucc+jXMY2wPa7ipJXYAYcxIS4mgPxealcGBXDhwlS
5VkYZkG2yNCMAuJN9bapVAxwSvw3mXL5AE/cNlowj9rFHf6QWLA2Eg87YbjnwxUP
XSYul88jECL45vmdwu7M9aoHkxZRzuY1MfUSvKr9A6amyWX8I1/7sTGnPRSeoKjj
maNHSbz8h7mG5BVA8glihtNVURlZqTthpbu6byeCsFull/BWX908gG2Bfe7be+eG
duijp2F5B460oAIbqNCJ94nKUsAr5kOT4T8ihJLpCDHVTGeEvnhhtRggwykgk6oV
SrHX+JY77y4/yuSBRgQ04LEQRXDYQVc+p5Q0x6Z+KXepazeBqqwKc3d2Z391G9kb
JpwByGBSE9OuSrPJ/IiIf+OoI99Wq9pp6hsfeaHCW2YVbqYhcoFK29X0RZD/GBzX
lyxBbqcLFkcG1HR61y5rV0JAjHaExcRjAk5UFYXeURgeaj3UgzuuUCuu4NSYZG1D
TrkV4X479f4Kqd/hhOb2gmeg5MKTyFKEZrwVw1rOSTkrHqfa4Kkw1nzpzyfTI1jC
HFxe82z6AhRc2iHMUaN2W3WA52Vx6q60D4PtnqzVN3fyRaPeWBAYb7fCWSZePUYV
Luj5x6eDd9WCQDlXjfFQQlf7Vu7Wkda2lHrA5WweWITDWWJfY8QUaIi/Mzhtmm8z
RGT8NzO1yQju5LE18n1w7kttNpAJQSSxGGgP3c+plsG5KVSwDRmFFa8MwGOR7sJF
GvfESOAoEtcnD7zSj7pliJKO8qKfYigkxge1d6PFWhad5r5yllIhdM6LAhtOBfUq
haq8ykNYs2rl6s8She2U0Z4/BTOH35PAMdKc/rsX9gzYfmZmETkAq9+DBEmqcyR6
JO7wGUjiaI2gpqrkJHJe77r460HRc6yNw7wbySKdeaFd/2vJ2MrweCOM5BupJSjC
yFysyq7j58ZIulY9CKkEoA9hED3LcBXhXrOeObr2bqmv1nY0UECCpnpN8mhd2JVJ
+Gjx8qZyk2ztRrctWcCZdmwuS9j/25d1mz5gVQnDvv/38ZWODhlkpfW3fduD8vBk
edWeDCRw71eMHW16xSXL75lMso+EBh4zRGJyJToyqI+V2H5niSl3g+/D9H9qymkU
YuNtjqFZoaULItDHDoVCj9MXvrPbgySlVNlhGZ1xcFCQD2f1N2fMeHct8NNT0zOA
pWU/OQChzyz8huNfzML7UamX5dXiFprYc+uNxzhwzI8YJCTCFMvDhx48+sjKqPGN
6yBUTH9tG15ZWnAnZ42djUpi2oH9RJXP/E5Z1EpMFutAMHJi+pTBWqmC7Wa/ySZR
/ZUzCKAQKNThb63Lu9ptkJPexHVIEwyWk4xxxImCa6Il+SdgwR2LTpQ6iXsRRQ4m
abHk1C3vkv7WqEJrPHHprjA7Buy92Qg3EtWo7RHEGmAS8bsYuq09pW/1taOvr1hO
rfwxNDAsq10U/2hjIeEQihcbBivQ49DEEJkHd94S7r5ZQGz/QdX9IKUu3gXVhZHb
di/QVHg52fR3RZb0fp3/a1kYLEUI8/PFZjIhBaH6a9gQWgGyTGSmmNymDixIMKMt
l1a8CGm3lVyh6MFGH5h0FXHgtrzDAh2sGIy6oBLrzahucS+RF5XIGB5zcA3rZlvx
jLzi+0Jr3JjOySDHxgnmsDwfrmUfXtU7Ka2mbgiZ3lzuGmYPWwgB30KNxmAK33Um
q9xju99ZEiAxKMnP2fGgspC6w0CMfKe1E/LdYv2rmwjuF5n78e/j0GQ0fg7US9dE
IztFI91XEuVHawGMbl2N8i1cY0z/6WF3iv88NmUWrz5uoy+EjTAIx2jqjSNVHgz2
dawSAsFm1X4T2nuGwnx/DsAwmRWlD49gS6QwzG1cZTC3Hm7IrHa/T9hpLkw7eZJN
saY2492oR3N4O8yLP9tVodgL2Ky0XK0ijJ9rNNPYg7XCg352ChRuhZcfjySTpSMh
EO80moDaC7GHNLjdMCLbEURffI5HzJann8xKzEU5gkSJ64mKihTsTpyj3HgmJEo2
x2P4IRhvftkIWWMRbGMNg7jjrrchkc/xwOhrezhSRogB++JzfOKyF79oV5Zksq+D
HU/1/uat4cMvJzrMc3rs8CVjNex1nfXSQAYvPJzIRoa+3VviH259STbTUyAnxN/B
tMkvOVxJyO9eUeFTY8FrkP/Km1kDbGHw62r0XStbffIeoatrNBM8MFqYHqiDAf79
hYfxVV4FmrOMQDxtdnWPQffha0tPGz2fLRes7LhUuNuDfA97bFDn1+erhB1vGurD
CErBAkDhXTLmH97DjWPfZ2wHOwe4yb5phlXXmH9NBRqVHGTf59ICxQP3i8o1ui4u
AIcmYXXK30p8jYbIIGX7JfzADATduchsYUiQ+A3TSi8guNFV6OO+hTGD2vRI2Po8
OP71oEDLDF/uKhIF4mH9agF/veJTbRlyvJcKX1Cns42psYZs1LvmVBUlFD0q7Lv0
TdRYRTL9bU+cfeaNEEcrl94MIp2uHMJhOfX+KQypXhACg6oKvNBv4KqjDFV+y4DJ
7fhzW2/w9bjpw2ivyAP12ZSxxlTbbw3TDdsP8fa6YVZ1J6qj5Xf0DNOUfxb62yj0
CRlI9E1gmo2ZMuOpVnA9mbjOt8JhPNgPJMjtzquP4cKpDIgU1iua6yi2WUlKXlbU
Bspjk02d4Cq0s2yEhrIQEV8gblqF6xhKo3ouS8sPv8iF0BjREYa7BymivZCON8BJ
YoEdAK/rxb6Wjr41QwiDasALeEYQD4azJaQBq1tyluM4kVai7Z+Yk8k5crh56PkP
bhL6M+lINsqPhSza3WUqjOCrDulirca7W+vJwNnAtTUT3/Xkb6RUR7M7LnN4/jdX
T/+k3hKR/04DFPDxqQdvEXD/IGaeRmu+tKpb1ilk+BUMX1HRE6FZWTC1UI0mf+l+
eO+iUu17wgDG+2A3mnCyZQVq82RcCVJrvv8Y5auYxQhrMMtvoezHy7jcIKY5ZZnb
xG6tlyQJlY23+mWoUWUo2Z2t9TKtgIt8lH0BGChdSr+DslqqT5FLZWTtfVUCr6Yu
kdn4zqED/cHdh+tRQuXzEBsWfTX/5zCIKaenjxvHd/dvGujux3M7T9a8zeX+p07C
65JkqyLDppS2k2/psgMEdtY24goHRMnFAYGrWmxyuvWI/8lPkRgEvn3qLKnoOEBq
tDFlU2c1lMoE8jRu6dcRHd61XwY71gdPBNNX1z5W//KDYVehVHjeTpcDrRjT38X1
cs6DCrEdGUjnUjZf9US/G4bSmljdhPiKF0n6e+lqv/hx8GT8S7RuofaEHJ/5LVk/
SPzarTCeJd/vgt2vSA68PK0BQ7Hq2M8tlJsdPIcIOD6t9jzRfdRhNJ/X4ODyCZha
0JqrETOPUoBRnD/jx2Sq6OsYpKu8UBKbZ6GWuorrXdrNz24Qwk5i2qj57PSnYcu2
TdVf7ADGRO8kEKaOJIrIr8dKjBQqO3wueBLhnmvPhsGvAkzoFcxEqoZx9rIern2t
i/Op+323W+et0S1499NiyFHXqyun7CecvY8EKCXowuumoGiflR6pDbU7vKAG3wjA
qU64yASA9P+0yJAS7iqRdFMnWRrbhCa7I1SJ3i9RNPkvKx+saZOtmA9J7JtxsA8b
OzsEAzPzefjjsS0ECIqMk/l59El9rK4ieN2Aq4zWxf0IXSMTB8JsP2MKq7lwbry1
nvpBlE8DjU0vnBawU8Ctxh+W416MiIhaEbpvw15dDTyiG9YQTym904GxhYvNdhcl
s8cWkUYuUYkjfnPBLioZMJTM9jZWJqodpcMTGK7o5at36b3gQJtXbfzyI8RnbX6D
gbUAbG2U+mfJ/W2XjTHnnMnhltWPU2YkOMtUzqNOir7kWrBQ47K7WTRDqNB4Yj+p
2GOjGVY+bkknhF9h1DGOPd4RWeI2+iqMWkNyzQ5j6VjgWHNTn4eDzWmWpYYyG+ji
BXGAqkAL2xe5o9DpfeeghGZ9PBreHdhNhvMkynMwxTbfCdnBbbmHGngGGXfRgtqN
aaE/JmnsHe7l0HAkNZ4t4RfWeHySlbmpiyW6Y2m3aZW8QguBd6n4Y3m9tjfgX8xO
GGdl/Ox/4cgnzDCYxLzmLVWWBpETwcwH+DpVRNztrbQzR9+tC8ECI9NKZJRLmSvr
5xLMFeZZpsmSTqOJRElQiaFN1cCwUKsh5nztta0u87RnYXE2DU8d0B2HlC6bjR09
se9AExvT34/QRJhkP1kh/ZVLua1+x5F6mEfWVf5+wHJh89xT5Sc2Jxb9nSjawytt
5YFOj+SBjWL1rpDCQR8SDzZwl3drYQbEYGx0ggh+3riUSVLpSWTiOsnLQx3k83WQ
WkuCYEzHxM8hAmcjHrCmdqaWFpFnizpxGLI2guHmGeSAubFcv5dqKFdRQh0H9Klf
vaLwJdWmLbmvJmgEGhs2ryijdPHJz4NfqM9SOZKYCGZU9SW7kkyYOFRadWM55Qhe
VshvDTKcclA/R59h2NVdT/JKK5bO+pWAb6Sn5WE/q2f4UkmPVE0kAiiZi+Zld02j
hzURbeojeuwbWh2lSeCV1AF8oXCiqYitB8EfS6kAO5zOSL4TTtSWIHQa/t+lelE/
YS6chdhZ5rGOZhdJxLk5jtqsFj+gMr9J7iaUS5ZFQFrJLKNqoAnAxogGANvjG5Dp
FUkUIYxY9H7MYWQWiwqvaoduwbtQG+0cjpz+ZTqIETnDKEuaUfE+xXfj3TfIPBoM
iwF5D82oJZVBUhYlwfyeapPiAonD5A/dwOcSRW+LDHvqftD/ou91ZQvYkPmZ3a8i
Edc9SuDvudeInye+K8LMfO1Az1t74EZXgKhjlR7p7yJVBy8xr3SKE/3pVVv4hxqr
/95wrHev1Whji6NnqR7ljDldWq1/LmzG0mAjPYnm4+fHjNQcjKRJ7wsBNXEZTAHR
JCNOHxg2OQt4ksZ+LwcKBh1c5jBPVSjpg/9HVgibzm1Vl/o9JUBQhdvWFLFQAJjj
PlhWwyTWe7EmpUPtzwtPF9JJzAuSy1WqmLAzCBu9L4zMh7GPMBHb3USJ1+S18FR4
qMm09ECWQarXx3nBO2v0IJMdwUUUvkIzMC1WT1wqt5fqlMyqK8+M/1oxajIAfDrG
sfv9+nlCYFFkzdTdio+tgK6ekQ9cRxn66JaW1XG2RLsDw4YaxOpHqBOU1rNbjYB1
qkj87fU9yPPE0jtDXY0NcmxbBIpRDVT7J+K0F4QrUwyNYjKpmpedApTMxxUtZeDF
KXNsitAo/+n/RMfTZ+pkiVG5GDSR4k5jcamjGDSAtOcLE1EREktb0EmyE1+fxKQ7
wSLti3wzGf2pdIom6VqGdeIkE/K02qYAGY+8mo/GbWwR1x/vH5MkO1fNzDdLAmgC
Ov+eWQq1Y07yAy7CD8iamdpZUCPjW6fOo9jEqNX430G+UFIa5TiXRPTcQxL1vtHX
dN/IFGCTVc7t/+72cAj8ze7VJnaIHC4wCVW3JKdMkPZO5CcHxohANhJ9med6jleN
RR/Bc3EjLCSq3I96N+9Jk0I5uUtdLljCBvIcjSJ5g2Na+As/0BvYrA5Ehqtg2SeT
JgYwQLhGXfY46mVHIbLCLTVhKbbGI/8WTYLQR2vPY7NEFWtMsFTY9NgEo+5R5Yjk
Txxrb9b8ZHkGY32TNyBe39PKSyBn1ZEygUbYiviIK9MuXAFB5lvUVSRbDGl02yHb
0poqQ+eVjlelgetQ0wf6AQrTBL8ELhGO6eTC7CqsDGGHzvhjd9Z0hGyJkwk/1QIe
PVJkib6433g+HsS4XkOPavOZ6heJOrwWSmqBoDMAgc4oHIQ9DvMiK49erCOCr2NG
B83EdNl3/eSzkQppqZNQDnKWiNDNjH7C1AkumLQSj+htlOkdFMJRT3UhRppP5k2p
bPQSNJsx4L10eMrR+KVFXmyh98EjxaRHEy5e1wT73E7gm20qTOuP9W6Ig50F5XRj
jz7IdjTYvzbgI7ahBbxu+Zh92gT0J0k3HoV0mpLWnb6naonquf5xj6SLmWBv9uRw
Xao8ApUeD1BTAm+Yw/8X1hSGSXoFiuwRyhvWZ5PTDYiNgYTH3wXujJWZpQs1Rk/K
tVWRxtCC1Y5pPvtCXKutayC+ipg6BfNwD5UOmiFUca2+nb9vk/hVjMteXlynh/oU
H1zFKJfKxQrlV8NOCdizMXvYU8GRo+JMOVF2uZcySSrGkBKtWDuYeqPF63LagAYu
+xqnOYqpcAVZaj9gNOG5w/2UxF1Q7Ze4YZeEEpIAKkOFkMR0ezIXco5F+/2KjcIX
rnuRvCI17LH0PkRaayHNfyYbLORlBDeFcICBOsh+ZcXymC2h7yrl54U1zZjAHtEx
Io1wZ+iT9F22+4ywatDBSNZHPonzCU43HzAULZjRnANk/oevqMj9K3ifloRZAcUu
hhCPgn8GjzqvP/ZXzByANlnSXf7lp2emwlxeTULT46hzTjLZdGN+FazBJPtSM+3j
ZE60GDLOhu2BnucNQuOjNJBc6gUIs/BiukGAJNejIpDtiUjfQ/zcshZfwwaoFm/8
hUE7lR0XvWYVgltfDv0cMZ0AnfTGobnj+7F2ud2Og56dCM4JemTuPJE6GMhYo7M3
yg3V/3NuPX/TeJ1kcfOCLDKN45jYfhOf8nTpV/AzYGeVea6hXJGya0LMIPOEYxTE
RqfToo+0S+2gK4APkQNJOrlIcipmHUXWt8HgPiUK6DIeGrwJNupU8N7M6sorHOve
EA0mSAPJibXFRXmFoQtEXzjaYnW7REYt26ARf88iZFn8SxkRtktVhnJqAteHi+rz
E8/RPzHUNJHr8OGT4/g5A7EfjYsJHT0MYY0IMwmALMzAY4HR8e15bBAwJOgYNDfC
bbMlVBf91cweD3cLJ8861CGwNw8og+XNh6NfGUt7FX80PrK5GwB3Jlg9LO3mdth3
aJEB6O1RiZuFmQzlE3C8+Dok2X7MkwPrUH8KOPDbby5DG8m5kSOkEuaAczTxW6o+
cnN+Mxok1lKLIN4Sk/zySS/va72dQFVJaMSeqTIizRTsDvV9WkjDXI+ilKt7k6is
78WQ7LGUDZDo748HhoTO0opOxZIx6v1PupLIgq3H8q6z5dZBAHuZioqK8OXngGbz
F3Cus+Evshvg/ucubwvyeBqUJFKbT+2rdsvioz7nT1GLaf5SjZqFeRiN8U807ZMo
iLnz0IjzLl2rJyfBfrrUz97mKvfGDHZPV1CJyOMNnxuC288bmDsCA+asyqChG9aD
QMR1TfDxyv5jsxUcworpnoykVepu+4koglcvNYzxlDB6rp3t2lzfLFApcQEafu/2
IsGM86pkozzb0uVw1cs5fpYBaLdm/5G1xnNJtkNMmWo3slLklf/q44kUGCgOFc47
n2K6Mi0QhypY+gi861ikaryWSi0oqUpWB2JqLW0BcdqvJs0du85lJ0bnm2jmmb6Y
pPNf/pephh7pSfJfT6c9gRejy1eG3Xut5AN+5arWBMFDNnNHlfxDshnCYf6+tIH5
l4TfzMX716o3n7vX3Nds8jX6jcb36rn8QeLit3sW75+5+DVB7RFVp625b28HF1N6
1nnC3wKfy2AwUyRwY+E4zbzH2l9oRXp2p1unBgYdpn2K9/0L7IEhgs/wRVlYnahW
G6VSZTlSpU6fk4lbzcqaVZ9f4IpwPGfqsD65MLyv53wVIddAcbtite/uRkzkoPVv
2h1pG/0jP03BbJ53wYpicpXGoNyEgdMcHrMghX+4Eee1WDnXDoeDd/lqTm7tupGm
DyPpHad11hognFZi/SqBH+pEYEaIbR/kYIp42EbC16qJSC5DE20Kzy1fa0xuYQlw
by5USbJEIYBdSLSwU2UPYjJxgrjmKFpDHOf26uqFsyyIq2ce/Jt1sfbE62rQWaZ4
llv0+dgpxU7tjAs2GFm1TQ1M8cZ/DU3fgA0fuluGIjAoE16m7p+SuURgFd/Q79ny
MpTNqLtrO6XJ44bZJj1sjZSigyfW30tXZqaGXXJPQJiwLQteHH2U6Hg2Y3qSPiHt
tkdIoxWiTqxNkcPV3t9OlMiyxv1ljf5SotnvzQZTMx8LM22M+P9A/7zGPLiIiUQp
CLPhdBC+KztBqYHGqqgB0BFUPP7VymrgfSUQ26OvgBedqe2koIrwFqe9DVaixRYv
9ITSqRu76Dn8AuaD52EWg50nmTKgjvCEPTgV6ZiT9rjH+RsfZ5cRoWRskMeJEkgm
Jy2y4i2zJL93NIxy4PqoH3vAceQs7DexM8xxFXeEV0bdYf0921IUHXiM8wiQ8oRO
QwEq0kdGBQl8+mNmZpaIh8TaiVUpKnuBOKXeUShQzSvbsVGQy8FWdh8s7d00JMTt
XHU6V5nR9YMpxEcyWgZA2FMocEe7SUcwiD06RW2cHW/Z3R9sUX7WhPeLDjDz2S3n
M5VfZWDIjYSQVEBgov1GN3/4of6VFPr6V365CzZiWpnfc9BsuNXaXF7ibri4bdYR
yJyMmlZSlUCAxwOZ43ESD4ZHGmNgX/o8so6I6uAZ+/1I7ws9T6qIn8UiGuEgMa53
j8PiHMe6i+1VnqWYWGBhCs6vGU3nAcQPA+/aS4kyjg+vtKz1Na4YOrx9soBG0GEz
ygqMAZzvfEwDGSbSpRw2w495Mf0+2bOr9ACnizC8XVg2668w4DtUCoyKRQP5piwg
RXgf565VI3oh1+OE5GdDLP8ikWz91iNJd78DbXNbnGZVXOcYfFBsuymunJn/GgM/
EVUAgpxZU4AG3yQEgJ/9u+tpJI4/ItZSCag0QmqHYT0s/XqmmsgQNyerUDO0jLLD
y9yKYMNE9z1IcNyjWyzQM7dOjg7cq3/XB+n2AHwHYIl4tde5Gl21gqA/B+oPlqQl
FgSbOtSQhD8fF5EDalRFQ1gUby9v/5MwknasaWeSk64vEGnGBkGh/fONXAMOy32M
Zw2rLWoyRMyyVpSJipNqbI6WGR93XgZG0icpfCFxOWumVVHs/ebClYvHfi1SZY0D
EvD+WqT4PF7OvijBiHILK+5vCFm2HQaDval/eSbCQF2X3HYLaLVGz6waXD5T12Xd
rGZZxG+JCYBqPGm+b84IDEwq6ha1B09gdw0ep7IpphTqewqOuQ65SEPDDffXBQrQ
UCuVJdgXTVR4cGDVTYK04BmOooqDPEYdB49Oei1JnW9HZJTgsIYAQ5HsAHx0tUFv
M/pH6p8AVhZH3k9yzQZxXn07tbs5el+pHBWGkKuBPrtOSOhifJn/TJoCZaUTGNkT
Z1A93yuECiyDFoquvABARJhPjfRjTa2FvM5OW2R4aAvJRkGOG7ep/PHjYCRVIZfP
HeHuZWTNMnFtF6nq7RJTTFW1rWcst7O2rkF5RDrI3Xk7JyGyCiMGZvQPYlmAMeaE
eyjGvuuM99xfL5FLy9ZvWYK3BZtklCx+hk13DpZOc5R81WNoDUeVPtRfqqhL7H7Y
zAl3iPZxhwT5L5ywlFsxBy+hvI5zdqI6rwAErVElmBji2dOVxGX1asysJDfKGdJT
IwfhmlRvshxu/Gd6BV7Ek+AhNKvODUWd0RQ6ghR0hD4DKIMgCHvt4fT6mpM9zsnA
yePakWIQtssK3aSrZzgmo7hvzShZFI7FGd4gkc4Yw53dvgOsJ12NzytgwIgqjXpV
dlT+QEniX8vhom0qHnfq6hjdvE0WR62TNrDU3r7sRnIx6feACmAXl3snU0i3cDPa
sFOXUHgwnKpsV4HqwPR1FJST5uejMXU1KrnzdOIxs29snJukUyBUu9zXs3UVHzRH
R3WMUGXdlj8P3/cHakHU2AJVWmLBJJ6eLqyjQCI15ynAU0i8+0z0wyCFmQVnUINo
fkhYqikExi7AfqvYrD9LTyrU9hR8oBRm1+8vFAZ6yDa84CPCVvHlaSmSxVad3+tQ
ypxsHXdM8HEV1BrFSfHTOJFWETb32Gd3ZYCCTFSk/OahkyvOR6ar1iiw27WuL8p6
ek2tMBMVPnsiR6wCaALWU9G6hTljYqLuTTl+432HPUXnrlVDxhbLYbqvynQGFa0F
bm/NMF+ZeshQb6TvRpWfUvp5pmTZAPXhYN31Ei+jVVXq3/klGaqtmJZvkySlT9Rr
n0bhGzfqbUxnK4Rpk87nX4OWJMW1c2cG/VBCKesouf8ChVIJylwz86frAuxENfx6
4VqQ8NAWysfIDqI2QJoRnq7Q1kd/fmeIAwl6W5dDEfq+mZibb1ykvV2MUwKM2kAi
gIjyTxbM7yNCdfjk3Tzn0JmYbVDr5y5QGnw+ppm7cmjbM/I2U8nLb8yt0BDHSuDO
/QcZbYAjZuAIEMpnK8DuizFI290HRZ2uLem4iEUQN3hQwGmGG2e18WRY2bOo5WeS
P/FUJUawnt9YMajFYj1A3SM3HjX7lWnHH3qheUHC2QxURAXl7VJ3ponOGOwASbnK
4W/KB87ZWQ9nstmRE6Z8pBw26UhBJmV25sM+KNhakVZ04lz/rhg1WWbxE25zuhEq
39RMMVPIm8c+f9XWKUWCRvcxfvFPLTkac2t9K+HDrB5j/JwUkoAn2QCbWEM+oSEU
Jtx/2d/wGU9hTarmj02qW+mk5WLr2/c7GNySmEufuYyJheq+9QxoLlh11kll0N6D
aSYeDkv5n1zCys7p+GcpdWfCBC4/zL2g3ZDSmObiYGhFnDF8LoM5hu3PDXa3l8wB
nVkOAfDzV521ehoFaFFoDW5F7Gg7Gy1BclODZXGzyjk4Qv6rLKVHoKX8EMGCB5PO
m2wW4GhB4dopXKLTbtW2vA1U3EDE4J9hGKQR9paiYtmZnSSi/CXHK0qRbX1dOYrz
+3EiaLZX1mYsS9TO4fpI+5kRbvUnebnc/7vyxqvk+fVRW4pi1qyOzx2Esb8ceVrs
EhChHOo+Atsql8SKs3s0DntbWQ472dWbyaVmtqJuY2o+DD1YnAFjQTb59QaRIcSl
unrFnVGh6NkwcVoCJGrTwsyg6fj2yUYV3SfPf+5Y7HW/36hrh47AZs7LtLs7cTA6
scHXfIzqHQ5bSlQlkfsNnQGwDawBP8kD2SRiyQ3lSTffulKcPYipU4lquvm27qwz
j2JGFmjfcEjy227QTX60mCNyA9oleTMC4Rz4mDQ9PALWZ0em+sU9c2gp0GM7Ub36
oEngmwLkzIeWZxbBYpku703UQa75KSgM98sE42y0fvMsni2IvqtV45/aOO8euv8+
mc7sdsJ4rfEI94UuRqBC1+r8PUA+HCkrAONzkIvST1BiGk4wWO45jiJuExW8/yZd
2A49yQn9e1kB3xLzBhL+0WgIvAuoEsvEQ8vPvi4ghHYG8Uuz2Q2GsvIh+P7Ow1ll
WKbOj76fgz7vF5lF0RIgT7SYVnsI1RtCP4cdpIwAODUYeYTM2pHzHWC0VzqEBXod
DWY13H4Wa10WtPYwWV94b5u7OZ7HysltkzhObMVrNW+vqB1QM4sIKyUb36vMa0hi
POH0aeaFLYtbfKBz1ocsqcZzh2Mz2GKIHz777l0XpQtd6mBRnQ9Z469qLJdVLdXp
qMiPdmysT192dhrPvyWZ+uf3IjAiCs35995Ig4US//020lspYOk/ZKu50sUPxJvV
jvwnKLCcFNd4d/WbnkU/zEUP2IooRbm4L5Jbicy3NQ7OViYrU0HroWzokWnCErIR
nuSOrvzFAU9IjDR2RsTcmJo3H97bMmgd/pxcd311rPayUz0pZqvkKh5kMMIalQh3
pKNzc326C3YVB5XlhjOF37IisNwc0uUeWoh3IteqjeNRpsK8o/7IRwtnS8z5pUy3
JkFZ1fAdvj5IM1QlasuHcKuVxbTAJXgjCgPs/4miOaTqRX47jeVyfwSEXkGva+/s
bVrH4POVJeYpJYwFP9mqeuebMkHVIvurq7JDdxa0bYiiQEQPSeZaaYAWFllTJx/u
IIVLqT4riigBCuhO/MKOh2TZozuSZ7Z3lifSJmBaiCt2+4/6+Q23sztKmZePlESk
puGbT5ir3Xp/e7cVQYTm+2BHIv+oVkTf5lbcxgd/mdDKcR9JlFFrsBRKXrLhqWwi
wMui+sVlaKdKBXyO6V0JjFFn1cl326yVLnjTeoWvfwwV90rWKcCEtZRTTITbtcqc
UVKE4PjDM4Z97tNVmC+bnND9vQjeUAa5Nu5QXOhpzXS8/WofF/UtjngLxdEaRjT4
wkEALJ0o/xNRcdcwmN30qpy0VUyWJ86SwHQ9HPvnXIrhxeqcu/8xe+kGEIXHkAfW
BMPb255BS76ShID0HySZWv7+7KQStspgCi/67k8t5MwwdM2ibCrmR+d6EBwMeqPy
qE1i4ySD56Madq4jmPcMz3hAG0zdlBbtMyUcje7NmJs7w8+X3uojgammFdMfPWCm
eSLwrjzKTTo/pJ4bepu0nmwVY6mEjAHT3wal+XjxR++0rQAY8W16hALBKpMZcGes
GxxkBZWZ5rEcGkrLpYWkpb1s7IwF1OgOP7YkRUtrkneUSHNwpvuDq8JV5vT30z/Q
7Jpa6JXDUYcitLmd4d9kCQCd9tvguja2EYrsv/LBgEyGM5ou7LZKEfIJ6fVkrqxN
1J/H1ful7dK7MIGfiedzMKeppNrehwBriA+A+2oS0uuY66P+hVwbrsmrPJMXE8nj
QZr1V7SZieOAPBPa7uozzwpbVQu9bv5akknjUdemhOZ5KgmeD9xoU72tIFn4Tzuc
OiaqKlzCU4Cy9dhl6CLsEAcnm8YWvKIvUV6E4WT1QHIdjTJYsz+Z1KXOUEA62N8A
V9iQutgL4ooGZZogTZl5KWoPTDgtHAZJJ5z65qcZA8mgeIxMj48SDrZsAnFgjs83
hHsX46x8oiTkAHMAfKr1lE4wObhGg4qkKGyTzsQ3qI3G0WHDOZKhVFk31Qw4axRD
Ck4VNlhJzBpDU+ODPwiUxPBEpC6E+UdRqeuIxaA1ILKgbAku3b00S+2ySLay4aiH
1pUj1SO3j7AiEy3wdCIpuGvyk0EOVQZE1y1+EupymJ4cE+XrnryReV3OFPbQnhnH
i9KrVUMUTWnoZFPJTRWVKIwUQSfjYoCprfL3Ofge3UygYkefKr0CgIZSOELdietK
QIFvoR4gL7vHjOYd0YV0snJgTtGWLMkeQ/vYwtZ4g+NLvRCju2/HjKvuMAYx2d7k
OMLyuzRRJuIeOgg4H8HAMmffOrFGiDdjUqSHuz8s0C1337rbQ+zmfguDX5X+u1uJ
N70ejvlAbMp5WRptwjBpURa01DMoc9gV6oe3UcUuSg0fHaysJM6t49MQgiw3kuZQ
E0I9YrM2lpxNRoI++7kwxsc8DOUDf8wUN5tzR0f8DqlRZ4KkpPCwjxbUJZ9JTo8+
wjYuwm8RDuRzND1Xy8uCj5s5fnz4eOFLr99mqWGN0CK+6h5lRSmM/6Z7mPlJ2rLl
KKkLzt1av8OgNpShTqAgUoFij/k4mb+pG7UoeDBS7n2u6RbhnMSCBrTU9pzNYgUa
MzFIUxhGx0ZcQ8+20dMmu102+uwYpur3LIZDFgv+VslkKxYieidV4L67WRrHRdLR
R8Lr6bUGJzOHMOJcGdnnpcGGIhn+M1fBehzzfYjlRV9jaRTCbosshlkPWISnc6hL
ZIf0nriSAo531UeCfL0Lnh8oZtyG+pdbCfrzd28FSyuHIQ0HftnKWmm7vbzXUqi3
EQyQK15ghff1ql3mdxqr8RXIgXaDMHdUP9teG2AYXGqM00PD0pxQ+r3BdTfFovTP
Tq7NVH1hl+U/AYWKCl96F+8vbH1peMjyYUhBis9Unq/8hmChNWKwbTJ7NAh8GKl0
rKaP0tk69Xdl7TJA/O+Lk83GFUozD9Wa0sCcOdUsnLAy/LtPpHHX6GEnZszBEXVX
amy5jyhwx9i654ukrQP5dcv1Na37k1GqKhWTYMkXdJcMWRS3vmQgbISVDrg/L4M2
atQvlT9WHaJEX3ey32t1ZAKkFa6dLmd7rn0lD+UIYG0+xvSKnIL9wxXYfloXKgZC
LYhK+OCS+CFzdeWuvGo47Z9qyKLaWib7XwS9ujYw7TAoqjxazWNsdwTaBD8wkNp1
F3kMmIHr8H7jMV4nV8Qpwv40ScTbCj8NV8i3w4s80tYxpkyLio5/W3NJnc1QPZ3b
upvlnkba+N3HLWsBHCpQCknxD5AVJeTkcDz8+SxCpRVT8Ld8aUvkfv+10SdiveW6
LsaCAkiYbBpofrol2xTZaf+a1eGWbji2/UsaiB5/3UXyVhN9VTuQMFAhK9+AhYZL
sLz4u5WFXSKxLTuNmT17z/jKAo2yJaMjPhjGJ9uUmRU4sUYZ7ud8bsclVGhlIvtz
hzR3gk83/GmvJM4cmojWcpXg9yOWJF4IOXz0ON0xkTPmCTrjoQe8zFqQFSBzeblz
I0D3i/VRFm0mQ9qmgR1PTT+HkAonJSSbr9HKCOnnp0keY4X7AQYfVkLo8ALPI0is
d1061h67KrHMg57NEdXRLhLUzJ+v5v8YiDN1JcFp7G/p5ESiccFtRu3alc058cu2
3XXvOy3I4K9iVooxQqixnHWSp08T7+mnX91AikuDZ+SXOh2wt5DvoLE4RzPxL03u
7ELNOhLaKIQAeFeRuOPpSvk/gj6mdHG3USN7dvXyOzV9YyFgdqeG3UVerRpBUlIg
SWXRRMostD/yZFvNnIwYf1sdKcCOWKJkv/eIpWdd2pouaiY1sJ/QUncfIk6apaaG
ZRlaUwvJXm1tOH00MtTCWVo+ISBzr4ExXjhqDz8CbKO32dlly6weAzNKvGQ0+KeD
zS98IfMQ4rcaJM1DiTF44qORTI/YNz5ayhi/grwyXY2/mMnl8ajc+8Hd1rZZc5/r
uSGFh19Y8Q+ATHPZrw0atbrPagXaJGVoQv1B8YtZTy+un728gHcIwUUmmra9x1fB
HG3AejJWt1qcK33OtgPlLzEHvjJo7BlDqSP9R3j3BhTGgDCH2Wc9vg221pIVVP7x
qFUnRkfBmBC0eJYVahzy5ioXADsSNdkts5W6sRI5fVuN/OlvCU7kvCs6wKjtHt2+
VyYTbFPYjcZxJStje2qqv9Zss1PHdlbeWWgDqikGmHF0zJ3T4ezo4fFWNfIQCFPo
llScp7l0stgx1VX1R/U0rFPgUpTqw7mf5LWDnoWmvRFL7Tw7TeMppvUR0dd6LzUz
8Bell8GsTHK7l/4PkqB4798wZ9uAYq48LEw3X16iizGKKjn7cuWLCNiE+sPPYEIV
3CgEowA+kRAwoTsi8mbaeH3FrYEXBBG0ne/N8qHNfVvWdbIHdI4DT2O4tJ7xg5+c
kC3+ElqqjgLQnndYvVZjjgc+VN6IddqRZujMMBzqSwSafNg56hfKDs6HsjnQ6ZX4
YRoFetUoI9Rxyn4S8qYavQxRAqH9Poh+xbIOqtqTWaCRUnhhF9NHoY8KIAaKYOzo
mDsbBbL37qL4w8D+bLQ9IGtZLdsOVgyhyBRHl7EW22HgPeyH6Bd1uUHxEgZTPLGi
umh1IMMNoODOrhWbQSxl3Swmq2v4LW6kRjLHz0N97D1Xa+CGu1iYiTz8NXaPZ8//
eNBmMMHVjx2cB0xkWbTD1Y2NnDqEf1Wkux8AIqZdr9ZY2YR8Xwa55LDxJBwx9sCL
//MctNd3ietiv+lgT5JGgR6gSUinNoPLFlkpufJJnU8GUFEAswzzATNdS04aADpG
WqWFKBJSZD2Y3mgNBwiLu4Viv+DzoSLmFeRpis1uvPAX8MlTjTtuuKyAwFBDjj5w
4PxzEO+ZmbVsnHDNxQKuJ6eZF9VeswcgxMfWX42JApgjCKu/Uwe7eN8uYJMNdCdv
KuHMIJmNDUeE8L+OA0fza+BqnZ2L/89tmp58WbpfsBs68DQcO2p5cxNRg1GxFOeK
05Ukcd2I0JotNXitfUmH3IKFR43FQ2e3hcE1fII5swB3OZTHQFC2YTdpUTZlrwDN
zJlYEssFGJ6tP3v3crykHYeZOV/sZbYjv/HUx4V+f2jaO9YBjIMClG488H090gkE
cB/lWNWBPmMaExYFagrdH5mYFItSjszwbvUV++vtSuBjqxDyjk4ZDq8mUbtBiW8a
pM9FznGNY2+RrIaRv0kHz6sDTRpKW+CxdWA7mJiHo9qj1oW8SMmYFDHixfTbHsIo
AFDSTiktd9f6smKwiIUvXi8vvtdMeQMEcQVvideEco2qasoaOHPE1tGhUsiwtYe9
s8wZcniWnfnBGersi5KG6d36XxoluvDLjMX/HU4GYVXBpYoDrmtiaVgqnP09p53s
zxSmj+llrSK1fYG9/CMQ9YcG5OLIzMopfdvR99VTiBtUvkK4gaF+ZKPpYuhEYaEC
QKgKTw8ixC2SQm18j1wJU6F3VAHoB2ljBDzgKg4f9MR4bmOwXvxKC/XTrh91kRp9
FysQxaPxjGXCxSiexeJIJEp3i6rRjnNX0Ywu/B4uNqSu/wgWK8M7UKn1WYUNAxZo
L1wBPZ7o7aIDr0WB+K2dQrKQevU8M+TC8smSpvL6/ypU88RetWkDeyCMyYcouyJS
El7fRBq8AKhMjfGuhluGIVScF+F6P2XLionyz8sCGpmL49qlwpVcBfECtqBxh6mH
QIfvOGNPDNJqGgRpdsTxiYggeaVU78TJo91q8jZP923Hno0Ukec5pDTBcK/1s4Fc
XJb+fiqwBH95KXLSPuGTHDdPKpinWVa4PgO1aAbt8bqJIVp64x1EbEwmPfUMMzzq
0U23RYda9em9OIUKgq5SFNViT15Ya/eLg8pXY399CDFRLB8vVp5BLcqFsYsLJrGe
klm3/+PQts1aLUhTO2Sb8OhufVL381wYitkElbRkN7WBVuGkveJh+pLjc7Y8U2aN
Cf/UQS0Nhf/c0iY9ecuCBYrsoZloicYGBGTacChrMJtqUO8EsFB2lyu0DqQjI4/u
84zOGcFrVrHN0HrHoaVb6hsOkY/ljjH4PVEvj/0lK61NNa03TFvu5F+EpRg01BYj
BcxpRlAT0psbqpYdT+fAVo8obzyjuBea7jokp9HVo6DptU7G1Ru3k7urKV55OOTR
KMjIsdbtvnXRIOiMifJ9J8LOt5yHt+aTruj6M9VG8yoMdv2rpy724/ckj5HVvxHY
C/fAtUNkx3nLErGa1oOpbeR5fdFnLvm9vA+GJNMyYWRruIF9M6XK4Vaj0oMeobZN
lqE66rkVkw4nyqL+kEzOKNXf0pRlaFbDQGzCK8JGS3Z+YvJZ54VJq6kyPUwsAUGs
R72aNFYkxjLcvxyKeoPEdM9yq+o2AggqXjhZPd5vhnxZf8HwHfO36Ci+h9rC47ny
hqCDDnkRXSItgnqES/EASwfhwbxs/Ca1Nfzw5UpFFCvb9iHwcIHxK8lXkKI9xBL6
LPL8CiaQxFIdZR/O9hvc4J5gYH+53oi9qvpFuLkWLeEYyxq2TRhEUyO2BQS5B0mY
cDWkhd+9FR2jeIlqC61kEiXak/vWpU9aBUpOYI8HYkcN0Z8xFzuVwTPddpYEPA+M
5/BZPyDzLFT/cdo8odErymyer9c/INb2in7IwSdvAadDevC4AUGhzXO2iLRdu3Sa
HcRozXKYNwsVgX129VqucVlO4//9grzHA+gAyqm4tLfwb3/tCi/U05qHQtka1df9
wgpqn85yxopzrnyxGrimCLmzC78E+kwWewtRr8DhsEEYSXKMI9UZB+L/sl4/nh8s
8aTBnXlWd06yRjbs54MaRwI+K/y/NEMvsL63ozK0kz46VjHeiFiteMAqlf7g1b4R
Bd32TV9mbhX3fEeqy39vCAV+/66vVq3z2DkkICR/XyT5pKsbxJRpcYllcc9KomES
QDGszFb23zQUDpUHiWfLOMoNz6R4+vs321sTmZheni73+FKEE10+WoU/SIYV/7fg
EoQRqRnk5Gs1kL0KzbzY8GYK0oMCi5L90eM2Goz/06hMdI7f6RBItmoUZq5yNTKA
RWBfDPM//UvYYrYLvnpIpG8GfIYSrFMPPccs7NxIK6EkC5mNQro2DTvIgghKIrB6
NhGia/LGw/dTHxctPayEY3uhuquO/IPB6F/scMalp2ek3rHk6Nss/LIfqqZFm+U/
EB8/Q7AeVWRhep4TLiN8dKHjjBQuX5GTvEA1f+lrpCbW9rlt/lAxtgaNzes718mq
NcctB/f911yF/Ep5lGJuRG6UfLXnalS24BGpZe5bHDiYv1oruRYMIVk2aPXOU/Sc
tlGqInOXuw9nm8KUf0UsdnLo/CIkq7k1JEo+DB1QwcdvzVKo1cHkvk2pzZRzd8so
WPP6TzuDQPOHK/oz1C6HfFDEQgxx7kD4Vbb3P2lN5xD1vKN7rtC46SFjheQdlayb
s6QiF/Nj1sYRIyJ9pisBCKg4KGj6Bjfy/2dmR3u7qj9hMxEjfGOFXYFIqS9M7b/f
HZZWpYIm3c63zFbH119TDLveqbEoJN08PCfC3mY7hC8Q8hAaOk3FCpP7PRexzPI/
rdPCM+AxifqWV4GnwYluKZ6i1GlJ2fGDqHpupY/ZF+NbptsOw7+dc8gtXMn2xf+b
IzPDd7/FEBawIdDVHrEPzM1o2VktGTTNRckoD0Ye2YTIb/igV29kldt4f04KlpYB
QYpkZaVwEdOqNbX2D4fl08fxFoYuXOc3CmBDj/17N8PIfB99Zi1AN1Fg2Is+33Qu
hH9/O/H/ycO27K+aleCLKgE9iL5gT87yiq+mbqvC6m1RXKgn6JB8wGIH0htKBXXZ
MpYK8d/EuGTR34kSg+BEliF1CjyQlLHCWnN7eayvH4zysEHcagKxwDEFcH/RYHAX
6oxAwdrdrhTb/xZ0/Rt+jE9AvsedBI0yt7LxUkACAVvfF8NOsPUFEI1JBPNmn5iQ
/l9I1EJy5a9qMirn49Id4W6DSHIG33jOIDkTRKJXNc48e+9dYMSU7qERPtVk2ElH
CNuPzpyPVu+RRcSQB2M3B7aLYq0qlIb6fMXkFtY3xNDKWZ7GhpZ6nSkEjyf9DSdi
uiuknBVpsCkRWuC4iEq5KGP/zbd9t4yXj+RCpG2FBKvwhYIIVHW7C9Mx7x4vEz4b
8W9GYxqYD6aRlZuq4WxdIaacEgoTBctt/jtcyk1X51KXHPbivmM+lmBzG+JVUtl4
s75SrifZz1nJmwmTEOWrdR/l+jFzhQ+rESoFXJnH5m0GYP5q+6k1IAqAf9834Dae
xyJHLg8fQOgjcr1H6XNqz8eIqD7qfHHmA+zMQHYHHvlaqDOpVvuhLFRw6cOriczR
+KouTv1ODjtKVBJsLVqk8eDuI3iRdG8XplKOjNAqZ7gOsz0Xsw8wlzB3uzqttPAD
mpGKyf3/2gxbtTt36y3Z1m2ZVL7ANaxNN7jfFqVFfxrhTDEcR/u7pef3OcwXrWiI
cTGxGozinbLm5VJp+a7GP/rSLLR2yJzUljrRvm/0rrOCi76MOgR/F6z1MBy/5LJU
fhQL2zMyr9qoanLE9ywFLvQQcbFqLj6VunACyc90EM885mdcEuZxjpiOb/caBgUP
dnEP7qqmyK6YaXxZG0q3QvJ7G9YARkhxVNkIuh56nMGUyjpHGHdfQCavVicAjZ3Z
D3CAX1MjGgTXX/rMGVDjs4OkZlihOW1u7sLrRBuAG00JZrw2s23aGhJ8WWF3dM8g
PULu478G8Yco8kbisb35RJkkfCeNrEtoUbz7YoTGSfuQZU+SPnCFhTgsj2eQYYmH
uxrfOTEDq/wLc+ET3RhYDlFkAiDva9nFO1JP3De/yNWbc3BgGMrMuBPRmu/nTpeE
cZ4R9IzrYV3LyThxNew9Rs6Cb7frhvP49FFKW+7C5X+JXdmy/2sXY878aqjee15X
2KM2o2RZjdnILHAvmTvneZjRx2wee3J5IO31vaB+75AJuXjBsESeBTlAWNaQFRqO
ybdJGiii4ZyZXHeCQo0RjlraB48+J7KzRyWdzwq6eUEAqeQ0K2PanG1//V77hEht
Gq/sL0M9lR/ECra9/uAf4L637v5IF3UTeIaEYPfU/9lrfK+7IvFLdv7e0lpeqUaK
mOrriSYGIoiJEZNxGCuaVaFdRxvFS0EWif0FOEHxdxWPGSCiY0cxNc7Q0akh+QSP
tJqUu+xyYzFigy5nkcz2sty6R7zu5PloKOY1xo/eGjcMV7bbEjBH0Q+Qorpyc6Gw
F3EFGyMBo2DrTCpFqVlWKhAlJGOmB83n+9sTO7Alu8qdLQcyaoRTtpw9jXrHl1Kq
Jo56/3xGhMorHzeA7sjitZECZYAl6VoTLCASdGY0Oc/mPJE+i3O/pBFPVAJQtKYw
3YbYnymqk6aKJ7L7ZqDBdY2X8UAVIadeJyunV0kO/ng2TpsgllfaYl0dp5njfk9J
2jxUyNfIOj9avQcfEPPu61UjeA7J503wuE4xaW7m9a4ZetWeWg0d5sSDV6BNIC9Y
nNdUtBs0WvkGocFIXnwIMkWS6EMhvQZTNUb5TREtHniPTA2oA6lx80OY35LTEwgm
1j2pTlHU1srqKVkvWeI0DfX1LyVbz1z4AAQa3q5E96XOrUpPmWE6X89kMUWHGMRK
MV6HHIfnTOcNDCdiuebQ0JlejCEhIZiYIzjA0HvmH5pVufNQnLuaeEqr+1syEVr1
JWHW+rYzSa7TR4NP2V9qrOHcmBfr8b4+s/a+OMh+c3s2tHRkyeuur30OSavB7UjM
hVrm7lX35jp7LB43U8SQtq9vTzaAB7FsUkQPrLLPS5sB+qjCRsF7Lc2jgqkqbrtj
mUceudy2VM5F3kc929K7LzB+58Ri/VBmJfxlzR152gkfZL6IV78by3ZsCE/a6Rml
6k6jx4/BApBtVS/lmoLEDBqC4ttjGRr1k3rHOIp2iToe+n3NHhMfvtAqjULghxGY
XNlGpacOwR/hfRgD0uLYjADKZ+VJgP6bShUW3QSyLQPKsj07PM/O0j4bfgOT8vJA
D1OZY02lfSNJAS+4aqD5QgWQJ35avxDW3WuGHTd1wabeNaEH+HYZcs5e+YWYf/XM
ctHygDD1DiN4eDA+TcqoN79nK0WnyIpg361riBaTFf/lrKQslbfbU/E72SKjkTmF
Dtgpv3V90eU70J7Ad2v0fTiTha1I1SmcqZLbh1oe0kSiqKEz8MFnajZV4cBVBB4c
bRw4kdtZ9f2thWWNWENspciO5aqvREBzNrlj5jRkSPCdVF+e4PWJz/W9njui2g5t
JsHaYNlIrh8XO3uSSXCom3volJRkhZvYrf3stLCmFQ3RLCvYyLwHRwq4VchpSr9i
DJuz0tup7rwigaUGQix1btNwt+PqAVSAoxPukaVFThdMEr1OXWo4ym+Ta1Fb9UDB
tyEgGRLfeypJH/uzIFOgT8XFrNjwLnRQTfA7ijZsSFYnUF0opGDTtlAQGRAkodJs
eOCtsSGOLUnfGMQr0LNAkdn144nxIXgBB2ffbUMqILT/dXk+T5XotINLgk5/HjjD
VzC6Y7gWrIAdWZ9R0S/3U1aBfbwGga4iTr+C9cqbFNkUR4nKsdnjd4olFvVPXfRy
GVcX9xx/pxlKyYz4n/dyVVMzLmPFDeETo8kCXtWOC0fp0GHf3ha238isLJJ8zGAL
k7TFlKnqYItym5FkeLYYk9UQfkilNxOSn8dO8x4E+Xz39B4xjft4Oq53SGPb20sA
UBdOO0LWTcI6pQqSMAkFGPs9HEEIDnWgjf71Rq6W0vCnaa7iskdOCNyQ1gfbJZPA
MKh51rch6PrM6tphl2SARwo2Jn7ijPUFNTh3G2OtVH2EmneTjYsoPZprPFewAGbM
j7XJycluaO5l6a9fii2bDQ78rJINf1P9reFxmy4PsNJQlAoKmfPJMSq8i/Iv18v0
sjqXqKcXp5fAxOXxcPYbbx1nA21ZmU+ZvbQ5S5K+QbbDuCanvfQVhZ8p4E9LQGW0
CfVOvhuyoPeEGXmOXxqKMIvxnSO1SqBXXFwrwPi+QK23m4vrFJBbTqyqQc6cYbth
tDPsv/P8KPHk//+xaPiMU67lryQXjhAobducVlOK6gjRc59yUqZ4flJUcEbCphpi
/t1lQFTD+nyui2ioJFy6Jm/5CXFbxTYRZko5ot+NALmuF0WeQ7kl4+Es+4nt2PqC
kIlklfqJzGFGhO3N2G7fDkJehPvuF2WRvKEcKFZbw4R8Lw2PTs27v2TB4HyeHiio
BRrz2xJX6bSmNwQia7wO6f09kNIAezWCVA2Voy+jLswVMviIvbSprw93CJNgQjPs
A5BCTVmnK9FjgJyiDJehpLWY0iCxT4Lu5PWigYdJA9HkW833UnQDhxeEjHmDadLK
v2XF5JmWZgTQi3WVJBoCClSIY0R6VUgW4hogY4DZHq37cWGNWeuVic48fSX/Je5/
jroqv5mFk1eycIKZYtrB8sKMguHg/NF8FIE7zJPjaiouqdOlCV++2X+Aq9iR3V0C
APgsXGHjoeAbS8VMEY+2+BvIfxHAHn1A+6LjkfnqKqZsMCGlvcP29w4rG+SoftxT
xi2XrIimx4SaeaWDT1Tbfpcd9PF80Sqm0SJK9vf6gTBG9Q1YYw5oePHao6Jh4SOJ
UZPINRjEMpu4/pZqOb4hK0o+54RUi7xSgNp0cUgBF/O7cEJmQj78aDtRtbvLlLs9
n3enn9sscODqvnG9xsK/muzyDjaAMuyJslHmrSpVXVf9Z2sMWHT8ZcBON3DiZYdH
YFPZe+3gHI7Vli/X2M2iXabtI/yPWl6ULHpH88NokakgI+GLtVDFXKZw+vZtdCKp
XhS5j4AMO//PFR7lZJ1Y1rwioOushYS/AnjzD6XbnmCJu5N7ESgoqHH8C++e9iDf
cC30nKJi85c/zmc4vmuSa1chcM6eFniQRNu+1IqI7uKzx2EGVUAJEyMXX/ciSYln
XSeziy/tYVSY+45zzDfQRMj130gqhqz+plJe2ZwVJ7vStVefL1+GDX/ammgreHgC
FdL/La0teBiR2f3bh3r5dPAEUp6bIpx/S2u7Ts1gC2NT0cBBKezr8fM+p9SUb4hg
avHjiwcYatPRgosBcNFQR/Kg/S5szQ0Ko/ukYtWayzxTNcJCgj/jrJiRHd6JElpC
/I7xLG7WOfHHSxsleNIoPI8hdye+GgfMIHRHnDIGYiZuMS9qd+DwrsTbCOTp4NYw
mEClQZl2951gro2qmOfRXzRSdN0roKiPFScpKbPiucLTZaWX5coepkZqP+5wNUBO
phsYU2KwQ0Q8naur2mbMkh4UJuJWF7+QzCGVFTiduZ2CvPVl/sMOp1UpxenPlf/0
r0TDSPo1xosCHw/66rLsdQBES2WLga5o7ct0QdMQ1qkqM4LawATu9JADYZSmEX9S
Q/uH0pZGysjU8UIA08T79wBA5YqVANk7HDx47CEm7wGssbB9+bu8U0FRxwsDYX8L
T0Prn0GXYRQZKvkn7cV99p7pac/F3i4A/P5wyTMCZb8c5aWxKpPEt4Qj6t01l4pv
N6OS+3Jx3LS6DDe6TaVGbTU0AfrQF0bsiFLyYHHFShOIXyeMFmg1/BQEHU8mBTiP
LsCm0vFbO26tov+YLidR2Ye7cZ+KUINwc8cb+dkuhOzMX2D50OCGij+avw/ZWtkg
5OYo3cjl1EzwVx16Ce8vOGDZp2BhphG7A5FHWlGRu0KQuhejGNfDdgT4OCiAvv0G
UkcrI15Vy4C/yK/ndTuTQTbMdeaSBQFPRr/joSLu1HraDr8djFN0FEO6+NY0i3jU
BPxCdTJ0kVPRBK4cspSj/B6hhE5ScQwZ8/SVlFwZCZAthgpe2muosZgus/TS2SOp
9vnJ5iYMg2yX2LbfErTee64tU5qiVdEbdeIwagkdm+Z5mqExaaz7dVxxamJ8TPPu
EPnMCkBInuZZYVDpPsuAVBNAHhbKKZyw/d60lmU0L6UEFq5OmQInI4+cboRc7wCn
XNFzBV/9LKGVtdhCvqKsSwgjCRrVN1MHHB2DghWu0si+1RxMpYWNW+KAtvnMygLP
nEIizI60MVbcR1kfxU3yZWe2u+aU6cN1QmJas6LVZ+KxF1tL6vnMmeYrLzFu4/UH
9tBb9E2k7wZWOUDGwdAnqlA3QmEusfUS6JieLo/8P/PDotRskiRrToFpVmEHC/Px
k8D+6dA0J20dBnaCPPMymIreAsEzCj00FT7alrDmkZ4xNlu5vnju/94XCFjbYfxV
3g8TOnlnjQZFA8Kx1a5Cq76EZmr6j/kDFqvV7sw1M7ZgwTOd7hfkMmmJiX6QPEkp
BWtA0uexJXc+z8Ej8q7xvFzwt+5nI1luuir5OO2d9Ov7s59+quurfqpLpzJFQyO0
Hc2Dx3ElC6h5i0DZb+X/MeBTOZz7EbTEAkpRFpDhmudRYMBGw5YLUHOIjwrCbYDX
cTmKbU8/5Ui+gxipw/yRr8G1SN3Ak5Kpx7UaUsBHb+ge0VPkMVOciAp4OfT6kESx
GMl2PvY+pfwY5c/tnXyf1u8fBOBrZnaQ8kj1zrc25vrd/6cm5VQI2aa2fjUsmQih
zv7a1TNE1vKSleobpI+sBv5rLPvxY9Lqp4AFdpq2/7sMnNegJ26lvLlCEK1GcuVw
hsBloIu9+8Fg3iZtvZ42e4WmzbgHobXLwA9FVHXVKf7P5J3eYC7F2GmZQ/CKto2z
U/NgC4Pats1IuGT+sxBk07DHfHVtEkjHz7v+2+7hhHS4dsiuclF5WpyNO92Ap3rx
CY4wplWqb2ERKNXTtgySBPaJADRWnued/dt5e42/01na5miBtLj+yuaBzk+aLemB
/FAiwOyH/dFzRLqo8vTqVUc3CGHJuf+9vU05Z91G32CoiLmLRAwthnUYnbqTBrWa
hIdCaaj2G/KIL5r/6TSMZflqtUoKQzTssveSrCnKZZW/OA9BgHDD82BvCRS+gG6H
isfQ6813Vn+idfOkff89XXuwTbD0dpXbg6R/wQ8jGQqPMI6nM6wNKZuFg7H8Qm2a
I/6cEvJPd/gGu2d9wdaQrQOYj6h5L/SZHGqJgyw7GetCoCIi6pfz/14zdrbWoahb
z52KMAYnHSD2IDna/RNgNLqtAXPU46+HUTfy5zi8fR1SxMPaznWvfF/C2wjasmvy
qxMZaLPE4CsFXuTXZKuECEBrWIXdkyh6PvSLkxeawHWHkKLlS/faR60rMnz/s71E
8eSoavbrH/Klj5kqDuonX7Hm6kx8zeRDX/urQLuydYGNQZuMEZmvPOwlMHr6NM/Z
mexjv0Xe8+yI8M21GhrzGqq/bZ7J/EiA2hOoT1EKw1yaNZEhjpiDD6PhczG92CnI
w1ehRQpPhWLd8dSNHKKn2+imcRn/LBi94kjadFKIjEJqvHxpiyXIMMnuw0y5AcD2
aC2ofT1dFPA6zQCxEc8zmBG6nUN5qAFog+3hkVR+WaV3l6MSVwDAI60WGPpD+UOc
11vP6W51BsPbsB5/iqZ72uekaHViS1p4hZf1oRh6TkgOD49IAQ0QN/mJtI8/Zcca
UL9L1zynAQWbqW/EYeV+Eg0DPLL82bFz179+kqxiYZ8AxY9WgFyLtynbJ3DLbSpf
+966xK4ArSfc2dCm4iGmxLHqc2qLo0t0FItGuyx7WHUVnPFqWb+TDc0pwuNgrA0I
X4dF/eXoU9jJ8DKUdn8oQhWSFdmh9KaXXijQ+jCSdtJooRyQx4pAj605QBTMSqUP
yXf5CEAxBehBDlWV/X6i2ZchmLQHwwFu6IbhrK8FxTKn8Ho86jDrWIq6+DhODbiq
6z3TzlRl+v/bbE8zvlL6wZkHWC+E3MU9dqV2hNn7W8ByxiswduxATADvnAyYtBwZ
JNhCMNV9/APzPFXBF+SXSRkZMg5RwAdBeZgjsmOGxTZBBJ1zjPgifF7mfjV2bL1G
+QhpFSwfKUwaYT3dRZCBiAiI/ThSgPNDBCAr2kj9oDhClffl4FK3hbtx4gG3nCLe
Tz3+lhIPHrDN+mV1QM2MNnJyrHG1/1xXsfavsvrkLtvJAAUHnoX14LRiJAAqMB3z
tGRw8RwZbKWxnXK7uXcWodDZZj0HJzHRAq9aDC34IBjjJWtGHhyvJEozpuVGxDDh
pnwQVRHJY6zX46Cmya7HJJYf1MXVu/1pA5rYvev9ORPrQZFQujJCq/n7un2+umyT
w7R5UdXcEOL1/rv+mEzGLo7F1W0ypLLWw5tA25J8y+eKMse/wy23Xx2PiMAQOHaN
qNEMvcCUuNXMLi+h3X7yLrdiSNdzJYGFr0YM011HDVZyC3DtbrpV75TOA6B7PZCV
gw/MCuRnKucX+r8vhPD2RqB1tYM/OYdj2+37XuPZeMULNGSUqyA9uVY9RizPnw50
WyxMr9xmuKV60Ky6cvsd0EnCJhQNOPDHD++dBOZp0kx53RQGkTIy9Bw5TsYN1YQC
rcubf7kgXuerLf+N9+gTS4CIoqTakN09rEmLO4jdGvgwlU1T4eFnd/8q+Wu5sGRu
PoGPM2+c9yMJTnjGTvZgPXCta3vTvfnlpeJ5vK3hgP3MmmzUk1UiUwDdp3jqF1PM
S1j0+ufV/jgyrvRUKpuOk+9q4z+FevxdcPEQ1jpIzddGAFz+YHUAsO+2oBkeOEzo
HYwc1MViF4iqvV8pwto0AybpGbICKOUffkuQMNyDOVaMSH+G33AgGvnfHVRnA6E6
uEmjZyxYSlIGfq5qfeHuvQKDpPknVxHQZ+85Y98jkZvQGyqq+4brcggj2ozdqvZC
iZ02MIYQKcP17wW8SoJogPL3JBnylfAptRBDNxHoTWYXfvkvdNmg4jSNtX3jms/H
ZT0zf4RwXLjydzND3RICbcLXkaAImBGml4KjW+zkSHtXDu4hSWnxiz3tHSSZljql
vaX2O/q+w6E8sEbbVpRER6Iw+W9J/hp5bCgeeWNdor69BXM2Mz1DkPvECZY4C6dj
TrzQFdhfZiu5xcKdjEuOnWiFxN2JFN5bez4BnTyRe6uyOX+LBiRPTAKq/SMdFo4n
uv1kAM4L1b13oOsqzzri43PmZ50t1ICz6xGxcthaAy/hTc7OEcvLHmAVKZ0N7ukK
OR2f38dzAKmW7nip37+ATrf07qRuHxbl+ADhh6Xb05CTRsqOrpj2g6nI6X6j9/72
TyPc5N/4K5kThNUrigikhz9piJTAwJZxIMUcYq/jubRrofU3XTnYbxif0jv8Fjqb
5XymDvHTkqkkYiagWAEH8PgXPtuItaRpZZPRgG7y1e3jq0vfqWi/Wm0ltFjdOJ07
6H2Z8rCKuc+SS2KTDWj4avyxhOCdt9wiV8Q9y62sgy+0QDu1f3CrzHQX5JRhRYYC
4TPNVh9DuvR5akYyB0rWMIcc1Mx6ThGY2TVEjC0tGMQWzDn4d8hO2LODUNiLnCy6
36BW2WMcxCJL9tZE6YwDXgLOIPOeDsxyt0jfokhJVvJm8JDVUqxi9Ty6139OSQ3T
UXanJcjXwEJkdiR0DOfZcr84IcoJ1l38TwTWb5NIbUAHjcO1mB75H9q6cDRwW84z
76Ad7k2BUCwssHw7rfXdeGnwYwTB7smlx8sIYFDmAmQuREWSfy6KBojOvRWqVjcG
EveiF9n35AbPrgg0oSgIeMcSVzVi9l7DDJY0HJ2FuYFQCXOKggT1ApypLI+X9MR1
gRWFv7gyGkY+JktWFuaB33xEyUCWHotmwBp+wms29Fh+BiPr0E/PvGN7GDUm/9rK
DdYcPBhEr1rUDihQ/Tx4DLCG3+SLnRMGnREmdGCHJpHF8CevJ+2MRc+vFJcPI+wA
CIt98VT/QRpAIDGN0XpBBZFF0tcsNE/hGNL+I29nYHlMw+WjEARMlG/BKd0FOJgD
W+KvgUsAVE7/gmPgBvVhUNDsXgmbJXchVAfofMseI8JW4Q8PIqRLCP0hufDiqcvK
NU9nGz1ezsv0JrllwEkunPh0KfCBsGwYzNO3+Lz6Rq3rUjYPJQzaB8ck3/ooQY5V
ELn1v4BaMsnu1bsGvXkM7tbLGxRnH+uxOxlVQoTDJMmDX5RbYrNf+DMkwRaYZBsB
yzhbMhNeBJTj7QlQjNwaMOE0PhTbtN6ml+j3txV2Mrkts7kF1BWp5POcx0xrHJFk
5uvFUWq4A63w1QHjTqCNLBG2jqJfwEKQp2oseFz1FHQkNOg8KKbW4EwLyw9+/Nvf
LKT2Wbd49j42dxciKx53/cUcRpc2hxeRxt+bOP11eXBNSg2APSpzGMzjasdAXHF9
xNC5vzEn0tg01KkUAT7QTE02aovHhH0vpTJTqFGztXatPpgdRKRBl6fJTzX1OR2i
fkFv+9xbVHJoDBiidh3tz+trvh+Zm+yntF9adshPnm7ZAnRzAuYfqD/ybnIcLqel
mjQSCI9Jky+2AyVNXkUpv45uvLCz0i0vCQ6Y7l5sM+fMRAzMSmrkUQpBEKmwnqLU
WEee4FF0FJ9wy0s9AM8gGIi8dYNnrIhWMfKKylizX6ScDJSOzIDkFo/0Y6nh+EUn
5rLZbkU0Yq4xi6ylzAtus/o58gVTkrSsaxroSy4krEaE9V3isj1yVAzgKms4TWlN
8+JIZo9dY/vXLgcboIH1LjZ8/XfQDZiLaKNLAf6OZxdtSRvJThS+/mVCa2/9yVU9
Fg+u13PpacszjS/QeDD4N7nmsMaXdfApn1/krw9UisEr/E4dIbHToAtSggGBmonf
rKjbWH5pYQ1GGN8ETBRXy00wNuK7jrXIvcGuVtNHn3R5q3f04ORfZ79bIOpFUCcb
XI13X9De8w+O3oJ0J9kxPZG6iFEL44FihJhvxwNKlnNqaAHpj01MtYRxNM61OZ6H
WYCuPFaqZLLiTKykOf8PQNeIa9wYNyiCgnyMyniPJPGdmxC4wSUopLhtbbMKmAKS
fvev6RyzvzIS3peS6KCB9b4NJx0WMXFGoEgOp0sBn2+yvzx0q3PM53rJOCFWW0pP
tEjon3LhESTeieQbMQOJVWFJVaKdAhcfh6846HI/ydAQKzs9cx2DDEgBxqWroyhP
pgMDu/OX4DIMlBJMpu4CK+l1zWsTL2kuY6FiXE0Ga394VCD7aDVnwSK+lTTCtzR5
P7R8vwTWTrt0UqkNzbJKKiCrQAcuR+GpOi+eSQsQVVOUkdBx8rgfthkShX637oNL
mw40bCGZEcKSniS/J+f05O8wb5mgDrfyFwm4TUay3QTgjQD7DcKgyloPmT+S0gwV
GjbX+EZF2zNrmX0BKAIU3mftJ2g1XOOseLczhbWZ8fQMnlJpPhy67IrzDRxegeH6
/bdtsV/nRVIqLf26fB4lrrdOnS+kibFB3h5RRBLgI4JISJyBUoyKO0U5Aw9oSu4P
NTTjLQQ1j4w+Jz4MpjumMclWAw4HAd7cK/gQml9Mkaz8BqaAWWIlW81Pihe4TmLe
l08WwKJw0VNhBNH6IuCFGiXfQDd0lY4zbY3T372kxzQjhCJx0HrnMKFW0bK8vEPk
OAEEWqJ1qfq7NOU+emz8t0sARh68nrwrnBxk5hz1/Ng2J8VkKDrvgqjaV8cpiB0S
833yBkb+V3CaJh1SrbyBHdlIilsnlJb8iaUnAgX61qlL+xJV8fRAYajT6xhlXN/z
eJj4sv7hZw4NTrcKzsuchHFSoT2/WTdnyjCKSORZ6+F6US+iBzSpotQQm+oct+Lh
ogcrlaFkbo+FJvrG19szvWa/RdJthlZiGUW/5OxQEyt9LeJDgaTi3CMN70VRz8Bc
2FCcBvwP/6AKXUhx35pL5Sojig0Qm3WkCY+8Cjcs6Gr3mAG1fuhmzxdJqKiTRyoH
V6UcSl4JSuukg9BXYE2P8gJUgaDEYXdZg2cY0rgjRJBgZ2EHFyk3x3N0YWluQYD5
eGZMpwyWpugMQ5/z/9FxSqcJmp3vtDwJfu/iU2L6qC8GgTWeNmsjfn9YKs8Yi8ji
V8VQGzVg/0aIZ2q1CeEVJuFWI/XFIcKqFIC1VS/wAadXHvvd9gb+KVpHdL/ii1ld
ugAoUlpMJZDvNJ22pBDi+zIv5hZfuUK4s/y83Rd0o5VdUL90n+wNpNhI+16R2uMr
QLoMGiQW2BBxb8ZoXt+B8KlF82dMgAkpo58XCI2LlIHAXw4Zcx7/fDpXVqbSse34
lpHuyRRBCkVjCRVd360NS4lACNXTsydkthZYsPlitPVrAZVsCuDeJiJfW7i05fii
QQhJWfVOAaMOm6TgLY9s3g9jNVqxt3JpE8mV9Wc0MSBqkSMsQiyqgS3DWFQGIktL
xMgLEdbs8TV5sePiraGUU5ND3grzHseZDjD0HAkqGyJ5HR3XVLA2+gtu5ooBJkNw
Qt8Y/dpdvwBYjxSQKEX7X0yT0iQlI3QhnsjJhZAokr/7lbIsHN4NNoyMouvqDgB6
83G6aDaHjP3Ko1ecp4RRnAFd0em2qzFwleTSkPIEaDXQwPfCYTMS88nTeVMI1DWX
o2/gKAUQK+45pWcHbprfqHI+YAUXcFKToxkdOK5ejA7x+C3hGbULGYXyKDxHhpC7
9G32H/tWWYUjznGLnheK0ZTXJBnJkJLGUC5b6RL2NiFWXf4p87FTD1ZYSXTn90Ys
a7P/mSiJwsdwYnjNqpAiVThuk78/fBoGMxeHGc0Ly8E6HO9Ax86wBlEB2SaHh99E
7TbU5qxCCC0lwjtW7ipYXFbte89qXSPYsdUvqAfEfWQKx1wvM/Go1GJNF+FNz6Nz
XA0UVsCptD9naF3CnWkwxkSRh04nJLt4gn8nUtL3b/VcOaGxnOqJMSBn1oc5bBOh
p6HFYF3GHgxyFCx2L+9oyEPkzilqxXAWmekEsEwS5LGcmb53yDYm4f50xqUSJPEO
dNTUDgXixTmGd/SHkFQ2ytSDJ8CGWyiNzYLSQ0JznfRo5hAvByZhGmfWiImxrqp8
EuhmQjG2epdlnTHecN83syLT4TJg7g9GGOwDOq3sy2xzUAhB5XmssqlUUGCggmcw
JWA9hG8KBuaEpU1iC3/yCFYbCqUaNanrU4595zMXnTYyOQ84DJQChqIgKmkjKp9A
4LdPm258ZKbzJzdy4ZxVBiCvhurbMy1g+/1lUr7kiC80tjIOsy92IflFsfpfmB7N
x+CEtO5CvSevUJqvxyQrJe+DeSab0XXK/OuKcAIKc0LwV13BrQ1MiVdLQbYxBU+c
xXDFdF90EJqp9wTWv2p+ZGT/kA0BXXWFBeSO74mKfZBaoE40A4iPAOhHeAGCERhs
U7aQ1gOtUzM7JpWw/r3Z11fxfIPyXHXXvM3j5ccRe4iTFcIrEUXqSKxtv1jEJfSS
IueGOk8yJfWuhms60luviokUku2gxeE0CQG0QYT7GDkEwdoww2s0q+i7Pyo3IYcC
J02i/D27y6n+3lThCyFN94rRMOiYOziXOg+UMB/fTOzSpRzKl/+RoVqlf7/4X65Y
DBwsK3AbDEe5KyDCzu2LQ79rbaayrm6SKaon+WagAeYizBI7dQTmM1RXNtfnjb4n
jFxIibAnqFGk10X7uOTVqe4GTH0HfyE70iasuIdW45Vnj6zGcoc9t4TQhh/aFo4l
/KN4Y/9jGYuKeqF8TvSe1BShnkAp7P41+eBWdjTyTTdaObPKKWSqm61u3hxT1lxx
4zELH//etmv5kiGvvJZrMP2F33KYJ+DyghOZv6K1BvNfOt4cUZinoR+ifRDU8aaL
Gk8JI9Z4DZub+Z9DWEq9J6VPCLauviHs65H7upWBIF1HeilM9t0y8wqWo+UypaLq
oB4QZQR408dSIxOFc9XfBDenaCRyTXr9eJGJHWL2GrV5Zrww4YZ48LrrCX0XUbKu
H96GxR77GdfM+fsVCbF89NJtSy3k8UXA2DmV68Tmd+ihSdUm1Wz/YsgveHDOhBrl
Awq9iaxYODiZdoJ1u5YA3iE33Np/+P/RHdx51RJUQ12tEW3KUODDlxeqayhJbbt/
S2kxn/NysTUV3lMjdawUOTdPsXrAiPwiOWnsfXMJX2znAF03YjNR3zF83vOmFutS
+ZmoqnuJo4Sx9iEDE0lxZgWC9dbFvy3Gx0pQJV1jS3VUVmRZoBW1Vd+XGvBatNOj
DBHl/QAtuOcEZ7Z3LFwJcZI6P4AW8ITCGZWJZ9GzjWhY1CpxjWdjnsuCBC1/2eII
pX3O24T49t4NI1sVV4uwLuDRPfkoPfVh2xJp7F9h5cxGt/aF5oHgkCFKwFsmUsVh
va2AD2FymBXrEO280gR2TTAyVpun7T/7PDWnsDDMCpAM7S6SDgdGtPOAuENmVZE9
8+KyY9E+gBTRokJKRTWpz9D0EODKxaLGCcNrD9MMmoHnyERTJEKEDQtuzV8esQLx
RSDRwqNM1z5gm2WdVtDx3M0aCp6rIzPuDEVWiYRg2vgMTnt9e+c/T4dBw+ZLqTJ1
XTOxrZKxw/P7Ul8rywKxrSV9d9lxEjn5N4NbnGo0RyXkScPr8AEQAPcFzlxla99l
9L4TAp3mO4YFDEtjyMCD6VVAIcto7OAI+egcfPHfoFj54DJ5PTxw6ha4tYe7ImN3
3yUmgkJet+6ooFnmYdhelGtlqThWqRa3m6NSsSTimkCm129Xk27rhNlW62W8L0Ew
Pu6HuNPoEmRYXNi8MDqlgfxL+jVFgjPyXDJ5EDUVV22oLCS+A5QX7neiAqyHGkjB
1qOydbN/oGgwlgJvB4Jn3r3y1CTaLcx7Up2wN3k93d7M/OHBDZm+J9ca9Ah/P7Jy
N5G6izbaKkqXaILGA7HMak4eLGt8bzNM+ggd0rFnu8zqUpXRbqgSPGFVGwzJkrl1
naqEi51vagbl2bEqEjCOTrh/V3rjw4hUDUDDLiycohNs82O+W2XeOlvWTjH9gjk2
7971XkJolFZptlJElFgY6tjJ+uRFgZaRcqsm2HBaUtQfByZgW4Ib9NQvz334mY6q
q7nbn+SzGdhIdbolq+XmFtkpl+d8SmKWizpAuRtbZT3WoOxEV66OR7kn0ZJmLt1a
02j+1WmfXkFQI8TN2BptAsBbc/XlyYWqCjxIQCw/XVsbu3+APIo7pwm7x5W19i7X
z3WI8ZhaM3RxpoYCMsqXmh2tNMEFt7yWmnS80MR5euyBpeMNKOGdo+KRY2HZul1t
movcLFzQxYwBHfAQs/QBESCcJLSzRF77Oc2UI1STuGy7jHFVM9Jowdu1mN0c+ZmP
Us4yPlhwOBeJEO/i86ZptjH98stRZ9mr0yNW8on4VT57k1NmTYPEGzZH0WSR2BJE
7o9oXBlZO+D5a+vXdvPTXBgXpRceJ7a0/FW61WRYcbZaXXRW8vdN8gXMqYC9cx2+
/WrnYj7y+gNvISD6GQeThUqakHMuwAR0nToXjN3pH4Gbo8k5F491EFCCFf9qZBjM
1obA1nqISIWuk+Edr1EnxrNKyHoZZNSTphnskfDPU9++zQskgd246wbG7kn9WsdR
8v6aMTNmmiN6dyV7I9pZckQ1ZDW0Q8xvdoMFaZC5gtFsIVjuDMStV0t1eZtgswG0
NXvh1uoxSYKqAF9vTVnPnCOhxUdPC8SlDCzFDHGbvL1GhrM3Ilo5M5JrRT8DgmW3
H6S3r5RVF1SbziUcNeEM0qWYdKlYoE9SsvgGdMYJUg5xqnXJ0ic33hsExpk9vHaY
DXVE7gbxhk/LzzmPaxWS/OqJHNZuoGRLUkK0mIj4qhQPzUrpKKFylc5wfwUSg50l
Wkrg6n8IcphOBX6KhRxi/jXC/7QtRt7f06ptjbeZTtNMFdTEwU8cxakCUKPIDglg
yGIzacqATfSlTYACyUmlf0ZfLLQDtTGR1ssNTLMyNlL1SvhURVA/S3uLuyM2/V5a
zp6MdWJhJFOEGrPTUUw5ByPcM2JCIrGhirCsrECYrdr131s2ZaYdRVfMr/DDyZ38
lgGWg6viBriIzGErMB9t9L6zPWixccqFrNK2ugA3ciZpHM4Oa4YfZENe0Ov3RMoZ
ZgIZxuU7g4A0KbulshIEFLPDxWQhuzCbh4u9vHlaj2dhcOZsBsMXX1rj3J/WPudi
lL5nQsDZfYlvDklDQKT6wiXLGs8po21S+bJQsE882OLGADsN6TU/44yTlZ54p9bb
R16fYE1Yxq1Wmj1/RMxaLk8AuZ3M4MHvpqFNhODrrbOh59+r1bkAvayXVzY0U8bf
qBqrsGKrtTdc8x/RhonqHe+ds7ZU0E4m2E5gznsc6/ayTge5zXMjGSxeE/rLHSEU
NT4isw2vnj2U16p1xB20SgNM3umMVXsKwpqVRNzD/rVPfkWIk0chhrHjdy4qQYNa
2NDMLD7nbMEuA9PxGrnauOzUE8BZJZsRpemQBfkw1l/jl2iv8QHcWx1BYm11T8B/
OrppC5Q5KSWnC3lLuRbypbM6ONxuL7A4OtiTxz1d/DJGpEcrG7nQkF2tkEOJ6kut
jkXwRwqs85sif+XDGW0VnrEssXO8wOrXbqe3FaZNm9rrxJtjexpZ4kXTKVmIjVio
bMeZuGvbkeW8yZtePHs5yC6Zc2RVsBzIRfVbAF22FctN1g2dX//YQl6XlqI9p5Dg
GcKiHjh12wDHZOUnXNGwQseeuf4NVirQfBEw62WuyX7uGmDsdtU/5leACrJjWMJ4
dX9HBTgdIm433E1gzMRxPCgiBV9pxPO0OjQYmCKpa44JNAQ+ekqRlJBYXThiaD1e
sGaZhKPVBWPB/uE9gANH8q3t+aYFRDpNyiMnaMQ/o4TCHvbKPKGRf9A6aspaO0UU
nwhcdYElSUvN2g2o/jUeoEIKUwHtru8z4vq3AFD/xectOOpk7pWqwbAgnt4VbB2o
hj84xE4CPgIWRpEJV1MEA69e80J2p4jRyf6xa5gJ/xV+pAM1w7zFxQV6Hen+QEI4
tkQWH2tHCAMuia/zK9vWRvsmTYIde0sIWu9a5N5/UMpdg8ybDZjdh/HT1d5e7vQR
+7OqwPaFsmKQsliJ6sC67y5USCEpPIMHnhRedLc4Rbt+WtcopHh+ceF0jY3VOjkT
1DVB+0GOdy4OdlOThf3iS7ikBl/7z4DBSkf1CkexccmJtM+JcdtPdA8HWY2+YBox
It265T+SY7YZsHj9y5dukpDrQ1KkuWxQIUunfMBOluYZKjUkG34F07npYzXUYzoo
TL2ZrK85qQZ1/7KUAqZbRYDK+dqWFQE+mTq7ZmMe6PQuhhvESxA8nfvHnSBcUPQb
8x9TIVnwbCFHXDgkLsUmclBLfO7DpfDR4Jk/tXUwgw5N1KkIoCSd4awZFBAFHhqg
0ZO1IJimSC6NX6Pn8CLMmwAP3fBzeP+BNz8Abfm9MVKwRV+1uevZXTPd9sDqQYHO
ggMlPpAhFgOupiMRFF/66OqdXe/+c4v05Z75zsv4UG1ZtVOZEg0ZznqP3Toef0rb
Ijj8TikhHocUhaCp/uXGM7+xMSUy8bXlTnuvMnaFc/oMnRwpr7Jw+NPPwXIKSSZK
8IYD4JtIrQFCkwdey0zkozArNF260ehA/sp7wc+Qshus90dZhE5gHlunXJ3jXCS7
09hfR82FLsz2CwK3kHoh/oOwELd+u2F2TRM4qpT4ES6nXFgP/mVwld5FHvBDerN3
rntAVr79Jnt+9EEpE3gyy/E6fz27J1MtZdZi60qeZnIEQymvDmhLX0hb7OtQtJ3j
o2PWLBhQV6CjgkWxZXI3vk90aeyixoYssgYI01BYCP1yVDvBfh3eoAoAHk+Q44Os
Hex+ClIdk+CXUN9RUTyZyXiFuSFTL+TfjHn9qqGESEi9FapwVnGn9DA3QpsoDk4c
70nLBqnn7Mw9FARxJkNrK5Gl5KenGyFrAyFN3ZNCywOuRCzBbrKwBM5vHqdR+4+G
jS7ShjUZ/8Kf1wUum3WtqlasAhKkuYteCncKMULiycaunQ4qKC6aBtHWTXC2bLzS
C4NlwayvHn7bjCLO5s7PN3yYtfK88VzrHXnsFuJ6wtnC2aoKDsI4jh53J79rWrsa
1p5Zbh9lo5BYjg3dt1N0LIy3WqBASh/f4cPFdtZZt7tDMvysC0sC5p/w4PbAvfwY
BY0EpXyALrIESJooBw6hbDAAAGiBVYjDhDNjlUCWKH/aJg6W0hFZZTR4NOEtxnNN
5J//7oBCk6FP5yX5N50f2oGu2IV3ExPF7VWDyXHejmmqKMB48aOfYXrmNnOd0UHV
lBEtLLPvUlDGaR6IhrYc72lmdjeXrdgcCCB2GbXXNfHXYffrfEPVEG2tWUeVEEhe
K2WUKH2OWY/opQypMBR/OmDNejwU2iEW4Puyx6LAyz7Kk20mtsl22ek6zpKn3XLP
frrzcE7QtTfkY+Bt+bhDT5a9U/8AWh+iuORxPGhmK7U2NrEUPf0Bi6UvneZL9zeC
vUb3v9z4fKMsrhdT1G/Taa098nwRuugi/1zaZQeqXexy7YWqDLGv5W47UbYU7AEd
A4l6TWFAs5Xz//KHvrp/oMihwPw5iMrqrLi+/QYskX25Kx2TBabomho4ychpdpmx
wMiQDmympYJx/a/tpVQ+G1gCCrxWhdTel2XmhjUri1G6iWNcuEUK0yWs9G4dwPko
lcVYybw2CpiqboFBToXdkrnwIw1ktRVTbs42sN0PKzvUAgmOOg8KIkGPCt1BJtun
v0k5b7Awxayrt4zyn6iPJBYcCwfHB4VGHCfhOri3f/pF8eJgwkKPqHMFgNbGnZ0v
LEPUMDakDfH2LHp9A4+HR4hsLz1vRu57lAnirU8zI9NUEWyX5/wHfRfyU3hp72GR
YNLU9h9qFXVPq+rXHDglBML5vrwwAGlQzh8YLKKZglrXr4N3y1IX/Zv153tLBmAB
LbZ9eDI58LQ7jI3A53jVzfEHUQ+vl+hNKqd8haJSMFWlaKwEc1CTmnpEso48vGGt
/4AEoNKtaoZ/5imSMmDuUskqKYo1Sbrq0B+UxiFmCjzLhmYjgBmYvz8BjnGb4qDV
l1RO5//6y5poqBxgUYH+hInRmF0OOpsfCUG2SPm357c0CcD9ZGSqYgVfo+Lkiuku
upDoDmdW6Mb0aqpBoFFD9tKlt7q5m5gh6aIW5x9zL9ojk+IjG7papXhF6c7eM7D1
fWCO067fPK+kppJqXqlMTdaULD0zlBT0mBbNLGx+UBdSfMaQYokPFHiN1QaAuPqY
xt7PFpWutn+VvNgCJsMVXhXvrmJU1G9GoBBjEagOjTe7YEFBlboDtYPgq8s1y3s4
Afm7KcRgXPyqDPdx42f/QCRPE24fl7C1ic/grUSL5f9FEuDyO77HlaAkM0aZ2ImM
+A4svV5tNufn7tNpUqeHN1IHkkuUHzC9gdlqgSQh6+v5cG43jZjQ86k1k2RJ1dMH
AQ1tgYS0xYl1ZkHUjRpUzJUluBBOSXrq4c6fB4QpW+T8BcytaqBi1tfwgioFklHq
kQgR6wa005Jr2q3ADSKZG9WYNQ/XBBbOwUHFe1dNnVnqqWuQXE9f3JUwSE95JjVf
+nL8qJKUYgd0dlV8NmC4J6KjW3PcouPOTuLA2MNEAwG2hWutGLRRatuFTRtzpjzm
NZ84CBsFfEwuOtBWDe3/PwJolGzVk7EfLeSqZRlMioRyRHg68HkoMLWU4t7wyytT
bfoVMoy2QnqC2AXITq3tU9fOtFOmSBBP/4VCNtYPPPW++114G2rSlOadrUl/ls1W
zi7OzEh8thnQxiOAMtcMdsauppoTxTS+ctzJ1hPtS7eeV0W+z/FLuCBmJt8pPEK8
EG60NuY7XdN/jGI7KkftrWhCwts0pNOUkXh/yKuDiI8Lk3f0fcKQ9Ba0Yb+z4v9F
u4VMoPRs33nTYxegYGtocp9o2Fr5d9nMMKIopzxaBh/BAxSlucU1dOG4U/3ygadv
LE+ukPwlv8Uklas/Ku0rvHoX4HRE6/Ju9QH8/FCE556diX+njfsAMz3qVkgwaxSo
fik/EPfXerYnwoo5s/k8HwtC6Q3x8hoGlqgDELeyWvgzokLcXbm3boORjgidXUKb
m6gTwU1LJh1R5bMLPl9DEb/9urHsnm1yF61CcgDtdq6n8WZ1mK296rK3ycNDZTG3
ivlJuslCVd25peW+LhUKz6NIo4xBVoyEb1dbTc93Su8XObw2/sd4C9e5JQyq3db5
BQABSapkKEk4OUjRxoRESpKBIRx1/59HX0PXYhDI1ZleHuQiuPapHczbj4WuYf6s
zyr3u+nHLXvCJV4LiSGnNFpldhPs5k5Hspoyl0tPN4KDgRDQ3JCdaAkz/PCnGxm1
dWBTqyyald0/2ywVQVa19uouM4vv/V+6ILFjF7gFJGxV43RaQrxyky7FTijjCuja
1apcW4QVUjvew1hJZ7VyceNqLM1YhFm32gE8hsXjyA/31JIxc9ntR0DipTbUK3ja
7YcPJHuEFB0xZCPtO9XhXR2Pe8tGI3opH3Qe+jzOn3IYUaLPF/FOYRvWIVwuduaA
wzDNSfBouuQ4wHCg9U50ZzZ766HDXQCIe8RJpyzJ4+xt5UdfnWexpAa3Vkz691Ed
3gWcgt1C9EevyB4T7ShivpoXeBqrpU/nMBgIKrLz1V1X+tILuOQwwX+ipnF6UIdy
QyPaYcNdbh0jF42k5u4aE2Im66mKGZXmb6nU6qsODy1WoRgM3LVWGp7j0HNep1SD
ogVy+AaujDMiQAHdY7z2W7P+9eYNqXRj0EDWXNiU1FBLIrjpf8Qf6BS51mX/TQZR
ZY1Iewm9+ZWh+HkyPK5ZyUaKT2lAfBNViCtiT/ACYJz36jkB1Ok2fTYRfddaO7gK
wYL6b934KDpfZNufucjB4o/bC0E8FlCoL14+O8KEVWtpFmMrsipjLKGWXAVCScEB
ra1rHud3Aea3ErhuJWFO3byqlPI6ZgbptHKTPOxHHU/vFk+bciw0GmhKIiyfW7OC
00JyWr+/toBlFnqw4WqrhanRDqFEadcBJ9hR2DylasBiGO4MtGkOT36WdWAWVo7J
2UuZbF+BLgqMDts+BZFqx0tHuAu8XlAPk708K9oF6gLu7UuD+GDtJr+tGJ3GZVBA
4YoQSyfwdO2qN6JlMfPYxhKTD4G4uEO0TqXOdQLCU/6StAYr9xpnpSB0KY5NbrtE
Z/JY1KUwk9Tt8IOvTzUR48GuK4R9um+bjvBtqOwjlo0AaYs9hE0Mr7MDgMM9T114
a09GZo2FOoIva+m51gIg0mkrehlS50KSyc3/bccaqaosZETmm0QVLu8XASoVNgYO
ePeo9FURBRg7m2xG2C7FTxYoY/RuQb98aZ8MsTTqR0b0sJKI/ciGrY8CyMWm58+x
ZIx05A9FPLXAVJZo3+zeNKVh2t8cqoKC4F/SG6zKbW9cRqkhVBAilo/XSwM0TCUj
u6KvmD6t8ffjIcsye+eT1TFszPg/2vcvZqsVqlqfnmGUkG6v1+ui2+SN0Ilqdp4+
uX7LB8nsoJPhuLEQxp2xjz6z7LfVyTS/K2Ohj9xajP2PON4gu7j/+pE4xidYPQam
/k3+Rtu5aoPkjjLxeCR6zgH2qMHt11uZ5ERLH+e/kbHSI3dwJvdmhLptPZvvwZPd
S+lYZTGi96OinmK9nNdlfHOTfg9cJIcf6pD1C4c9nu1WT/MjAaIodcOZnI3Ack82
p/Dg4FftLly8oiqQkwbWXSXxZrwCzqC4N0Aj16YnHPRICPUtdzbjWfbmU4yJ4ncc
sgF/Jm22D19Izx3QAhETK4xx8YXY3hS4tD4qx3OOeLY6jRx5DKQ+MW4fG80YlOP7
kwIaTYSiSmO7R3GLew52ol/n1R+A84fYzvLdRfugrGST+EUH3Jl6NZb8e5ZgPB4t
3BYuxHG39uGT1UQ/tYI5N0ZWHrINd2+CiVR+OA8oaEl/duOEwlS7730OIE/tmNWT
HsoIrQCsbvZhr+BBgrJyDHrdaLv0nVUR76wj+KAybLO42MwBLsq4FgavDrlVDXRY
8Sw1S4NFbPV7lSi+2a5sH8E558dv9zkBqpoiijcxa3iQXG/Md5fQ/7PAAd/zzKIX
enOaBuEicRKgIOsiq6v0TwR3Rbaq0m+iN5l9iWg9zifxOfCavo8HK56Vz4V8Zfjp
cH6KlDeMo0cGgOemL2VjkeKE3ZZYukuY986klvazINc6nzaOU7KOkWzPH0p3VT5s
ZOxWHKoj9Z6YNGIf/Y7xxwQd7erVWyQTpii72+zCimS0WxMZQYe4WSK2ycpd9BGk
XK1XasNP9XLg//GCAyCVz9hyudGKgbNhsTLZtFt9D963vir2OMFFSIsjZ5zzvlYI
nCjHN21acFjys4nOOZdNsL4x6NpBL7NCk8UZf7AT+iqMNYkntw49JQzbTbpztawn
VoNYtSUP9X6Lh9MSDrOLsbcEQp3eMPrbxj2T8Pe6tonyuSPnF2JZIyRu0eklwm9C
3occyWqL4V3T4FPujbNuYrFwEK6gZirxi8vbSIFFGpqkihrdJ5y/38E3Cu8iY4z5
iTGD4IMaaiLSODU0pwtFfat0kvJ8VIoQ5+Yt0ws6U+i594DTuP5zDAI3s2a8nQA1
NVmJMV5e/f3rvvWOtMpaz4p3WHVGb742jQpCOyCouT+KfmZYLT2wldrUFstTGVs8
DdHhsa74E8/GGlUbQtsXorxy8qea8Nx6a4se++TFbXUk9d1I3oL8UwlrqMKqc43n
mlu4IneRCmU7UxjxGZxUGiJqAEnGCHcKhqZTVgkMoLnl5oDSrgwfW1vp5nC8kB7j
hc1OAVjxk9ASwXnhzACaVkPTDZMzW8KlnQ+X66sPE4/A/Ir6e6JZKb8LH6sw4vkZ
lSOWTzNr4eeg8Oo+ZyiTX7ShynQt4Vur7LoY5N9MSDM13tiBB53rvDd/jHtYXN/a
/fOFTRGduBIsOyvcvzFiKKYJ7RZsDZJyztpSsC0ESNfCZ1r2O6cj7RS13RXHQilv
k4kyfSzh6LusCuDypenKxoeWFQiCyE8qDRbvalL5n0RRgOcp5jhEb12JFFNI7l5/
E1O7+Uxtdcz/7YwKrcJFhFbpuJXvqn0tk4C65W/suBMsS7x74789kKU1Vzm+mTTN
6RsJDu6x3hmpV1dH9IFm8+iVo1TtsWps+3sOQdtZm6SFwJ0i5yrivtPWpfAAOmhT
TASMdWipC+H0IFz/W/+5Udm3EXYkupb/8y2cRd9bK0frSyJqqN0JTktJnPrIrwE8
TuPqiijDk/dA3JOwU9Xn02xF7sSm8uEBqRZUkxMmCqbsOaQs8Qd55V64Izw24JTr
/AfWiqAOWcame9GLH3on4KYZGSkIiCMfhQO8OgLSv67Ai9fBBiEKB+DzA1qJxfmW
SNix1Zxuqvi7IUGV01gMzbgJxn7cY1qrGe23sxWc8WrotxfRbeh6yBLE9NDtgkFe
iKbFC9ISlWhgV/FcdlPQ1JwjoLzduSatpnar4irUm3t8/P+bcPx3W6GPWZ+lIvcC
YaRwyEXE0SiJwE6RuH7+ANiqJSpFvwebdaQR2efxUxdZFSu6kVcHoVsfeLe1uJp8
UodaywT5bOMNCYiHAZPwIlHN+/G1DFwXFOK627dApIyRCyVpGUfjKyDijCDH26t8
bfA78ijCpvZ2fol/HGB/IovfsF+XL58dj8vpgi+xNQ7+Z20PQeTTpe88FXLqj+AN
HTyZ/+WUXoStQkmOcLp9oF7kEdl7BsZOE+KXs+m6wB/+QROlttYIlTHKGRTpl5Ay
oSxi0B90J0HKQfc9bJDBfuw3zri408rnDOpLfBXVpw+sV2V5O3Wqic+t+MQFllUR
Hd/TfMD/hGIsdsNdOFuNu6Ff+iHeb86Z3uW7/Uky3QZcfl8CS3Q7RSoT4SIZwhWr
awVyEKKKyfv6G2OlFwlJxQPO0U/7xkbEJYaT8yA/nrhtmmx7RAyKhc26AYvk4pBV
TSQFdGl1Nufe+oVg8BL6Ri0RoHYz+TY8dqVXuq+MxlSADI0/RR8rbqnzyb8LzWaz
Y4/ImONWKxwnc+8tm2Wt1qkz0j/YNVNsYONEqMA8E+1nFw4P9kKvdLn6RPqN5BRg
2WfjHX4GRsjFazJDvm5VCD0GI4qHDxGowau+kHBF8uEYsPMwOcNRitDlglcsCIcN
FKEFiTFWHnC7Lq+TNLmFDUxLN+uDbgxpKiApjRb05s3ZbZmERsE7jchzCk7NJf8c
cDD7cHLQuD3lXO5v62I3+rT9Dcv3OmnFQ+8v9NIV1f4wT5MTrvzo+rchzg2Jx0Rz
I+03r5rp3N6tF7qlwrZ1SqLTiLVvk7aZnYG4p+17pKpMMBLO8qpIA2tYf0zCNu1L
WCjOKihIHD0eK+U8sguNvcBTfnTqJsmDO2e9AUIgRYii1Gw8Mhf++i0+McYrzASD
AgZd2k1CZl63pBJT3XMinpXmw/NKyzkvx/aDs1BEPUlJchbU5ViceCNhfjgZi4tv
/G+HN72Ozwi3+EhWaGMYcXenVIfdk5m5G9sL7qyjgfWgUm3ekqvEkRfVOo2AmZ4o
q+vRExt2y8rplYfxnAJ9CIkZY2tgpXXxK7ohM4U5imVZeREJi1aCnt6kcyO6p8+R
7hF1CgQ729xsuhfCEzyYliFak+FYv4uaE0RbDkR+JpwmgawjFWGE8I0ecdm1Syjx
MZXilRFPOss7WFL8mYQgRrixCEobgH7I3unoCOGcL6RQS2o5IUKtl7gf+HzlI0OM
PuWFd2V+wOpoH7Hm5mBRH2tF+eqVFRZHl5nkSy+MvYVSU6EUX2VKkLg6a+nr3uuN
sNZdFPuk04CDOsABrbhRRphylws+1iBer5+HmtOalRLnelG8mB8Mn0OPPOEobxIw
79U2x6oQJ9AG08vVQ41yFMDsN8N27ulPJHed3mRCkJy0dJMZwT79hZaN1IQcGZ0T
2/aZWP8k89tyMZ0lbrJwcDl80v9SbZZKZAdiGfRdsjTB6+XuJ06ZslFqvKHo5wy0
ubFr1LK4PT9UFq658UL1dD8rOHDryYgmxX1roz8gwCOdy0xRF2WAJURP7iZ3lvaC
wCRCGNNIF4L667F0xU2JiRetGcTdmHQnU0miP7sp0J8OcGytIFxRtlBFh0cg60Kp
J3Gk+dzL7OfGI3Q3BgDa0XSrOLgDEfveEa8kLZztnwARrKmeft5Mr7rkMYuCzD2x
aWrJa59UgePvcLr9prGbYMwAG7JdAyo/gJsh5OQ1QfSqmxpUD/dqtYfoh/irDuTi
SHwSgpo4xbefeGXFLcGkp6aNkGqAub5nVdKHMtrrBpWeXvnFbTgy6LVPJvC597Kd
NIGIYVLYb9SQCvK10zshxD5d9FJEQa+Uiq2+FcCmzmpmATZIKbOW3ddGA0siCwiL
iOsrdwwNYA+pwnj2h/guWuNQ/JNi+jatJXSzZtsgaFZ7i5UDIHx8mj6l6S2hwi36
rZfS+mEcT82bLfJvpRfD5teYA9q1dlrJAdzwpoc5y2rXtmZfu9Ntifzy2QpJQ4kh
RAjOZczFn3HqSbTAJ/fuZaCqbGrSRxqzl8rC29kUaKwC9khxL4wQkgGt4wrLToQ4
dl2Vh8UlKVugyl1Hj6WK4qJGJHOLHefaPiXefc6Db/FPjVk4ZajdcjQ9jeK514nZ
pY7HQOQrWbdKcPrD6dnsNV5BNqgrfn9ylea654bkkxLc7kUhL5YayPLClqTWs0Hz
aF6d73hezEzvy/LSg2JLyVjTCvleOeUSoqGTO27GBlpfypCNA6d8IHUD9xtkYqp0
KQBczJ/TDz8Vt9TkREGeDrUngBhOdOpdmbRgbSIhF25NZbyOKAjjXAhK7Fd8BCeR
/+/tCyQOzQKjTznIrSq8HhtYx2Qk6uC8ptKpZPsFw9DyFaOSTH7pf9+mgY3sKxud
QM1bWlLdvc4uQTQ6TfJe3e4WhXWg/ua1TiKW5v3YJbeph8OWwY4/AM5xEEMtFR2J
MAVAFLrqupFiOWYDsagWV8L4NILHZEfIBA2iT72Z2jIpW2zTXXvN1nna+ZtYHdqg
nQMqnbk1ionyUkaf6z4AMUoeXIWzwcEHLarVFEUvjXzfv+4zplJLmOXqVoBr8RxV
A602yGejyFtmNoqZPAjz6GmOPbp97JUXKq2V8VXekgbKVL31kNUTJU60Tb2eAiCT
wgPp056DOAHIM3HMmZtgnq8HcBgMsAIxEb0bLUEQjFA3ArUKg8D76PJC+bOJsR7R
sHp335zg279IsJVWvRpLXJU9C8ox/AQXHvyeejr7li+5kA/T4HOJBL8tJFaLUS8J
pIP/27z0KNv/A+4a2vDpDEti0WpXNOUv1XfyMqPfW+DCWO5jR23QXqQmqEJ/x4XC
MXFmQJmREW/LYWaxoshrRnNOL9ow2+YEaKB9Q5WEplRT2yodBJ96KuaOrdhd/0rL
EQEkgT/+2JCzvdOb3CCFhSWhITHwZebvYdNKFtxVy8eGublpxF9kC4V7HOTLe/vI
ARJH559wIoS7y37QTPUKbaxgNME26HZlNAhtz9fS3bIwJS+W8sDi4b78HtRdHIpm
BaEK4aiWn5PP/b2JuWMfFN81TDqfOBT/nOV4fqbjzI73w7Nmr9CLMEB6XYSLEmUt
H/1uzKtmzoh96FDK7IUrs+w/fgNLIf0i2vTxdGKMtbywJcfKwx0gAGr+rkV9cb5l
xgo4Q9u8iLemTUDy/p5+yOBbnmLs6tRizc0UZqq/biuX5c62L7MRsLYainidxOvv
cGFwVAYOUsL7RsS3H25jplKlqWQ+wAnkdWXZaoKfpecMJtGve61gBOn3N4f5nDCP
vAox9CCRhRT5aEmz7r5L8JC8q7g1cN5BVpDFhimNd5yjETcXIvStQ+QPS8lRAf1r
LLWspEHUWqOZgqY3VgEkEP13RX3Lo+CWG0+UEgcBszFAY7fq6MHqlRRg+PyYaHGJ
lGyNX24E+JgyAmlcOU3j6f7iV68oCPGrE8Lug48ik6Gpjukwce5oLZSG6FdlHuL7
n/KokL2JmqG2CdPRaBUrUMzs0qeAeu5LqtMsY+tS59y4DKGCh72t2e63/GZTUC1r
VqklisDB3/nnyB+hrfbMHty8dtTIngJoWEqKhBMBRXbezUDB4KOLbnpV2gTd6xSM
VzOEK0HVCQR4FH3XSGzPJj8kmLcv5o7cknvUJHeEFxD3fhljFdVx7cjFNyg4VYAl
Cn3AkLOyZX7TBOmUiro+Ph0b377GlBkZWGfJ2cSrthDPWVMBJUtJRL+Dp4TQLDxD
zswa3McxXeOl4p0ayxZNzge03+rzj6HQaVbQZz8b1YGvd+akPvKLz9sCCQWfOqAM
giS4AJ7hjLJJQ8ushZ6d+nhgqlz/QK45kjRqKRCPxGVyge6nCD6f0k0rlEEm9PHC
qr9p3MPN5gpWn13LC2jtmQiaPLV8XVYjkG/uYSd8b9UiW7ZdfLEicAvcRyB4WFst
HRwlz+cotCX+rLWLiOZHao5I/K1MuRF76ItHBFMTAvCPm9svmBEeHlfBuZOA5UeR
AuaC7qNPqpSiEP7e9TeXn8njCJCgvWMjBE6L6vs9hXoZI67jrxOp9prbWfPx1u7K
fZwIbYZvvzYCdxQRflc2Lwa+XjW7ur+dy5yd6AEEBn28nvtwOOH8J2SSp4pBTqDs
RwjgrEdN0zydGkA+CKnI6o8/lArbjCrobd0/NJpvmdWJe0eFHfCxBHBfpsHfHd60
GbUWX4kslUUp7Xr8RpDFuaDmzhilUdVdM8ifmMgXmfpRLc0kUxPTOXGOlHwKcV/m
MpcLyRCrF+9SoR5I3TFL2/3AtKb2QclyCom/7aSuOzID1PG2a2UXIeV86UCq54aM
8rgBhiv/+qbOLUlScVifA5P7Pd1m0zkJDOpdJSgK01Wbxq/7Gix6vsO0gWGLN7k6
5rbvTK5I0XVRXhl89zfBMo7jozaPb64Qyvdd8EBTUoeEkLEN/vaO4p3VfmExHhkn
5xjJMSdIg9WvDRTMBT8DhVx/aa/xujzQ036wE3B75cW+F3M2x93vroowaDBmlUIl
09UKN6kk9QA2GWpx26EAh3YIyX+DFUwtVXMBHjagNfPGL+K2xAj+oFv/HbIsQJAl
o6YJq7vTCuwL17CC/BhWC+gdlveZb9EY1asCh0CCr2GFFd83GLLQqGir4FH1PKAG
b4L9kOMPS79P7hhVCTs9PjS+0esMrAO1dplOCLCuW0D2UQuSNUCY/Xxic8i1dv2S
Ei8FkK8ZyMUoYZIZN14M25u8Bx2b3ckb6CEHX9z7STWuSkwytDMst0DEZgx1bNSB
zfnTpH0CZEy6U60IsD8PKol+5Q7wF++rZ053ikeEUl9axExt6LWvUQXtih47Kd62
CvrW1zLCIJo4tvBALZvMY6xJALzcaRoGr7ZlrO6T1RrmvBtx53wuX81X3M8y8GcQ
epKQurgN5A0JXSRcSBdSqWYk1CNJ8DBqEwyFy4a7XsVELf9mlpuEYoEnOIZlCrna
nAqw8TFWKwdD1KlysGePiTEjXISmiWq3Nlzxx16jAoCR+lvRNs+A0G6aazPNliaV
8B2EKE0R2ubYbOHv79u8a+buOiOI172bYCI+r7PNMCNeCiC39K5NHEYgdkP4AHzn
6dat71YhOb+AXUNdDewMGlWqcaAK+N3oR8k0isDXi0V31nTPnXjrfpDEfcTEW2tG
UX3KxZmz1d6uAWZBuHjJV7DQxMKQdwIgaOMlMeeAcqwV/+doOpMJn/6AaMPEY3mx
+SP9KnRvl1r06vUrSTXUijONx57Gs05Ij/ilY9j3samZCWz/zkt9SrSUt3ZncoFQ
xYNE4BlOt88s7zqKYu3mgkNJguxSkZ0duKmQKlnv2YoIxMuajc9jUEp4Oaa6+Yom
Qw79J8Shw98USLcflXDvUfD2GLxgQW36jOcB/qvVSfcX4ElcdOo5g0PxGCfWkH+H
C1c52HG8nHzc4JtHU5oV7DwZ4tXB/b9HuGeK7K4fnQ89v8FB0gV//XQxS2wh9kWC
72lGhOxQ5sz/zZL8zZ9UxWVl/SlGDOWNsiqSYUHT1QVCfzACU/6lCA6XjHzaPb/l
OHdxuKixco0eIr2v6Cnn7Lv+A/cBIr4iKNPR5LZzarcc5jSP2HWFQUk9tPhW0K65
LJxNwF103NDMPTdoHXWP0Ys75PLq73TWbeptqG44Sci+L3FWMOksgh6czuOfYBuk
ZI+xgsLrTCN/MdA2+ExhKQwAgUuonLEePekH8kChNKIYCUkB5OM/P9wTFFppcdzD
DHPnET5KpyD8dNdEAa763xDZCvCj8IuiyQcPXBNy/myOTLBrRs954KRcefkFLzO3
IJ1nq2jiT1Kwo6NtaoLXjZc4/X07zRf2LXTlFX1DbD5ODxhE8HZMapEOoZwm9Avr
31Q3Y8iWVP1u/X8h/OwMJNT/gh3VzTcUV/bIjdvy99DfhWrkaUM8TtLkUibfgdH+
YDEeOToMP4shB/yCOp/+94FOQRe1CGv05UbUoXr3FWaWrDOLO+SxwlMKlEdPkFTl
9k/6QxLMLXEpe60ngkmDlVpR6j6H+RgOkLHLf4rJp6HbvjxngHCTOmXEqDr3BO0C
PEMqGJ7/9HeqyhkTYWKXJUygBfe1hGGh3W2aqhGKQGyTZ5mvKabCqCgXNZin+Fjm
UljvgSDaQVlta5jc/yo5BP5hueQeMj8mZL1rCnbGtetQucATnBAgiV2epfzNEnyv
ZovEnSNvwJaAnCSsNo8mC3In2ReVN2hg/aO1DOy4Bwz+k9zkoeDs6PM8mxIiTEnC
qP1UJyrgAMCV//nrxRiDfcNxpo71WMoNS2ynqnR5RGq7JvJ1odf0AW4/m0cZPGg5
tXt+SwwwgaTsjPNJeUJ3NaPnTi/HZVKpiO0I/vC+AFUeT8RCMSUk4bLILikx8Fet
I8d68Nvb/7BQmdi2Mud5ySBGvDNL7mjKWo2euywUIanegxC3D3rSca3IlnR+CZ/w
2Jd7vefDZrT7xVt2AFP6XwMyYfvBG77SxJGTo//P+pJOo9IYHB38Zub7gemy1HDv
CknR6mVE6jFpnghBUE/L1pSnJpjoTZnDUMuIHhW+Ix2q6a5FdASw2JA9SfcWaZSp
jGWKhHdIYFKbV8++6upgoRQSIA02KrGKqKV7Va2SshH4VHNoPg5Ny2tlUGy0OKl4
JjI2ewmIauqI6w4BHwQVSxCaushznTh8NOQNxUjzB0uohplk6tRuPJh7V3d4MobM
cM2fo+gks+gNCl9wd01YZVgmMDjdoW4cuiQR338Wfe76ScHgGT7J2JgPuZP3FRWC
IJSshKnfx7na9BP7Ocim37sZBxvsFnp5DgTuCV09Vn2ZSEV5Xk2B2yDGyKulMXAT
9N76RYBtKURDPh1CaNQvZFZDu+9GW9qpS4qJcGW9rZJuQXtZyJ8B22RobJyfj2z8
HkfEjtYDzWkfVPopf5JjjkS/M9H/n4bctMOsrrPtx32AG7hADHgElYnbivB0dl+z
5Skpgxf/KyDg0JniUwuH/KDLwN3ZChEPRDS9wX7QUFmbOv7zGJlGuPgZveFJFr7V
NxZa+IdAOCPD1pM3Vtw4wcy15WyKW2xmsr3N5ejb/novG0gov71mhxz5vwoJvpZn
l+pLOL7v8upkYDnQ8PpNgiNO0jnDGfXX3W2M61zWYc/TBT44hKe82lN4qyhwQ9/Y
Co4b7MUhROnaJwLqbBeZYBKCZV3zy3aB73LT3QpbvdTgPET+UukWLmBqPBNYRqwj
MbxfevwHWy1G/sRYfAR3sxxOShSxJ9lZkkSn7V12wLPKG2ovSJXFbmhzdP2FCbcO
Aiim4/qBCSAfrmsf6Y4a3i8q61TWscTWmR5982x7k9G9NnfzrPydXYwpVT4vJTAK
AE7DFeuLYaX2Ylae2KVdHs63g5rWa6R3ym3rx7UpEkTCLZ3Bu2arWCXJNS6xHZ4+
cKVnci6R7h+j4kge4dn3jCLdFRd8taEo8woAp1njXM9uqI4U/Pzl0YK5aQ37vqlU
Ve1mtFuKc79gJlRCfL1CPlLgBObJ3/xp+fOyvR5o3EuC2pEnrKTJVhxpM6g4SPhk
3MAb7z6bRJnULNo+VAO9mTSMj1As5vbRWYM9WNrQqy3Nd0Q09EmwfpPePpQXwkxP
0v0buHEy1gE+NJq5pGbRv4jBLYCqaNWqqVkYE7+a4MKc64c/nmxB5ASnpG1X4k2Y
QieGOFr8Jn9KGQOoNlnjwDVmdiRHnGbqa4xmoUGbDuGVhcjJc4TVUwyBnkcRml1S
+hr3QMuVhmwMqBUXDxjhokjLnNVw1x6D1exkt/sHyCtBTybSR0k0Fy26XCLw/6PS
unA4m0X0vGQVrKgKyMfQvoNgh49sr/rhVE7R4RU4chlXXPF26hOm5Gfxd+e7vq8d
+Qmjz29+aj+GYYE+Gxfkz9fGuRvEmcxXAFN0fB8giXyNMMu6I2m8uoK3We+exPtt
fftLqEwohXrDlabDgSvl9ZN2eNu/OOYDqe4jkKK/u9ErdRBt4/Kaug8Q601ue8nY
rRiVAVMZK8baTSv0Y0vRPB0nuOuddtU4N1qdLsthRVUjqtUxHkRyt5O2qITKj/QH
dYgOuGwdX+VgYeTxS7GCqe3rsPiWt3G1k+Sn5aogGUu0IzRzYgSxphhV16SA3atP
jsbvzGEhBCyqf4fjjs3A4yLzcqRJHtEU43NQaGinZ1mkVoQlf1eBx+lztd+BkNkD
paABgr2e7ImY5llCj5YM43xv12lmGyWsjqGTXgT/i8B/YUDrXpHh2O6E0sZZHw4j
KsSqV7Mu11wcwjwvaN04v4Cny2ADrj+IiGbQLSgehY3gZ9NpqJG7SgbvLuxTwZow
u8QLOGdtMfi9wGCi47RpWBYmA/EfhaZuznvoDZly7w3qcDMtEhX8Gu9ax1lCG2ol
0uJMz3IrjpSMTXGwH63fJRLkuRxkGIh5+DHKGuZve1QvK/Md420Z1cfflKR6tztj
XGkhVv+nBfOX3vlS6LphB1BteBXLKA1gayY2daKGC+1iJs67VHo6ciqIs61Z5kz2
I6kqadfVHCkAFgCxiHBH7j5SchMntlz7RrMMjmit2GdTtVrKdi+/t5H52EGr0R7B
7kZd2ztSo4cc7AdrbTyxfq7WayvA58fwOlojkjB/Ki3LzS1qStcsS3BWslo3FAbi
HjY+z5uIwnzdmAZS4ftaqOucJE2zylliyw2kn63/WVIFuHiA0QI+xtmj6r1DMFI8
hHNC2ULGl72BkZjp2wpFpLYOi572E4rtDcKGbQ1o+rBYu9bhfIRstalpSAnO6Do4
yDVN5QWnGSV6Mp3EvOZ/+ZcRnYWrTUSHigoX2XHOtPUP8sBRk4ID6wOD6PADeuWP
m77nFGsw95ei5zlUyr3AYjszgCTKN6fBofTBsdGD38zLZz3X9BPo1grqRPZrMua4
5QeUba13C5TwoDpf92r3IxSQjEgRfg5X/v27rPoDJHuX70oPq90P4UZUh1pbWWxq
fsYXTR5IPqHTjl1zKxxl4ZH94BVMEqVD/LUxmQK8hl39PaggFCCzDgDPUCq2c5Xz
aJzZdDbqA1ub65Mkds0WDFaPexdQUFIlod53OzC2pDeZ3wT+4zuAdXDMp/Nd5lP9
1NY/dPdFNacvdULA67EaY2wwNtnDXcPOnuAMmc+5EpsAbBWgO0J5enxKiQsFTDW3
/0kwYJUYtK6l1IXvh24E/1sjlGI9JrjeptGxAhHazrLtkNlct9O54ic35UaLuKRV
ke34HdL7ED3CSkAQqU8zTilFjGlnCCgCuvwOmLUdEX03cxannUE3yJBV/O2vZ4XH
5oBeJUNmP/Q7eJifAXrqJKKVbEPt22eP59zdg8WCVHeUSfr5A8/67yfIdLJl9hTs
O/od3HEPWUTWM0iicLJUc9KLGu69qjxW0g57pjTZqRfbV8t7QbY2wvzvBaVExCFp
VQEB+g9Nw4blTZNOXfvulgHommgAeyDOSSOY2EKX5PNYO5yxgZY5zo2AgmHNOJ27
7ESsXCtdpmLeLxTpbldrR3o8LQ1DHhQh2q+8kcrA1cMQi1V/mx1DXQTvzIDc/F/0
7PLhkb6pWgLLtSqO4j2HnBRWmdnYJts5CszKA4S2OYgmANj+bIsiPqlVXMHtVKMv
TMaf15EG/Ms+leBU1Sqt/an3K/3XHemkUfsesbATsyENzFRtq/IXB9Hfb74lfM+B
/DPXkBDyEFZHlhiscpNCEDTKF0ggVv8yP7yIxHKd/QvRVe8Nqfq72OVr6+a/oH+4
Q7FXVpwAeCV1FHMRYauK+6bSJ+Mp04njO8WMLYds5juRZvY7UtW2kc1oShUCEWTH
FEZwdLsWAxRDuaisYFfbKxfes0XMs1CbNzPffnBjcpZkTUqvOgKn38is1ebzxow7
5Q0ua+U0PYJ8wXrQztluKYkc2IuVpVbTthN1yt3aghXFntzZbbDx1cix6NtHswjU
wDCMaXeMqWZVpHNfSb4UZzywaYDCdUzFouEY0bs+H9cP8vkdSHVS9O39Y/so9mUV
MNfTXGOSwpG9C8BpxLu3pC8+3GxSbeQ37J3iMjsL1P7F0Z8OXLB6u7RfwbpobHPh
YSRc05mzQV8Bv86dhznYt/rVlHr2EphUtr7nQ0A/QUTfC3PvXuHKYMLyYgNvi/M5
exv2cbHOKXk1GGwG2I0+FAoXksH7iWcBXi9oh5l65U2YCxidTF0lDNGrGw+kTAtI
86sS8W1fS/ex8a4xZjgOVfX3YfjLzZpoT3NGkt5QyegSe0WQe330zxXwmvpE/ON5
KKPecWTY4Bi5cVWApKdn0jy+6S2n3914v2IHLW5cxxixeWaW12qi21M+skzqdrtJ
qh6MBqPJy5espDiYyY/+nzA3t3g4Rp7hmTPmmH/T/K8rloevCCI2e8YOUJEDmRek
e1HPw2EcQbsE70ekkd6BSVEerozqDqwQ8DsCJkandON0gZahBjRzToNhAeg6nDHk
ahrvQyDe5OHLfxnk194wbUwW5G5Ejaa2vIQYre9nFhY/51Tw+QcBpyev703SLwtC
Fo98FmSKa+KyP6IPJxEY2IqcA6x0DRmsE08CSd9FjniYIOLD1NxEGW1PdDBP7O+w
cNmj/mrtkaArc82hkgR9os8Kx/eU68p9PhAEjwNoZd5DAjt2/fLNbaWTtN/KxUIC
ixA8Zpx4HRT61sHAbRBqjyZA6tCoKXl8cfq4gB0rUgGEhsGGuT3MmM5pi+s5UTwM
nAj8+7IDX7Zj8RfCykSZmSkIIWYQ6lfww/iwwp8eli3epUVP5Ai9G4Jva/mT/4Wj
9JUewi+bFZDshaW+oHk/+gy3B+iC8fCXlcbSpvcmRDPUImPTpSBlXqs0mrTaGvpr
YtsInDou3eCiCZqNWncxCvW0rMRU+AuCMwFiPj9z4tulPneFWYBs2OI/cXmQwZaC
o1LZkk7IsmhDBUaZx1qnetRvNXpaaywGzrn0Idgsro/rcbQHXM/dIRcyMZzX/LAz
To2SkHYAmEULmTU5FI0VH1p4/yh5PWEP38Thng9ZWYIid418GmhbfQuh+BeySwWc
cEFvjnxSLaNFuf1kBNPZZ5uWtuqi7LYePx3ybjJSA2gmxBDOLPmMzTvc/SxuL7od
E9uLsCeFZ1Wj7N2lI6Dvhgafs+hNJf6XENRD0IhcEtpTFoQ/vpmK2LKLLr1NQ7pW
rXw3s2VI2T5OpEtelSmZWKNN6WgjyXBlk5BvOqNuVIEQxi1vJkvDxeBkSeEsjNVS
WUbKwCJNAXTnW00xZhApRqIgpayxW8baY39/UGYnN035vl2RqnyXqpwzhWkDd5l6
IqgHEqSpHr7gKoucbibH7H2jyIs8AXMP+S/fkTTPqlQVI8oOQxlCX3NEECZJbZx7
VwFZiE2hGl5k8VPAlUMSdpWvLn1PqWS3p29BW4eKWThF1TSUjkTceKi4oIyGbfON
JdzST1H3ogstUmG5bN2HNbUJhJbsWI1efA7on0MsMEajp00r4I4KKC+ttqDo5FCy
QeZEOJ10KVzCjkHkoY4lZdclZo+m2KV1ciUo3ENslXsvQRXO5tJz9HZD3fSqURLR
ZjQ/BlOaAviibNLesaGBH01DGApsx8BTbwlJJ6Cou6Ob5kAXD3ZE4oy89mB6FHR0
0+eweVJsHOK0AlFOCv2uDgLWfgAScAG6y6PAm//6gY92wvXZtXGBTwdqIOMYktzj
r02E4I/XzyIs9aOppQkEtKMoV4Mg/UP5YEHIcupLAZc1CG4cuigkyHG2UJFeOwdD
kZmLoeIO+ZyoWMs42IleEo6UL5ZMr/InN/dPRYiq8z122X6vCofS4+wc3L/w3btx
iUXxfKDhIdr+f37f26hqU+ZXawLiRGYIeJQc4eXC2Su52u/CIcNG/aC/PjyTv4AK
0BiB7FA4uNAOpDWwGZIoSWdFXhc329KApYR4LTa/xECznnYAOxuI8ld3xWhMlaGB
L+46aa7T/9tU0LtUSOqFf/skGzulmc+vsN9hXU+y2/u9KmZpbpmYhxWUL+1PM5tk
sqf+sSxMovDMUt8jiF/pn4pTxU5BeirR//1ik7FDLF3KuaBj2RguF/0LfeK1J3sI
EE0wn0NLeEZCCaHHKWJO73FF8drlTByHz+Fjw38XM1NC0RcfW4C1Lfy+kELu6TQt
lyGsl7drZwT1qojxt+EA1kZb85z8Du3hyOrYUAgvU7Ses6DI938PfF3s5oZEuSnV
Fmwc4r/s5H/C+zlWFqv0ARUrMq/5jl3OEl79disAiZIO4VfOsdhGp+myVsWaBMD7
ba5BRSGVR4goUXabk87NohdztimwJAW9TkMv+HDQ1dovGlhlMogwdKGQmaaJ8KV9
YtGx0hOBasRK/b9I2sEcCYmS+fhPQShSgOALkEh9/8BH2GItQr1bj4Zly9cvX0q4
ivwpDV1ic4i+1/in2PSNtsLmTwpFuYZSLHqhaXv33oQpdb27de2hT22IhOsWZqow
FXkLJdo8ZZyGn+c/QcdLmUQJxJSheVa2fGZbuFXEG5yoQetg2a1QTkIJl0O9I2MN
40smbxsBtPgnaYF/kxD5iCIlz0/IfRqlVnGDvIXVVVVVeLqqD7Fl5vem8Xc8BeJ3
7PMJ8JsGRs6gr6gi8ZG1mWj2qF6dd3IW0Pt2iucLXZ0hKuQNeEJ0vXQ9sfPSMiVc
gkPtF+SXSO8e/fvwqzldLcMYpmUhB/sM8Zi8QvOnVh7QVBXs2UWfZEfqyX5zAqUH
I1NJkG5Z0kB5A+/pShnf66WtCYpQ3fksdJQgK02RKZcIRRy0PzEkBdw3OjFtr2WY
35RYoc37xBevEZPlNTz0+LbwEomtSYvcHawu70woaxZM0gOUToKPssvYNU08CRMM
KOJIJX45LXTamfIVGjdh4pyEUYL56wG3if8+UE41PhfTleMG1kC9rg0SP7enkTNA
ojUeNwfqL5OQtD66QCSy5bdF+fv3/bPTm/zjbGtUVXOBabRdfRibwe77z9zYeePV
cdaFAlJdjSS6JSZyDgK7UtBPP5x7xnxWwLJkXaKHxHUVhI4g3bTfv7ry5yYuWntR
4M4ZhLNgeOGEThmomHx4STnL1ZbiimLyBrq8VQYOuBUHEDu4PBn3iztlAPHWjKG9
hyiWgIMQitVlVE8ejKqspBcEWWGdIJ/jdHPWozYppEJk7egqTrQDI1ctAxwtJKZM
iyRsRQsmhtsSS89nCn0OhJ6X+9uP4V6iEQsP5IEMQkshpLIqHjvSFc1eKPOEb1FJ
4Byv+KOcMCUh0k6GHx0t9z5/JcU+lVpD1BTLtpZsjo9soa0vHqmW4hygrWbR9Emj
H6srZvvL7kyMfs1q07oE/xzOM2zUZr7s/es+0U5IV6CLEv5cEmWij3a8x/axow+J
cg90Bf/WYNZJzm+SvSFmA9DvpPCMTFdKoJ3lAEz50NPilDH1vFOp+w0icr7Ic09i
UDE/GeBmadfHp89ZzxR1ey7EZ2xvvmjBylSkqnH4xr1I5dVMjvsuBYafHWNXH6TP
2zF2YaTmYhyQCB5d+T/65Dfi99/LaiXY9uWY3lLO7YnpSiiCmLCC7CBsQP4E8ViG
EiomVX8eNNuvoalSl5CjWN5/PR0KBdczso474Onp8Io+BAwC0RW/koVurgI/aMZH
pA4b3Y7VkoQCiC75EQGGdCgvqdmwvTpenD1fW9WBFxpGwOzhald1LBSoKe4+QDZ+
YdyxhWAzPEyF9kGKNVPtE+w2fCPm5H3eZGtokQY9eBkX0PAkLxhpuEf4BacIjPSm
wzAkH+CPbRU34RTQPIvnEZnQ1DRdfLc1xHWbctORhhpUN8LhwnVX7dl2bWIzeW/y
YcIr5HR5XfvsGC2qSIs8UpKXdn492wd/Pu8iogsaT70T6W5xh0xj+uCGr7ofi+Gj
Oun44sYxsjBN3U3D7atDB9xIyCsPyiK2hG35jKSAkJ56ISUwBMcea0KADCS2QVfT
rf3tzfFjhBh058Z9D3/iX7iwqEoqcVmGfULB3TiKngctYaeionIncl7GbdUtg9IS
MnuD5k0vfY6h7qLObIrPuIfIlRIGQfz9QrwUPR5SEnbCA4F9lN+JjISoXuRnQv38
+69ONQFzRDMvlC32lvjlgrytd5sJWD0WovHQVdqsbmekkdxinL2tOZH1Abpy5cGt
s3gMECGHZL7R0mSvpAYtz4TVauyafA2U6S20caI9rkK7c10f8fR3LsmxmOgDQmlE
fYjWkO40iyLcKnICE/Z3q/+InE9cnNFUCeIy6TyzsGm+4T2M7rWbLOcR0VAUUJEV
AqB4vd6mn9AwubMabvhUPzw8WKupeTJl7cIq0nVJAfUvQ4Qnbl7g2fYzAvXgcgXF
o08HWzPYWKnoT1l5M1GrOOoEGrWSQ3IKEdCCCM01L6ENn3NbXJzcvY8TDNKsBCgi
fE1XYBW8vE8JLgGSlx1Uzr9/af0bq6RKXbFkPVy3621YyWLLgMcYELElm2aaeUGc
92A1jaKzhB0aOdXrfHrc0wcMkP4I2nbJM/TCUodWvRCWn50/rhmzotEzN2olAJDP
ki8L+L0UZg7DgcjQPLcUmBGj8fa8etnlnba0cKs/AoaLtEUq535KPtraADMV+yaA
CJ+IbOHPmpRLvrbRr09MOlTvAQVjrveQlWhfbmnBvzw9ebp1OniXWybOAci6ZSeS
oHu+ppkY/UfnNRwzEjFoscUjnx1JHQ+ORn3AhxMo7vv2merIQELJ0Ork6optVQiG
ImfSn9hx5haEiTn7eUSPfiaGdIuWU9bMMnUtWUlxvvOe/vLEHNSefI3BkWfQS5Xn
8PIb2Z0+K3F3qDHqXvqsjh/rwF+ycC3mSMwGN5KbZg+pKcLVQ7QRYEuO0ZC25tmk
AHohC1QUnUvXR1lwquXX2nt0Ky1+JkrfAcFA2wM9+wsoht7i70ndCLGr/xFx1/gp
6J4Y0vvDnSVZzRpGLuNckbTuuewld0qe1Z2u5qZMzlsISpPdoUPqKHoIHBNI/o8g
Pszz2TSf1mY0esvBmMVoYy7obBc0vNw2P9Zpwk/1rZhQg7QmdJXe8TH/6dXZzFGU
XEJNkOly/5v4PovN4ctCEdiTGPWYesZR7sT7SfyzlrF+2iZ06ACT+mUtZC2vgBCG
DfbHsS7lWhAeELgCBUswOlgjtKrP/ViFgMfJSubg8vjT8I161Kyy5Q0nPGJaBAzU
DHo7xFLEGu8JVtSwdEWJuoHXP25pOnXUXQv765H5onyRXSwYp23TOxrPzKFUh/kR
rJnpOb3/Kl+p7ab9gTnwFzkG0nod2nhKZB7F0aYrlwyofgMwNTM81vLRZc0lJrEP
Ysd0EOScG8imQWTrQkXhpDTQXxMwmGj1wntg3V62ZKkZ8zOWaoafJfu8HxC8Xb4G
VNiFc6L6UyxwMv0KYtQnVHPj5F2hrIXZvYVgDBoeUMikA6c1kbSk18Y/owEM33vE
c9kJOaez373NtfTqc2uEv+hVCoOxYNWIzpG4n6uHmyvwIdrew/q9W4jl05qNrIDM
LbwL6CNZKhH8y/aarvUvGbAK9XMJwuzc/tBgbhKGr9HN2/YeKGR3jVM4Ghv3uLlF
mPSjtS5XPyoDVCpMhP5nSDYtnGw35pj8IPpvuEmvaRaThLqlMbYy/pNuC+N1r3rl
8witaeqRltlcbGEqvTL7teBa4tJOo+I+MlU5IWySOAABZYxf1Qnb2Ip5kHYdNZK+
rBGiDAoKUh4F7p42UV/vekzvArbo1WYapDrzv0vowGHXZIaIWUqxiyNElEOSm98z
Y44ym9FU5NIVM6gRuJzxe+fi8k4nHhKEnlfP/v37boCZWHwbToJXDxsDMQGzWB1S
ZOGcgfCxQU7kuZwoGa+nhqL6QQX3eA3OqrjMbx/q0PMTYxqapWYPsdU93yETzzPu
+RG1SL/q8wXJPaW50G19wltISLMNZUZCVe3bTl0ZHE70L+ypvGVKFeQzzOZx9Daq
1DX/aVV0jHmbMC3YnQWkHTRyfmhFWOzKD0rOdtyQuYbBlDXEW7iOqfsEzhpouChO
a8tmPZfLlyeBG4ieS7KnePd2oXBX2COUNwwa/8k1HmcNJwpy37VrXqC+uTuBK1n5
DUciXfs72bYI/VZCEn7EScNXyf1ATO7pCo4FWmCZDD2XtuEZQRePLfHltXpw2yzn
T3ff6uVtYrs1ocgxj4H5vIphm1mdv2vBfzQ+cGbVL3V/ieG0+3zS7xITml+4Y+jP
Oo9En7GfmfxjhMBkoNIvAG5CjAmT0TtVKKFsOUclWtev/FGlUAFMedCtyfVGoTpt
8YjGAhCKv1uv1lJGHtZkGGGniBF3021mXZQeOMtXTD4Tcz3H4atZYlKV92QSDUf2
5k9aS7OZ8UlQAO1/V+Z8NQZ0IpYfKJAMRgRIXkxbehKufx90ZhW2tgvrEvZ2o3TV
7lrKgMHGx3nIefxRfULnKsA4PmuNLK5F9cjVQLHp05e3FQHannJjvpO301uOv5MB
6uEsQlQh0sufaXYVSLZSc7nfkhz74AigVtx4yTrVvSCISe2vqkKezNEfLAR4abXi
AyeeVOIAOBo01XPvUTRDcpLoNf4D3uXf8ydFOFDsjwqwb/Bfht6Sh8c8cd3s+xyV
/YLHY64riSI47BjwsxHcT1iYJl1UxyvsBPyhtmp+GSb9UKH6erEZHm57wJXUZumE
JI3jxX6kRBfNrcmvISHsW2gdieyGu+Ia+VpeAhASQx/vKXYtHIFXBGIYFX0NKyMU
HLDrj/WQ/YjeHtDZf4Z+5E3oV+swmac48xtU744WV9I7pnq1lOgU4vyMn4yy70Ik
m5+LNr9TzoSUATMPVObWCNnp4UMNIcwidtrArFfJvOkOl8oACuGC6EQq1AM/Vtf9
lfMINLUwMACoJ4bw/pub66zOiP4lzji9S5+gj3gCa+wsVHlbn2ApvLZCJ2giVbL6
TS+ZHUAdpYviR6U7aKhK2adRUr+XEm9CnJSAMURer24lBrIp3tbkXG4Vzsp62C1E
6S0aZO8DiDTFkuzzJcIMlfrvC6XhnFyxqPixNIebs++JbhcmNVD6f9tEBJ/xx65y
jf9PRu7cAtLN4yitgbCAZOsuA+CWGafsYONVyq82goK9VNasVReSms0KeuPFnim1
D0cKV0FNec9QLNhaZf82hirH3z+uk8GgqQp06KP3JL68C0L7ZJzOBW/9kzaMn/ZH
y9LkkwVZeJvEAZerCEbnEE+9mylPsTbRHtpdEt4/EYtIXCb3sFlf2NdTpw8w9px/
Hq27XNmBL5myvevdI7U5/zRhyXrHYYH6VbvrctiKt0y6XK4lJZJxn3h4kp8onqwm
9bYm2/GOr0bPRrBz+L6nKQjIUdR7oL+Ro8HS/kU5TmSFY2HEQvz8NBKOKz96oLou
2l4Ht4/Oek66hs6cu6+bFdvj1XgurBHCKOu6Px/v0CtRzyQqQcbiItiExJK3CFJo
XPmkEQ/NYh57miS7tFDf7vctYYL5iZLp3GVtGntOkhxjhz6872CqzmIfCykuGLF7
Oe+TXK4QCbo8BPgk+W3s78KnUsIbtqgGCFRyH2g6n/TvYGrW+DdJCSQqO8RGz5HN
5nuiKuc0x9/xLCcio6tSqMVVKhjTUiTRwY5grOU4uJNRXfqB0seXhCx8D2Bw1cTi
1ozQhqhis+ToIA0wG56uZ83moqkCsr7wkANZ4eDWIkYyAHj7JzTzanK35ILFJu/T
mX/z7kO0x93e1WSYn3mvUsUxHaL+9cEptUJYeDvBLgtyHDiMg0995xaca7jmpWpU
ytJFltV7ZVoJ2VMHoEdgmMLth8aMMgP+ZdnI9c/Of+t+qg/T33TPUCH+zgZD4X53
8arqz2ZSrCpohLvCMZQe2KjNMs76ZtMQ01GQL+p3rHjRl1qQV7+C4WhZmgqCecqD
T/QeNXiQMsEwd7YbsavD3vJuK+nwVluYGEB9cv520vD22AoFFwug+JZfgEzgSZJ2
qfDW4UhMaDUjLlM630p3d4DDhbT+yVxO8LyvtrHHhq9ypmzsRk0259u+lslGOzqD
9Og4xCif67DbUGwHqZY1AflTrf5CRkiKo4QDkLeTaAp5+p0C/kaJUfYZ1zfPdRKk
ckwE1N7hN/rJMJSV1GM4iakHvgPkFLIx1gpOMvG4w2OIoMtU5yZ+eyezPFAPFlWS
DMXu7nLLJgFJRxmx0iVSuoBkb3gX1pe2XwqSyGDYZCjpk4DAq6+Yz1aCAKzcx2Xz
D2uTbh2UKXFiDpar0bWBH3MEUmPVhQXGZY0oAdeZR/JNaUk1YqwiFlpD5fagF5Iy
xkVVlEiuCycxE+dppp9auZwrJ3zwe0AcMErC5ILrNvojPFLCNZM/qr9lBK4BhmfC
yMV5lHhg6oT8Au7tZsNdQJ+sGyordJYSc1z9Kq7nRSqO3BSIzmZpbHUhDT1SCjLg
pj1fnZpa/lPcksA4uq6uVFCr5GZFhj3m6eF18fq7SDh+kS3xFDHY5ecI3B7NgS1b
bO+pNQoPZW5fPMIQwASNeqjm73Tqhhqku16SxPfR3w8JSq0VDMRRVhZYnYEOFURT
fgXgVuYbgA2mEVdFcUBLWagaDaWH0x2hD1qieXTu500/aUFlYZQTi+obIwvrxk8p
nBnSkxysvwrdoTm/rRcEFPHt/F0oqSgCz/FiWcW1MdLyf8hgWEsEaWsBjliwUq6C
SDXRM0MXuJjbc27tT4YeSxNVPTh2+ND+LJdrcqK5+z4ldT8mV/MEP6hbAnIZivfa
RP+aVcb2dTpPj/htpUIo2jEhFrA1kC4I+T7K1s87HJ2YOAno+8yOq1uA7lng+av4
7yDcqY4opi3wpq1xXJlOsuVvuSqu6YDnrGtDFfGubWon7MoHVQHVZaVxNMp+Xypq
6tgg1GI+ei22VYM041slX0GrrZSZKJNy8rLrHbvJvgqDkbNMQLeBnZA16ULOFeft
oHR/up10HcvvfDj/aRrcGbEhthPdL5XAoINPH/PELh260m+MGqBQ394PBiSsC7IX
hQAIEUP2zy3w+e3ezpzkBsCfK0N1bg1hlPl/KpLMJNeD0iGperEu8jFkXr9sAhng
PFhlxES22oPHXIraR2vCgvco+/zCf34zhIbXoqMh7H28ovBKCRV7OFZ/hDDxAG0G
4BUOSjEJudTiuXPJjoc2nqYuX5sl1MtQdoa8mQC6bjJBbNxtOAyRxF7YArlK/PJ4
/J/85Y5MXMQOCRRzKtQF1HZ91SrZkuktKn26ZSKrUdBJ/+WkYf9ws46jDxOvCbtp
6SA9ybSk0uTfDk3aHLqmR7+VNJlkdhXOVHRS7O+hhW+k9GlAN4iIOA+7lzQZQvaf
kYTu4DWCD4dqqVysKOYuiPFbfWotH+FLyqjB1TnG0X+8sH7Eq3Avq0RDttYJil9D
vJXhclLnDme2oMc6MUUHGxFcMEC3SsJHqhB999DcD+5iPqHQmad1ZJtm2ArWwfsU
6wuk95VSMulSKxq5lm5KHjUUVM7u6FR4QcOu2uTOmUp9obvLPbnHeLIEOW3DpESK
CYXFnFia8K/WfKbQzxHwbNQdSqR22IFWjkrZIOiTU0KxPatVONdIITyd7zUqHmSl
8w2L1ljWXU2K+CWZ5cagfzKflGym3U47IdExNqSXPMhoD6fD/vCwS5iCAsAgWJBN
xrV2jPY9SnvukZ8f+5kWDiWXiJBxVJ2FXcPWHEJ4hZhC0OB/iLVhVa6VrTVNjXib
IRkpdzVLppqSnqJk/HF2uVZkU0rDNIKaBun/PoRc1EvZ1sxmy/v575jp0OZZZeNX
+RQBnyUeNXwkg+FQc+ffARfZEtAzYr9YBOrIVRWGI/a4mromKBbXSEl104Nnq6by
mZCjEtYDmC8w9ekKgjATRLdUvqq4xkl4NOY1g2XATAi7DYALNdmRJpb53Bt2NfaU
oOMP3t7I0pChD+PluFX3J+1/7mh5wOZpkGJSb7a7h9Tzi5ebuUoYG6aYSqdjAzU5
OVaZ8plscCGXOIDDaCgq6hej7XPyU5Cp/GABMiptYzbPmwFpsOqItxEtFt1WCMLq
442HKButKH1HLB/faAUWR9z/1hWNkrdDIEZXgYnsjDHlu0Xm3eL2MvJGN3C3wzSo
tjjwuaepDFtCHKd8utjzwchkVQfAr5ANT7mgTgQSH3CB60HmpOhnGS1GbxFATrGE
EsVznGQxAVbYktRYmsiFTI9VRdglKmhFQeZ4IKs5TI1HzHYQE6kWysM/+C8OszYk
AGOmIz0NmTOC6M+KO1uUsAWyXMXIQvZQmM6ISDHcW3jAbCwiQ9X+N7HDEg9jqeuz
Mdv3G2MnYvn6zM0raVyIY2tQ5+GcFIbxhJdouSNE/36e39/771Gz4MEAp4O9ae3x
FNriZXEgfN6GXv1Bnvs5RLwtUe1bFGCPD++O5hcSaApGWQRH5gcAudwwsyTbJake
QCkIICuFlDrax0bFDCXKWHAZnudKbM2Sn9npV7WaOH7RYoU5+JnVW8uxmXhlDPY+
8C7hLtj3kJtgb6PwUHwwYRwb6uQlRV43YTiD7QARI5DhierHJnzu7WiWW/pIv2n2
AQFt2Y7am+dyThCDkVgU9UN4nLK8PxSCqDiu+q1qX3DZa7p0xaIOlZS1vYHFeKzy
Nt2iy3wfu6GBuHOBEuB11Gf6w7DHD+0xpJhzDSh5F6jjDsC2xwYxguuiKX8eGWVp
RY+mgKkMKSOEVajRL0gTv5bfKaLaBXlwmJiotx1ywciLCHsHmqUnANAGSIBqHs5l
7IWupbVZ7YMrx4kUIklH6bw0/VkuR5dAcu3Ms9QwkyxACY5b1llInJZ57YtxdnzD
IrGxL0YPxpj1eG+aTMtSfTC0v9zzKWvFWcrTel2NGeeSa2A6EM++EYYAmTfoBlPG
omkNlnJ1GDdO6tRxj59mZ5sL0KNQcPvOWkjIeZ9mO0gjR84LKXIW9sahjsXBudHk
hdhMKWsFDrZhkPAfEIcKSHMAmNzLOemmcH+hAqXcSs+30t/RhxmYy/a1oQSTj7OK
4TjCO17t5XTDJqR4AYFulW3YUWRo+YpvKWzNp8dErLOBjJByB/+To9sUSqWo0TcS
wiwK/BEWgo8lAfMzgIXOgMSv3KTRnam2xguvRmj3FD7h0KzNgVs4Neln4Ey5Kx4N
kC1t1FeD93j3HSx6ttJoGewi+CaGL6omhHFcWG26tsD5hkRACEFPv36wHrSXrw9V
jl/Zvj7Y8nLrhnPUDRwgeZ9dDZ4usmZu7RJhaOyJt2izi3IP+wim5S1IuaQNmHm+
d12DJ5MrwVtEqdP9WnHE47LDufTeZgHT3AC7+5ZsaFc4rRlVb3xSKz9NIakFHIId
crPbdQl1QE5tLRNciD+ctNBngLyd/RiLAO90jl7q7DVS0z9fGvSMlDGEhVMB3bMQ
WVJmx8sfMMTmtG44MbtXcJ//L1tZVh62qkfdTd7yFflOZ1/DnLYZmuLU+1TIWHT3
PMJtTw9RCr47MCBRvt56bhwlULGgd6GVMBuGzqyNV5KaN2KTBj7PySXYwrfBerZD
sA8sm2Ty3KnvetX41o0oH7LCx5Mv0GGouDmSpnZ+MhnABLIkj/B7EmxK4BDnv79L
YbcfF4bqUJaymghlUb/saiaeBzgJIGQq+HxBrnW5WWcCzBfoYN6SxhKd//owqkwR
QUpcNtX/OAIbIkK0jz5jzA3vPH4fQ00h8ugd28gvdAmNKyY0v1jBo6icmpFyFZoA
XiTfltS1/5AxC162jxdrtxw6jEVe37u8fJv89eNeBkPPRWwtd7zo2H83CiYpmhYN
4mIgucIEsidLoPcjqA9L/UcJtSrk2EQSgODQnWAAQFAo84A6HJjzpNVEuP0hEubg
ga0dQwFYXSQe7Ik5tcFr61QBDxQ4nsrd+hltfqU1d7Dsp1BBoyZwfLdnaxOhD0bW
IYoKx2ZMWzLpEdyW0bglpOQHqHXhx1shFX6WgaQ7TToaJN0DOmNQ3qIdgSdjEdJN
DFBs9QjYFGyDyjk1QJqxOJgFyTl2OpRdwFEj1eCx+MyAPat6TPJ9Dow9chBN6Tlc
LnelEVubPQ5DVOA0nlyH4sepXF1roX3DNN2wCO3apuWUbbVpUoDpLGoNd++dIyrX
21NURnsnExcOVF9VidwCjwM7m2grvQl64e0vDIgb7wx8JunATYB3/Tv/BnHD6Pjf
3Uc4QNlTOTclGUufu+/ke6oQQMeeqs7HA9ayEWXAZHTlMI3HxqVYZxToYV4zQBCY
Lge6YXpYagcQewNu+q9VQ3dh5vXlhMTiktsBWqXUqgl1ZImBkRILetSMTGEfncDd
la4Z5RdvZwqXevZ/YZX4Aph1HbWHeP9tINtEFM4x0nsES5ohuO1XtEYH2FTdU/WI
9aW5SXQsuQ8YMDijousI24HEaNq4Whoj/YrLDafojzjl+bBD/vJHhmnSDgtBzclV
Rsb5DAL/cBYeAwT/q8BB2c8mcbBL0q+OztLJ466yvq7wmNAD1i034DQ4DILTQScr
yDz+K9Z5ggD6++tr3OMop2UTB8yfQgJh0cvtMvEXmBHq5AjWVo9sqebrHfEOh3DL
laAUOaapU2L5Q8BP0FixfncKweI+cAuNnDTlgdtybPOLVTJwtcA6+p3Te5J+p+JZ
On9hhmyL5LBAPlMmTY1l7tc1elYTDpDqSF0NOKqPjFmMQnmGDC0YLATWYmgca4L1
f1CtS3jbNF/EIAfGBFccv4/Nzgy5D9PP/fooOxYM63ja4MxRf2OpP6fXLTKyY13i
mhMEIAQ2rIJA9mMTaZWUtkHoNWQpd8kODFfP1z45kZ4PCW0OlZ2RdW0xMrS7QXty
5sRQRKypxDWhf89BClWZ1Yku45tPXWDQu1C9jF/hfJbRtg/YovOHosGDUia+hBSW
GHWPGqgTEiUHImGU8LCy8UDzPok9oD7Mbst/AlMjrvE/Q7JD1zulmOvSKfPJiz7D
tdzUjED5cQlQjrX+wk3NH/tN8a7nVAS/OkVDPerz5lGE6wf80VxTEXPs2X54qCmt
LnFClS3je/kFStUp7TmsrGxn2DHAb3K0PpAg2tyaI9mKoR/JKyRgr27jTQXnuNHr
gmYSasXplMvCxkzs0U/1SeOruFVht8wZs4K5BBdtk+/2v7AvW5DBcWhlwnHO92RQ
Q3IkvCose6lgzGyWXw+11t7Ry0PJTXEsWY82rt50k+4Hcdb/1rGd7RCGPr7pYC+9
V73jUNJBhMJ4StjlAHEJ3JSQq3VSzZpoAhMEbyopU/53xnkEp65WOdAPTWfMK7KM
2FgIEMmw9znI6EzAyxDAPOptGbPdzbbAZKq7DCyqdnrRYDbgexOxxh/4GO+puXao
u+MZyJ7THfZbncBgJiwE9bwICsHigaP2ym1BO6VT75xSxQd0p8pw9Yyp3Sn+q5sT
2/lwKx+cJKQ1kL9S8jDe8KuKOqI1orFP7axeyJQPgP8BBUBidaSRGpIGqKaBGQCJ
ufMHbiKk+ijqMd9FVAeq3A2n1+fr8mKg7aTJs/6hlxRPP8vm7xUrHiQ3pbtA5lsG
IXu7hXTjXmSCHWKZfvMQqG1gsELNrLSiFyjXGJU9dFGRmGgaymMFcg6MTYZFtCPz
kUtgG1Cb+HkO2uH/KrnEJ+pHRqkGHp0E2YzPG0d28OVH8DvX2rbyO8k/gF3ATRfD
xS1I1GC0LJLGmYGiqGm3GFL9tTmFwM1GsaI8EiY5wMImEFg6BXocUo0CXd3Or0aS
OpsBnWNRMJ0/cTj1kHvJmbQTiT/TW5ohu4hbdnv8Y+ce6zul3Sey7BSbkCm+9W0n
tKyH6yC5XSsvC5MwMk5oE+KU0scEJAox0EpFxyeWxaGNt4lghQWxDgO1XXGvcpZD
dtOqT/p1AucVU407nnUXF0Hz/iAW2hD+0UadWP+CWl4G9D2MWlrxTs2sTc+Dr9Cm
y7M56U8CJqHckAy78WqrEpLZHquK7+Jc0bQIvPpiWmxFd4bwc07rb0pI5aCv1K36
HEfIszbn+jqo5Pv8MBq0sjiWk6nCXFEsGYEz8idLN4AGHTCAKqFZ51W2+huwPpjm
bOfT8XxlUPbqHRNHhT41z3tpRSAkP23J7VGC5MpONshYHTpQp2z0f7fc06FK2yuZ
ceXZwkwp0S3GhCeZoCglcSH10YBJp3/Ik2NWPCWNbTt5s8KxjwQ7N43ZIF7402/j
SDCHx5UblAK847eCrlqvuiZLMMC9pBEAqd408Uum7mX1Eq1FJ30mX9PAnjmjN042
EuO6st1gUFlrBjjxF5UnRK9xTeKLlxKcMfgqryg+I86u5FJ6Ye62GzjdcdQ4NW8Z
5ojLaBhVTuFbeBE9NqsLHQT2w+IvXmL+lC2PhRt3IL0StM43uv0U4beXSmVoFoZy
9KTNFN0xXOvUC9zzWDEMCHwFl+sM3yIy+2VaAsvt9/EaGjIZG3fsvaYkG9bCuz/C
h1nkzmgVouRpwoou6EynB/IHQXb2MZgmxKlgR1o8Q0BDHywifhHG0iyzJE9xUZQh
mHY3jIK+RCelh3ufQT/qTP63RI8Rvakvt2jIDNBmGGvHSHr4Iz5X7wn0pyliH9xN
cKPw5DlAt/eORfjoYay7TnSbva91H+/YGNGSfE3p+sS9VILpiaA9hM8rbp/USJ8K
qHNpmxR1SWQykrimfuFB9n4SOzQnD69JWls+EvzHrvWWhnwghF2x9XT2s3XW1Lqw
5K1zX1sBt0RaJTZlZuwOxKjFimWfe0nUQsrUgvbsoQaAGyiHnAqhHLFX6G9AMgCm
8Dckbluny9ZzfghXbPtTd0oS/D5vKrr8R2D2ySFLH4OwLmXlxoXICGTYEaj0OdZU
h3BogeyC6XgII1Bv+YVmhaOQjWSiKC5Fk0A2obR02iygY7uYzlO0W0KL3aiDtI++
mpSEDwVHKeb9v5dSfkKc7MQc1Zaw0Y9uQqSxU78whTKL44iTKwdOnJZ/pT8PU7Rt
nYIIs+rXuM6K+347sf5jtyo6efjQqdxJwRV2SIYECR7HdygaW+cGAJsg6BeLHKMs
5/HBqpZkDH5pB5BOo9FxH3PVKmeqUrHXHGVT6FmVKzpSJs6ag+IOYzeLUtUYh5Vo
G5FigUaIEk7cTt5nSH24yTRFC9LO0NMH13whz+73rqVXxYceZZIXaZEK8vC/U4Fl
gPyomO7sYZZ50Zt2QJGXTawDsQ42uEFOl470khVtY5rD3GuXxmlYHQIC9zN/AJTk
AHkxXTQi208qexyNsi13dv7JGkTRIqiLapmZRFG+avsxK/aEmQWj0kVtn+Ya1y8m
zouoI0otspJI8srmD4OJnWtC1thCzlA/TUyMiyF1vf5ghenxAV1rElyaZNZvy1XO
hCBPsnFdZLifMj8gpf2qEeijvFU8zjxt36AH/uIo1HcmCqzgbuRfVKwEkag6LSJB
TyI7z+IwMBqVDXhSWC9BzEeyyMgalygdw4x5aXVdL3yMIjcgNXHJR87lQp3kyivu
uIrmljXJdLs9fzg3xgDqd90ARmp2j99YKieyYea05wGZy/u4Pe84gpvnnuekwVFj
gnRiuw7tDw8AiyYxv5rSaRLQO9t1AL12GD71DF5lahOXWDOxHTghdhJy8GHI9t7L
MZrfTmWEul+M9sVi8g9evFKVtRBFBAXgQ/es/PK1hQ5qEyyRrVTiu30fYvGhg60t
mKM/h291Sey1LepseVD2l0x5BjrYJ8kC9oT5L8UBdy6AiBq3PHW96NPmGu8/alu/
HQNrj3CnPMnjvaNQw0xYAMWveouzDelxUb2mAICxabYhcprym0MSO9zo8MM993Uo
LE8T/JGK1+TcOeMfS0h5PgLcAULy+sgOIxxbBPup9ghzWLN3zYXI3paxkm2fuWKq
gQtbMunumzr9ku7g5NeF+7mDJoxRfJaFoa1dNsbf9jOvOjZ7Z9/33xZJgcV6ETri
NCTRNlkn6W0rOD+ISBxZ5eJbKfdRDXrvtxA+B6PEUnadOjse6lG7ys+sp6eIzVpS
kps4eg96vaJTZ4GsIodDsp4mwL/CJJRpRoLMgjB6lTvXYsMR8896s63zKgptXiL6
uEBrUJRwmcl8DeH3jxmwf+/K1wJwUJtJoMpsDWLg3RLgg1ll2nQpaqu1sjEAfkCg
o3NErByNy8QYmjFTpos+auTuaN2xaH6Qigjj8kSbo9to7Vty8Wfw5DffuYXm3o/x
WAmEZSUTVgheCih3JwO9yGKaXHWZxBi1NZF2z7US5A97FHXZ3FtTyo5OaGwoKeJR
vfiE3jbR/G8X6AvvT0nW3t79vyCm1IidDkT3W1kWn1t1Eb1uP3iUt9yV3132jCS2
tvJwyvhD8vMOu6DPBnLJcTRcoazZhLeEayhji32AfEqUjTR4ZbFroYugkXWV+pIl
jF8x8tP7YlWxllT+nQ2U1a7DJPZL30wKUZ73hmKLT/vjLfaVhaAg4g+gy2PPyMo8
GIgSmkm/mgWdc69dTBJci7fVSq6aHhOg+xngIwNtjNruYXPA08LPWnL+Y4anag2K
Uw7VCA13iTEsXMi7QkWB6GTmcteve2ZKd7cPdY2vwYWNcXD6kLD5hgJhErLOyfmT
sAuGcKBO0Y1Ar4XaQOft0ZfFB/wFh6XlHAJVwjB1UAKRj9T4XEpw4xaOSarLIY2O
Qv7VjemcUfhG2qh02e9MZE94+RC2z9O1++fAn0WTA3qOrDEJIe4+3S3g6klr1+Rt
sz8f1k7Z+OqLgN8ZZqhdWALc28aL3nFpVXVxCuopk64KU12SxXjTt0uLtpuup5T3
uVslKgVgHzf8L/xXOkt9H9oMpSOTg0Np4HbEDR5qySvmXmvJmGerDfSC80oOxXxa
fDeAQSyQSz/Cw4rRfduCUw7oIUKI7DxWlwvAGIKZGBM3hStIVY2xwVlY9Vw6JlVg
XNEk+UFGPOHdsxhMNj3vBkov8dRCtuRjyr86pENTN9Fd+yXnjtdqyP27QxmGM8V3
41kGW9FfR35CE38kMmAxDZpzJaXH7faqv7XCV586CELkmMmLMczmclQMeg41v1iS
hqMFOFZ6bT4POD1UeIAiUgzzYPd9YnYdXu53shmFQTMWZTxovkku8cRf+bT4Vwpy
Xtc0Nz5khmKhNkWDztTZ92sdf4qr1nDC8KQR93Jo8LlmaYkTkKVem+GNG52tVTgL
VQh5b2CoMgXEnm51F8YEZW3khHOVc07HsWh1kV79BvxCdXlscbuS4tt6F1dFY4PW
7XGBHbw432i+AwnqsnMgf3Uoc7XYZrjqggKrRu3InYRIBgq4SYG/Ls+URfHFy/Ez
rwHRgn7C/ZHk2HX6KMSg3kcQBs1AKda5b5ECaR+0tjGjKiYSRWgYgpch4LRlwhLa
smTeGjy9vXE3zN913XlrXhRZqcBY4PX90wkIxc+AXKF/RmHTqKrNfhPc7CJSXWYH
zLfh+WsPeLhbjblSVL2RmrN5XBWCtyA6xaDuH+Sdj59g9gMygLQqpbrQabO/593Q
rtoY7bMRpvAdMzMXzW9gK5ROETmNlBNbNXx0aUsQS4Fepo+9k+PWwElR3ac7Upti
HjF7osEkg21xcHHmU4G9FcPnrPiA5a0fL7gN51WQpLvfy3IAl1TOtS5MSgjBe78e
EfZxAC1xFSu3ysnQnLpy9LyHY2H/+VtXpZwBNKnqK2gvq2ummhbeh8OHb/PLZEee
+w9OOBkchgFr9hRkZz5pEnIFUTIhToQONhDZ77ZomaM3j89b6Mt+/cOxZtlymKTu
XxlJqr16sC+evLNjLlRNhOaPaO/XX+alzwRoB5yGZta0UT+vS4YOts2ogvO2hjlV
Hd5i9eBuethAFE3cfBzPnCyMBQvAw0OhQLzUkuZIyylhODy7Ox3eiuV1ECtGfry/
Y0m61ytwEwhW7mm0SJLnunfXusE6+8A1mZX+yE8xjPBgdxWig2Yj7/VgPJgKZmUu
NPqAQ+vPQHO+z+r7jyvFE21Vg+2+by1zjQsR2NEtZoQbvl0KkXfqg/c0ZEkLgBsq
rsIgGnjzZaCzI4EGaPV3SymT7QKu9a2Q6HcEVkbBgbIc03icSPqtNE4IEfs+vhxg
3wh3WiuB2EldjzEKLt7Tv62XRF11q7xNDEnmSoa3OeFKFKpgvhH4XID8Yytcp8e2
SjzRtZUoXQ9nJpW1calMpKzEJ6k05L3DetlQHCTF8AorED7szhAfzGhGabfCIknt
ooudKkLUg0JOsArRXjnFos1LOks+ODDlMI3hpo4MZMJQCydbOLjo/qpamsr6jfbx
pElYvc/QKa2r+MTNhrwLyZGYeU9UJQ5C5CQWl5Y7fcpAmNIQAlZ8MYGMbmknGjlx
A1bueDBz1LUCXacQaVmaGMdyR6cqbfiY5AS+865Wt2Kj108HBNEfGkXFqK63zezy
3vZb/8Xpb9n8lDwvqM62/JbQWhKvR0twkxGFIyGAdmFAK7ly28DMABqAqBmqRXGD
zVSmqyTyT7FQ30gdKZ5eDSkufKLG6D7du3UQcMM6H6kiZlif6pMxDjobdjjSQazm
SmDAHyRMS47kuymRGSU+f32oezTZk2Ox3RNgkXirAslo3mLR6G3Ou3pacnwZ8LFH
dUul1zUAB4qdnxHZquGLvEcQKd/YwZdAqoEDCP5WKY+Blpyw9fBu3QQyvbLScS/N
7ggtIGNZo4eXxrUtDjnlWNLvBT+xK7FuUKceTeWzgV5UsQWsA3dKXixCj+BGI9m4
s2I95bg16J9VZjT5GZ6ERPAVRGIWSiGU/ad1rAf+ErMxSBAueMpgbYJi73Xs+Nj5
eqqQVXc8Hrp90+96Ylouz0knMCB7CX5HqsOc68R3TSrojEWKAgzhLfgFbz4B3/5Z
qd+lNVCDzOtO7L+xnMHy2kZCxu7PhJ5VNz0jHALNe2x5rvnun8qdkrYHXCDSMmGM
KPcyNQ3A5ChbQSZondsY6Z8vR0b+g5EKJreLTyrEbJv1vPvOKgbwuwuNKhXSuJ5A
Zy0khyreUK06FDwk4FN+8GKtj48l7TV4m7uzHPcqEP6oRxwBZb+Al2Yk2k9UvBAP
5mJPsQVqqhKwrcsVTarsxSceUeYbR+4xUFUJkufDgEhPybhmIjHLyhD0n4kU/ATH
8siWhKojwI0kIUBHBOC4sYrIG9ivWxWfNXaltP0BrjdMn7uRoYq2ICuIdRao9Pds
F/eGnnhlzkgoi3QjBk3evrhOmaGCUIub32lwh+6R8TqMmZbFilGkOKT1fXh9em0V
tpJ5gqbtNXo7v/23KelG/f0mJbponPuyskJlKC6YA9aCu2tCfyXizgOjdLVHftnD
coy2GPw08cEvSSt1CrvIT5XAWmNbzrro8H2RB//WYtelGEwACRNmVDTjPPDegqqO
7EE/cUJTRJBd0SjBdHkSNdVUDV+LVWoP2fE8TOUd6XhfVf57ZlD2mNOYmOxyEimN
KTjCXa+JlNGroieUVhbJuWH/WziTUnOobF6g9xjVpnJELzmGZjHTmfV0hqWpX9Kr
u1A7mTMuH7rSo25WDKW/7+3CCBSJB1Q2/n7vqsWYn6A40HWDhD1UBvpPJcSLnA2o
v6BR4EXt062PE1KpsTTWziNJc7CA466G0FWpuWypontqBjdER3nB0+ZVPfMfBLQB
TjKxm1c6QEFnLKL5uJFkWZRwrBTkDKo7LV5K2YdgfVvApz59GUxUzPd+FhAPGlHO
mfbRhA1yNVmdQvYDxH0zwbNDyw1IHqwX+dzVc15aSXh0pR4lS1kAWiFklSx4NxjT
PeCYmVvF9TJ2QBEdgJA5oSbNqs0v+B1z1Sm1byYHfTcL+9MG/SGNdIpQPQaOTz1h
aBkFbBlMi5Q29RX8tZz3zk/mXg8qSc9BVoUWVo+NlmakdBU/Ur6E77Hx6LuFyV1Z
LlYrmE6MjzF8c1BT9FgtZRHdiBSedRxOcrDg6mQN8Emmi3rzrHWzfsURF5kFAWsq
Zh+9TWh/FDn5m/pPrnRSlQ7/YH29d4zyXFMMoWpPy2f6oF+cE8UvSd2c8B33DTyM
vU9SxK5/sFz9YNRPIpmUUWDNjNncR9UP2+OAGzDfx5ZrAJnT3z31ZLcpwf21TEpY
Ol2C1hyH+zhqlfxREUbUyvtKEfgbA5oGasgvVx4nw5or8bK7/cU/wHrGF7ZJuI2t
AjOkFCQ9SrEul21k2LfQGRZQh4dm40PNPC5Y4U5y+3UmqhhYAHqTUVntt//i7pTr
N+hNSZ9ahxsEqet4FSHyTpas3acRW3HIks9jxMfjm43U/DryQt0WCafHLX6+B7R/
TaH6qhMYJfebQLf63D0cLRLBhAAFGPDMpzSxeXeVIj5wywrMVZMwW9/ECCcon2nv
xL1CCOs2q3cgZBWJluVr4/ijgPm6b8U5/TpiFRKRKnkg2AmdZZwtWEvwarpGwp+j
KjZ4EvlZjFni3bmIaA5D1Y2IcTRGUbM8ygl2U0+SpaSnUbhx92xM2LEauI4zbKGE
PM6ZlCPcLbwt25GBxdDNU2AUP869tsEI2GGoKn2Mm1XLrGwn6PhL9J/oYpNsrW0A
rzn1s2dSmj/PkU+g89HqwGc5IE8kmD+xJkfdFdJ68Z6y+apVwOBnsY7hPJtZBhjD
GlFoEwNkE3bsSXALH5v31gIJD01Nn6p+RosvbV0pxTbyUDxYhlTHXA+cxdb3HY8k
0GRjPovpRx+m2x3tEvTrNVRDcU9qIacE/LIpZbEePT5agFEiFznl6E1SOo5gzR6c
dkVi45xEC5fRaZP0EUpb/esEshfhdkAguvkFp8ysGMe5ReM/oMxdnXiqOYBv30a4
0I8yCEP1IsDd8Ak9GQpIXm7Em3AmkWfuABfGhJ7qqk2JSpZsgFvNJlcaOeFdPSHn
OFn7FDRRubWIBJq2t8ifbPMgl9PfVDRrbHn4/HT1m7pcf+k/Y2QD0ukY27NzymLT
gTk4ijGa9Q82d7we2lb5DxK95hh+gVJ25yWLszwiEbAhnIuuo3xvoDGlwrMt4J7F
/6gB+sEOpe6VOlY5REJfjRA4b55PkuS5Kfj7/jM1f2DKpbfdeXuPP+hMqqts6nOS
Vzz30gtN67c3LCraswm9XCAFZmbfFRrKjZkpobw3XfBxgTlo3+DrmhQ+GtaO3nNT
/urpyFm+QLMVyBvLxuZYvZyodH1vp5t/+tEbjVP9SqH0mJmJ7mOX5EMFtGqgftGS
W/gBsLLWnsFrhnqjYGVxr6hmscQrXp+wQYGWNVKvFZE3Q30DAQqQP/eKANv5V35c
mN2sG/0O2uYB7DD/P6K3n3N/MheGRc7wv1k4JJP5ktEPOuZVDszjNCbm0ndKPYC0
btAkwpflsvUtK7vPAUDlrUigNp70ulNQa04FNqZ4IkAsaK+YOgB3CCA/M3E6D/rb
dKUIzpz/FSr21MUAywsGF/Age0F3hbMIVz6ySPcZrxeODR5qGbvvs4jlJ8BbLoCu
QBFQGWcvE+/NciaDAn9Tl/lhy83G03A8C+sHqg2Lx0qQQtcoi6Ycyciza4CKwF+l
hg8IZgteDhlOlPal1XWeQxGwLk91jzTJWwSeWuANjURLUH2MAw1aVfKwvaWHk+e0
TILFocTHIN1jSbceB1TS3Mk5eCJAMkWH6M6pkwvGJvPUh/IEu1uDZnyQx+xicY54
cVdO+ZI4OEuXFVdTu1RGN4uE2vRlvQZnRp8DESndV5J4/l2uWfaJR1nHLKQ33FCZ
LmCzVTyTIX0Vn8LViEOfiwpyngoZ+SKerfV+ekBGqGiOH0NrHLZWIiUGikVJ1iNs
GtkTn6JH72O4Ag6nux06aGLIWrIAoUw5lkdcTsDVYYZkRyS1G8mtb0a3lk1ozEoU
plgn5gqQy40fDvH43y97vDSJzsEG4vVar3wfZMSKPEZDe/gKOMgjNBkES7TyFVip
5mwB81UUlWKYupgSbrCF5uUQCV0utxp5Vw50HPv88fpnxZkXymc7uDkYNSIJRoXT
fk9fypQnhqzJxz10Z215xnFJFOF26FEKwzO6te7ZdTkmldoz+SScLXiQ2XYUGVlK
vnKoNDn1QAIaloaSYLTZGz629lGG9uQXYiaYaCxj87jUP25QFsvwa0LnzgkYd3ms
O3hJenCSoHi+NDuCiqUV6zNadDHyXyo2fXXirXkSv6njO19Eq7YG3NdJq9bBj1Uk
dxczY3MwU3T+KLzloKaGTWpwfI3xiRKPGKM26s+GIyq2QBm+xvcHoEgRZrw6CYvs
emKJveFqJykm4DF5gf1dqk1CtJB8zq6n7VWPnY1o5sWfvTCPR+HOO8hxbE6kX16b
IYNEEO4h5p9ZX+6YyBg63kJYU+InddF4JzWhaGr2Tp/w9nI/iSAeFH1e6BnWG1eR
aryfkC/iaAEaIcug4lCCvzZ3sJ4pfEzPBsfyi1UAUIhnjvgOEuyHj491AGqDJbjK
xBGLTAhuVfqXrhbJqsTZYVJS+KeZ7qbmeL16oSiR47rthQPFFi398Ka5aGbTiAQH
8g/B/P3XCNJhVkwd4WVEgTgbfssQvQo2Fo35VT5rLk3u2DkiEqpmAbwmaDKkmAFc
Y6hIpx3lS+2awWvuwjnmsYsqA2OMIwvlod/1qi/g6CVFL/wbRLVg3RW+jp9QU9kh
d+0x9YpQKv5gXge4xXEzEpe78tC5JblEUvQgpjY8QRUnKTlB4zdud7XA+IZ5NGI6
yw1XjORRm2NjYmy2GrEtePY1gpkzl4cqn3AeisowktPnzsCluZuhckQrTjlFFIkL
g9Vdi6Z8GCJf5MxsXTPMk4etEQB5Gi8N4bgn134hNiTYeFkfdRKHEXqgi2+H/vqV
/i36uiDZFsyRigdVtxH9ObQ1Xw/jocb+UZhRvP+rN+Gbpn01YJx0xkXMun1UW1MT
Zlsjo8N3iaKRkQ0LUceH3aAlMCGGl1MPAqCP4oUfUIEktKuZBcur/Khfa1YSr2S/
YalRziUYq8Mmoodp3H54jODv0SHQx9AwIaGyeVsmVzhSkm4Yc5HG2C0MZKuTtjlm
tr+EXeM45/maaMv/A5au3O18ybX41N9cmHjVrMukgwDN97i1IH1DbizCn2ndAIBa
26gbMN5vYffxfnURAPDwfRYOh2ILH7XvHuRjXESte0o/XR338mT2BlDNcFTYSmW3
n85lshqpeB33C4jVnDq4E5xYl6p8B07bo/Q78JCG9rWLhwPz3ranAngSHc78uauh
fKEBPPCXGxDUyJPnB7nlgBMdsPCD0kXMaK7Q/fIGhNdRhRM7amncimi7jYaNiCet
X2OovcTlnlJ2QAoPbkMkD1fdW/jKpy2rbfd+3fV/X2CnO88EXCw6I0Cuh4Nc6ASt
6X1ekg/AW7/HqKrwM5JxQdd8vGE+LMfQSrcJFpWNmgbSyZ7cJtSHkb42dOTtBBZp
sqPXK9/7Whfo+SgE7g3fV95wMeq5r1+5coakaiLsquQfufNJ6U7GcpXaCq5vrpqg
MMfD7BFAw2AwO/ehGv33c1/cV8JuFi/EZO5XzO5XvU/CqHoAqkWEtbEUyTgiqUnb
GHQPcrNCy5oJWV71eW5OJRG38i53cuFrbODyd4WZWnwzmjGh1kcpLNNlSpxx0sZr
eKXLoVxx4CE+VFmEmWFjXB3i+HBlBKm+pjuZOqLJDzaVKFHw+eArzK8POczGt7Fj
e8z461YBMKDMbjsIAnRxqPjYwmSYEfq/eq3AMSUf4+iMqf1LPKp1kSIYMCg7uSv6
8hUrbukI0FSaMgGBMsFPQE9HoZ7RzyKCXPohtoDCp7kCTj3V9ELu+EFExsddASCJ
yARx2jE3jX/r3M3W+wVXvlrFeREYDf0Oh/qtlPwCPNHz4iQqpSrTtv68Is567PN/
/NqVFduTVCjqRhdGdwuoVHn4yHPf+myJnkkmPjksGEMZXK6I2oTJ1t1ID+2E+AZf
RlCDOqu1UbJm37Dm4pl8Csinqk78drvAV3fof6g5nPMAiVknDq5HPnNtBBdYsFiS
w4FdZa7xlYqHeXNUPSpCkHQSHleG6gOthuR2a9clnOBm7vYOIo0qMVnsg2SOioNA
CCIfrw2SZCVBJez+QBWXjpEWIwJpXUr69x71CENNAun4BoQ++++goclVTdnI9UAD
nWqKJ2RkFI6ahXj6EsCgQSf+SuosQtwEPp0etO3oenbWkM1AuVT/yT5x15UKrXAg
KPPNOz+8au/M4rTWQj6VYg1SkP/c9tAiPOP9RR9BuuL4D2I4IBJQ9OS/RypoAtfr
xRSLRmrB0XyH4pnrH9RlK6A1C4B7/AW8EhcOXS4k42T2RVWkSc34dlKP2x6xzHpU
VXj2bpn59DAp3wF7Oi/w2xlnY67E1bOenK+C/ealXtZciOrhTK58vTcIRJ6SVQkc
f65xmeo+b1uGiT5jhB4sOcyZ2rp4LSzork5+VeEh9A+HoUNh4t7rEAsieKWZK3bK
Z4JCIHfjKfZ3fonFPbe7AtRwFWG9fit83znxUawj0v/Llz8y3YcbSvquDIAcONlG
pEt/DASRpM2DTBjo2mJh5/U5y96JP1E+Chp8nbue4g2kkcWyOfl7XQ+6iJgdpWDB
2z+NOxxvkzZxqBRktyqLo5RLFVYsFy/ZoXbVDOcZ2YCUooQSHS6w0733X1zyh/CZ
OvRfF/KYPuX6CYepdzFStzqlqRgndU9GR4DYQjw7cekA+HXfjdTIKBgnHl9UudZ0
S+HGIFJfeJQJbBcCL36DSLFWqBKgMeQgdxkZHnGic1BOgHqvDek5K1qWZocTzLiF
RRLae7YYtgbwfN3nZoSdwOg6hfvkGp24Nb6LOY7h5SVoKOHli4nCNA+hpXKzinex
nKYfdmLrVHdFknrPhRIplRmdVhmveVCoyI6d43rGssBeTOOdSBe7bO1sMxHJZr//
pj1+f1GsRd5n6pxLSNoaR/XZJFJzbQkjw9Bw+TLvNtfAlpQhndjFHLBR8QvjvBHm
l1B/T57O5dDL6E6xqLyp0Z57nO5CXRSRN7Za3jd0d4/xPylcM0mR3qvjnVkH6Wj4
W/xxtGgczh8zTrQKrrGoKwBJ+jt4TUPfl7dHz+GUhqwFmaLAMEhZxi+IS4NUmx3O
fk78U4IF2dTEvelV+8PGGBm5saCoiLGcJAK4qVDWF3rPBB3N1G1g9bFBK/FB6fGB
h8Zay8N/gH+7kwnbFnwcRWJyTNqOHLytktmt2+JvXhckHL8XjEiZ0cBIPyvFmUO1
CjV05ceyWmQKryn3w2c6k1647NMSPcjC+f6ZVkKkwBe/W9T/ysabE6uuN0MnNgcR
jToem6SJuQeKph4j0ldWoz9PnIrS7vwmpdmAf6dQqokDkbduBMvrU7JXlFj6zU4f
nLUVpUGfsh6zxHptV/bhTkV1EI+yqpJepcW8X8G5pnay1R6KStxQMwtuKpQlso2r
we43F4grVEGVw+SQ/KpFo8fEo83gMUNy+GDalpa9DkXnJgRTDtU/Nnbh9vLe4e/l
ux2loVEj8lgFllwRp0hiu0iNENmPuRj5QhCB0k/3ejGD1Kc3rO8qIhocrhpVGUws
JUHAN0TKGZ7ETp0BVSU0sP+A2uJkVveE4HmWkf7PhR4w1ev6BOlzK4BDUo/iPh8g
xvBCdizWdayCJ9P+kTSBHWkpifW+wxiKKQyGP0BVsR3M6G06TRYbtDYRAa1Nxp1g
dOwtj46EkAH3bPDV2fg8zCdS36YUpBNTYTPptd5XdIb3Zmz/ysRehieXqmLRXSnQ
b5h1drLzlVCugso/wpof3wbBzhfnaQiMhbAaLAya+gktELsQ7yZlCzHLG7J5Cf8k
q1dmGWcYb/useo+farugbvqd64041w+9iMmwTH5PSMD9VE0IqIqxi/pynPk1+cP1
LInzun+nCNikxC5EjlhDcGuukCgXQ6VzExypgEVQqFEQU+sYG1fE48infDBAWZrI
bYGaGJdCYphiMdC/iripG3Vbkymk2qdieYlKonJWYsc5RxOuPLe/XgOJZklq0IJV
KM16b4EqEJKqUkxw5Z8Pf8Wr2dXD2aEKgGro/gKh0mjWJzX6u0DpgmB3awWIOVVr
UC4IvUUvBXV7qJ1oM6ubcIZzv+QarRVjHgz9U7Za8EPYDDIeyNckdSa4FMYPwpNz
gWZo0VZDAsp3bQuVWi0W3vq9B8kuf3eLf9NrDfl+G6mCSmffRJt/1LL++AA4DpXQ
DZl0fQu1gr850YoBnXII74Xq5JTIMEjI/ePtr/feotBodUcDy/3Vugg3uZhJJqaV
knHMbsS+oti3bP5VDSWnw3yAH//YLTYNeUE7kGJ6WTy73ltayLHRTFO2QQL14j+y
SrJiMldFsO0v20MrrcEZcjOiWe9YLmm1wH42mloG3SsW1MoV4ups19A91HWCy6BU
hKL3gouEIJLC8sYgZF21So1UNYKDbOdNzv+AtlyUEfb+P6wr+nKNxj4WnMmgFoYK
6te6BMg9+Cpa2NjGS2hkPkPSqIfudmn0QaXIk4FGYdkyEcJRDoC04cgvhZ+1Zutq
Bo0kiJfHsgbuKEA5+RrxUzFolBaihU63bjNSX+wbhNtcDBQPL85aApQiYjp/HFd2
ucBW3xXrZuOpUgNM9wK3vv1baJwUe0IXeXgHkObQlI0mh5NZS+jc0wrTP/sVaB4J
XYWGsNmeqvbFIZMSMgQpSS1kpyfwDLgTqz4ZpO+t5jWQf2gH7n7EaVTjgHkgo52Z
70OoIqACN84Kzm6qJbN9RidyWBhW6PnHCYrHtVlHEUm5nLukkcnND+9uR9sDh5Rq
xqdmwv9SSkklY6ehw4NhaeyjV39ZZgbvy6Bq2UoXgytSzjSSoHWMSZDhNXrmyZ0l
BMSst0qiJeGN+gfpalo+XieWhMYpxe0Lb6fJqJHFa3OcSsGUHH+8Rnt8K0iYN8+I
wfgt3m1YOTmPuZCyl2g6rsYYoHH8FkGIFZm+ylJKc63AEMK9zFBERKCgrSqsf+U9
dU0acv1O6zg9ATU9PI+Ntn1MYc90fywonpCp/mp3iVTpnE8YVycwUzzEt029pnh2
lvnxcokHcLYZg608lCWnexsRzGI1oPNKA2L4RFGltl8mMdAfzlMt0eBx/iBqxhvW
Y1V3+JNl031DEarpvzYLKsaWe+DyEPtQ5DPp7T9hzsjjxi7iRWaorFjFRP51RM9X
EoqXYbc1SRAKZYpFjWYa8vgqJezcmL1+L3cTzqBYhQ/ZO3i6y2JwcyPOJEGOtPm6
C1KzEJOIl1WXsOdfaz+ERkFFKjCb4cdd51X118vIYIYtGUv+jdo7IKeiTQasd/wc
KI0QyakmgWng8BJ6lFzZgJvKjZV0EjTPTL+xL6BVUOKNOc240lPk3YIRMrKPagO5
ug8RVpavI0poIItXJcR/mwYYPBw0U69TzfuzDvMd9lL5QAbWSWexNVdq8UQjddvb
MusOaJI+3iCaE3YkslOpy1aRveSvPJ6Z9tuOv2SCoaMAoGdAzcla+zYKzrk+gRFd
E09hXl5E2Iygr1ALONqSucQL5ypv12Rik0gtwdmCkqqePl2DfT7vU35ZlV+W/bhM
3AqSTSPVuOXk5aJIYbUOnqGMgqBFhAYmGWwV1VD0tEsbyF5N2D6Foc0ikT+IRAp8
0MX95F4cZ4u15E+7dQrYAEmDsyCVESoAhiMQZMrdKryUi53MtbB55rTnpFSeN4Pd
dqFXZCQkZweVMwkcj8wQaC6Bf7itkCiYjKoa5/J+j7SqZ3YsMUmtKkDRFxwHK2Y6
jt4hwLwf2Wuzaz9v/8FcFF54Z6HSE8IWeqgIh0iySUMrobSrCtVQALE2wB1qobpz
lVrxT7zItjj6GpO6rNO+1NnqyW8wl1QMPf/EZfNKz6Oskygsua2YvuuwG/SZ1ecy
B32FIhR8YCDeromWCQtm83yqVu753lrifspHIipd7kw2Hv7z0wVRjYyv14jFENYZ
Cd3ZOC9M6BAUzI4+Oy+bhSchMr/iEg2Yg9/P3Ia0RZ3rEGegqKbRZKuHKqURGpcE
feuoO7U4YUMGAVpElfFnz5Ln7LsLwln05ObLqa2yv2JZh4ObPp4/JY0+qQlduVnV
AlEjpK7/4ZSINPkHK9LFblXxKstNqSIzifF8qwiC5sSGQo7h+g1t2/GnRKsnFP0N
gmGI+L9ddbrK6OErt0O10FjWCaKv9unPW4qeQqEXKawTapp1Rj4L2srV4Foz3OrI
2qf5m81+3Y2GCaQ8VCRvcZBEAn4HAd2swkzvV9NKG/ebNiBH+3Jxhaqn6B76DKpJ
Og5BQ31HzkMjlyTM4aLO+cuH23wXRSSxlgiL70UCBvKjlP39JSRNkarf+Yn9mcWV
ziJgNVIc0fI9Qgjj316Ps48/m0+/1a3AxAEsVBCWBQXUWAsPFAETcCxE53VzlGY9
BXdm0m/oDKJgdOe3g2LG6+3RQR+bclxWVrEwt0STuYNQ7UbZyvQV1vGvkJXFAq3x
EqVrbC9CJOhuBvpm31mbCJE8LfRVd0rnZ6iM7Ex2MjY3wI1/EUUv/i4BOr9AdKQJ
LSPl8dqH/CBExUQva46HJgcXfFUR+ti2YgsBy2xfpO/f4TCKn9XMWDumO/VbEm2t
EEjfscGnquZxndTwnQsu6yA2h6tRzwHNFPpO5xRlMdwsj9TUrOHTdTHR7MtMloZe
11EcNF6eCjhBNPU+1X7fVUUntXb9k0AvB++GtbYgrNkdHjfOFI1ojnYf7L8Sh5wZ
A/vaI1DU9eX5ipoxbtMueKu5ojf9ZuKLJvoicggHJi13swLsGxtpcLcKtDZmE0Xo
aQc/29JCG2Nmrxql5wVTacR4jcj/Rx092a5+TQqeqWmlcW6sh0O7VzclyDdT4VUf
FNpHYRbZ4/BHtiHzNVxI8n/J6yzcw37/HK+n6EbGLIkkmLFLrwNzxjKinqBJYLyk
tCIlAsRnSIrkEqUOM5sE3yPF/Xt6re/MMqK6EC4W6QvracUGZpKnSvaW03mMPmve
GqvkbN9bdNAd9VlBlYp30rbS0LMFYebC+6N6Wk0kqMWalht+7xUqO5GsucIcTZTr
Ff9ZSc7edwcLjxVmcjMdvUp6t2Jsm7H2FawIySOGYDL9lO/fL5ZTnIfQEwfOc3ma
6M36U1V9NP1M4x8+cxlRdDHhGX/S1y186uU2LD78XQvMlgZVzW9Qt2Rrzkfba9Kv
q+vhQdQF4NukEIXlRwJOZLoa/hEiIKnzzUgaV0fIZqmOLNUg9wCwSZmZxu97QWUe
CtG+Rqa4mjmwYY6z3OzHMRrwv+GweY7EjNOog29K8G8w8B2X29VdgN3zv9dF5vav
RZYXzGujohHZ6YOpKkYb77eJuMxtTlgmyWzofzmUJHpE7qOTlT9YrvtujwKsJOLv
+9/n6TlEQV1AcXORIO6N/egkwseTYKPYKvhjsOPSozqIn8PAiFWUhMpUiCLZSkCL
jTiu7F9S4LA3xXuPBBON7BiSWqiqVaVpwWvwSqrRH054WF++d1k0963t8FJktdhy
N7UTGBwGPImoaTNUdy5s43UuDSe4bU8dUOu4vfvJsHpnNGZYBrVh7doQlPRWkkRr
4+6IJzzuUJcORymHM7MQdmCLKfoGJxCFkZ9qA761mhM0H8ZARJ2N4lPo9fU5JxCv
xwFrXuxlbkj4RHYjMe07NpmKpDzCPKhKt6/Sx/KyidvLc2jZM+mqE7R8Kv15a3kY
InUkwMN3M67DBzd9LK8KpcRN681+L5wAIbr9/hC0HY7gRdcJ14Ss4GBwEtFtYXRi
eodIz9NpR4oueck7DcNx1dh8WZ+auDz8c18b/WDhGYy/zFNDBDDKcl7BanWSuRbK
4Gmi42Ib9oPVxoEF7ZS8UJiV+pBlFx45NIBvzxOYLaHgc4ND+r97HozMCE9xnvwT
haQ2EcrxH9HSMJPDcmC8WOX7BuDKI0GSjzPmDd/gwi37B1jUfauXcdyxEQpb7tuj
znG3EpJbh17l6lmo9yoAFJHN9J0iiUE00BdcXNhyxn5E2acgSZ9FqzahoBHH1rmO
B19d2TrDpm5VopBx/twr6Zv6u+dyrLDTO4RumJdFDH043l5AIPgsM6oNcQojXsHb
Kg67it7aQyBJSCUkcrcQwYWaKxEGwMcAFnf1pV1+BSjdQMAS87HBLI7Hm6hFgXJk
9L7O1wZwJ/Qj2a9Xva7TarkTU80hKkuuydPxUKXXCWPkwlY+cGTEghNS0WfT5ZkV
P2A2Sgg4vLnDNNLLzMeB0M2GRfXtn2iwEQri660IYBxYE36Jf9ymsTvng4+KsJPX
V5DLBk5g3dvwl+1YRTXpnc12L3pN3mMCMbUIRKGSAiZ6SCbIk2eShkHSz3Yc/E2l
3Jfb0MmgGFxPnPR6wTDiWUCpx7a3WPGRo0x6UZRKKl/YlYv+iXNCExbYwR5JMMUd
2rFdYFjvDpGCyGYmdOTpNEmrHfDG5yP+EJWW08rCZfNUwbt7h7PwRjsOr6PfsV0i
WU7+yjSNT3IHDn5Z6wEFa7Zar3QkTsRwrojohxWYeZHZU2Ise+rxYTSBFyuUQDTN
CTYKhKRYZ/cPxRZBXFlNdrdsl4fkzdao5I09Vqr+CGTMK0EbyAIyYgnb7wiaLwok
EGqVLR4nVVrJiFzqrmbbNrE3HzJT3Xhuha+xqQmcCcLdbHu7NusX9nLtxuSYX1W9
Z9OuN3rEO4SbG3lfcqJp66q9il9Ea2xN417pB9P8rW4t7hSgkcwP2cLHYYM75iwd
9wq4xNSpWVsam6Fmht+obzXoEGKPg6TeH/OGUpHg03oBq0tlKkANXNhqBezZTg3m
hWEnZtt65IHpDY6W5vSD82w1FbrM8PT7qZQbNUFDAlllaLn87f+1yZOlx+MoIfBq
DUWoDdciL4DF9EUzkdc/cA2QtoyYNTW9IdbsExltKJTEjOXxI5Q8f09chTprbuxX
gGwDF1cNecereBA0DZJvaAldbqsYjBwiQwk2+cpE4vhLlgS7NYykny0p2fgBe8qr
omr1PPtpxooVrAKazvoIRdP3U/s1r5tqquMRYhE+RwgccbLhc6O1ZvE5vs2oHuX7
qc76/knSdXMKg7RkbJZhMPVWhQGySZ5/vSJzYcSfy/PED4LKeJ7kch5puxOrr1qh
duInlqCH8ccEtc9FvulA9Op4fTbiXsxZdfSnT70lQFGqSMZhrlqFQ1RzXOzLAA8S
Y3/Ux+8XSpRO2CL2j3lgoxzv3J8sLZfm02GTW7lUNNDnVABq6P877stgP69n1C2M
aILoMciUARBRx7z3bX0qiidkvsz2Mv0H9Agifs+W3CAcBdLpxQxJdhhNPLPJLvGs
GsGMwdLWCHeytCmUHO7Fr8nXqmCgSK6kvTaIgX9dr2r964+PadzRZUByXOJmanfG
l+WlfcnYh+GL+tmc+aZTd16nGmoAMVNTRkM2w+aXCdd1k2j8F9VW0Z03/DbDB0a2
VBXqYiZm0UjkayiN6+cwX3x4kDzCdr/Qc6XGvR5xEYb7+N3XzZz19+Q7phUygnpu
depKX5D5kCbAgIdQF6HiH83LEBqKmHDYiyJ2zEozc6AuIaKzjw76iBwzLLl2Zcq2
4haNOaEV0qkazX7OWXZYQUP4FiIawbYX/IXZ8J6lNJReXhSQVZfbX4ApEtdUA3jc
nfNFTUb8rD5XYtgYsR08BAlNrH2DUO0MVfTjflaeEwDHnudgPV+DTr6vlbeMsEt5
MHtJgqJEbdrta36vg5ntcN5Ti+BjW5wh1heXBW4yu95q25dA5GiM+XcQUnt2SNfi
Lf/Ty0zjBZnMBLb6UsyGpQKmX4kzvLvwWKVFPwnLJN0Txn5VRKLzvArBOqhJfIWr
4PwQahikOyA6lqhbDTNgf5AaCFdm71uZd4hl0d3yQSAsXR06upkk1yb7OrlSIwQb
7FLDnfpsH17zDQT0OfZJpmEMuftiLaNbQQoh24ZooVG0Jd+omXounzwt3qVGPrKK
BjmGo6GkcRcXSab31j4GzUbnk8wGG2F87xX1qqop6ooMmvZ+wXzgjW0vt6IFgqJU
FCY1xdL4RuHpvEGBCLLphYw0nDVmajORmv/VDzt9ocWTXz7cYsUlJDe6CcPSWtld
XQqRQvMhpXYE5M5ftehpvLXaOTK0BLUS8Whf1rgNxRdDHnCW9MLUvIDSM8kfDg7D
75wNjKhdvTNleSYDXKDUPjzKvI0nEQbX05zilx+ptwkK/nXaMKY26k23D7q0Vq/D
sq8cZ8ky4UHIJ4ZTrkvfJINFHSaqx+4mnM0/hZY+pa5P9rm+CxVScBitKV5wXR1q
RIJzXyfecXfipyz5NvxPYZiL4pkU/yzc3NOuhcbFdPCOtaEXPy3Ro9mjSYp6JY8+
j3pXw3oyHnm8OX8Mh0X7+i8xUCv1hniB6quQQ4U6N3o+E3cUGhYTKoUAUHMI7y6N
EU0Wj0VZdrGzbwxNu/CZMd3EVA5jW6i/tIXGPBf3YLcSjuqjvOX1yPVB23Ry5cgu
kOqH19+fdVtSCQLOZZGEsmC9a5YkSg0FNA6cn3AkBJsWyzlkvo81LoYksKc3K/ki
xftbtatvgCP0AmK2ub52XaDEaZKV3Y+vxtx3zXWpCYpG6365Gz5rMWxvQ+LVTN9W
lWyXCu8ed9O/H6SiFYzJqmTTGtaXGRWJcl6TBYuV0VH6RY40WJxlEejJDK0YfVnn
VodHhn4sWLxGRn5/CG1UEA/F+xhIefr8xBis0U/J3dTT9uWZAbrLx7b0ixwNF0s9
ZumHPYaCdNhwC10cHXKBBnGZYME4OqgRP+XPLxSA30adYLgPTyFAR5QLQwGvsKP9
obRkGvXWuhJj+3Om4YK+smbsVI5Qj1t4jeUluUBEtY5DDNfE/yn49fen+qMZXC5e
EbmXKL78h1HbaQ0cQuQTiwFi4Xabd5aE5FB6pIiFHydwr2jlFwZRDRLrAW4wBr08
3S0q0kSyJpQWkAIiCC5HkokK6lQO1NcNWgHovYAPqB8YtLkWPsQIVvuCNXK9gflP
2EZfQlG8Pcf3LUNotfzVJsSTxhAtowcDB11KFpHP1PqrODrv4t97OgNcPWOH4+wh
v1xlKWaomRqTAyuKbC1fQDbU7apr202D2ZJifns3V4YJhg1FRLIAuaScOm+lT5/e
dOghqj2ypV4+71Fun9hyDlDaqj5vK6qCwbDqBP2jIfSSaJtYMPAEHw9HiNMubE5U
dmfvnW6Jo0vQpavD/4U2g26f6DUm1bVfRy678C3ioHBXUKTbc7SyiSC2GRZ3f1EQ
d2waGarFwOXzJnNIMqN8blJhT++do44hl6DbmSVetI7vSsZSNuQKGn+cLAXgqQ4e
GicV8hESUcQ3+OWgocZusUJR0kEYgfMdT6Zy15hIICQsGEpDjdrXmLrsvAvpFOwg
h6o8MegJx88ck9MAv/Iwm/ab71wdroCgQ7FjQemqxwh9HH3rXoFTZh+6VL51tCCH
pBv5GvUnBIWDVJSUdttDkV+O18aqfavBKzJf7jkEDbfKMCCpJhHwrX6LeEISvi4x
hB8cV687m8uiad0a4vy516BK4qDF8jSt0C8lA25eTWoY2tXy4XwKrmQGHSqVaEKh
Us8avQdXOxbUa2GvkD/je1Az8y/JXQiGTofgWoaSVrc5laGzgELUNIXpbLWseROi
QJ9o3GOU67T9Oo5yea5NonKXvBtt2Ojjp3h5CJ1+m/zke9fWj7FEENDZyDtvCc3L
mABUTj+hnmOckr8SO3VH6/vf92pg2hhvurwJLGMDCyixQyca8BicKIOT5zPcm1ne
3FVJ4eYxPL5V9fQ1F5nxKY6JAUlAdh54TxPTnRNOvMtKkGPTwU0sYLGFY99FVNqp
OQfKwSyh65UFsgeF2LjNicXM4CXLmRJ5ljrkWnVmJ4u4BxM3MdevRI5wkjCHH6fS
TCtbC86CxrAwAbJcrSHToYAPc4MKCjknkazRI9NYgSvjaD9FtTaI0YCMfQRYwfDD
3qAFH7iEJu9FQaibToVlOMbF0K6GUZ9ojHAnwRKo81DYZYp0mfrtw/EoQd+tNbcm
nx7d3aYwiR35MXIoO3SA9berFHcQ7w4Mq/rvmiX2jWIPQrJCy29jJPkTcp7T2V01
Q10dnX78Maxbvh2eYifPlo5BLMhjVb9u95oYF88PlwuVouyhBbjXpgcLagQTHgGP
GrkNNcAWzle0Yn6WfqY04IAKWaOVey5C3oyQxQrU1ISDCscxiqHKJ6kvO4uTGWT5
zRhqUAyS22pyoP+E+T+htr2E6n5f5XahWzRIKdALA37VoECzXHDqrZZ5loDLJ5Eb
DKEOaRUn417C6S2/qTs8OF/L2WfgbdD6T7NLJhPH+S9ZYgfljHyzBag0psCCjpFd
jxtc6nNh9u6MwKFluePqZqhoL+JvyjIUTgh0Izyx+E7M35YRoPo4k9ISEsVyMvJa
Le0almFpvSrnRKp/+p66WHUgY0Xy38bBPd9jLWMdy94QqLWIoH4Eidn0xW0iwH5i
W0pkXJo4FQvEbsn2BPzRI1k1Cw+uEITB/JkLSlRCVqu2j+RZhCGbdQWDX8sB0WYS
UK1iSL6A00zY6gwcIErJXmx6Lro9EYGmqe174NJAJIxJh+hM2uFWY6/5Vt6pvj26
5FUZnZjdEokbSdK87G0doPRnYRtzMWUmLq2IKWsR4UiVnRm2Aa7KJt2xUAmniKM+
h9fI67GAI+EYpeBGsH5Z8XDiEwlUrafAkQ48zQQaB993eaB1KaRxaziSZVUR39An
i6rKQLQZZDZ/wBfh0LXFFeQddSq5t5HjFKjkZtdh8+LM6nEoWJDCr3eNMFpHoOld
bNjqnZZhwK6tJ0AGwsJv8NZmu+U4LWCIQf/MKHJOo3mTFKvVS0qYPdjxZWJfcZPQ
L4Z/GMc6OSVoAEHXxPQOjhnJqc5ihWRp55biKKBbEUrBCsvQFFnjtvMFYeuRr9U1
RnFYltJBAyoiREsSkciMUkEwA/1l3duEwgeBxcPwuusot6Fw0ir4MFP+03FtrKtf
LGVCwyKh4pKw+1s+OqGweIsuFug7TdvIfsRBtAHqdogpOQR4uOV0977FghCxy/kF
P2k9OsLbu8FzWblz3oJl4iLbw6mHwhz7Y5ftTG/oscdcRwerUnjHGkI47QR9Tj0V
kRzWozeQyYhLhOW0oQWN2klCDTOfjCvML6w6k/s4wGT5v7fS8zBX7BUMRzhu1Cuz
9uAWGdSgJ/DQ/USvk4Q3fjC8pO1pRv0cO7HgDv+E4G5pz0Y+I2dUIDJP06YsW/8f
p91GjAuNJPVNiANdFPlqld4Zn30yXA/anC3Qt8SOHLp48GTR1pt5uIs4rvAexzEd
wnjphH2hjDMlpstXolCtewkfDtKgo2NDKUFjPqjtoETiUycNG5zVoZSzyXNDCLD0
mA25ttTARkUNsJpWzixoAcEU457itARJI+qBXczNmievRb4UY5YHcOZgzzJikOqB
MTVD25hzNkcMH3WeybsbKJnRQst87R90RgaM0DWlyXYSE3A5vz7TCy7nlDpL6ayf
ke2ImljXCPFI9Z/HSHuPh4b8PVAxSvFKiGQGZyLZvG0J8zWh85tW9/pbMXW4WIpr
BMqn3/gbKb8de976N9MJnuDpTo8D5wYGwzp07MMBXYYAnr5x0wwjl4+GwQwuEWtg
ETFSLPvwsSIog+UhJM/tl/5T0r6DY1P0COMlTS0xtMMT3+rbQOonpHRxWuH4C1U2
8Gkz2qoPGbBqyNUJ5r7BHRrtdCZ3RuK9l6875QDAgk1at1TTGtpVE3QozUcPJmpy
PSc9wowrxXsh2sS4Vnho1i9V0QJWgMCriNrTbj/yX673gRtOqKAVWTuWEO2b2oW6
6tHSaq9p50VFLyHvMnWo7US2zMEUtHV3T+4XbAkt7E13aK58IfJSwRXSxiLnYGQj
zASl3tcNEOIksdHGkEfzjYKvMPSRl/yfibXkBRNxjQHqtm3ZuGYN9DY8IXQN6DSm
ykpBe0KsHm8GIsGej2uzu/ItKCkuZTrzsgg0KewsIBVp9HrTS6zw5R/S9/75chJD
eukXQ8xGb7Dy7IY3G/n+vH9+TXbMQzb+UOss5FHCiOU1u4fJuX45lr3YFICuwnMw
rfhN3jijIfTCB29yvY1bRCsTMr0s/tZHxEdIKylP24BR6xQ7WLd896jmyjXruUeW
K2aabykYnmKWxBU2eKQEcRPTUkX+tsvXer9zK7vAmtrxgNMDzVKTkHKG4X2Sb9DR
CSMtkp8TgHnybavQazLYoJnzzhBYmh0ZXxERUVeTnQapi2sYWGnETRWV9D/othC0
nK5jk6KqxHxhY5cul9wWNZF+XWvisRAXfE2BxSCHXxURJTTwjb+Y976Ej7l6j560
hRGafdzjhma/ySZAX8MIP7dV0Idl4ysSAwmxWXyk8ZXgcHeW7Qb1nYNpUBdE/Y+l
2x8bveh6IcIoTWhE6yEwdh3Yy/Y/9YeRxNKgPPEUfm1emQRWNqYWg4eVtGckfWP5
ICh6POT40fn9vfPHy58Ny99tlgstUS+n953ps78eMK1IlspPRrvj6wFhDXUOqzEk
p5TMg388sE0TcPIeonT1Uz4eJMPFxpEl819VZxiJVQ7GHobFaS/RcmtLkrzy2Fvb
avMJLjzZrojs/kAM6ppLxTCMSCjeBQmFuemg3MrQOS108YMOjewxPnXtPW9GB+h2
3p6r69dAVb4krLVBGsEEgSHWouleoTWOG4xIcBO0uVTYj++vL7Xbzof81znehqGn
fgWKBHeK+3OfBhqktyBgoZcw8pgV99EimLLk/06vc1yD0fAwJrJi1o5sIp2PMEWi
XRjkkllfC5mTUlQXGh7yQZC5UEtaIXsHW3dAyftWdvf9Uj55MOfzIeLlKLwAlrwP
ydu6d0Aav0W8r/fZyzgbo/AzZi9fw1d8y2uJ0rOHU2UIewgqeirfNybMBguPgiMG
7v6UNnDhwtJbh12WNbc2Y/PmjaT3cs7X+CFb0R9a2Y7fiUY6WkZopIr4NqS1L4B7
nmGbTyVT8jRi8FbQaCozytnjYRtGKrqfFjgGn7SYX/WmuLybl3DF5PHUv6IYu5O0
GYbCqepu22EOb1Id/4wliY367eXIuOQdzyViThWXgnbFW61n+IY/+FAvlX+1MRaG
QSngYBXECDCKxALvW7IaMFFFwg3SGxorbx6fziqUNGWEo6GVJVJiI5S5OXk8LQQN
YYnZjraBYIeGa8j8bcfufBM/ItChMfKcZYjy5kf/wktHkqY19yOV2ZAigANl7yoS
wOrr+bNgwpEI5DYDXcOrPbRk3tZWHdk1/Hk29teoqp0lrt+eLc1WS93h+GxTSBrz
4tSp6ozigexY2hKmTZ6lhveWGWfSxtJI01gD9lHLxUbcJaUPpCOf87A8hgOa7/XG
IwPjLAOVjC0+RjzF9v57WdvPU6ij4+ogw2/m8Oo35qLuy68FjgFjYs1RFIRisF4T
CnW0koc8srCeQe+7b8ArcdgHCu5L/nh4J9V0mChNrELADWt4N0ge5Z0ACO30PwZN
fVmHOvvRdfLsK8KLcpJRB52zirxcz1VXWxQd68lFkVLWjybWqJz8AG3Z27gh0ZZp
qkwsL6nkYGjzigX2sXIEtSMpn4Gcv9nrzBlgZmpxGMCHdsVJzQNY7uKtA2/14wC2
AuV3E+ywJYjti7MQsAOSXMkREGIaYnSlizK98WcgXlW/tHDuhx5nkrUslco2F5B1
TBKls//2UXcig7JxbTZUNQFUFnM61vXsmPh9tNiSqxEyO33yNCgou6BuoAhk3DYc
xhpJttoozc8vJH/CuEg24sk9rxRzD2ZJUn0KLg9rFzRTUtXz6Lql0+GHJ7T1UwQQ
DHsNqxzjw90ALayFGvncxrXsTUrWpwW7EHVyVUCM/UmmEbKLMz0LXXC3tsnE2rJW
g9jjN/5d9EySMHXdCNYB1iwZu3hSH50ij33/FJJ8NIFk5q0jzPWbyncqVL6xVaDQ
jZE/yViCut6IzSpkKcIzYL5DtFcKmTc89ASlRyOeqxhnX/pTGlGAugPhXSUhh3Hi
GNi3maXutsa83NejVaE6UeSv/KtHM/HROATCv0hpUiLXotSDCgOSe83vL6UuZjFQ
zG7i1U0Iqw63ZgFprzanj0KU+H1kD10Mj5kn1sSuHOqUy9OqiP+dGwESsxNvU5Fv
2zCxVOgUiFOLRmkgcgb0x/fK+CD8M0fpdfIjNu9RuAciLf9hF1MCU8nUE2D+NMOe
k2hzKOdgtQMWEe3NLkMAmOHOc3cLcc6CJ94O0s9pgRDDtEgrgWvTCw74gkTse5/k
QN7YYVNEVt2/FckYBaDZE9T2fBgrW7HTM2ZzrjpRum3/mtxxBdPV9qXy7ytDeYK7
iiYmpEDbTDyOV34XBVlcTzg9fzQZOh7v9QJr7/4p8Cdkm5xu/k2nLKmR7IADSsDz
PhA2BUhamjKdd4L5B7KPn5BfQODHLMe8aQ5pHS664BzVYSMazCaDhHhS1aUbeuo0
MokTgd3Sn1LkY7L8898B/DMx1KsOCPHR1JFbcAMcaqixb0K4DBtsGgzPpQKmuFGs
apn7SH2UztQ1x/tecN8+gPBRNtd2qvmFsc/LMc3L4ozaZTpvZH8eQQKqgDIrWCP/
425I+NelczVP12wXmNOQwzAj4Vw/ZsTamNl8hX2izvh+QXKGsPnrzxWcwlKZgc/1
mQ2LJVb569mxCVCQkGKvJG4YoH2FZ2QogPiIiFJba5i/goj7/0ocbhYFwd2TQJ39
Y7Zvuxq5vYl9Pl5lIegchZl49C7L2Tj1WDXigGMGsirfUrfcxUvs9A/M9sSS7A6I
XuH+3zlWOY80P9klohr3ikpmj+NLghlVNFtwhRpo2/HiqhSolwJ5tNmq/QIDFqIi
RSz5c1qyXXfQFkdc9jh3gfA3cBbPFDWfF8ZO8axOSr59dLSCMRDJebFl0j4Q4evJ
L4Eh4PL9NwnK5WBHxQnw02PlB8iv+pD483+XpKKCFmpvfKcCSWNBpR2+jPDGIVU0
28Hsk1icq1x1ugGlIdFJIE7jlLPraJSWNOirEeaTi105DmfhuWY44YySdWCsmiKj
+ISv0yS/bvcjqAVQ9LKgjFOeYmIEUKbd6U/rWn9eLYU/J0bwgd/4hD8TNuruFRNG
ooeKywkHc6p07tMpBFVkcCUm2aHfFgoFHzUhCTrZGv0I91+Vr7rvvqcZjSinE3/F
jTFwiB+ETEn67btNIzzo4W1d7ChF9gOjpyMkBqO8JheWzRxL6ELTigYHbpty8KVL
oZUgLhh7fxAuX1kCAfp41XbqJFqgDCNOLf0q6Hs5fwnTwi2y5/8WzAmGpAWLLElC
Z+95gjwpXPYq5EAWW8HQTsKsashzDj2se1UYBaAyi4I6Hxs7fdRrrHjAo/Ep+N5h
88UoeJ1xGbq6u26/AfaZHjRRNBRFFYPJbW3/qmUOietIZGF3uPB7if3ZWh/yT8W8
FBbsfzmRCn40uNyS6PcHcMAF3aIoW2ggHwRiuFT5XPSNdIyvSc74tI+MDZy9GkTo
omXwOwasOvIJYCJOrcLNoLzf7bEpJTTXctD5ysMUZVvpgEBrO8eOphQwDgaJePZP
R3r/bipjuHUrQVk2qwN7PEGgSED+vuuqLn8Vw0iNsDGcK4fLSuZkXrQv0JABSYSd
GOo6A7UWUrAX99uKYSPcZXvgcq7wYFNBJsdPoAlJWsCFZOCIW0u6hPrMUi7srHS+
QLpXD6WGvjFc6RGa+qrX3LUt+urQE+B4mJLtJKx4hebp9VwzmcUU9GXvmOBDrM9d
WgLbvyrUIUpfLBqvuDXbIhmw+I5TWjurC/NNHfiga00F8jn+ZHP7aHtpvkVqOdtX
S/0KV19AbqA3pmyn1W+3t7FXSV6vKtZldvOWlMXwcv/BWuzJkWvhrpRvTqwm2n53
aya8KWiDpSJyFILR8v9qaX13NzxFgVXg+UIHHq0QIq0850Fhnfq+De3SMbMpew3r
200iqcSYV0CJOshvCU8RUHxPS0+pbInGYct/7PZ86X6PjecneDFTUS0cSZt6LMBW
9PUa85DhOZy5dsq2qh/qqz0hi53PRw0XliHyF+ZAeuIEEEQl+QkcPs0k4jwtvpSZ
YxS17fNVpq6fKpFqPmKearPD6+AjBatUApPe0cPCWZ62lkVZ3tQqT6EeYmKoX/qa
mAzSoJlE+V3q8iFjUC6+7ICFn3aMEbotjRVmtFF8xpzaYQqLJfjRv6H0/6IHVLJT
PyI1B9WM81M6fepAkRwemFE+Bt0vfUFVCnsxIKtAeWnFAzFR47DDPPgSEG0GCtQJ
sHxSY+Btuww2oJ+2rr0CQslRMosSzQB5njrUbnkFbyh6iQI8Y5k7peA5PwD/p3EI
nJOQ8qf1J6veTzwZeEtVtGIJc1iAGbEJZ8LOoJ75nesoHdRl9zBoHoJkNjcXBCgY
2ME08YP99+mC3WIwQ1jde38tKdRKe4tM+6SaM3LbjC8Y6j7WE/rcO7Uw/RM3UlfA
kVrv+OE8yLz9H7k7FZy0Ly0ixb3iS93/53Ag0cKuOF6GpWemjKlsi7SsOWDGJw7w
0pJiNiQv+RHJ2JOUTkBWpjqJnUS6YESOJxgqqLQnhnbBeJh9AR+EFMkgZREKqWXq
ofat2yffIK1TTqfFftEhPgQKNWlIsgCA6n3glz+fDT4Wvly9cd7GkKrE8O3tlIJ5
l8hJjXHya3mNcIr18WK0D+1tXvH/Txb3UuRKCBWS5f2E7z5upbnnwyM/TcYIS527
8GJQRD1YyHhF1mdUbYa+OjT3eL/RzDh6VZql2tIMb/QV6o64ieOC6OVn7ZEi94UN
9AUZnBnWiX6k844PvnyF/ph9wO2eU3UI6hqv72IY/KQPen2cEMLOVMrZBZEu2wxa
TsDXfnaF1R2oP2OqjnoyOGkEI/Hbtymc9UE3fh2g2bpoHjOH8L1weHy8Y4m3TP9s
q8MEi70+ETfyqy1U3wvrMwAcXbyP/Or32n1L6XxFGhIWVq3u9bueLGSLPpNwR6uy
xio+vQWfQ0uTYSZSB0H9fRAzkeiQIHj0W9pnBrGVUHD3G156D3VbXRaIYVE0Rzij
NpSXVbkmGY5SuBrQyZ1D1nFnLIqbFkCKBWSmo5PscFu1mHwrh9zPJuNCk7g9+Ucz
iAYFjng9otko1G8Y5BIYRTHHK3niSuHulc1D1JAEVwKPniTwx1zI1nrONHQbKqGB
ntEkyCjzcj68sOoztw/Ca4VZxOLjh5jffMAv1ETk3CfkS3hiBsZkeQkdQuiWwRZI
RUhlUxo58PN1QNS2CbfxsHHgQ/PqhEy6GjfZtwUtXErXw6+0lOLf1D4pZ+dLw0Ki
xJKtkLaRVMslujR1x9TQ9xGmXvnnDNFui5rnl7Ee7ztlZqL8A8Emtyaql5XBw2V9
esMOcwIO4PdUzalIcm/BxdsHzN0XoTQhgoNlgj/RdZ2DJGubanKrzBmny0s2E+bg
vxSvrIteYQ7fiOOZ0gRuUT3m3abkpuPsiMmXTo0ucyz5gzwbAsrygtt9epA5HcpD
8HBvJhj22ZQHop+pAVKb+FWiAc/LvKuyAuqklWho3w0rNBWJ1LLIXxIlmooXc4mD
j5citu0zHEU5g00kkLWs6b61zcTX4kbhp1FbkXYPSnfYb7OCc9gjWMaWdVGT9RNX
LlOxVvqwE1TLpe332j36DUyJOvgUt9lJjOGqMHlIt7IeJ/hPXOyVc+zRU2Vzxmgb
0l9q4Vp5RadEaJCvZOlAWja+Gbw6dRzYpqWndhsGEChv0PLBcQMGl4vMPDueOWDI
YhUEcxIgMP2IHb1StMvb3zCwvbND0T83vSO2gx1Lx/T1wK2GHcKxudqn6zVkjVU1
qtaGq2AANJ4koimXNGzwcqh/2+eGj79dtmgKigKu7zUd9jesh8BaE/4hQ0BAxzAN
LYydohGv0dbzZ+50Kx2/9hDImGemi55CCjgVcI/mrAxmHtyLt55rnTiqiwjPmh1Z
sqF/rPFZz2qrCq148QdV9xpX/9L3SQgr8bbzzjoStpIB+Y57RvefHOeI6FY9Bvi0
vPtZlqRThQQbrcPb5mTuczJ0naXapUcrMmqsuTGK+wiqChBxGZ6kdhixAwgVH4Q9
GegIQbpMoM0kcNgYFj6v8TtEkcKnmAPYlu1CflIgWqzZVCgzf3R5/6dgGL6jb2SX
YUraPKGt44BpMLUCmWwudqOQJVl5WIbRSXXAZ3T/9vgvWRe49UDbAXd/c+nK9u9J
B9aG06yM+KqPoBkWHFZ9+0Q9vmWOf8BAt1aqwvxTOBtA7oZlYlAfZboiELY+ps4k
kOsDKdnwXyxz3pdXFCwBhz3wBnxdJ0GI4FIR/mLMSZs3hu7YsnQvekVcVvi9E7ct
aMSeTkQlM7oNbXc6HYG1qNilL+bA/DhZtRolYnggEmSftJuMeYWnQue12UmuM2xX
16nM61gaA2Qz6iLGej7ZkgS71J8sqOPgL7dK5KdWO+cyHG0lhxTe1QOpjLvKvG9X
DUUC9gnZjrJ8HCzG/In1VPohMKhShbIMTQiW9RDQbC5BBDT7m9rz546tm+brX0gs
6QztVs1vGvjD0+i72HX0X3km4b3QbR/26Fwo4PSXdK4dZOzIPxvenmGH14TXkISt
C2xK0hlOkByQb5N5q4MWgPbGfAEVc46KBfLn1+NRDRpJ4Jbgli4CEGV2a16bJIUT
bHiyL5pVk0WjB2rZ9HvpCcU+GAGmJiHotVwMh8WL0GYM0jg/60JMTbr6t9Fh/4Vd
TxzO+6VSYNNPWmglOWyG5+SiUS+pmcGUqZ27PQ94RYjkBLjktV/oKPY5x5n3u1c9
wfwCZqDFHjZ4SVNxaEiomE9XL9SVwgNRuU71qhVm2Z/qx7t9ahY5R6Gg0x4ARTW8
ObuPuW/4Fdu1z7DbZ1XJrAuLT2nrK50Or1MNvSw66KEAu6ZuGjRoH6MHmt+yBZUX
tknQK6/Qh8z/9Uk0apIqG0lWeGDrKQEXVyY9ejFM1NlwDJc/+y4L0TAGEGfUtN5l
F04+uhzNlAhqEYW1dUSiJrPk2W0O/OFkcfRXxXd8HKSsk41lPPWfm4IQg9XXyFOR
0TPZYX5MKcxdYAVvXjxIP8yLBhGgEN3w/sKa++06Ncv5Gyy9qB2nEEn4nKefpHf8
zlQECfou9AKq22ePoiDANTjcZuBwA+TxFREv+GT+ijYnKeR4a93uFFFE+2GBocY+
ekSAaEXAv2Qhz19aphoNDQYGGoUHIbTAoK+gqqpKGFyW/pXQk5v54jWjR48j+358
16izs4k+tLky7TzjEYuF4qXAfiRBOITuqaeW27w3rl8RhVdbpAXRjTNTBI0hQcue
zGfqB0XFebARhsY4OP+1/7lEKEbBL+hHSEtzsWF+IBFwdmWMXH1H48P7WK+DD2nL
/hEI6R59ROipqGMtkACOBVguq+yt41rDwO14skFUepWrxSscfgCfc2c4HOshZYUl
Rw/4uCm9QTdIPwXWkCGpsPG9ovPzsXjamI1BtRpgWo+7xyx0L8oL/QJw9tgRaRbu
cXa22cHz+RjmNW8PC4gG1cQEW7PawMAIeer3Rx7DaUQBjH5N2WKYdPHDzY2xBkgq
VGaOzH9wpdkaDNMU1sYvPSSLXcxkkGLUVSNCZsUPJIgDB41tpnVoEuxrIpi8ZtRS
LZSgOpqpc49qF8EP18B9YMBp6HGui8Wtfzl920citj3pNyytsvvFimzxpENjJk+H
EGbTj0yzQYBdGwFMVny94VTT/ccbjYSLRsCN4fnZyGJ915TyIAUYHcDVUfS5iOGi
ikjGjxEzENcthW/ieemONjmz6MisYAjzU77GwgiJY+JJbiG/7OGqbkLMY09mlKff
XXvEx3fa7X4xW8xBpr63YXEvofPGpEp/46s9YqJIac8V17leA6b4jPDZsAo3nmEw
+qXshLkWl16fWys9jdPYgNlAlf36+FUy6PFJtRgqPKeJi+6A4Sl/7Ndb3vZaiGSy
Fd+wj4jpqeBJjMBs4+9AVQe6ssCDpTg4Xo+NpH3CxI8zoQmXE5JgxhcyYYBWWo0M
W8OyUaRPZqZgD0UrAVUs2/7aqhHHuiepXYBqX7tCFzMO6EAdaik/GHTibNT290NT
1edi7hE9pwSMfsl6IgRjwU+IU/9qetByu3TxzuOhmJVcQavdKTEECXpeXxcqULqp
VoE04PPFnIv6HoR/ZMa4khQOWQHqxEDqd4dt1AgCW5OUoAKHvUC0PV55qDT7USU6
41BASbBkNuOtqIx0o5hpqw76yA9n3tpa5LhBsJBx+rGk2xRnYfWXQDgOiFu2EiOd
gqmee2JDdhKS9aOS+JdmaKjRpG4Vk34WjT3Gaon9RHVPvMSxMzxEAd2r+w68a6dW
vFkLfaKCVCdcinek0H2YY1PYgP1ruSoXpFuCetL4ZnI7xf5QYb8uNdyGFhIJv4F7
gMzo/9ArU7b0NeDxEFUr5PjC+7yzm1mi+pKvnPti16vHhrbzOF/o+7tZEa7q/c4w
KrU3FlQiYuWrFO997FUoRKDbdyGRNX4ca5b0uYAO/UH4/er8nQgUEgOx5wgLnEgp
Q9XylkywtBX59S/We6jdaOeHeV5V9+Cj8fjmWcHgE+AUDVK2ZkBLFuMnHv3bP209
mlu5CKh7Mum7I9LV/A/UHTj6QiCzq/zD+z9vvKCySi9mHuhXntXyCywMADuTVfe7
Ic13XqhTkF/i9GxmXk3qHVkyg1eGfbjUt+5t+EWE1voMEdwZtHG4smP+8/1gyZ8g
40n1PGjl4J8J1MVeh+5TgJT6SwN8Kb4KCFYI3tDn27ylfFFz/QdyzzfYU93VO1nI
Iw6txag3D1DVkJXbWkF3tjMzixwaahrB5Csbl78E+YpGaJSt/gGglUyfMa1+gtYp
sOUJ9A0frQFbkrpxAzBLjZ5Gn2E0srGqXyHwY2EBwlNNvFEL9LQyt/xpp07snHbd
lKd7cqPPQp84AyNQP87B6oJyVa6qnq5kn4QpKuI3bf6zmKm5VgsKezcJdYTX25Xh
h3BH64ZE7F9OPqVy7hwuRZuV3kdfZOy1/Bt2ftbM+SfFrIDD2ZOHdHnS4azJEGmO
6+M7sOVDqPEUrq5W1wekId2S4v/hYuVPSd/kcD6CppHdo8bcEwa2rTbRBULqs+Ai
OBd07b0cqt9o5qYXJmx+bMeA/W0eIrsrQ8yT7jE7Kj3PIS/h0rD6OE2hZ1X5be5b
b6aJm8Vzu2wnBU6Tm3dNFcY3xdmi09Y25AuGCZYeOI/NTmLGQ6XBzfWsaI4W2pb2
UblCoB1M5xcQQjBhwI3+uaDeRjoG/ynes9vXDFBv4qL88HDhgEb+C472KObk4cW7
YhLdBCdBXLQw2VVVsIGGzCYBTd/T0ocL/keDb7AP8DUMLSYzrBoa8Q+mH3wlD/ia
559La59qDkmPEnUPpq0TmRVSYIlkLoH8W/CMfN7bX+huwuq0VsEZ8DPMo8ffac9c
eQWpbsHoJwthkYKHIAbrzeurEMxuz4FMYArnsm+sIHV9VnKuueuuL1rNFtwz5q5H
s5iVb/Um2DvUUWczqxiPXswSCa5B9+QUuRUR25bWlqY4+PIpnNkCMmJUrfrZuj++
DpzpJCI5HRvx9wY4WmdedMyAb9eAKFB/bDshaDhDJjM182RKKyMiBPKyaqpAUE+a
SEMiTI3maOr6PTWxnwS8tnDxz7pjR9hhJ2IU4U/fN7ZV2Ov6q4kHH4vNymjRBxRu
trFY5FpkWuNy+ds7S2CC5wAFN+7LT2E/08oYRkPjdEbcKp7cYvcKky/DCwrwlkps
hAdu5eMnTwwW6ZMZxcwFF5WaCi7PIln/ewKRHwBTo1ERuWjbmkt2cq7uaRYUnI8W
mZL3S0dedz95hjklIOQBz+3OVENzVXBVE0cfKomoUfih97HP7e9MPASULUt/zqOz
3X0cExKDYXZz5o9bw5/R16M7YtcYmEVuvIQfgVN+cFwDfRyNr7cwa8bAnuPfX/iV
GA33o0wqkN0o1qV72MMLLMp/tgw5qqTt027Xev7ga5vxLuTP7CvWbWnG2GmAHCph
MKqqs8qFqKsNqipVZ0ZuoDpR5HoxuZpRYqVn0T8+CAQ+6dfX8GYpkR9k41bjRDag
t+3IN55cTYNoCPxPKqlI7J+snxpFoIkpV47CFIxmYV2XizCSML5W/VBRQb7gscjN
CNGWetq6sOWUNVPR7rN90crN/7aM3kp0MsCrItNW6XckoSyPmPano6oBdGudmi4Q
J3zY11H+E0oL4hVHR8HQk4dUN6+xmZpqFJMB6UrUpGRKBePoib90xD/aIjGF4uUE
BuUtDWg+kQDmHuJbSxtTrcOMvAc7b9AFougH/9AOD8/ETs9UMdUzZwJd54TQNGzR
a2FY9AXURevoc52haE/30Wvh9gjXsDDOCV2tPlBtyMC5xe26v0s4X3q9zRejxc+T
UgshhgVMu8Y2Td1bTaF2IiYD4otk0eOLVb0IGfsDlfTGBasI9GCUFOPF7KKmMXrx
zXAs7WWYYDjIQj3LsL4DBScdmWmxsMKGT6qMoG6cNBVz1rAjdQJ6AjayncmxY1NR
QYZoyJeoHU82/ZT1bSn+l5HRExdskELKLI8vQoFZ1SkPqxbCMjOf7BLw6MIO4iUB
VXtEjR1jN1YEspUeOEkxsksnFAtIFeVF/XEaDriZg4CbOIlf7JjhJL4B90qBuYq1
YdC4l/DzOczHSsbW3yfg30RrsxEyCFS45s6vkic0hHni7nKKuar/1KcJzunrWU3X
2ffZCNvu5Yr6bWlyl68BX4n7SfgCtbdw3fXR2gdIode19ckVX335tsaYO8VJr5NE
NH/UUC5+CyeFjDtF0MRB985n+cP7H5u7YNXeSjzKNae1DpLFoSw6U9R5Q52NzZE2
4hsqGcQbAGlWd0d9ZElsvU94EAmxdY1MCYouCUHWvpljt7lccTOxDMZqOh5K1yha
CQIjhyPkpYLvdcBD9dojY4PAvISmfAVDU5uxm80aB3Ke7GFRvLEt/29BY33oztXz
eKkxQigJ9Pt9aF40lZFWTY+m3ShCFzRHnAglGZHPlv1ZeDG1IjnxWZotnK5/qbRc
xr0o21i+Yls19SAjZDrtMtVkEYgomIYffOioEVwajZSZfBLKs7mRX2d67zI64wrT
VBhyfHAHMTHmfdraqUHf6SdxPCJtBiE3wtPOCuPfRFcbWD3sF4VNFI9uR4m2mDT+
TxX7uxKoLmKV5XLuow3dddWzhtrI01o3VfnQf1t7pjAh8P7qlq64eSVVqdc6Te7q
UUveyzXiXnahyuwISBamifdTmkS4dNkHBGzfP7uBCWA8dzFaA75wzRWAYQk/CqfJ
kRmFdj2BcsY3On52ncqyTzmCthdRbsSIWFcCt/9EpeKoD10Q/pPL1Ef+HH/wX0eO
N+XWywAQeu8Fea+dcZk45U55NsBgeOVGiqwZ0N7ceocSTbYbleL08OjDZrpL3Gb0
rVHc+xEP3ACapUU7rlSjC6v8CuQqk6n7erFJ34oJoWmBnXbmzjvQgiKCXx/t5TWh
ZYYqXgfmYY2B0l4/etuiy4E3QFT7DzS8Jj62qTcc7oWkeKksFygGnWyEK1Is8dN/
AlipZ8cg4dY+1ImMEDMWocaAjKLKMKyjxIWdWieY9QyK5MSrtkLqsmIqdEj+dQ0L
cGXBk5X4+e7QCBkSf0+/NF7d4Wzk4rWU1/GM8pgG0/sZgQ1fOi6WR//KnB061+vm
+BEwYlh6tFeAfAyX3UO0U3k0BFtDB7j4LqIe4YpkazPQhIoEjxakjSk/d0fYt63T
S6YmCwIaE1D5oM0X0mHer8EGa1f3vdmMPjQDVARxM+4JsDvL0q5iEKFcdjy0MNLC
QcyI4XXsBmVN7RoeXga/348WjB0h+hgkggS3iBe1bMW5i/ZVPw9GNoUTWms7JFal
ESW/OAe48NMy4t4O7HxlFuT6FsDWmPDGKinQkKZhqJME83Hb3bdsvn6cmJgGvTG9
80OG7F01neM3XhQmRpr0Y8FTMzH5dl2RazHNG5PI9dp4yVbCysgYAUbWKCFxAgBK
iingP0p4DI2GQCFhvXaulvWxxtCg4CXtVOmUZcsa8TyMI8RNGPuIxD01X5xDO+QQ
EnIkep/W3B5dbTJruuIgberU+rY1c0EWvJwWxFsDt0kKHY7tlCANAJ0jazCUmk8f
a5mKv9c93Q9TY6nmFI4UMe//e4pUzlFB9aGhbe1Ts4VG2F/ERM7Xvp0kQRHx067j
QbTfJg7gCDHOHtQKZfvwJUb/Ukfqs/eOaQaebS1GGDR4WqLz8nBFMfqygHterUcO
O7AHmSuvHsMdh3tR+Tm+hyyznqsCEafiY89fGc1KewypO48DX4PwlxXep4vJOuwi
hcsGIFrioqi+hQcEzzlSQAOhWezcE6DmX9JSo6Q8C9AKCA9Pb8tyHgUvT23bHW4n
CqQWWfmUkZw+c7vNmjqbZQajrcEqYHOR7U6Vc2zHlPqLIzaa864nrTDOJvR4OiIq
bu2vgoUb8gOHTmw3OcG6us01/Xx5oR8cawYaXUhUg+Rf01lYtumurzSutx8VH0l3
Y1QKrdlgj2hIJb4lQQZKChtCLalc6ppTIdR/GVOQNuE0lehE4Gp58Yr6RgDBL48V
4DXaTqshpwyBWi80A13V7EFHbLUHhoGxORBW16d92+DC4rOsMGM/TKd+b1Vkfg7+
g3CqG513smTch3QrtWWxvA5OgE9oVUV1/JK6gciqNg+ISfJ3TTsxqVD22lnmNLWi
afGeYpsDTbb3UXZgqxfS5diPj4r0iaHUSKKoerQQciTMGCJ2Gvfmm+mc6v25HI+C
PQykC6zsUu+u4Iy/Wj4lxjZdf3vhJcbgn3V9sIiqJJG9T5bXpCZhlmXDgqxcURxI
PZrrsHCJoLeY3cttUfuzC6G5kHgJQB0S1X5vluL8CyTyXRfFQ684T75uON9yojIl
cdESxdj62I08r+A2M4jUOZkNgjW87dSFQF76pr/gR7roruXOd3EK3uuyz4WUHUfC
IA3IhNc6W1bmPM12bw8lAcfas7iXEPwIQHCLh8LGdc9xlyOYEvyhoid6No+bE9Tt
3gqTxNTs1lwPHfYRBfs2wql0D1ZXT1yll0siMeetILGnYvglyjwkywozCiTnljLK
Eybl/X7TUkySDnttJKL8QQwHA1KVfAtF+iA6YfkBXo8p52kElrbYYEJ+BR1as0b/
7JFyFG03y5nvYsrMUDxG2AF6/GUmdyJ9RLz0FJ6qENn2I8gaj00HeabT85kNB4Db
zt1dVGIQO/JjPDGJb2EPC09y0DoAqWhBQ5trb17lAD/p8C70mcvJr08I8uCYPJiT
33jicj2URm/G8/iZ5WI8gDNx9tPaGdfgccqA85Ejz2xA/+htuvReXLsKCGcMIn7J
lLuRpYxlxpqlrjoI2+i8YdPLwWfz+3+y7shK4oTR8XvZ3SYWzM4y/kLCRRpSvJGd
fi3hMP4UWVcCCz7HZOqvr38CKUybzvl4iCs1zPxALd1sgpHmQJI1F369MUxT7wQs
59oWEbjCKZnrgTMdiamsmY7yJUbMj5v3vIltrwvbcCRmXlSq6+OLCLFGY/Amkw+O
ObsLdc2LZ2/wc5FuZrQVbKKJ16fI+ywFGKnI3NKaHShvjj8h8r6gDfCQM9GNiMlS
oggOE3zq8/1JfZdnEWbOOMXcCBbdGpTu+K7cGAtNWffEz0iNYFeo2FylzvMIVZ6w
/LTmsaIfcMba4qN7cWlPKEwg2qhmXkVzJMwQvyW6NWuzE2cnvQbAlPokDKBQKuR6
dLTXbETVUAFwfI8sUzN3T7AdObkqtYNZiiIIyrCNmy5WIKz4vhJOTi+OSjzgUzPD
t0Rd3GjSOVvinQDvQ1F5MALvVDSuwJKx1gYQiE7N6H06H+pe05JPuToEZITdyPBF
+2f7gS4jeylc18O53Bcw4QYyrjd5NaconjaDNDgiff0DWNTp+nFBFwWS7tQC718y
pwmBOl3agw3OZMzxulmH2ytMiYJHmLLN0izTH4+JfuVSd9GrDRGgZedfg3Rxfenb
Y+8aF8Eeqqn0wrNLrqScm7ExER6O5arutsbjsQl213AcekXhHZXvm4PTEki1pPX0
qLfiD0RM2BUstRojXbc/kLva0I2SwiVjf3s6gU3uTIE0C26DQji/5RVJt3xaMLAc
Je3t0u6G0fAcaE99W1polLFjwZEdU2dsKMG/o8k/VzDI7btSO+4ihZqy59TxSx4C
nGJzOE5Z2dySPiBhjxH2kkyysSFgA1zGd1+7jOUsn96ciJ263y8A3/4ztwu+Q3OL
mGGWExQthvWxTAJODUH/opdhWiHBmIi3yiVEwa8H1dtTGZOKYszitE3ig9cs8+b/
fQXZiKsugBTwCvBwQRguQfNBG3shDFxEdmickClDozNrcqjBv9h8w/oyhDBkBliQ
8mnTSWRb20p2QB/AeX3Tnn5FNZPp7xBv3FwwXp5Sf29FljHhvUD/ri68JVZ4dioy
y/GctbKhKaCczpSdgDZ9/NPTlwNcYtRtdEa36CqXdZrDsXBJuDbRYJdS6gtLK/aR
qvRNQU7d4kn1zKJ7i+yiBpia0j4iT29MHg0Gao2VVbUHM2Vf/K54yPKpB00tuIGf
6d28X5Y8w8Blb4AqXDfrIlSgCYQRWQ30mv1mSpVryCGCP+VzRBeWXpTpY0Dwrdxx
BgwKHJUzu1X+AOn73vpH96TxzXI4MAQtx0HQxOFtU+su0H9ZZEGRZV7WDPzR5Qos
h/yWjaqrcoOxO9UNNAvcuoNLopzykpjsYz7op0IDpCHsSKbABeMnUmBDap2oQz6L
FAAxUwm8P9huVqAXVu3w4hgASmVL2v4sZrgvZKfkbArrBKIAlFkdwY+mOJqLC9jo
tmwxhzZdSqudlsE8/YEZNCmhUVrcfkhDK69QZFxkz/GRS1F2vKQAfGzlU3IY6m0T
WedD87V3zHpGaEw7UzUmZaZEElYvHLEfpb/B02qv6VCRtzDmoIfetfn+w//Lm1Xq
/eb+YGtJqsJZm9YhPJId2GiaUEqHArKGP2IuTmlfnnMkLE/qFa2HrOKuTbE/JoZO
4LQJew79IRzLFw1iSRzD0qsobKTY0wYGLmz7Tt0Yr7xt1ROHSpt5CwZSmCQnQaT9
KN+CzP/Wzd54YB8PgzHg3+LSbQaRaCzJPh1+kg93kZAq0U5F7CH5PptCxr2h54JW
2OA5mBEiDc2oMhOWPvUP4kt1KyBq8DHK9RbjW53RnQJ1hUcuLXv8ZsaCqdhYEPoU
kA+LU4YKx8ZyGLIPxSpMSlmZITXxlMW2LwhaY6uvW0nL2Q7tsHfG2rYTwo9o2AQ8
8s99sl7LFcq80D98OHZwuX+048aiTJduFnsIszsjYVR3oAouFvjkK0bPIyFlaQRL
9udCMRKKaxFqEru6mmBz91csG61b+H5uDnLwT2j006oeMEe3pHdvUyX9086+W9mx
TgOSHpjZqwy3d+zEgrNQe1u1F+XUktefLte+0FEeCpyJP+mH5P23aA7VsHVpqu6M
Uuo+29TnWnVSQiEs/JSa/tju3SdSXnLvp/REX375LpNkQRlJGwJ5/Zw/4SFDbsmT
QZ8vufFlUZjaxObe5FC6UBUdBr9WnR11k62HOrYUO1TMAfS3t6a+nupMChpBFJv4
f+DnzaJPSyNHwWYpdSXdWFdQx9zaf7zsjsVBLUVrm3Ka6A+kzKm3B6nvk7FBvXjU
scnZ1jsyZfst4PjcjbfgfPsjjkue1YoaXM8CfH7QbfpKbyxDrD2ZAK7k0Ig7gomF
Pdk053g3nS3M9vKrlp16VPPlaFcQnx3SOl7vyxNUPSnA/EPHenBKaMpjC+HeMfKf
rBn0SWsoWSaGp2E5GJP2c/2b+qEVP/tOx8d7Y7kjlXTydWnWXM4djCwup7osUbD3
wAjAHWEUqTG++OIaPNMMrABv708QUJQdE3lderDN+NnjE3AsGQ7p633umFpmOzuT
zZXYSTjkHj1WCjU36qtzqCakmRO53E1P4e7HOxjgBDnT8Mfi5dYYaB+aMJakQ7JZ
RYDliMjaJ1Ep//mLP4tY2XGku8lrx9ADWBa1IxgmpEHmEO0NG+fOGlV8bN5cMIUy
2jlFv4dIBQY5h3H6uNeRbh615j6MzZLYeA/63HTi+rDo2qmgXHBhJDvq+X9tkojh
einYhFdEnUiJvEYOBT+deOWMzlIlbjbWPSIMz5DAJg9B1lWz89Y/Dh9XIXRSuguA
nYQtJDbZD0LpzAKXXVDMhVGlFEpmnJLPGyjQm4YQ1+MoRXv7nZv5yc2NZ5mxkaEP
pDcXuNz5Y3tqH3UrbPgGRqeOW5L7uyFzerXmxtudlDSLTJ2l7sJeWxTT4asxMhr/
5io8aoijpUvnWubLA2D/vTJbU08UJEXCpsPnynMH8bNZh7lKPLtOnb60vK+WnwFE
kLcFqRfDknJVGrHOcGQyIWPve7veaNENdmSDe9E3PH4Q1EyTH7hbJRC/oU7iTmX8
elKrfhelORf5jWZgM1ldt5hvkNylGZookPfLZgO/bcLRso8KFIskTBCUwgm/vKXt
QaWAQJSgUxOFYVdBLQtdPXlx2uqm4ZCHTCqx0RoEQ+DOmKcxFUHNZ6y6P2/3XNPz
qoWnOfJ/rE2wngnVExrQFmOG9uhGjPoGpg+/8f8Xjt5mmGRywsWUV5GQt6qX1AhC
q6pXGIm4GgRreFRUxJwRvtKK7SKgwqK1F3kIVmLrKtOMKT942Jy4JbeZn3nVS50Q
v7UvElIyiJx9QA92Kgw5eSp4z5svk4x/GdfMNvjRY6kX3KcXOFkpc4ysR0NWmCx6
4At/56uoQvVcvs4rvSJFgCLSwO5JmnMhrNv4BLjOfVLRKbn/6FhW4XhzqDaiS8vP
7JCg8oFYxXtlXVrMo2NY4hww0ZTYbQc4THLz8q2F+8rTvaKULAyfxctQeYfqVwAM
MCfoXiQsQcJwW+b97OvJWlLk27npkCDmS7o8tcGgakX77e1dI10+rWHcmxgxf72h
VzSH2XJFOekSzXSKuLmj2gtiMYHo40eI/o7kDibPchiTLFXoZ1n9GzOAtzIW94gJ
Fy/+vCpXNYnVg1EvRuqvdW009xmq0l1K7sSexdcAcgwAga9V2xSEUC++23kacl3x
ekTE1p4Iagl253LPp7L0r5l75X4tGooinYE2prtsBwlvlYfHTq8YbuZCaAch+ZyS
WaXRFRigdTsq3/fwXV24PCSzJavtLqzg0f6ck0aAQRiAuqZrK9mvWycfoo74gn9J
+Mo7oMnUCfsF9A1LNg7q2bCAv8q3oP+1nS0gAq1otqF2zRU67cfXvQWzp+fWXqhV
l8+OAod9SO1LLhhcURqrGFLskLuOkYIvHjqWPBsPWatMF0ApTzxY28MW4T4ol1+3
S4/VRMoapEilV0zfxZd/d7jl2Lc5pfez/K98e6hL8xcDA9W+RBa3sKqESKlAQCQd
dSigyBU/UorW0Fwh5J9zyERGec1pmnCYAsjcEjzMQ8QCs4PGX2oh1gLjDjkTVBtP
iGglRONpCqra4aQSYaAT7oNhtOeNwoFn2qBYYsg5u3R+6GjkZ7oNdR9u3QpG6DoI
a34pHdkppQsZ+Tl8IaOaYP008bsVuGwbvQRXFQc4aNyM97bF99be43ST62DA23zw
4uuSC/EPCMibl69HP5+8C1S82h1wB497Sy6eK2amZW+HyhXE02fhvJCfVJVEU3RM
DOqIV0sSxkrJRGdkJbNrF59H3COxkFSwOmDo38iNTDuQlciiuiPgJDaKMVZKWui+
kX9M2/5S/lLgUiCc/b51dMWSRXQAc8rqdvWIFcGQab3u+lxFeOMyDftFW7K3CNhK
cttwgwev+0WT3vxrZbykbAzHlLcFF1vJE8iQ+wM9yWz5myOz2lcNMJ0d/f4R4pAW
m3dp2jNVHAVU6/xKheyexQYvP5BjxnL6+qxwGRRIq20HcGwOzletOs+62GqCARz7
dCW282S5Eu2VKjHHZF5irSZBRnukMuaDjVLN6SeKJ4gxiRD0vhhRPl+hEz18+0D1
cEJ9JezrJIWljf4CVMGH6mvSGwKMApPO4uA9mkjk4mLaxGDTldrYlV7Khqntq7ot
c6ejzqEKlFgA6JIPDD7kWaT2g5rhJIizJJwG6WpC7wQp3TvsJytFFZiJkKiWSiR/
PcGli21uLtGOtRuXLXvvIN+s5qccioKGw5P+2+8qbXlVyLpdwK7wCsbrfggwMvQ3
gei6ckkzo8aSszt+lMsfNfZ9luRO8Cfbt6EQqjOLnDJgmrF/Z5U2cpomAUUxhlfN
Z5RoUeWOGDFhvILs3oNEPx1l5GgduW/kzXlLgX5KJiv1DiQ5NjFNWQNXxdIgd86X
ptezobBVwWBE/1IKz2ZKQo2orPFxUQQ5JkwiDFpWAKIRHLjyKeXl8HUN3ZcQH8sz
YrHcGYfMU/bdFVMn8AZjNJexdXC+RqFGWvXUJu2vQNQg47Sl6uDKQhZgzHW0MSmZ
lKmWdqjrCA0izYQCU0mdj0AbmX8PDR4wqZ4dC/SqZrf39BmqO7Pnm5AIA0GucNwc
Sf4BOiE869TglGL0Soc3OizXCp+L/sXX35GYXljWgaqh36yB5kpfjnho0TVmzx7k
sgHOtP5wUcPuhr6NsvwGZ6uBqe5cC79EnhOV2OUM3VoU8Nd/14vwJZ6XD/CUmmtc
v+vycUCZ258+krXYuMckUtFtWabMRJBFimlbNDXv21oMU6XkS0uqodeJlf+RCiw4
5S9JFSPi7mqNBuFkon73iUv1ZJ0ExKgwx+VZUj2yZXDPaMvp3wRWpe43v0RzyKtQ
Er9zuYhWovlVLnnDWJ00J70ap/Pd2OVoLVfBoDIeLosevVPWG0jatduVc7KB3q52
NruBIIARPX13VWS4S5wei1Izzvjrexb5RStS/KpEPCvyd44ebkoUR9EnlteGte9r
B74gBkQCJNLmpDS1BgV1Uo9I6zMOtSbsOOaJsDZe6hRhNXGEobqH1xtykPvNDWm1
IVeK3NeFLxaB+0BTh2728zvi6Dpu1MZXE4cWP1uk/CV0AsmWXkVCBcjYgSL8hTC3
gtAzli4DNNt9y0nM/pCmDIXyMob9yI5xKuT+NWZXkEEs2AhpBMMb7MQ6TPU7Qtj7
QOUJshOcbO3JpGxGh59lFs/TPtW1EtiSARSjHXmrcQd3oA76i9sqcEvieXrDKru/
qQiPqSKG8b+qUQxgZZ3euRoJt0KnQnjVxu18m0qNJG/cKr8+NlKI7tgBg9ZPjQSu
NEN21AtEw2Km2eKPpkWx0R3GOqUZnHuikdiI9wKvVAgrhmKYEQrBGl5rzkPpLcE0
uiwGlYtTxTSoW8bMbQ7T5g3k+5pASQic5ZexM1TL6WmgCDyoZIjkt6+DtTSTuMBo
lLwHcos8vqHFkxvFYe8d8NSqFYA3Tovcv+2rHvca/wVAVYkVl48KEY2EqlEe3fkz
OGCphi+HlytDTmyk3Q0EUzurYdy4Y41EtFdob4gpHpRBumrV31umh/WSnEYZHbNa
NUNmYjvYtuanTqPDNKDaoqSLmvmtGWp61sIa0ReC4LEG8U8s40L2+my6LQgvZSZ5
B9F7xUSIzTvCxL6Ej8EYmntCslL0zYJ8HXyUVTQqryJl0ahSIZfMZrW7ZRKALc/o
jSJo3iG2lX5xjlFTkyiB+yqsJtMiL1UANtlcm6R/OqilmPuduksy5KFi9cyy6o/l
Nc35wNeEWqRrvHsWKsNnnY1DtJPeVaJklL27zyXt/XGTD5CM9lJWbphCoIGh81Iv
zPtaAlzl3gJ3+ZD4uNDO0ciKmxYb50avyici+9RL2CFZuJjqme4+OPgRetERnaWG
lGvMuU2h6B9XQQiiix0I3lPKOK0k84Q51cIS2vAfi1iPc32Jf8Hmyh2g67EDaWKT
KNTo5QUairnhcrqPS958aSF2ycJGTIrpmU5S7RDsSmt/GR2GFdvxfbBQ6Yfm7i+k
aRs8WNvnfAEvqVmnVYNaTZDkDKMMubCCLslOmy1GQlxo0YiiHrIoWR4NGlrXXPds
7aAx+uRMngwchcZQ3rlmtanaoPEKvVKHrtRgrGTuYJ6IYD7j8P4+7kz7oPgh6mTG
JdWWN0wSSTQFbsKe2IiIIWPiUkep1vrCuAdkxcPkHstbgw7epoigLrQPY+ztZP1Q
VzQ2tgO9vOGLXRQSgAvfsVv6sEcvDmJ+e20jsIZxSa2tvbRWNr7tdxo8er2jBvg0
X09P7LQM5VOK7tuNtssdsHJM4lqNNP9WKryaGH+0E9gT6YDVWhqvElC6a5yPYB/J
/vGGTOOWA1V/xPJerOwMjc38q6uWrwM74cSK6c6A2LKM7WVi2sjlWrmP0PEVwoXC
gXDGFD8WygAb4enuImbz8WQb0u6DbvrEKEVFUMUgAgK7EV1GZyqWotCi+rVfZDg1
cnh0F2tprvoXfY30xYoobqDcO9AP64NGzpQMFi8gW3QyYLFSfAN4Knt0HFXx5GEE
Jke/sLDf+RtMwyClRyQ01PYz5EbeWBrGBUqMDxAPyz+OfFxZ243F1EoKpbklobZ8
S8Bszw6UfEBKAXSBFnu0ITYAW34sw2u2sFdVHk/6rTKaINr0z9sb+j+Kj9VRpTQy
OlV8c/vJoEyLIS+ellBNmahKzwZx9xhZ7qbb2PzHBtybtEMvV/8KcmOP5gWAmhMe
x22QCcmqgOZ38kQmlXXIBlW36seZCdU/SdRYE7mHfDWXCTElrm98v5ICGPNjBN7e
rttz0mnfrw6cGC5nCLp9jWhIMp0qEcqcCy8CbE/oZWrJluMcZfWVeyJPzZufzfKZ
QKhbRQw7eH5LSJX5lsOKyAJaGwBvVemL1OmBWSqxqbEBcRTXZU9BK5d70rLs5X3K
Zu6j0fKgvyRRJdWBux+9cucZqlbaFfLi7ed0LUKu/JNiiE+v+2asfMmiwa8F9EFe
MvW+2TfGSaNX7IPzXjb9lzNqBK8Rlz5zYxyPxNS70+c7LGsbJh8a64B73uPNEkGu
3JvPmJWnxgJVHMksbWvDSVfM0EmwGHcKHlIn+j7U+dTNRL5OrBCVRk0APWPZukzG
WJ6IQkDxioJWaDNr2uLJ8Opi7qi8aT2jESDg8a5GfBQOViInJ5GXwwpr8GzVQfAw
kt48TBNDCM15Q6nA3MtezqO4+tjuYFWpIj4XtfyqKe3NOx0EUJav33pRZupHW+AU
j8iWodX6k7t9oHYqVoLmvBlYcle/8xCS0H9624TjB7zZtaDpJgl2mIAlU/WX9fcq
hrXfMOQJtawvzp1j7khH++MmgTD4AAFtFxybjpshe8lhNzMglJ/nPd6n6j0BeEl2
GGSQN5HcjlqgGanLfeDVO+n9dzkIvgBd7Q9k4LFvk65FXFvC7NWwIXDtnxTi+pnY
3KJy5LoaJeefEqNq9+wbVEZ8dJePH0pd6lSMdP0oV7jjc3X0dFM69pmcv2zufN9d
OPUJXrRsEZcwCB+3wacFwSq7xjzXtZAFaqU2KuBgO+VyJR5Du1s861v91NLfzwzz
5nQICVpoSc360A2+unCX795KkXcUFEsocuN0+tBkifg4SJ5XLXXaQ5tGtI73pVBi
7GpSkqZu/xoLGHael8SUHLpXTgxJLLSwIZ66BJAhqX9hJTd1k956aRBgqThHP/E8
HvqBp7U5q0RKUXZrhagO0izNX6nCdSsqWmjlnkZUAAAO5EhZPYXVNt1g/65IX/6w
Igf3byxEwnBLphblJl3oiv9dtsnCYNcfYG9ih54EDUZ4bNmbOmEJCkyXvw6vBLCj
hYFVakaH7Dcfb6e/rGXsvKJdoh6uSB0KefkfaRZ0mI/totJ6xZyjPOsP/NGxzXrk
38grWFZUJWWnY6mwaGMWSVA4CVfj/uAdC3N0NstGOjBIrsZAJA4COh+MpqILwOyg
sqAjpR8WzmpQ4s4bXsZILNCa3w4QQdH+MqEmEtxEdHG4wuKay1A5g8QNt/uNAZpU
TgttAGorvJZON1iA+n+8NbMJmixlTVV2bFM5KYJlhHzW+Hhiv8RC0yTd5gxE5mcn
ElKd/hOfqDxi+SC43fqmWei45jiSbxIytfVVoao4IHRPW6S04gCWTD0R7XiTEA6b
OuLtq5iqua/ND05mj2iHaQfQkD3mParYjNLY7k+rSrpk350R1jWKPKrbzi/5ZyDt
A6vzeN4Bu/juBZpGXRqBzwdNEN2Zq1yT0mu5/AQKqcq5L8Zj6/KznGa+mqEZiPrn
i+agUF6Vwu9D9V6KEc/uOrMiIeGB5/3PGiCmOwhy5ZC7LKXTHb58NlEM0Qlwnv4r
jfP7DICv6pgR4AM1VIbFZAgfm8CkPDlXvfTdDmc19TxjyqjaOSvZkhVFdp1AwwE8
MkNHIcL8o7+ohpvqk1cPe3ebEtt2CRi9UqdZEh41fyhfoP5ZTM2fAxg6VezAqTc7
+2LA4wdefSQtHPEOZYAX+LcezpDmHHKxW1tnlE1MZbEcVcXJSiWVF2EIPOdy84tH
6ISJNGBsLKGI6QicajefsHnNa1nz2xrQIy81gqZUA81duLJrWhdoOEmRUgEMNMsS
bxnlIgi+U9O5704uNl0Kv7GhGauxI8Wh4f81b9mraYXiEIJrfGSK3vi2YLG8v5nG
wAxQVuKd/isJUP4oYhzkIIy6b6HszkaVV7J0Ny1NUEFWvX0apsXlH2Xq54C4Y59C
qm6BkvNmxlVJhF/eKjraqDRUYkGl7nr9k8I05WB7Px0QeH8kUaUpHL66Zwy1cgEq
Mz9Bfs9NZlLHLPKk3hCZNA5SzlynZCSHY1PfCJlEofdZQVX56yUuGLr/OK8rk4Ew
wYTc5q5j/hRRMt1OeoUNNKHBl4WU+G4p1vs5cOvdBxWhLtvNjD2L8AU/xBElA2TK
Z/tlhm703oygjX71Ao3x2SqyzkRSFYUvIyo1ja/ElfI5Ku+Uo/McNZKMFMDGkt5J
dZd52BojGWYIBnLuYAsbHwkbodNDiZ7zvwwUEfqNPV9rl3uiau9met78LFlQYpYn
HiLzC+4/hFQn6l3wzS9Am5SPxCnu2HkkIY5VfVGjmMy/sLSQRWmSIii13X5FgjrF
H42h8W62Z4JO0FT5tY+NeUzLHBoqbzBkjyIBBqcoQrsxS3ujQ88B8L2xy2hwOAfg
Iis7M2qAPb+h9BP4N+olpuuacCUCL6tJFB6nBaB2fFhxWZ5FbRQMZwEun0oJjuRR
dLf/2zEgoYS0a0PSg1eFX09QBtFc6AYiSjc2wZp2sPdNCdo6/HY8EWhLX9LBIPId
nQ8qMrlNgA20Oz5vJGqh4gvsYCK01YcI4PBTiCrFaxI3MtTNM6UpuKL0sfSAOwm3
qcKboRb64vElf96s5oeX7Vv5iCmckKS8UT/zqFQLFuP/IM0l69s5qrizRI82T2So
iaA3BFpoPZyf65UvVrXYpZ7dp5fXbPTxbLvww7kbXoIRDA9CDTPtet3k9k+lQJ9J
JIEPLILbXA+RHwR0TtPuChTG8JrXLsThtzbECJuI2hH26Y2ZYGeBpaWnYpPPknvf
JKJVqI9xJwA48k7GjL9J9AcQbYlXb22Dj3b4CJ2YaHH6mnHAnYYAp9I+9Twvq2qZ
hOy3D2MQTNscUoc1NniGDE2ISIrGPUsFAiYg61E5voS+Hq2qIzttDcFtciTz8pR2
ddv6kjj6ppsSwTh6KyE2cpTdW6K5OWxlYfFFak0NAAPeScXJ71ABRL0CFrcbKABd
92Bjcz7lSyNex6Jv588SgvgY3QcX7nWLZFS/kgr/yMGgCnnYpW5eJr8Xn5KyV78T
DZnDrSoSBMcEl4H3FAXjX0/hOpc3KxVUvwMCWkU3XH7XhDR+1lbm+cZ9ueWBVyu5
qeC1BIoTrzGDBwnmK3CiVBQwwzv0PHw8S7xfrhLBlI6thRaUpHgq1XBHI9oR6Z5d
/Vrab+P7KqLtKZC6Y1lac5tHb9ji/VwIKQ571sV7l6QFJtn/eCU3G2nFLK/qy2f0
o3+DAfbiPNcPStUjgxJ8ZAsEJ8qop8par5jXhCLpTmHsD3WB1OHZPM6WJB9+0VNI
6SOL1OC+SodPbPHTvn3WuQlTrTFASbL0GPzAfY8xuCuSQ0TTy8Cyx61OVzghGZqj
nQuTlJ93kIW09FX3ITnfslSkN8Ie6yDDTsIFtDF5ajuciKG+URenLecWdpNWwg/h
wvOEDilvqFWe4EJ8Nd/QGdbtyzz5WOqpKD+dvXhzMQGvjzUgjsVahNIqK6xunGas
iFo8UnEHScmJreIBpi8PiwUIpNSIx6miRS77+94AG8/lLPCzEeY0EQSEKNRhhqep
WSzDuKThTwHV38hYEPl242hxN1wc4Bulc25SuhpOZ+UdPKzkT/zEuxrRO6AP9f+g
kbAJHHhZBWZin5hCLDn2XMzMZ6Tm2wm5DRfO85BHgDjQkJPrxDQ288w+3J71nTPI
3/qZ5lgL0iURsquqOfpDz+HZxD5Z+8TvPLbw1oggfyqIg8va5J0Ff2LMunS+Vt3h
gLNbPDB+u6mFtKXhlk4k2OuJNHmlE27JDpnHGEbeSaSs6dhg1LXmafBkmqgCSO6h
QZsrfRzqKk1v+uRhBVg8yZP6vS5zocAjjCm/UeS2z2orBSu2ufJU6nGqUnuJveCg
GebcYu8TEVyFa5YpXSZf9NesClk3guJRk+a6Urr7CteQJuah8dROmVgQu54WrnqP
7dam27ugH9caoqowv2A+bc+lHa2F68Jgl4lJ4AtlTQau+K/+zMfyKWtCqQ5VSd2/
DTpMg6gfcGTdHX96+gxbVd92KsPCXK2CaaUTeAGZz+zZK8hXRJlciruq8R+y9qLD
9nQ8jwd+SNy0HnGxRR+KmRcBS0HUIvHFhtVcMdE9ybbjbNOsiQGBQ+unwOacZy0o
Qyt3IaJnuYEH82w27gtJknmtpXAWbF9SuTMbnQQvMpKyUBjxyw14LJrOsoMEgqLw
VqFe1jOvJZWVNHut7EsZXb5Cpf/XzdGNgFaWJsuEZTAtwBVyX+VSStJ0w9QThfPT
SYRIJgr81vbkOlAsaUKLsL03uQ9kG0+DodsWFcvHtR6UKYqa7yOMee98sMAovKgl
Fb6bYQRLCkmmGbglM7wBzhhQ4bBOLTDNMkc30RQxDecyXf0691ssZwfNQq/8EPXt
oCCPQJhFVUMrS413CoVvN/7SWRgGcvyNVSjHgvO3J9FPNXyZ/3PcOVum0+Y0Ps2q
+Cn/tTgGc7gnWjNgttyTO/xcXKJDwYIWnDvrmtZ4H1y8yJur6n2A1TflIPGMttyH
EwcdJBGII691yaayogqFaUOFtgFhIXJEusIR+KChKn6oLxbGuYCqkocEECyu2e+T
wqrI8QvIEUQ/vBnCCGcfP5J7qpLhrLHX4jqELaNOX7ybA5Dc5l1oyTwL08S4E4nS
JZDIYWwaWrKa26NNsEobkov6BOWZJm+2ZrNEiWLgIFdZYbrajzLDpwLpfj2fY4+1
EvZ/Y5usHONK6m1XDfQ3uLXNIzV7awSiPiQDZb+1kV1opD3hahHavq6US2qR4cTs
f5Pt4Dbbekv452W26C7MvhrjmuckgY1rbbLYv+VlTQeBi/o1JAZboHXO9juq/4/4
GV4evVmfNwQPToBpFwzpc05VTwYL++XSJcX7PXVAN9B+uSJRCV++GXB+O0VpkGpz
AXLrj9D2nkaswgT4UJ7DSgnaIhIH66OOy6gdf/HjZcTM5IRbYBNQv7C2Blo+5pRg
2wHyqoayV1HH8HmcTdUqfHVi96EyZqW97fy2xJGLritJ1Ll67yG+h9vbU1Wmg2J4
5PrwR+FHTShAzZ/vIK61YFO1X1Aatt7Tceph+FnUVJ9Mxfy9KgOwcxbDWiPjjzRl
hrz4TEmaPf/Q2Oqa6ECvJpIECTfuHPfk1UE7kTm5ZXONklgAtKsNgl3HoQeaylHm
s5sMh51JvO/sAXcMXFnjwpMPex6TdP3vpzRhBrii7AAFGg+wJODMvQgVjY51ATT2
cis115ZZxkemNJQG3VRM9Jk91c0hguBRXSxGGziMFjigiQDOWue0mz4LVZXkoGOw
/5MAizxq00ZwaS4QWtOYWO67q/okk5CSkqNwTdW5zP1TJwZVaLUjsmKxG1FOtzm+
qciSHrDtICvdltb9L/6j/Xrsvm01LehgjN3hkKbYuflfV3wuxXq/c+jIVa8XZan9
wMSbt33TfqJ8U6Gn3bXb/vAxcMXRyTIw2V54o9L6PFewzs3vQDo2zw79Bs9/81b8
LrfeAOz4QFPpQn2xRB11uvSq8+o+o1RhfkObs7dtaOR+gpIIwEO2Heexw8kZqmux
xXz/GJ2MvSIuYVzgArJdwItXd8BPf7QjjbN660xK68fa//l9k0XNPWVhC4iOR+xR
bPhJUFvgFlrTx316hwflZGZvjXjTMykXHZCOfl0OkG8ynuwdVxohM/fWAQ8YhWCy
Z6XRhukId1Neg/b5CFaDVob6f/6rRYfLARfXrAdmCrJYDOBjXCz/1ZT+nD+Pl269
R76kOAu+ekrVORJ6+XgLO0I8lha1B80MAXO+CVfrKSnC2zwECK7D21fYJHe4K4kf
3yBKRszNBE0DmSs5T2w3obV2vQZbbCw2b0k3orol214rPdg/78SUgOdG9ngIbLzP
UaISwIkxtUrKHojtxvqgAeyZdxM9Paf1Ygl73kiowTU2DEVagKuVIP++EyF1sTCP
TDBGh15CIQcdgCCsdv9KbgD7ZyL/7eoxGB6bwGuKeG3tjKcoZJybL+OE91tgenSO
ryUIu12le9OT7UN1Mtu3GQxzvNM7ohJaCM7qZDUhrE6Jp+o71AtvaTU16Ogs/v8A
PUsighLUDYS6KQEvRiarXxsTUWAMGT4xooPTS1pp+TLioxMAu4TrBw9EZt7uOR7T
zXwF0x0D41JIVjMneigqnXexctWrmKzBF8PeL3X1+NHhTbnELRU1H89yiS+fZniU
FKxnRBuDGjsW0zufv6Wd/am/hCX5U/iZfihD0fn82UuHQ02iE6LQZ4PoV8/lYE9r
vgV7lgbJVsPf+mWODtGenaAbTj8YuDGkLoHhn70SW9zXkw9SvCnDE5xKr9gGYIkH
bnYsT5xoTXCcH99E7gtjKGQEe9CMpPc5ZmrxqhZJBFYTgKqttYqmL1nqj6Lu9sed
NpXu7Yo9owKKCTYJK1YsarGZv+VBU/dL0arEuiwulF9cu1OGyi3Xke7+FDulcY9y
GXcte3EdF5H1uKn2igyQhgBYxxu+ysKqnxRSHv2vWt3Cg5G0nf9lduWGU0FKRpcX
Mf2ZK1lzXs6xrDzhw+v5YiZRFEKiquu5bQ9DX+Y2Ua1lkuVfozqNt6Bgbyq3+HXW
OYh7i5rDsX9+mGOprLFh1ozRHNig0A2rTcvg34cW5W7yx2+wJrxbqwOrGYlp8bWG
djN5zgUpycMxHHbMCPBYbgotNZVi3ExvZ9bnEkQ9pJlKBGCS2ivmYGubYeRTpHiR
2dXuYhPZz4J3kTHv10IZOf+9vCLXUzzQGOhyQQlCMGsQXfd2Iu8X+vGxDlX6Ji/p
68ohvwaKl6enbrl4GNKOrJJcs6eBfagsKvGz/9GXWOpKVowZS19ZHkRcvE9zT31f
ZcIhpdQO94tESlKPSTcHuaR/DkupFUuxBbud2tm1Tld0TdBnUPQrJmyIg6iH/NS+
czbHYwoKI/iHZx5hI8U9RBrY/nwyMM7mTntI0mobMC1HfmIPJlwABONlJQ+Kpj1r
oYPeb7XURKIcvwrecDUKy/03EPNluHRs+OZhUXWCNxoevLishvx/RTxRCIsSHHkr
tI0ldPs+kY9g7PXmRroJXMT48oBq7Aj1eekLTR4H5OsgGMIn+2szDxVhrJ53cmlr
IJgT6H3sHfexqi36f048oK8/NkSiA8m1fNwx0RwWJ3MZyXDRRGoS+SRoDVMXpoG7
J17P2Kr0kfkAvAoGLBRp356vylTB7YMkjrfOeRCXpbAiwS1NXwT5LIUZYswct8GX
IxIofH9//iXnuOsfBOzblvNjBfxRfzfUXIBTba3KN4II0SqM6qugo0d5ycm9NflW
P7ItBqwofFLPbIm+Y9giXrP42sEi9wIQgXKt+PPhqj7in2NqlAkH5Vu6qS1c4aNT
Ho02/7Mo9IMOzAcTjf+VZ+WYlzKtdQIYv6725PkjviW5nRQQueOIkzgMmY5Y836t
kJb8o75Keh2nnx3m3EKCNbI0v69zSWvHhQg50H2eNeubDHn6ruKT/96UhBEnmU7y
rh+DYeorX946OfyTFrF5rh6KiITIu5i3Mp8gf7rioLcvUP+ZFky9WUMtEsxE59bo
5xdMrnnJ0vcg+Vvb03vEHgnXJU84Wv4hpRlpta3uFscSJ437YcpkzMq1ZKVfHq+x
VdJxbYII+sEMiOTuPv5uWzCnW7cb0IGK48YaHnInZx77d1h8r2xn/xc1XKXyJEC3
ip8q/NJzwaxDLRvnibUa6dNyT3U1Wy3NxkLA0x8bBCjDgzeCqdQ1yncxq1BypA+x
W9lfDA5afgH8UETX2RmMFxW/h3BmCCvftP7ZMJljvkqx6iae6pynaNd6DUQjuJIx
QORWPVlcXFFQkTtL8leSY5yRo9BLPrQMsZgCMJpOsnzhGHStaU0O+jOyY2DPzLSb
KeCX2ID9IJmufqZhh6oB4sRaaBV3WMMUh6Xso4wA8xRR+s/mwC7DAIuLvlfYEMwn
rQ2QDRxrwFJmzc5kwvO4ww52Llyevco2FHmVhVzM6kdlVvIwJT3tS+lW7EaPM9c7
LBEIGrucvXUjYmHBeJ0osUEaO2r9+J5uE2vSnoYkgLcuejQaeskTNWie8Xl1/kLR
Lu8o0l9vtiSBZwd+f0eBZqmfY/8b9fKrZq24eyFDcbRHCAW/Mp1VfmB+7vyMHgHX
OG2IqFt+Eqbay8PB2+w8dim8w7NW6EuFcsY4Bvk2EurOUY8eb4EnkFGI7vL0GYl9
4LK2U4W8gHG5vhtpx+X7HAVytS1n0rySZPCsru0RP3Nkm8JlwKCuJPk/MeUyKdlH
scrlCKRuzQQUtsSLPH+qfuSFTcm5RidyYUgNeokiXxz7NnW7SxIlAnA5ITvbqD39
X7x4CQF0CRAPe9v8bftsRmH6m1u6G6buDJDtj8GBrQTBHzCWaiqTOfVbIrx5b50+
k+U2O1lg/axw8s4+ME1ktNiXo3SLNacPi9ZcQpesAW8fi8MLf/JSnW071uFu25m+
c4HYUsXeeAaO4LpBIhVRPD7BpfKESqFe+BQ+ROFvgYwXhQxzJGxHbzOGzVi0Q9Pq
pigvqQkUPZjlXLxtEEmINw6SgtMQ4aF4NwIuvlj6pE7OZFEPvnTOA1DmUHjA/eDP
As89ETaPlkIF9DW8WY1KgeITgNRUBoOqCrjSVRgzf37iAUZxQbXklUImP3Rw7NPQ
VYBkmRe8HpTX1TbUBWpPhLkXp9JoZi9eq2z4CpUwi4F4zBCi4MAN0I25CXwDxX7Z
73lIg97xUkk923CILx1WefRhn8khk/DtmxFzzb+JOJVePRznQjfwF1QJrROXdKm3
9UZ9hLh7KH3ftAr6cyFU6+hkfwmos4k1Ig37iJTpvb4TCIQ+fMu83jJ1kvJlT3yN
ssWkipxLL1DUOF4g1cxXTYB4X8FV8jon6gQFSzmXLhJAtd6Laj0CetYTGoRrHHJ9
Rb51V8Kb7uTfeqhS4Cn3vDE/POFh/9DIeYhrdDNxNFj05wtVGPELKvoMdwpO7xFU
gkvP6CQlfVoSbZPIvSg+nqSZRgGxc72UB0KOy2vIKHqj2F5opga62g+uL5c+fHVn
mM5Kai5vjGD1CkaK62KcJb+9KbiC5fMzruqAs31uajNYo2vreLKuXRltn2B2VB/v
1eGcSTZc8O+ivBHEyxIB4O5UtUCLqjk6ss2UhbYL+P2+kueM2T/WDh9q3JD9Xfno
bRE37Q9LQJRR8I9Tc0r3hTzYCkmFp2q1zwnqa7MTF+79r/h1172hxfmzlyRukq/J
EpZX/tj1ODGm8aqn7S2/vqStdgVx8GIvwWccu2uNP0UoITHoQkfFlZhyGhJgV3v4
96H3a0Qy7e4pdbxCFaGRyRO1gAOIgnHjbpWIIe9b6NYxy/Aua2iliiFSsvVOmVak
doHMjVbh1iJlh/wUSxlmHFc7bhMCm6A52iijerS9fKU6F6LlgJh5y/fusHbe8iMl
B/5LdMnelisN/T8ZZvT0vABz+obyu3E9A+bxC1EpJwOXFICu9f8nfsfgWLhrnxbQ
zcOLY9Hwa8HOsVvaLRxZIz/k+WtalC1uIRbJMCySDYfaC2U7KzZE9kBYrozXTB2x
JX1Ltd1FfIisD6P0LGLfXkSFvcbLBOSY5eJOCwkjbzG5a8MMZXAx5bJS/Sw8WMB/
uU+1SOVqYpfpS23pr0MGb0Rbgjp+qDiUT7xgvJYg5FrRgTuFoFagvvggiuPhbo9p
j/O++j+aBwHe8qek0zx/y2SmptIMzUomoA0F/ITh1S7WaVdTrqw/YWZvbiln28MJ
P/V1TQ0ssb3vIWGNcZmsQV24NYqneBIQRfRo9y4hkUv0eg8G5I+h4MaFKkPHKznA
LQnNZKPry3Qh3Q53YyjZGspq4QfEq8bogFnbF3IVzzZw349KS+sNcYbiFxhyy1zG
EK2jjJgVyxOGCys1wo7ayEdG04kb98hamY5Ao0Yu6jc3lNHEewLgqTMkWoALGwOa
Ujf6y/xJMfAVe2yDSHXwBqxLy2cmoveBhokWwzXHHQ5/ep19AAdfcsikrxKQe4n0
nOXVCO/R8zqkMDGXinzdFZDivgausOKLQu3hll5AvCEQtF/G8rzkbolwLoRN4wsT
z28uW/amRni2LL82gElJ+Gr5JDwN12L311hOuvl7k34IeeOvbQS+E2I3oGSm0Rkd
6OIJ7BivNlRA82pGMFvgqytnoExQTWRYVx34t+thNuDVsS5au0fD03Se8+ULZ/bT
hTMa3Nj2/OZnEzW/PDVXKHwBkDdlDSA0x0skixLvRql3R9T/Ivt/3Df/UfZ0IbhB
q3UVJ4XsSpafAK491ZLgAW4SLdJmuNy2UdDB+hwhAf9zO+M4HRjORCgoaC0/GWXK
ex6RIepXmxMUqcX+O+yazqR49LfLJlxAlKAxfeFo0iBaINNIr2q0MwieFE4kkP2j
nonb+U7It1v/zdvi/dDt/1yAdJ3BrqWdRblwQde+3IVfl1S0PF1ZQTfSg/mZ0wMC
3x/252bZbH25//v4F3Gma9ewSPIS4s88Fn4cxVVQhawceANLFS0XCbpKKW7xmwPF
mQhlI1Lz12Xtv9ArOxE5wdjHyKkZwYxqimJcc0no6Pd4OhKue1kXRDnOXUmnaiLF
09taYwVX7US61dfrIp47g6vWBxtoyMqJEhCfzOhJ/BQvgmvl8cm4uUFYocrLxVnP
P1irWUD3aoZ4pEaMlSdPRDiIz/rqMD0xSBcjAflzv9pungwbk3CEnzry0tXLtzji
wY3hFvmObsfgKwcQ+qGjZYnEwIvzYS38F4T9NXw1eYIKwy5HrVTSKg74F8DYogqS
kDH+2HBdz3pFdmdbrx/TPw3P0pgseZSvWSnHy+XTWW+ewJll7yXfqhQCZiJYT5y+
4hzuAA1ReZ1mUpnUdwAIZ7tPqQB8bL7+9uijw9iEj4sWLVqLOnNLiM+JlSc7s5So
OStP5XUQNwljroDI9os0KiF7521o220oLNuEMhbj/82H23J4QKAGAwR1XiAxkiCW
6D1gNgI3aJij+NUB+y30HtsWXbuCp/4ElFSBYfgs2Izdfjpf9wN+a6/2OjYmQF2J
AfWNv411Ho/+86wgSgDpVfdoJIMHOTmv+AEAG9Zsl+pGIML3i3VkVpitrMjxMU20
bb6WOuGBPorYb2v++fRrOYWuckmBrZyXkpUtPorCNsQZj2q/SXOUp+0QCkfuZUBt
KlDaQZ7/pNCenFHW6mlE76MsXvzJb4QeVlVskNVMlIqN8A15NhvevLOFBRaFPru5
LKtWq16tFGoXpMVpRRHRUH0HRpN2jr8dtss3yz8iAnYyHyZDxgI6CT98QW55WLEO
C20hRnuYngjgYa5Tm026A5yuT0eY0kqNYnklysv5q9SA9ZwA9h1oG7T8WQtGzFW8
s3UpqOVFhmL1jygJUpyXrupA9s+SKgiVVzCsGbn3tkeYHTf2QaptEqpp4eelanWg
2unF2FQU2zUELN75yWddq1vtXsPHZBD3prPHSAUXTBpleQQtMH5lOytA1KGXx1Jp
npYZKj0XyUcVXC+VONDgEFpI7QKKWnzNRXdCHYvse/yX5XBrnM28N0P6aL0ohC/k
tB8CLd5vD6ryKs8wHvYKj/9KnHMQaOkpVhlv87yYWEi4Ra0UI5qegrUnns/Vd5O8
xina4xPXXuaEehqvSTp6q1nxJMlhgrEp/T/ss5OK3l5n2gCoi/qI3MBCvQUsD1vd
TYR7DsU9jTQulHshofD8KKD5tK6w3itVFgPCwZH6KZbQ5M3OCPy+GkwxcDi7wtCr
YhcjdZK/wnJNgFbS8VRcU77tF3s5I0gYkbJTtwsjoZPzzo54dg86Zz/RVMxmNwFY
J3UkoIE0BQchGWVRddb9s/dw03BuVY+8CZbv3AqtCPxQSBH4qH2WqEAeFwQ6mfcR
+Dif9QtTOqTTMonNbEn616hSNjwjcyg/P89y2udw3nINJOfFq36OUR6VHoVljdd5
x/izDedDaMKCQest8Xh0OsE/Dk4MMKBl11Ps6iMwzflB63Wd3bu3jwD4uz1GdOPD
T5Srv2smC/JwQqjRMlSqoc4/vGNzIdFGcSHa+9vzCcGyBlGfsPQTOm3Et9B3Ytq9
Z/YZxzGcdKr55o/yN9pUiDgBoenwYpcoPZF/9JSfbkUjQ1KnBZacrS/tWk2QqC+d
zlOmuktKQznsx3WIU5Ete5j4mtjG+7T34oe66T7jCgnTB0g02qGx0rvnYBHWA4tE
kNNtFIepqigbdEkRZqQbaETFs/PVg8qCyvOTGVyd2na9kG5CYEW8klyxFmQ19NZW
ezYF1CAeZxJqF4wecKLZUE2EuBdSyHeMvGgLbfQJgpQAjrbLtZCK8Gqjo95AVg4D
ZYWQAM0WYTYCI8zbkcV8/0yJqNLwoXlbYixhHwzgVDBq8j605CV8dlfsxrzSueLU
ATt737wgCavsf8cpmDj9WQ2ITl8ulKqG7bGUZYPVGNC/y3EJxYWpd6VeYvFRIRfp
+x2FYaJeJjv3VuOBq4jI4Vz9McBo1WgdzsRDpzdVE1xj98v5oBJv7oqTJ4aF42OL
S8Z6TCBKF1dEa28VRlks5hVjJk/e9f7iausk5LRaNq2VjqXMNy6TmVbAUXd6Mgzf
yssJdWlqBUCh40IVOMIPMsSSLiW17XkJRYR8dj3F+QIrSQ2S60UQc6dQ7URg1jQj
cSggicUFuW16rAMh0SKz2wNNTOPHlRjEszg53vSmgYgd9hose3wq5ImM3Phhgc8Q
QssKy3Vx7rkzAhT6v2fk0JU69NB9K80WaamMeMGDCuYPol4vad+MVPmMfCxqbF2L
9n2MkV9S52K6k9o+2lwf/UE8xoYICIpIpgdl02aYPOKiuEp4Ya/gw7GFsFAvNOWk
BVQOtnHjTKSgLRbWeIcAo+1binkK49BZXxO7b8c/H+YMHCygpl/avUa6YfEUwwin
Wb54yIyIcgJE1Gjw7gU2YPhbmxiwbzb7swyWDTlmyx9LVoHAN2SkMIbgxHE6SWC9
SY713q9GyGd4wUi7XEukyjcI0JaB9hTn99d9yO0Ct/jUWnm+7QVWoptYd0QOOiST
MWpeylD+IG+Zl3ILVjNmlKXqFqHRUAOXXydcLhoOWEB3x2GF3AyvxbcNC59njZuI
2O966LnKCUTAE1KTvGTaOvvf3PSBWOJ2onS2ffVqU2gm2/9aIl3ByVDWSdqzA4Sv
lBaE8lfnkRPVGPmFjiFg6h7+EjQtZRXPVaJRJL+7XbpY5F10FmqgNfJ5nwgCSwHn
uwaQF5G5Z+Oge4K9HjnDkwbbtT6HJ+MQgARW4m4ggczdMkbybP1YJK5Qj53HikDA
5v9S0m2tAZc4cnTIDBwljGBvQsjsBzNBiq/4qloBkt/J7qbyAnMFkkZNEH8D9oLB
ep/JI8/1cii4GGkoMqYWUref5S7HeqrgDqjwoXe74sD7Nuhcky5d4seWpZ0N4Chk
rk1We+5ztX6TdpmyxsIOI0XyTizf+hgBcLQHdg1pmSh8gAMihjyLWucyF/maB7+w
MsXO/T7pLhTqRC5J1LwB8g7OoqRLBqoFxknA2uvl8r/uDd381l5qoUT9wCz3ppcp
J54EegIXfojMf0gISWWGbW38mTEB0RK+ucYoAkfqzTmYbv6wuXb9yGpY5b7WEtrO
StsjhGuGXVBpvnZOpAOZ/oSZ5M4kzRKsZph2Zja21AtKf+rDSdXukXtlhU2O9D3s
sELe34PzYxrMujOJmmISZUlXucGkDWHDLMosnulUZ+c2ciC5G7DikEdJxleLe4Ka
MPFq+SyBSurG3V9Ceums1LQfwCpeaSrHkO9i2dyFXwuhUVU1L0APRuD9FYORIQ49
KjxYSnYRLhn14Qqlx78H3kR45tBNQFt3/1JMhk+dy7uI+Z2VmoqD5JJVRdiGQ+gX
0nBGtvDwtxIoG3nj/9NNkroAD/S4WTx8mX6WNvAlzaFr00ev70HjbZBy8p8qNOxj
snfM9Oi4IaoRwDvuLn1u3+AFFrIRGFRTy4pppR8VckIylkdv02OX6PFii8ZfkBMs
0JcW53b52Y+wOlWP/u0jC6Y/IDzkcyA3AZovza7pr8RJPdSEBpiTxb1ib+AGryhR
A2DTU7tiDZ27AvMCzIKxsQq7exYUQYu3/Msv8o/gzvocMI3QNCoG87MrtyFz4KRY
WZfpNpAoqnCBDuXKZGObdsit14I2jRlialx769yjloRQsq/esZebsBUa4oxwdtEz
22BZX0h9BzbvQx/tBDHWs9q5Y0ZmkR9e99A/1OGgcJdLm3ZPWrPD4/vb5gby8TWy
xf9XKKWxZfFNFRlpasu6NfS6SLjIdjP8+S9ELMZpJASTGOvvkq/o7vl9EEvJE8Ky
prAVpDyIQX/qo1D9DNJlgaMQctgpOnCS++oP76fc46Y9RMe11j4XxLy/fbzuDCEP
TSmNOj7nucStaP82mxU9Mc/2y0lTdteR33To3cVhkMx5nCSLPTbYVnILZd5SFObO
D3jJxgxRhblT7VeT6P/D4iOU2Wsh+FtzP29ABPcO3EoWjyiHWeUALz3CLVcE3br7
plKbVhqKzRqd6I9eEl+fCGxPLOJC6MrOoKzZ8ymOxapgEzd8+eBLOxb62zdJsU4j
KYIZhosHqABgqIPN5hPm458Xqeg/NJbEuWDfZwkR3Jx25W7JhLA+c8xZ5TQtfg6H
ytkXY2CmKcFMIgEOqOc0GkNi9RCAIVYM9BcGHictGUYTFWM/kgrrwme9BDaIJDIX
C0QRiqag2/k/9ALIXHbf9t2udFHD4MlQDtW8d3jfhU7bXLlaUfdsBWENgbPEZhpu
/tE+RjS6xrn6+e2ZsUFpL4GhbX+kXqvuisa4ao/9MurziukalQcu/R5+X/KXTciG
6AUnCg46wdPk0tHdILqgUBvBll82Ajjh/+gglO9n5grFKsWfg4fcMbFkgYiLcKLa
lv80GOUJ4HJh7Vb6Ev/v75IrFYjzy/Jftdbxf+ulz+FEkhDRLaozHky9KGuoldF/
bkaw2FNj8aV8GMyUtKetzS6ZawYG/BAqaaT3vwDbvBBwJRgBI6X4zh1VKIfvG4b5
+h+ZGhKU7Tcw59u+aMNp/cFvylIqATnnG74egCB1rXLVwilAkDs39BQzDbgGaKuj
b35mVRcPC660f5D8VJ0ZSJan/Fhig0mX8cttxfnT1tRLFWySpgzeRDj8/p14nICl
StfGUJoVGFqbiMBOTsWym/YtNqNZbtaNdjuEIHARatgNYiZhK1x2H7vcnuUKlGUn
cR/2QW+WOog2EI88eB8GlKqLKZp8j/bkwP/hR3NYSfWxD39Ki4nBoHmjF9PrMmKq
7XbJjc8juN8L8ScD9gFJk8EOLhswGzNcjqyUh0nBtzkxe0rndMsLCPI2dG1cX/xP
S3Ua7rZBS+BrSduEEaaN1w06bMgxNUCAJj5OSbnjBFQgspy2Bt6TnxYeHCUoY9Vp
vgMzsLG1TbamqZk0svJhGRIOzdTwZa3nntKGJ9MoaTxO0OOtrTz2A5wxK+GX8TfM
a6t7dftoNdfAmpyh/QCtcz1z2HehTzHQqlcA+MTw1kgjiW2JwSOAnItWnH+X1TM/
2u1rbQ35aUzzICJlOebCDnGL/EFwRTqz2aXJPOoEmIau2x2NEb6595FsPTA0EPZT
lGTR6xznb8253idhuURKGWkMiw178BCdAd/7tVON6pNN7Taq+/us6I2t5kEq8odM
sl9t4tlVzZsDgjseBhKvXd4n5rMYEbPHctdHHEXrdYBvdvE3cxoUhaxziu9Iub5r
xfbKJxTKCWaJwSxNq1+L98IkaVNbKN0VzBwXmRPAoo/TfKDe/M+xOKvto6lx93lq
zCZQd+JoMESgqYCiICUlBtPywIzoaVkKW/CXGw7K4wgFrD33X6I5obZzfEC1AC4n
7hVj0F4sR4TDfJgDRP9lB47hDmQbTypTgw2j6pqYlA8hGOzxsetWEJvYda3CfG/i
26gPJMYTUFumPAwZirgmSdycKJYWXyZBdSSx/z093CNHYvkQ5+1bYT7J8Pdhaytk
mOcaIcvswOVSR8wJRQLs/Ha5XLy7yvnoiJKPbJOoymFfG/ZzBFB/CUqANZSMiBhE
lwFR1w0oHvsTFC3kA328lYIFx8s5ZdU1GBRM4+dX4uU9cBhJ7qtTqW4swKCVaDOW
HxrsoQ86WE0hmEbndNvhnSgYwN+x5yvdp0ytkSmooLJV6awOZlCfQAh0rFQA4WWa
z5HDiUjjnOPcC7LlTOloZKUzrL942QnLmUVli8BsMl6TeuZoCwaE6GYZ9tOtePAD
qYW3OkaJEsgB+MxJs1IqiBdKwywc5FvO4zfaAP/Q0Yz0mV3vuxbRTtOv6aXnL+mI
ugDR1LYxWqRkgw+ABqBLggu8VD+nrahFzkl1EtLZ4jJ7LbH3agKphgvfGaOQ4ImG
O6opM04cJeNWWd4ToKIS0HwAitB2fn49dX8vp5//254Bky4p3iYXz94+Ty+tAZEl
RaRqnUscNBGKgY3o/Nk301PJYHFZ1cn1t8GwoxQWqaLLL1jlMByCAGHEJlA0Of1g
2BEv2MUismF5gOHASHttLQ3MshSC8nZuXVsh/FyW0ldke6PY91zGsKJ/fuaftpwb
AIE3RWX7eTrUHOVHzZQSJJs88CIq3lOkorierYLDncfS/aEG+ndjwDHj8MYhCFX0
kYikBCjM87RtQJyUG2KeCCt+eYCcE0NUILvBPL8fSdRWZcn9Hx+DIx1HKp8wSXu+
h9f//ANf6hZBNQihtzADF+DKEOrwLhvXcs2lhRCFPt7I5Zt5s91fW/H2XTkYBnrQ
7y7pTzvCsbXfdAGUja2mX3RAKEGJCqF7/V0XWTsIeXgFZzz63kVwyXxazsxCNk0R
MZZfY1OPwXrd1uOyKNU6WmESPNkCsy7sqi/yKjhkpjhCR/BYsnI2DkRCKrv/BJut
VpT7zGP5zE/39AMYHGio6Lu9Qu1jb8x75ZLxIGj8k0b6HTKfqIv6QwxMIotuOoVw
d+keC9ZXfxygCr9E4JKwHPFcQNR5iSBXks/mAqnn2Uj1IrZL3ySUEuuDmjKri8CD
wZUld4IW9gdt2VMAyRkh8oM5kluQp+em40Q+FCIoJkPBV7aZlnjI7Rng3RQZ4c1E
MNArINBYK/02TuDAz70nt4gQ6uIZUEijDBKHnXqbuTlmkC8VqGg6BCxFTlNtoul4
7tY5NG7MGZDFC20b1haT5KJv/DUetsOEkXhlZsQ0BjDvCQtELZlcILGHPy1LX9dj
vpI4TcFDvBjuVqVV4+mNaDyDbj+p3EZF2fLHfGa52kzhh4rqwxzPvtmFyI8Fn2aQ
+/dv0N/CIOJNTt7nLejul9Q5tWGzxBq398GLV6u/6B7G1+OSnK54xBNI66q/rzVo
xsn4+51O594ciVoTigFMElM/GD/F2MdHmDQIym9pgMcv/ksLM1TZuHXJvNwa1AWo
s2AmAVWfSAaailyMIJhQ0x4CDLnkb2016nHUHi1Q1gENicuurY+gShLc4lF9dcBe
lK1ymI0j1im/AUHCB2Yj6X09gNTqgxsm/CuFrKIROQUycFxxkevnrnEpE+nccGbT
HCsnAMq+RN5T5QkOBtybBCdwlsBAb+sEYgU35l6WdcXHbp7u47/iYBl1feInFlac
LJhDgifx1xB0wYmpJe/d51nhz8UMPxrU5Kdkmv6J6ckdgNxAQnYT1B0VOMWudcE5
DMPSsqpWna4xPIlum7tegaUnLZnj7teypKEboTGZZbwrxraCUsT6uBqYk8digVPk
fzsP9pB8gdreeYnqeXSc7CRxVKUT4XC5JHhmiUYeH2KFCvMWMCKy8+vyAoioUay3
0H1M9eSUXxfjDSjhXKUaHT1JROXn85uten4qUgxzKNpmfEBjbJJLD4t5aLYvbLPu
vKg4Xl15YX3fJLGmJG0fuAypuol6xgVoJsjPxkh/VuLuFc0+N8B1dUf2WTaJSiy6
w+8B7sxdewqqL4MmQ+aQ8d3NYovUTtQpltkV5fQox6rFmpFPyyrryY0DdwcEzf1o
E4uIbYi8D+AVei+TlPSQdaHQ2e+n0S/s1Slljre+/uAuJmQg1iEJN9CA0+pJqnVF
56RMJMd3dcLYylfpsuaxBgWtHSEOjN1P4NYlZjNqA+USHM3kGudC7f5wN+GAIKWX
Bpat8oNKPnvoj5630UDzlhkmmCWDVXnYLWCHMYH+H07S/ikx2Zqu7Xqy5HAR9Cl8
jmN8bW8gT5bb7J/nH1NXVJv6zI8LXNVkx15tRKLo8ejvwuC5f4lF125P+9mED+h+
LgWJryACpRvyjFSJSbWn1BG3cQGx+c/vI8cOb9Dr2Kyw1QvkOi+btPOwmt872oEf
TCeR0HhuKCs8BdOxKieB5Z3Pm2T/DcjraIKYfMVfg8f6rpIu82h3IqEDBOyr6SXX
b3SJFXUXYDJAboCXv1c3jQqn5zJXL82bUjrd1c7hcIqQXHUnIkZyr2b2CZkdcDCy
dPlSqR2mJVwTqoUYIWMSLM6wW8gBdtcnSl38gWYKBFLIqdQqTzhIoPkDrZetM7Vh
PCwWzoDRY+KUGGQuHFGPxi+i9b34BHC9RRRNbfZz3yjIu10pAIUfRRTxI/MDR+2i
WOtVxjZPb+wk3fahzmu/3KT/CEabn0mHZzKo5+7236Klq3hVaSkYqEcyizKiRZzG
FS6JUrXHporjGIZQehk7tpZNCJ1DTPKE8uNowgQoUdvwGhvPwtqpK/PyMRj755Ld
EmOjei6NCN4AxM7fjlbNKCYhsl9SD1mtk1D0rcFch4rB1W+VhZeCuT2g1bb5q376
E17DbMrcxDuchNrurqvu2XIRdIlOzOp3vA5ClWz2V/166Qg/27XxUfCLTzjhJ3+t
1psuouGF0xnb0NIpLv8R3P2V8LWz0HNxpUDHBII9YGOrZFZJipAnzUbTFkFat2aZ
Cdd2WUyrywB4XjrgrCmyFBJqDUlieofFesqLeEuWIVE=
`pragma protect end_protected
