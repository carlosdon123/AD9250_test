// tx_jesd204b.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module tx_jesd204b (
		output wire [4:0]  csr_cf,                     //                    csr_cf.export
		output wire [1:0]  csr_cs,                     //                    csr_cs.export
		output wire [7:0]  csr_f,                      //                     csr_f.export
		output wire        csr_hd,                     //                    csr_hd.export
		output wire [4:0]  csr_k,                      //                     csr_k.export
		output wire [4:0]  csr_l,                      //                     csr_l.export
		output wire [1:0]  csr_lane_powerdown,         //        csr_lane_powerdown.export
		output wire [7:0]  csr_m,                      //                     csr_m.export
		output wire [4:0]  csr_n,                      //                     csr_n.export
		output wire [4:0]  csr_np,                     //                    csr_np.export
		output wire [4:0]  csr_s,                      //                     csr_s.export
		output wire [3:0]  csr_tx_testmode,            //           csr_tx_testmode.export
		output wire [31:0] csr_tx_testpattern_a,       //      csr_tx_testpattern_a.export
		output wire [31:0] csr_tx_testpattern_b,       //      csr_tx_testpattern_b.export
		output wire [31:0] csr_tx_testpattern_c,       //      csr_tx_testpattern_c.export
		output wire [31:0] csr_tx_testpattern_d,       //      csr_tx_testpattern_d.export
		output wire        dev_sync_n,                 //                dev_sync_n.export
		input  wire        jesd204_tx_avs_chipselect,  //            jesd204_tx_avs.chipselect
		input  wire [7:0]  jesd204_tx_avs_address,     //                          .address
		input  wire        jesd204_tx_avs_read,        //                          .read
		output wire [31:0] jesd204_tx_avs_readdata,    //                          .readdata
		output wire        jesd204_tx_avs_waitrequest, //                          .waitrequest
		input  wire        jesd204_tx_avs_write,       //                          .write
		input  wire [31:0] jesd204_tx_avs_writedata,   //                          .writedata
		input  wire        jesd204_tx_avs_clk,         //        jesd204_tx_avs_clk.clk
		input  wire        jesd204_tx_avs_rst_n,       //      jesd204_tx_avs_rst_n.reset_n
		output wire [63:0] jesd204_tx_dlb_data,        //       jesd204_tx_dlb_data.export
		output wire [7:0]  jesd204_tx_dlb_kchar_data,  // jesd204_tx_dlb_kchar_data.export
		input  wire        jesd204_tx_frame_error,     //    jesd204_tx_frame_error.export
		output wire        jesd204_tx_frame_ready,     //    jesd204_tx_frame_ready.export
		output wire        jesd204_tx_int,             //            jesd204_tx_int.irq
		input  wire [63:0] jesd204_tx_link_data,       //           jesd204_tx_link.data
		input  wire        jesd204_tx_link_valid,      //                          .valid
		output wire        jesd204_tx_link_ready,      //                          .ready
		input  wire        mdev_sync_n,                //               mdev_sync_n.export
		input  wire [1:0]  pll_locked,                 //                pll_locked.pll_locked
		input  wire        sync_n,                     //                    sync_n.export
		input  wire        sysref,                     //                    sysref.export
		input  wire [1:0]  tx_analogreset,             //            tx_analogreset.tx_analogreset
		input  wire [5:0]  tx_bonding_clocks_ch0,      //     tx_bonding_clocks_ch0.clk
		input  wire [5:0]  tx_bonding_clocks_ch1,      //     tx_bonding_clocks_ch1.clk
		output wire [1:0]  tx_cal_busy,                //               tx_cal_busy.tx_cal_busy
		input  wire [1:0]  tx_digitalreset,            //           tx_digitalreset.tx_digitalreset
		output wire [1:0]  tx_serial_data,             //            tx_serial_data.tx_serial_data
		input  wire        txlink_clk,                 //                txlink_clk.clk
		input  wire        txlink_rst_n_reset_n,       //              txlink_rst_n.reset_n
		output wire [1:0]  txphy_clk                   //                 txphy_clk.export
	);

	tx_jesd204b_altera_jesd204_161_py6ow4q #(
		.DEVICE_FAMILY            ("Arria 10"),
		.SUBCLASSV                (1),
		.PCS_CONFIG               ("JESD_PCS_CFG1"),
		.L                        (2),
		.M                        (2),
		.F                        (2),
		.N                        (14),
		.N_PRIME                  (16),
		.S                        (1),
		.K                        (16),
		.SCR                      (1),
		.CS                       (0),
		.CF                       (0),
		.HD                       (0),
		.ECC_EN                   (0),
		.DLB_TEST                 (0),
		.PHADJ                    (0),
		.ADJCNT                   (0),
		.ADJDIR                   (0),
		.OPTIMIZE                 (0),
		.DID                      (0),
		.BID                      (0),
		.LID0                     (0),
		.FCHK0                    (49),
		.LID1                     (1),
		.FCHK1                    (50),
		.LID2                     (2),
		.FCHK2                    (0),
		.LID3                     (3),
		.FCHK3                    (0),
		.LID4                     (4),
		.FCHK4                    (0),
		.LID5                     (5),
		.FCHK5                    (0),
		.LID6                     (6),
		.FCHK6                    (0),
		.LID7                     (7),
		.FCHK7                    (0),
		.JESDV                    (1),
		.PMA_WIDTH                (32),
		.SER_SIZE                 (4),
		.FK                       (32),
		.RES1                     (0),
		.RES2                     (0),
		.BIT_REVERSAL             (0),
		.BYTE_REVERSAL            (0),
		.ALIGNMENT_PATTERN        (658812),
		.PULSE_WIDTH              (2),
		.LS_FIFO_DEPTH            (32),
		.LS_FIFO_WIDTHU           (5),
		.UNUSED_TX_PARALLEL_WIDTH (92),
		.UNUSED_RX_PARALLEL_WIDTH (72),
		.XCVR_PLL_LOCKED_WIDTH    (2),
		.RECONFIG_ADDRESS_WIDTH   (11)
	) jesd204_0 (
		.txlink_clk                 (txlink_clk),                 //                txlink_clk.clk
		.txlink_rst_n_reset_n       (txlink_rst_n_reset_n),       //              txlink_rst_n.reset_n
		.jesd204_tx_avs_clk         (jesd204_tx_avs_clk),         //        jesd204_tx_avs_clk.clk
		.jesd204_tx_avs_rst_n       (jesd204_tx_avs_rst_n),       //      jesd204_tx_avs_rst_n.reset_n
		.jesd204_tx_avs_chipselect  (jesd204_tx_avs_chipselect),  //            jesd204_tx_avs.chipselect
		.jesd204_tx_avs_address     (jesd204_tx_avs_address),     //                          .address
		.jesd204_tx_avs_read        (jesd204_tx_avs_read),        //                          .read
		.jesd204_tx_avs_readdata    (jesd204_tx_avs_readdata),    //                          .readdata
		.jesd204_tx_avs_waitrequest (jesd204_tx_avs_waitrequest), //                          .waitrequest
		.jesd204_tx_avs_write       (jesd204_tx_avs_write),       //                          .write
		.jesd204_tx_avs_writedata   (jesd204_tx_avs_writedata),   //                          .writedata
		.jesd204_tx_link_data       (jesd204_tx_link_data),       //           jesd204_tx_link.data
		.jesd204_tx_link_valid      (jesd204_tx_link_valid),      //                          .valid
		.jesd204_tx_link_ready      (jesd204_tx_link_ready),      //                          .ready
		.jesd204_tx_int             (jesd204_tx_int),             //            jesd204_tx_int.irq
		.sysref                     (sysref),                     //                    sysref.export
		.sync_n                     (sync_n),                     //                    sync_n.export
		.dev_sync_n                 (dev_sync_n),                 //                dev_sync_n.export
		.mdev_sync_n                (mdev_sync_n),                //               mdev_sync_n.export
		.jesd204_tx_frame_ready     (jesd204_tx_frame_ready),     //    jesd204_tx_frame_ready.export
		.csr_l                      (csr_l),                      //                     csr_l.export
		.csr_f                      (csr_f),                      //                     csr_f.export
		.csr_k                      (csr_k),                      //                     csr_k.export
		.csr_m                      (csr_m),                      //                     csr_m.export
		.csr_cs                     (csr_cs),                     //                    csr_cs.export
		.csr_n                      (csr_n),                      //                     csr_n.export
		.csr_np                     (csr_np),                     //                    csr_np.export
		.csr_s                      (csr_s),                      //                     csr_s.export
		.csr_hd                     (csr_hd),                     //                    csr_hd.export
		.csr_cf                     (csr_cf),                     //                    csr_cf.export
		.csr_lane_powerdown         (csr_lane_powerdown),         //        csr_lane_powerdown.export
		.csr_tx_testmode            (csr_tx_testmode),            //           csr_tx_testmode.export
		.csr_tx_testpattern_a       (csr_tx_testpattern_a),       //      csr_tx_testpattern_a.export
		.csr_tx_testpattern_b       (csr_tx_testpattern_b),       //      csr_tx_testpattern_b.export
		.csr_tx_testpattern_c       (csr_tx_testpattern_c),       //      csr_tx_testpattern_c.export
		.csr_tx_testpattern_d       (csr_tx_testpattern_d),       //      csr_tx_testpattern_d.export
		.jesd204_tx_frame_error     (jesd204_tx_frame_error),     //    jesd204_tx_frame_error.export
		.jesd204_tx_dlb_data        (jesd204_tx_dlb_data),        //       jesd204_tx_dlb_data.export
		.jesd204_tx_dlb_kchar_data  (jesd204_tx_dlb_kchar_data),  // jesd204_tx_dlb_kchar_data.export
		.pll_locked                 (pll_locked),                 //                pll_locked.pll_locked
		.txphy_clk                  (txphy_clk),                  //                 txphy_clk.export
		.tx_serial_data             (tx_serial_data),             //            tx_serial_data.tx_serial_data
		.tx_analogreset             (tx_analogreset),             //            tx_analogreset.tx_analogreset
		.tx_digitalreset            (tx_digitalreset),            //           tx_digitalreset.tx_digitalreset
		.tx_cal_busy                (tx_cal_busy),                //               tx_cal_busy.tx_cal_busy
		.tx_bonding_clocks_ch0      (tx_bonding_clocks_ch0),      //     tx_bonding_clocks_ch0.clk
		.tx_bonding_clocks_ch1      (tx_bonding_clocks_ch1)       //     tx_bonding_clocks_ch1.clk
	);

endmodule
