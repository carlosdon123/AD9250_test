// rom_port.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module rom_port (
		input  wire [5:0]  address, //  rom_input.address
		input  wire        clock,   //           .clk
		input  wire        clken,   //           .clken
		output wire [23:0] q        // rom_output.dataout
	);

	rom_port_rom_1port_161_iitz24a rom_1port_0 (
		.address (address), //  rom_input.address
		.clock   (clock),   //           .clk
		.clken   (clken),   //           .clken
		.q       (q)        // rom_output.dataout
	);

endmodule
