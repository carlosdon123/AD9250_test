// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:20 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E9RSLK6jBR8NZJobF7oKmFoQRO/D8ZJn5Nk3rV4hT2ujZrewRBwCbJD24FxAOGNj
zlS8RQ2n6zPhXZeOOPzouT8Qu8GoBLAFMVHFlvjr9Hh90zEIGhSmUgqy1C346kvH
/LrKp7p1uDePQX8ZUslgSCKRZvQyQrcE0Hp7mUGQWM4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10768)
wtoZ2D2YPaeZLUdoLzuLGdlRGj740RdNoNQLFcZJpKu0uFaqX95oTOC8da4CAGLR
Ef+vHuGAFGofRwi6TqCKPXUOUaO2oEUEvOj4HkIaq+Bv559caovzBuSkgzP5p9fX
q7+E5eWPhlaPOqD+i9OxqgXwn3Fz6GPIDnMOUCyzQXgb9wnCxdTFbww+tlg/hLrU
gkJ2lfIt8qQQMNLt+IPydhLmYgLqBCwn0OlI1/Vqch/GkTw/qKCk1MnCE7z4sNum
jWZDTGDm0bXuhOnOoJHa4TmnnyDeMF+LBJtAi9l3fxvr102wO6N7KzCN9TEEjqLS
1MZioUrjAy6zlApXmYAkCjFR7/FYJV5S/2iivV29NuHPWOZ0dGuRCceXawBqEMuR
GGpvkGQjd2iwry6BSuUr2HXBhof2QW8TnVl8Huw0wehPdSpsl3CJBRGML/agEYee
EGfERQtqUjeyi5+s2dWiai6KfwX7gl//WQtCEx8R4Vsa1cdA3hgyPrNqxmNSdJCW
3xjvepC+gw967tRdb1GCGzW7zF82AHTz9MviyhDvSi7G8ogoz3EQFfhJf6pZOSlV
JJcPDHtGESLXl+mngQhRGabGbbd5ZDDYIyOwpx6qS43+ILhGvld/tGOvYOrFlsq7
9s8XqL/3OC0kijXrt1l7bR5uj3CpgO9qsl2Xt79DRgY6V9XM/C5SJRCYJGT83k3C
S0tqqjfBan2PvzSSC3KJy/rUqNHzyf+GzHUYGVfYC/nlVpw3mvS71dG4fKYVwCLx
XRgwnfnJnpeRAcyJkGUeMr8qTZxTbfFDaG/4QZSirSfSxVh1UKY/KxW0WZCTR3DG
BOzR7pWaWDjv84znLUryplpu+toBBAWbchBOCZHJR+yENcdeyRSPQJB2Cbk+2Orb
myXhLYZUAoAGZ6wsIWt8AnPMGe5jPQmPkQkUV0sgphcfhDgf2mfUjvapnM/BepKP
ZK6ycNpFrhM5OpoC9mN15UY3nmBIGC0IpaoEyI2NoCu2Pfc4rZ8WiBAw9eIZtyNA
Le/RODmFRVcgFfsje2UKViroqx0J5cXLOuLJveKe92isEuAdqrk+yzWbk3AYs2t4
DNrDm6CZ9xGVUh89kcjpaSeje2cHYlwxHYQWyuJsvXeIdU0DD9eZyc3U5YGg8w6K
3R7E9IcjqyCIklBi52HdkOLoOoDDJLuu6IixF1+X6fNjirknU4aAmhckza2VNz8z
qxcwPnZOUM4qO6wHBOsYIGfGC9vcyH7LxDlfRYqZFWuTz9UEENRjRwQhE+ht1EnR
6A2CpBjQQiebUe3qrg0NkvUoMmgDQChi1VcUmqo8WvgkIBF/RR2ACTyIdicSWYhW
72GTDEBLcCCdKfApytUvRYmYFGOA4Kk7uNSTWaw1FgQdLuDOiAsUxoTi0A+2aGrN
Dlwz14nh/Hjmfl6O+k0a/WP2gnCOM0Id/hnPftxoILr/qV7R/JNJuy9wY+99RAgb
cX0wuSpTT4tqz8sKqgUv8uAsM6qHl2gawGG18lEj3jmnVI22dpywsMEG2plnU+Pe
2P6MOG1pmPVM9PcYqwRyyx7Hm+G6Fuvi2WKL9Gyb0UCu0QARUuMw0OrmNoY6XAtG
N2znmjWZlQVeb8qvqi757WEjJpHwCJ0C3rO2o6OXrpP5Q6+3S5/Qs4FrA4xoRiH7
idi+eIbVOHKx9MdnPyH/K3UB762YdiMOpx+KQ65ThViwzOL3YmjevbQsrdhUfefd
+aUPyXlBMtP+0j7I1nciEzTJfrmdGRVvOo29VUMdiaLWxaHvcswe+sh+FyV+NJ2n
lWHCMIz09Bttr3Q5vd104LnnivMa9KfPwIkoYj7REZsXQaTd0GoGekGeHUnVSGRn
DBoJ+i1o8rg+x24fitdWjjVLhEqFPP+WNjPqfG5TGQ6t0QNytzz0TxGhG1gGx5wn
zuSB/IqJ7L4eHeoaXQd0/25FWCCGgPTKfbE6yHZSU2yMDI9+XSFibvyOwQLL7Yzj
DcFEq2bUWAUb6CqZaHRKV0dnsVid+qntR3BSFutR6Y+MUPNnsx0YDo6IDXdF/GFb
yckIkQCYPalRRlOw2CpUL9BM3Ulpi0kTdTeAJJnySWcwaANDgxw7raQnh0dWdJe4
CMaQDpOqE1wKboQjknt7VCiriPBow5kV9+GGgvrJRhtWKS6G5VtxhoJ/+5iztXRD
jbTRX5PKK9QV+YfI6Uib39QaLI6YubWpc8K/oOhbCCfd49QQQ/iC28S7sk2HQOp7
wFnXO/1WuAG1C8Mw7esGz4WMovFn24cTMdoxe1Rf6pIZ5Q6sSLykjEFg2sPM7DNK
uXpX5MrV8IusosMqw6ZvwTpv90hrx74p9VxbRqe4Z15aYv7Gy9DqOQNDHOG7BLOL
GpQ14R9Jb2/CMOwB5b+POkSbKD0XVuJJjouaoWLMEVOrFmepX9HfkWheUA6teEIM
ugtaJEwj+UARbUxtKWakeeSzuVsePbh+HEKvKExNGIM8WbiBoA4Qkk6prOE881CA
6YtS8TRCsZDxUTIAbMqQkXH2IpBoGSdoFT2+8KvX1yoSJd14OBMpZGuiGOTt73C3
YoLkxVUjUe8wE/PbnbZLKZJt+S1MrFFPXBZzFGod1fDaiSRr9HLnoy1mKJTYSjtU
d24prnsRKHK/umdKRpBo4hyFAsz40i8mHYVkcvTl4AimY1XdQyJSg80k+TW4eWjX
omuNjtIUOtSSWEjkLPlszvSOTKST/lQVI+WJ+x0941vwxnQFiR0ZjmdR0enTd0U4
e3rpPmt+QmQAtyVxnZQCqhBmXfnnLacPI2x/+UgVT7bRWZZjKTf/z0VwnAALk5D9
1LS1eIIeNnu3gyE/BdxtuinA31hgzZ+FRD9y/jjiYTtvHV787x6AWIDPR8VthSQK
tm7TnTpKD7adLsFNdFV90aCKDfSRBs/ufowUCkNJ66wCNg9HEYsv0M1Ue0ZMj/R1
0U7+O6MkHVmz2sNEFKKFzOe8y42sk9wxhHmSDt55Yqubi6+5E4lr380wca7TtR1i
n2onjRHnq4EupBT4P2SYvwX3+2c0FhGNoXrgKVxgIqgXfFfgZPWPEJ/jbu0FAGFm
67+h8TwdawTO75CyTMbijmZWAGjhBfPPrGQxIe7PE+pC+/EGZar/bLTuDGQexxz1
jGpG9wgZxdDM0CxGTYs6Xk06IpNWwhDeYGae7jjTyVy94986mxcqqDY58zjRjwOG
sVcE25w78x7+K/34wxUt4ZwM7SanHm6MX0MkCoxs+9c1CHmbCuFgH6UI5N0qDVdt
Ui2bY3brV8BlrzbM+WuC1TqWzy22XrE2MDHvjttVk+Y6oHADjfDBPvYdGOGA1iGL
TbGiQ+uBBUkfHbT5M1ld0CV0KzrBDdmRwbUK18k2jHiIIPR4Xhz8+Ya2530AtJtB
cGUUn0yGzIotNTXNrGw7VW1wTKRmhiNZBLpEY/rpei3t28cUoAkMtu9uKJmjosQL
8h7w7yFY8dMS75bUorDHQElIbgj2K/j4FNST/XdPcypiVxeu9cbjo1+PEuZKiAVh
m4fQDRMb5lUBNFB29EdenfdrKep4buT4k8ID3fnCtmj51dhoaxqbqylixOMevxFq
ghlDGQx4wq54IMQqJ7CHMMRTx9iVg3Ng58BBYXtuEgynZH9TCOY0C9NZ4CpB3ghQ
nv45jufTZ3Mo5dUFxRvSo9/GzE6JLXVPM1N+6Oc0o/KTYd/BQXLWKmzlZTeUQeOo
wC6mPl/phko5QWD5Gn1ZJPtgyA7Ps3ZIZ4wWadNQKYbMMmF8U7RCzENLiQi0w5rL
96WZ4q7whNvbeevMV8DurkbPqESWlHq92yupPqW8bM9MhZhJjoXGwEksmWxUlFV/
lPb7Y+5OZtR/DYug02y4kdmQmBtDPqbjHDhrA1e0cW0GqalwQlUvdinwtoLGhXBu
OGuG25v86VqJE9vzb5Yo/Kk9IjX/efEo8t6DymX5I1EyaA+MS4FMX7D4w1f6ohkN
XG/ZPF88t5Uq1ElaX2j779MRrpwT8FGLcDwvJuKmJ0kjyAwj0BkQ7GQRTPdSM0wr
kwGNfXK9mLpYl7P3f9gjbMb48uX1KOEKo24LcORtdLWuBbrpnyBISkhx4ZGaWcuM
mXYb8c7F4HmGoPYAI14P4Ov9iBoPwY97WVVa7O+jy4RKpyvLs4E3hUKJve9fLxev
q5W9V/f2XgfS+dQBXQYtu1GtlOZ3KMeiS/cF5/vtBkiW7CQlyPTsxb13uGNbEYwt
5M6sH4I185sM+CCmiF4boDDlH++DFgQSGwEc/cm865GeMuwJpi8UckBbtUNJnF87
ISBdsuOoHEaix81Mll4hVi5jo5vypmlvxLllUs8v81ZM3HJNcXgXuvgzudj/T5SP
i3Q+my9i47Z2Nskjh1mxm6appabL59mVujJLXSDyFRQWU/2iu7c2SqF6FD+Y8yRK
A02gGf+XtNni1fvTC9kyWl5qy/aybzTKUCPBMJhJVR7TOOxnjO3nGYyravkNs6wC
MjgkBwH+t2/0tG17464Z2Brbbhw7lNF0VIXTCxRjkIU5pIcHto6Wnu/U1kQ2m7Ih
fAgxXKSMJ5mmaYVD6VVfqnfuDncVjLapdYKqW+bd41IMt6XEq80BAZbsksdGIMo5
qikYXQIboPUzwh7NMkbV8U9o1+exOOlveNCwizzg2ifCY3hmFYYoCrLLXZeAzDUw
I097D4x2n4+VjVKSj8DkBI6Jzaqgx2vLG6HK552NCB8t/sEghhFTA6cR7QxHhTKX
KTwwF0kg6RDLyZ0Sr7FpUKpTCXJ2Jtd70PqbPuY9yMdT/AMZf0SWVB4xm31VOXcS
arES6WVNnr64t25A8VpMgzTNeWoPrRjK9t8L9HFbPLe/24NNI8zMJf8Nd/E/sP6c
Lz081tNh3kuKyJT8lg7zX0eDMeu7olI7GyodLyDXec2/W/wY7/hc8WUDexWf4+jp
HBtDxxfyeeCEShLIdu2siiL24ukFu6nxfZyiow6OtDkArAu3Ch7Os7W4s84yeN0E
LTB2cpfRilPR/DlkNMfPxEeolK5GQSmG3yxMXSKXDjKYU9X5+eUEbH3UG15j/OJG
QS17vPTzOB3N4Nejg1k+g/x8OB/OfLBC6Xwo813Vm6vvtJj0tGZ6QItft9TUHnuo
12O0JXysr4cbQhktKyQbpCVf/lbRW/gGMO56XZmZNRI0cWGM0L7EJSqBOa9iTGXS
h0D4YMbZ8MMmUCQlg/oLSEglQO+kRr5luuNY1UdanoUtOse8R1uRgFLd0ldLXypI
wXP9LySZooIGFyDzU9Zl4XMturSpL2b32AsaTwXa3MlOokAKk/qnDPzTdSI9WYqI
OtOr0i7X7eBJKtmd9/M9zEp5GfWyr7EUBA8XyuPDx6hypgVLi5zYVUCXXrBGq09+
8f2hyDMbAWRS7CFzrf1+hXyy57AQCwhXw2JLWa2TqUj4Toa/DjP4x+IioqYr4LJA
RizUvwXQRCdyoCzzb6EnXfDmYSaoJHwuKcUTyIdae3LellFgjwM/8njN1Kl/UYHk
j9ou+9+RVq5hlDpMcBZYtndGuLKZ9pCO8EGfrID+j0YyeAqtZrWzCgCbSW1l7vD4
7QZWSaH1tw++HTGMJBRe4iRUTb4gAjrYWLtG0Muv3OHWAMGBWWPs2LIG8W3trnsu
lu+Jads7mnzxSabc3BXeI61tT9nE+h/3QdBUV8X4Xug9zh5sM35TQUYROUk0mP+I
0J9RqgOSBlBJQN8Bw8fR1MoflPm4thkITCJWG8fKE3k90oQ9/ROX3v5tWzWfo7Kq
bXWW2puxMItFFSfjyURAynCcaHDcfE7wpLJ7riVejPHquXkuVocqZhRi49X4qkKb
mcry0nxVC1O/JZQ76YAv/H/BlpTI2WrLMLF2e2+3DUzbHY5i7rAzc3a4K1U1s+S2
jAnoeYZNQORGEx9QTil5WbOcxb0YMJRFHbZTqmQjKVa7V4g+lK2EfsDx8DuN5fmG
i2O+WByTEE3b0AnKytwqCtNi3UTPAV8ikC0qydo5225zTitqSin/UBK719fIXyv1
hQnWFVuf/iVAAaQjhHHaU0m3fVs5XKGpiUCh1laHE09VyrzSbJ5gYlDJwe1rrNEL
Xs0/iC5cW5fNioBvt6UCBeZ1p5WW+zMmIDYpo2L5gBsfFwAXtYGHvjWcMH26EdwH
qmbg5jCR5tl56+ZodDAyPdctXTFoEMDJvD1117xEGsXdRl9LXopL3UPbgniFp9Nx
+StMCcPBQx+E7VfwX/WcOnmeCSrXX5nW0H2WNfnVbwJSG5c6dHQAB3YAT0Ol0arV
5w5HB6pyjKx1TNrkN5kyRfCj81ze0Db7HdB8cmM7iKn6CfhVvTPHMjK0eETiYQb2
j7A2U0qAx9tzPjlUa95VkWTt3qnt3BMAgMYzUzHAHg1KGCm2KkE3Z+AAB3D1Kp+D
FTIZY7CYjXO6Jo1UnTXRUoROxjvcDFxdf7tVB5ixWILGHqaQ+pZwG0nG2d7xPznk
WqkvpCjlf5FpMpH7MEsPy8kZ+4pC5662S7TALnzsLX6PpkeoG1MTen2lIGIiS6SX
04yJvDXuruxTWiisT63CirWQQYujx8lWtaLiQkNoKpPsXS2GZR/XUfEVm/9OyNMG
xqHHTHv9TKDeJEDfXIWw0e+oLdjCNJvE7TTSG0vdOfnyO+G/2+03+zUm72Klljx/
hYdxT3nHrMfb9bW7o37ST3LLgqH5MFTtD9Uljf9NBumCjZD7qn+myBByLc1dDl0t
UrHrFksLsoEOJwl1OXCYO3iY9mI4OIJxhuYQ/4R8bhFIqGCkktLyMCDyQnytBzdI
mE3yEnCE6ueki9a4RuAbAZ04ZoUvz32JHhaRM7KH5It79jQSfxCZz5LpIfJcle9B
oT3h+udrERzXJFrBUJe1Fl8RDhK3tFA4GIFBp2YBISayOLW4tz04mPwZJskDrEUM
Cz4dssRBfsRAWZ+oBAiMn4KcxnVHJbHoOgN04BbyO+S6pQwK3deOdyyClcy5J+fw
fiigtYe/CMFG7354imLkhukwxZa+bgvVxrfxGKneeJq2kXr63oSqMjK4Yu7aqUiI
mW97xjC8OUMt9Fk5SNPVuJfXIVtcf84terI13aDz9KnCE5F19qyznv9ziSw4t+Zs
Nj8ED528UXsbTL9lyX+j5skfaCFWT7rZJYTnN5bjqRGhHibcsH0gvxyHIC0wUU8I
QzzKz8SMotWMlbXprUFS6FYvIZ8tNrSOh5V11JojmG5NPGIa+whRRvY5ptF14dbJ
5jrvIDGAXJApr2umaqtL/h4euWhDxHlQB0kKF+G4e4bOlwL8W1kYs7AMwBxjr5df
UdIgmk5hhvvOzCq6lCx5pACxStbjHSsFLiwSIXN0I6Yq5sMY5rDIFQLt+bFB/CrT
l4O1zvfrUdvWrlq30AnP/zCK8TANxKmttR34hR8xpe4F+8E52PraXj/eKo3ERdUx
/0/MWjqNLg1AoH+lPZb7Reo0pI35KKrkP1eBmPE+5LO5Uiju3t4B9oe3/KMDlPth
rrxZp+N+dsUqAbw5qXO3e4Rp+ZEyZREiN/R6oDFVhZzM1en0xvzcb2JBr7nJwN5w
zZ5Nwvud1vBCEsCDZDRD9cFkaru7GHVG48ANh4hdnE37m8yW2HSy3rD/1h2DLio9
CkwS2SXIhMkivHMbBU5MU7cbvXzmASzNxfG0taqpkj2rWdL7amKsDzGdiZL+SKcy
pmIBSJmYOSCR1X4mwvjOO1id8Kz577i5QS5npEJX15ZNz/Tin3ySIF7XkqILku0R
MvLOuTp21SXgk0SJOv0cYmIoTB9J+IxUBJFEX2H/4Fhbu7HiKlCh411KGnNoaL4E
LTnV5WSBHWUI3Yy2emCkL6EbeiRdz+Y8erD2cXQES4rjjYghG3noZwdIns5V78e0
blne39akeAUJZ8Ls+qlJAPhUmDlj1R8TLIo7/ru+F9Fdqft8C0j8ctLXFLttzx9t
g9Wh1QjNi5FTl4H6Wru3VFyEnuu61JXHtO0TNkirPquJk0UxxUO1H/vhdYkI2jJe
883DJTxFNjrbo1Y/SAiErIThNYagW8L6YTdwX5cY8EOBgV9oeM+Ua5TIlKjVyUJf
u0fkyKJCy+Ckiz1L8jQjq+xbIZBnY0qBNlL+8JxHn07SaLefIa/3wCcfqS/kKBNu
i+uxV4ns1w8iJvv8McvAApS0L0FMgcqWjHrzqSxjuNygVBFr08eZ4wEtOwS18OK8
YYJ/Ub/cZHYzMalfYeFHuAR5/BY7gpXsC7DTQU4y4oWCfVzNwip4a9giinSQ7cYR
zjQQyyH1Mlhc82tcX1QsvcriTPYu8+NoOaB6/Kq/gwXEcY3nfm1gr3Zpt2DOMi4W
1BoPeWiwxRff9XxE/uPWHGI+U+mE+QV4a2b948CyUJMG7h75IUxZUW5Hk5/2ZPkh
BDQb4ljfZRa9zMopcUJkw3uAbl4GkJtYSi3vtHdjufDixtkY4enoyOqupX1LrzM/
9g0P+HUnRTIF3Rcc08PPJT0gylFxKxEyXnGkDlA/AXz57/RkowGMMInL6fctYpHe
orQOsLVUVhMjr44ytagc89QN0OvxKfRpn5Gc0I3nNfIwzQbJa15I/ej07K9hwdo2
nxvb/G0LX5UjTgXc0jea9CSGmAksPtfTl3ktkR6YA+qJNHF9igfj7ZUMXmfutyyf
SqI5Q0PtlAHg8HaBmiL0DDEPnVEChRyxPkZnkX25Kj3Fha3AYZ3SHzu+a395xupo
m/1oJpLb0Jg05pU37Q8o0AtU3muAQe0N6lpoo8FRSc1a1ePJMjP7GQcIJceL6U6Y
62yJdOSKX79mVYjwUMckpSS8rtVK8t9PanKMnT1VoRI9my2IkP/H1NysKxB32vv3
SDJ61pyxtBIt/YoIDT3+1gu+AqdBbzkb0LOLacer202nmoqWq/m5Nfu0hayl/Ypo
qw8rE487jNgyGBM3oP9sm9ePLSbuLaXQgDBQ+O/VVtKmed+ePVu3StB1J9UXiQIQ
O5ar3WVe+3Pus6qN++7x+qZw5OXrXaUen4iDUSIqIQvlK9zJbhfz6kDJgC1dS5ST
ArfrLq16iID9FmROgfYgUwhJG79EXtCNDv6uCJMWrGjUsR31Pi4IZX8ID6ZCko38
LQ0T8889FocWUjmW+sS/FYLXTVYfx8CWhDo/Y5cTWKyiEJV8QS9XZ1G1ToDw49nu
vjsQc1FYsSsoyN5NTV7uQB3I8yaN3qPeEkhq6kIYl9UNfsI56Ew6QK8KwHn1ZLZ+
RcY+fzpeLz5TYMMI1wnfGYvbEeg70ygF+vNQgxsnS4wgb3UWCEAFEK30TqwXxn1G
yaZ/IAMpSqH9mOV9oJvVWIwPzxWDOz7K7cnhWZ62gsTxjWO1cM3pF0nlD7AdYpuj
mE4Kz/qyw6GLQX5Yfi5LQH5r7yjvG1XWP5Rsp16Nxext1BstgZ+24Ok9VV83MUDw
ulPCngDMSlUhVg1xe44/ldsmn5cdlakv+a30FHzdq5u2dRuS6jxT94rpoZSmaMvx
U409DPXg1kO5X/rtSLCJmKE0xk2eu7kXrJk6GusIM/s/m7RWYSszvNLmRtT7h6oB
zD8ygsIUeMLuxLchwmK+JezsAKsMhPUc28IeNAs9akEyq7bToHAgB5S6DXg9029y
PX5A9k1bFAX2ZMytWXl4Xl1zlikoSYXsqHXvmBYUYMZ1ajtZH0wWfo7+ic65syk+
IwGyI7HJ3a1Y/uHkk+9kp9nzW7E4bnGyqpNkQiP1ZgiP3I6e4r6lc7p82E1gs7OC
59VE9NPol5nljxNo7csd575wzyjXaA5kRu+p/5Te66jr760JyqK0kKGPjOYG91a1
qrZ+uFmZm+zjtAedr/BGM/iThQ9B8q53cY4FRDncniU4PVxHXse1jZLxFed4wdWT
nSuA22lSH41vSUFCFm3fzIZOpYMu6CYC+ULCUWzp8YqXkxPYkLyFhLFUjYmTzbEy
5GUVLgPgGCtom5LIzCpKXLMViuD7CmkNJY1awDzO5aADTvlHzIWlHsJP6Ka71qa9
VwRssd7Vd6oEvcPGk3BrQ0ETdQQjSTN4vU0WHYBLeml2YzGZVgRuLQ/xhgnjWKvg
xRSiQHXTFS6w2zESeq367wdBZmQPE7STTycGLBZNstUuWERi2XRIwW8LGgJVMjVg
oLwjd+fjxAmCDE1JYELHDucSPy7O/yW6QXhSqFNHMsdkNYMxeTFYXJkWO9x0Eyb6
E0jY2ymj+Y7yIP7X1fFAbQV/Mwfw0F8RJhNXnBtCOpasnoDlRYZuiza8TnZLhBbN
+96m/8UVW22mO++FVUYiJ4qKAoZarIJK2Ir9DKn5RSyVBCvymBPJZq1mniw3Q8xf
EkT7C0v/dZ23dx5n7e+e25Nm9EcnXV0oRnRztdD+XbsHRJFzziap6zBSAduesFBu
Sj2Uc9tz95JyM6RzLlQngLuhfGmJUiOEXuHrxWhJjVTVRZ3jORdOgbBjZAFc+l+2
bBFemxqtKGXqrs+NIhT7IRFn4LzFyqcj147Kr1Q4RoXO9bBG+JLnh2cdYcZhwZ0/
i9gw1Chy31zyqUeP/ejzs2HS0prp8c0ymU6WZ7czchS036pPGXuvhodSpW9VKWFZ
060IOxFF2ahogsh2JSnORZgw7vQcLQYOgKefV9Kyr0dj/KM1Q6Vh0R4Yivoh8HHD
nPELEFWWk/sqYooYPBqTASUIjNHv/1D3E9NlgxADd9gJRD19jdzI+ihZdi3edH+I
DLY3I724M0C2QnmN+7U1JtQB1UCdCrmsVfukSPh4B9fKI+v6OAqd2zZlgkSPDiXf
Lqx28liDEj3hYamZ6hCxfiMmcR3S/4/rf/WbwdsKKcJwYAoPlftZ5levV5s+kKT/
qhzQbxZaAtB4urT3n0BQtpLYSFO2sDM2JLRriyNA6731GupCXHovaSsVXu7jZpdq
8WQWqa8yemTGaj0txm+PlHMDhrHAdco6IRIVQ1cd4xktSkqIauthRMgA/wygHCvr
shQr6/XE/qAnpAYYYw1jX3Pn4RSsNtJ4eA6e605cS39QAjSEW+6q0Oa+TgDQC7/R
r4joGqetSQx4QLadf8LhH045EXN4xTv9dpX3Lk2MyT2ni1l59zlH21xhncU9yseZ
rJV89T8QbtkQMbY+trbpN81sKn18jMFYk6cPebprimA06IcgT3V3s27yAQUeT8Ul
kkJmnVLreFeklwFkq56r3W77Olv5AguP5PODs5ndDaRCOzMJWz6+klpgChz84zvP
ewOdg5043gf44NAqmejvhx+RKuxxb6SWuNbTrzsb23GtiUI/yqEuCQd7DBhk4N9v
ifC3PJJJYwqBItbhZqShctpB+erPI9S435bkcQoiLM6ULq56U1EQ3xfjnJd8yAwx
5FGZkI7D2sY4EXqI2hDMxSGNqoytHrjGb+wkM5/24hxYHLl/Fp2ncTv8Z07FwL7l
izzpPzHwOG2yJgGHEoOaWYJgSDdOmX+B1pRADHXtWsTbdp9V5Pr/ioQMDzM5V/Ey
TevN/h9uRUacuvkZNyf22PbuOTTXbTjcGDGot8N3sh1I8EAnEu5nhM9CjEmncBog
H1nw1lmDr57Cu77VVBfs5aYLlr+wTVNgrNWNy8fK8Z9MmRNSuv/fYUz74E9Hgqzb
wNMV0iGtdVp1D0aMpkDWWhq/O2Ar8dSr3gX2ponHOHqJtRm7Dz21R8LBzig6p1k3
rDG99acMfDP3sO7GY6Fd6Y6IaGb2eFkUP84dxxl0yV/y/jBD7qj7+cD/os80iUxl
bbU7PqNRr4TsJRsj40OaWwTbptb2hMzFBsd9m6GU07L45+t7v5V4TBBUQsM4p8gM
399cs6hIJjx47sC8aX1isfF0IiT0JcCiYffgiZm1zAl1vMIg6CkZAnm4vwWpuLQm
LBmFTjXRbOZ8c3TmD2Hy9nCwgQI+kiHNTW6KXmwaULNzVmu9PHnUiQQMhyocA7cE
qAtyWv5zOkjp2crxzlcnfyAutc9CzGGUf+Q5S1OWRCmKdEX+3MCnk2m/YxV4RBcG
irzKd4Gc2W+sj0W/Af9DGeHXx4rUH6KlPM3smln7bW4/yoGsgsVvfnirZeOdN5Sy
c+oU8xbyaQTcy1vi3gGVCyS66KlZ8fACZXaBA7L/bUuI3Tz+4DrzqdFIyb2R/pCr
NiMaTP2HNBbopQpLkgktNu9l/eQu4xc+oNhZ/Mf8KNXBTNtkVdyAqdwpmSJc2xji
RQSkbMDP2/84lzkvQTTCumBuPS1gNkiGsOwgMDM+uNVMEKHN11mUG3ZI+PZoNETE
JK2LzTGvsFnLvo9STYB9dvlKAZneXNVrWqejsJWq8CjrK2CsE9H95EiScRE9xvbt
69x1kWfDGcEolHPaVepL2O1zPBG3DdHzUfmtBcoHwV7gSBJffnOzMWJ8P0sZlKUb
YszsUrDNKinDojYfLMkgbvLiZR0H9Wigo7P5Y//ncUAWO3TVmR8rOeHdkFAsrR3L
kqKK+hfgQ4Qh7SNLCB+Qd2MMdh8Dr/B1btu54oXoH+szkSIhtAB9RxCOtuRSfR6F
LG9VSPPZd2k9kOx9jM2lYq8Yuyf/gOcfKq30k8IoiAyGIm1T1MVrQYftrE3j5HMg
XdaB4m2aCDusScqBn8SopXvsna35fP3skofIL5z8BgZenB804dCoLodanrrTigSW
TrXtFLRqC31Z2kq61ygz6aG5eo0aRucLTOeIsokYgQdPohGADTUm8lRqqxrebusS
SiyMyXKPJh4t+oeiPzAYrOxHfY8QDyH2ZJ1FGdN0Z9thczUp6yFOjDJdANQ471LR
vmGvbKLmLmd0oFdCkkF8oyrXo6XmelfTHzA4mSrH/BADoxobSMRbW0CNAVSFexap
DwnkTSpWBCh6bnUIxwse8c4HYbwC/OzV4er0Z+nwkxm0ndy4Pq9rt+q72JyiO0D1
q28lrYVuOsvfH9+l1ff77ZHrwqg6apk4hMAmr/hrF7iK63Lw9evsuKv1MNy5Ezoa
c3lCh2Ka9wvAz2Pw8NqDmTeSy93Up3o3sS54y0Dh1gWRGKCBOb5KW3kpr+nzS4aq
TNSTtIqYpcSqyU1TsBJWhx+1mjJWMSpDM+P9qDmlJPc7/FJfi3zEqFlNgOHlNBMH
biFJ+Iq4J1TlFeq5cHPYdGsoo2Ya2WrPztIKiqDyoFS/lucPgkJCkxlF9gEG1Bbc
TN+YhBmElyWpA9chu90ajTnMBsT+xqSuinXqpX5IiGRrioRmI0ekkzn2wDWof3xT
Vr2zGj0eeuJ8Qp8ThFFG6yk/N8iM7YePWT+Ey4m3c3NzKtYlgr/hPxEcuuBlQihr
qTY4JT/pe/yTJmbME61/9MW116QgMKmgT9mRDvd5OzbkZdgnPESSJUN4VOvj7c60
pCLqfvIlChxtDTkH9d3kbfO2nvrccSqDhL1fEGc7iSJiL//gO5nJAt3pM6nDKtMF
FzUrJHUZlW4corbAHLbNO33WQyfdVGX/zH8k8pgknKv3mQO497Tp3oSS3cLadlZu
AQ9HH+TlZDbY+bGI2oYZWvOMwex8kPtb+48jJqQkPDMHfb5BT9Zw2RWVDb29JAcr
oiYXWzKm0WDNMObZ20UTyktJZLwDxXToLrdEP0suAAsg/87JVghs9aqbueBbI4Vu
FY509v9c7Q5JREKSFPU099ERx+Zq5Wykx6wO7QuXV2H1sWyWd4N21tOinGPXFv9s
Ad0BCYIzWvVsbcKEjPL+cYMM7IcrwbNwA9A5g6FzsYPhcXtZb9NboyMQj16t0hOH
+P20zGGBdBKqNTLtvaqENDLD2NJCLc23mOaQzlajvTWvxjZ/FM755W9PWuuhBIay
IpRtVRc1Aaiawik1k2ZfvzVH7MKVYw5n2cJLxUoSM2MnTSi5HZ2bFdD8ZZj/1qDR
xB4hWuouOt5nLaqUQNJq7qWVFF1vw/XeLIlaJIMJqcuESRkS87r+zanOFE8Pznl8
jVPP7UmOISWuR4efm3qWWNnY6CZTkKszxyRSI9pAekSgrh91gO9WITwGeiAexUlb
blhUN7h/bI3yxZqsULAWQYb52b2z9LnpnDMnE6Eip4GtZhD/2iejM8VA+DYxwGZX
54LxYRqiAtbGpr400wvjtFFnoKjyQXsi9ji2NZ7D6QaghlEI5iGUt7Uzj8v1vnlx
KW7IkIOHW2LmAKgCz48+eQ6yajwh6gXPucbPnOgC+01YtPQiDUKmNEbcFnsoKiVC
QOOah79XNwMA7xYWgP55jsQnruXOvhm22Ky79CAN42JF93zTXFABkZxJnOV4+ghz
8WljsBJZkRs1psLzpwdxHfA3g8ve/+zIS+c2X26sGXM1zOMY8Oh4GJZNPUa+APm4
P25Rr79M2f+H8DdQQYsioxhw6W6+tWHoz3j6cAO5RLijYvTtzGKcM6KI5fxGYFZb
gjtUOgKEjHkS0Q/S+1seUw==
`pragma protect end_protected
