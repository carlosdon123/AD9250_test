// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:22 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QcvJ9GIrxnFRo6kqyMtG/tEkS9vdL9mI7ziKqq88HkCMmx/d8DDexJ/pgJyE/qfZ
utqH+hAeAa8/Dvid5JJqthchAdmIba2NQf78S5tFbv8qoJWmBpwIqJ23t672CGuV
fRjK7cFGWRVrnDPnWOpfxLHhZyKSbOU6jcpxvipal70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 762336)
XqkI1uqJc4VmM6RWeQ04Y3yzY3zz6hmAN3DM3MKA+cSZ2XJ5KrEcw92m08nqyehB
+pUuiOiqe9gflIBuRxN2tGkwJ/0rTRX+I3uEU6/dtTgB26QwlacTM9n3BpuTNs3q
Ns5M5/GuEN6jYj6bV/gM75Hc64YZKQJZDK0iOaEhusHCsSaYvtzHtPw5o/oEPalZ
QzuM41Yw6Q+EUH1v5c9luSJAR578vwMwsKWaSu+K1EvHn2xBhl1KoFSVZC55LuaU
onBmej6VFdHV7ukZkMXJPn+1JMgLArZjLNN3R329d7CFvJ38I9/XzoaT1ZopyzL6
31ULPCQZ82vbt1fT0b52pqOgh3fkDbta9sqom7iQPBGcxJppE/uFJAT1fTPfv+jc
p6TXpd1nWOHMQVRYv0FTS+OPYXgb0XKWKOEc/y/YXWFg0qcHrD14Q7EitzLgVKEP
+y1CRyREPW9kXzLqizzJUNEMilXwWv3vomUJpQVeYr0C6nc5W+MwGkk1LpBA8f04
KjL52I6lHI6aIMGOa5BNtsPPEYAyZiVewuo7tus8xVcxbwq6ej2wBxEXgGafLTHp
p4AgrEghTrqp5eZrHvsenZj2J96ilFn07qYVytErgcCdvbPWM1t2acfSiS4cI/pJ
5Fzc+xxxAEZqaUGKfoGFXOiVclB1iC1XBLvHpIGgeziFw8jEC1Bv1+w5MWKejrai
lO8PYQwNFczYB+L+2xT350QxhxM00Kvd0+pnzAK5SgFWRW4VGg9LXUQVPhdJCWnb
m1/q0lBT8h7/pW8BZ1nFgRlwF3XMUEoBGXSVaY6ayotCGHrDsLDZAv3jrC6cEq6T
FlPfhRLn98StA3QZPqnsZ6gCz6Yob0PfmSj0v3FY/HQK9Mg1g6iWLr2EGezLHPaq
MwXhLOjhGYHoTwWoEkXr8+cEGJB5x1COre5C8Q0OhaMNKfHGxwGlroHAARy3ym9X
1aJIxADvjNoAQrRsz2J0UbqVDyh1iTF861bJ2nxcS7r46tvN7req4FP9kkMf6t+2
dAM7p589Zej+AJQ/NG6DLs9QpmktlIqAaw7nArWM0XtBgk/X/H3D/+TvKmAhLqBb
UL3bD8fDqvCjVpBV0XDWarO5Y/+hX+Td3DUw+d21Eq9XyK/jQuCDyAocPavtVy0Q
+AkMSQXn/IGuVwhRMEEYZVIKzVTRCW+cwVHjKJzTxzWQV4dIgg8JE6b09JaEWvdb
xk28OGeppXywQEfm+HNBUqIeCW3w+lwmlQ6xvBZjFCp/Rgh3Uh5tKn/4EnOePAO6
qICVRJqXGrZR2AUFO9UDQJMbcASTlfsBQ5nM9iFazbkOMsM/OuLf9WkXUUyo9Y80
Fw/MzdzVdyaTbCrsgb6KV5SpjaZMJfJDfKcoahbwNi80UNIDdtdffjh0XQK8tKBH
4WUxxjWYQUQxDLTPschvXCllE+GcuGbUJwMJkfFmRZ8zT18lc96jF94fAQxyKavx
qxMS6DyKXgl8logYIRNU4J0SHoydGGafTOMbqarPUXcy7viU6OEfbT7GqldWQrRN
x5wm8p5Qvkjr+hwZgjYT09UfkAAvHK4WVenTShwsuCigRA99BgWzl0Li5XErxfvU
9NY+Db5nv8U1TiX8rvbH4G2LKmMuF2BVcEGeWDyq7mRzrFhGyYQITIA9OH8S4rjd
wwZVX7YJksY+6OZPycqvOuIcPDjU71gAPsmtTZSpXg5ED/lZiUzvkPxiIdjBbroI
SDJpjDSarfARwk0kj7Tf2A82Cq+nfm4ek3DHimKyfCTGh3rzPjZgQEjA3jOlO5IN
WFISQnA9nB8JDbFAEv/VrMELAhRjqaH9jKT5S+FD4jbcyIR+XM0v6+nSqj4t2jrV
qOClQMyTu2r+Rr/50Uo4MiSKMTuQ0KPa8KdnG5Vd7zfof1cAvW3AQvHQHFVZAk3+
uvPFhAfZqzOeOwgtcy36ubCQLOhZGoWxCGtN6M6wUPwHaHCRAo2qkzSUFiQGQ81w
AG08yEF5K1xpkWbUltb79F937egXIsTARedqZqi7oA878w0BSZPRYhnwUO9X9ZeD
NrKku1IGIpyUjWGOs0d92aEgF9xDNv/8uYc7HZatFusl1MATZMdRgb0/bE5hyq5G
q7My1it8yZYAKnLoedrrAiMV4JxY5+duIEU8IeCsvSe7sFKf6Ji5Cp7ya5dz7vPD
rEoKBEoUNvOiPpmydlHCc6VISwIBnaAAuIV+vKjFAdeUJ3gHjuuHo88/RwEKI6e5
t2VTdtM/BwUb1FvglQZ9cX4aPa8QNOcceN4271oiy3VkfaRRq0ZTZvSQYXtI/fgt
WMA+qbaoDytA4C/R9lHiPnPji0nCRDP/l6HMJIWhw+1jbGMl3GZHRK1fRMeOZptV
IzpETEUlQlIQp8uAzxC4/KE1nt7YPdc4LUIfjPjkJD+1EO9iMRQt50UCsso/jBYD
k9Z7gI/Y4TO6HjDu8C+AQGwL4JGsS8GzDi5eRA7RgPHHp8IooGqYtnPBdJSdeJ2O
MddfjVZV4fRmx+A4UHmZe1Qbywyru0p8VhFsqWIJASwLNxNIQKI7aJeJkgbW+S/j
azu6YWIo2/1p1bRa538lD/bR2pUniSegNZ1wVJASPQTqPRoUWSWa7jaDsqvi41WD
B6sKmuMD9Yy5gZxLLB+jqOrY7aO8u8hhHLAVO0zuR8HTe8y//EdLe/LSonL4Sid9
LaFOzZwzymrQnoaPbaVIah6FRHVXvH6O572kopeJ5ZBTUAu6T0HUtYGkWD9ToF8W
Pr1rEco0K+A6tC3JOJGC6XFtnc0EHdE8EfbOe5GqcMoRYaGZBTD1VT2oUKyNfQrr
QXt4otpiP3me97+OFzIK8ht7KRDb2bLI5IouSljcvtfADcmwKJX86fb2HliQM/Yd
QcuT280VqaZjnQQnNKa3yM/mXoWLYHdYavFvdVQVQ5k2OMBd7bon4aaK2hD14VVV
oiqGrAWaKARkC270bzFnIf0ky54YHRBDcnzuk9kBY8N6lwpwoQKXdY0BQIlJnhZo
lK47i9PRfht2pzaLyP54PpHxOdv4pyqmQXeSRGG6fbRwSl4hJXyjOQ+NwC+pHELV
70+nHTTaqSIJMtJ/q0Lb2ekrb9jp9N41sOw1zLn8Gjh1XlV7ME2jlUQG8MgXj77w
1CNVyW7FRJsqV+S6bWde/uAPg1XXQo4h0GWkw4q4tlGyJlRlre/P+4JYPxUcdXg+
bcr2tD/loJeh+VGsH+elVeoAvplxzgeFsnkYtAYIVLVcVpYi66Z7O6ptZX9R2hmw
WdMd/WYgtRK+qsUH2t+FYyI70BKTBIUKeSb8Q6j30MHw4s/4fLv/ePcgIr49gWO9
Z1KOZ0+a/mpIXOwUc85nh7aXk6myiS8gTRY8w0OXQDCcuFnZtUTJjbKS7+p6Xqvy
ptqTh/1R4x347sLqws+3hFjmgm/JH+m25B9L/MLfctIVKZCFIsnR6KgUAI833RDf
l5numwREN3/KyzIICx9xmtMdozXj+1UAt1YVz+HeAvWecJ9/SxIZ4Xw0fe5r26+0
N++P6eCvM4hp2mRhe+TgbjuULJktGHsVFEK8GXvuPvHqazch6LSSckUCkzRa+k//
0gFGzZfCwHlydpYvuI24ZTdSGm84YX+1gqkFlS46M+UqnyDGL8mU44bNHf2KQvWb
eXXFfMtuDSSoik6s20qTZ8ljXA6RRW+0PEn7EFokI+wopFseo4mEX6sct/1ABnOU
gV1R+2bo9ggGF7/GQGNhzl2Z/L536k9VAqBEFm4Lk5MhMVB3E4e/XzCYgBDti1zC
c8RyCPZg10prweetKZLM+CUV7B6bYQNo5Qa8pp/K5lb3ccHCt/WXYg1kdwlwLaHs
KdiVJqVPG+QlCx+HARxChF++/XleXimgAkJ/ND4TcdwK4lFAlFvl9NSJY1AH61X3
Fum4vhVsXClAJarTXbXTe10Fjq+2LhNMTv3c8Mp63NVvFc04fVV+VLA+2htkEsVZ
55heeVeY/Pm2jCkbbYV3NQVYZaulc7vkHsShhvNBEnl0J8HMEF3dRgwJXEKgRu8C
X3f+cLU3UCB75WeIlnefJn/7h+JxkLtRvM94q4ybcKDmAs9X5/5f3aZlW9TIs13A
H0U6a9Ku32siMcOKvJEKAV96dO4CSwXA821/+6pQtEWl8rkkHLqYhyU1lEc7QYIX
V0MPsYEioP+MtnOKSxyDdYtiINJQ300d+I1DCFp00ENYsqzs55VsoeDNEgm0t/Gk
xlszOdYVaMQ3U2ITLTQqk4B24vJ3kvLA4xS6t6+RmLwD5BGNVqWubHwM6hR2wiGe
6S+oN3olw43zRCjT4VSYeCJAZPBjjAniL6UuLOBC305oAkj82T/IHHyvUzL5Yzwb
GpvWkjPzM8V5pNSza3HZXy9R3570VPu6edNWhxjdXpbr3FHKpll+q3nYnDF0Rpav
7HPFZRagpaCaWDBX176j6v9c8zWgahJR/TwQWQhf9bp+YGwiV0ZRlK/tup/AHYzI
SMh7ojb4DA2nwDcEufudmdrbx3p6gUgy495hx9CxAnc05yEe2kGX927ZO+pjfOM6
PL++NzdSIxwevoXVDxxCRi+q4FEARFdFnx4ncycaTb3JqTCtvTlzIMODKOKeyaKq
n6uQVnqonwAKelDljj1gggni1UIdWonZ3EqQygIQozVxLrZinbFh2hmi3FvNVp/b
zgdJCyO7SEV5emCGJ2grpY++MdUoJWW9ycQZlDKPEqEbZtNX6RcmzBdbRZ3ZXR4j
knvTdfSESWeEhHxqjRc/dbGXeg5OPZU87QwSLV49KR10pYUJfXHg98H//iNnoQhf
St/n/QA2Opzh+q0Wrq14FDfZ0YmyRzsOMpQMBF1+BzaHf4g0Q8IMG3aV/Y9wOEpf
bexGJPg1y2Mrjx5gTK4bg8M9M0ZdE8tUrrVMsJ5dF5E/Mjlcw8v16/dcMyf4/gno
6ZuxZJWm8UoSzWwHwP0uIrYVEyOOjXj3fLQdCQCcXnnIoEZc6bb1KTD1sOaPZg8f
QTkf0FBk8dIuN0vSXLcfZVildlPrEubL2FYImPy5Q8y3p6iI+0KIerQLQTKnxH8y
jPwaMA7KR+IX84P4s2c6ghvYaZ3uJLtmrzoL4aj4T+gHqdktYWAr+mCd/h8LShJ2
jVpDl95rTWibelHi2ue/Km5h8gjkIjiE8VXpEqyDZ130lqd1DPwX5myGEzafc0HH
3WECuhfEnZ5SiUtN0oVGWUX9GVGP+805EjbGJ6YkESV4saymCZhENbD2DHcMXnFS
plmEHHaZXWE0tKsryvPkCBSCjE/kQBeVECX43WU1SXZS8bxl9H/skHvcIGqdGdJJ
/wPaaWGXLKTveG3FHllLPkKIk1M9h6iqmkt7OIvJz0r1qEOTEc1faiKQqmm1I+51
pNR6XK0UKB+BSTmgZQM2CA/bvQsxIJsElV5zJOGyFuj/r46g1te5hzRYCy1NcBez
/cHeV/2C/WU2tbhSUCSvtv/9tQic9QOJxXlHZ2SpaB6JfeC7cRFVx+ufeuyCzrjT
RVosTRFsAGeVT8UDC26znjj61sCg0X/kKK0kTmR/hGzyoM0tsN/pFoedyIzxsQ3n
9ORQ2hToGQgDBb/N71gMHtqvQJuaMMfMM4aFOUOwsbHjHAKyERSMHvIQDODeeiRo
UAcHg4QWQ3A0P2rsQocVRFiSGKWc8riA3PM+qneUVrFuhZ2CFLgzAhAZYYx3PMmp
2UH3dJAsv7ikiFUqaFpUypxh/C72QaRChKIWVwJeVkIW6z2hzVoGImx4B8ju5xsj
OvLytzm6ndgwCZlatKeCOQ7vxvXQU9TvD7SuM1b1/LJeY8/r5JHpxq1ORPwBOiVg
7JExDv9LOpAsHwuEbR5vPwxw1k/V3JOX1CzWYQJxkpMkLL/NYOftBDTXKzQoQWc6
9xqG2bcu8fGeTjtR75xWfF0JB+5smF2Zmz8Fivq5cVNxtdkfwNpQD/kvyy/f93Y6
J17IA/+6G0t5xGWlgNLMl1rcOr5U2/QkihE5s2alRD951td81qFLi/GCHFD54Evi
5cg7HrJiJdVhAU33GqkxlwAphAe71F606Mt6yCk0BRMUH8P3RcZlYtqfqq3jLUzC
BlrMcVeD/zMgNk49j5Lt7MJjnIlugP/uvC6tgLT3xgsWtv4aagGamcBggyIMXtJU
fyGd1H05TC4kSc9AaXW1tUb7q1aBnwJj75aIfvt2hZmqtCaOeTm9q2NIDSx07cnq
H8ZLP8EcrxcT0L5DbL6E0CoqcxJ4OhegA9v7X5EFyiSubCxpwX6HdlP3EWCoxRhJ
jvBWfD/8hJ9PtGqJcyO3xwJe4sZnE8g+VipQjKkijBZT16KGUoJFliEQ+meWo9lN
L9iVifSHcy49/pHIy3SnDsHpbujRdspulZfV7krl0T2Yfu19sUqFH5KYjajrH+jQ
3LNLLW3p1dg6YYuGJV4U8f1BczQKhBjHr0qDFHt88Tu5uBM0uPnxUNf5YBk/3ig+
MeTkC9pXMewgWWVQNehrULGTuR1B+Y9xSd1xyAD6+TbC3rHjM1MJkhcSedfQA1+R
9kdFCj2Y3KtBRXj8Kv0JNdoEAFgohEszLW3CeX7T4awumGx7FNKYLNwUq30rfm+S
ZIjFIyBESzOpUUMpfVg1TpW1twFWOwS2GYjtvyUGkowgF5KDmqZ+1PZK2jmhY8dN
OR9lvwoGiVjeFkwCj+WPAbo/s1r2NIAUkvBD5o2ww3Hl/zthUo7x5yDX5kexK0HG
HdwYGV5b5QGG5d68BcBwBG1IyAuy0kSmAeBU2EqhhlvP/IA2guoLPX6QOxfpqTgh
RXgj1R9ghqjQ5iMBDaB87/QPIek8pFpOGIub78Av3yIyVyjVDkiq1KmWUtuxusOY
F7WMS95bUkP1hA8sniBga2TcuvxGfUkkc0z5VUsJo8UOFe8rAK8F9LImgA0FWFKu
hmAM67ogJV0j5oJqwPxbp65D05XKNsyJ6MMnhU+BrR6uqtQbfH17qQg16eaFej6V
X/udyh7+ZxZAVNEEB2KNMZFuT4FCRRcz8rVjU1qQ5QOidHPD1Us/gol5YTzaX5V3
xGsqkK2B2s+AIzcwY9YMo5AI1WOk+dpM5s0afP3y4I/XfssJcJYpFCnS8KwP6sxr
5MUunwIKbKFUT3OsQalWMRqp8oMiRAakRSJhjysQY1rsplrld9K4dgMBYcLH60tY
IdkKVaCs7EGWsdNke+qAoLtndnPg/WX6oYv0s//HHqx2l7sREdGM8diR9TvHXixr
BCp24GiwD2SnxwU+QFzD8BUHSgezl3g99L1x/H6BFjMHDmxziHxtbwxxCoGvubUM
Vv90olXbM2wHrlokqMBnAMIoCWLP63qJlQXJyUjY0ow3/FaYDBYu4STkJ1QdC54q
lsGNFw5c01537gDPWyFJQ6retXgLJYyPXKCQoiraJbmnKnmrQNooUj5TGN4Aagb5
/EjqrpUWVMdeuutKhxNfkPywTSXWvcQzJ396JY9khwOuxTkd3p8TCG3SNwWP3dlx
a7bfhqjHhseK0quBr+v8+mYHyynDEv938TO5OuMybM/R/dFh08iTImV47zRcpBjq
sEKQUdc8oES4wTz3peq9UIfugli9BPG+rRztWE3vjfiELBxGgbKkpI0hBbKh50Za
4QbZ+enGAhrokC6wfdEMc7fPVwcFLwUjct1K3wybUijW73eFBLGA0Y/qbXz9Lkiy
U6UVLwFO6e6L9YffUuH9cFSVrgLvTZp7u03OhMz1mS96JHyZZlJNdAZSYN7ibvlX
nFH/rSlNMJMw3eIJGc8hklaK8BOdqEbzDc7L6hZBo0jtMh6jPPpM0YTzuFbJZ2te
K/BUPNbjPb4X9etvBPhzJVWZIbFtPW51L0Zh/tOnaMYE7l1wksnlVoYSd5kg3Ltk
3lstCDdoLeKo97A4kojEzGq9NP2dFPpSuJqlYzaHtOTXD4tO2JD47O9WUPQlJgRH
Em5KW1XxJ4W3iJ1vnqIGMdWys8XhqlQRAGEXnHtskcJGPLAZnhr2hlCgp1Wjff+4
/IMceVSjXm5zDNRNL+6jMttcFB940N2HhPR+KkskT9Y+5HsSF1CqOnpcn7BrOpDt
Z/jX0+0k6kddkkYbyArpTouSfvWRWSCQXKUszBcPWwK+x8et8BRtNSZMUb/SvGOE
htIACZQj2f8vulkneetw5LPES0ruYVceAXKv/jcW1gGzMW9z2QNtUtKa/SGEnfpP
fN1tAcjA9zx6BCxkbL48t5EeTUQGDy39cC3uvIzIK0QeY4Oa+1XiPQUYTfxz+/6x
o8m+PV4x9MgWyQ+Mlul8iLgA7kDRjZ19DH6drqYLh8CHZWuZtP4IjkVvhKdhNvKs
XKBpz7bObNSSeWEfC9jmgEEWF/6tRZNP8rSiZ66o1QbiTwhJseiZ0yL0IxYVabpK
GRz1U95O3XOBruY+RU7xFP+VzNsueRDDRIy6RU3v7RePu5ew77ay/L17vMyepEeL
JBRN4IHf3X/MmmWpH/+GVOuF0lX6znwaY50XGwsthAqCCOAogYk4cQVM3wVo5gji
g2aGUKyN/OMqttoHEmjhlf+HmV4kDMqgQ01h6g9Yf9dR2eYzwwob6IIWEwlgSxPd
BdFWXWZQkrG2J5n+QuxyIeOoH+zeV3ag2CUHAzd7yGUy55fXeIxLSWZCoszU/sgP
dgURui++y1Z4dTGfGLBRFEuaRfQPniDBtHGCaDSACBNfha+fQAGGG6j0ph4k3ttA
R8uUFmWuy+uCL/oCv8bH6/2SN3p5Igx5HEP4y95EUysrbQJ7Sz29LhnuP8nTfBIj
aRV/g4tdb62JhKHf+Xf61c3N79vYfUILkuEGGKfBMd0w+y5jCx2hZPlA664AfzbJ
5GJL4YVELCElX82+GbXyTj4tQUaEaAjYjLz3vh5lEPKqGkBOUHhPvurBhiXVSEe9
RGGzz1RDWU2VBk8NIxbThB8jOyShQEGe0kfiVCFRv2iw/YQmngH810OHVtIyCF3V
IwFhWEggD5EjEEW+fYBGezPHTS+IdTf3faFKgSjt121/F69mCtDeGU5IPhOy8AvL
RG6NTQvLy58GmbiGs9tSs2rvsP1t1Ywg46Ki+TPRvw57hncZuQMqtW4uhdD6mkVw
NPwY4S4iWgmHD5S0oMx999YCDY6Tn1chhn3Gq1hBv9EoHAtHkoRz02KoED3gNO2r
dPrsdMWMSpFCAYggXkMaqhccGVOVXQ4T2jg/qFdLw53zCoLS3/SZhV/jDx7l/jmt
/5ky/2g1q8RGvDeruwsY6dvMWsraooTN2DVYHzI/7BHhhQU2l1f5jpp7nSfqJcMY
hid0CLwhlRlFmHLhN+YfFi5GZo8Gqs3Uz/bdI3J+XyemL94G5npHtjGQkUnwFYsG
i0jx5VOMs0Kxq4hnZeWMTC23axFnFoJw5IZOi/N3tmonHwNnGrlosLZSvSWSjj77
N4oOLhX42BcM3lifaPPl3pGJijFEdTX99H/hzoZGu1tZ89vSZWTQ9OxsaYmLY3XR
Gsjr9TuQntuvwNe8uoq5zc6Kq8vvybdB28Du63scL+KymFuV+zlsUtX9m+BqVmRt
sOxdxmkNb5hUqUzd5VstxWGrYGZBIWVK2mSmFYokmjAEZoJE7pRMSkC6xztFHM66
RjW+SaN8aUupf0SotlqpBPXgavm8m+2k/NKme9jVx7dJ6XPnDIgfTqZsgbn6g+Dq
wj44eKNL8Qdnqz9KeXge/JyomhBiEpROeCSwNoK6DJZLEVnpVTqhguda5t+KfP2a
U2BYhAeiTvC+G2saOubEF5HfS3q2o2GjQrsJ5BWvJRNOk+ejHXsIk/EAHHv78udo
KkjQ5g+cJ9dd5NuXGrCGdPs6LLXkWdmXNirBGQK8oaJUbQcioJXYItKim+IM2sCQ
beTr0WbZV+9SSZcszYndWjCjHJIiNCSLsZUhoCVSETVe6rqBvXVZeuQmAFcxq8Ob
NPyJX3nxeTfzidTsnaUCQsSlDRkIs7yDo4BXo6yyGF19pBn48bVQEv1gMgB1oqg/
u0S4OAlQ7i+NmAxAUe0vPcx794dzIPQaJOWlzTbyo0n4HJGCugA+nHhXYYbJp9Ea
1t+q8KfTGnduQuzvpyZ86PRmeAMVlEhRKAwM9BTkyV5No52eN5kiuaZf0eEU/dME
DorgbyLYb9elwwp3gB09jIeSG91YlZ4Ep52McQABokNP99bRR1wx2njA8oiAlkd+
sF33Q4GrXeTN3EfgMctE41Pi5zupd3TC9e1ysV5BdcTpd7ss0NaGQw3OZlZN914A
ceCqqNjHMEaTbK5yx07uK7DFc7wije1QMOi4xrbRhka3MzwjsFbEgGMjzswrNn3n
rNSu/rn3G1Mpi6esM2coO4dGDuYds4FgzpUEPDY1cDLyZiIwV3nnJHUArQCCPoui
ZFPlhJbZEQms6GQZcJ2TgbrYd5A1fFbgg2Rcugq+J8w75oehA6dpCo29PtTy5XXq
5GBPWW+n55/PjwzU955TTRsahcBBjFahG3hCfyBhJ+bWM8wWVG8Aefde3VwtZrlo
F5vRHj/9IcbMcjFwvdagSFZhHlCSBBugOTFpSLfwSNJQgJc58mVI6PU97MeZlpEH
7QEvtMwlw1KC2XobAzejcjx+c2zL61wBAbUz2hDNXrjwUa0OXrHEa25wWLM9PtZR
APrGmbEiV4QnYmZKO/w8kdpUqIofekQ0kFZzNdxDFiftPT1WpZJ/nclDhuZP5skg
ljpMUQJTGieaSDnP+H1P04O/u6At9CxgnlzjXm3TZUpnSFmSlpncPJPTcOhGdc/d
vu/m2/8ruvkgpRDt7hopDDsdPniD6ztxUeKXnYoOCRpLA/+jeWjkv4uUzRGiCcaF
wiYeoKKlTP0dOQiAjcwYfHyZq/gEiu4AeTGK528gbsIdnzI+vDDcf4DvUomb61mo
NaD7jSLQVPGyHPtMTEywtjbr/iKnxBQMklhqBBNtcT54UjEKrophU6ybPOcJpt/S
b5pAAuCRNorFkpGTaAoV/myGttgCQ+LjIhIwLCFHEmyg8wlJ9cqAEN9oox+ymv3N
PTr9gJBbuwkq6KBxTb9xQcFugHd2nXbC0qwvNYwr6cOXoqUxt5k/53sHEw0VnXMM
r4DT6PQSi5MeZStEljaacoVPwBotB3o0oY/iUDUzvYEEo1vRslY8Q9J+OFZfH6Hc
LLNi+rb5mpCEu3qnRtPPtmhhKGRjb8Umfhmqp5rQCKiprzeNy8ILPup8mJxCPgeE
AxM9ol08yv3BK36cjj1VLz7GMhR6F4Xd7NIQngcuuzaNOwEYko0UNGeEIezL836+
JY+Elp5NmiydD1Pc+QP0VPIH+RV+7fkjM2vTR/3d+/f2FVJksjJIS5lqCir1ie7y
jlhMCN658WFFBGdT2GhmLDSJaicdssfPEzph6OyORoEEcaa/VTQBPo2PSiqj+27x
0vfMr2NY61AVCQDNcSMTlI3QzDclVVB66DGTbLasR2TVBwq+Xoior88WBnf9V2fG
/1xgYJdk/RkXQTF1le0VWA8UHfPqLfcxD7pfbVgi2/+YbaP9gFw5gyf4j+vVDfLm
rf8CbRQ1S0nVhBXQwu8UvQ2iaEPxiwdKHoMqvd9XJHbBRagm/gBoS3EWm/N+4N5M
R8kaxIJWeP3LZXYt+tly+02D1pPRGFT+K/8/cb6tegJ4Mo4sVWonqRicFXYxrV7m
qcfQpl0f910QTKY4RmCqSPGac9+p91BiHiBeABWfTzNVKu06DBX5RiKhdgtHG5J2
yvnnkQT9L+lotFaqzrOi4WujTlj6UaO3OS/Ad9S7d532tZ+PPZ4tdacUgthyCVXO
zQ4liNGAN1XTSb0Xx0uhup/VdbjmH8Z3hOeJQP4zNuc1FRzGVTF3jqHns9KkzUTI
ZAFX0PR4LFudt1mFuzyNzugUoPBOrKeiHW+vNwJFALC8Q2vIfOXrB5yJydShwV2D
CJfPeJwA5DmcIKmU+DSkw53WuYtQ8LQOZBOFBUUTrJVHeb8jnxzWBCz/F2L1fVut
WA7jeGRJ+3DB6afyyTkD1inYHj2stCZyMvdQK4LCL7ZnZ5MygeFMilTpWfXsER0P
9U6GLq9ZUtsxRopOfKLTnrqAs2NogyGkuTwqxno6uT4GRgTRpUhOrJD+4pe8Wbnb
2+qMUteKhRRb3hS+GLWa2ZKdMlLr5D9wMimp4hZh9CgpKbmCTrbWpEqHjdKth0q9
xz+5xg5Hm/gi7M6jQ49nwoniMz4eeMw0xqs4QRcqM43dLY0hsZxYXkFKMlY8ISxw
i2oXpekZp0fWRgtK/J/AfxGtjwxGeei0H7G2iyPmBTZbUVRkRHlwffSUr56x6aS2
6KF+YXLccT2elk8NW3wHL3VbYADUGxosuiRW9KTF18dwzILlhZdCx+sGVPSg6/g1
3CNh/rOrNZxHdHXZHGIccj8P1f0Zrd97/KkkucbQb6MT5vLiX0gxnIThSRE5ULRH
aTXjHlk6zlZ9oujB4BvmhojRCOMidulE7C1yQl9ztwuqC2S9W8K2e7yhFKLF9YSZ
38W1fOVSOj7wxhnKmUzzKLtN07EcGLgWxRl7dqHGvW3BHh95PNiigVs7X7Ps9VVa
yQLCs6vjZs81L2qD/KqqtrauS33MjdJtnB7XT8jPZTDeQMLt7tbmJT7BVm9AK96U
J0z50yMEnSl0fMCp5+9CfvjzmDBakUDbvsumVeD3v+aveuuiPt8DlYPmvRZvQxtl
7picxmIw7g6CqPOIrQQHrRyG19LZTXDyUEo4q8jgZ/TyNnTLggBvcvnNT+k86+Y4
6eYoceqZ49WX1QuTtsNKiYH/zIigM1UAYtNb8l903w2AVvHqmkDABf+vK+slaeux
vldnoS/5JV1cp6YsEOPZoaZ4AoY794kv8ljUBb+GcJboAACOuvCJ0GJs8kt8OrFQ
lzElOKZ1VEYB9saNwrNh1Yh4qjLkOgCgro7RwCerwxbr2I9LRrrh4bhK0BqLRTds
o0PmiLyP8ftzTiT2wqGwxh3uhV9YeXOi/Yc485Bd1VZtJ2qxpn96T+RU/YVt82iL
KPUYsKMEkfHS7l1oBLvPgpekKjCHP7qFzpw+hj+ixuL9NXd2mZybsRSpa95Gt4kk
zygJr1cx8OUbqz3+HBUGd8aUqu8fezNvCfj1T1mc7DhaNOKkFNs5wsq3JrgGdrU0
q6Fs74BiuxzNxv3W3JL2HT5FMzqIBrcoA+dKtZaOm38XQ5/Pf/yaK7LYSF1Pousf
z2xtJJdIJEADWXkC0iE/30SO5U/O5ZyQCGbwebxB0auaayo87zrw3TZ89Z4M5FpH
tX/Q+oKZXyxfqQW6Bu1N3/iKe8KEfip4Z9Ki3zehdrFTG6x62b25TPRPkTMlHPtD
ShX49n4fchkMmQrT5PT2gPCWvQfXeyuH3a3VwnhKTBDMnDSbUo7LDi80ZpGbNV5R
yE3LNNzBlb630EQqixUaKViYIjRoDSWIF1T2T36Fe5C/gpYpx6Zut8b8+IfX6l/G
Vzzfbze0a1sEDdGLjh65RDtWadGuculxANDWR31c4ObBy81crEcE3DUZc9SxMCbS
FgugbAkapx2Q9Usnqd7wOozOL36iXV61Z0OQ3HNmSepV7kfr6why2xHqJ/LwtwPJ
RPPKr1Ay2145ovZzV9PJ/LSkmcxs1kodRqZWd7v9i+nQclNGOZyZABvxP8lJkC5U
xvThTjJIN/gZ7GLvJIhVP7QGyJLS7cuel0COFmG23b44tVB05mP8pLZLOHDWyltQ
A2snS6v4BFNcYaRosfWJmvjv9jFLlMwLmNHzKxujP5W3Q+AW5oro7r2K2A0hX6pS
hJUuMr05u0v3bxlSTNHWBYzGvLcqfiI2R9LJLnxHrcB/7QUrGoRgAWSglYbAPPCC
bsAL3gAHVT5xpBIa02it9Eescfy3unnnoyzUDDs645Ed1wCEUxdOWDvsp4tmtuCh
ODNU75KS2zSsQ5/L+D73PXeU2ubNyme4YIfSTFh1ckq53+Fr3m5pI2tNMnn4EVsJ
GlZyLsRtQrijNjxeh1eTgyyf/pYRXoqO+/SpNMsQLOBT/sGURvWecRl0bw6xhbt/
RiqOil+AlUgYXAhbIRvEDraTYNDkNA5tUb0/3CGUbga76Q7pmv5SvPZdNpYgI9TT
hz7FEzRKzlXk/NAepoJetW5WZB7OiMfz1QwLCOK5jEny0OlFwiMCgfGSsdbUwIDD
0/QGhx5DA9MMeUrhv7NsFdID6O5Jh744qvotFluk7tS+MTPEwTEGjQbbp4c1axME
SRV4vFlq6Ul0C8UN8Lk9nhO+I7pN9Hd42kQBGP2HqeadMXPGVa8XN/gkQ2n9FYAZ
Z80+qHlLDCAOVtVJM0xUSlZaZfTE1fZpAzgzkKEE95K2Z6EkhROc9/JNplRdOwi2
pJ+NhL8+uis5nvMSae/wyFLFTSPF8Jb4Sh44eAuwS4LV0GwUCIvslDvJb+j3+OxO
VcBCIKKULb8sxBzQAsn9cnppnygdv+Tt1VATgXu8g5k+WcAPH0CiD1WSOFx46zQ3
WZDJJBnAp7Ak80G7JRGdzQMkQstGOkyMTACjocGRpniviCImQGI+cxHcIsiRCbrL
TtvvkNY557gKUyCwWCyuTL8a785IQX/fyhrSoc8o2+u97UyXHy38UhfRRVZKm8dW
gH8N0r2beprBda8xu4iT9+j8Tk21K9oLhdVuogPpAJ94ageQ/z8babAwkjl03Qvg
xWSsSIF30LNWQdJWAy66ApymQKPaYAVxt7r8vhOT9CMv7IJpCqAWZCvpe1HwydEm
3SU2+gt5OeGnlBry2eoE++PpPD8nO+XRmjkzKa590g0vg3dN+4zs3xzywEIOljOp
v9kmEcgQDMtwDBUwNA0xaD4N1od5xMqQM8PyGPvLANVtKwxlbBQysVmgYYv1a9k/
NJ8womPJTki3Y4GIqtQ72mBdF6Wz+5PjEB8bMazWdl9E2xFbGpykl5fol8XPQvVV
9XglR3kTOUvhgdaYnzkzt4bgI1g1A9V8mnZwIBZPigxG+GUxV1kF0uS/v4CbWfOW
BYlOpVH5djROkeZsZDCBP3kROpWqwfGE8hhz//sVcMjebHLlxm1e7GHwMjCx19/+
1u27/LSSzVmhiL77xXfeep9ryQz2pJyCr6LRUniOf5aTbgWiIRv9LWD1wNYWpvZM
dE/0TAJqF/UmrSh1KIGTh93Ef/5Rj9KZJn7WnS+Y+GW8yp0/C0GLPUKdfsuWCK+6
svOcI0ZZ+wYgP2mvQTrbF6l50YvdBDFD9t91VqaI4T1v1l6lyWlr11ZBHfrgh9UD
cvq/2pet3fhRcmH/b7A2H+QCfP/7cuQfdW3OylgCz80YSRFQT/G1vErYFdiFlpdl
91nuQm2LgTNv5Di4vHNhshIZ0EilXYMNKUHrvPKapMMNiQE9fSDQuR39NCLXK0IN
FODlAw1TZYQ0dc8g+9ZGCKnAMKHwkYLY0I0hzFtaqV4v53ybhWgjn4QD5S80Q0q3
9SUHteUMnRNqNLLR5dU+7MZNW1+/sTLelyyEDN4L6FqmNl1d4c3S7Vaia5KmAbR9
v4xooFXXqbtYtCB4qhe3ML/tmxMpfqFLEpyhIewKuzhjLXUbZNySU3BaLMTt34+L
BvC/+/C2iIz1gtg1IsyV0kDbF02+0K35FDxPthKfN8tVHfdOxIUR/q7yZWlrNAlI
sEH49TYAwYxMXRIncY3zy3u7UlBHI2IAVEt2HWPUT5+Sdn+gIzr6Bqx/B/mLSfit
sYFdB/X73+ss2ykWr352ZzZi6BMz+Ra2ojsVJmsBhLS/wswi8EODPyONvwD17scy
OYWj6eX3yCR5ujjnVcEttb+R6eB3Qb9+38+sDBo7CgZKl4c7Vw6jQjF6uxK/2GzS
Yari9zCvCVImg1f1/RuGl8t9ZzSww8XRBxYZgsx3mRhf995rjBci6xKcwmKlBIHt
yrHvCRErzhynTT3K8Mb8h+YHmjzOg3+jlQZaP9TQuM0wg/R8eE0gpzhb/qLdw5co
SDRGvn5TDb5OnyCbMUDTTao3S+2sk+DbuQ5s3blwRd7WFnMsUSJGPobAuUozq+Lx
suxnQxx5FwMNKr0/sXeRa7cYQy4MSbOoovMSMGka9sMAZoQAmIHTcbsK1gbsUcI/
wVeFK2b9oXhaYBL2ChOnwVcRv6GYev8QVLktwthqcwu3UATOmGHFYIbbf+sA3g1q
Iej6orkGxS5YZTCb8Kwr6iCsIjMJCfGy7mgjJYY2PvVgiwoZe7eUIIPx5qOMGEqB
4Mxptwu9efQhjl1s6v5+7lKEv+BlJzK8BLwMt28W9QJanqBj/rB7SgnSZwFna+Ds
uFrZhrzEbwMHJrGhCfYBQ8hZR4CUWKgLOmKRNW3ddY2MyLvyMswgrAExZhP2EU35
rRsIHe9ktc6Muh6OoKooJ0WVTcAs2w1E9aG4MiBmEooSPLdGjgAOsQkjEJlftQ66
s8xDXLO2pILna7lrZdiocf64vqbcpFJvf/O5T1fBM9dhcZHWGP4FMCJSdCSituEo
Lb4nUO1TVuT7y8WgYcPJMgeM1zebjs3iTSnKwahqnNKRZzYwyWJ8COoYoT8Opmft
i2cXe6IuT3GNfgkM9/Yor/YyUOmj28I70i3uuzVCQ8zMc8qAY8Vq2+mnvJgyeTeC
eZAAU8UHAqvI80MtD0M+O0ES1iKOeeAiWvHAELpwJrVm80woHk0fJXS+6y0QaKry
wV7UettfHc+4uT5ynkmwG3bNKXti3o90LcyXVNIVmWu9iJQ0wkB2m4hPjVTAZUcQ
gc1vmwVkFu/IlUx3MwQi69meQw74jFdrfq+IduqROFE6cEq4Z2a1mmFHy8MSrfHH
n/3C632V82+vxxd6fZFB98PH3wRUpfhgG8efAbbGBzN4+dSxxvas3YB36/Cib83x
+MkrryH5IpXuRLp1X5WVU3BfT3ZZy+ObYX2NslIGM9nLRbGFZ+1eDGyyFCQaemFS
xJ8xSCTAIj31x3vQqMztSFMuYOHoIKqh8gaxe5f8AFHLdURvNVXQJYAhUudx/fhH
h4y1oLGh71Dj/Y6RvAP6SI77Bqz6Sw7NlinufRF7j0BYp6RDXlFprWZP5FQtQFyc
prEVgS2LcT4gZ7VwVZWeKYFU5FhV0FmI3vxphEAPaHq2EZfi15pqcsMjYuf3W57j
3GWPcsRgsBKZpAGNNJ0P2+XoAjl+IBALGyxZL9LzygVHYA0yS+J54o4SBqQiltIn
0FtlL2ITqaizndORExhrMH5VAGs0lXCcGJXTYV0d9eM7E1PBWZZVvdDUydO8OR5f
qiSMkKJoLJpRZcZZ3hscSAYsWy1igJ3vDYwtFXRfRtZIJ3HtvpMVV02KLLAN9ewW
2iQQ4a52EEuYOAIosJeGifScoxhiN4Zq10XSQcI+U/tGasCMBHkV31H6uw2qCeMS
sdt8CjJpy7vtbJOqrAOgWh1AH0SmtUpksHW6Nj3xFiwScYWOVBvqIkU15C51vTlA
t3/qnHQngxVvtPgXXuvfZU0WYCDTvGjBSfvpe/cnZQgRUGGLDqoJkRdczyoh7pH8
pMfDo/HPBtXxoAtHLIUCDFvoWTrmYHM0H8rMx7bqss+jVBjD7tNrbiKen6KAG32R
6j1Cxwu2W5RqZV0B5xgaRd8szwVgm6lnR1YvzlRxb+yjDCdsYl7ZtjhMTRvL9EwE
TkGg/YOZW0r2R5BEFWvO1Z3Zj4CXzZTx3oKB7GPCzrHPZ2I3tiV91PgopIhN4xtr
v5m2UsCHDrh9XoCcBIUTBikUfaa4/6cxvF94yUnPmTCrXA/M0l9YkppTHVsnO+wt
k1vi27wz2cgWbe9UresV+g6L2wNMIQK9u5dEofRJlpydvNm/i6P6FGrWuAfSeHK1
SRh134z0cpcqvcSHCHBhdfGC7D97vIW9A40vocRRjQQL/Er4TY+Ob4pUq/0g1nIG
RwzsReGT9hgcFNOz0BAvcXJp9rCIUbGN7GOZzlSR90PHNfI4CAx1EQLxv4GoLFUb
zUAqEUoNy7kD7yV1X+/oEIMmTTG9KZzYkUExV65s3SJuMDO5O+WfAgxLoqMXzP0w
2NLe+l442JMp2OJRQezd25Shb80AHpOd167acQLJAmCerMPuDLKU7IicNShHvJpe
KWVsSsdCEtLcfR5MstrX8FTd6NFx21gb1SIEAA1uYno3YoKvLQeAOAptandd03Th
h0FV5MDT2/fMlG+OI2WxNygMXtZL19liucObz2w8iBnCllbBFHqnPe+Hw+fyZwmC
a4AU96ZE+YlWjonjqo8v99mELIKfpXK+UTm5bxMbcW9Kh6oSq9y12eupJnkVvArB
oSuCMh0yNNYkfEJb4+05IK+aGAzKrWPCW4H4gB3G3ohS9WUxt+CuZoNVEvFl6YtS
fVqmhjN5n/kl3Zic5KjSE1eNXUUuk4XI0jdABBIss5N5HaemjwNdISlljxMvrvWk
9+NHhLFnK5bv1BqkYcS8CeQqeswiOBxYJkB+emeU2czy/zLNeNsq9ob3wv0A/XV1
e6AvSULDQ5fwSaTSiaKQBQM5ZE5i0y6dSrhp43dHH7n0ltdIEs7pWdXvL5jzsYpS
qY9aoCMJyd5VT/NTRHuIEeecGFB234wdHDzeMZApEG5Gs0BDBfa2wDubT2aKJy+e
3dKYZ/3mBAyqk2Aoa7jfL+TPrT+wLzu1qb5YCVxaWduIJ6w4zGq0LYZF8Nfrv6Fu
nlLe9JFhqKjbAwqL+vSzFTyweXkYjjc9Uxm6HvaTRJgmQHedWq5CTmOxzOx0w7in
ub+7HgwSINixMDg67B2m6J6cdDuWvwBmywOCLWO+63nyawCEq5DgiztJu/1InSCq
WXdFgNVKmmtuwLePu6UMTN+CwnREBnrTP8vKrVQsd4747lm4R+wshmjojk85l0te
U5ChRxUd74Re7fHSoXbnPFA8bB3oszwbfyZTOQxnR7sqTW6VHxrvU7e/ZFZJm5+o
fgZec32j35uuc+0VdvHHp0G/kUV8hluw/B9ZE32frXw3BIbpY+GCZpY0JN9xCf0X
Ca7rVCmQKYcedFYkZsgjGlzOSHqfndbSs3TijlQ+4CSD5AiD9R84URc2uSPXEqlv
QgeQhl6XjPnLYQcq8nDIbYGcYwEidfCcdhiEWKx2vCphSLvYYzcFgb+6tM3rJkjk
biX5iRks7udciIo3n2nG8JTAMgZSV7EOtImzV3MgxFU5OmA0DWGxdTlAxCp3bLpB
MDvvjJ8dmfsejWbOmvzNqEPhzaRuBoZuN7rDrNWwmqPJniu8yoD9aVKQHklJcLEO
4aGmzfeHdw5lpMKQxpwPb1bA4jfVYnQBoxU/cggvGfPYidQNGY3AtL0ka1kT8PrX
ZVbSvOXN9j3t8IdRsD+hMZE2pczGV8wODkFewMhjblY7coKBouaTKFr/LzcgbqUA
oQjvQpU673rsGQHJIgNpbl638+p+zCIBeaGt63cIEAaU1xvb4GD8C8YiF28cle30
LU4tabARjiGFhphzVJxI3COt4yplTN2g353X1nPdBMYjh8/iZsYb7FgQIyStTqA5
aDY6lAaIrqeXDHNS5WHnBS8jea/yxIdFyyVGKKNP9hHm+ds2dQbzSkuTg2wxgKQm
LxxHr5wLxg23mrQ3HWrDe1pA0JB+Zqw0qthWZc1IsFtlOH7f1+bFAYvuWlEjVo6i
As427xh4vQ8aQriXsLYyc1pvJUxA2Ty/2sxj2GGtELJiXJ7cWmKUCJBiKQbPNU6Y
XRUsuWko+d1LD9EQUf1sUlGoDN+TRlhSKSFWQxtX6nvdedqkCeOa2Xa34AI4Oick
YiWFz/QAmFh8GCG9L3v+2t4gf20JcDrTpp3O5X7EZpObd/pPpHyuz9i7zkw5qD9H
8xjkZnrRPWh+Nzsu1pXxTmmKf89T+tr9xfTg6m1jFn/8ziK64/g+qgqmf66N4Yxq
hVY3ppzJlHE71AXhIANcEKVo32S/E8/ReT/uTaVy4f4huOQigycxhkyauyqbz2Th
FiKgDuIHrnR+XpoCC07CZCQFkSALOk4dGGf25/qyYI2gWgJSKo4ArfltURnZUCZ7
KYDIDbmqCj1W6bmBqsOhnOacb7blaoGsRRJp6LQbVUIpXJxhjusnap9rfPJuOXK5
Qa7vLidEE9+opA/YuU8z8GqMULWO5u59ErTmbLlGgy0SS8oyVrIK3VSEY5q8ToQC
prtQqCrScWl2MWAoivvzGHnDTLHAdaIs5Hf1CoMMlBsuhfQsAD6Hvb7M8bN35UGz
0+H0zsdlJqaFTaio7uNFMt7he0Ht/7zez0K882QZr2d9m2E5LSRQngHlZjunUK2m
v6gLMRPHNqclX8ZBrJ44j2P5QdAekbsx9JII5YtcgopweVbhpmD+u/KShSe1O1MI
X3HqE4NBjFuWh1qLFeyW9tCOZtsQXNQ9bE5MuaSCZPinI1Q4sgZHLtiZpjglLNJT
lzsjqIS75FAohDCBcOnxBg129TIWwXrUY3I/c0X4LVDhufNtKvlGrYqy1Hhde6QT
8ZOjCGPU7gE2FsSbDAHSUUJeg/HfE7ZCD0EQVOmvf+1j+QgBnHo3wDiBoVcg2ALM
83q7UBJNLNWiOBh2P4yJukRgJQefjUi7wRf8weAVt0B46/VWnGrIVDG6QI5MIo1b
j2Sj7bpgk0YuPh/4esdtQjvqwLukzIMTxTjoHzZPwP+7JEBKYCKQ5s3a3cYZ0+sq
mLVSlPkIFGa8dOpuROFDgYzLlwyR97g2emdTxyaFNPPg1JBLsJSYvjb4PDyrQBR1
U+rodArdcFcliDHchCgrurcz4djDyffDe+YmzvV8zWaajfBztvPFsY9tIikI6jeo
1xWFFOXLIQqJyhvaOMwo7yOYGYS1b8u9LfSLYWFvnCMnDCkErVtht3FLtDTsHrNx
E38kwBmV0GVLpz3R4FOYA30Tt9YY3kQYSDGx9lfUTvMXDc0i8sVXSRErl+PoOhho
H4DpTOWvKAKyU9jQPQEMl+ai/u4HXcjyxErNtTK3MYxQwZEoDGERdpvA+AN5R3Ki
FiD7stNk4UbReTv/5EOIsLSVh6qCPQBnREsq8nUXiPLexeIvjydLuuZtDE7D4g1M
RQl/HoK/FNh/dsPhArR7b/PYB/ZWBl+uJh7QnxCARwUv+cCgcz+8cUP4QSqbAKs+
uIFAdhrOotbtb6wGe4F7a1zfIjrT0uxqFSjWLedcX6bscJX0hwug4FkgYSkRqkkY
U2qzCX6F7/2d43iW9qMpz+PZXwuCB8H3eVF47BeS99R2sgteiBRb7scvRcRjWbA7
3/0aLgFYoD0LScJWK+U7BqhxC+5fEBDCQPzIjGxX3t/M1bWyRWpK9VWQeKWp1Z9I
VCtA2JTmRgztsAKldsJoAGkNCFzhFcpu7UMymZT/oCqFj5IG2ynt0Eer1rdPj/yR
sS9SI/E14BDEGvkANk0CAHHbhZRo7+v3uTkLhlDZEDtV8q9M8U4nASuskQ2eI+S6
K1JkrOy4in0cma842tk5fjhViOVwmV3dWaaJye+uQfuHn1/wf5YacIKW5dONSxGI
+bQ50mV0u32PUKt2tGXHS2iPoJ28fcRsDN5IapGOnkynld+X9thasjFopKvRr/wK
i0a0NaqYjAKtafkEo8QNwVH6SORCek3voPwAK9jNUSRgc4RJQ+82+5LsNDEAYlsK
DcoNeoD6iB7Nqk0w2kUx/ppLxcOz0Jzv2jO1rWSTnLWdx3LWclxvuXtuUsnh6qsl
qPSkHytvE7KqAvsFR02F7CUPSkhSo7cZP0Z40ym9c8v0bMX7m9a8DS1sfGAeaDb6
2PWj+mgK8MXHL9Qvb5WW0SskpnzrQuiw9jSc9HjZ3P9fjg81WKeXdc/ZPMTqb6Z+
NeYBhbgknkg/wndPyRqE7aRUYuU72ESHpvzDegpB3LFt1OaViIcO6KGvng/1E8bT
XuXmsDCvkNDke6E+28wZTR9sQYC+p2Vw2AcPaeMaAvzJcr9O10GPV2IrqNbDD9pF
NhRrDDbYGzcUqvzGyPKQGBKtQ3hmAzaP+op53uB49NaAk/4SOyjEZuCHNN70sifx
ikpUMDJS/r1q3MZxBgjZvNTHShxnKgKUe4pN4D7YvzilgYYhnZ+QZQmJtTwk1e7C
XOxCrLzNMxe6YfZdSQR2sa0I2TbJW3OF6AzE8AVmGle03HGds6VLzILPinWmbPlq
5+VnXKcUsC12/ivTe4NHpMQIXsi/7xH9xqsiOJW1czH1cVaRG+fMOKuyoxolGIus
/EBGedr+2ycAAXFN4/KdWT7CVBdBVOaYUZ+Eqjkpgr2rZywFm4YfWwNu/1PjpdVh
srw93hVMyRNXaOA/TCSvkNHUCsAWCvVG46lEHjnnpIH7qHmDS2h4emJtzcYfmPlP
o7yi8VOZF4lHhA2q8zDOHkFkUiHVCQpbK1dDmyYb/P4zaRGgSHIArHGclQQhbvys
bEtwBkbikdChbBfahkExcjLKGe+MvxuWvZ/ye/tv401abGlJrmxFvxvTQAGniMF2
oGSC/aq5r+0thCpuwsEnTE82aWIOsNlSvkdE+yU4j4GMuKI0+p05UULiPs7TuN2D
14G553hsb397RI4xD1dl7sKMvca18yr306cd0rdOnoG62zDkQZ+6mPbUEzkYQXLC
ZpR9aK8jrAjyvOaXohMJZL4UAbgGChDb0E7jTsMsY8S9hYYYzVXJT7KRgovmOsa5
5hntyT+5U+OKMn33bgFJ/D5pN5rCCggxyRWqd3L0QutdCBEAxmLgAvxOUmFTaPyw
JVSFA5P+kJ2xyPBvj9rgxwM5ecWz3lekzMeliOpRsEl8kpfpVLzf7s4mi7Lcvrfh
cV3l2XuCuswQQ7Hlbnj+rBwBIcP5E7P47bYLVFNMXfoFt17CAdCk0IJJBsxfbOYV
toRc7tKHAr6qKSH7QYZ/P4dO5z5CfdLNa9Hq+ilZcVsavj124LtCHeUvu/MDnja8
wqWrSTb2Mz0780PvLazwfihRavpOgyib45obezA7bECMmCyJtXGy2bDra+QNUldI
IssfrxlnRxbgZRFwP8u9Zlrin6OzN1sS+OhzO2GfexjZ19/ECmSOoyF1dtalA/gA
7u0z174aruJ4LxeGoN3DVBHGJzYxXYnJUKYvmD+suDTDhLp2orGzMd7uGl6G8ppK
0v7mqHzfKqvZt4UWxaVSRSncwZd1NZFiB3JN9cdun/NIjkmwkv2zWy448/ZHl97+
6KJADfuGXiNCb8kweVj4RAvZvyUXJP8EoEKcxkZKzjfgqrk0NcsOfmAABgoo/FXv
DowVve5OPxbUmEjOKQ0pzckruXcTAH/84mV56TLi3X+xykgN2UxymvlFbwx4jtrh
bRd/zK1MJL23A9l2p/V+68GoMa3beMcmssR0wOpQggpiUiWPu81Z3rUbK1xcuXYo
tEOh+OJHq9rMmYam5EhnuOoziNXBRHV9yupcNYYb/mT+DF82sRWmjkbklv36WT6g
UZK7dp3faadj8c3AsKcQOj3FTbo+VF4fdxp0jCwj9PZtZ56Ean1YoKEbxMZjBj1/
/J5Kuk8s05nzAczfPI17zsFoqujBjO5ZJShT7pZKShgWOFctQjTW7bBQ3FIJrw7v
TLNjNPeWOHo+bDdsLGXpEneMjK03tWcoEcvyebYgDvbWUyNHHx2sveN+TAHSJVjD
XEXIDDHdp78fO9mBphZNt/kvwsw5XReCxsOgXJq0EopcGCBsVAvxPHlpTaGoGpJZ
2+HNzwSt8Z7AxAVCSW1hpCV6nweO1hmJILj6+NiIEHue/8JFdhCAzHsMzbPhngM3
QZzBa3EjY1XJBJr45jJIJatyUYBA1xMYdewOIWDCVpuC0Im75Kot7Oij6AAUeh0B
XllTYm7dfFg34p2/d8755CXNOSweab38V3JoZGJoXcSV/ucS5JcU2H0mS+ThZbeZ
vOqn3Pz2Yh5GDn8xiPMCC7U4vdhbyAXrVAhB9w5jWU2g4vPCW6UNv2hxY+0FZnP0
0gY3YkdEjYF/qsB3w94iUL5Xp432WdHA9Y1wjpzSLr+QD/NpZW8TX6IUF7j8znvO
pv/VepC9ImGYO9ebKNi18QkmihEo5wG5Lww8jarSHXJZMgd9OWdxBBaGdU6qcw68
8MtOwX+8DRXNR3T5ilGdU7dbpAnyiJGaVzafJwBb/GqEn3efcM30IWJH32DYC5tq
Uvcw8uSqvXAAe5vY4wsbCVR93/9dlAI0OvwEayGmqOgtvAMSaQtaheicME0L06fN
hEjA5T3TJ7j2dFb54/UzOZl8ApOkOTjMhn3JIZX0eF2Ys0mCAmelQyDqDWx33AcX
jtqgXTS34y2u7jfBXifpHP6bRvwhku1Vukzv7HjhVIbutKHhAGPNhbfOvBNfwIi/
f/pzkIOm5++Z0ua8coGpv+RGYLkKtZ4PDN4E2Mjk6junwVtESKJbDzWPbf0bY14j
JgJRPBs1o10yJCSpn2A/fJ8/UxEhcjhVfCZIhwYWE8XpV2ITtIU91wycQezxTXEp
b1Qwrkt+5ATiT5r03i64e+Q/Qtk1bEGWNOHtVmsB19QisZmmEPly7wrJntbotbDR
n4uRoIfDDx78/OhirSG5UcvbUdjHHQI8/jwnw/nCJB36sslwu1Ma9r4qtqMLnfax
o1Vo3ZTxoO6y2VFYTJrMzQALgpcNpGBwiCvbpIqvLd1whju9uXwbENbPPaVSuqSx
5vGpFi8gQkDJY35yMqDyDOFBLAlXoSww1hWpR7l72yP8DLjGXTXmysb72rCnCWwy
YyQy6PEO8JDokJMJes6o5fDbAMDfJv/hSuZ3Lk50kdtixj8WyioUcivxr9DPp5z7
oUpaXm8WwfpM4atyL+W+LEMO+UrIjBH/H4mFDp9Dk//kF6lzqkRD/fdb0QR8ou5c
1XoPxhZvqJhaG8ALlVeTLE7UdB2a3Kdv4PA0yZooQKujqh3NojsNfl6aa9Xd1XIz
G3d99Hsks9jNToyTL+COuU0c3D5w4uKnapUjxfodxODDoQp7Gt0fKSSCpuxXbduW
CRI/RDvbRjXMBNGiYdZFo4r/cK7gzjt3RoCZ9zM4Bs3Cg4ExTHKk4o3aGS0GKHBU
mrDTqg6vKkrKztmRoPM1rdSrcn6sW3BioaUkuv15KXmKROt1f3REL1/gdqQAMdTF
4HT6RxBfn+33pYO13IVW2/JMUbMfpgyc+PG+04Gdi1+rj/tzXQUd18aSXtdAGYXd
N93Q3d8VrbhuwDHWKtpSBP5OQEPAwNf5BDolxyW0wA6ZZoS9WXIPchqx5DzWeP6t
zQDfIQYmrKga1lWX79xywx0DH2Yv8uGo29QXQ1c6s54fJVueFV2N6rsTadC9hlmL
b865aqcRgicQxboBi7QQ84LQBMqTf9p1cN8cybZVakkvwaiB1uGwzh4yo78BAJdQ
BThexwyNsjZiGWl54sWrsXlM5o+TLZlGN74e8v5GDC4EFspvjDPjKyVl+EQCZU29
Xp7osI4S30KncLWVOaRfxxuFuv5sgyPM+q2iRWNvsvSjNfgeZqRkxwTr5wCaNaCs
pyFm3h0qKfSzyMqR6UwA4nPmswouZoJwkvqfoIPCAKumyMuK3pMywqIncFCQwWKy
0YW2bKnh0zSmn9FhfcAhURVi4wX/k3wup0WRHiQ7ncqdAkeRveo3mwDI86/YLo4G
NX2YtwOVNl6dB0ncSuXaPB+y/ecn8Qce9yxqCqLCKXVpqFXr5D6XwxaqjeYhdcQ7
tMaZr5l18Z75IFYzKGxincXqgLl3oueBYMlwZF0XO22mIR7QC0/gBxmOMpe0qzlN
G+Q9rGWk2s7c4na0qnmbb8/YwLx7P/Cu4E7yMJkpPke9r8KXe1GAUY8FuYBRJoIf
clh7tiI8zSIkNNYgFGueSh0KApfwxNElZM9nxaDuhnTud8gDZi+KmFcB+P4FP9SR
iFpyXVCmgcYKKEym7UTAvF5gbB4eqkoTH8xUvRQdgRp77mLgEtl+Wvah0rWfGWO3
BT2cmy+W9maBLVSZoXwdPlLvnPOVJijfgiAK1N47lgKm0+8prM1DHtx/cubZvHOE
RWt77xN7scMqNUCvui2TkteoaeIoQb+d8sxM0io5DeCnlN+sjMLvNLJ0fFNQOgLM
1dId/K391P9Yietppe/PssvcFfi/frem8AUOQ/6/ws3lj7ejkKmUCCeMj3ugGfg1
yu3NuQtJlXjm0c5i3jwNY5WxU6Eu7htSYgph9flhqK6rov1WG/qRffdCdFunyXIg
9sc8EKtkvp/xP1Fb71bcC8/eXRB7aiGyb7ZUWy/rTHo0DSuEqNJ+gdN+wX9MvjKg
rgoGwX+0Rd2qnykx6X7btr1v1j2akRKv9UPCU/42OTSDwxHkK38boN6Lznpun3t9
afW8sYiK8iIlKAf0AlG+IvYu/C/Y5dfjzJJ0e5QE3BsHl3XvHvIHQVyPZ1F+eXt1
Oa0GZH/cHyQrZOMt1ENveXCthyGK7Qv2B2zht27UpQvU1V9YP4nztJqNfq0kqElf
dp3nk1J2hJzFTEThu7/e2BwMmkIqgN+Gu9Ms8OlGuVmHOtQsu/JSTkxdn16SBAOt
fpcjazQQD1Ct4y8+2nt4mZCfYAekKAN/2B6shM3AzQcXpvPgG9thY5tINcVfJwYG
KFBljMGAijmX7jQpsxciwhAeG3KnPt2WD+HDQBFPClE3SM0q15Z2W7/KJeeb7uG7
HTvNFV1vSll+A8Tcbkp2Bl20eO1olrOE+p6kY3Lk24fLLmOX8CNYMGSy1nLQEnwo
GDS2uCNPn1lYxD1WSe2r7MSJsVAU+ArBtNc9kRXbxhv9gZEYPnHW8N3iU0pM0g1H
ZTcmnmu0lUMkFt1rGPVU7jQ6I7tgVCGXQH2Bag2KbESYxEZQKhlDC55bm5SP2Zc+
BifZEWeC6FdSNOpco0g453HuqciBffGEfGFTbZW1ExJiyi08GUFPLNc9lskQ3+bT
4mdcNLCpZ+O59xgA7uf+z5yOCKmyKZOWAkIfFaxwnyf+GkYdbPeYDoAvJTlHKDv9
ubFonJ411OMnptdJaG+6LXyuvGolv9ftusmg/fPJtTiL7gdppAWRt/Q3PuIq14/j
j7T/wsgd80KhRUE4zGafh9qgjqXyqnxgilXLtS3cSEkbrE3N4ZipoCcSRI7+lHRz
DFLgO62HYMZtMEYINvBq8QsTFkW1D+N+u9ps5NGTouhrpT6zRu5nRWJkzGL5LnCW
MWfGnucvxvaUqL33G10eThcevzBJ23/9JMs5q9fPoZZh1yP3/z1Af4t3ceMfnZKU
Dz4ivhw1qzVCnK0uk1aInyDX43hy16wrSs6ITJIfDLBmnFM4XDeUaL6ETIzO/VvI
wisraAlEOa4EEQaiyk6DqNVV1Lse3iinHlQ+K/NeOhjwp96eK2fSfH6f6i/smK7T
YRYOOdLPa1qdyHkGjmMa0DV4yVGF0ZoOrNLuti1NQ57IfF8XWn+U1bjPAAfYlJlE
lCFI0otClWBiHxM3gVcLtJwtf88cm553OB9CVm3y3GLt1vAKDfp5RAycrh/cI0XE
zcSywb1mjuaj+ZcODLO4JV+VtjhZhb30o9KPXtQm5wQqAbFxXYtmmxESVMhMhb2q
S1cUgyCiLJhVuO6C9eUpQw67MXahfScUe0DCiA1EnyyUqSsOJcR0oprd6xPu3515
6kbdKB6drsiNoBqb5KQGR/stLzN8hPwZFV1XyHyqfCZKwwpW79UEhhJwpnacfuMt
i0qxy30AqFHyf15woyLh6T5Hg5nD+Aq7ACf6rK0y296JMIdX2ewwl2xEijBYzJ12
pIJcih8Ey//sHn44KZKrSa2p70W5Ba/F0GcGzJ7aI+wjI4LGdWKh0hHkBHcYwZrH
pGRJ3QhE4kRfCBqqvuhW95tVi7xlLugxyVlvPO/k0rOG1PK7URwZ7U4AsP1Ee3sF
+uEV/eseIzNJQ4ck7CwLGeuimx3FMjCb6Wz8bOc+HV3iSgyCgQwJXzoMepBs98+J
3lMNHRZ9pXol5ABNiE5RU2xs8GMxiFt2AYl8pKdR1FC5DOSUw3qjRetm42/USc6v
ZLPe6uC5RlUIeMcYSvTjpJENcKZfe0DBdy+wd9CNMDdHuJMIuM1erjbKhNgf5XQz
eqIKmBiM4p7QshA2AVbAldK/x4WbpWWdEKCJj6KRqew6AYC3MIA4JM//akfscXjh
SZaPBu4shAM6cjlnlJYxOFtT81S1yy3yg3+H1mLGXh8CE6f3My9/Yj/4KL0L7EL0
jPkN8if4tvP4B+en31aLPSqEFJZ/Dpsgku2zA+MP/DeiU0S12DU50sZgLXeFRq3P
oR8Xsv2y64d1q0ICv46yxDjtxCaTevMqvTf/hcR+XjlyZvHEKGvO3fWEubzpoAji
m7mIa6b4+8CgOn8poCGa1VLAmDotCRoDQE/XavB/QKpSZZ2psfdLKCCmUhLSdYg5
nvaiLouMnDJscJON3BRn3LGt6lFYtGYheoGhrW5/1h5InAZOA/1oV1k0Ld/bDoKb
26+SBm8RkJZUADWdhSJbVTgTq9UfGSnEm6An/sNDAWxWLqShwEFwz/2x9vQGQqoS
prtrzLmA7Ptp/n6JnV9ZJfLgeOINDLJv+9nV7JG0D+WLsjwhgQma1kGZ6eLNXpd+
/jtPR9vHzxizgDdYMOdlBp2rOzmzbgzwuOGmvos2NCj0tYvgHj84NjWYnYMDurvM
R3eSZZedmLBUbTcEcCuGJ0eS4S5qBe5J6sT8kGZYAbmeSrexB8haaLQ4dB3WpBz5
AuF0F4ZIZGbZlKMiFGtHoZOmLIiaG45N960CZh2DSA95AvbgelQdkG5jJbOM+e2n
zqGT7pCsJIMXp79hlbUKdHTWuxqxN2xMnebGuVUtR9ohd89PHY2wJwv8xvpFSohj
hM3T60SjxIvWenRGurzHWtSrve6619eI9wmXa2NY2inOyZOkuYWuZL6BF/odQ3Jm
QT9G3SGirjyPWwa4wxTZUBo7BXHQW25assJ6oO3J2p/u8DIJ1ADWjEtKQxrnZko3
Ib+k5FLHfCkOXBKQMDHknXi8snyZmOFJ7GZs9RZ7N3c1Tk52LKEXOgewQSp04eZ0
U9TT5J8bqv4bSzhpmYxdu6rOmlgDQ90P0r74XQ5yV7K4M0SqtrAlYEBOWw16R8sK
pF+SJsXf78VwJGjP8U01hMA5pb68TE/xzBMsFX9KJDPUtqYFcf7anmX5PeZ/NbN8
FjQ0lYlWf+ixk+ssWOehBX43kabWLeUam/V25Oak5dku3KGeKU12xowCLEQa1tXJ
wTALma77Rv91Z2okyMoB9wEh+iO7i8riLf5FL64T3vG1GbdyMxxxeC7XppqbAO/c
+P5NUrAnPco1k7JVVdaEHwTqdbiZeHvbxphCI3RyFpHwjIkaqEqiLRuCfJioKAnu
ushaAR16ULZFtbbM9K9hidPm+V53BQ4T4DhIfemG7PZyTKoOJ+FtEx/NzsCak0LH
TphhljNG8hlFTJDPKeKtEsRUzg3Pms3oTuNeg4zrhxzUQFIRC4uhqlq1PzevK4GA
ZyktGHVlpv0LogzCXGG50x0LBhMMnKbykb9V5ojbqH90N4kMXr9EEdBoDFh75QBK
Pst7gQBU5gcX1LYacQ0ac4b7pf/qyxVspj4CImJlzEyHzqX1mixfu2557WLiOiiv
Wcoy+U2U3QibLbXAepUUch54dMijSHAs0R7MWEyZf9KRM2qMgfO3cuICEoSKjVhM
nvehDnXepPpV3cFe7mQmpvAyaRFMJSzZhXmZF62i5gQ6fdPoZh7mj7jk8PiKz1i6
t4L1Tv+WZ9AW+kCWGiVE6LdT1GleQCLL/b48NCJfjZk+HgnQOerPkLOl/cbaMqVo
aBkiW31BsOs4XirqzA9E2HXTTPsL2gSdUUEO1QlgoknyaRQfUAXQyKrcgImj+hXX
wpR7VnYS3oWaaQ/e5AELFSTsgCO5TnDSE6rEoxGQ3pIvR8Umv+voLHkwj0csNIos
x/eEMAaJQ9xAbDyg5WvvgXZd8BL7dRk8ifwLnSVSTVn2KwXhbFVc86peW6E78NDs
9Pw+pr0CfJ56EfbCbIE3QRGY9V8p9dPgEq947pGHiLQ5sO50lpthyJ8hFpgqx2Fi
c/h17acSwLVpC/wMrnVaBuqT2FZzv7s2NdGteddJcaKYViISYS/owqdRUv4XoqBB
3EMgF4T3WEOZa8WGRvD7KZTgYmE6EXLxq2TgMdpPtbsMzj3XRhtk8zOvUS4cndQ5
Dc3w4XpF9DVU+S/PF1IsNi0CSuOcEJAsGFB8eloT7tTsVbFFms+RKgXftSU4uJJX
h2zZmtULaPNGjysXQSZ7xtdHADs9lCE5J46vXvnNr+Cdh9Ud/a7CMdHVmIBgpvrn
0QPXOYteBDhJYpzDNPTRQ0vTkR45UKorhAR3f5vbdstoFn+TxZwknVqnIJMQeTHc
gofV+bc1CcKZkPho0fmRN2/XMB0pSKwSyhfV+jKq1q2l0HCh5Hf8Odqn+DYSsAO8
1o8wewRYuFE4gF8JE3YSryVTtD24chzpyXecpsaVv6vlQGMDACB457/N9kLnpKN2
CO+pMy8Thx+r4HxAkqjTvDyRU6rBvaMfPptJYs6bQZGVHZYVmDXshLNmzcsP9717
gY7hE+lmTh3Hn7U0VuE79Ewhx05XX9olTW9QyVaUu2CL+BgVXOe59xBxEPS6QeGA
dkj7jnfaUnukqbQvrCj80Y2ffMEbc2M4pIHNblVCw09NXYNvq9frUzJs+XeyvY+z
Icnkr4JeCXxoZLT7by6SVChf4V6OLzEAAGGK65zacgMlllkvjMkQKPlmqSUD9vEK
uU0DwxDAqIIm6MIzOtnkqVSylY0DSpuG9aMKGO92kSBHnwFb99+nr3c2Aj3QgF2H
HFYnMcVtAL60o8rpiP/OVLNj5p4t9n0YcuStSuGzlaeCPj3bQzpTzVmnt+b3TxYo
wl8y6elhhXYasDPj3h87K3Srf//0uLb7IoPgIa/q+bNA10fr3BjBGV4gAOrQg5N1
nfKVibqqz+D55ysKr/OzKMNqwHGI7thxDrRrnunvYaX494Im8GjbXWT12t1nsBf7
GsUb8goXX0tfFPAVgr7LcFzcFGla6pzxpIpoGBiVmqZmQEMbRWsvdT2omzRGvG/z
twHlHNI8nM07IVT5cJ06FzcZJlcMTh0lxGuSqQweBVgJWEvy3dpdBTsz+a8D9Gbj
m7qNTT8WUzsfmPVjCyz+SLyuLLYHZ8HPB+SHs1KWIvXXZdUBgj3jR3F9yzv55bfw
72Y58hbb8gT8iKUEMR+6UPsHOTOlZ2sP7x5DvW1iM9zKO9DGqu1H2rLETZ1Yz5VR
HC38AXRsx8WX0Ez0N0uiLDNZEESZJAqYoP76IRx+q8dg8//lbKoX8u2Pk8qGqAmP
IiWhIa+FXSfJnwtJDGneuwJQZ/VRr1QixySFfQzPnhk7G0+UJGzCmqMJ9BoTddCe
UxscU5ogb1//OXeZ++eK7IG+azLVCQYQp0o4KQJGtMELWZOJI2nYdNuV9tlJl/Pi
SDXpn4IOt2Zm0INLEnEURBMgs6OZds6hMRQGa6vD0/6aHPfzGzC5aq/N22rbDPJ4
K60lv/LsVErlcepEl6SPSFsC1JxTsGGmAwJZUTmku8gD5PunwqIUNupNRdbKlStE
GROClsV4GQHbQdhANm5dBQKOEF3KAlPm+I6v6wfCqLmYggHgL+hjro3LCHTcTiMm
MJbZg5wuwMfldQ85fSAdBhOH55xb93oEXyd/yBCONynxucxCsBq1NohoA9cR6gwD
dyppB4WwA3c3xgCX7sK6goJ5izYi+MONm7TMp017UBhUOT9qKtb6WdiuwoBTK2ie
6ovS9nfe2cO0cgXjJaK7HxI0dR4rSlxe3o2qHeOb82Q2NYPGQ1VF/fE3wY+VWkNm
71YSbvLPmsFCzBzQsqoCMH8L0oqMflfTaucLY4lTFXkGs/YKq5mKM5aOS7jLeg3D
j8Eq9hsFVLIX2rOKjkiXf/wyUgNVEp+PAoj/HIV0eG+pllHuKXsFrB5G7MtIsI7h
4tqrVeUkK/gB7GSmUrtvNiolpFoeA99aS03bvjgdV7bGgEnRjC5wOJUezmiY4L1I
YLuyKtMBmxUkUNRH6yU26X/bipfZeLkoyquAldYdF2tNR2mCiKSybzKkjuMYeeYu
T6KrO349cJ3PurYCSbwx9oLdeFJx5RKm0WY6DqvRXnOzPdibBuuoa8BRDDwGJ/g2
jjMxCpzSGDqUHtjUiLzykhoSoUrFiO3p1I1+u+U2pHyufiwi1lF0Zy6sACzy6Hq9
YVcVxY2FEhtC4vWWP9MDhy8sw2slUvoLmaryir4R6/RTrGAJ4Gan3IW0KQdzEdz2
GjLwcIXY4zl0GEDkFKC3JNXTlpYS9WhW3FCQKb51gCh/sAkbQMgRjpmzsS/9dfcN
1ZGzESvottZ0VcKmS/VK63iYzETD/UabzVrhVPH+AML+TtuchVPbKnmzDk/quCOC
yMYLvhCXwPXBzVu7k3pWd1FEzftJWyz7P9DK2CgASqSqp9HYt/C7IqhfjxhBrky4
EnQCzEbDAuDfrcRkP/GauLOtNvxNEMbM3Dm0mAm2GT8Mv4QB1Ix2SgDMxx6Hmm9G
RG625fAgUnG0Igkmtb/LdkxKJIAp6BH1G0tyHPiezK7LrxrUpnLmOSZP7nlv5S1N
6TOeo8Uvqa6kaDI0qi8iOxSy1wWEJw6ABKH7pRF9F+eU4F95vWZlCUZ2R7u2E/Ux
Xi+tSwA4r9q56aQO5Gq2aPcMs0sLx5rq858ZjI2POjTTNdC0bvvanrPwi7NGA2pv
8kUfeC1PKRJN+qPUaezvLV/pIWWvIVDcxh7h46t7jZAy+t2XT3CkhHviDRJjtjVd
2DIfPe4D+tqaQJFupCqK8TXFFUpoorWEF3NwzN/Org/jXMbO9PkJ/8OUxMLv/YFR
8mrUyVfF+QopKEmSdZ+FGxPXP4C8G+ibIKf0U+rJBCU76+/rWmI9Fy3d/aIMPaVe
YdUARKX0FceWcDRQHMojHxWIAw+a7ktusVw1XIuu+9UE7S8uZb7Oisguhypzq10j
sLosfOwto7ESyo3BHvx+Ps98mtDZ7JTD35TY2tKd+McDks1Yk20JJ2UtFNCVgEkd
PAZMplAacXM5kJYckellKmmnBOu/GADBna+g8FWzAwSWllhVT/oqVRKfJuVuc4/t
jOWWAFCgmkRzhTTxMWicK6jXkERshCZMtNtgv0PC2yXp4whzEizgV5pZyHdAQerx
uxumiR/om5HUVVU0KGmdQj2sCIzImR/0OMCRT4yzwShzspAkpRZ9bfR6DzyQ1EXx
tJpsBCGpSgF95HqWYbS2FtA8BSPAADJdtvKtI8l+boDoLndTzAzYCBR+YqSrCKuJ
uwgxDH/Lz7hgRik4mAkADPP3r1oUsKf9UUgruJ8dATioEPDpoL6jPfYw0+qrFYxR
41bRus16VQ15yNyYDNkMxkWlEvORghqUItfFDOpU40D43lcisc5CpImwtiOQm6SE
0r2W3F08/tAXB87/Q46G3qRqablxmrxMk17TLd8dgo1qA8EKFCAxaz2i3JuyduyC
cteZ53tkkVAmnAsGxojRuxGTZuvOICRDe7cnTpDi0hTzEqc5bUex2uD6jUEhTQ8+
vZvfkBr95Dd0YBqT16f09h9SKr3Xzj2Ldb73vOj2+NL34yB1GgnAIU9FaJ+eVmnC
VrfjZTpCRh5mojNGJLqYeOjjWDAizK0I872YLgO2xsEl+UGPkB7C/pk2TJO/b4U9
YKV+J5YDyWW/t5J2cntYEvlY5ftMFqkt98YaBw+cahDJMGq157r1g6KYypMntzr3
Qmmr+QiMmnbA8c6V1k8s6pdfptrgDwaDuN/j1Cg7alHAVV5+7Oq7SukNn/ot3GTc
qkKYtEXMsbxfSAJC9UpL+n6MBNVdQWK9Ug3N2idWW/VC1Bky5SITVfY2QaJHgX6l
Gymz/8xbsxLjXsR/SDor4bUbRbfY5yOeaJ+mxh166CvfUYWapfSvNcPMKDfcchEF
I5D6OiZHy06bWA184ym4d4+hRJhubiFPIFb9mPiPIi9G7yFoRAvflaJZfUv3Nhrm
nKAA6n8a+UDZeW7S3lz11DzqIwB9FLx76Tjwhyv6H9rzQxESntKfow1wnPRUJVz4
0TXf7/tk228+zgIVHZ3furvGdqE5bJtGSHWrlN89b1gqq91jDn5NC+MWncpsspon
yZTT2iMBZcKJw7v2DGQn7Uukqy6oGccPzwq91ygPbHIROQyXwy/Cq2YfQdlEkIsx
dYlA6RvRYEaXJXxxDXJy3edUhlpqsMZpED+y4bZIPeXT7O3AeBMeD0y25PwcR2/6
c9ulMbdlthbPLMf69SeTmNy+r5q6z6Slrpxzf+iaW8aYpcJRbanK/er1BAD4DxiR
sLBtmfMdmnaM6Sq2CdN0ZPVvmw5lmbDp7BFCt35OlIUH/k6WQ+re1mKWNP8qpa9Q
gIrApcc0IVPiIT4rpSjsiTHmm81SqFxEd6Ym6EYVD/xE4fOatCwQUUalF5lYa1qg
RjmSkOrl1/hxZ08HUmOMKhJMlEbWfyX130XuUtEDVDkhcYsdPv0g6BcBwxsYmzgH
sgLj68xZ1lwx/Yv7so41lrl0+Tvh/juPG9QdWuNUSxDLZN4TBf6m9DYnXUO3fnQI
HQv/uGWmlNP2icC+vpNETX+BRZ6m2C96ypcEs6PV+aeha9i0VwdYkn6NN0wtBiKO
GmdARFGI4KXXyMkW+WcCRIFqoknd/qhA9UX7Vj8Y8i0OozaxFj43yFSOGNNRdkLL
OrKfPDDQiHhe8ZbHggrt5WeE/rYy5NbzidrzQ4pL4ZFEypMDdDbOMn9cf3N6SNmL
ZuSaP7KaU7ESmRxFtJMGBbnsUhn0ph1RmV/fuf70JwXXPzNoNnxl2N22Ef11nULw
TDZcMJc/uFxmyIvoND3nZwDBqymRyn6Ptzk+mFmKCYrl9Xk0gcm22KUhvp0DN3jj
0litabwyXwBC3uxpmiXyQdWo4KKQhHDfKSyPEj9yqdL4sZY+ucTWiRyLjDi65vZO
OxIrW5yo/1uxmo7qEIupNWpG4IDKntGEntUqOvZ4H6COqIfTHP4YkHoX9RBOy72O
nK9fTdzv1durYbHp+eYqZplrjb9nLoNPrPyK6cIkXTVMO8SBJkVZV+0OasoY/c+G
cqOTI7FpcuOPIm5CN4jAvXPiH/NbcF2ZAMWoRWBpPiQywrVh6dBauFTZl1lyqU2W
m2prSXH226HMMLsD39bMHl2kFwCtFlgfmcfMWYWlwzMqlosxld3j48tuECB0UqAJ
XM63kpAaHcl126ICtrx+YvlLTYqBRCZhXefi35c+u+U6NHo7dDJp5rsxqW3EnOtF
9sf+hAW7DsGJgN1YooQCNu2X49+0O5drBT/vIswDhvwDLfNY5Q9C+zlaDflbD5x4
oqDxrsCmYXPVUmyheyCslZdDlD1rh7vynXjnUn9HAdsTAQ1nF8pcZkCJM5w0gqol
q1T6g6LHGHgWnj8hoJkrWJ8t4sJc4Sox7eXxHCK+EdpNLprXSsfxnxikR3zBsqYb
tnPBOcxoqfappqo0wVMKk57185IDS3ghdfZDiiTecBuLYLNTOuIomFv/j98U447Y
mzI1TiBRmepA8KS1gBQe+zaxTXt6q5nhGDy+uqNBJL4mc3XhisjW26W4rL58nSLI
yxuvLsJfa5CEVPWKaF9OdMXbAR+vS7GwjwdXOGn2M6YNIHLbuoKX9C78PBTxfSu+
Z/8PKeP+PGJdeCdIQbYPO4XnjAwxn/Zv2nb32krOVKPz2AGVzIXNk3yQRBCHT4OD
DSgvHcoRIoNqWn4IpahkD63KXaTCmS+df6YdPRGZjIF8qezAzu6hoi4BLYpfdmUs
MuMFZd0uwvhb9ejW6/u0P5p/gne7GpOaQI4Pz4j0gx+xEJMrceASwz1DZLTJKh33
gjSTBo2gZfgUwFMQameS62M5+3z5mdalVCaBosLfokj2U0eJ2qmlIQZVLJqw2j0J
7TawetUGwuzZmuaPiY7QDuGkOU2C5Ap3A31nEWsIBCYIgwbiStycL7olEVItsrSf
WEKN9nuwgiGQ5QRh5R36Q+pI5bXmBnyKuguVSQrDdu6xaXc5XCVktGEfoZkcgb+o
fl6cLyjvOa643r5bWFr212Dwwy21ejivIAlDaTz2v3qwgJh+uk9BR12cPlya1Thw
/B8DvkoBb65FfLleFo0bW2vzLZJESRS7x008E9MjVfSsZb2L1y1aiodfsOIwi4uZ
JhkFCkhVL9QTWKOQ8aPxdGQeh7Cxb/vCB/YWOk9qLSjYT8zHUNPvMj05M/08fB4y
BNZMF/AKyVmLvxaESk+TaW8ovI64z4I14hwR1B0dP54AsOFldgZyFkx9XLEOmRMY
hoeXLm6MCHDjiTBn/sR3E7rvmO60aw16SkyPj7DngXfyDzxvs6ALcf+4/a9Nshak
YZjdS0erlp5FwBUGh2iBVQQbL5F1zYw6Yqk8D3EL5cl4qMqTvJYLWT9csVvsh2U/
bA/pUFpsVpWDR6dPiztzUQVWvhFJBPBxSuvVGJfIGWST8dP7xFQXswhDR1BlMXkx
phocKVxQ+siC1AP/m7vrzocFa+WmmhAyECi8hmX4hE6elho1y+82DTRQANCRjO46
Is+TXMhGKWsuMxECONsvEouyG5pXeoEKujSn1PtjM+Q9Y+K8VTQeYsKngZf9WQJ4
Hs7y64O8DJiKRMZMCe5xnqoyfmLTEscOib2ZP6ocxiih/KS70Zbw7iUGuvoQRLsW
dK0e4D59UertzAoduTEitmbB5VGqXOGLZYBmYrTgjCyDnzD6AVf9j4ueWzscWwKh
u91DrMXo7k7kUPe2RYJqzUKCnkBIjGy/difo/wF2+B9eMug8WgzI1ogN4V8nrrM/
niZSr1agbTHVuIKzJgcJBD8iomrB7oADXJ5gWT1B/yzK00VcCieDcWSyIPoJCZj5
xmieONBMDAOv5HwAcbcKetwafB5hvWAVzLWHzftJkB0mS+0dTwOBVq/PeZBzGTGs
UDa+wqYmIzsg+kCZU+HFOY9kuQ1vpFJXggF3YlmtdY6JgC8VZrDK/cPndsTqJ/e8
gXy2ug+rB6w72sWQbOc3KGUMjgJb9P3dS1f501r3Ou9UqJdpdbmKThJ3t9UEvchC
6WYEwsE5uLrPos6NMMEXjIwobF58Iq+dnkHia5sPKqEP1G+AlIAKRnt6KOCGe36U
7fdG+hCCrJdr8k9jhJZIKFKCGAZhF3wh0QfrWU46LZtaEi74D9x8xc95qIFUg+ed
QnuruAMZIazSNc4MvkBPvL/y5Ma0urO88ZsYhuQd1AXGFZ5HmbAN83yZ56FNjLvT
gs5YtLIsg5AGapaQAdeQqvPuk3zgtDhhHKHpWNnblw7KTBDITynBewESoSgYLGaC
MJWbn+Ee+0m7hZwyyntJeMofMhXX5gSVzmAmLezTyk5a3Jqti0T+N+Igpr11j2ws
XZdKsgEA96cP3zG88nsKDs47Vhe49WVrh9iKXSaU8TG62HFpCX/lTQrJyMz+/Ctw
vK7teOehwyN/J3TAmtB/FcGwLRyBem+CvZS5yIuWSdVLS2//bJaNatGKRmBFa8M5
bC/oh6f9Vq+0jGzmgQDnur9hPYKRn5aKddTut1G7TBcFMBVqY7Q6AwAVGolCKmH4
LuZJBiLZGHooWgxm2UJAggGMLThrUc5XSd7BTXjzA089ZUndGy1HRFNArwcUNCgn
ycY3/By1K9zMdC8ias3S1+jAAmk7UAIkJl39mObzSkG4pz3UEMZNPeqcg5IAc93J
TcHLg1EgHk/+fxB5pHPcjLY3td40vkaioFZc4GcOqIUzrn5T1Tfe7Qq6t6DuO/4h
jBy0aPXCvdNp913v5MZhZgFz7+ExoK6YmfJuJTp3AFaUcn9wgHlpQX4eK1vnfjO/
CMs0rfKm3+99I6HjDjCO13h/WONecddqlEc1UncH36rGm/2ddhm2MVxVqAgcXM93
IxmYNAFGhCVrdjO5amCi3+Y9RLps/K+V6gLMVfGmMejNOO+6gl8P+vty0woxtESV
1L8f6HxUYygSUYxe2J+WELb+lkKhygHlQdvcANmid6ps0xl0omo0czAG/7W2xQsB
AcW8++41TQX/jB2KFQYnsqgR7ko2cA9D8xvIAZWqhxMmib70mMnrTBAtaVvbBXQ/
tcm2QVJCHbwJb1vHwwIXwzmSWlMKkbSsJBT6pJ+FsptVfI6o2YG82y2AoAClaND0
pdaQWieBYOyIssYW5gJXjhcE1gq7JVHyII0PULBngZchE40f2CVFcBHo0GUTviQC
rfjUFX8lz92q6mUGtrxtz4BewLa+8FvBY3diPeCwmN21ymqGnoeVA1tPnc+nqcHv
3RKxFR5+z5kKt9iEzb7Z0AQbdH8RUO2XwX2YPs/c3Nbu096Bp0NRzcDh5BBHguq6
9vKYiJHnfoaY4aMFAkJfAF34MRgt8ynmIT96dFMHlcAHMp354c4gsvEr6cBDF5Mk
dd5jbrCOIxggEAtpn1NCVSLr+9Q7IaFgu1q1p0zh/PG4EXSyoDbV73clP/JmaSg3
07BUfdMPltjNpAK3gW795OitM7oQ7kj4+QKJettDz/0lli4r+Ts7nwr9z3v5Qgeg
UH/F0D3JWEsYS97Wh641W8w+rbkqjeS0wFXbyuYKms4erx23iJUz3mY7iCN56fhU
WxOMrLEST3bM9kLgFyR/37dupHKouHE6KQU2QxvkIVPPBul3hCkztvel3pKqjkKa
vxSxkzqj/niJQEJgrX+a8T5+F8KDRWGvvEetq4uTUaydZqgwfy7XJZXVA2x5g//y
uSuk1ynhFJxRWHo4E7jLFLtTvA6hDZCEo7DLzgALdD1vLCpyo/SskOC6M0i7+9i5
k0MzJXh5R9e4rMarnTV0Pdd4/kbsj8GXTqFzo7uvlybkegOiTnckgPzla3qcE9Rd
TOfHbC7jXXz6njEDLSXlwFabtXYJaTFdtAul5LYPRhGtB5EqqyzcAWEbdsGO/p4X
P2fsa7GVPRZWsqYVW+cRTc6hbINTDEQ3pwKqR9byELiyOqwMON4I63v5CA2RTaXU
PsFliY5MWU6ut13qFhfJBWoNe8ZvPiC9S+rQugbwRwBp9TtxkhpV5xahIvMcPhFd
Af3yWXa67la218LUzgYieCFTIKg47ImnKNNLt1bNKnQIGmABTBr3AguR6JKgh9aq
MOzkP6sVVbaLPla6taQiQH1STCLB/NHKsFcWEWDWI5ZZB2LTYdBCZ8jAuOh3/zN0
KZ3K2xnBh57mteu5T1yUftPGlitV0D9bojywWh2BbunYYqFZ0BUSYXJUgGXoWFkH
LCTM+WQWcmYAq/Rq1JHPXTc08WCuNWDaNplllE2QDiWk2KEAYMuqGSSnPR43iH19
YwCy46hOAfSTbtVaqUDuysM5uqMk9CHLGLg5Gt8Sq+UkgznNWS+hN76cQPM8EWIj
KoTn4G7TLktGiZfqswblpQumdzyahreXOpax4LtnXLk+pp2GgsFObmEGdojdYwSs
x5xffew6tofmGklNRH5gIdxtvDijn8lC5J1ucczAvQqBEO45TgikNVZWpCtBoT3Q
hPZrimCm1nlyOQ8H8oBMbO7kfvlApae8Ft1omjnwtrZsJc5I6Wp3a+2XP2zktmAp
QP5q0BJUku2nFKW3wWFSqwOt7MD0n2Btnv58IunmRcQI/Tk9hmYW9Qj9iMK4ux8d
ZbOmaNH524aiFbkqGMZDTAQamErhz1Y7AAU04jnsyb99h1swWXDP8K5XYhPOSrTk
6NmecDssiRilqfL8IGFgA0/WRPYy+s8nluIX5ylbJY9YOWVJ09YnQq23SE3dSXzB
xBSzcYJYaPIkN6Pf0JPEAugu5axWZGF15c0r1OfAjRJmAeZp3TYSU5tT+YuEnfPK
EIwWOk0trqvYnzGVSXhNm17BAizuKHtRwzlDBHVvyjspK5/LLx0RoxlxKkuzgUxL
fn3LFz4fvH6vyiI82xAD2u8XVILJc8GuqOASZuPyzqEVV796KksOhlkhgnqN7jmM
1v5W9wtPm52bCc63pjIQfcdYwMYXUUoNhesDGzUvnzEAkVE8v11agAAAcLESz7l/
5LKXKYJG7PjRXRHEARJBHDKoed+o7t2kZh1es2PDue1UYZFLAeBoySL48dT1F1uM
Un2+LpdKWq4T0cI4SxqmAzf0nQZyxizhtB4OnEuFB4mPliNHF2pW9diy5dUfR3Kd
RkkkWKKvhGr/nbyTmJ5wxKeSN0e378EkPKsMUO3XF62tZrtpzUPbUGGqaetBWyKM
F4EFqf5EnZTGiCHBXsll0ku/XcC3SJ7C3KaSpxK4pI02LweT/oW/C7/F9jqgpHeE
Lv+DIZqTPM9b1YpeQP74Wxxbff+jouKdT4b/JUZ7OKhS2ajTlCdl5kK7yytdTTfA
Bh7svTptjUSNBx5PjSZXJFet/29x+s0R4jBYz4aVikRveQQAIlw36ZBXSbRxuqc4
HlBEKdVjCr5yjReBcDqFx+b+xM9D4i/jyNeM5vsX/bYaxXMR4zNPnZYISMYUMA9U
GctCkfCtlcBCIFYudiX5wKGyZR1psLdo5WT5Xkz3gMvzZorYaYKHjNCnEHOsvyNM
/TGbqKjiE/j+KxwTqV6J2NJCPtzSsI7LQAeYLD05HRwegW/l6RNlgxyFt6y7DwIP
Drs24OoXhYSKBwEfLoQhVcb8tO62bQLTBolEFTDicjwQQw9nyEPAvN9Fsb+2LMq+
L5rn3lsuJ/nhZ4/ik80/WHpypi8OlRQVg/fTVzfXVUKXsdmYFBwptuFtZ3abUpqx
8M5fpE18igJYfe3fdlx105Hn05TH8v7mm8NBEnVyg9KMwob8MHDWZd7n+k3p7gth
JybLC2W+2eFSGO45JLXJqDnehaGZfSqrZAgz3anotPrsV0iAY5+yu5q7lu1Su9Vb
i1Pm28XdDVgF7QQ6ieGCRxQImDnIL7ZpGEh5zFKrkx4NTn3c0tlorcIsVATPo4H4
QyPoOYlhiqEs014cplH+W5vkgvedZOkL1VD2ysbWirCTHjdKs55NeKgTzK4FSfoR
fdLPG4/MtMlaiqljxO8L+tdNHmmAw43IfAB52Cw5gYyvYemxlSycR7Xn649MH+x5
Oh8DcDdS73td2evXfmqypqvBf/0rjdRch69UYj75ZbWKbfd92feAgL/UGDQou1GQ
d5nUi3PUXW2KQBvU3iMoWZvlUHmvom/v+yupRdjgcUQXK2uZF88slWnjcUdG+Z2h
iQ0A6GbqIYpm4bQF1VAG7MFFAya7/a20X6cGaBgGEZOaEl7envNy+wrlzj5ORRd6
CBu+ax+FYc+FUz59dzFfJuyCxaOsKUHphm6izr4ceGObhcm6/BJ5SmAPSAJpaQsq
1sWHRpxKrQSEnd87cUiFHffy8iQIQXGYIVPpwfiOBAldbu3gXFGfOxqGFoCGKaJV
oFYMXSTikMd+lUUxJ81bYXBwOnuNqpEUot2d42oCfv3gKC/l4p610feb/mlc7e2n
Vfx5M6qMbVv6RYiOG7dHo738d/72MXjlNqK8bWAsQr598wM1ywq5+S8KS8VSZqs9
Bl+r0MTXtXs0ugRG3hSRLHOMppD2kcSMTx39cAqaQ5uZ9H3R0BZF8HSGeFTTTN28
HR1NfC2197HwMjWNIrMZkVuN27WDlDMocYnlpy7weDlynoIZGRcKauFYpNwYl+4b
j7qngibnmCbPeKI8YAI52x4aUhkPVa2eomx3gCHdwk3i/+DnSzLUquo8f2vF2HBx
5PIOeJLJi+m1ll/cYBkOKusFiaImrkqn1P9ykWtLIIWPZGA3tSA/ZU4t9q3XDuit
vmUYSi6kA23F5iQKuNOwuHeUOijolGnmjC3NgXvEPtjwbKwvnpdON6HUcOAAC2G6
/NHJ88v6S+BPOqbQhAm0ejOX11W0BLSW0gM2iHtxSH1ajSVnu6HNw286zmHh7DB8
YTAwUCuCnEBUcYLHcvnW1XXnPj7hTZ1bLhkh8W6+Ys/7Dx8tb4sy85u8P+b6gfvN
gy6xSiQn2Dy9CxLr8xjXy+pUP5UO8vkEA6+UHtcU+FVQiCl0r+AKL6jBqRVpUD3+
NDdg43HH2AhEr39dw1P5ldQRP/O01yjLEVD1imGmsyNnIRYlNKX1cQWyptFojIqN
0UEGfwb6x6wN33DOMwfeJ/L+C70LAHd8Zuk61PXmoPgc8NV6jyVzlPlB25t/3I5f
GWzJV6Hqg6vhUtv9NMFO9e+HeI58XaqEpAvhhrmbUx8Z6zwAWBDYfB2/A32O31EX
aVbxw/xvPRa4CnR4dAsUA3B6qpXn7EsX8D4Igs4VGXjcMy5i8rgmRu3Fk2grmW0M
+6kzsXWKSCuZwMMnp5LMPY7nScAmO3I33Yfl4EPPtx91kuUXLK+V5t9Ex6UXgAdh
91EMIcrM+JGGlsla9SL9cQQz/nuG6jC95TApMc54jBT6oXxjjqvlBa/1I9GzqhPe
1RHFBSj1AoqM/wVAO19ftZ00r0M5na3FhdRBQHKVIQMFKfvoNR+egLJmbcqFkKnO
0IZ6nozR1auFzAdYlUoO+YYLBcH+daHsfWqfDzWZMSGxQTVOEU6GjJf22/OykxIx
EDO38TtkFEOxBo+WZH9hKuEydzZYkO/ilFylEqC/Td79zsPduerI8fXhPzwNamrp
9Q5J+Z0hF33YlIvgavF8U81LWVLcbb8jhXNbSMNMaOf83hBRsBtW4ed+FxoG08ZF
CM9cp4VVMLsGvujrbJD8WJYbna8DaOSLAlpiB/rd3e6VkVsxpsadxvG+icR+bNsp
yNhK5yMymAfkL4Z8AbepKv7LrthKcYB0X2DC8QdXDRqWNGNrhqG7djE7OO1/KDHd
hUgH/u4yg2shbsyCpL6XmkcNRudwT0EHYX+KnVGuuUArYacxbnaugeLVcN2eBYHj
seJ9jc/A+T//6N6aNCRMmXDxqn5wNTNqqT8lv9uZRhU5nPVgdzEps2T7jci4TqCA
Gmn0MRINFqcKVKjYyeldb6SYc6AmbwNjcYUkokteuYp2HgeAcVedC+e4esPlt78g
hQiQgthZt7smRWobBzCNGL77UQURLdxaf5XrUCutJP2xGqjaB1ifNIZVzr6/+2Ao
UwFCXqDgyvkKNR4mUn2JAnEMW1UYxkgo6yYjfrVYTHpOPrRBOKAHemAf0ygB52G3
wxT3UC6qOIfW0K6Nd8/0EJbthHr6zTYiQVCELp34xKa07bJZWfo0oyZ3AGVktjM4
UywT0XNdLt8VG2oxagTkJl1N9quOm341p+d1ElZ/aCtX5+qMPjwpOE30OLnG7HGy
DYo+u16jds+RmKGnLuOTiHHCmQ66kJe5iiOoYl4qPYILay2BIQIdiXAPqeJOLWXo
POic9omMcLDtHQn7yLEntMMeDgkAVZYG4hQqnuhUMt9tlzBeBob/G6PZJyUBsSRm
xrs7JMkUyOT9FcVRdW72bbEnhUYj20qos8A3wAmKQ66Mjc8NUzJf55fekDjWuNsO
jEZOYwTjelpsv2WTuITQA9qmZv3I2r6veyy3ks3Okk83w/n0W7CDDVAi+5Mz2+LE
k3aU1k7yUzpfTj3sNslm0w/fVOUMB6CmqqVkwK2ElAQjs8tYR+V7WfsmG2ZCmlWb
sKBujqtuU66qwWqcwAo2tRaqVKQENnq4jnCFBkmv7kB4Ns/HmP7s62ArEQu1rtJq
o4c60oT9WJ6shDG/WcrfJxG6XEhi64Je1eBWk6hceoGgqm/ZaiVBVPss0dZ/wHtX
4k8G0eKy/LKTq0lG1Cx9HOPcAu1S8I3mWNY7l3axlgjXccPALFYbcpQJ79f3sQdN
ZxMDyJ8YfMBn9XHv2PGEATzmeNf3PNkjcxqKvmZBoDTOKjMC3a9q1+TPsNXsrY7i
jpP1OI7FJEKZb8yeEGb6iYoiyiGq9wke5LwLp4HZt9K3WomU8swRXc4J48lF1BW5
1eBGtVYoqjsbuhBl0zcPaI71xQe9S23QNbwWSJ8um1JNu050pj72ojtDvQEhCW7K
jQXKt4wEEsvha4O9ePwWc8ZN2ZQSFiDuGZkMe0bQcsHXCTMGamUUKP60AA8fBiUt
nU210SlSS3JNeEvz8lmn7IVx0lSj1XKDVZDPg72nw20Vy3uOW+1k4cAdDZD4yjl3
2H/asFNC9CUY39niVNPu9HD8EnqFYFsAslAvCrfmWJciY0kRVZw2VbLpJnlnixcO
GXirWZRO571EJA1WHyagjrpJsKN+I1MyFz6IvnLE1jNq8k0R9VoiEh4meHAQcikU
ASgJgyrsKvBYEvevAJ2y98BHzoL6FOz6vOZONcnE7sv86cLhqDDUgoekFGrIEOFh
rpUT+OdUFSmjEkww0hiX1T5yyvcmA4ujEYASCGpY0lG8aV70rlnQCMw2uD0cK5d5
mYPGT2YpkDvtP2XhUDdfvR9pMO2JKF+9WTvg31vVny1wou0ltFVGQ1s733YrOx+r
dX4p3aGFtuCkl2thel4GWRoJhcHAT2AsiG/vuBwZF3SXfPYtpvt+OK98JPr307Lv
W63FaSl27KzpQDs50lwIzzRsWusoIJjpb2ljsooN8B3Nd2jr3Vw7cEsh+21e9G9I
S4SWJvUM1Uh1JgZlN0FPUK+xUVktE6FSziH+lCVfNZpmnsXY3I0OMbbKulS0tkp0
e7c8cMi2VRGeV4T24tal076PoXSk5xtfpWhVvmf6o7UV1dp7FOTrsCZ39zmTBM2n
6aCf2udip6ODGJLM+ehbF3I+UQEgciy+Y4+tVpq4lldr8TlJDY+aV3Mhe6G1KNBj
apXFp1mR86XnZU+atDa7yWhIjNyA86vNZQ1ZOCQJMaxpRB2e2VI5GbJxFvItgyzs
GgrmFbjp+CZIaAqgrMTEG22TNZL2ShLIHRPX6+YNufUonuVfz/W6v1K+xUHlfnOv
iib+9uQ9jSE+oe9SNrTbsXlDL0DqXX6P4diAZ/fWvpTjEgREku7hsgmEDkhB1MRP
RGd6TQVS2F7aqTEjcTxJbgsFw4Ep51XlWM3u6K39kI8HAesM87+UAEv977DX9pAr
YDeOLpFJpk07+K1JpJlQZRoduPbV39zs4HEXkZ12ozd4OY9yW7YytQIqPUACB9a0
X8vNty4QgunIJPnOYn6Uj3nodIxsSSROaXghyTx3MBP4HLfwpIud18tTj79wdY31
jAnsexSnAgaEO/1OUA78Wz+irleaXAmfXp1boG5N7Vpzt7Cvcqsvnrw0hhlFJxx1
lGnV8MIVyS/Eie8mNYM3r1JGwbLoCIeBvIvqAzuRHYrgjHMG7XjVV9Mnc3iBBHP1
bOEwV4+yCYJIPpybiHnp8ZKTaQhzUkNllgX2WxOsxjDC0Y9cjwP2hUZvcjfaS6DN
kHxjn+efeDrEDLtQO5Obgu3AraqztyF0S2tPIe/MxrPpcIpd7FZv+2V39Qhu0lAy
xIRprCNEVwd6qgu69xTy4tLsGjD52ydtyp2FJ5htEw3Ydwijg8CJ7NeNCYx54TM3
LW8Ytpyu1JqgXsl24clux3ng0OSQ7feeNVjmUSLjtlrhIEncU2qfTOuMSitIBpM6
W/Ui0vHj4mYBzs0GDtJ2KvvAG0p36EyI2T3v6RxLwlsIOoWGzxwHTaQu0lINUWHm
L8spNsQsXMTbbdH+i6Sgd3egH+7OAUM44qVGMhVUivHAVasQZX/5mpy/wN3Kx16V
WjvMXTXVxVpLuShdNpKVrtmU7F6wcHzvmK9wFm2XeXzp4+EQkZM4SVl2pVHl98+v
NIc/MjSZYNu8d0i5D1h272iAqJTleyxKqaB8rdPdPWLpDTVBbLkGDb9bSFPsSxQm
xLhpLz0iHVtPrq+QkAralYAYgl73ixRJ/bpQEqpWPl8RVEfMARwa+4f80PnY75/D
I6yZ4lJtjT548CUsc5ELwQ0E8TnjnnXzEfQhpDc8hDGzkUroQ59WiEzXFQQck/CU
svv1tTCGWGOr6VUUjl/VQPAQ1wzfLZHI4xLKgYDUoJv7PYs8rjeHJjNx2bF0x7QB
s84ZBlh3QMoiw7iOQDh8YUTWaO4nD5kuoF4RUDvrU0BrEC1FBm4oXrWEjkV7ECaa
MHxcD5ti/BdQbDnnWKY8PirCsC8WWkq21K5h1NstaoGwkEB75ns0kVitIkmmgfAw
kc4mz5LI5qPvXCa7oA3gXC3mCKvtkKcwfdhDio1IcXSHN/jpi/Ah8PHRbX8PZvZq
8K3Y/lHt8K5VmAplNW/RL/bgVB/1jfnj5FZ4Tzpj5NHwAkKXnsdKxpcpD2xeR9aN
rBzR4wmhxSM+Lhx/p/rs6bd4LSscg/xgbU0wtU0bpz1POxVy4uyQ5qjGb51mJagr
XIK71siRe48b7uy9yls99rYfIJssEAOttacpc0FV3ROz5eNBaiqSEnUzrEtP7JY5
lMeH+tHS5vCBKLtdr8wMQU0CYI/nccFPhc7iK19tna6FlsqSFh02lQaqhu6/VdYB
MbDG5mCdFmoMTFQeoI1ckUA8QvWJp6lfONKykUSIraOEMDzPjuUVIEuc5fPTApc0
ZxIiyyBRDibrdYH5oFSwHc6q3oc5aryDNSKlF/ZjS4UkeoE3mRZkwsWn/glvJdNC
dNblO7xYF6dakTpLEoQyiF1vxUXp0p2isSkl+jFv1kF15Hn/wI3WOnV7xBO4TRJN
Sl/ofbPwDKAlX9/FwT0mg4oIe47AUJeA9OvGWM9j7zFr4fnkzuNHmGv0nntW0Iek
TjH8TjGy+UkNvvhCpzGoEqoPR0N5FVfXZbUDcg5o0R3/5iahOKOBneAXsRW2VOfP
YIJPUQ9bji5z49ZZbm3rfW5D+YpT084X4g72L+AuX50tYG19CpssIaPFJur1gU3h
Kt9kSVj1DHLl7itTvERdZFhhMbk6N9KVNj6u5mBn6miRWA+utib8gLklKTM/QZI6
WOG/yv0BRfeMh/HRikPhjyL3X31G8+7i3aQxelvWXaNelLgdumw6oGUXDGd8Br3/
heEcYtzaZIMWQyKPLD96ttAMiB36qNUX122Vs8sPQWYhviB7qEXHN513g5k/biq/
ex9doBpXLF3id7VrrVPg86c3YBoJfzfVBCqMitjwb7bIzZjpqFkRqZYQ+ZZWCPsX
Gzag2UE3oxzatVKRsV7dBukAW4lTIFlIM/gyfjEJovOzFK2FX1uOxMd5JPiPhCax
C7IuO5RPomjObR67m1hCJn6ybgmV92ANxGLxqWIsJpHTcFI6eiw9nP4IB7gTMQiz
n12glJp2dOnK0eZAYmlxKfwYR9jrgaZHvNJe6aw1RgB+SS+jECyb9jlg9SFoC+jr
3LUkTR9lod4lN34DKkcFtJml6f1akcZO8O7c9QEf+74nvoWre27wMjvUQnMbQDUe
x//DaboruPZ+yW8kFXbO5b5AEusRFP7kKgufqMiztofXKKWEpDLw/Dn2VowzQgnM
umUDMGWRIOvl/qb6QEIJKkxNMty77jd1OtLcGLWHUdix5KK29DWyVLmaxzhQseGW
rS5aNnQhTi7K4ey9Es4wPLhHQYp3avQjl5fPAXUjaWqhIsFVFZ/Q87wtTdgshHgw
txjaQ5BQ26/vadXbL6pF5UJ4NiINYuED8KcUloFGcAm+VTX16YOvrP0DwPaYQkzc
3usRbW14NiIbjlfM4rhrqdAaMr3TqzKZ5N0pniJI3RtsRcjrZqRR/LrZZEfVhVdr
5MvX4ZLhmEEWAgraTNlS8lK3X/bT/vyqfEwjnQFpJ5z2Krvjm5Dp8ZscBip+ZmfT
tcxL8Uec8grs58GoULyAJE+iA7VXg8Ea9Mv3Fue+Z3v0OV8iE/BkdqmCZRT55qKJ
F9gP88PoJjVaZn3jRprCpEjc6/0LbMIlctjIHt8JXF+ylUBUFXirAnl0KdHEZnDc
/KyivwDgFv0YWUMhJdZ/cJbGOiTmNTBtG4WmFw2ZlTbJmP8pr7984bMzW8AfGeQj
FIPlgbSvBMaOdrolobQ3lOis5nZdy3Sl/yLLrtyMM1gvXCFzkBNyNxdqeuJYuJWW
hXoAcFdmBmwgvEgu06C4T937HDLEsBoJMoHw5PGVaTYMBkMQxJ6rXnIHPdEN5ovy
GK4Tg6NafqqzNp/v05X1fkOgvb7+tEYWWMN1+kBNF69kSzVVKyROvwuF6ZKkB5yr
foC6hujNRlbbDcyzYnsbspLN2TMK10fbpcLMc8n0tiVkb3cECuRJfKisHD/3p+PL
H1TNShXL+1D3qmTanws2/DQc0twmFZdtZqFGni8z8RBpN32XwCRzuKLe0Xg6iZP4
rKhlwq0Oggn2MYPzAUPwOATNZgihTLkvsVIwCGXEZBWQIDjIID4OoGCEpRmxOE/o
Rw5zwDQB19T6X6PdPPViEVIQcGvMzGA88u0KXI9bzRJSijSl01Dfl8vhu4crwXE7
QuEaq5PlwO46KGOSMd2sQD9LwwKU+3GSHSz4gbQyWxXHaNlOse1SKBcyGSuOJrdD
ZUPr8fmp5fX/v/T7E9fFVK0u9/flck0wKF+KUU4kB3wOzk1bUxKQP4C6mIGm+cjY
QxUjxQO5wD4oglzOkoVcjrG1wn/rXrp0ZTOLqLxkEOA9rhfoITR48psIIwCJGm7Z
a531Uo7mNS9d4lsi4/17xQaRM8Ksm706Pk1tjmM8Y9GOQV9KRMWjF5VSFGUez10H
KNXhhziKepB2T6BJLroeInMWjCmkPi/ecmRdRCqUuqahYhde7cUVuElyd3tMq9m2
XoTy6J8QnqFaaqqJTIzgG9ogdV/CMAlLMJCBx19tEDq7eqkgLLmytqFYoykarDNQ
7BEqdaJ4G0TppeLt1wfz6iw5uR/4qYYBN3bEp0ZGmoyro2l/qb0tj42Oi+1brBtx
NHpTdL+w3ypVDXjWTRbfgAWzt33S4HvloWuZ//n6MsYNOQ9x1o5Msp9sHp0TYNXA
N0Zt3yvYXrHPoB/av1eNZqAVCenmIZjOI1BSaeoDSoGo3y9RSpEe9GNlaYXakANI
XAY2q/yITN0RLVhMcsPjj3GEayW6utZEPY0w+wWUoPSc6queSHaugx4XsdA4ms2B
VddRYEtUgXvHjUDxZjS10ZdBRaNcO46CFdaxc2LG7Tn923sIyEQn5gvxW8dMih3F
3HrYT6MRWQJWIXe2U3Kr37seR0+MwydfzbP+JkX4lNR1tf8gxN37qSlTAe7MvTHW
9xBWGOEwrnMZda2PjLJTYDI4Gk+HZ6Z3Gpj4LNagXg77hIKWhk0qDrqphAoyR24U
2kWkh26IUb+67C2LydT7MzLKL98OWyNFBNhwSEWEdYw3rQqyt0H5Md/QCGBVUpl5
VO6Lx20k7sx4lJHoC1xEmvqPMR17QiA+3QeCEViOxDQRrIqjALLS7hkwmAyQrwY9
Nyk1rvJ+3FYOvbFV09haATP55YpRCqHZCyadkUJ+kV8M2son3hmiUBS2h6OX+8y3
GSTKrGrgx8uw0bgHRVGBkZw8bc79MTzhnusdKRIbJxfaUlWW1rdutgqkosfm1AB1
P9wMgNT0VUEHYRmCodFQZflAK7Lg0kneQqsEqJkzoGx7wxJyxuj+JeXIFzYO2Svy
Qn0OmHwcY+OO0bpSiYQ6gbwPsgHkQ2iukeyqWTNA+xX1LerLylfPVUmr5tHte5Q6
XPV9Pqil9PfEt7NPtsfv+fRr4rbaX7Fer1UkdDGvCwO0//al0hkrQB9QgUKOYphn
gaZs2zbTWEWrVRhK+CVTcVB+5wEUPnr7ZA8PzTRTmhWlbC0OB+lWX50dCFGm0/lI
iqXms0zy/SxWBOf6xZKlwBe7CcIrtH1nVGKoJit8s0ngC7K7mDzaDc4qJ7QN7CGS
r/crbFOCxkKdygGH9LLWKFMXiTncJPA+96LxZ5hkF+89/Fma5vk0hOjZzuHi4MGG
4iDqX3/3fe3IULuVqivuYeCN+XpHK3DSmusQhPn6it4Z//agTcFyz1+/QCeGa8Jd
GOIdJTlilJ1UNVV0CDWgpLAF9CqGadPojMe4eDxVH7ddujxzN0Du52Xl7mAa7Lg1
ABFin9QWWZAhvFFvX702J3iaD7aimgAo1isjsNurigi2gov+tbv0MOg4bXojfwx3
NwQIb5i3aNvcADx0yrApgOJYmgkJT7IOUWmWtgKFJWJKim3xQkX/EzRhRb6/NPDa
hgYZgYv47ID+BpFQ1t2Uo/gB0T636UP+cSMK914grjgfn9xMU1RPJYJBWM3Xb+Rm
lviln2KoIMeqGu0LIHS4E8mlZM66cHDmCMChVGvSp7fEeWuZBMCfpYkczQSqD6QQ
p/QTtv/DGAY7GTV6+0Mj/rn2eLGICiAzcRWDnczh0nmoMxgVnfDKY1KbH0aMKJFa
Tlqt9msEc5w9RWnCrTBu3O9oceGLtclYTkUUKF6QDJE477IaIMg1nwfok/Fae9Ua
o+saKLUKWKBaGS+yEAVhYNnB10TmDEkxeDJRiDEneypHF1JfpjFqs4xkJ+LFniYK
JTMJaGupYnAZXlXaOUzhQi7h17HIEz5rpZHs7Vb3BM6tnz2E88kiJNP4C7jd3rck
NMmnLTt0qQ5MddxtccPG8RwnGD9bdDVB4RRet03Ev/W/ABxWxAh89u9ttSgjGycL
8JD2hGRUV3qw34lo7ARGfhwGHhS3Wjt503C2ZngaZSotgeXuXbyKlAvUtq11No62
dwgdUxnlmiA0CaiTt/9QTFVy4tOeKl5GjPncghwhh2cZT2AjRdGDcnGOERAomrRY
nXWn+1P4ZPzxa960HQyUMjUxqZqPqE8pTQzenahyUjlpi2qIAIewSB7RMvOPAJNQ
a7gIH+33M/GhVJsyaxWvKDszCGqltXw4CGUsj/gD7x6viSQLMmt37S5N26pTb6yf
gWcQ0sDKdEjL281YIaJHRTDhO2OSXejiFDrgP9ayKit5aC8ZFEHLu/7LD7HUgJyL
UNxlcmJGqryJQJCRM8jDWK5DAviyvqbcObIGx/2mLaTm4VKzwzhYZeP0F1Faatqy
uoIbnhQhu2PzCBcE3RjnPS5SfKrozL+VuhPim8H8TR/HafxVKyKW4B1nHEmPQj9H
qK1j6tg9xotfcctITrswDT9x2n4o1LRyvgMgYUgrmNHdVYF41aUt0YdIKxfKKsbp
xN3boaySpc+9gcZKyfrc25uta8hsk9sOOTY6O+guErB3CupHOkaqgbdE9SDUS7Dw
rSRKT2bW3d0KUprOxxu44xpYQLEioAkFsykL/qlhQ8G8auLOK2VZRvKCb6SXYzi7
2Z1v4cXqWHZLhIGfW9YmtqDxAj5o/ClbGqO5YY9yVKckSQjsvFsZkHSSQBRVMcMy
hthfm1/gj4EETc/47p1F/F/lyEUPU0RCQ7x//6cU8LAy0ONaqQmKVocjy3q1Szrh
TjZYROCdq8QJ/jFXs4VZ14Arnipcy1rqkE+VPdMtHqwfhokmxJ+v5ZLvKtkkG957
J2+Z4mjKrAWdaJ9NGRjfGmd+cbDQujD1GsIAfDKMFsTF5uUttldkpkLAA4eYBSE9
woEiAuV1L37pkQUqiD0bphSWdN66DfzjQ0Wi8IITbov5/zvt4lVoRnOP7R1QNeBT
MiHwio/nfiA6qxEKqG2DRoh2c5u0b360S24+or7VDQa0Z3K08pr8/xrFsGUnJzQD
hhUG0f98Tpb0EoEJcyFV/X3W7lHqGHjFSzgHUFjwIsEWb2J7vBpewevaxhgmE28t
VP5szoXGTeq/MYN+N0H3Elk/SMspLuXaR5QdXmLIs4F+f/JbL6mA5LV32kl0RXO4
X43cIZcuLlpeDQj93IZ2ggBnM9n5cgfACG1BHbMlD7WvL+q3tHp7Xomhob5qKTwi
CqqgNQ734C6HCPqllDgZFy6b84Asyk7/NGQlHsjaoPLoK8a2w5K+ua+DsFR7/4Na
XRQtCo/NU0S0ZFkiF2cVvjZl/2YlnZOFWk6Pm7hu3+zxUuMGi5D+IGfhByEv9d96
XZB8tOlz1JKuWVNDNB0OswRYn+wACgv+l85XVRb2wn4IgBa65dLMb0W544oZF09U
L/NMYLX9+mkaHLiUUe2bU9CkGEUvPph47IrK5odXzbv4EGwKm2R8pjyyb5H/1Z3E
YZRxrxde1iHkYho8BlYjkP8d+A1kVtaLdlL3NkpzYW8jVRaHrljupHVSEUOvB1JI
TzBgHFv6yY1OStx1juXPpVrTcyRC3lg3qlmcPQlTmVTA3AJI72cKSgP1oCtIE/lq
YFZeBJAPuziMFxdm/ND5SsU7W8kujQVZX1RAavVU+A0tAwzTffbeyqRoEA00SxoS
MPv9YJ20q1pUWXuGPizCGAhndXE828+SQkmWL1Z5f4tNHjU3ZHW8bQe78Jor70JS
bWVzKjXg//SFyVOHVDLB22purw/Y5Nt7HGtjl+4uEr+GuXijg5rvzGsZVbBTpHJ2
QvzS6rgdZhCF5CSaVio3/0+1T2DsU8YB8L9aVnBOq+sGZvPcjJma4TiQL1IhG9gG
ccdY571Q/YqyNxRaJFn2djLtTwX10+at+80RoCLHkaUjn9bPbPr8WmLM1B05WuaN
5ZbBh31MLdknFiKG+nGyJkK7bfcFOKqECeRzjiQ2QKyPApN95xjmj0lD8uyZvkQO
56GoNohxhWSmG2ZWJj/2+AjX3DfH6OTBnqQozDn532Xqm1j+zv1wYfcgnrSp/xdB
ZUMkZGzQqtaQSFIgHW0ILYNnv6aQE64vTCXWRPtKm4eo4MA3dpKo2BW6zRIIMo/8
raLQVrNPekBiXVi5QfT8QcMwJKsQ9FmkFemT/WoxPvjNqMNyDjxB29CJz2GBIkeR
Opc3jpy26aREPwx6Ar+VNGyNsDSGa2VqSxTqFLV9rTU3bwmeV4skx/7k35kidBK9
gXdEVgkYuiJJaPV1ND2YJpSnu5rrT04dPZUv51pf8chyD9j2XR1qErJHSPxSG005
GWagQRzu/zZ93QRKv9mt2ppojbCYm4OoFF4yk/WMVVeMNB7bESjyy8IjddzAVdH/
GBW8CO+rFvOKx/hhGDWKRHmDi2Gd8WVAt4NeowBpfQ6pJe+Cx/ESEe0BZLaOTjX4
s+HvXdUjTpu3b68qNajPWj9J0CctyAW00FVeYGhOgzknnKMQI5/ttnHhd4DBgq2z
GVdUyA5BnFbpgLlYMkdxxauEXXKatO7c8F+8my4sWFofNIEA14iobBxt16g+Hnz0
oLZ68LWGFakdUGiXC4fpeSZbDtEJrDiIWdyzUxmVBGhKem74/DxxUJEWLshai+Au
uHf0EEo+wrGl57ex9j6VaCPVKtGd7WhdQj/cjnfK7iAQioEuVfSLJdd7f8vbHlFk
ZN287x1GjQJp44Qd00Hz7t//0EwgM0uKCKQpkztDN6dUQOwgOleju6oQHISy0BQa
gIVfVIFFKUzl1npfjoWItJP5mgEh0vJyFV2G9ejY2SAMvwTqXfSbRgUAbEJCSGNr
blugdaJTGvHZouubuAHRij7Z54EDLfgW+20LuKdg4Xfq9tX1q42Yyv5GS2h4CVM8
h+rU7Y10mgYfVu1SgMDSjcw32ZLBQaz30UTkzeQjiDkvxR3mynSCV2FUizeJGBy2
cKCWTrsG59gcMk/rwMesaV8ExSJNpDvoV9IesmU/eOT7uv5L12I4myyfwNMntkRO
Xi/jvh1dQgwBaJgOR28SYUpm1RAjzsYho51PM4RXS+ELWwGVI4BA2biXDbKQtkM5
FMFtKjSndY6ZFqD0LXN4I7lQbJFmL9+nFSMi4/w63he00Od9RL6zl4LUTvOgWsCc
rHU1jpezaNsM0aye0xMPr7l6cc08sCsBr1/AdGkYnzRdEf2YemBQcgVzKSFvZNkK
O4GRPZk9YBlFywxr/ufbps+biGH2madLwP/tleQKDpIc0zNLzDiNT+tst+35wRhl
KEB+iWQavwZkHqAeWdMMZjHWAu1NyL/+gciwUdUAyL8zJEEsIcbWDhQuieIzz0Z5
n/rJzrbghCtilT+WCn/WEz623o+SyigWu2FjBu7v7aQx56vgBBOab6dTOaeCab0c
adhSWBCbZZNjO09nV9+oBML12yEtvL8HHPVv+OQW7DcwJSA02Unw6WwC92JPySCN
mYBDe4UTJ/FvdmgyNkHjQ8+XtdEaO8+x0ceLU9O9JVujH/scCj2Y9US6WxzYozSo
mzcZqfMhpF/sm9c/t4wclfw9lHTNEBOb+kmp+iQPAzK5N0Dp5jHJpgam7HBqiNkN
maX7Xf7U/f4MfqfQzQZE4pZhE7qxgVovQs0aTiJEHLCCPzGHG4mOEVvsZzlsuDBI
99FBvoYWubVdQWi3c58xxeQotsbZ3LgiUWPGWAWO0iwMO4EgDh8gRowjp3iPwUvm
UXifM1YWlpSK0/tFTP3nsNXhV5jQVyMipHZyjSQyrsTBnjgegsKgrTdOyt1Rfz8z
nQKpAEmbl3PtjJKrppq4Aud16ENKHmvJkMltfDmmbGWwRSR4/6Vrj3PZDDJ8sBq7
/E6X48YJr7OxGPrESPGPdFLKNpsZjTEVIroCeJVG8lIXJB3QAu2jtSHsgJ52Wr2O
C31U1Y+MPpJd26V4TvtGtOBjnD1IHj1UF8P3Ztt4UX1uznkHvklIyhzcwNdiwBII
wgB0gfa+vwfNTfqxig52+xH0nehWILofkJEbdleY9SCeB1iayofTy8tulOw1yij2
63E3AUqzlWGiQr+nOQYSglV502GyyGV36/5pGtnunFwqr/yu0AM14xUzYsDAmGL7
qPazIAr/VuX8XTCTdvG8rdGv9+LPJV/CKxjcFLj8mAXT04cH7oUX2na1MPjWSi6s
7ExLdU7AHekWN7gyX504cjPVE8H1IwmsgxJrf+hN9b2fNOSv3PNX8SkQAoGSnILS
RBhBtZoJYnvdGZEPSu0yG8UccmtuJwliHk6MxVMUXROrGotR0oG8r/GyvsF5FD/+
YdV2T20NRMVfSjp4N3hQNlysnqSGXj7fzjRhatbLBjWgWFRujVAuuBZMrxyYOyeS
8+5TMap81qoCtnyt9pGUnshWeJP6Ki0yR4FMcrQ64CiO7eNnchX52k7EyaXhZYWV
xJXPLEUtxq372TxDcemHR8C+I7dsM/dAdVsbLvqoaFVV5P2M0OIpvd9UIoL8+Fdn
gfXpuHi/g9wJomWSGelRLWdxkoDhcD03VVX/VZZIx4bxCeraUF8xzA5nLIwhMYwl
M+qoJu2LutftyEAHgfvEZ6kE8vJ+RF3q/ppTvUHt456cHKVIdfrynCS0GApY250V
l9KfxK6j/wLLa40Y6kHKw7xYDd+DhYaYHDc6XGVch6UW+wfKNV/GZAp0TX4EyRhR
wxTbRnThdmNBrPjb+SLVZpXbTO/Up8oe+6Gx9tfNFeDnhZ2TO6l5pVJhnErRo+Xs
fJ4Qhz5CVixM0WYvaYT+DsiyyQaFTSk/Z3kdGt3Q5AJ3jmqEkiCTQ15XZBtnU6hk
eVEmRF4MVzyR/ZNqZ39DFFKEfDimlowt6WMLr6TNmIefYJV8xq6Lqbyi9N8f/UYv
6BKrpM5kTEGF3cUsraA0z9o7nSqcpsX3aFSQyJi0faUymLvaQlhlG/98w0VBflem
SO9mLqtRKhYMi1f6WanwNcq2962MV8PxRiAW17rRP8yPHtNNf4O9lN5XXv2rC4pv
4fCBvyJtqjWZCCLLOEoglhcPBOWQUNNS+Ccaehws3LvNpRZ3vftGaTvTHeT48UJT
Ghyoe5ly6GuZLSH/eliHpJ8eeqC9jI3gQKzdUUoV4OLrmgWFavLyQ3Eo3gvATt2p
wcs0/yY1dg9OYzyI85swBvV44no8gDf+PBW/6os1vInrrujYde+o06K9BOyiMKIb
Ra2YScaIm4Tr9EzqaYOy+79JGYo+MRUJSciY/kNszDStEjl4CpVkx1a68fP89kLH
rZpehg0/PgroxzNuOlcJuImLzlg93brVz/94zr8eI6/1fSyw5N/34m4oI6Evuob1
rPnDHTpmgk0ylF7JoiUke8aBpHVnrBcW95uTHK2J+QJAyWfyUDyyi4OCikDyvI9g
ZCLwR4RjtuL7qsror1rPcdtbfvSeWMlIRPqs5s/nqp7ipQNGJI2Q6vJU4qXBe5Ia
QuomONagY+yPm7Ocmdp6kyZwOfPm9nMcWFzu65TZla1rMwah1m6D1xbhR6lpiSOl
sYXKkqL4kbSStwJ80fazPCppPgTrTzMXOrPyVV0dk2AuUmaB80AxoU87mfVPC8bl
AlDN6VhzKq5DeuFanIZxPoWrSx6VOs4LEtdVXQaVOhyMdI2i6b1cE0PvV5J3htK/
nVXHyQwdVC0zwUp3YNmjcZTFv3S4sPMgG/xvAPCv4RdxFpcFSFPzm5fVDj/xyazh
XquSglsllBsINwWElH0/ChLzoTFwdeNyce6Xx20GhFxwjBR8PMDguwhBRDyWycmH
rc1TS6oFQ18u11YwuuS1tlWyiBzqSIx9dvZUWwjEx7DlCCy6nG/8ezwqvZMagfI6
ycBnWYpyDhpIqoM95KoT+Eq5EocG2NCs8xiUEOIUBKj4EeT5kO4VauDxkK2XcSkC
Gz3F7ewLCwFEZ+IPT1LS3Q4tRrKFz9MPwuKMC7ZHB1wlvUxfP5CRJ1j4hjClEle1
Px0a41Uo9IvZX6P9CrN7Jw1me4B/iiR7AUMuVxPmuMo3xZPMVyjGT7DYLj4wSjgR
RQ+AhSItXrCn4rGoArvG/SQ8x1mN3oVYd8B2WNNEXUrKnufeHSC3hAv8+cxntik4
+l6XjxG+AgiE0l/S2WNuuPwDsRn2uL+Zof14fLfBKqNGBJnVLW5hgVC3Dy5M3jan
HsApzkUHe/EzL6vXw4/yZ3wOPjekmdUjD5ko8XQCpmDwzLhG4vXaN+rcyG3qsp5i
VsaIem1DTqyUU7TGXBcLSZBKRDcdl2kgqlQQkM9PmOhcowraEcJT6PYiiwUuMJKj
MrgPjz7ehw3B/S9Y5alLrzGYptHtGWMRLIdV+Yt1g+bflciZNl8G5vlmegQk7co7
Q/Z3mw/PJMgt4cpGtrzyDhfq3LyTAitaio/iZPRaFBp5vawy9GkuAith0z036oG2
se60DxuWveE42OIkXSOry2hyFAfBMLzW8N4Z+gZx8CyuDNa0EWC4zZ3c1/MjKIpS
SBD1cdjOAJnQWBIqbQW7WmSirtk/rZhOSbMwFlCxGIx1EhaJV2pIxbhhKcL7fh2G
sDNGNf8KxjsITnoouE4FXmHhRi+j617Ks0fjCKzGscvClWvzm0KybL6t/nDFilna
+eA/6+u/0XBzGuMZXVMHmVtXfZt1luaoixPA39Bv9PPtpFW7NWMqfU94yQkNnQGe
haR1FADL4KnjgKFqXK82YJBKzKJbZoLKAQE9Rh0Ep46zFy0ra4S1APgJ/6wtQeMq
dC4zqKR++QXL+5oCB9zzlSlxHPCADA3fboF1aYBESf/ILSn+qYgs/Lp0n4oL8dTE
iAyjzw0rrha6V/aSJ+qIc93JKK0zBM9l805O13l93iJWqdWEpciTKMMLD6E8BLpx
FnFTmvyHt7gmkkNI8tXVnX6mUKNLHhFOGhCGGei3AMmkMjgVymWhNPXkcEHtSASk
KUf7kcQzkCJhJ1xgA/z34dPmi3fe5SLCB7a01odsrzzUXZppzB1F5equkv1moRvi
oRwmN+QzxugrFpz+SLETKorIr8QCbAPZE9GN752Jw46h/5G+142+ciYetud5hjmu
5uCgjNLTYT/h1ypgtWJUZcDK4LUAYHYnYaZah7wDedfsmY8nSV4m0XAZMo4SENYd
pR2KE8Wg6FFqX841/mr6AVM2h+wwaEq90wmj+syVGWFH44RwOumH4Ap2epnIVt+v
ImT/XEfl8MeX+C5o3pJ6Gnz8jBkmOB/szktVTH9uQGFAeAxSu8Bnjrm0yDr+2/4N
T+TTuMS77X5lohoIHe/eu03TIM50YI2xzLf3kUzNXuOF+v64X0ERCLrac+5Wl4rL
iGsJdc4k+eqkZUGXkQbNmYNjoaI4BESfUg+KrVqXH2fFsCjPSE0nsXbR5urQAnAl
LnrQ3xRNVsuIGTHhXOKQD64DOuPeHdU7XEKhBjeNaSja27qAsQFhf3kiePdOA6D4
3POrWp6iZ2e/oX8pQbPd0u/CC63XaDUn2ty3SvJBj3JWpimjPxMIYGCFI4S9WBSd
0VZJkcNxWkqylGfMx/meIdrzsBkmlKWm9P3EPMkMtCkBMMjUCWD2n7L3K6vaDKYA
yt4pheu0KnGRNwVcalm9dT3SlbIhqxWBPjEpZ9UhyUpBCp8n2QcjhILNuRIBdyE/
tigIMJQFPxJtsHLyHKh5avfJz3Nb0SZ1hfYxReHhv9taGijrHbCN2anmF09hYjux
5h+Anm2tc5BdkBxZa2hkSWvqVxknTb2rrmBymmOnk/cqSFJ0MTKRrE/Y/qI0KDrK
vSnO2JBMF6Oa01uNy2NgctjhwXeQzRkpwXK0SrsHtzqCRa7DaiD6l60M8mMsy/Nv
f80VsQNBhdItqRXp4OiZcjVPRIZ/H57zNLC0LyBAdqfbotw9YEFfx7LtO3O5fZ9H
IBcpqt8Ezl2tUhrEo91C6d/hDZ7cKmxlolqfyJJsshOxRq73QAFBUQSuxdvDopPj
dcOW1Y31cd7yNYV0T0r0p4B/llcZL7SCHn+AYwR7Fu4uClqvvAwehVgcGUbZYgeV
mo92Jr6+sFNoCH8N/pVAMsidB9ymntqh89bU30UoSoj1BbsTvtP6NoftleJSeMZK
/vj4Q9OgBgHkQB56tF7Sb6IUblNZaL4cIQlMUIKKVVk7mJ/dyIJ0dZB+7CGLw8Rv
xC9rdmwQPnnseWNNDGjJxGjqstTbu8cLWTjszeepyzn79rSoRpFfihhkAYkLP+n6
p26DLeeqGWykWKFYV+q408Z2l27nAkz4G1gId7Xou/F+UIgsHGuxwz3kItwgcTpL
zt6MoOKCI8xAvz9n5UfhrwPAtzr9zNefzP4tv8eADTFgseecgRz5uez+eQTnZ2gt
Jrx6g1HFibodv8tZ0/zFFtjtqtJ51CJJrJAn7HrfpEhcsz+moLaniavMz9ViB95m
sy9mW8VDbp+CIunvxis8Y8LA+myO+6iqgyB1RnN8DU+rhhwgDBs6wGCVoHsrEpgq
Y48JZ0wep1IKMU2Kl5tATdOG7BHIGY9KILXkfLLa4IkQbory30VgPtbgRoHrTMWT
DqVMklCoXG3UPIjUbT/oKcWiUIJEx8bgzhy1KUizAr7ctLXEr0t/7xcB+quonOFR
nACSaQ3FU/aqK/JMWTb0kIa8buocKxjvu9sxBRlsDNa7TjGY2ZnWONjZcdEnoUxA
hDyHpx3g62pjQmVv4bx0o1DJBLRuXnGijTzJGg/fHPIEYWjiCHvCp8Uz0sGbqi9y
olopn5+EWpkojTBAEB8zbMfLeMw19vOxa5Tir187OrOiMAiavAy9jFyS9Q9o0qXx
ojtwLsjZ1C57BKiRbXkn84KIXdafPELaX63nuU8tRNp2jZaTYdwYRsc60a6uaHJf
o1f7gcmcM4J/tu5LY4gk8/HgGj0sXpLJzdya0pUOFLLEqcwSTJVsMYHL6OzyN9rs
7d+0s9+pjhgvqTiGjOe/2zkWJtjXKA4fBcVeE5GhL+dHBCvRojljwvPAlRKfIyCG
N6nYTgpnQGM/YMgR/nblu4d5Mk6R44QtBEqh8mHyGB0Fx8hKenmkS7G6tRbAakRk
cO+glDnuuKqohyE4/eZ79l8HRECAxG7ch/yJ7x/rfYGEM6/9xqLExcLBc8+ohwfN
ZWneiTYziPsgGQeSZAoxVEuGnloe5Zz0cgM6lnuB+OtAc2VpNCV269nfUV+t95jE
kDyXuSXfXr//Xg7glTnDWGbAQsDA07HzvxwgzXP3bj7GZ75XfR3D+EXYRNnQ5YU6
m55qH4/ynXs1767GP9o3gFWlh3oLlHFCafkZ04sb17/GH1kdnl/bOee08k8kJG9C
zbhC0+wf1fgmp6hmQNT+O/I8NcrvRlSd42N5Zosxvq8jtxZbx2ofpXcUrliy5SXd
yKT5uhdFqq4UsCHyqYDlvXL8M9gkdV5wXv2quX3wxk3tIricS285VdD+5Vq8ETe9
vQlzVpuXh85F6dSmzehPnVVaAiVOoPwrp/X1Gq2GqwUIaXV77SjM0w0BD46vhiSK
GFy5tskzLGSWusWzrX6Bii1EJZyBv0juIvaNfWJGuayr1LTpeYcJydPZja4mwjLs
yb3GVN0Eisr/txqvYvKzUNuYATD3+S8L48abRZXZpQaM1RAI8tVobw8sn7j2pTDm
3ngxnqfF97yXZKg1I858r0/75CDG1CdSEFnMAAWmD1Ph/05w1scA/1o9ptUoVgqt
MftcovqnHcjm4xfbLLuFfDAunKGmHO6ugwP6QukTmV44L0poNt8RAV16EQ1BJgsa
qw6X4pYGyJ8KeJir6t37+GmdIprfuofhHT3ZsCVLGgOStn8uSjF1XSZqMPAcQZ4R
3DMACH6p5AOAGJrQaOzfpuzAMnINNce45ue54Sqwsx9n5I4tG78ETCVWHkFeIsJe
ah4Yu8JneRnyPu/CvL3X4WI7jUiuBPYwBOGm1xe2XRdXi01al7c63qYF4XLuh8nj
mLGS+BzPjWk4arvyoR8E1KoRS9PspILbe565YLD4e2MoTf4sOVjKBUZVChzR1vxb
ooH7HKEoOcHYBnfV2FH2tSvA43LvQtw4ndQotj9RN8nXd7ncbGN5jy+24oyMrBoL
MA9Hb4wEyX5hUiM6V7s0ZVCjJ5JkeBc75xRatlOvzus7x03DPGiKq8oLviTS/Rik
rgE7ocxNyIgn4/FUkjUeqtiOTB/sci3MYcZb25NsOBO47CqjmufMOe9w8iVBGZno
//WrALoutO0AilpEq+4Qo7CDb0nAI+SMxNi6uvczw2CjEV0YX/ma5kgMmr7INEX9
N+zQrv+si5Ss9RHWRfjlSl5ikgHbFB5avTQFLFrD0IQgFSNmCZAILyvYAy6xDD9q
fQFLZYABUlh6bhwFbqGnTMhUJ+rYXwj2FGEiL7MFA4CxkWeO/kqtLsQGMxHqhJ1I
9XREYYFngk5687LN3kOgv6DIPXLSuV0nrLX84Zi6A4haK6Sg7VJYK4F7NsDo6FLM
gpJ0EyMP/oPYL2NsO/xW7LEVQwqbtfcslgzhucU1C6Pwo6a06+cwx8fbP55ucFX/
jSl/0HIsp8crvZu+dkiUbRZ0L8l3yumxPq+1khSbjc+8BdW5pCLmShFIl6uRHqCH
HwuetbiiIbmkwGiqMkWMais64r4OhXEZdl7rEFMQ5G4u0u9BpUoypjesZ/0mpqqw
Ehh6jMm88Mf9aGfVXVOr1yNEKiQTVHsL6WeON2OJeG8VBZ/gf0t3vDiYCLv0t8WA
o27r2pDu5ZILAHLliBsHQW7nG5tXvA0H9UyXhSGqq7sJJC56G5TMOxOXItAnRDbQ
NOQNX4qqdMpjGbGYfZR2NJLri2p8OydDb/uFQM2CDEHRF626Cy5YRYkIyXBgx9/1
5DflpK2A6vCp/ZM6JTKSp+xfNQc+aD8DQVkRQE0dPhruP1knMES0h3spBjJg+gOx
D3ykxjKCAMRuoDtEedK7LxQ8b4niyaTArxK5ZzHuAdfTqCT2hJcC9FI8soaWXsc6
knpIFmJ6u2UEQ7q4B5Gp2XCIOZpgyVSkEudN/45E3urgx2muRuPk9NDZ6Crx927B
3RvBC8xaJ8SAESLzKEXBtW9f/Hma2XRbQ5G411RH1z3jjkYFxfL4V92Qzr7E2acb
MABgiqQo2qDOTLJ0q0Ly3PNrNYKuTTRuiMEu7uwxO2cBzgQrAhJHDe/oRsLlJUzT
OlruXMe1IqxAKu18m4yad6BzqB6yOpJlj/fnhiNmb9TzFu8tEkt1ytwbBr2VmLxT
mxMtrHRtvI+botNGTPiusx6oVeCXIF9VmJRnwIzbMbZ6RFPrUggymtBoLvweHMny
JjhMmMe8l07G6o1aZoS5YMGyQe0i8Caj6l3+znD4Ve8tbRgiM09yCu1js8RR7NPZ
UQhNycgtAHb7/YyM5zPH1lPNc0VW8uFwRyt0MsRTLkxyfsJKXjxMvJhJdRfBA9/q
HSy6JnMcfUaag9aKCIy1gvhPnZnuybGtIhCkQnM4wmPfzAs2bcdC3kPQasL+sBnQ
TBQa/yOv6Jz8JrTGHGixM57e60AvLZ6a9Oornw0ZGPCUTuJV+i6os0jUNmfmnPtN
urCkMAkCyr7ek8HdurzwjzWYDweqgPyr6dxA0we8QEYpTLwfLbstT098Hha9ipjG
zYXq1Sxy9eF3j0Iv83U4Tt62sqENvPrBW4CY7bOYQbWGWsLFXhcmK3yOuhRuDdqN
DxUIbBJTpCU1vcHtO+iV511qwVOeuG7h2Dzmobw7EtEVdhEw97hOjXc1uzeyiuae
D+KvzjjDt7jGXD0Q0y6CUvgMuegNVCc2FFYf/pohvBaWEj3+8ZntV8C2+2aZFupi
IUgwev1HpYHFs7Kj9EmpzAYqJF1qL1P8+rXTZoO7BD3Mo7IOZaO/r4W1UIDVDzzs
Q/wF3ORth9ZATvCNAfuOXfhqzzADT8MbGhTq3fXsGcWlhoTc2Nv3MOc7o/XBukO7
825eKO+aPAUb8QWBfypb4VRmGHshMTN9ryLxYjRYmUoOkZT+nohFXOO1eUqHU7So
28mUZ+GQBUxAjaJ6XtTGBFW2gxcRqs2MuEhv7wXwPFrNvW4C7R6PRd2MJLb3dgeR
Z8V96GqbNZB+WE1+bLxNJJSsEu+RayrdsyS9mMyGkxdvRyuuLFR7qa6bNkFOaC5M
F/xUdDs+C8M7zO+k+8T+wDR7LA/Wk/Mx8XeyrPANo8bFIELUNPrdvDomJSG5gpHC
wnw6k2gqTeL17Cy2uWDvwNVvouP/g3RfTfQPV52LfNHyo8kUHzrfO1iROkxAhlkZ
X71Z9ocdWp9oDOaUJqLF0zs1UFzSetBAcenyNOQpIIfoH18RxrjPyUqdCOt9SLWV
tLiGzoe8lcBddEFbqjHmF3XLIKPQF0M8J11sIePPNEdwj/gYpkxv3QlexnWqpcxD
Lbb4A+ty9U5DS+I2kEKi+fgd/4rSUxEG/Xxy0V9pIPLqdEgyBDUcawoZkxSGqcsN
FZvAbtfSk6cCI2Sgn0hDayrmWIdFr4oK5hNS+1033B7SZzKRbH7P2k2ehGXqXlAi
UtOcsxzpM/0oNmbvRIP3qa/v/HVq/lnu02FKtTuPQ7vYMJxnfJUQ7TKAxtUZgH0H
laqkjPglt1n67JmJGIw/K0kGHfTeR9idH++CokVpnXlC8vJLjHpI6RxMxCVGwsPQ
cF45UI7GUj4uV1BLjklBqEOkyWNnFr+pPlsKheHkI++teAsgbpgqoOFVAxZBLusF
1YnkSJ2VKXrj7WAP0VY4Fo/v+Rn3npt/A1CgnrZJkRaIeqRSqWWsnVQp98j65zpt
HrtQLTLJ873pLiKUfhrn68ToixwTcMRDLpncBNvtduFShkqBwguYguc23RgXpfk+
ZPHru6lJI9na0Ibn8QNtonkU8zIwONxHuUVbW0ojWYjq8kvJAvVW0nLurDPXonrb
SKgvdnZEXnWNOg4OU7xDCLwZPtIN5HlPx1VyOp34X1crjk+DtDTQyHzAgPoR7Ekd
x/0pO7913l51zxX/XSG14IQrz5KuoBSb8BCWYqafAYS/Qah1SS/4P2LaxUpjUixL
cMkmanWmUt17jJZgvGAyJdOl2eQI8dpS5InWWIc5uW6PtAqGrug/sbzdth6g4Qoo
DHK/C2VM0Ik+y7NC4R94uZyqjEuPJ1XupBa/2/ahmS5BiFT9CG9k+NbMph+lLQpo
8C6jlXe43+NROxI6deMWRO3nq9X2FOEwQHdF7Wd3EyU8zdtAZPuklN/6UH8PLUoG
tAPVOZf+4af2Xa4LyuV0+2pReR7nbgTO98FfyjGobC1TB81UsvmQF/SmJmhFdIzG
tAXujUGK/s6X5wycMCf8UOEkGxnmc5S1qfhF5TfE+Ijy7VPr9GXeGsaMdMtlzzAF
yFfAHKOBqEZQr9UxcoPwsD2Cv6ZtHm263CVSTKCYRfjLNgigaIPKlVdGgihUhWh+
IF8YHOZuw7YELMDJyAcLs2BHnqB6PHRTXZClofwL17IfHZD2Cat6uJwU2RGoDjuA
pAekCGf4jT+AC51zJqlfa9UqvQZniHOZCKzLS6p7u3b9jVrsSs4cxoWpXBEkHIDT
VDIeyHX3eKmVuX8zjkyXsUZ+2SvUaGHH+m2FCWMmaO8oSmPiTxjbv/G01ofKArFy
Vt2oz07524/WG+RW/crz+5TIw51TkREKCBWoDfSBexBYA8sEAZx0wf/xF1iJyDPV
TS+DZn/oxINWsrPkXUeMjHudFOSZC9gNgY5c2vzwM60KydYgKnMbZnH3aZ+RIMgB
hwvlHyoY/T8cFV9I2sxw3tCwOSSkvS0LCSqiOTwTCukTmP2O5bxXfwuhT2DxupAY
EwWDnZZmAePy4LntUKxTRcQgM2V0O+gGgPJvgLGD0MrtHrfCZh0pbDqcqdIqp2DJ
EXxzv62yX+qWXHHKoTWaPAzOi/J50QRjjta9Oi2Zf1lNx/qhdRtJ+C2TKPQp+jpJ
wKt0D5ZsKRtOYmxnmyiuJeFSkkdx7KBR2lxfPch1fSWBOLktC3TW9OxRk7SK5Sj0
V/8HWEp9JserFLy6X/ObN4yxcexCLO/gAuai1dbrjxiPhRS+6vcm/IA8KA48PKQp
KCPPt7nTS/4pVRnd6L3ht0+vLxxhD4zfuY2r9ft/J10Nk8dbY1hDx4hObYSicEpx
KMhzCD9L30E1fALa861tIgbVzlGgQn8JLF8V9tVUd6A5dibZ7oK4NzhO/uZbyAmh
0PEAaKNYjaXUSdnrLXQCE/hIp5ckTXpRZiBpNu1bKUzleKaVQUEVaVAVrpCeQs3Q
fW3Meg5WuxUMutwKf1GA69AtOQzpXrxwaADylUMdC5Zm1//m1f72ZVs21B6fF7va
1sswSGZMaZtf2fsRrSjCvKP7jANOt8E/IGylncE9rIeUaNOOZmyj20g+e5dNzqgw
R+9zBEqf2MDGhKgCOdqH+RZ+RXpzXi6qi3jpvOfm9y7FZNPpMnr1UCFOKrOCZnsz
e0yg/bUnbJn2KyUc0bl6C8G1K/oFDK4ccpeOYYFvy77d1sTdlag3VOydTcf1QVCx
gQFYzlA+VedeWb1QQGss4WYpDbisbsbNUg4LmWciPKanrOLg21tEJXq6iefXJSrj
FR9mvv5wajpTKWl2Rowwy7bpUDToc/6DAMt6BB7NhlVDmN3d1rUyO+XwQhHDqFV7
Hp0lI1V2op5rubSiH92f7z2aagFALHewfNk8U5TRlHdjvyY9nhGsdtwYSLol/7sH
MHA3W82HCkv0v8yR18QD9aiLPMbSsl0SwpL36Lo8l7RPL/BLpawoRYxUT2wjLiAy
Sarl+XMmjObEBVM1MrXpF8viL7/xbpaAx1eVv0KeD5SmlZXiNtdzbZmFIkThgjWe
2EL2gRHoBYCsH9WVKqGbd5cXAPMxHjjlltJaWvfUJ/ZNDenusFrMBwURTgKnIiog
u6NkTrsZYy+HizeG6kgNxo8O2W6nQ5fa5ItCIHVAvzFgSzcrcdFxbTU4I7gYba4S
QLly9XHBx8rxQYwah/60xyvAHENyZjvEH4uixnoQ1JTWpV+g1Frfr2ouqljbh7F1
KXpCt1+8GbCRaJ3GTxRwlrqUA3rng9ubWKOMDvH5YGmoYk/94SHR9KsKpkzgtQmj
vgiPWwWKV93W5pIifp6JNCfSgYhHq0akbDEepVDY66XsenDOe48HyiHet17rlTtK
px1ffC9W7RG6saOlrwWmJSByySl8gSSLmzYqY+gdwJvCIRjgfEp9NYIAykm/FE4v
JcxthHXeSecXK26SuGOe05xMmwov+5XPnd3OTGtx1qEPTtVFXPzf3V8q9RuETc7A
XDx3u6vp9FXxxnjDmH9eC6Q8WuXSBbbQ9iEIzMxO4xTvi7G2aOwjz8+vHkvyjWbw
UBsAZaxxg692JVWTzFZjcbz4+JPpYRrAIR0AQz5zIEugpfAXecubDeHMi10uD8JB
Dfa6YwCLJDrU/8W5bPBDXSZ9YJfnAZ2GCRbrmA1AvbikEdAjqjHBWfJF2Z4Z/uHg
eZrMVedAcaS1wTT5prG5537SZCG6DwnKD1vvpPVfzAYBZgggXU3x6WdV280zhDiP
ccHGlEVj1LYxOVkzZ699TqeKZYRtQqQgvRAxenILae5wtAR50yjxYpVFEdoY+DGm
699ZPYTwvThUcZVOo9l0vNxe6E1UTthQxRo2CkueSPWSqZQ8/9AsC8fMvu7fgAit
AFZfMIauyc305E3jB/ZmgLgSbtM3enWnYCf3QYr6T0h931egG61mi9gBai/VCVBt
FSu6DAVgQIhwM8yftTKivC7p5xAnv/vUSNLl6aP0ufvXAiktN3t5o3GAiUxXeUWW
pU3G58hiFxirgWQa3Alhz9uXr7uqYDs4ntfYJzIkE3nNsgWvkf7cmnqu6pfIfAbE
amAUvFX19/M0EAAJmLaix9lp1WXNzM/l9onITvh6nBGCRmsPDRPT4T9yhzjczQDY
QsOBti/uPbxosr5J2/BIYzPkP1plGyk6+xyz6emyx2D0Ai1G8peAjeAz4lRdZb/M
j/6kgzjwnwtbFnZARFKQYczmn8UzjGN88RTwbAQXDX1+9H5z+ETdm7OaltgtMctZ
AKNKMcNTUGxS82g+FLci1LybkgKgF3bOMws+Rtd9z5fNNFXzlPbTeak8JyFBpAdE
u8MwImRiE/vbW4Fs/fplZ/oV0E6Xx4saufT6+JonIr/jDt2pLZ4HJVcrAohdVTeO
rZ10FSkWj2zKjzgjWTaaQOVq2QAPuicl4G7EIxYJyvjZfa9BA40ay8yU2kaO9k8f
KUuNZ79B4UXkwwFbpjWzRPw5z0WY7fHO74VoZmO5iGJmVpmECS12XX5h5kT/lBHQ
Vc48dzeUxiNA2rgT+dgJEo3Z6bYwGpEIwPDHTxNNDiFru/ZZOoC58R5RVomu8uXw
+ZkMGdL1UHtdYwbmpSUVo9TkzI/CKiRxnBdwI3gihrLiZ1Q1ReDgqtrqN0InELfn
a6RH5qyIgzWyTH9g9Z0gxBvfddqkGLoO1xJ7MAnvm8xFksKD17md7S4a3a6FiLVb
m+VzZPyefgwG+wHX5Hj6Zuro2urYxQeGso1Dhrvae4Zl5GriHB1BU0wtN+KHrQkn
+ynh3QQDTI81XWou+Qqs+Na166uX4ahd2Ewz6VVQmP7UoYiZSY8aiXWvXztPHuzs
oCS++idsEFAlmkS4p1tNf+vQNtH4iLz6vjh20Rey2V2JV8AWwtzY/hV6zDfMcz0E
Z0PVtuljwz78cr6sRYSr0QtNF/qoOcRVnv8+rViZ4YUKHTd7p3F8D6tmv2BBlRs3
6A/k8IOZDTsCNww7PCEh6pSCDgI7Fj+NwmBu4+vUeluOkSEF/vvGk8yfpEuy+eQs
6xH3a0HL2xU7/piwbI9FrSzBqrnph259evPnr7bumtQcdDWD4cKuE8YQTqooCJFX
e4qnvPxm48ofNec9VpR4QU73VFim6NJh9uKswJjF3e6erVvYxfjSgDnmjqYMjtUy
BKV8GjeDrBHtCEIIiDL7tvLPnL93fZrr2aEWhC8ToWmnXcPomHIOEyFvM7hupqfQ
qpeUL7fwaZ5uW8TMpmOVS3gb2qQVNjmZD1III+HK6Ymb0qMuje5V0K1JNkUbSV88
zfHspBiv6WCI+xcpSg9Y1ynXws2lBWzA73NThplZEC3oZWnBC0wKtzxRpmW4VYmp
c4Qxg50Xlgqxax/DHr8U5h1vpctOtnGK5+h0JdPCrT9jBd588wsLQ86Gcz2eyt1e
Tg8UWh+duJExJUjSorE6HaRxsGxNAHX16tk73NeDgbzFcKp1LWYdOORn/n4+vPdL
u/IxrhtkrbIOn5kr+XRxzvilK4mYcTtKeb5BSdE18ySYb6ndyWpsw8bOBvKPG4DP
SYGKVk2bSYqAhBf6z6j1zTVlgce7cuzoJOWxxpYvTvzq5e1I1cQpYvqUUakXO3vw
3OBsNWRiD2ge9YUlKRagRcItGLloPK//C2LHrPXWN761oyDcTbyp/5GXk398r11v
NaBSdKNSyMZum79tcqQ3VY3yOOdLDt8rauolgR4jTlKmrxRevvfsRmE8AZN/Aqb9
CM9QwrDMDTgqto7XOkMGUKvtZbb2hY6641NrwkXvxqyyFcMtbfnATNrmCMqIjzxb
VoSlNN1Tf2DswZe0/lpLsfeNwvAl3u+AzJy6skdUaJAqIteqajxAbkZv+sIA5qTU
uebGNv7CcI9FFG489Nuf+atrDsr/1NOq2KTatBkDZKckqPUfeDmi66zcjXBfStVt
Z4CRExXqFSUEXx1/mSo72Lnib9AFIOQDdr1KXu1QUtIzjX5239zvz4RJQZjDQkWp
+m6ZlKmi8A7e2THw3CYRaIBHCZK7XkP35EXhGEzP3rOCNZk3fFWdebphtTNn4QuH
gIzf4ziRYMloUaLYuxZmzC0mThSiUOBJRsq/kUPP5Ot6PhZ8Itvo5HkHhcYqUHpB
T4mfwCBfkc1O5dDD9tAKiOr9EPiO4KDhYqeXV8yDVLZTHCg0eXnV4LnMxHZx9sgd
ZOHS3CQYvMLiGoB8sGN+fopqFgkVruugaXWEetSxx0QATlOPOGQ+bBF491QlMjVP
QfO70MQVri00hwKLg0G9AHJgM+PlDNK3GbvGKTqiacCEuHFDIbGVH/E5TyogiqYq
ib5FYz/VnlnK5zyqO6P3+zEn6EjMJ3808hWzdIdDrX4mjzTRYLgrxF3ge8isGHQp
zU+IX5PyGdpMPgYRHiRQpXc0ZwbAKYptI6u5ZRMWfPWW5ZfJJjv7KjNHrzgbgjMk
8rFddLY7VW0Q9uFdy/PEXCtCrdAMSd8GaeTHvZQlY2PsHsIqcDIRnCrgj4Qfys+u
dvdjs9G/5Z7NCVI6LiFXkmnHzMKIySSYt/U74pOi4zhIAuzFpI/FN6J5X2/GPhPF
asjsQuUC5XOL8GF9Eo9AdbvT4+bij4nQpOtigDzXLgH5REg0XzrobATsXnQBcBQV
1QE86d9unWx55b5FoIaFbAF62uv2ihs4Op8uSaZSIGFgHMBEuHOzRIxgthBSF5a7
QfBprhpa2VNLfEqnoyPWr1Irqeql5eIrUJYlbDoOEzEqE2v45RBJ5Hwc+ErQ/7GD
CWxZ4U9o960vfb/fdLbOj3yrlXQ0jtynGYdRkLH0hVDAsGz6QGwYRTGCNW4ZFys3
TyNlcV9yR91b2lk+6CBcg2vq5h/rJVA//9TtfKEtAkgoiIbCali1hKnfk1OeNU7V
QWHMopDB/LANgCTFbFeYZotTtn2dJ3hOiZIhHqwtfOuvLrgRtRvU17BOurzTZetI
WHsNhsv75uOm2vgyckdA7W0pbJnQEQ2Sxk/v/GCu+FMNoLcriq4XrsxkCZHeNZFi
jfUrkeHIqmUra/5SCKgpdfznH602uW8YfT8LDAvuq79mJCIlbLrStPhUWgGycpFs
Z0/I6s47FiqY2Oy7zG3WTSvcuifqQIA6TyGBO58XOLBLz2Yxx7MIJcOOZXHGP0ZI
0h/V/jmyfRygAALzeouEby5MSp38jvh1qymeUZOYSjZNmyto1viFTkRi+83shhTp
ISYwJRGUw+CHdPlszeYGJgz3DGBvboxMTzRom0lKXwofoY51SmUzr95ihfiur4EF
gNWLI/P03YrroZWx+tn2EkM0ewoEiFRMxrNK1qEdFw5k2K/WfdzuC4DB1iXpibjd
LKfwW7hRhEsw6GSUXLc1sN4L1qQigqqChJMvQJfEjaRptWzVvHqeHL2aihmf4nlk
On+k/lRWM4wSOrKCNqyogwaIiG+fUHcIJZZHUL+b1SpwA8tGpcs7bEl28SCA1ppY
5htZHAfRVlgar2CUxkFNWO28l2Rhuk1xiHyf8XHKCZrDF0zXjLAYYXb2B6IIiUwX
wpa60Op8kHpyEHKjsUwLXB6uCUme9zaM0yNJoNwFdppGH1pyMW6EbKjMgmbTE3MR
toGPAquMHLOaY5mrf+lmHrOUY6+7twetbaclPKpi1rjzSGzsdAX3KH3AVxICBX7u
QRGcairKPOuHmnto9cbcG+WOGeJ6LsF+YlmCs8w+w7T8hoyiZlt4Fa0XAonlYnEy
YiDBS4s+qX3kIqgn2qZqgVjw6coAt+DgDu2PlltIHFMaoPZ1j4C8ExaQwzVemEz+
sLvC4aut/31fd8wybQr1HbaOIRjf9+8CdsXlwbyBLuKW3BXDXHqL+0GO2nIbteRl
/20umBEhUQdTsb9idp0Y5UGYzGRDu9bzTAyI4qobfx9l4GHHJoBYwHeVLWl1RcsP
jSNdMiuE5UKY6RbxzjhzgZclUeaYWVIZnEROIEFfoHxIQWy5CY7ahYoauxwlowA4
HNnxLp87Hghop5Fy/6mpAzp8TVt4UIF8I0DgewhaJkhHvbvKhSrddgsELnYPA7yu
YzF8I3pAE4hO6C7wi3Y3C5ZJXFRAPm2HOdaBB9QmVPmhbPdvQZehvuNrTJDGzGf7
8IyMAINwCPPNu4lrWV+1SVBM8cAt1C/f/iZgeFlXbXCY/eaJr86H5wAd7QiibXRk
lLCVBEL6weI1an8Ll8ZuPYcz7w807BLx/OKWuOkWy29uVwfQ5Lx1ebcbG7N1+Duy
waC0hKBT9vsFRkdZ1aTMTeQP7xAyUIt8o26ffepknVKPZawzjq5m6fbhIc9RvkFq
ExOPEhjvmEgdaBQQe+ZbeO7mrAX9d4jD9AU6yZLz1ImWmlxwe/rhiaQEM/lNdYtz
9/IPqb0GUCtUg4NDwuK1GXNUz52mv0I54/wbU3o+P56U+q8ai1tI2ZLXvoX+T0h1
SLWvsJOcaS+6iCHo/iKAem/SGS9OpfHyq0U1dOZEUgF7FrKquxekOwkQ6nhGWRP5
ZaeGHoxwg4L6be4dZGsLsl/B6Vexjh1u6+JT4zdgZ1uZ/RkOyyxkH+48pkM0GMGm
5jqRQ0r8Vcdxk6RTqozvI6ajudzIBuhupeXPJ6SdXZ7M8JHkObt3j4aHO35eve3x
mIbEApiyBaqMvnYeNzjfzxODYIfCP9PdcaIzlcyAqGzoUkzDJAI1rsBGwAS57t66
TeURXsXK9OLqXrsr9pOSSCEGVtrA6BT1nD7ZnDcMhJUdtpaLZqPj/uVaul2loxnZ
I1rocsYsi8rSAIMKfTLOVUzJwHQV6lJFHDnDi2LTdR2zkxybgmzSdqAv/dqdl/1S
4YU6xNmJzscjhlrFdCpcJXa4lUC6sPsC2ypnI5B3mvGWf1g9K/BTYDMrfUAH+YSP
edFpbESBZRqJaYm2WfVUS9HZa99PPK+5aScfd0x/we/yWksp79jkP91mpRQ0fGwq
2DrrXz0MsbutJHWGaXZE2+W/2mHQv7esL4VjOdlUWJ3lzOGqj7DuOGxXFyS5XYgn
cpD4DBTgGNfdvJ2isCWk4gu/GdjxDZq3NL7YE+58UrhtkiVLMQ9DXBvXUYeRUksG
ZirdKaF3JqVNpreFHW/0143FFWYdX7Em1fyFtg20d1GOFVdggU7Q+q5Yd/zAhg8i
fp3w74jPPFlEAVC2gUWp3ED24nXkCUH6Uzj0SnOB6f9K6TVjo77sz4dcgSG6cVAc
mbZ0gGBFVZ/11PFvXqLY1xv59+5IhtDI2Nzt4eaKL87A6+7ol3IEiP8SvGoYCw4W
xzuZWYRK7w8Dz+En2/dmMiaChMy35ILF5Cv4CiWCIm59XhsK7YPEI9CJtAH6yPje
aUZTwrWsjocuY3dFdMV5d742kNkQmBYkiRnE3kd2ZLhOR4HhdMmL+kdV1pRZoEwI
/hpsWzSNugNgQ0Xp+mDG2vrGkvQnR7FuxTNnK5NSP0ZN13QUE164AdsjeBSksNfH
VXwm+4W0f3bC419917i8MZR2ZZ40l1T3qzOiNwdXk1OoUdIo6XUNeRcuU3oCUis+
VQWxOg4fawDgZSnalxjUyxzeX1MaMODjrDYs34sOEQN7wV1/fasXAfp8jYMJJce0
pbfYec0yrnBtAkYI4Y7gd55Wlo8ifAqFIMYH0L/PhBcr+9Xl3ruetx+snViYAqmE
W7tqN0kWnZAqftkYaTz99ieyhiYUqe8h1d6TCD+bkrPcJu8Y3NDpKhdN8zkRVM1t
3//k3PXyttMCNGaAgdhP6T2dzFVxOQYb74IuCcIXlMQTkYzEQph7grtBrfYzQVdE
T7JIvVxUm7sNFGmMjqCwUrvsZnwfuhg0ABe4k1yir1YRnXf+jgrSxyXlEE7cjdND
Y1I8IUMYDYYL7BCoO/HPFiNHEg/pLL6R0UadT6Lfwl1cIsgUlkVBXTwLulAPVH5D
dvdHcJApH05TDclKkA/6W9fepXSqb1/C0WpnETt/BufZl3TSP0a3/h4mVbNDCOtN
KOrTJHTL/yQxBDTWmmgJLys63Yj2DzIFlf7DRex5zyI9tbwMdTlvq1blZny5Ytab
dyYkiE4ew5+/45yPjiqGoDlgs3x5TKy/jveMj6g11VyJEca9zO4sOEeTCumTwnCW
BF++O2bS1XK6/jWXpJoz06mdtUw/4Viz76wx8rZYR99TzthJMUskTId3agGSambH
9WmfmgSYfSLKSGNldPpWgbqTyxypJJqeuEdARXuDfxpURscmPyGncMNKSVrjPsBL
pJ7DUu3FIB8b7h0kbsQkMi1yneMvI+E3yrPKcgfdj7H/dw/Zq1TEhQ155eZmNNE8
6XQGs5diPEzRBHuNOizPh66t3sEx64DC+AKMbhmN+mc/DT5yjW3I0lIhfuEEmm2S
9q02+TJXPnj3aOmouN++b9j1KbpFfsYnGG13SVq2HvxJgPa2sTK2aMTTw3ElHd6i
5xlNY6bt35tcH54zJK2vrcO2XY2B44S7qVhaNI6wKjhjFF17k1KZyQ1SOMCzA1z8
Gjqb2FYPM5UVF84eb08QJ7aIaCdGcoQLAVvCAH2i9ql4AfDJl8vXOG48iyiGLUvu
119lQdkmAi7DaxJ2EhvZ8coQu7O3t5dxr1mntzQQmdxCQwYosFv2ra6V70XzNcmh
F5K0aDrpCSn1IU0XLTubCeTzzZoOvX1cZ6BhB+JnhNvxltGZ9GBMLQNNcI+OSdFq
g+kk19ayGQ6s7uuz1XR3swLKkqFOEeObo/nh+THca5b6R78sib5Jfpi0ZKxcevIf
8I3LJWj1JYlvt0i0wEefSsgwoZ/FK/thXY3HxD1UyQS0gkhfwT7pBub1ir/8tY7s
tUXqjn8b5rpS8mXZSP3alQ3HIpaHQObxTC9VR5hBZ7gw0ofDE89DpIRg6qWe+ssu
YJrFEfRLM7G54C2X3xRQCJqo5wsV4T5MXYWwfZ+RzP4u5oM4ML3IsObCyFqKFEIK
iS8xJCVZBtOC98uUVMMjXez35NhWzL8DJSKvByf2qIvsKh6ejuw+na0JlQAxan85
5zTM8vJXtG6rbetEk1K4tM5kuKVDNzbYBJ62e+xOXZuq+P799Jdq8x/tSsysgr6o
4SmEkOHZ0buPKBQqrxqjGc/f4i/MOwhpLu5P6nOd7lZdbwqTVCW6UQGXTOHrdoZa
dZtNNt0iT+gYLMcMWJ5sdppwbYK/V+Ps7NJZaEfsLIcZEH5/zc6DlpVdE9MibtbA
kCoZHJmC6fFfJ9LrjrWUZi6TLQb/ubjOJen3TbqC113ELQwvSLgYvbMByTH8Aok5
QX/wXraJYgpC/EZ+9E8OnFtrAngtAOVw3DVHdhnhuk+HP7SsWsMyqaRLPr+vTXZx
U17ujGgqjaGFB/IFtyn/B/jy1aI19Eambqv5Eud+O6Jc3jyGBupxBXtcZ9Swf025
X+bCjGquPGWsbQ9X6U3xLraWE5XpielhlQcl3OPAi5meICqyLuZn5A5pOBRR46oP
qfZPnoMtd8eN3va+Cj4lKNqbqdNaLGOIdbJGB8GxwHmGw1m47KaDtMt2P4IZTPkI
PpzTgl4k1sYZyTqOsIpvr9XEDqYjgbYVPGbrKLfJHbVW649pojz5vfAFETkptfyi
YgnbKL5qPJwBhZ51oEEOXI/WXUUcaCYQKf/GQSkh6N6onfhgNdSH2tbHa1z05MiN
rnCKK2ak3hviX6mJz+tbFrcmTsVKS1PX3n95T+27nthwRK/JOv0ztaD8ZWK+Dlz/
f0f4vgdUl8O0XMNrC25FvuFRM1Lzr+wkZnAq+bWPiWPZ1stTLFLpMXA6mIjKJwRI
yesvrW8y8YVYqB81tPP4WIfddtFQekqWw7jbHsi+eWktalZKEVFgx/7fOC8VrtiK
rFEr+Rr6y9gWAXZW2FJBR8Y/Axl3kzJ6pzC8DTP1Ief/FW4QutQB4ExObEJe1Vxx
/bMfun8OcHH9/1MZuro9w6LCpGhQxhrdYjsHfI9Ld+LOgB0hBwW8gwWrs6M2oD1h
bHP1nwa8vqHFftiBEG7cF9/oHQOn8L95+G7EohKHJKEq2JHQmlyX5qKJowsIhlbL
CRVjRfnoNHYETWsHXCBOk4aQxBl+Q/0qAAHdYXwOUUAislw5L5xr22zN3uGtOuow
ai5anCHsxB3ESvv0YD8LCYxeoiqtcjDpAOsFayF+/LZz28WdBFvcSi660SwwbCC0
LNEkni06LjfZq4oyeCR9umGUAzY9PRgrOhJWBujbxiZrtJYB/FCSZtrzAj5r7gnO
EZEh0Wgix8OYNRs30zaBUui13qkNP74BDVHhGbIGhBU1xd+/g69lMcyfjU6yMF85
DRRzb9DVjgOyDNeAkr9HrcTAo8Yx1zfMivuNjuZt1SCqW7FAxEodyJtW0Oj/8LtO
e1MCXtyhJ+4n0ktHS/RNY18XLWh5JvTKQz/POkTCQ/zGoTdUoKOnK2fJyqh12Ggg
P0YK9CoBIb8Dq1seYwHIqESdocq0AFd0v5nHuybGu7xoQIU79UvqWth0F4Z/kLb6
d2LtVOfOrbf0JmUVnVDzkf/Zpsiz1Of+oK4FB0rC2g5TFxVkC6jV7IP3MoneVId3
AaZ0avVfU3rtFq3kTfnHkM5rk4uCroLozorCjmUS7jLnnFrb3Oqdj5CVndjO/MRc
xO2LgnSiWNEYQGVlsd3GsyDW8clSk+TkwJbOPXX2XQ6MeeO01qQSWKJRgv0QJnCB
o1fuviJbYgkGENIWhVjT/0PgZVHwBnUk/VS6xRr+/FxsM7o06rFOcr4OeSIOuhdG
XWLqu30QXCLBo6Cdhtm/VjEv4pcvu77mFmy3YnF/BWVeP/yVxvvp0H6H2f1VZBpy
KE5W5PGqFtnamIXQXP2rGAprxYqHw6NQFU9tZmYXeqzVVdwZqNPX8nb7uffTWP7J
kpW9JPdo8J6A+PC18B6wxN3DsJDof9Ie45ZbSBJPiP3DGdfXuA9fPV+3DxH3fhfT
CTmuETtZCHebv6HKYOkHWdX/odxM7q4IgCz8Se5NGDISpQL2UA3Sv7g49/fMEpNE
W7+OJSj8/AMjHSoGAfJzs5iTcL3CenvIqLhJV0rqLA2p0cBya8MpBgZ9rx4tznwg
y7JrOfTCzT6dKzYX/N30L0ekxmt0Ht+pXb53BldYM+S9dJ5d7zx/cXjCI3/ir9AD
M1jVrHXQpnWSTWV0GC8IAwZ73eRvZB9WiWentLakiRv285cgy87aKcPOiuw1KA5e
v3Nnm1FwN0wHrIffdlxJh2wib2exz+BOBZSX9WCFsYIwWRLX0jK3R1LLMn4oazQu
4H/GLpkj+826H6nsPVPmXmyG3LCTpxiutTN4Wd26JVUbVthla1ILC5EJcYULHg7Z
4jHAdG8T/5YyxR9bw/EOsQJk5VF/XnA/+Fw8AyXPRwn2ujVZ2HPq/kWOXdLqSCSp
KFlZxqkGjAVe88qW9Czho0Vsdss+756ID7tVUnRfHGxamiGfT+gi407nB8m97ncn
oPhuv3RNlPHuWT5Le2vtj0pSrCeLIQm4L3FW8CXNNJjb+j8E9DczfJoPC7NGQqqB
mpvXAqobeXd+pNkvY6KyrVkv4tNt/IrMeqLwhHwiwEJIeEFXckv3sjVvxFScgsI+
rTTCt34IaMsb3yTYcUZktM3Q1EO4p+TBhLKgta+4cyPbupE60g/HDLBQg5kd84xL
w4FTZeTIHLzDlfs4Y3+YMHR5UfEyPv1vmkLnC7+TwsJY0y5WbvEObsW2E4cND7Ht
o4jWEZVmr835kMhB2bAUIyhXlpQFNxqu/7SqkjZ8k7pFC3lO6GOf9IpDupe7Bs8C
fi2mjm0Uzl2I4UYa7Cvrsg+EtdJEMqOHBJDhjmLnaj4x5hj6oP2Ov+mlXn6wMIX9
cwhySYxsJ2lGXSY8SWG+p2BLwilna6uvK5dx1hJbAtc1g909P0PIv8vKnYpfwPop
vgejE6M8yM9Cig5llxoGLK7vMSyL4Cfc/WnvVM42swG9dINp2YN3Q9uChO7f6D1g
SPV8WOkovXpGv5rs/sXUFycpdb8bDllh/Gw5uT43KMZRs9b0lh+UlvfOW6OYvvdc
RCtG+VJ+oB5w4iksuqOfLLhCG5NJ4P5WBjLC7tc/cwNWdGWISipuIhnN5dfpQE5c
l5p2oUGwL2IEeLv8QPBhhDrf1fefTwXksDEYl9m+FQLcIC01LxgTOB4hwFmGfzyP
zNYDtah40cLRB/VqyST6nGHRxtblINRt1zvplsNYCuBwQJWkCvb71rnn3OWXr30c
o4NFlM98qzqTWYJd2g4RNFc6oHMxKZMQISkUOg4asTprWd5Fii/rMruQp7lcDNw5
WvN1w7kbBJbBuZPw/8p74nHl6bfdAAXHaar8SFWu/Svyc/U3HoKPWLgCVx9Qd3vO
ltX62gVZhFXs5Iw/u18e4dSE8lqq7T8Ou13EGENzMSCbVy3I3+5RgnrsE+tOwUMK
XlWvzOjufja7Vm36El5akitN5PY2IAO56hh/RdgLTc8dbFAOqqpu8wiRd671E5uW
kvIE8+8A8ZE2jE9gNxnZ8b/CGQuSyUD8+QCUMsjCwT0kQ9o9oQEjNTfZzSB8qOmM
Xny/gcRbg/da+Pc8+sn6qB3u6relQJCG6CPfh+i8q2GTqzaGB+jSKwXaHDqTQ9FV
JcD3IOfDxLIXh5eLCXtHcQrrrHaHDNwjl5D9FbTD7trUSISOZBKCiNLDR72gbnfz
MeZmVk5D1cCq1DD6QKT8VrOSnIX07WWpbrIwBsNlJp30kKeNladFfX9GU3jcMhr3
aaea38PtLetbU3wzhAQke+LfYYKEWu27TrfD39SF3h6fGCai5h6bENHlh/Tp1vzr
sg81mYmainWahEMYsv0vdpH88mWKZhQqDNWZ75OJAP/fc14atocAlY6oE4G1SxJp
o4t4n8p1jPPAxRpXWuIQCw4PcZ5nxwlscBmJGF+7C6VXBZ0gb8tVGpBm2PHhUYRP
+lRh2C/zY3fsoRePf5/AnDLWCTY8EElbA2V4q0wvtJbNltd8MvfM8VHQg09mvgFA
SypoVJAl5I54D1yTYAOppyhyKWHYevHagib+EKvNSpYFL70pThIZQBKALocUUWag
FcMcQWoNgMz/zJUaZitsMBwv8sl6wsqOIllsyKYhY5X4+1rIl6x7l73eZse+oXfn
gjP1zdBaJIsrcAMsbIF0z3YWEiSYg14J7tnxbUVazOW0NLT6bnCMRcEHEy8+fCZb
vFyY/0Vc5AoP8Tp9AG+AWnSZ8lVZ33sdt4dlOCQwpNhSjqmLV5PBJPcu26U8PnHO
C+wnZu1924shoibxrEBHE2GHi4hJMTBayvwNnGCebRW7WUc9ys/2HHSeUOkZoOwp
I47/GsMCVKmHY9JXkhrRHf0PclVmM+ea2mgf7eIS/pvj3rwqImh79Ah7sRoGII2u
neHXN3LOsMPypo9JkREjQdTWyUpI+fM8UBZdQdLOevD1Im8B6sDKVZ5pLS3oYmKI
xL2Yl8Ia63faR//08rdSGI0gLPGGPm7TdqsOSRGeVYnhLARDAU4LYFrrVJukY6wz
/KwDTLb0Se4+R1waX57Cf5iwQ107F1u6uOCiL9I4R1SyP8LfwDiczEMCLm2LKaV0
igvdJ3jpNRkj5qrTk5ud+vnJLQgbAQRyatZ4ALWCRuQg7ir6t0S3B6HaOgmVWo5i
yZEnFJHcyjgxSQNpFzNbuqqpTxb3+++2js46o6tiZVk5IuTmWXTiNdPJkarMvsIk
q7Wg5CA0stXCQ9IrjvyAsMCCmzILNHbqktTO6RcWNOb8yRdC3thhOSkkI61GR+1J
JL8espP/18G2IteiLBNtpa5tjNkDg5i3Wfr4JkrnCbRddTiWR3iQSrQaG/nlW0wj
KVCVAD3D/VGHpKnM3Y+/NYFaS8jWmbxlqewZKXxZcckJSqZxt3yDPTcRkicAToeD
uKlcIUhBVRWWVQriC+XI2lId0tubQjsDCYMpfbIw/X8wyS9RbfV2JqZPMrgnSeuB
eLdoatmuQJ4Mair7GnpGwwL8Z/gDPRaW3CX1ReHTyFLZqT4VXXNOAgw9Wg4wwHwn
HPtDKZm58YvVPM+21TDh1cKrl48SfwPy03ZDglpTbyWZ/AOdMuDgNEGPJm/hlDje
JMxQIfmgYndPNYNo6aWAgeUJGJcHi7Pt7atXuAdYFYJF57b5/W790zgyhrT55IGm
rsIav4NB2usLmhxqAN1TS7yAgfx1sLDWxk47YDx5bIRCeQQ8LXPJHzUyLeiOFYWc
7KJupZE71m3oVWepugxgF8I6FA0gum0n2A1UrUmpwR+IjnwVV1kBierT/9cPRxQx
oJDibXy0v/TyDQJ1V0xUjEvdvLmizjoaGP8S1GGoXQsL2TYrZONQfuyH0KgjWX9K
UsOoBR/HhnP093BeYXqGvmq9fmUkncF9fwXTGJ9siPteI+4ZsWqv/eXeKDsnRej1
AhsIv+dWHIDOZlsrCEA4oER1Qf63N2Bugg+WcWWwn/NLlDL0JGsYX43Ri6cU7qDS
8dvkAR7Oec5vyAi6rGn6j0LBMjYd1rONTp4i3GLrkopf0dnHcDMaGGhjmbpG3UX/
O/qK1SpM+9703XJaazi/17jrIgcnP0ZrPSVIctCN8psmp50jN8mQDDWChTJLVeTC
AVYDp//gdt91XoiSOLOTGapq3nGLmknB/Qf8I/PCgpMtnG0Aj1O2C5lR97cAEgTu
vT1Md76STW96KLXuYozbxcXf5O5EiXlkPEjhGtfiY71EVJxFeowHQocMAhQjUGOO
pQ7YbJhUxP0I5toivtQItbEERpVYyVfGzGWCfkDJo+1iq/qECd+2+JMl12392ykv
9EiglNIwCPJcbp5pKpd9tlN5pL7XU1dG8D2Fx1xKl/pCsJ9Iyl6JvchK4f3OL4GD
7hyU1kOW8L0s/FSBFrknBbRf07gnZQjy4dTz6Mq2ETGDh2i86KWc22AL5cS7pK1u
xFL7MuFEiWHgLFDJyP3/jP5XOrgPJq3D2kqA9b/YR6djKwdtSQTEZ94QpuvfpaIw
YuClves916S+9OAv3xbNUX+aHocjwE/mlJy9Ky0VrbsZijctcwghPMP0kJg+vV33
gR6rxIsG36wSPJp0xlkGGOhPiF3r3Djd6+ZpyU1kCzL2A6sjn4dWxMsmrgqrQ6Mg
eZ5p9Q5lq6DXS2v6gN6m7hqqV9J89eKgASU6QbKKEZqOCdN5NVeiwQXlvkSdZQcu
9YkX6T2VAFRTwpGsH21wVxvgiY8aKlrLSYSuBOxROUZm9Gv4y07VR1UOcymt3niD
uzuHQ9kkKIJ7/WZknIn9u4CiqCS6DRG/BiYFrCQdrOOQGwVMYRD0zYymrcFO1kw/
g/fLfMdrDT7usI2x7T0hQKb1ds+LWjkm2AK+2mH//Mpw0CljOTAPxF7l7Bceiq3W
4soJnWY1NTqhO/5/gN3i/L0D9Vqv+0zXZi8oL/mLrM8GuZ0ssaYJw+RED44aTi0/
UODa123wnQmJO0rnHDup/BvrcteIRi+5IaUGayZND644FNeV22QV9HnV9708xjDo
rEYObesVLgDX/xPM2+AmHSf6VpGlntIimtETBnkzfge3cEbJ6+25VzM/ZGVy1dq1
ZTKFQYuIGuQqvoVHzCJvquVaTJr06X03ZkKnoTzHMlQRvpwSsJGZyfr9SlmAOFcW
UYyNdUUVJFj1jXuhI2HTcQC/H0kS0U7FbU7n8aB1swEKQsgAoQbD3u3OedrzUXVT
yr5xZ3RAr3tM20nowQru0tA1fJ6SQqNTpDpepqU+Ffa7aBPypqpxuA7xFRoYx6Gq
sy6ksCLTturJ8B2DAIMnMgpjGYZq1OphLT2HcbfJzgUKlFTEP03BncBenF5f+uYz
rAsgBxsDgIOm35WpYUAHikbyvUjjpvs4ueBLSqEHdi5TZ+6skD0NTmqTe5asP9jH
1q/HqT2/x3iqrTozhDDoKI6t1I0ZWoJHE5i5T81WY413VNTeqinkk4QWf5FtL5ji
YXxm8gJhF7DI9nw0XVdfwZtGxJVao3uYi1Zn+lko7NKUU7W6TkxITnwqy2Zp9FZC
WWl39iki2aLBZJYTwlsElX+ebeKXIiix2WoUIs+btQNHvZE0AAHrA1+hRn/VvSW4
fiM9mS0LDnQZtb57WRQ5p+4tw6aVsQ9xpbwejP74Z24WlWx3+T5LSm/ryB37+gfu
QVIGqfW9SH8BOFlS8gFE7URzmU6lLQ1ZPPlrqNGD3+aFlyqK1xdB+QQJfhQQOYAx
ueBjyfvOnhxSd5fV25Mi8b4uGEgGUTDxftNpYBIoqJ9owe81qZEXctL8HDFCMEwf
Pxk4qKucd1y966vs/Z5fPoWBAyX+ltFLH+PlBzOPbCuJuEppY7k+wCGZgbNqsYAW
TKzs5yCVM/ZXNj7a6cliDSs124SQ/NDzud/pDGC40rIN0AjA7SUuz0CgxfA/XUY+
XHuInMWbEuU96a1RAMIOqC74rXYle/6D1OzuQ1S0kZq5Qv5OUroROztct9+YcFQQ
Lh6IDwybe6xMuuQmDKEIVdjHauVdEFacFsBb0U3PNRcilSnulUh5UWcsfBURMfgy
DjnU1GcgqRVUQQx8jCViE/s/nzJXKtyEy2whYgya6UPKQ4sp6wkveIMSIzVRpjoy
WT/2pEHmGFTGyj13K9OgI3vZZbmtxLqyaR/v5V9iRM0E5YxMBcjXMEv5F6sKYBXu
ucsoTwQtXd/1rWhxx8cC3L+TplxkNKABBMx2ynLwOLHlDD1PixgOQ7K4srzBbWnS
PSrb6elzDyMdGAkvAVWZ6me8hcwCwhFb7oTLTx2HhDD5B0dVRxApfes12DmEYpfM
4SkcNlrlntAgS0UTg7N76Ei6ifaTU6Lp1HUNhnYCA7ZuvddjKBKEBiHxPVj6amRY
DGT8XepRL95SlPuW+7oqLaQOGIq5GFINVdA8WonjCq32a36qGxMw6d7l4LgKVNu3
mzOWbuU5LxFEO/0z+JawzrLgAgMi0LtMOe9D7ItW0Oy4VCEOV02Tju7xyKfl8DmD
s+cMuQxiwCdd7Jwcg8TauSZvGRR2T1JNH5XMJQrcQ/yg8MUESpl+485NtWNd4kWA
jLcoxlKx7cjv3yEazd/kvhTjJ5maV7Zn/g8EiaBdVWleUMWOoT7kbLtHPA6K/Yeu
eRTNEqJ9bP9jcQCRRGPivxa4vTqmAhlkTtmRhbPGbe0//iMTtkE+8SFSx9/5+Vid
ucm4z/8TIKLSQ0q5VK6xo/v3ka26DQsppU8Zd9tUl1S4nVTbq+X3YT62H5+yaDPh
0GkZcNrnsLt9NdSNrzgggz1029BKrOv+vXFPeK6kZpKirvFtpkWWlFn/G2Ub+3fW
bps457AjfcljdlpePp/Opu2+qfPKghgselDc70nXifK14Y85PQNuxDNQ6lFWtlfv
WV8teLF9LzRgdRXUDGafzoghVO+gN6XnXI4P02C3kQwm5VQC8sE86kYMc0VuwyDA
J23x65UiTOEb4zhh1DyW1a7C5VzmsjcYqc5hfoZ5c6aDIAcIPht5E8ePCJ2F8nF2
lyTQbvOMNel9uppDhGEupFT/UDasgiE0rva4g3Hin/k7mVFlWLoYMz5IeEkfRR/9
bF1EoTJNqHP/mRDT3050prob2ag5c4VrDQjgzQ3WyXjoLtV6cE8g4Gehjp9pcf+l
lSR1+L/VcwSFWsyBifj8DN2k3v8ne8JsPhZcd/La+dedKgMONp0k0Wi9ebMFXKPN
0T7Dr0BSNh4PMeSjMDkw9ZJ85qkbRMGcQqg3OzaEXEBz0OEkfx4YUXCSmTBHN4eV
zKljws3Hwbtnx53SP5QHIFUkFwOiGZS5yfLzuQCHg8/EWvtLFdkV8cXRKGjMsXv7
8phRLpAM4xP04Kd0WeOOjxt63kF+Zv1onH1r2vrJmcKxL7fbgqRq+ScQAV110m6I
oZDOV4W2Em5fIQ7N4TvenfFfbMSzAIgcpEVIBFJcO+9ClS7EDdIt1L1vnzxFchZF
PnmPN3XTPhvYlRG+PtKEYl8qhtKRuWT3x2NdLRTLKqtE0kF2bWwZaCvTqCRXq5r5
0FR8d17r+lHVf4HWwCWiKIy2oXoUZwuWwtEjYEtTo3d+gjLuYtmoU0+arB4APzl6
rH/g9umzAMxlyFpZc4FhFBMuMR2LatyTX33LQFYT1emk8jS7cvSM3KuZDMZSsRf0
WUwPg3Bw847ai6B00Mf7ewyWpZygsepivPC5ewB5ZwyWRNl2onxpLQaSNC3G10Bw
+UPOTxjSd8KoTjo1VTPBkqL6qu4zQFieGxkSb+qzhqLB/IKhjfJ85Oe3ksY5JM2u
9AIYPviacafxbHdoooWl+okKYSF+LmCtn6b4s6SEt66HuOQXMfslCVtC0QrnA0Ys
fcwj/MDv0Mvh253OWxk7wGbpyITZw2xmJp3K9cY0hlpneM40+jXpxEASf++HSKku
SK9yARrLITEtkiaAbBpNuP6mTqU3X6+aTc/LAKaS0/BMRhtcMfMVgRBT/skvQihW
zh91DTUGJVcmNEn68bAT0sCE3pc2dXRgEun2bCNnNw/3QqeyPoKZEBG9T3zH2lUe
xJm4SNGKHHp961vTNB/gx7tbIvFI60qXVLZYHcOfBAcaUu9xbxxrwZ2Fk37GAtKf
k6fFV8W1CopTv+BvjNL9eGGcDGsL3/YRgxORCeX/ct++f3fXfTI0K3cUfT6IaG1z
36Om5QZMcq70VQbZE4oZrHvtiUuQNixCoHVmBMuNzZpNB0oec/PmFPvN4XUjY+7m
smannXQ7ImUyRvlIVU+WM7qMqrdSIu0IpEM8EnMVZ1TldHiVucwUuHOtCn1AT5nC
4ULwH+tqoa55uh1AJ3nzd/3xisbxxKuJukl2AnM55QXOY6sYk7zm0FmwztZ07Yrr
YFWYr1fYYYbYb1U9uoaKnok5Fxo3vv3SH0pxYQ5hn+q9ujZHwvXvWEcOXtflVVrD
EMLjc3svn5nVF7sKBhhaoUnDzq9eJ3L41eXuqf2iyuUKlmHpEnoDW0YOkHQrIezN
sSRtbmuiOoPtUd+Mbpf9XeiOiC4fAgWmNsMQi/M9fMzdTIGIS7Cp5fvJ0Vx82hQD
IXRy5Ep8cGYd7us5ynTk/uAO0BeI8Pig4H1ZcyBa+8B94vAWnWS7ymRgC1SdMGl+
cp8V/Xt/rXcrkj/KfRb6jRneIbuofLztXjFn7F4u5uDLWh1DDjOSZLQwMA7c17BP
/Q/N39POToCgEdo0Z4UMqrP1+0NW1R3MaNq7Y/7/ne0gZ53b/K3qJmR7QF0GByvu
eDNPoFGTJ9JaspyTSUE4MZRqawdzayJEy1dgoTsmWoiGtPo24AP1uhDqPBeHU2tn
EmtFkg3KQt2V/rvCty3FpWo5l75REZQnN0V8mxTYPolCf4V2R34kn0hXILPlobnX
i1GLLMPvrrSUQT6opg9Cy+xOxkWGf+4DyegskyQeMZ+OreR6HbbFnFsnxcUlQYGB
iHZlny0XchKsdfJcLwIkJk8MIp5oUVzes2X1HAtxlFtEaz8axcEEanXJNKHpi+bg
GGruMHvMAy7Vb820lXh00RLZso843pUzXprgQRxFHh7W08iCnMd2bwKlc/5unnii
SX+oaCryqda7Qd+YFQeZo7Ynap/RXnuYHmn7zkHP+4nSPXpsjCWHqpnUDEmg0fZU
bUvsr0FGAyhQE7BmacZz0CA2tF6gmyuENVV+UwZMQ9aHNdJeLvQhyEl9SZkNzwg2
FF4b36pplUFFsT37Uw/qYsAbfIs6cE8rDBiAhoWyFz3vX8sooqMqaqc9arQF+UAF
LDgGulxKUqOnn3WjXdWenbOHtBel6Ms61FGFmK1WDp74l3ZwwG6m6On9k2NwMOV1
RQrcDS97VPJt5rhqqBO6DMQdEWOJcCMZp0LpcHP9cP2C1Ck3d+VK1/VvnLLRKCPT
efsmsRuqtUNJtv0JjxMo9Yu40H01JAXNRyYKbAMY+HZSHo2NRhFuNzwbKZ+t6/je
sFbR6HKrREYNzSeBZ3yXkavb4OlIV7c2pVSQin/ZncEPO93F7ADumwWi1F+adn5z
ZkiK4m92febpYMV14D9EGMU/OkIhM/NquSDxKApgOSSAphjVDdshtGyc8Fpydkip
SAtrombRUQuE+QBGdpwZ7lMKrRQl57E0D0sT0LcGkEY5vcZhoIeW286oNCgHN3Gg
JrX79XLamMudJ4B/71v1RQPxU+rt71D0sYMsGUDi0W3tLerndqf6R4W1xbK5MOug
hGFA4OYNLMWveY0yZ4u94ycquuoK0ZrdZk5UFwvP/jdlPFsGkusWF9ZW5hnC6FmY
WIlEkhIDaLp2ma+ylF/1pXpi6TOIDG+6geKTQz+c04POUt2gHXr8GqUD4PPP/j8D
8anMvlK2z8xdh1PuI2CgW4BUIkL2jAf4JYponxKVIY4RSFctonP/h/Iv6RmeRhkO
kIYdwqi9+IwN/eW+bg4DOzNkhio3uyyE4jAArDGONoCWEq/3V/4ErM8o6TGG+Ui6
YO3DlrIx7FE+BihOKnawBt1ub1TKHLBSk9PYZ6ZtA3L7IgGKUBLLGFwOAIizsCuD
pcduQp7nni0YQT3QRKwrtCdrVxbs1rh/6nmyKai+uAfi0hpIbRDnbdgO4FQfkPbQ
rBJWW1U2/BOHi70bDBwvAvoFJNIkL59e+AyR2+dWEuLNvACKkoYEAnI9sLAYi1/g
qHH89IJH/AerZfxLp9SGiIUdaIzymI3Aa8NSnwEPpdltC/gfJBLLHqVf9+Muo8Po
gEpzVKj6lZkQ9QY1873ZCRgB0WS/+NFW9t/I4OuauCM5TKE5xjYcbKTRU/CbI0s6
fLn/DgL12gA3W572bvxR7MpOLjm1GAK+/LvhCnmeINEL3yAua/TifRdtZa0xMlwT
qreyFs7kXGMSBog0PLhvqPi4+4MgXEi51D8pO03kmW01R60tY9zE8h2qC3vkVlGj
MkFTi1LIf7YFHiVPmWEXPcJCpz793Qk9n8oKq+V4LLC+cQNkBRRakaYrGW06YQvL
o7xR0r0FzdpjjBOMCO/rmvVgm1FHa2Z/sY2Oyesdf9X42sVkEc5IoocM1J9vgqRD
b5jfEctaQogMqse5qVl0UQZwlnJoAfECvKTDxvc/j76ID6mXRUS6muBN1kLRjI8w
uimaSlWsyTndJGlxtZD2DuNDhIJM+DkqD9JwH3i3O1jV6b5jmgXtYicZsjPLnecR
+WHv+KrcTnw7sb5Gvy+AYcq+3e8kDEwybsZSUdb76Ak9a8DdrmZpSL3QOujJ/UBY
OaybG1fD+4SEHiXP2sIEyZRL5VSL95RuvzxR/TkoFvuk4w5sLKibHWKkV+hEVjgG
zoj251KjN7V0fbezL9S6f8vjsRtG9BN6uyZIfvGnV8ROFdddn+02Z1npAJUn670T
z5G47NV4N1oPqwi0zEApRCT+ZexkDiCDa3wvwF1BrMUcGQbVRywl3v7dDl5KV3ZC
8B+brOWHrjciZuH3YDsfZJ+D9wyVyLL9S0I6DgeGUeZp3M2mP/BtPdXj/4fsdZ00
wRb72tCSKVCFuePaZAZoO51TiEWt4cnjSMkloRm6zk2pYJNEgX22DkOUG3WIc+ol
liGjGoHS2lBoJOuNqHvGbVw3pveeu89GI5J2dNbsCMGXM2dEoz5n2R/k/AXTg6dS
7sj6frowSUNTc8hlYxxHL8Uo3RHe4F6Z/WSreuhYB51gjcz0XiWi25Lob7MM9SrU
ER8tir2yl5weJ/YXcyf7hWU2GQ6wi5lCCotxNAjbxFRLJivypERHBmwc1n4esEdJ
0cK/esFMsYalZqllJWGPFhVkt2qb8q7nHwGkC2lgZTqbjnft/tHRpHxkPZcyf0uo
LCv9NzMLYqhmmt55Hg5KGHXvvLeHFNxTvF8GbLclrihEcQCuFI6FozcLg/jcMIcf
R10VcesuY1eRaGMbSB9ThfcYCEhctgs9AtWnBmKy6Ce4DcdRkSfVOWYD1HVGiAhR
Y2akjx763ekuwK+39F3x2GOmmPbT1MBxImwi/HzcutePiZloAfU7pTMh2UZwPTvo
Yezru+JxQdoQSxohl9K/xmBHwLrhihvENKTvo9sh51cwC1F4IxQchUog1kao+gz5
sA4fVkxOdKVYC9A83ebSpqYJp0iO/mde0MMS4j5REzO1RLTZc5GnTLAf0j4psSUB
jtSCfL+vKAwIXijldZCfw62p4fp5AkGXPOU7oMUFkVRNm/lHUc+DjjO2y78ks74L
lJ7zHL3fyh5b9oCivEVdd1wHKelgSC1/2wvcz3PElpU49/DsGxYpNWxtP9Ozs/ya
Ul65rCw3P1vk0sSOcH+En6Ji1OUHFVro0XClM45DGTc03TFNvr8WuXrCcf/6gFau
NyU6I1lRwW/O8MML0kCnhmZXzTreNm9mPMatIo3xDzG6MO7+eggQqj6KVq5vlMhf
cAFQSfA1+kBKwPbcW36421dQdkaPAnBVlkVr14APLxvQud5HpUk9AiUVrlBS61qx
H0tisvaIX8jLld3L0M4asofwMfa+EzdhZTMIm6g/L5AVLxfjKC1Z6Kq3O82sqZc8
VkL9pGZzcX4XS50zWymAfnvjhnZF2+yzGpP7k5p6Qza4bHhwgVTpcP79wfi1Fx6E
qTwaKeEAZ7ePNAN2dFHI0YLvGAof9z3iQlQbZLO/bc6ZSOJeo/L3A5hsRy+Yccmb
1lvsII41LMe+Rd4jFbYdSwf5gaYXcwwatfScfiilkR7mQKVOynNAOUuK/v0x2RfQ
+Bj2ckRE52euIXri/sJ3yvZSNK0uojHe9uKokwcQN6ZguhtCyldAGjdffjW6iPA0
vHI//9WDbSUap8kT+E8mNtC7+DPK4IcVrDThFglpkBgLRwS6CGeIx3OmyHrQhb4e
3ZOEkeFGgyPtKn1qz1LBs3c7/jKQtR3vCKozWfBp6QdED1NKSRh+JjRXkZAvCZ4C
7z3td9YDaMwoEyCoIIh46EMUSF/nNsIOKASTucANmHlzt6/M0ngiY7dz0gDqh7ze
SGf65pU0lF/k9znEJi8tyBUdOV2YK2CWfASibudlICRvJ735e/NaDbBo+O+N17qi
L+0knC1GVQsqyfTTeSGkzOJq3dP5jOunOEH1lw54aOIbWOUY9iIFVA3ppxiX6LHm
+iev1Qdy5g4Y5lAMS3KW8Da+kzJ4CTiuw8+TwUVWvAfIIuEcMZYWHe8WL+r5Xjwp
fOD+W8dgKt1ii86TsSuNct7ogALoa4uXYHJxup18Zqxnsq9Sx80DgpTHUFyP/puT
z9NzFI1wNZk4Rh8vYOhtsOrrGxOeHo0rcW6GyAqpNIg4jVr2aVh+uEJtzvXzbrIv
uqwc/VpXu1tFzJ2UUSDtyP9dbLPTjKbPRZ2THsY5Xt3xlKlX3uB3lmbWnNP/kZ2k
jA19P/jzyOmJFYcTNAHmVvB6aBnJp3boiPi69VBvJkuCx28NUp3zIzgIwGP6h5AP
ggw/BfKRQ0RsmL4HoXypI4AIMVtdnIEMKJqIkno+j57Z2r4XlNHn+yr8aj1chBfV
ckimL+aOpo9Ds0glR5y6PClMj58hNdk/6M5mgyvzeSMvam7AV/hVw4GMuGV0hKIH
J0oVnS0N4Atop9WWuMRjfHxdMhd7AJDUeU3uGqmLZVqCdHnYUPcz+8i4924AMIvl
iO43cx9sKAu2Jkpe400ccAhae9TCrZg6pOcrwxhn02SIUNQeyv3SzyMGOxfHvJ9C
iJdfA9xsgixp0mDbupQ4wS4MoHjiYIu2gZGJ18FuIYcepIWc0YH9G0v50Bd2TLbT
P3GTvh4Mp1bcw866QEerur2rI6i01cW4sBumceqfVYolgacoiL/qncgs8RoC0jW2
CBfWXasNMitLnG1l20KZWNk+vvK7IhL9pP10G6KfmB63BHpwVAgYsNAkjy/CXb45
EFT/UQJYYTLKRsEmTzQZmaH70e/JtFT7zWv6CyqZTW1y5kgYZAAuFuEZWHENyl8s
6nXG+pMav/K8eu1Kl4dhzxtgeiEU99NyhwUI5P8aGALDKeO5YyZDpznz4Ye2AW/I
yqHFgQklMdNVZEfs7PWADxuhwNi4UufcZURUwQ8+2RYudLQm7nXQ3Zb9lJ1j5pjd
0e19JOpOdK5ztiON3/x8mGVj+0X7vQ7iiCSB+8RqX2J5tMMo9Pq7re6WxV2EDx/O
18uceji2BKbzg99MhuWv2ng0Frup0NOxQ4SGnphwV+hk+37aBSIsxAJNO0Yc1kh5
CCOzr9R5YNMuEwR4pTc9+ajEu5l3NaSR6YpWzpt69nZDz+YBUkJ17n7aFsy4bkm/
lY65Tsmfbnx16N9FT+R+tA27msYhFlG1ggqn/6vF/GjXqQBXYe+cqSedEtjlGClW
mSHa/J1LRMdditsKVifIEaSLvL/2amJ/aRNLOPNZd/ywa3PsvLWhw3k36WFukVwQ
85XxppxEZwjKdfuEaszIM3iqfbVZYwoXGLc6P3J+VD113mnMv/Wo63S9IyajR7I5
DHBYYqyKsNkFUgSly9enEx4TN4GQeuItBTFPtnlvIwTI7sBXStYulDHrIqcBi7Mb
jINv+Fv2ceXxTrtkmwNEw2SfHs79aSvCRiW0X8HoWkG8Ou9lc5OmYoHhyujdaHQu
IuJU35q5BWM2TU2Ru8QHpgrpngG4LKn3XDgYBuW1hu3D4qwDWcLMIZ1JpnwWT//d
cI1CkPoyCPt7/FoOBc/RMBYsUdUiG4PpshQWxl+i2FG0FluN2txAHR63vm4OYQ7z
bz0e8TT03vc1jzXFIQq939pCBrkQFe9yeclkOpd8Vd8BylCgxh2GoyglCqYYlVN5
lC+X2x093PNLCqKDNDHdGrBtWF1hUa/JXO/6pgsVwFEgqbNKxPyn7EAgD28IaX53
p18iM0KIlznU+Utr0mWUS12OH0GwyOIiCZFncE6iLunsavCyYtY5h4yAbRUBqBh7
L4N/utUSbatOPQ4Yj/3Ao+WfgzHa/VbFVht7/4IQX1c3p/Sm5nx0ePAvvmSV3/1x
ZWo7I02oT6LBvdobFPSWWPiu3jTIc5UK94YFg2n9p0fMECZG20hJ4w8UHvXR+DAt
scSfQlqj7zCDpj8CpWRPGTAME+97Nuc8uY5lBMQq8E8ifB5Q0z+chTDtDsO8RjvU
6Ato01I42kL7KrxI2IcG68px38IeRTMM+Zp0SNJyDST9/Ep6rV+IKzUEed3SamSo
B1PH2vMaY8Wky9rA2u23EcVnGMViosG8iRCIUUp1h6vWeEqleF5AWwic+H4QFpQe
1HQu1ahvhsNU/clDYT82k/oWITKNxXHiXahK8y4rwstQ+CvC6b5JCI+XVQL+JQdX
oHaAg3X5fpdTUMaskVKkqYQ63iiqJfpOzhDgqqNYb87ZozzdVQ6qHajhbjE2JWXQ
vr8L5eHQHisFUlcMwC+dls6syYgBfvseyAx7LI918v1rcsJViZFXNX3pBNOlxOGc
nDQ4iafI5QkMiXzIqT+1LYJMrdAFT1G7LPcjtE8rbsRXiL9E5GDRakjUBCYicmy3
oJU+gLYXY6mORDBAt81thgjSYH9sP/ioBAtJfpRSgfkb0eHLx1fwqiL8MeFoFa+e
H/UnF411lgC2/ZrK2lRJaR1Pp/nWIrt15FtLWRZVhq8eAw9pGozNqzB4Nhhv+VX5
/h9G3SoCQieFa2WrXBjCyk6abmIuTijm3dfbo0J72XWVGUM6YWBt92ILPCGa1kH2
ID5rurmpGYoT6Y5koQ7A8YBxwIhQN0SMvxpa38yJ/I0YElpYhy2XUYcpfV1B2SKm
dTZs4h4EA0l4F7M/LP6xQlwoe2mPkZyD04ZUmPKjuF3KYKhMOi+MdFsnpXMrMuw4
BSgYrQgu/jSIFXgYumj7nDfOYmp+vbqgKBKmAQiirdspTxGh0dmzJYAs0hPZTV9u
L8RtU9RSudNhqvWhiex3xXDeasYLgL6BywKnCx3r3rBUxagMqkPiCsYVayNigtti
rQpcffStDGNV6SwCdmeysfgpZbTrTRxWcE2BeEt+9r9D9IKeAJ20gLDayeapKaFl
MzjZJQnkgxQY/S43JoJfX9HCN/aT+oNAzID9AJ6wi9xpptC+nZO4X9K1TkxZ9WeT
6UGhGwitH9SrEiKV5gngSeG7z2NcFuJmhVZZG28Ix4qL8pWnlWFfhRHOwFn4uzdD
7QRUSWewn7ovYKV8L7HD3pq6mVGHGE8NQoVxcX6XOq/9I+XR/hlOy/Xayx0dIrgG
CieDmIiYzfM8rdMuTkNjMOglKMrfoh177JbugbwKXDU9Nu3XtuDsRYku1B4h6iFt
q1pNc2ghb0ouMroc9czELBt6U5rgsG0sw3zzDUH9PsAGt9u37yMDSVzlKh6at7nF
fovWQsETJ3yU/dYC60vqd/TM91jYrwGiToayskXYt8tVVNcqT94qEDW9hMynBrkA
EvCsZ3CRgx6LtrrUh46rpeWjQtItf/Qvo7cKJeAp59KuThWyZSL2l+V7wIiKodeE
r/6KdJJVG0ImBTW5W8+JwK5g5XrJNovp6zZWGAQz++GrbNiolRykI2oz0ZIXRl4W
cguLgRVIXlEBt1IQsPVxlE7UnORrK96AVp80iof++DIuOr9HqMFsgf+nyqXZChc0
FEp0QkhfscKd2i8Y5KCqWFKc+2LhVMmxxorRO+Db0dvehgW7OVjNyIIFs5I6kuu2
Q4QtE5p0xmtwVVZE+//HiNsfwCH3oR6hwm1qogS2GYtAmgDWxIQJG1/+GfgZ5/Sn
Bf48CvwTxkaHGfWLdOIvTJGinyj74Dh7i/1a+wmIy71DPmxWIPJWngLLWfa5BoIS
QF9DGn7QY5Sgh2dqt/nnLvziOb8YKpRnlAIvg3WT2WnQII1jp6KjV4LmZ7ioENr3
ytuFXaGRy+Q6GicFnhQVVV+nVr4xi9xgqX8K6nanhy5+vTKOTvG8sIRxaHGn0PN0
ppS8iGLy14B8/O5UpytL9hzdd8cfkWKJGw2Sl+4wx9oSB/7URf5irqO+WXJCcMzF
kRImo3mLnoL8/zhtzkVfD1RNv2HIgjEaz8J75wTmryD9zwA9GeMcTC6pFfJc+r4j
ptu5BQrBcOv1mzAJNLvEM6HlLa8UhSeY7pTrntU86zrGSJr1xjafrvUrgm+MV7X1
zPTuFQfgKCvkwlftEm85FsosatlYXpK7F9rM9qGPvxdyQgp9H2flvBgfmZk33T4r
ok+jYSEp7RcPMuC2uDG8FpUsjOQPJ1mw4XcxzAupE2/YMIMeiYEBoNWjqGS14tUC
DJAT7EAX3eXdsAm2v9PvfK0eEt0Y/tiEjOj3gZ6HIw8cU2+meBoc1ZSfJ53L6bdW
mx6lIYhI+GJlPVmheBZXUVwxh6KdBGTYKhs16yvMwKVMIB29/qIP9BM/2ZG9GnpY
GXDp8kQkYGbD73frJeUHJdWSWdtwP8Z6B/xBq/Dtu8uay9sLbyd683f9lezp+SXA
5BI+putkwAmP6HJUTRc93sswA2wRwnC3Zij+hd8IYqfPbABHTB1tUeiGePVG02QS
9asaoElFnUB2ZDqBxnyYGHe7agca4Ryu06mkn3Bl6WjzjQHk8qxz04FmkdbeTkBn
8ght8hvt/qDggWPSOYXxm2o+gLCULat/Qzk3NPwxlPqk/ZSwVBKMsoIyXgPCIBGk
ulFFKTIh8oSaXdYu9AKpDFByM8iELDpBR619OqQpix1uTHgpu8YjmYexfByUG4Bx
nD9g666WVzP4Uug3aHCQnw8T1Df6Fo8kvc8zaEycL/uT+E24OvhamQ4//skLsuXL
q8nAu5fVCVrS+KQ4zn8S5MoSW9y/yvOqKXUST24h7Qh5uFGkwCkIlDUGGQYEYHYZ
vdl9CCA9FIOwaZzSZV6aoPy53Im4/myZ/bA9TcOi96aJ7hFiulrSjVY2me6AOmez
20go7tTWg1w+h7fvItHPfBdoual3znBssMePTigcERlLWwtZjCJgOJMz/QEkH+b8
gHrD74Cw4fNsOnWrhfjkmSNcQFB/vbjcgptBxor3XgWHViMIVR8yF1BtFn/O2Gsd
DWiegOGQ/GTFpjjcEqOBNJvZVK7cA4smVnRslSlnm/v/IRdXrbc1SmzsQW+KGMCP
ID34DhrMz1SrWpdMrEiL+gjkrfkW0H2RxGF0RCQ7y+8BrA58d2wZDWNqQR2Dwyvs
S18aTkR4Zp4089PwHafb2Uqrb1uw251jHjENoYp4Fnl5nujX1eRQj4Hi8HGgKRCa
kyCNdLydEBYJ959CkinBbQPLwSZTyOBRXro5717HvNgDiWv66yCoNIUByVRnxtJZ
HAmFjqJB+d13ErS4xdwMNNVLz2PXZ11ZnIe1/illRtGkZGBKp5W75PRaMKX9FbRN
OqgUuinsiHhCOruWKo033Hz9JU/pgxJ3ER1G3+kGK3II+hxwMxf77qZ6ZqZwkicY
jivZ6NoqFRj6srJebfLXzJ2AgfqbkldxX4fpNYmmP5yfZvNTLtdKVU7E+gnIJzX2
qck28roDPDr9S1BEluJbn4kHt67ORD/aKlThite1/XKH1p95MvP1JCVucL3UCrvC
mR9HcLgmxLywMpWzj4Sbn3Ld8IQg3COL0fSemb4g9gzj4N2SB/lOHuMe8d0ofTtf
W36ZfqbP4fghvzZjCrJN5w+aWyZ3xB838NdqPglDnSXPlFn7GIATM6xG0umJb+Ca
H30W/9dSSbFrGfiNR4gjVzekXxeX46XSiOcNoeU8q/4y0ryNgbkY7633Ri6Nvtz6
TM01GOpoTKUBVB88eUYLLTLcgLCIOBD6dCfmDwz+HRGj9fZe01X8Abq0+517846d
plcOoJ1fi2KdPzjdpgWXzdySQm3mnAx63zpPi5BaxgaTrf6q+lxrb0m4f10GeJWf
Phlj7wah0Detd2GIyYqvTMWwFYH3Wbpsb1Ehal40k9QxMisfmJTUVsfAyOxxH6u1
W7DsO05rbGEoINFJxStW5lfqxCOGPVx63UYIkafBVQmz6j7cOnnxyetUylhl6M27
4bFYgK691YgcmN5IaGbnL02dOk0hEDUamO/E6LYB5l67R0PZLzfI8mp4Y9jgDf1V
RZEQSlosP9NeOrgfMat5Z/ETuRovwTnxLBwwl0YecaOz92+IL290Krl+SPmlRdVP
EC1nfjjoevSTVYdeGgLGOr+C6heatgFnLxBNkAvif9Q2jSTFdgVTRudEjompmQOI
q8ytddJERk9cwged14eFUSsTOvf/oxcJ6YEoZML0PVRNMcFRvPFqQCb767RTaDTN
tAVmxjIivRkKNe82FDadYPBs0JM1bMJze2OC4GH8bym9KwVjJ3iSbC86YEvs7WCC
je5Hj7Cd2YithRXyD++N0T5Kztrv6Fr+uwen5qi4XRy6zoblNdLZuaj/2F6MThx2
hYtMSUhwJFIOBdu5eXN1IyKGNATYq+cEMZucKxcP+DPQr/0q9kzXs+zsEhnltPrr
caPaIgWbUDFOgtHjD85rVlbFbeT5HTwSqP1BxDLD7zhwxEhGxOhNtWtukk65KdGG
U6VOqj1Xcjoy5rnm4lW3A9gUazLV+YA0mXwmEQSupG9XuufjXojO8WPzmlPUzS/e
0aeg5LWRqvUytXNKWdXizmDVbl/UnFomn290+Oa3YBq0hajQuVRuKdjbUaDBUAiZ
K7ZGhkW5xVkdA1u6NHiNMB1VKfYmvxX/y5zk65Vdr0wztWOgm2Of8aOopQ+jfmod
JXEA4ROu0B9vECDgc6GZ31EXi6emsp4mfWgqNdYSRNFVnG3MkoNnyNlX8+PTSHxG
ntZ47DSC5HEj9R3QejWB/AAoKQf5/KuM8hK/6n+Uj12FO5kb6py7UdKrYfgraZpk
WXcg1orAH3/JeJloMnwF+FO0W4kX0Xpasildx5XcpIQ2wBd/fBdpRe8piep6nBkf
bsdFBnaS01nKVMe1Iv6vVrYgvDBhJGhsSeUuKafgH77td7nY36RGZuYGJhOCXvEs
YUjF5M8Mzdxk9CRn4oGXqDQ4J4e0D0kDolhz4FhEzJx4q3zSpO3ueQKWei2IdYCU
uIA8ZgVEHLTPZvDynew0L4Dl5p1QuFSW/xtEQqNPSdxUOAlkVaZ4yv3/O/tTIpM1
OY1TCFSseksc00O3pegNc/zC5JSVzPT04eHh4rPyQxisfA8c+iaZXo8p0k2ewF7c
xdMlYq7NQbJ9bAoMXjbHKzUtKAMcM5l0q6W5zfixRzmDZTKTQkfSuraKf46xmrDg
51ewsMH9bwo6vaxchnjjXbpoLgsJYP6cae0Sqxr8PxLR37kkAKloOJhaoxk9Xte+
2E/GAhQmEime5vWT8iQKxFqbMDTJ9IQHZYySR6U3A/KOIi5WuRnjRDTQ73NvSlfb
Bd+cNT0njLL+PM05z0/qEF7TMeTRb9r38gMEWrSLhLcWx0Cq2N/x+rUni1g8wobu
Jp4PjZQKG+3dSosSy24eQJDhdDM7AfGMjE/hugROQZETwj+/ZpT9vh6vjsUgIw7T
LbnoBrmdrGdeeNyhkaLFjP9pnj60BxsA9LYjV+8wIva0T9fhlG2vPlE+FPeOTtmS
YixEMj4EhzdfaHcru5XLk+D1ZHzlDv89PNFuwTwsb0ZP+//dun3IiZmU0uWRc3sP
WxApjYWbbePOaGNaEqR8zr8KM7R5MAQzmaoDp+lUhefBDO0cs+1CQTJ4SoCVQ+/A
JpE8RNSwAXFgDEKrfOVALA8I7Y5ZxqhfObd5uwycxsgntozuOvOL+naF+C6bQwQJ
iM+vp+YhMpl4d3rO7QoN0Zr3VKKENAp0AlmLLOuim8PQGA0Drit2FY2WAu3xn/lW
yx3YSK9aaYCTgDFGeL3LCBbdIXEmYV+92dusNjiTTo2ziSlTFx9Pg/D18SPHlEBX
ipLNpApIKgK0C+zlnJq+XqM1z55HH/cKzx11BESbsQeGfTHVK14fjUx4PgW8oqax
OpwQR6r9SiV76lbi+rCLSWnP0r9PXi6TDWJ83ZDTAFulEw0CqGNwfQdxLlceYufC
f3pvihc8lg4M4I14Fwk9FN4ocwQVrDaDF6p2sypyNX/AyuloW1kreY8u1xcXxFNd
QqVQYTn3J/iaZr30JU/s0aSXSMwgHMrKiVVvgR7FKhiWNAu62A7/TJruiKyHc7AG
2QDa46zTK4rwaY85MVv7Ew0beM0d+G0HUfDAGFZz8lYHRa1fUb1ny7AGn/8IvdtO
LQ46UWbdQwJJKH+qUN60oGk3WHdQ7yFhjtC6ntEJFbh+/7nBvP3JcxfVWo3k8+bl
Ottguuw2EQaKbTPAILvl6TRkhNbu2esW4yfihJhNbCevZD7FfqFrNZryhYtS15T0
L5ZDe1TdtpSh45Y0Mh0iypdJ70eWsD6aOhlu2+/nNegmBnFm3wWGwuC26+NAyrWR
VMWwJvAlbmI705kKeI69EuewlwP9Q0bRWiYyoR9AXAFw3vA8yb4y/Av8VI4iQpHo
rjTwMyhmpcutr7yJf3vaL4g2ZjRkxZST2vNag5cyWRlComC8gjq0dCkri54bEplq
bzhGODKBHCiqgNldPJeek42X/WQ+bhjyFyPP2Qj+LZgIUuubMpdHxJik03x2mxqY
Ntgz460NSKAkYZaagieOPKdyw2LgsbFgbUPhPP5ZU2nLqNKU0PBrt4kqXs8X1hVB
Qh3EEWMkd5Hw3hCClLHLB3JvjL1CPiXtVmS3S5wOpntbibZk5tViu2U9/OhF+0HK
RuwXwMu+B4IXvd3zykzRlnsQgmUhcRD9p+Aqtn8j6lyLMcc5mEDXuGcZVqErF5q2
j5yxOk3KpWg8cdNHSvRGCdqKpziSvg5ivzaHsDEZCmt0FP5WAYXNfQ2/UJGgnk7M
fMk+lXQHQ9MWd7MXDjfCwiT02d5wLCyeG+5EqO99pyiqwMnHmLHYwKkFvp+1Kwgj
0P970IrOqv9HC6gROBkrcuPz8xSi5AarUzY08MkGH7Xky6ml8BWAxrGZ/FQkGN6v
n0V/KLT+8EB3amaTu0LbCHgXxklE8Zy+rQtXkGldNpQotWIQ5JfB1F91S1A7XZoP
nh1UzhVwZUdJ/Kfk0fhhNPi/+7w0BanKebCW3s8HkeTRrdFaXh0rG6MeU9GpLt2L
qYhlG31NAR7q9MMf91GPVzAP0y3lcM0qWEMW67QouD2b5Bet37eoTp9sEd+isJR8
VIIHWKjw6tdaGMyT6U418aChV4NYJZkfIG3d4wmw9AMzM61XRnP1Wfd97aJBrBfL
cWzYWNCHssSZo2I3qpHZ/miMLEocs3IcEdiKeIIGeNXbSqQ0LJQskOLe4EcltYY1
K2BBNsgEwUhxqAzYZNG8DZWjyrR6GUKV+9S2vLDhH/P6ILDDCPoQkH8XDayHSCxr
l/K2jBpB0tJiCzfsCrvtUsEhiECDuuWdd4RpudIMRrtuhKNGjx/pNZEhwSWNVj5A
jqm2+73IuDL+gFnR1c1+4X6oZn46UwzhhBzfHfTaEjbhM2vTbQIhZtf5njlYdQkc
3h0fVztIv2SXBp1h6tzA05TQoEzZQjjdY7WmnfeK+MJaPI83uKd9csANhco2D9dS
1A7GHbNBrQxNkEsulL98fnUFQye9rWMv2t+yanoFSiizITyeI/dpXDfdojDXI9jW
QQ1RZN4u9StBJ0dH3R1XsRN9lwfl6I5OphMfVxkWRhgj/umEjxv3/o5kmm6abFMF
zNhD8ZSR+sVIaXDlErVcd/jtODbZtVhPSzDYvs5KE/nf89UnujKHSXeAPvcSw43o
tfKZR8Cvt4Q2V7CTS9vXRHdlt/u6ZMZcEKcq3nksbC69weLXE8HfnZQPCosEX2Jq
powXuxub7N4dqWfMz330Z9JPmZZ+tINTjObUCnNhczOnec2mJW9BLFTPQQ+ctr63
aTVR2i8tOJ9wTilCJHWipAKvYL+JysR5466sUdtJ401WpwpnJ9pncQniwQgvJ8/q
A3ItJGE1wft+Bu7poGn8nY3/0+1RHAPLChIsc0OkPRSMcMUV7a/zjy0A65ZPVJKE
b1Silu93BvdbipIs+WHqgTTWwB3G1qvcb0Rena4heqvvRuP4MVr8wnVxhM0ArwO+
R9hTcwHcHnvtlSBsWmAVjZJpH/23g4fbq9n+K4J6SnXlNvSkJQ08I1fe5zCCwS+F
xKvM2C1aFzSbogKqBWrS5YDFomNnU1eE3o/ySAYxkktHBRLQ163HAoH4dNhMHJGK
tWjssUMNkujFnLXZiEWuo4DZ6Ci7WFR5n3epoHGem6uo/GUvxcOJR89r0TqnS9dP
hARzSnh2RBtzz236eE5IZUHjXkh3IVOH5bsef2UaojO1LDT1ZuHnFVBcjIXr6o30
9TpzYyNvFBeGfDxJnoNdXIALwlPKQMtOcqF1TU3MZl7zv94+7UmCh++5POZn2R3E
n0OObMDGJy94HuO50DbL45+b2/QC/YKIT4D9vMZWQbE2T+i83PCoWJiizIAV5vPM
39D5nJjtAonn31OMUTWWIDfPGHcI9ON45DBvmoZJp/Q794iqLuy5ncSxPcbMhkH6
a4xuapBWK+SILwKB0c7+/KDu+41KOIkoUzVUBoBxnrTC2b87ZlAbclO4wg/IEI28
4NSLUxOYyJSA1slZ4YGwozeS17MnYrg9vGCOuriHbmAz7EbUcbi+e51MT9sR0IDU
1TIwsjpCIWaVQ0xHitiUAu+9NgfpTlIxrEhfnfHkQu474tDDneZ8XX4L8UB8EM9n
LCZcEgbgsFjW5I/4cyvCo81arKcdlqI6EvqUUE4em1NyL/bg2pdCqblB5ggKGH6q
Qxcuw1NEMvscu/fU61hU+AwltLvGU9NpDasjORfCD1law/qNtx2nmSErQhmvvaw2
flHauGtXWkzyE5Sa5kQiGJwGfsP070nVCFkLrFhyj6XP5BtkxbNgE8Ztxpnx/4Bf
zHsL1iVco5WTnol92+gTOJXU4kOhNogiq43VDffx7DwMZgkXuXQdUw50b/dOVDol
vOx0L9jp4dBltJwqhRIl6jQ9PWLbJAxzwN4Qx08N6hVhX/VRpmLr3daremAwom0x
iJMQtxJsK7pT2x2fXbmvpIPxmkb8NOcUUen/5PRVeC+Q0TdPQmwcqgqHbUvmAkhC
CuDtez/4XBv5Xax6HHAVcp/Z/AbUyYSPoNJPayjxJuMYf5nd169NRHWkmCDzXy8B
kFzKrmHuYlTcJf8DtEs3C+osWbMdHJf0Bf4SfHJOo+RauHAXthYTxLU1/eLOd6Yp
69EedT29ZKM6p1pu+oZgp32l9kC29srALz4d5SLiUwS8/b+Z0Cirk0+ywo6AXWaL
adqpGhg31BRJInfY0vjZ9pnsNoKiGOGcWpNI1pooRZpPNn+dAOPNTzPueBcdxu27
bEVZ/PZy9d+mogeeV+cjYb93HB9Mvl5FGKcv0txN9ynFwtFyM/lLsP3PJC/g6e94
GO/AM+Np3uDQ9pSjv9zoFTUYZw2CLn48x6KUFfeBFItKosJE8zsb2W7VF7LU9vNf
NIp0FqiJ69It85TGgo7JDrS3DkewOMMYxVWMT8t+rAHHn+PxWA7lAG4WZWFYMI9P
IKM/V2m+xjpb8Bh2UVyxyIyb1xcS7PEEes3b+F8ghj3X6kYlr4nIAbHmoTxOczVi
hmR4QArAw0WptQtaocNIU6iDYC5tkIZXJXs8cRajHIEfoNTLM5iA3ock/2BdSbNr
ODih8lpV0TMs8Es403PLP0oTIvYg1ijxZMKsl2N4CRhkJuSWMTnWySCoYgFHwlKO
9AjkshezHC5pcOSlxRCWLFqNw6j4DQ75GiqQD42Rg2840PykI4nRWp2dkz7hv5RE
2/z1DUC9ccbsKwEJv7dCnLc7jNYzmbNowxcc4KZap/v2RLV2N/o37PjronXyQVXs
1MWYNKTJzFx1km/Th1t8PQ/ga9ehNKL3x4wYQbe7HjTq9p/uYRU1vuS3bl22PaR+
9lY4TLY7Ro017WhhlmvDVESNqce7nLjpN7GSPAnZD7vkHATGJwCgal/xZH5chhVl
jMgnWGFZ9s3cCIivS8zMczL4aHP7qHP/JNFikH9VQ/tHTZ8VNOxOyR9ibYycnuZW
1T9wCc0gyw3SGfbExAs+JFJrwLpFQOVVxYMAPQNptDcF/7asGwfFVSaP6jZ9sNFU
B5hnPbVLGIdM4P6oLMLY5oGknD7Rg5ra1Q4IIdQAFgaEP0AbJ0nqN1CUE3a8NfwM
uG1REMhwTw6rKZmE9h109Btz/6JFQwb3MbQ/RGOd3GThiMEryQI8F2hlITgZboP1
lNs42eUn/U4FjKBIgLbCjXu2lj3e1cdagUE70ggrz/w2vc2KX4EPmSFA2Nz3S97A
RPg84JDd8FmXE7RGq6KJeY9KyHdGgKnKugbGVSDOqYCo5B8oR/BRjT0XwrJeVAIt
qekFAN9PxrGfq/1Nw7SArCRLao5bLL+qghW5MTMKbEDrgebwWxTgCTh+E6nJ9BjD
dGCd3EppbZe+yc/VWsyBKqjX/TI9MCUZY09N4lc0JZ4+qTKqpEJu3rk6szjkgp5Y
gZG/rIo0/4F65xoAvrEo1pzjFcrUjUEV46aedXElHhGXlKWPQ23B4/HoBgDf1WXj
mY79ybYxly8eP5VmD2arRXyPT9Sx+Lv1y/d8ORQtNpvfkQgFjW7n5nk98Z0dUlqm
rGFVgiQxkdnraLM90pQYQuOHefvApjb3BP+asLv+QVc/DWjapWVAb5vtFuBC1Osw
9TOHkDArr2uV/aLTFSCNN10o5hjGlwxp4+wqWWmcUknuWIbRZ6APQtYYrbAwadPV
kZ8Bxjxk4TGRXgqvpkWANag3OOqi5HQkVNh8LW6otapnG7Uq8/8axq+1uKpwIRlC
/6IfccDI+VDibyY7NqNezTqWXWzfN9TyDkIUnQUOqD3tWA/Y8uNtthTXpHS+zEuC
vChZtwLoInQllpbRYlgJcOQGgUhc6vBeaSoKABg5S35URldLfFha1ZpIKNeP0SAe
H9IQAkmwa+WB4kYg0qIVwFdEjDamXk/pDePk+6e3SizT/AfWbQExs6YCDdqZ+PB0
YZUIvep5oP/Wccq/Foyl0iBpEPprveU4by/e3BuZXENieVvwMGKLET3Y7MCBT+bC
AcsHPMPoH/cw9dKJrDwhfRcwCSF7LmH0r6Q/OCvP3DSGTNnFjYWTSifMqrtlONe5
ZuvQrXUBxiveEhB2ogaBEY3HJ0kabOjrF5i7pZ/gJFKR4XwZYzOzpJSbU4gOF7i6
8huL4vN39nnbyFiJfx28hur0f7ROKOrFo64ervL8YQAYU6TrUfNF3s+KErKtRG0j
LTVywLCUq2pncj7mt2+PWfSquEvp8H+wKugSewwEslzeuvCd5WWgG15GVVvHJF47
qUpXRMCjZSm1s2NiDaoN8fU3S60KTs2+womcRskLsegNlrzlR+jU9rAZ/loA9qt5
aiP4J8EMfNxsmjUuBd7B1VFqm7lorE8/z2gMStQFXR1dYMBra8BrcP5Ra32oCIs0
OLjI4/Ti1uDpZWNesMgYzUAn/Z81CCMibwdzV6uma9eQZkdZk7nCyCb4SXTPdJjx
hh+d4z1mZc/CyrgkVLnx1XOgs0PKAfhOlVnb2/cWs3eKcRHxopc6xLefhg+/+wT3
N/k6wGxiyiemD0ZWas/fPVRtBMU+mxLvianqxk1FPo24hgDk02GGdrU6tgZdG8r6
OlXmNxqpg+TAsJDy2NXhdPJRjCtrcXApCsd3gqeTDKTkJ5Q9zwrY94uY79GQP3iF
q5wbpC4RzmRcnNoH2KpQ5LBiygLwUx6zB35o0S5XryiqkQhVZk7cE0ty3LiAu+pp
LZmeB2JFGNbG0Zkz+P0IK78zHs3D4+ltmoJqtQClrHS+YTArFvMPCcPvQL7Xo8Wz
WU6g5c0/6LoRrsrnItEp/0lJrOfXI9tlsuGPRWBWaoqFw2SlO2cErWEYZekOtT+P
S+A+7ZEXtXfIJ6Uej5Dz929Z5AulTVQQWzWq9NRhaYJc9F4KYZtywjdkvDTCyCzP
/yIoOimI/4yefye/ESoc3ZsefwplBJ0AoORZechuKvMlQsZ2aOdHh3Z93skFMejk
De46j18L+VpVoXDmOiXY+Os8ZQZPaExwpnJMK2k90/Qm4EBOQb8XvJNsYr0I+kc+
UBHLBzqd+Xi3LzjRT0dzf+lysOMzGvAZyU3F/j3PRdU5EHjqSesTpjKiu5MLaY9E
V4rWcOxIKdrG9rpsvvCaYIaoKQzipGlbCLHpfjO0JryEqrUfjdc3TWtTI94K6tp+
SfvLrYSPUE8+nRIDCwszGqAJg04thCJ+AK8rbrRkCid2lZ1KCSZtcGibNeDMar5l
ENR524kZGXpwKlEwe5+zvVmxhorwj6xZ+BVhb80qJU0hfUrS5iVMeVQa66IEvjw3
ybMmZJC1YqNLuXs7/2wxqYgPGnNuQvnLCvIeaHvy352Xyjx/6qAldMFEBvIUK5br
V3VI7EDwoPDt1Bse2poOSeKimQAOBc3/P2Hv3MZrYGB268hG/rgph7rFX80VYUNb
+sH0EQMKukzpsH5Qn1DYncfh6sFh0T3wo3Hz+eaKrbTNJeSr1hT5IA/vwdz2cbnb
itkoyi1ZiUx0BPhCSqImFy5h0gJaHSvVQzjkPPDjgcruJcRiiy+x/T3W2aZAZtun
kjRjlgyuIUDbZ8RRQ4vkXKzy7ij+nwipMJ10/IWi/x+22AqKNIFsNULo38D4jyxu
6Chstp++A2rZRZw0zG5r2Vf7XYuEt1iOguBQmFLhobEp/HrNtrKsRv+gyuSEBYwt
vgm6bJNooQZ1CH0YI7gv6XLO6vJJWyXw/HnZXe/6ksIJTij3ItBLb/emlEY6GRD1
ayNgorZoHW58qDxU5fbjkI7kNbZMa6UzhzLHEwiqes12ijKCcAObZ7HdOjn7xkqc
E5icOpboNSbOObato2qnt22KivDZn7aT3HwwuTbOadHvHjaCUXVo+TRsqh6NGewy
OfyDuC5n7HE5A89/shXZabxpmLKxh9fMWwqCkWoVNqXlAb9xxPPGnfVz3UdPNUb0
CZS6hy43kGkUuPxlfHc/CU0oACsj81x2BSCG677lfIvmqSrdySnpVnuoQpDguo4w
N7YNfWTBW06gichDaM5m+R2U0yZcZPimIyfoerM+wcyc1f+NVTijWdijLhAFHw2A
wM3Yusdi27mYXBshv5m6e/DizBh9uiLiJ7Gz+83/zEDn4620V7hAyL5NdBSMGq5m
+zStJLF0S/bNn0LTTV7tWy8ELObbLAiI8FNoBpB5Ge3NO3efuPCm9qgSt/HMghkt
tL3VkqkiuHT5YDmOjG/cwsyUoOnqHd5lJMhG7ImX8BMDdHHwVjinA72/Z0mZRpWS
eWeSgqP2QFlntSM0gDv2uADkdRKHBc5ruUc4Hduj5NMDTuymfQm4LRxrjKks0Sbx
zO1v7TFwLaDwMaFwo5nPZaT0twxxxdyW2PsXpQdAF/Vt9IgalH+SmJBLiLES/LKY
H925WmYCy2hsOrQDUEXqYwcyH9cVzrVUkunHBGo63n0uyqXawcScXH7EUMfexmIK
gJzdvXo6jf+LJyRvI8gHM8ASo6n3nTWCTgBdBr0MqdnYvHoH9bPgx1Q2klzwsvA6
mIm6eJeWhH9wvn91Oxgkl7Kc7kKyxozWJab0069s83LMd2p5BPlDhDDWZupxJgTC
lerhs3pehZ3d+YNSHBoYZdfHMt7IlmGmS1zYCJgTqfJjg0Lbb6uLHUS8BeZqdkP9
eW+eGEOkvc407nG/kTWX8IFB/kiSCTPqj5gOjEov+c+iUedqNz2gzwRcaTmHrTi6
KAcKXDhLHJ5ZWcuGYYcgQV3Dxh0BaXZyrKhWvr3TerfssBI4RX+tsnIB24KLN/xf
SRcj+2ILlcR5VfinmHJc9LSAgVjfXby+6nJqT2kr3GLPEu8AHkE2GU4qbVJaoDbu
mGo0ZgsdrUDu7MKQB/QufHbCD6sWGwAU17p6pYqilYvnUT38+P/eLEIV1SdYykEj
ywwld9aa3oubfRyDBY56/Yws8YqHjfe4EK3glqnDv6v6flxzNOEvlb+X4xwCsdi1
8Ri4AMhAPmu2h7g7S0l/WwqlepXbmaPKGh9RCd9dkEZRYj0vDsOSRkqdw2Y2beTV
ofYKLnd9KbT64jdBLw9EzHfb/TvCVN7bwqMhlG5MFavjpAccL5bZTRU8hKWn9X4G
a+EZv35Kr0m17OkEdgYEVGXW4Lak5xL5x4xtDlHl6zcfKTHqp/AorNOlkSgCCe2z
TGGITrvngesYfFvTshOwnsF1FSv6lIcBfR6yU1JYtTRNJOe5rUXoMBG/OiMu3vgB
QSbh1p0pRLftWuvCqOquCQLAAEjBSzukXWY2OXlu9wutdA2GWytkLmM7258Td9JX
65I+izl6Q2Dj/0YWMquzRl5rbIBuQN41tbiBwAxtSZ33fYP7sS+X8ucy2X5oBiUh
Uep1yqRG31L67VEryPQbI9QjdIjixI5Khx5LunaRlAu3Ogz/GnOAPTHXwjgfToro
6are2Dq2DNQZz9kibHXXTEYjlOOjWA/W3oyHf2fVE30dLya3NUUgYF2qHlffVapj
QkvI1cNYKmeJnOqY24KPMgSzEBl+0sVZW+DEOt7fim3n4aNR8JI8i0CZQBYIYYms
1bDqA89ognc/22qgVcPLirpTU69pwTDkcJMwnovwN4rs975GslU7EFVY6tLnmAvJ
Wjbthlnlpjwlkiqaa6rbVP0ifZiERTFMtkRvYbL4qFjOc7M6T30SN1A2RtF/7a6b
BIWw2DccVqiJtgYkvBKfWzhrRetPX4I0fHpEOmx7oybvu9+QcDY7hA6lJ4gxsRY+
kyFezv034rQaWF0ALpn87Vjbzrri89WvDe7hzcEaesiJP6NwX5DGi3G3OeUxDTG8
U0G5AswwPUOmEXhjyr+hoySfMS6YZwRe2h1PmjFoVkGYwp9mervBmgw5gMUpm2JJ
76eMY5ASWWDAdmrvQ+ARl+JQprPfury3/7YvJsK/ahpidWv0t4AcrJT4p/vFdILr
2KNS2BHFv1vMDv11SHjQOeoQqQwjiNo3ggCONKYLTH67Z5TLaAosoc4X2LUSQYXu
7y/D+qwHdUylO3iaQ+MdxfXs/050+b/V5FJUqmmmco926EybH3FL4sPceLK2vBK1
EwF0CWHGKr2+PL3vjRyKI89BtiCPrqGPZCXeZ79IWC71SoAjeQXVetewiAkrmQOc
Leklg6sS11g4hIa42N20tkjojszaVwsuNkO964C4nVBjMNMwrsEdq68uTQy5sj4d
KyVKe3kzkO2j0bCr3O6gGpU78Va8icH3pXO5uq4+QfP7ZOxSv8HO2aufpFyYPKQw
2qKLFkAUL99nV7fvHbrnrc5/aeIvbsddWUHMxDhoYhVNMAqk7QIdQJ5qmlHnqvoI
TaG2nB8DfS8BaH6Z8Cn6ArrV+0FTNY0fbN2YBNunm4DzVxbRgXcfYv15bkQWnZkv
d7ys52hO0tKeWKTMJeAl/Gce5/XFLWKK0GBMQGi8sahCK3v2hU2+O9ynIg1OOzcc
vE19WahyhhjiL1917FIQEiYmmBR41PiULNwT0pMiNV7+yzSZIvyYgYkp0d9zKf7N
nGfRnkd3ieTyQoFyhaVE1CtP959+E9vBPjtSF9zuVytL8drabepSavw6Rhm4gOBU
UU4FHNoa1Hm1AMOIXLW/1L3CsrJlmSp3VsJkyd6QE2nwWq3uyg+D3VFYJwSIvt2m
J0/F2FPoZ8KL25w6REPtFLJIkAlDQKdYDIce+3K4bA6vo2t3E1E352iCOXN3T1Sy
XeZGiP/lRbbnmD5awEWG4CvM1x3pv2JtCmAMdTOs31Yhmxvi2eXO11R76+D6Vmf+
yQxh73RRpGfz0sF/7e4SPig/udcMJBW0vzJW1ofAajC9qEeyXIzdSV2+NM7JwfYW
2dEvrUCaySb1/uAKWGpkKP3+etd6IwDSXyqidveVHdgTnKLnY5iyWNpoLPAjVcR3
gv5rQY7GyxkkwIhsNHqu2xhlTc8cZ+ZHc4ngnkdnv7Tg5/K1qilC9tWrE/r7PkVk
tZgIOSofxkpkFSoranXgKRbBLHO4rVlfLZUQiQ+X84Udubm9D5V2ae0itV93P9KK
JOD4Fbggo/1vlKJG4PmcYR+UeswUx8mDv6d8IbBGd2snLir2CXw10y1J4Hy+wBgA
ofO/oNLJHEj5EsrXWmmni8xHadMpUnqGMz+8yv+Q/wnm6sP8xq7J7DaHbK6cuo0I
5fZEvRnWvJJIlf4C/BgIYlIvgEIWuERqqka5JopE7dC+51XCODf0oqojhUtgxMrC
WoEqIDKHydlTruw/hGwgFZqV46pLTdSFsLMEr/Ht7/xB2LgDByqm+/B26UbZIkgM
a/lBPfpvValatcrxwuE4Bu5Z9k4eWM7dEB4O8CxgjWiyQ6HSZPzjnLD2AGm9BsPm
tQ8xvBuNxBP1QmyCUlt6h07kWw5HbfNpYU2pSXWJxlkOpn3td0MMarm9pbXV3I4h
gCfDSCWJ5nwIASNKDob5dwFg3/ASq8Ano1smCtgnkuDJ7rQdn+j6a9kO1FVbncgy
sMEu6GM6Lyeu7I6v9dujTC+2Wxy2ZPj6ZCg9qlDYTpgHA6Mgw3b3j50U7QIfPQ+4
koc9SQHbSSI1xGib9Hkj1ZmFQS9c52HXYT01B8gtSMFnuJS7wMGQc84iNpFjbJfl
twDFm0KABsQfD1Y9od6YEXt30bV8s/JNvrL5WdMj1vWN49JmuRYLeHymKrdNhOet
EEc9LPTV/ir1cXzB8klXKeprDPukYQI+9IIVRJwC8HGm947F92iIOZpTAOHhbg0W
0pUccQlHxaGK1Qg0KyhujLjxFgvbmp3yPNAzr+4QUzeReGWDxXhOYTr0WVphMV3j
QSOz/qfAIM4D3Rr55AFdGTRD+bdp7/FrFbCMF2AOP1/25oL63JncfYmKIL2IFjsV
xbej86fzAZ8zOvuUzrg9Qc39lWwNbsArK5h8VfF6LnIPki5J7bm1JOKjQfIxSMyR
l9kicWsMSjHMWCEG+6WlyXsKKmSgkUzQoAiEz7WEbzU7TpDZIASE2DRbkEYxpEHi
2xegDcPH2W3U66Fvw+7C4byKhmNL8K/4oKcH9C2TwZM3mtiqCUNQU2lrqpcljWlj
Pw5oTv+pdca5mHZhyztF6nVCNorkPMy5bLWNpQwWSt7MLjiFfJCvXbv9y/Gm/wKH
AaVStIhtS9NvQ6X3fI11BTMDtgl1r/a69QPT+6j3TydCq3yCHablY2FkwGnEbvrH
3Je0iiuINJjJsSAim7QpHpetA4gkn2SAipKMCLMIld5h+af3PgnFNOHEdYasOoAi
jNrr8Y747gi5UX9mTdOeAK7FsRC6sXM5PjNEMraNiqx5Bh/S2YQReI4CVvk2+FB+
gt70z76wf4Lk+4NyOg/PkHGhMHlGp6Ix0Gtx2tnfM1Q3J+sgXWfrWH/zwZOEu7wB
BifUbCrN81pFHlfsV5js9n+T23prfPrUl+6oRVhgaWZeqzsjC3QXIIvEQjBhPlIQ
8+rDNasdULD1OxLJ15CXF99FKJvgVgAODkdy2oL3S7eRCKe4wwqVqm0kKXjPcHJO
yBuGopI7TXnddkHgG0DwYVcKNs2qUg1ueR8ZVB6jI4zPBoJcdFc61hHPIN2gWCig
YtAweGfyaFm/6jb78eVpp/ska2vjtW0Rs4N1r5D1vHEYmKivm/x9aQsezfgNz5xS
fvj8EBO0zgh8QfTA4213fFeuyF6DLSnUZ+e6MQ7uSxKRCLq0HFzn17dvq+2wrXHh
FCjT6LIazb3T1FkwvWU0CeBXLdnjtQBhkMjAz9xQG4YB6vo+LU5eLN7pe82B8PcO
haTOPjsdEY4UYLIKdrV9at8uC9cjaWBz6My1EM82HYvC/Exwg8/QAad8l1gDzdDI
BiVBbrfWHsppgW/ccP/BVLcsuhMb+qZzIdsGn71RromcYwadqZ9HD90CY/fkksUA
TrlOJ1Tje4PCik8yOh2XxvNqXR3y9YP+Mjw96Rz+WWYZND/Fc19RC9W98uBWnliX
cZtlR7sh3EeInz0UfxTWPK2Z129nQClyh0QZWZYJ7vz/cZH85URLhnw6AyJYk6xf
EPVEvkIQ7XzK08KT0S2w5UhOWGBrf1ExMPG6zaPiv8Hpc16xt2TmrlqVzRpoifya
Qe5LPINq2FGD18kU6+3TPy/HOXCA6PaIxF4Q7/2E39lYjylW8gJYYse84DlfCRig
Wn7FK3FzlSmREhtej95jgoIN3CRafaBXr7Aj5yhk3ydBcWMNPFi0nTkD3uJ3FFVR
CBO2LWWrHgEfJKXbp/ZLD7uw4JnzmJh0N1pUL8ke5nJKoXBMvBDuBa30ShsWyrF5
TMXd6jd/6wTt3FqpMpma0tjnUrAioD8HUG4PU3/5y12VndRKlP6/wFhfHgwSmiK7
KsCvF3pmTgNU2ow+Jzxle1M7gtUkN9sZN94XpghjrBJ8qq9ie6t7MGbMfszCyQa7
dTfR8zV7RJbzdsQLB7rFs7reRR8PzbHaOT1S46JEJ5O3nzC+WHKk+eA3mjyvp8IQ
sK9Nrx4Ek+tJN3NYJ3U06hHrnRnzldLWKxAOeXlV8yidy02ZpogGd7gADtJx42DQ
vlzMgpHeCkIo0peSZzRAlgKsSIhtYuPrAXhDBuxwbW1xZY1zS8XiAqS0UvYmaFA4
S4xgfnPeysJa3V+H3XJBMV2MBWwt/9uo17uVWO+NuTIGPWvfigvdb7BRCzf2PaDt
d4Z/o/DhidYa+Yh8zBg8OGF68sDVk/ORaRjWIdnPffJvdlBCDsQfaMst2G13JTLy
Nb0EVek2vQnR5yFsKTzAbXhdPS3VGfnM3kVRnmY6ue2grHPty392mygJPqoI7WBV
sA3Ma+LYJ3IDvMjIN3MWxXcQG/p7sjaFfjtPfF+3MtOsztjOXezN9rc8/mh9Rnj9
0qtR1sgYoYqmpWP7DsrTrBbJ7mLRZZW/bFR4K8rTDGaxm3h4CD6pUcSj+JX505dd
ClvUQJbh5NizteBwfnY4q4Gwq/dVn7AO+lQuIO16DqISD1OfRPOIvlOeSN+JBaii
wL3sGC/B5hCyihnKMBkD0PKjgpzafI1l1kZBI3b38y2dw1PHbFuQX91RZ9gwKb35
k3QmOpn8Czb+th07JnWtBPA2JMdJs3VlszdXNm8BFn64ODsxmTnZfWq6/yTWKmtm
jWUDgbfNKKh6b3Yh+4fxz/BBEEOWbzcjOfSjBZy1obXP93k2GlgAD+S7KEj5EeSa
E753zrI1MVbtnInN7l4IE3EMeWtWjWg+lW+YyJs50nQH1BBT9AQTTdPswxYbyBDl
oySuyPPsSDkBxyx1+OJT2XwFhhqo20WTp+s9Hi/Sdmhs9sjQlS+rUVH/CQ9IojuI
2MmscEhjW80WrnMIKZ1ThI6IaqFse6UCJEnB9TqH3JqIVChrc9BAEfKXQAOcP0sd
Cwu60NWjxxqNAC9Np8vpk8k3zIHZsKUDmEdIhBe9Mh5W0T3wzPtbEaSc1+2bZak2
pdBEA7ZE3n0UTRB//blXBjkyBpDgT4omnI9iBW/v6qInndRE3NCiBH/QGlu+Yq0E
5mk7Ibq8bpVJno4Qotc99wRKDq2zIIKfUKSt4WvAN2l5hO8D78GiXC7JsgRpbswx
N6+q0VFIhIRbKfUd4nk6SGjYmRFSPXVz2a7Lm1jGaj78U6dN7RFpz37nJezN0pPF
GWVAoeEaWPSVbAIEDkylWp8xZbFIg74ESKhWNdepCh+ZC9nEU64/eLsyndz6GbJ/
9Tb+LDeAL+p55fORVUpckhPXTptcTC8CPE7tAmyFP4i+V7Gh1NSuL8FOuEpkf+Qn
zuKeSyBxd0ZrZuPtWdTbHrNctgDlBSevlPZiEVpLXOOBSCFsnmLokusxdXAyTDf5
wNMxbtu02lqS7SJDojkuJN30GNewNyTkzT89m54Ushd1Dx1nOn+ybr6+3qo5i/at
Pj6wzR36v68YL6Ukfg1b/iatkFA2SI9nziOlPImyAwvNuAGC6GdoRHJN3n12u5in
axupLGBPD+Yg/VUph1853iXsmMmvqlvoy8+O6rOa6WNmyaiDfhTywUkvr+xZa/oa
aV5TI2t8Ai/eToBZXaPVsLSOxQEI7HgaJdAqKfevD9UBO9aN937fx/+UQCYTOjEQ
vFTBNrW6sOu7MN/cHxI8lvhKh1pdE/Ci29TbjOc9EQTfbpYsBXPNtAo1O0h7IGR+
hvsReFkcwMsVPRp6IpHIiJJUi6yU7S+/PPM9ojoxS4+OSw98SNFsXGriUJzHAkZ0
BqsOXY9LkgbnnFgC38qRnx3IMJuIGmFuLuJjHDteIoCOLHPkmkTyTXjiDTodPwiN
G7a8RrFn9Cqddunx9cI5FhAKhva2fRFIPSHVeOEDKCJGFQsOlZu3FU5eC3JxWDRC
1vosysNo3kw6lXxWo/fwbFR30cfk4mmEKzXmcg9mItwLvJeJjiWJY7rjA6UKC6AZ
LpuW065MHikBAecvEwmvm/fqwLURDMbDXEFYPue1nyPYSWBLiRboEekrvRQIYDvO
8KfKpny0SPNoiFAyolVKNT1P9sN5q18Ay25nQor8TKkNHG7g374s1TikK1AyNoWb
OKzzn28nq7RL7KL/acedgALRcPQTJhrapNkBTY52TcVCVoXluktwGa/W+hEB/boH
q3giuB101xlqQ3C7VpOn58usFAHBWZ+06ay683dUCTcAiVmhSsNnjT2R7CzNDgjG
IBX89q1ifHkL9dbfU2ULrEQOPFBc4G2PJtIA+phj+7HyNFjnGPEtBtk8ELcK0f6r
eiV6waT7bzjcOh7xvG/qHIPfWogPgSB/jZrrjfKti878HKLXxuOdnX0ECe/5SiuK
0sZ2tw4DN91XxR8tO994vCpNr4in+J9HJG4N7+WKJvDg3tEv0fj5/IUNvu/pH3t+
y9NTAmsmITwnJjJH0b0/7DZnUki5X5PX3L+nKSdV2fOPb6f80cMfmO47sJ7bdn1w
AeoOVfYfVS4kcWuvvJWd6LWBvD9clc0wCaBu5jD5LdOqUUhpsiukzO10Z/q0NGb4
lPI3aaXh/PUCtnFG0ScCk9Tx8gD7pEPZ2/JmNZ7KgCgkpqs2QSVxVRHm4WmGPVCK
56USoL316D/9dAaQ99KywkTYxOvILnVXWMjwT4vmJSvbn1fu4nkB9dTM0DEl7hXE
1fDjxn+diluSmUg2u9eSxDRQph2CL6NJd+eeNsJau2CLVZkAT5gBiNH3bBe7FR9e
/3hijFqkUigp5aaEhMwnOX63tniP0dXnQc/aROfjOWKtyz1dubUOeiNngIqifgv/
Anifkm1nCIxgQhda8NCIW8OGqnHFv6HfJL5sJ5Cjqfk915KN3wd70pX1pAK3Ld8t
jJsfvj/CtQJBPCZ8fhgo1RyD9gxJ0t6KGzOAKN5nawWgYgInZCssJHRoctlsVaV1
XZi+RgPHVzrJtfhNV7n8ptUwDn4AXugorVyTxn6oVJr+zAHMb6yQg/6neuc29KDG
1pGzH/3BE0NAt1pKXtbGIVIAbZ28JUcLsvpYxwqfB117bOhouFSfixMGcwZEbrKM
dEaHgKAkEwOM3uFYLaBuR8EfumzUcngk15LwiNfQCXPQp2k9Dk6wjuv+GKx5lQrX
eIZSRWH7bpwPFsydha3P6dRqZeJeKeiGCzSgSYELemYeNWlwbIGLtPONcWfVmjXv
YtR4fPCZBAS+3HDmNtHE52wQFz723Q2DisynlkSn8MaZ2UwfclkuXNt8qQJxSzoB
kMDV72uppf4zyOLbavHYIQG9a13kR488ge+MA2vx/wmci+FqdZq2/O0ec3Yc3zeF
o3eh/MtWTSe/yj1YD6GFBMuDuDzh17ual9yW9PVeNGTSQ5VDd7ykxhqeUr8VTe5w
9JDkybtY1WAyQlZtUWuRn8BUo9KrQARfrK8Hl0v2GmbAx4yWUBuoQDjygzvZ4jaR
imFWiNYJ9XL94COttb6jX69S8QWVMvOF7GV1v7OYSX6eGvJ4vCUZDLXzuwP07i7q
EldcRzkACSeeGbpzFZxLzOFb7IMaGc05M+S5WaGbrXB9rHX9dB+dMUMpu7UPg1Kp
CgchndPQ6UaBlrcVweUTkEQIq0LwjGStEaqwZHwD2/XszgVJ4CV+2QO0AoarX45F
4gJS4cPILCD/7VUE6UCTAbkASBe4pWGkNQ95mexUctjJBkNMz+IshKSoXpKaVT1V
gsLAspbrUjvd058xNOu4Y52jLgAdz9Q404vlZPIjoMA02Kb3H3QcvxuVd4Wwu9SG
68hZy9Zxm4ztTUxbCv2rBf28GCzMS4jdtXlU0ypSupcBxLuTmhoY92gNkve+ee64
Db2HLmuywpOMKRuEqfONm05Rc4qd39SD2LjzzDuZ2sQ0FttTCYBSg6kLgGfjTCTB
JWqZz+T8PYn8KjvAvkekX5TA1IP9hjZibDk/WeDa7qt8GXZoDXKCwUmvp/yf22ch
392IdDBDdoOv7vPIRSHPKBMeYT4bKmSwmh9b++1qTBmkmtGlVeGMUE/iG0kxd9uC
ZisvtHyqo49iPf+6/iouZhv7wnweDai0iH+TndycFAEuzSUBOegBf2vkfx4cfHdt
kmoDmiRC2zQCKI0q1yboI113pQoIR85262aKLvAglQvIHDGA0Sygm4oxyIobLf3X
l9GC9RvWVVM5gfJh4k1tzHfPSYpE5yEGL7omfLTLM8xB6zSnvKOFUQjd3LMJrcBX
tEYpw0pdpgj0U5fP2yPLWQwsJ3GQPzTvGzbNESlTSPjsXQBpUpnxDonNL/+zsAaB
Su+1kERKM5yO8TUtjf3utMVhH/Ccvv1Kx9HGBsXapw6rnaqGuNIC/z+oSmwrnoX7
KxnpTfedeRSwCKrZpLVgnIlkLBAKhZK+FUP78P7E3QZGoZSV56Aoi4BHwtgiH27F
e0Bu/WVkP3ST2E+VhaYrmlPrtaekmwLlsTzIcAdwBPIlg+Cy5Qu14ZVoKqGA7FQB
lqLNC+su0U+Vu6NHPFrbpulmPFdpK+gbz8YNUYOiHRet+I+41uG+/FENbAb9Slju
sNsAVqTi+njvJe49vouvHK36VsfcYVnhvBAdP0OuUaEhQTvY+y5zKSssRQoO8dly
Xv9C64qSv9x0BQCfXnHcWzyibkw1gLtmTBZxmBXaE8MxGzDpstxLfSetq2vpxwyN
aRbjVbXj9IsmIRswn5GxlkXO4mgEGMl8p4y1cPgFcNY46NH/oG+nPbHBLQGmAUV5
0FxbF+nFkr664Vf96IgcnJHE4sGoBpc1Z9shN0UJYtEE84yJvI4QjmTPcj+6uE8j
/UI/GhL7CqhfpkRAQjmHLrmXTjjRC5tKf6lPuzsEPYijEfXhldXShSzdKhS4j95O
N7ccyVpXqdG4VuWCD8cTaXfgLwp8NRUHrclzD2RaX0y4Ubfg8QnC4oN3J/MH+VKw
ClWlg+jEmP3DVPbYOUsx5xxrzaADs1+SYP5C4b+bc3j0DKazvOByxjJibqkRtvog
rlD6vmpCh+q6o/dDFoCYibR8etDXNZqrqhY3X8JL/MYeKomd6yUAeTpvSr3i1Tiu
K8br6QmlAllaI6vz5CJmAqIcv8M8fFDnjUrK5nTZHq4kIe9c97gQxihQZogeDaPh
vXSI2Nbv2KBuo07enpp/I1QkyJgRRQjOV4QMjk4wK1NX4O3unrtch1gN42zq0eDJ
yiZLmI41MvuZJZoN4YwOipzjeZRqFYlujWe3QKxQBQRPSCQ7XOh+kF/XmnTI9Sty
dNfYGtV7Jtbw1fxAlqwKPJoDgOuJ+jqbKTI086BTZvbOLDVCaSxUYVs14cj8mEQ8
z919w1onQme4ZQxBa7fd8kIK1SGffAlGka02p+g6NN9ZD/GYZfjvxU02D6nqxyTQ
Kq7XBNOA4eBNuClFbP4oIOyq/oFWUwlUPYZvEpmYc+ziM00Aqo3ZnCcZH1y39a9C
Ng46slk0GrksnCikec2VmFe5kJo7ua9VxMm/0TtzrlXw+1nJxJlj4TgAD0pGfGYA
2KT7lqIwS40efvxIajZcWd/RLaS4A+38CUmCdhHru3yOTV3HmgtkptDZ6i95A81f
foDWA5S4nlDovtaYPwkXej2mVFHoPkY2uKO4jfoYFNG1HqGMz/CrqqTCxu8oiLvW
USTZFs9K3Jz3iTxBsuHXF32JmngQjL+CxxPWgP7Gp8f88odURieTfVMcpTDoX0JX
PK2K8U0q4aLJXwxwdP/no3Zj/lTUwtO8k/ArPcnMCnAgZyernMSFCIT4WJm1DY/w
ZdOw5vWeIOf/yiogy2EWXiPxPW+OueufYLSoFvSR/TToR8n8/5rUnsQxmAAs8hLQ
N9B1yGfrxo//uHqw+zuKVTELKfojhDqiDkzBS5PbY+2+BG9M0TRL4dLOwq1FbOVe
qFicIjwhdZPnXABgMjb4skuhEuJTlu4STu8Fv5vjB7MnKElhVaHYH2JE9uZ5QIzr
L1eZhYQyxdaZlRgmxlThK/wsBPw1cCsv955LXQvkFDgb8Vf8Eku8icWwOz2T1j56
zIgESYLKK8MeTtvbRIKfcvt+5zcv1Fvbrd09vF+Pi/jL6p8inoGGKoBzZCiKCkWH
Vz1i2vHMPNjHrPLNdgVJKjEOMEuGlnBH4WDmcI45sCy4e1qB4nWh7FtTeAdXNg2g
K9laG27wn5uUC8zWHW2wcxA+7P42zX3gwpWgYGEJ3JLQTBwZpjKA7f8aaMgJluPz
Bck0CseUqQHiBCY791mVlfl+mnJ7CI4OGNREdOl5Fx84P03Vb3DxdSdq5xhNYVit
LsQyZbLSQfda61EJ5zk3DCWjLpXmINiCjSJ8lUdkGM8Dux4uX5O9urMlmP5PFT+K
HbEFdl5+3PLmRSsJmYoDIy3RBSILODg1A4PLIXbFCtU4k14NH1533txF2U6uutfQ
F4s+6+OupG5alwpFucx+XNVjrO5DY58Q/uWqCzqPpBQrNRV36F8jfsceBSLKxaaw
hQcNVWtgLGIdrJ8/Ri+HYo73QPD2cYrirdmm6G3NbhESKh52doRJQm42QF0cyadT
437dQHvhrb3dk0j+45ouWa7jr3MJaThE03LwczSfcWJdrH94HT9HRzTf1Mmg8/cz
8NcSAbZRj1aopGuCVPKz8X5G6Ro060XxlAOaFJ7OzMDHxFud9vrcBOpJuMjeftdO
q4VN3qp4luC8dnmaRoLr4oepXMKR6QybY7igA3NBFimocXFynNQn/Llz1EI+eSWx
RiqEjXHZwaheD/UYNdzTj/FiNil+wACqYyo8hBqlqaTns10pJTnBGHoQ8aOOvmDw
F6aRJfItdAJAk7j6S3CFAfar284rnuIHeZLisnPzJWdo2NM0V9csjwZarWRt4F0U
eQpcyR4FgYIWJa7If0q9lRtceFicDzc8RpJg4hH7e22QUL6GS9fBjrcX6HN0Ql0u
z3Yspe9SceEuXlJk5Xc30mP1xOjXDA1nzD2lpAVpdwr7gNJFEIFN1GTdk9TJ+Y5q
ni0WOEy1qSSA8lRCi3fk69M1sY9g6luwq/1XOyKghXS+Q9EhIt6iwbc2NxsByL3n
/XoZ0kixaKCwW+ol4EqjBc5dxtDLp8TN7IwMFrVeDXkgEP8Q02/VmNS2jpwrw8qn
cO5Kj/xhELKSJbLy9CK4CzqvRntQ34Hp9RDpYSKMHOsqqQCi+gLzAsbXuc2hzK5q
+TcTNUe7DGJHmD92De6YmnviqCdtyhNdsU2JLV/zaA1J250wsuapTS188+fgn68M
DDhdHPvYtRMThRVu+V8HargPBClj9yxpAV4fUeIedl/IP9sSF0ahcxso3+Ki4CJW
C8bU1KM+rX7yHYjmwsqyccDVE/LHAXA1IW8pcWmxDrMF7HVsfhS2+Gem9tXMCAun
Pi/NW/bUiWwjSpJPhut/+ATmYBCnsIiEq5zmty/i1Rp3V6B3G/jqpFRQU+1d2NR2
EXGpFSEvgkqdx39lcvowWPlD4+q5E0HvS40iu4opMlf6zUMwzY7YKl2CNYZ/Ai2J
dFj6+8yvBzODEpRJD1sL5LUHtXNGAA/fU4HmZG7+WtCce22WAfi5GNB+dnnPGG0B
UYQdmCOQmzkWx+F8li4sFAAkt1CXKQl0YHxP3pMqT21DHcQ/Sa2GjmYACPrjzpBB
ELN+B1cSr3oxug4fR+hyXi4Q+6VbsQEOa4mAlvyCNib7K59MmoMslHYwYaq+kdpY
dKBVS7IdP0tdQkfnlI8iSLaqkBm14HqmRZDXwI0orJ14t5lkEWZNjbidrSU5wlxW
XN881PydrnyGQLcXYI555aOX0JEoWfJ54/4QDYST8n6TymFFVKgZRCCoZccJkWls
CJWRtWARGSHie4+QffRkfEf/2luT8NV+7m7VxIlimhkAp7zo5QjnOWtF6o7UJQy+
fpMNvTMYHAI3YKer5mZUo8vL2fNk9gxoP/j9pdldxlMVsPYCAU8+YfOmmiP2/kyv
NXqBAjL//wSfzVDEn8Zd5mVPPFoxKZSPZXPhoM9V8gVw7T3GbhALzb0IEMxDus5Q
pJ/zZBMNC1OOzRc/CNnLzyzqKjGelyOPKpP6gnT1MO5k0Xj8mpnDYSvOvO6t4H6T
uSH+D/2UXlGtmzGFgfDOqalOXXItdmW8pPUO3X9zkj4LVAqmN7c6JhEs9Z7I1gMp
Yg3EjRRKEEdiOu4C2HswK9nO8S3GI/hcPXoQ87CW0hZhXn01PW/kTg+oW3XSnTG9
tXHYYJVVfwPDFqp7ELoYRrD2WPObnZ2hiMnJeLqoEpOiNs2cYZlD/G3XbohjTq9V
/9kG/DUVDtbJNV5X/IVbEy8lMg2jAcI4LX/H1xM+VYE+pVqCY6M+9P5WWPaJ2nlh
SAABt6mxI25XILv4YuQGyVRRa4ONajzyLQKocRF6xpQQZAZKThtkhpmymGWZVOyc
fkZ/i9n4F1U9BaSirbimIdVSmJQO/maQ3TzxpOnjqwC+X7vWXGBKgJITyFQUOBqB
qwdXCj5ZkDRuxQW446NxvndbpJSdBQpTjXW9gfcxs8ckk+gFEwZ/gCuGwTXWREsj
RDUS7pnvanlPDzgclRdxvsowsJQZ6/f6grtSMOBDyTZZBXYbTUlsZx/9VMVIfAMa
L1euYwQsFY7iVAdeWHLRJIfz29SgTYlAeXlXj3l7/z6+3yXO7e5diwU5ODqq3W1x
moE88LWAHMrPSJQOQJrOvIXhQPrhiYIExQndChdZl0i5l3ZFIVL/zRINQI2CCWL4
+mwg0AIWhZZNPkcY3bj3WEDX0iOXb8Asn30dMwuMZPJw8ZAe64UFJe/HRB7WTu9T
DdnWzdqTIWE4P7S1J1a+lBE1oKru5t4Zej6h/4nkVPxHlTMx7ifBGsUfzowsiSeJ
9O8E4yWPOaI7nx1PmwwGakczXr4YwANZINnjVDd/3Nz5pRZNN9m8/isSX0pyrL9T
RItK3OmnRy5oCfHGfMGGKq5QFWAyW74w+i/tS6BQedN9EIP094EqKihyl6QtTwDS
/EyozbVF5geiXv3lLbdobiMJ7PLV4X0OOoy/YCMxnBJAObHeQU8YKRdOua+F8tuR
SfITPyw9tfRpzPrSshtFMgpU3wzjirTVUTnwbdF40qFM9Sz9SZ250JOg0+xvkPcS
yj62sRJzHRg55dnfYr6GNOAAz9qZhV/n5N7hxDL8v0kVZdIIFlUjZYHRE3dfR+vV
84mE1ve7W3aCQDuALdomRBF/OZ8+UG3FD420ayaY4ESCxNBZyT0TNL1lGSrRPDPZ
rMI1t2dfN04glnIgAletf+dbXhQA0/QrLk1XWF7iOJUGH4Whegd8BAVcrqWiS+qv
NJva+Hbotqm0vnp6QQRrRJZdiJ7WcLRl+kBcMFQ/eMqCIFVmo1hJD4ropt+WHors
ux3LsF/deFZk9yhoa52FEtwklentgGXpzH0V7CKrqgFJcRp9+pxPC/fll2KzfThh
l1f/ovR8nQcqBM5PRgWamO/WhhAKYhRWtCzTmE19OpNkXCoTrv7ONzNxgEgeEHbf
Wl4PdMrgDg5EZW6gpsfFuoY5NAmYmRv2pL0Qz8pPY+p0I2EP7n625tOi7x8q3+PI
/pcQ4XjXmfxeWPz8OJE7eTv/1xYy3WXOpE/L/KZfTfGePuGIesb/PuWLTbnCbokU
93okK+bH5GLDGFZUYkjQx81Now0JXQcyM/UdCDkISjOc2WYskkoefGn2rgqQm3od
1FaeS1EX4aXaI6e60xvVaHXasEWlsFYb6eexdwjAV8kFIolmuDE2m8GG7GoZv2Wh
92Iyfc9JcXkQpB6TtO+BxLYEugbMCFQ1X8ucytLx8LY9PigOfxqBTAZK+II/RgLb
Ao//B9Gk6P0y3hoU03nV5Lc7X7UmoDe3HmabLTc43VtL8g7MQPM8XNcS1CGCcq0n
pTI1oKQ1VyxMWIMsLKkCiV5NDgEfs6uwSYOvBOkrlEQ/2IuWhoCRYdEJadykPi13
6nD2dUO3Na8XZD7caijiYnLTAAgg7fObdZ+FVBzfT9HQrtqOlESriz9Cf5B9Zkem
od/vlYO9wz/VXS6+FZRkBVBCO4MOCwE+szFM52GIs1w8UL+J+8U7SRu0et4zUSAf
RiK0ywBneRW8iM1FRBeTFiftxs1G9GuGIOocR0s+Dv/Ou01QqjhFuFdivO0ZNSWX
x6UxtEOxpAIos5rjfpDR5Cjd/YLGrpWmV2M27sntu/zSm60PWRnU2ZqSiGoCGycZ
ds0QJkiVfJHjq4+13KMgBxgrLrlu3PoWNz7FYDg4BbXXehL0mq/b97jLdRRzQJT6
7apWZa8KpgUUCUX0fp3kyqj/b5X7Iwe9oUV7fwJLhZSg+HWyfOO/yM7in5kXTZYR
cugzI45P5MtRT0sCLThquErjZfuro0eysFi7+S4nqXlo6hte6NaCCsfw/lXyxUZZ
eindMUBUMu8TtV71mGi5i3VTw5mn/4H4xe/+8p6p8lQqBtAz3rpX/IDTeJ6DGEr4
hfNLIynGEfb3PWWp9rx+ZcMV3YizYD/rPY1KXiMwHuYLOM7pBVuJFb9NpnoYBuTW
7QqP7wWD6z819PNF/VrOpfNYneE+rPkLq2UWzSP1vHoyVfrSLU/tbMQuLw10g8gu
7xkfeXxZbqtGufht464RkRjE7GQV4yrfdSyk+DCvs5FvtwYV7uaTh9Cqfs/WARdb
8TLtLa5YS18Jix+TZwd/eTDp6wrLxDQ7Xjh1cIlpnHedT1D4SEEjvRQCchiD2c20
1VQU8ZepykEkViSGupnpfDEXESZmK0fIZ6u/KMoTzXZVUKC1D4vpdjE/9qxCqjTv
RHG1BaJSBxoADBgTUx6HvKP+wbKkmRaTJVltjzOb+yn6tlLqcMtFmijhUHLGjTv8
pPcCy9+5pIKlV9gr7n2nT9QO7btT4rvNnyqYRD/ts5dzcEM00ObOJNaST+hlrp6F
Auk3U+gBVkNAchiGhy5hBWPA7nMHbUBhm/wFUU0nsiQnWluABPpG1XkgpC/3I4iN
rRkYrDg6/8m5NwWFZpkN9Ej4tg4MUXTXl8/89xxMkH15/wO6saXkf/lHg9sz/TX9
rzCJB19fZCadYt+SZqXADzxb/rEMBYpaAN6chqF4zDTTZAB3S1jZIbQY6R4Go6OJ
4SUdSzX1UaHcZmpf9xCOtQZJ3wbc5tBOugq3VFv92KfGjMLRnYLWezbBPb/K/RLc
42xcLJiI95quV7PQexc9mJ83DH9F09214jIXAg/UP+YYUEGD+TUBPkci7XSWBmZ5
mcTJ80EAwsnFv6MQeCcyajrfnSdooN0XgyWWY8DhQhwbE7wUvX/u89Ih8GYMu9vW
8InxcPFmHJWHfz7KBIQv9t9e0azNrAhyNtXkoUi85mdSvp4cT/rhfK21AJcak+0d
OHzybh49E02wRlf3EZl4ebmlAAjYUnvngHR2LiaJ71jpdNZUPXkYknnFz1UpWNIl
M5Js27VfdVTCkXhCpAOSyUlScaYVywc3Q8jDhx6mRtxlY8Cmn71HqaOTSdLs/Y4E
miJTWe2U03ZFCc73UZHAY/C2w/hKr6kVoUPaZ7AkRKBD7HU0oq0pxq5d3jqkrYg1
ce/l30w0ySjfMNXYb7OVKWfQIWERMeGJtaGs10ZpfzaUeRC686vy4dfqID7VNEj1
H0fWzESmNNOY3q0x/2meVuj/WsTITi0IsufRHSsPauNL+agpataOQgoBn9F0u1L7
xalwyPfSopCP3VQ+DW2NBDeyAiCHo6gCh+Ln+GKkp/wjZjru5RDE4UYCMj0NB01B
S7VjuCHnQOJOr1dBPhdDfSTaJFSP9v495vJEOefMP/5DnM2yl3J0bfKb+65cuOiT
z7+PgkPohV7IUDv8UXkus3WDhqrUlyld22lUaIT4iU2QZE64HghXhnVO1KIefZV0
Z0/L6vKuBGI2TV+rLBmYjIf9LOraG1WBMq8lFebeIRsT3DKQUCR1QUbzxiGw0G2P
vP4VZc8PoajZczULTzaVIMJkyqHkDTgh3QAXo1exnmxhsCwU6D26xbtg1jKtJHC2
fnQWUGBOZecaBTqHFn3R4cgnP1h9Ihsg7hY6/Ah1FiVOq33N+6+JtV1F68ot9jlm
4z1sSWIykN9mO6FfZcoo+8mRrutslpOE3jFfEvsLB+JTK2XoQkGm5TtEiTGWnmFy
x4tMozfB96l9hL6BxnIaCPa1Qqyu28WoZul3n9SlF6tEVD32GIsMA+RU35imCvFV
DJQXLjlRt6b2TAb8nbhjj/F7sezgkkbsCUOfa3z/OzrU35MRSJltbfzG2VP9EBGU
IZB0JyN9inEGeEPsDus9vXh25Fe8bY6PH5XJNPWW+h8pj2DXsBPsGskyNjCdpjUe
FGrfL/tmZn9krRgNuHTwgnEx1PzkdR/UVaXrmfB3tccFLEhpIGSy58PttDE9lVNG
ArnsnBrM3b8H0jUqCfVjeXn/hH+swb3RhuyQU8d7MX9uvSY+r2r/eXjLRyZj2HCS
v/vtFctIg1YdZ5Q28zfyDci+aLLqLbDjHQ60dsCDxcY3tMSfuLzOeSy44/UuEvDW
fs0bbE/8PgYfzBfE2UK7fbk1LKI5V2eI33YjojCmFe0r9oAqQdBjreai/HgT26u7
Xslb3r0sePSLds/eWkWe/q15KfJurEs2NFKMhqY0XWM7hyFCJ4F46fOQdGS1ZMuo
nwiGbCH8aDMNK7quV+r8e7PuLZENSQWQK92GXbXllrkoHdA1850HZqVUENbpjDi5
S1JUSri1Gphl1AHyfzuGMTk3eYdC2gP8F/vxWewmNFY8BP7KQfMU/xoehgF2OtUV
IbVM4P1gxoc/XY7Xm4koTs4ILb+LeTsfSUU2UX0EKottvtO7l7U1VifLXeISTyrP
KHvQK3M6AQnflErAQkTc1Ibi8O6g4XGs5p3sR7Nr1KF8esIfiiQP95XORVLLdv7U
X490kIwF7fswZ0aVtmhlVcFbyADBTG+ix5+UulH5VEWTlmjInnpVmdI14y8OJm7K
Q+GT3H/M39vafbHTgMwQPJ3EfLvTb1hE8VB6CaBXhZL7P2XXHIJJhwP3MCQYeyNa
Hw82Y1NrO1Tr+59dxqXP3jLKkLqomyt2aB6GHyykr1/CBxQMQnyEKYtI59ROJSEH
VDiwQtP6SJ6C/gjTLgPit+2/iVN/RimHxOWCfg83CYtZifBKFtnrX2UCZnpWhldV
LjKAnwe1oTP3ZtOXX4ws9NWg0OYIbIcGpjXwyfgkVooj0KqQDx1WrF3IsfdBl1UR
vOSvxu1onia9aI8+DGYni6RyzK7isdSwtPI5JICRnCJz1Fr/XRxSaBEx8AgG8b5z
To5GbadeiHU9opEgd2NdZxWO3ncmo4lwIsqONKKslHSHXQy3DWh6hWo18+KA57ZJ
947/uqWQ6qy6I5KFdSPSJSovGrs1yXIuBVCJp+3R5PcuSB6qO892va5zxIe7VWCN
9fyOkKub+KUwDvNUCt0omqRIXvbOZICyJC/MPVnO4UdBzn6RhBASw8nKY6FxP3Vn
FHpqg3Lm1f1Obv5On4tLXkZgrhYyMNXOd5jcXhvfjZpvTom3vOOxJ6IIiDtbvGFR
u36VUHOfBvoVrys9rH3aBmQ9A5OcfY37TzcQG7DRna9xWxyDxLKNgUNShwVxpS0j
NNMUMKc9/DrHSyJM0I4t7+95yxi38Wn2kVut7sZlFzwokxYnlhbaRNjOF6GEF0sN
DY8nbbdY707CqYr1Dr1Fy81UAZCMXsBOdig4Ekr/GzXBMf5BqxEzKyNwbKijyvYv
11UH+vkJW70Frc0Jpavz3xwrG1s0C5kePPVxtVgIOFqJHnBNuICLrj9uxG3A23jY
2IJAKld2T2j8xSqnG/6b9vPHkxXwVZOWbGn9mEazPqYWSrBLu+8EhwC09H6M+aRW
IvhUdjuvoEVfXlTr76qJEWS0Owl4HOOc9V3gA9eqgkmnn1/L2lg17WJ+WKqIZMjr
CK2FQYiM1lem5lo0oJmDW3Rvk7vKFkhhzKJ1dQUmLKJoJxHLw/5odtXzNOqQeFDF
ru4w0hQF9IKWJsUs62Nqp/sxL3nu03DiAzuJLGgxqDbFFQA0dR9cUhlLB3eIilWy
QKHKgWp5ILyX7Eve6BUxQvumqcrHiPJBm+5b/mDSs3z9X7TqOPvu+g1o73MUTp7b
uDEQcOxXu7FbKIEXD6Xs0KEEGiSAyoqgPbJkNcB4YjwHl0Kr7EKocIP4OkVe0EF9
LvR0RcF2hlmSDdF7CH6yTR7Z8X//ab8Gm+ReqVMEihTFtXX/z7/W4ZI0CMMxg5mR
kjhuj94a2ZNkF25iNi+nJSpvLwhtRMV+13lMF0UPju2KEO0HPmRpSFmDi6A7u6DV
5LmxUjqp4tGjLZGwL4TfBS5xbpyOSty1zOm4YCHwn7yMeDA7+jbw+7BspK0eS2aJ
sHTkdcZXD5mEs3ZLeo92wRlRpZQYysL9/UZlMZEWJL4blJlVvj9/g2BgIuOt1uMt
lQ/2xOfNR7eg8Ld024ORpBVrVkULjxAtd7jf++wXTT4HeqeZyuuCMQVqKQwhQLF4
bscdXdFWpZaFp34zLHdJ6lQ/5MBVn2Pz3vuB0URBUDnMw1QsNqDSkb77tdIVeSYL
u5nypWb59eHdfm5+VRzc7SkOVBN1e9+Ii/tDqbrZFYNHIWp/pceXyI7ayenPAVxx
RloKnPNIGCqUIwH+AnJWNErAH5VtZX6XNB6j3j2sIaG9h9leWt/Dqd841xWBTARl
TwrjnNURQcKRADXQX4XkSNzbc7lES/H/uLjJe+BJ0OvXq6SP55tVvR04axGF17dy
3lfNE/SApEjQ+fIartUh8M74eCcl1dy2i/48Nprzuc/cJlYUnj0B0pEa2s676H98
aB86ZuXMv2qsd4Hsh9APanxHYDmkt0ko1fSZ7CstwDzYt1S7EjGU1eGlUVjEqDzj
ypv5seMGzR2FkPAqd++t3/nB+A7YlxbqmaFslqQVqB11dBCO21W19BOkllKm9RoU
RE7s97NOuOE//0zO+v+WT2nbmcSrWrJm9e82i9n4wYwvcyN9a417K8Aeu8JGS/xF
ngqYoACowDNn2BdrUhgyI9niaiIkFyOLogQL9YrMwwhAEzRCQwiQkxeZPMbYxrcS
pJkCWPwEjARqQ9y3PFQIaLS9UGM+qoXWasjepTuEWi2JQzhiUf9GOePPJ1oV3wRX
CUviu3cSPEakwmdUitmrjXIAJS52exHlAulmJPjPrjmc0cgXO5Wmb7IfMwV8hcHX
jkzkD10OKje9NnnYQhHwS4BX9YAxmPbcN49KY1dK3DRfunj1Qu3iE0Bb/vVCzYYK
0LckLb3lIwUdlD08basNCoAgNiIhQgQCQOu87swycm2FVE0fedQu8RNTtSqLacr2
LqPmGIZuJLpZinSCpBqZZUa09M+OIGjgbdRO9bJ8ozS4EEPr2HNG0vc56+sMWXU5
acL7EC9KAsYHqkFYJa86VLl4RXltp9ivPZ6E3VmmFrCF1O5VqJSEUwV89D9zcGvC
wQC+3zE0VVkFLblWJVKDppZITBBh6mq0wYJ8GTN809TJfblk6F9W2geeGEet89z9
xaXXZdZPXO1EyyJa/NBUdg00Or1fQlCUXZ6lLdNVt/57PTecV8Usr3l5oIsh3AVt
t3LhLzLkMW9OYcUcQV2zjhnhXgVkcFBs71PlNSilTFPHekWRShxdcWY18yrtQqdU
xTPxbv9OIgwrJnu8fgRAnC/XZJLOVxNub2A7RBQl1BbtM5oZsJBdZGHSvU0a3Jma
T4XZef2LiIaWLW1jLE9C8JzQnUf1h0GQnMgCKSFJKcwVgxVCuCYlAAf+lc0/xSye
qi2LBJVN3jcZ6GQO7X0MQ0UDDAoyUvPut2q1aPxSyEhAiAhEAeErNu3pJNwfr1Mg
ewZTi8kK2a568jvoQF87eUJRLMvfAFVSPgfw0mbnX1rbZWAPtldQYUbvDGS2tZv5
5IqFFNpsruv4lykheIRsp9Z1FJBueg9At+3dDV3f+80C8GH0h3djMUBPcsKB3sKo
TpThK8SQ/bNTVZ3HE9VNS98E9T2BoLvShlrRVW4cicO07zAOWudbaxcfAHxCIKYZ
M275ue4YJXwSlG+Z/S0+tlvRx2tdCdvC2CShcDUFQMe7+1RIO/g0mOSraa1iiN+E
ElOcJ1bkDQINYR+RO3oeSvlBwIj3I6bZuNqpLLSZhPrbIBunsZHFpgTkuIypmIyk
U6+eOPM7CD5lTmJTdqtjUcN7bigDTQPhKiPfYRfWUXuLda+5dc03hVGIQmlVpatX
JBQVpHroJNh6b4xpmdAHQ8j/x57zjuw2Ub6EeyU4alYX5UwHbX08ibwpOc5sFxoU
aiPGxPI6vUlGYpoUdfHgVGZmdmqAGEwhXDuvEavCLi0B/D6j0wFKKvJmubpFSuph
D7PhqyO1a+OO7svR0w5ds0eEiUMAy5kpHtK6nE8pduB/zTDnRlaohXDTAxEBPrlv
HjsOehyjV+SO85gI40w/kqefXDj8fX/nxzJqFGzyVuk+AnQkrQJj30/C4u5kSpBw
hbxC/ftz7waldq64CSR5QcFxB2uUAXwsDOSn88OxgUgkY0Z7029DP79Eh769zSzx
lNjIssMD//L/4/NPr0qrC6qWTY0vdlAGoiWJn834bmOedxgvXKok6fG7s4m5Z3PX
6TUYYhQVAbwJvgFPgtsEWHX98672wvwStzgmEDP/EJzhlu6l+NdIJzCHMmuf/FF5
zdWJk7WUmyVtvJ9NPZVMrwFZtvC0KEwiu1k3Ic4xeKsxNhiEnZvZTCcc9JlAp8sp
m1bQKSYSScQbhLbZ265G94pXUucO9Zi/fZMdupOZzHOSY73UdP1by5u6q2oi7Elc
bMWA0rrwsVRiHYHu9eavJRFDEZardYiqS8F3grSIuZNc1S45XyMoPg1627qDpm3l
rkASkKchzLsQDZUWI4taGiKag7QVvTH4GQ9jWEeKh3fuePMPdfPbcetbGleIZ/sk
B+EWQjToXeycp7FSNLfFCyTQIKfh4sE19Ft7Mn5+Q+er63DWv4lDazlwssMJxnVE
cOmXMsi9feagXiTC8X7yne1m9cjnkcGtCzaXhdzFh1U9iZX/9H9mlaSsTdAa8pJS
Is35m3BobDALQRcK4878A54z0NbZZKQLTW08GTqf43hO/x3Qr2S2/QzeWuYbVfZD
N3KQLg8MZ2tBP3kWWiZ/17qMi0d9R+uN62WAg0ezIquyHpZf8d6KVqjcRkHGmHwO
SlSFdrWfQ/rKGW22VyFiNOK4YawHNN3uBZZHHh8MHgv7AogWhJ9q+l20JC9U+5NZ
AKVZcmRunMfMhxpZj9ecgypftqBGSkOblSo8IAPILGqpjbYjRyx2FQHCAYRcsiXx
P84dIM17eWzUAF/XjP4rBGN2g9AFy0qjskHg6jF1Px9ENGRdYGV/g998ivBZzg+d
bG3K49d/r1Lt/5agsCOGHdE1h+qbCWjIGPclPFd7CCB8L1+0ttOqkgK45bPHMVr8
KNFOcs0GJ2Y9pe0b015xEVN7iW6rUB5hHeZmTAHyQIt+VNI5V3+7PAb1mvVDA8FX
dkqN7UuQgc+O70FIzDPw1WESjgfS7Nka1nJdEkWDlbafCIPys/d/SMGnEfQjOTIL
Iul8uVaNN9Pjp0Nu1B2Ge53o/KVPwvsjBVnRgVbTSz1NnVTKu1JwHVIQRqQ0m2r3
GLdlu4Bd1l07/9sVjoDPL6OuAvcXd9ff+V9wBQxi1BI9vgzjXyuh33p8bSqAOnuX
TTbaf3deBxSV7LrFmvMm8uB9/ESx8YvrKG7fWM9h9gb5sBGDXWzm4s3EreUvxz7/
IBp+fEzXvwdUmg7CCZPPyZuUCdEacX8+g+eDUu12jkEXu/uztCJmCJqiBnWJ+CdI
mFfQ6gF19Vs1UYyVCrVVvwG+yGlA1s1we2eaLvY5C7/7Ku54Y9vdDTrnspvItLyR
gmmISHfuzuMNG00qztOIlvDLaNchF2DnltUFW4rZdMmUik0ZdSybbg/bhI5oWW2t
CVem6WMNUQRWLyN/jfCIn0dVdMYaB/nwcpk/lmKLOCHAyEd0384mArBBbptdn1m9
U/kCxT0Qq8viIBWQEdnG+J6Nu9K3Vam5VTaPGiTz6danK1E+Rq25WkvTmJa0cJHA
hVh8Fe/bsAnc4ldVCHSLtxu7Ugfl3VICcKpe7aq4w6XpzusxWJcYXbNbHNVamUZD
uaDFmof2wQwBnE76RZesS3brrbDxEDwdd5epps7J61qXllMWfzvWeXodS9oTss3C
WWpZzL9qAlc/ZfUmwTTHDgAQZ+lLbGv8Acpx0sNrTY4VIuGD1cOD/RqLgLv2x+A+
cJnA5SMS+qZVOqQsaZU68XWUkIG6CLVPSZZHSSlL+FtaBsVSa9ovDYBi8+xhGB7i
keoaMBtixUlrJ6Y1se860L2Qfe8jhQP33qFv25D6pEIxfrxRBRQFPMh+gwCRASy/
DPDov7g+qz33y76Mz5dwpuDX6G578+4OEgfqBt1L03A95fbbX1gaSrDjztyaxIZH
Hdl3a957J69NXS17XAtQvwnI+MIvR+OZrV15fTea7o7FmArDWMZj9ndMKtv/Rs+w
Sjc9uutoVaDYVIwq8pcml5e9+TdoYD6gDoDYV3/jqMxogh+zX8zN9Rz7FGBICUuN
LO7jhWNc2ocWCyA1oi0/Su6J04kiD3Btw86/a4y1JzmnjnZIA+HdPeWba6lWF87q
UUEEfrMJzB1/Ulj9OoDJW4F0pglvL/OP/1Skk7rs791QEka+nmChdMHdpw2KGysy
s5sSkScI8vCvIGAUeMbmB33GEkrprAPslu6TDQ8VBvx3HVIyeW5qHR9Kf416KZQ3
PmC72uk2pvCYyLbQN1XBlwVsqxo030rAClXvqON1ImNW1KewQgacllhuhDWCx6Cd
MXhFXr6tB/gefGM0SICwBBq6Hudo9txdSPFsIRhdy/sNVkRfptfCA+b4G+M7Nis5
RA33tJV7ZnYUcfyOmPWov0uT6UC0J65qzn7epwp+Rok1cIWdZljavvrGoh8t+dR5
RRZS9uCpxQ/DiaZT1vgONvBH2wqTMmti9JCVvHEAimF4lppVCSQNNtUgF70iFERA
Lb+EtCnbXId0xPt7tKo/cWuqVNsBNFrMOl/bXuHoSXZKoHAmNbRmX0hlInqOIQhT
WQD1WWc5ffHyeEf58PTZK1/QQYctiyjXTiKi7F9raxFqkH2I2BjietPrugRttXu3
zDWcC/VVxiseIGbttNfA8BNmlyd1btoy3ft4ajtA7mcpWLOslJR3Xh63MLkScmDa
k3K+bCNtnMiKWavkaip6DnAqOM9fdnHV9DOM+GC7qelRbCOPDOg5D4Rt3akjVgnw
SfEzul8/Zlhp9asmZDTv+VEZkx0ynTvS1t9bob01zvOk9qdEz1MF6XRMVKOVRMK0
FjVkwO3wHKNfEy7rmUEcKlW2/ZVLrlf1gkJ2NWjumUuz7qji9zvT+ZSb/i2J2hVy
tbcZ2NaIhf1ntT6A2sjIjqto2twFBlzE6aj67sukLcq9HjwK8cHeu7bhZfg9cWZn
vANhdEr2l03ER18xzFzfW2UZwWApxl+RLxJOVn/mwUph2BsTjBGmpMLyJEg/cInT
TEEkTvZfZZnNW+Eclkc27hX5emXpg1LJT3l0XgF6LJBi2ojhWLouPG4lmmUD52lP
L7R6FSCzs13abOcmDFHKcNXcl2oBv+r3A/RhSU9Cq6jGsokitdZX8okyqlgBfMgJ
DGMHlzMY1UMvvN9S2vh7oWP+UiJ6nC3trg6SK8HoxTb9wEWcks1nEfcre0WTuqVJ
doKsLMvgz0Cpr3nIERzVeOBx2Ghatxt9ClctB18BT2wlw5BZt18ClXhYLUys12Cu
ej5VnsxxUOiyg+9DoQE4fqb8I83Cdr95d6BsBazm75skR/2LG5PQUdXprbwwRUUo
1dOuKKA+DF41EgR/I4z0DhTl761yyRoqhjkd9lIvCx1xdspLUhcBLCXR7z4RA5vJ
QixBNS2TG77T1itJgrDZN6sGvhGp/qwk++Gt2hhpT9XfRGXfF1VSCIpc0vW3RUg6
fIFxXxDwIZ3RMosjA+DzDDwrpNJJtq0UEl+wnnkr6e4Qhc+wlRCDW40AxDcUHbFE
M9qniUyGS4ZG5e7AArq1U3EB1Bmxcc99qaNqcXHjLfu5uF+iSKpt7vu1ySIZg+A7
kCAh5mE2vPpUuZkTaNZnD/AxYoSbZnEgb+J8worlP+qzEICUiN/HtHR5kqcEf4lG
h7R2dj+LtX9hWDs7NNbbhfl7NkWYBhpRRz0540B27PGsV5myQESCRLtCPOBSqSww
wnvOe3mIJXrr05VnvselVOabFSE4NC5LAMlE+4MLIlmTLyLVIjnpcGKflraRVERc
Kjd/sBAopVn3YEhWARsJcDJ8ZZomW4d10aLceVeo5BJuVwFiq7/4SwdgrZIQusjO
YhugMjHNY6XS85JilyOMg3++sl01XdtQ0q/yi/WoQ6AJNhB/QMKS3CrTpJklHdCj
KAQ5ZmW0D2Q37WOADExiwpMNjQcx89VPzHxqITbbm2J7uFtK2BD6VA3e+y7Lkrn+
3x1Kj3jdcX43mJj0ECPBQiH4hnfBMSqL5gsDR+YAN/FsjW1p/dj1ed8KzEz1b7Hj
wAM9G4D/KBig1CqGme2rWdFz071pfFyMximVPO8MdJSOYHWHoQzDG6yWAiH43c5m
4bXgu8PlYb7JsfjlyJ5l312ZRG4yE+exFzreQLvorF+oRdRNBv4YHdShxvLkXcu/
Ja7AoIdZM4vvQtlW16X0t/8wxF9dibucS6+kxVP7tIdvI9Q3hIeiwaG0mqpxO4oP
K/4VAAYgd+Yje49YuZPFI/LB+Kx6NVZQ1JKHtmnrFe6qY5OhQohOhTLjlQp7XuYK
12MXgqLx5e2E6Z2sp/WJjXIvcXmpjt6BV9S2s6zyAhYZda3+CovWOgwRTDI+JMNw
p1SeaQDIIZ+8YOdiyYCsSWGZ0qen6pFICshyIATbQRpXF8UIFI7qF4QjLnQHNkVs
MH6lSaWZBlErn6MXWPXAgRVo4x8ZZAz/6HzgLaC2hEkXWRf6QEBVK/f6p1W2wVcB
L80RJ7ZJrAf/2Juvfhu7LSyqweh0uXbeFjeeRK8kir1OuMgwk7y/KB8qJnHk9/yF
NAyejnC+Z21W4ubAyIMq9asTRj86qzLktcLVsNV/GJ+7wVhhYKe990JHaMV9IUlO
eb9qHjP6S2iStO6M5biEO11Rw8iqR2bUAuqlFQ/cUE94bYeNx9Aqm9D0xaUT4xXM
0a7GMW57gLG8rYjUp6HGlO7/XV20ZgvlDQH6VzFwAbMGvGKnwCsB/0o2EZBuHpwL
YNTubH4v9Fgfk+b+DYgotdWb3aIEhibO91PGiEzEAYo57YHji3S1OA/zAxCFVoGX
cDyYxNAh1D8OJvPLs0nyaaXtAOIBwAK5emzrNBOZ0SN17wmfPSDSVCepjESCwfqn
2gYc9sJoEQW+ZLUrLoVxSs/QLvh5XwIFj7kv4A6J/pWG0YMjj11Fe++//EYz+0BC
WRs6nvWWSpj21KmFfsxPjWCcskrWPyBRslJQ02xpBqmYS1enJYJVwCT9dKOXHCYc
YkUwlDIh01xnkGTUP6SikNi1Ho2aQHvlfdwGxsjt8HemNajiitfb9lEKYxmNbnrm
mt9tymx8dm7PqkQwrSpFzEykIjLXVsGVQbpLMC2bF+kLCXcTAo8xZUFHqwNzZsyk
Ksh6fOsKlBwxCo6RwISa1R2p7Krm/LiOyxHWbWCc4JeWu4mQh0bXT2LAeyMOl+rh
f9EZh6UobYHq+GkUxnyZna1hdqU1VTwdYRQnAtUnJ8FSmCeGv5RpXU7TEg0Bd8qP
yv2AHMLxv4Atef5Ka1ZvUmM2eZ120cI16mi+priwtZaU8V8niIRT4hAw2vWyXeuL
IReIMwplxSac7tfd4UwWUGvfY604QpO8nFd1x/45p6VARJIklcMc++lxvtrL2w+2
+JsU1Zy+ZaPjfngDjewmneaPSBFYYWw6JpavxWyOfUTL8JwMnm6VCsxqNKhcHDMy
QWrjSlJvFHCG5dvl58mv4ofQddaVuA5n7t7PKVBWv+dZo84aTe2AdtkGRoOdiw6U
EHVIR/7p13dokpMPhbvS1ES18k3mRt/XNPXsbNoKSgP/bn4lisVT/iaPCb6zc0WD
SWCFm7nUg/bVZB4FDhHeLZaWzAJ7AG+zBAz//8EVDa6MN0+VCnyxxPaRsp2IplMA
g5Z7EQprVJpPaFOoFr/IyI7AjXchA3lu5k0O5epVyyH5Wr5V2aVuQUi7AQw35fyK
ChsZrBIawziH4UVPJYLBylMR2O/JtykBnlM2q0qjj476aRYuqE04LlleRLSawzp3
LYR6XzT0vbkgJ3UWz2e20ZPIN/omWZhgCzpAaDEJ/L4fcQZroIi22BI0kE0QhuZc
UuXhwbaTkRk73vA0d8WAqr8+OVtpFi1oPwW7VNxDg1/xp9S/WTRmL4dmr5lbY6o+
iR375i+NVsIQ5V4cnXEkZAg0kGEJvV0nRWttmjp5RXWC6e7U/5Ax0c/JHMynjtNs
AAtIzqgwf3Z4XbmArHQljeCSp07Wnxuo8YW/0IpuYLXK1J4vFu1GiHovZao3isFs
hd//YjafltT6ufH7iDDV/TYraJY1BLNRU6jSFpI6iVw47W9LDN3czcEMxsSywxDF
AUjpz1r9algVANF0BYHjCb4nY5CtzuNaHasEBYVLOfe8zU+6tO7ovtLmKYJ87XHh
TFG4pqCTJwTsW4s443h2sP+qqdrzqb55d5MD8u/tGl0KuqOjTo6A4yO5KxoO5YyO
Ub0XOj62O9ydydv61XJMxblU4nytWFmfdZjQPkOq7kZtPecfrzSUxhlXFw2wP8jv
h493NLqH3GfyTzxaOQszWKQdwkARPpFvFJClFUVKbpPQD13qYWciKArp5/Z+m3HS
taQYrWhQDgp4Omy4QCOGhFCegK59yYGUCf8o5sfIHLCD/xlb39RF8SvBmaru4tvL
mKsfSlhDVBOd7sepMksRX4WC+FoxIj81/RRhfuPwKfFHt6faANHxfmUAPyK4HUWK
I8BnJjyZM+niUktJiHUDWg1CCX8Tb4q/RTRAO3ij1LlvfYGyeASyjiHl6rkBi44j
/GMDGGQlIxOJ1bvMXaJyvxOk/+JbOrOKoMKLHuTHd1Zr1IxF9WyJT9bk2o89CHip
OSqODmg1wdQ1g53/Q5qtXJgsa1n6ZvIrqPXQSpVqK6iZSNQy61a+NDO2YjmmwQPy
zZgPqNLGn1GE/gzaMgV6BV0cGiQadUVHK86/f8KeQ7PfM32lC1gO1x9pGRflMMe4
F+A/6Y5O2WQDHLE6JX16wEDq/yNlIkWD2DgsaQGvr3XE3l8SBZ001g3ETB3QTxYw
/En+bm3Rm4cpF/lpob8E9oNGRgLH/Gdcr1RePDS63zFtSGZAWkPRgvgMBpmG+Q/T
oO/ECPyqWp7BNbF4AmmG8PmknNTqtrDX/vB1zgHkFlGCer/gJbo/1o5nWEuGoWcg
OI2dSC9q/D8R/qAvY/GEpfRdMOplHk+gGhBXv+rwsw1cKaQ1V5xYLsMckZTqIH9H
+pBMu3kDoddYduwNz69zqT+4p4KaglfT3tiGkWLDhqpQUGb/r9ys6Ju493KCLqcf
+1AVO56b1Qd4VJohoJ3Se1w0Ri+0P8u4uu5LwpXnq7bX73pUvTrRiMmz9ENfxWJW
UMpA2aDZ3f+t0AFlE3ZsY/tOW5v2ERr3PscOWa31l6sxUP9MnxmivhE3u4zZ1Adb
xxxqrTlfAsH44Wk4hZCAvGQie8VTdYj9Nbs+I9J6PJtCs/ZdX7EZ2ZuhLuFlxuY2
Oehb3XAQAAcWEubDZPj3FFHrr1/aHcBo0FeMHPCmWPnACtqpcDRygbQU8YskWEoJ
P0tT89NJi3256Kl2O4cN3vI6u8m9F8Fsqzl1uRTngOCoC3lCxWAABzDxWiEHvGMi
BMQZ9ZCp+5zgU0H824q0cJV8j0SXuJGhnVbSvjFMZXMVtfU5kn9hIvOxSOVVuxOP
yq0dj+fvfn2qnDDR4D+KRLP8zXkmqXEN8O/yaX+nd6RbII/5qwquD+zpbpQ7FbEB
QDK9isXLRS3siWDFvgqFcoExajjR6UWIWWUmSQbZhpEudlAQghMqzIJphBznzjQu
yQl4uNVKSaaHCtvEqa9UdrBS3jsjyKrtKLpEUxNNd8AJwnYdGdeTpLpI6GbYyON7
ao7Y0NA/HxPXXsXsnKmwhDxWy3Rj1nzJzZe5+O3YRwLMPwZ+g2RO8SM1nohekgsL
swI90AjV1KSQmoBDSvlk1s1ECkaxZS+Z2BYoNbZnBTVDTJpPCgOzRrZJJqqan/Cr
CBEHGmDPXhV56qa5PX1/2W/GIDcw+nXbeOxFQa3jJZ9uPzY/2jvWu1t4PJx8Ghx7
74Fyvmlp4G1C4SLB6IQasFAS229iHG1uU2nibOCeEeGqMIJrkswER0C2fdc/aI6v
8AuFPFB2H/k9qXBQD6iknbOi5t+bXn/AjMCaJta4tezIEa3fRyYuBIqLXCGQpZrj
jdRySrZ5HhOq9cizxE2H8a/QKPsrV+O+ZdxtjKSigGmZWDAYBrZqd70qiXwAEh1H
hj8EmHyHbwKRkoKg1ZjpXu+vUt1bvoykYdxZMQq5+8MZBWjK9iX2kT2t5lWQpYdf
BVY3996uuGq7f6xvEpAkIvPevyHlItcQygRHJhq+DwQLyiy0Ms8GZzDKHEvtH60E
3Con0yJ3DntrfXeZQ23M1UouzMyAlinIDALIqoDKnxVX/ofOcNOYLMxNpaeGOeJP
XsGwZyX9c8RO0OULL/b3sWnEuY9UOw+BsasndXmLwvKPfs2G+vgD7+Bm574LiLvz
f5UdPX6Vj72sqx7BRPsJUl2o0sQ8SqMMBE5McZalr7C8ev+Lc2LhZqYe0RcJ4X4v
OaPAzHFjdmwKHjzfA6hwB+XX1om4Dlzeazo05IHqJh4E8OxHQvAbTJAx1/UZRFJE
0UU5YZfwIiK61P6PFVomC4yA7Ol7rmygu858Ki+A4/UnwV/ZzgXOfMiox107PhZB
lTgrHDy10eqacjUVqqxZK7LYhBh74eZfQrMbHCALHd7Ri2dx0OxXLNleNnQ9smi6
RkPRll70hiVZXkfW+pkXOs2WAhGUkD9fSxFUiyh55RcvJSmPzdsB7uM+qTv2L7WR
RQWnT8TIuyb5/Y181kpfhqULlACVLzkGdG+K2q64MnSSW5EocBQksmcWUHWZ6Y/2
ZVTeo4cLS+eO3+xj4crDM/CuHdruvToyKoDTq9O6pBdcJub5smlmLrSqSd+LlDZJ
XbYp2Ik/bHqVkYdtIE2mO/9HTRK1GfCzgANhhdvlmnwKb1gIuRKjecgf9GYKh38w
WCpZW09qbRSQPUwCJ+Snd7lfNn6S7k4kI+I+y/BIkdkqI3pXQSAV5FKqLECn91yq
plwAfMlIqiKZ7r21vxGI0tqE6w6mBjx9YV7BPdyr92wappEk+qXjsYLaFQoYWkb8
r7oCjy7jgaOJXi9tv+EVtokfxvu7HEYTe2yOzddofMgM06dH7OUyheG/4GoyBr38
uLbuMpJ7+QDp5t1XklxhdwaYnEowyRAkjjTzDFRPjuzFbT++CatTinheqltAKMbI
eFVmmC+1bR/6qeSkY33PmzVp1uWbEKY1NUCaHFNlrmVqKi7sNWoYtFJOgpt6nH9q
M5Pf+eumN/j8H5O0BxNiz4JPs5Q7Jmbt4yj1oUaEPMSGO7cXTd90/3agEjzp20Rb
zDbt95rZ5Ki76gKUKJwRyhGDwQvdx2rsaUrhhWYHZ4bMID8hEQGWz5lG7qUKbYTZ
XP8xwwKZDX/MGXJCpHW/n826s2pQxJsBq8hWyGQUzbxAHwGVD6tKqX6bKWOXE5k+
8gOsgW5LtG9MqAPGYbDSs56PT/Glb/6MAOdN10Ij8MmBN/QTjHzkGdwHpe3YcS37
pY3oOeO+yMRhBHQo8GQIgWXm3ASAe58+YlecOFmLe/eHRn9Rgwtyhw2mm1O6xWQV
9uh+1nMaAHkpZ2gd7rSvn2F2+PXqlWM0RyHxuMfRvWTYtkFug0+xcqy59+Zn3Mqy
Gt/OQ4fO0Z6KAUiAjMGa1/QgM68tr3EOKoXOK5/gm+4Q9GWvHWzCRPf4FN2hLQjk
SlSfeg2uljzuGJXhy27Vss/X9NAah2ZNb7hKlw+yEcuVq0Xh4+VQJoYLeNAcLci1
TvcMb0/6BjBskI0/gK73b6fLbhvu2tn9PCCP6n2rpDmxWwvq07Kob+6yIifItmq9
Q/llsj8zJDscKxfWgLV3l2swDKv6xzeA6mEeXa9vOg2xeewrOpMwyISQBcffZWUT
Cti15QYsPchMAWVjIOPmfiDuSN6jFl2ee5GVH4FHVwPgz/32bOBHardJTEEjUAbl
mDsFTRPsBS/CmVLokPL3vjwDMgpFfl6iYBt34vqAO4WkYDGhXwmBNz13abnzpFR2
hNQrSwksM0RsGIWFtrQJwuyXxjqXr/k1orHnELyXVsOS+hUlnaUFspOUTGIpQ08Q
b3KsnvvVxY5bYNruHsTbb/MhgKYOCOZgCi7GPM44NnsXiraDTDDseVjKaui7wkHJ
BTvSgWWAIQpFsb/vCatNcQIY7L4pWhlcvRrxXyaaBf7FKNsSdd67mDiUdSl+Ze4P
r8nO19j3A7JGabGXbHk+DxNFATKROV1szf029f7vML0Shk9EXeqTEGKIGsBvXk0W
4QRjZ8JXMU5vKtCjE/BumFa0/4KlWDvX2RCMjC+LnZ8D12ooFrQUW7IWx4mt/PhN
SoaBnM8GUh6qMLFIpH9PDR/Z6+GbZ8NQoINLwmasKJcWX7B7us1TFrgd4GZ2Vivz
UD5c8YPkgd89zqwzvajiRXsNkvLoxrAMVB09u8Xeho16yU9fuxsta9qPg9zN94oD
6wun3EhG88qX+NdKR+KmyBk1DAB5mZkP8e+b47A7y3U78BOpXoM0WQx4BqpO40tB
SHRNeb7rPhfH8Mm6ayPN0MnIRkrMWZ2abVm+GrOgXBAtmpNfGTfoPtKdVOiQUe2M
Hfgg+X3IRWbR/BFMD4rKP2gHmvZe4xNH6kLzsDcT3otZXuRuXdhzcBSpBZiBxEwN
KZKQZPh2PyXxYAXO3b8OpWXm9fzzr1IRKihMcHgP2jqlwYFMMjnndmlZx+Yv4poi
DtYaTSQn6hWfAlPwQeVpNfyyLCUTISzHfgclTH2B7sBUNYExZ4sZl6tTEKhPcllS
hv1zHHlZwzwm4W5tX6eCsNfWDGObp95wZ/7UaMzeSfiHbg19acyHJREKCcnf1Dvz
UbXeB9F8XsJSrxoJ1QU633ku5fIo+zUZqOKuAyfc+5NXNVrN2KjgBnZYudRfyTB7
QIdUMD+Ng+weSDO7aRclZ7SSiThKm1vlBJ+CXCWhezjFA5tRZlefhpjcpMzQYf8U
0x1WeEOkdxF6bWbPJ2OnrcaRHkcxDKUDIRuWInG1xBOt+d2yCAfGij04sg5/cccF
d+8G/hh4WI9RmWHEyVkxNKdMgipdcuGVtYTH0g9zKIh8P85NfPzGF1I7emePROvQ
HYNkmuYDckYEjRE1K3KNTyAuCZ+OgI4GrrA1p+7qg5W3UxdN5Rt4p7dfPAxk3MHM
wGiXtqiZ6KhsotcRFZ9fqF9fVaVPMLHyaqcU2SISd+rPQtVd3zY+qNvU+FbgXloX
rBk93lERRJ9VFjLT7sGhAJrw7RCCeF2GqSOsmfTdagmgSwNPxcGRV1fg2kiPwsxx
5uxZDhab1zEwmPhbdIZflJ9dXdjy1T9LOQvgTjOoeaAqmraDQEnzC5mozjD8RBt3
6f2OaMiiufhD6YltCB7a9mMcUveMmbVDvCIIFt/OAWCYbG0wRCln1cDrq0avcaTa
nRAYLLyRBqQJh3AdTdzNg/oWyjSuQ86my4nDs3lKFXv04yaAJ+nLaKLVNel604GP
jPIqt+p/erFnJFSRmWKduBujfddBEJfYXwFVDuH0BfrUpJF3UivuwHvuJdqO4ZAy
URJqn3GJcVdoMalMG72hYEAHcFsRlG/VBenR+H/W2+4qrD68gU/qTDI0tWEgyr5s
TuceADW8s9v3cXgUr2jUeV8jQgAMAGFBXeehkPyA4d2BuW9QvXOdAxT4C73V9PQe
YJKmTTXNBITlo6XS4/KuuoyCCOA4fSEoYGrDIn3DgPo9uIDz/3NLuc1gJheUveBx
oXuLctu/PcP7rEGvr0AkVOF+3GeYOsLQQnNSNmX5TGBu+9Uzc2aYGOLQ+46giUW0
q5Ss3tueCkfSZz5EXKqgGIOyEn36fGNTfEFtrYPqXoG1ae52v58xA9M3ztCFzl6J
i3Kcy/PhyPN2V6LMzfTfXiltyZcHG4foZknJCAs3nkDt6FWk6PvIqfS+ab5JZRXH
Mk1Y+NYWV0kXZAPMH9EXfL2WS3bnoyf9Bl2eXfHutSccjcEhz36ojqVQaf2aTa9S
zI69wn4qUIWzsl1VIYNmMtSz+sRIdh1qTdvwSD8JjrTEGdOpKI5mMZ6sW6dKzo/e
JtPhX8EWCAaJguvZooZE1I+uHXHkOi+rc4TzWXcLYXWORSTjIv/2GVUWn+O3xHB0
0WNlhHV+nij9HIsXf/wwAQUZmAXQ2QC+oIAHlBy9kns0AGXaD39bJjWUFoSraCjF
o3PoqFjwSiVzSyXrgIm6iGDITQFfztp+I84VTGYlWW8kh2QvegepdCMh6ac5SrMr
qc8mQ66VVe8mShT8VYLwqHxM63WV1ESyWF7ex1YHKwXaS+7ue8bQZP9oeRiFUqQI
f6vVb6NJeNfL0jIoBwK8y0KQiBqfSaFvbCT4wVzB0230iYfp4cFER4XiBZYnPpnN
VeLkCu9WObsora5zXTADoUaus7GbOEAjHmMMRxqPSu6o+phdfwg9BpzPJGvHcpfS
1LOSeaw+OXKdgf8N8aU/EQw2qwPjmK3j7kLseGjTZCV5Sa1fPb23kKK1YyqAb16E
YygWmrKJ8SWyyb4kA0sMKTdbIy6GC3xyy9FMZopk6NihD7tDL5RQR7XPnAzX1wJD
ZA/bPhzBs3BO0r1ZF3PiwFdNgVvlOUzs5Bd9churejWhm7twlzbrIVfRKYkP8XTL
tOhWxKagEMeoz5QX6AmaNmMHao9I98hI15AZs/apnE17zOg6sGBne8+8T3U9Uowx
Qw5oKmQVpy1bmVITkDHLyadXmmDXz7C9l4bJA5kJfA1f+X6e6us69v2tv38nIdRu
P5h4RtvL1lVUjyniU3uwOl39ltIAmBsLYpcbeZIuyoaZ7ynt9hCo+WGnXPb1iFNx
EWe88d8ZXjACnpOfUvxEgRLhS2Y1MTXZVRcokxEHFNl20cskFWUWfWRGQXXX+xVK
lFMLaVXLW+eaKE+PYytVJQJq5V4fhIeYHgDqTfkeb5SxUR6tfN4sWxGuzNOSO2RU
Swr+mgY+up2FsxAYhbo4/KI9AoI7gZxA9LJ68LHisUoBlwAamZLE3cpW3bh8/kPr
WaaFiMFnRbmS/j1Owh/9ZFeN+T5/8mLJOjzKNW1QjU1BxtWR7TTt0VFlJ6+70lbx
NxJDIVaiAFPGzDmqWn34TDgYjoo0tg4xd9Mx0Wzrv1sEk27gUN9naGYdyzdqTuyu
aDUwoFJhFQmcuK5pdM7n7fKu+dtrr93+Ay1oagMc3G0ZWH8nTbLtgABash+jS93K
pTe3qdz7bVLyoIIN5bsNzB3tDaLKI0BSHD7vL/ZoAvgZvIOBZjaX05BVLEamnQoP
k8kVa5CfeP5qtU7xz7R5LtkQdhbkNjM5dHcUefshj1y+wn0tgtQ+ldn2nJIL3huB
lT1Tdw7jR23zpERbw9GUMK3ClxC2YvK2peNzSNE7zyRu8sL5XpaMeiq3KXmRBHs3
6Qee3zkpVw8t00zE6EvP6PjFToh+5qhWidxFiBWj4wnki5HU2JH0DySIVQcTnQXr
cuU6Wh5/Mk0uLTIAKOu0+XzG7EuCBrgXJYksHtlPm2dND3jx79oeNXjMt+wNH+BT
/wKqI6ML+5mHRcVnB7Vp5EAKw5LYBjfK5sskMjVkwsUXyxw2WBgQDWdUcwwMbzF3
cV1k0n1zrLfFp5Jq+OA/k2A0TEDfVo2IZzv2y7L9JO1CfWJMJj5vYKvzOizoy04h
bMTgKN0HaH9Ft+zcV/z8KjOP/iTupToW1ne/0TvFBPOslmki6WbEEEq8lm1k6Yej
bCWS2kY4Zu03ygCokrM2KQ/7E7DDcZ1dHcVOQ2TNU2vl/ptcf4RYKlagwUGh5fmG
Ogn5bHNlRpSVvNsRpEuqU21ePXSabOorFdIfAKNZfb+mjvU05AiD563csKZbnLO9
z5+8EW5US9ka9V6tjEjVKndQgs2if7sQIGn54YLx1avGSTy/QGPBIkI8zyQs4c+i
dKyecNVZGmC5xWVYbDTL5fVGNw/pGk99NwBmVx+uUCM0JpI9kUB+KHhSLx/KYIZD
TGFs4rZCUGUUAyczs+x7zIjSJ8jjGbGjJQqHAJjFV5PuGryu0/o9FvS96UX44ELV
0XZtsmegmq66dNPLQPQlF9PIOzWh+oZ65SIHGTDIRVsXJ0UlhBVZI1+eu/by40wP
Tlg+ddVlwhJtpxYf9moocle6nHwO8o9EFDp8P+5V78Qg1BB/6OahCOH5udBjRvuy
JkwRbArQvQO8fbmPFfOuupjC5u0UEuj2O90OKXR30YFY3vrBGjnZl660CLR/B1Cf
qQcH0U6l+ZYxIBv+r/OUYRT4yvxYJdx5D19JpdriTBdf9ZJv3Hekj7siW2mAWbwD
40z7c/8XyLfphRZUB/6u9suHPFYZZK4uf3fi+Z8AZ5+BVn4cZ8Una3n34xniXHRt
nzO9E2yxk0c0BdYCo/iE26BkZvMcezg8UXUdPxg2ZYKWEyH7spKjeWKKDJCIcNKw
crzNK58EMtcBCYGwtCSyLG/CeoXMHqy/E3KonPCi/kOqI59OR0dGLWXEwyuUaVb9
Tzs0Hahvp7qT20Kw1r7O6hbJDfeTFEYF26LAwzQDWmt3SDsieFm+iurDaWaMECVW
z6ZWn2irBdq3SoawScT9mD8/AHxok1pRisCJKrsZXJr+cMXNysd2JKeyXA3uFAue
L0joVAsfSCR+EHzgRv3yryrB6w6PYO0v0mB/MBET87GX1WVNSpIErk2DhyRLRG7R
Xy8d/b4OO4hruFjhI2pUn+SCK2WLsDaFcyHyfTFqqBRLHwJnf4YhilSzeOcdS8Ra
pVDvpUz3ujuaqKNb4Cg+htipF7+LGCBNHJbBzraIfn+ybhPbsl9lUIVkRvUSe8aK
0jDBAjJ3NKpeyHX9i1A4xczNj6VmLrlhpbZICKQExVbRCPkjrjHNyCf1uXMOY2O0
6dyKdP83cK4j4/lqPy9tGKGRCEx+8PUqodWhWV5qT7A3J6ANjE89+nFQNxCSnja0
/nwRYKCGrRybD93USsSX4aBy5q0fRL3EBWawU4+VqKgjuFlqYMGSIjvrTr8OxfLh
3NcgmbDMO5nT5SQdvi08Gs8BfU6NvL/qzuTw5hWqIVqldvyTz+L4p+a+PkAxXedQ
SRpQ+d5/lha7T8OroQKR1dOx9kS0NGvBXv8jLvMj+5g/nVXh9LhCnyjdIJWZ+ChX
lhk3Ks7rGvxqjjYEwpZmmjUW+kM6bGGUnDvp2KZy6FtON/H1TD+VLSybXiWFSNdd
P5Ar+ex2exMlN7JqljDrBAadXpUDHDJgQR/9m3WFqxmWNJUZ/tVPGDX3U+Fsp2iC
arqK+oqfNc59reEB1K2EtYoafXvqu1TfFPzwUBPSlt6qLBdYFz0pAikHHP7FYl2P
kXQjZpSddNuR/u17XzwfUq3NBOutFF8Hs+V151T+CnJ+O0F1mtrIm/peDaGwpz+G
7ikJywETk4QupNwATKf1Vp+xB1X9b29cC+PWrzR6xVc91d4w+t4OjH84fGFo5bqQ
Pm1yNNr5jF9O2c+yui5eVfTyd0RJBFS99U2ez8NGse0vfWeVHzUZRTWg/PHBJkmS
H0XuYiwUkSZAQblYUU1a1/t+bClPM1tyfQo+WfiwSUMAlS4YbFoVsf+wYPYavyh6
UcS848rTlJWqGiE3A2RraZTSPOTIsrdIKEhQHVPxw57sWDZVLyIlngyJwCAo+1xM
vmRNU4p1cAJssj2ES7AFJczEkzF8wo/wpSCgJT1KCLImUa8a0fOaKd8b/z56CZEm
Sw5vXhh/ricaAv2xjWZvoPZheLVBgOOOo0umUMwODmzq1XWPExav2KybIAX/TE1x
aEZDSUB8RBFNHRHe8agTKw4IW/3f2zci0mxkZ1JP2jdo+IEtAZLLUUmvt1dPXHUN
PfqXxumbv5SsYnv4M42XMH4ZcfLaK9SQyG4q3BhoCtrQixrBTSa6OvtqMoaFbv4l
P3mtGV8oZ7dvwmJR1mNkDdRRZPgy0GcWUl28pOCXQLpoJKbRpeeFjEO2US0GPNux
cW1qqT4WVr/uUUzvHwZa4tBU9S323BGF8dy5IURWG1sc/EzKAjGu68myM1kMxIj3
Vla+41r/kO8Ajd445R0BC78gD9BskseDVLrUL6hdItLTIO0U5oq01CtUnJUnpEgE
xdy1DbGCAjIzx5lxtBPQivCAOEePJSwj9gNJr1jLuYYDyN9dkvfnDcJTT9gM82fI
1GsQ8Pd37hQrQ5sG2lcc8UpDm55QvDDVTPKezbmGpnPBOr2mKJ2zDTIs8T1i+n2p
u8RT6s19yo8zFjkPt51HEQiqqUnM6HXeBN30b3bCohVNkeOYqlWHqLTb0CKqaDLG
QCuNmW9shtcAkhLuXhUv9dQzifwcWgiiKxGDA0hiiEhIzN3gryhiCqF2vhbVqvlH
nnVHQ7U7mG5pmIzbhSNqh+xEKK6a0VwbTJUPGL6CtD9e276/gpAj/Q/hsDmU9gv/
9krudiNwbVdUfgAcwKJQJA3oqoGNTJwHAdOrZnl+eD91Qa8DF0vRqoUFlwxmudDm
bMp/nEY4JRcj5yDbXkYOcWOCz+KQUyVgyZn2clvhkXhyTxk2BANTqJkHA0LDA3we
ssaLWmdVyx4HdCRCHZlyrli1LZohqTaR1MGkrQ8wm9IEyl1FhU7tsXdtCsXbTwE9
eehe2Ynj0/lGBqL3B12E4OBF0dToLPTBlccc7CEw6XM6vV8NAOizfLRguUZ7YSG0
TA5jH4fPzcc0fbJpKVjghSxPR5MnM2N/fLSZAjtGDGmiyX0Df52/W3zSEM5OhazN
NxCx5Tf53uLSUw1ik/VZJ6vuVaq2cWNMDYd82umCz3Pkcp4zXSJ9Mr3/mgbYJe4M
O9B5EEKOUC691BqGpUiQJckZVLj8HRPhbZYpcfIdRr1938WAI5UG78BsI6e4YrVD
yHBXN4ig6t50RNP5H/AiwGfS3S4lhmQeRyD5cCunqJi8zCmE5rOToaFNQ60CcjMU
Pg+AJizKtwmIs3jjWoCs6N5IPYR5gTSstIawDagyqds8XzpnRUljtevG2UccXMHs
jgLB1kE5nzRWpLrrH9oOkHalrK9JgFas4Fd/CAry+iWMt54YI9Ayxi2TwNIDofzd
igXlE+RqpUoLQ0pgeDWCW6GZnOScJ6TrNzoQwfYw3+kmcFcz5J890TZdobZJ3P+r
+9RwVHpTZw6pd9axgQTA86dXE3Ef32aCTM4eJV9AY7HmGge6q3+Aq5kZavuem8GV
cavAdHSMedeGAAErk6jUGBzKNLAVLNdpT1aipiODImHcH2j74nPXTYYEa8DnAqiG
1y2Ka8DL5J4MONxod7bFGn+pWBqhJfVWxW02+62Ji8ZAwdexK1tYGrmW/oggnJQF
aOg2y2GyQz0PZ74wD0lv0v3LqC+/REdqtibAwPrnNCnrky2fzLCS4ULFX0e6Gcr9
WMab82OAvHz1YEAhMPb0s1Col4M2RTx2tsBlo3hqZbcd4R39eBJzAct84druaQOE
2/HYl8ammdICZZqnCYIIKh+E2Byis9ZaJux8Dp4TEh0C0qUddhZBr202Il4+TWUR
fzvR8sil+34EDb3BJwsslHQndcPEo2sl4UKUaVoDOFoU/DvX5vcB2msF5f1+1XzA
4pqORp5tXtYgRMfSFudhHVxe1riqSUMQk90/GWpA6MoIrl2OydZid4dIrMJv500U
wfa0ywD+9GwGUUmB+H3vMzcuNn/j8GDMe9GeuazH+GUyT7g5aigSjEe9K7uex1pB
kte71dWM0rM9TpjKCAbt2WTDSPgMx/Cc8JhEjgsfDDYhLQIUN/AFpKALH6XTYCDt
JcMajlgIbHyTejKvjHGACjY2l+DSHojJHI3Wz1a7o1kHmapw3mCIbLwl/Kf6eMXu
3HF7r/aER340r4Ahwjy7a9aDaLQTsb1BMQHvP4Nsoo1CA8fO2rDACc5bUnutCpVq
waLAfo6xTRPRQ9sRV6rF8qDkmA/LSiIgzfP3e43gKiHL/LL0eAzGjncQpfmhyfRA
SZ5iZ1ovNIe79+kmFh/KVlSJWcuefMVn5AOaB3Pyk333/YppJyRYOwTfKMpP9ovX
TWzHF95G6dRIcdc7pEz6rqBnLTDD4GJ/fid5H+qb4HyJgF7e3s6OWnPyxblhtvWX
4mMxeFCrnLpUtk1gBtItdjhQum9QIbFBAvyPUjsQLlywOKOO1EkNYfvxTbZJeRBA
oi2WpRlOUjigDcZRa4ae4YjwjjWfnklDK06dxG1icwz3UEeg3WfYS96YgnkoTuW0
uBQtWra12Zy359+8PfrhoRh1QxPq6OWtEFqsAyDFuzi1hT5Fm2C16NWzU5VOUKUZ
6GrGCgwzOjtDlS0Bue3+32WTur5J5BcgYn8mIl019hnw8DMUnf4uFxPrq1kCL6Xb
GtL4kT/8eyDp1lwu4c7FW1+OOff1JmeLEWFeIhch/tjFGRDAETgz4Af+OSurujxu
vOQqzBuVqsksUfk41bDWdCVtQ1LMCv9dPzdWEP8WQRXcfVgFVyXkxIIgPoXQBk07
fSTtsqlOOErfM7ykJhGfIeHmgBQGiguNyna3xp/tGXg2Ffq8EJfkrX5KYcPSMuq2
n+Eax/ArAMD32rUhfPbcA0oUqV1C5jrb8m1saqT1RKLohfYm11sLcY50EvR6KoOW
qGL8tLo9uwbNCW8vQMBw3UCPR4+J8oql7jsaJLc5PdSo9w+EZzKZLas9rk/x5dSa
Zyao2nkkGurFaJSDQe4gwWOZQIb0TZR54fXqzwifBg6eKCMxyHg5Y1y2Ow1n5AI1
kGXAT1h0PeozYtbg2s1x8wATtMnYP+RC/e3TyvdUKEhsb/7+29sYSMoYK0DCWgK0
rTFVx5R2WVdmNjhwXBKpIsffLix6HFhKd7TomvwjPLBvoTpIHuvbwCvJD4+Gi35s
QLM2H4Zdcg7c2nmsmN554xXSkByh7yAwbszaz4mx3WVZqGPzhmjqZpORLFyEMvDT
fRfv+WG+2SPhhO763drqD8mDGIcgJVSHYRx+LxWXNbxYoehB5Zh2owDK3+Yr4IsF
E+nj5jo9Lp07ACLyXMl3Fz+NtAhdHiyGgrm7ymy4mlBnfdfmLAmxqbVRKixfawKq
ybaGg6SXImISYwi0ZQgBnL9A6F72z1ab2C+iNh+1Zxz3gV+2yE9TpCJUvAxc5Toz
tbIjtRcAUo1Gxpd7bpujIsw/E0mUzaAoSVnihMuKlR0gsabpO1yVBhHe3JUucqUK
AeZMZr9ShYft1fhdLxkAb5/HRcfaiU+S5x1WouKIT2SPXZZ9iW6tXWw6KYuiTWgO
qkfZGMqpUvgZlTId+p0KHqO1iANLd9aI5T82TWqdBmDHlkXeisNYo4TOe6Xt1CUh
t+u9PZZwIvkPbN54UENLrY700gXKtwvK/Nsgw/j0HIlsSntoCbPvZSLVVDUnQDgo
y2q0QmupyJAqvs+X16f8co0syznmvLBFlRxBFRv/7FKyct9/uNO+JQdVLWVSJvET
uWBcvo8ILZqxhHn2Jwzfg0xJnTy4iqZEr+YzxY8e7hu1Z26B+2l3WZ8Y847MbEHo
ZqrBzj1tdIjqbYlqSQlcZtIWIAHCtFt9T5ZfIS7JtoXNxmhfhMtZ3Z04v40OI+P/
7oUXwzhzYxstEiGKpIZQ7CLJvVDATHKH23rgHtns5Ts5r3flET/6pr1uHZY+Z1gF
ETtUOT0N1YL4dW/YIebEEAqQJlMRtIvnDRrjaCIi3pATtsW8YdnINs1dxf275XLF
jzQD9mfoPCYLN5Mpdi8DxQG/QKYKZhs5TSKeZxzZTwf4NWNb3PHxUPQlj0B0DUnS
jbFmA1jgI5I9Loo4l8URG8GlPufP3eIOaaS/QNfZ0imY1XNuk02jxqPA/gOPfmmo
YWf/fk2YKvaKxw/d2Lj+eFe2rnuN7yudVsLO7dfyv0MSreoYrVfdR6+Va1kaoLEb
sztIMA3VsTgM02HlRikOtb5E2Rn/73Hj/z24Ex2kQYcoF+ntx89a8qcIXruh0tw8
5I6V917JxdualmOymDnOkD7Cd+UrLHlfLnpFukCZq/XP1My72DAfAhcwVKj+LWsc
i1zvhBmBLNhwfD+5WJNyLfxfvxmirdnFo2Cr0jdXdmhlnmqZSeqxCTQwe/RY3w1b
UAGxcsyhfrAwY2l67+97g8c3T+6v2+D9hb8XpwscvcEpng7hvRHW7NjI+Wi20NDE
C2M6U3PLKBcxtngNhUTVDvu/x0ZG3MG00PB43wIKJHwTAh7mcsUlLZFbE9+YDei7
c9OjYKzRPeRI6Y9L4FUSlaUFrxItnTywA6OWuMOkE7fWlqGp68RA9uTiygjJtM06
6NbfGAmYc283Y0o6KZhAYJ1h9i/UXuBxFCS9yM6hGEk+uUscBYiADTfT9Z2wySyc
luGqcamnBJElYiuhjNBYADb+TF79f4ojQTV8O/eVXClFGgOSc36b7EyzJ6NdP6Ck
yLptx+nEkLGTrHFmR068iSnfsMGXmbguv01sNgWsTput2b5ZquszQnVixV8UDuSg
J16tHiZ4/GitjTaIBi4XRBV/ZwbvTv/89BhKHt3zIe+gyi/rYrAbRQstZJHpXvkH
1On52XWxtcVvAhR//tRgfe4L/AgPmOl5UVuSjpwrJgKHsHqs/rAEbAI7uQVuIhuq
F0GisyAaNq/4rbSmVRUcYDZwwYTo7uibfetOJPJyPYt7dkaIXRtqsZ4sFjr6Scn6
M1pcKaoiFxBe+SksAg5qwpUIi9RtmEIPPQehU2wA4XK1x3xRXM4T4WNP+I8tMwx8
F6Lrty0nomwbzIcGatT2Lb6IlBpobQ/uy6X2vpSY0ErEPN5qEzxmfJQyNsK6bhpN
J0UKMndSskDGkRswpyNBurvopjD+3iPIpst8m3GDP2W4bXiPZTAXLXMMRfeGRxOF
3/2vtoIRF061K2SfoMuaprH5CwzTskt3b8rk8jaI7CYCUok8KCSFsE1MgH0bOegy
oCj+/IrqLnYJCMfzo/l0JJhLC+fMm8lBmBdxsk4Gq3CxbwhJHsX6ruPttFBKAOVf
os4cFJbTtXojVboCXphQIvpFC2apK+Dg9/ljRwa6O1Fof5bhFyK7JoliJHZKMP3D
g8aT6VZ5kBzD7DXwKE9EA4FiEEJ2moNVi28ZSUHZJAKdujx5ESVIx9YdHz7EyQhe
uY8Wf4Z+P5quz3a25yWzf0axYOnsRrYBtbhH+SVMMQ8QIYuTs1SstydXLoScLwgh
lxZ370e88b3664NOfoZMX+R6HsKw4jgN2U4C2hiiiy8c3StK6zdVGVFLx27B+QS1
yovCfI6nST7qCfn3uMNDxhlXByNCiTPAZkdb0gMo9POqzGpmPANtDg4yD+XhxyoR
ighKi/Mbovi2eaZMJnyuO/aMgXZokQXPTR5aMxJDsdlSPKF5IUkOk2vL1iSfApkW
5H+fmZlG8tXExFmJAs1bhyaYPPSq91F+WPPxz2INftqj3n8arH2+Qb0usRgZTeSo
lNKgJXsLFZ8Pfh7YALGTIknGpXmcvhtvS2tPfPy9gP86RxfmpuZFte3FkvwO3lhN
GP1EZzE5zPoKgA/3634GnJbwTzd8E1+H1uHYnCuQR1SPgnxEXOU3xlTLF9Esntb5
2y2CV6F0AZLhc6ypIcz3fH7GwHh+wBoDyn+kLwDPuNIHop/8f3kSUwtoLNRtURNk
3/omw4gOBpOtv0RCXH8NUFwJliz+bl9r5IkYcJAWuxQ6vyytFXE86qwH5bouHBiz
eIeopSpKXR9gvUGLPa+5m2Ivh3WXLZEY2TeUoG1AgUUy3FCEVQgdffy7WdD4XESY
MJwHqX3cwevlNbbmwFGDQQQIEIhsDbOUHpy1gGEKuEE7EWt0k9O5f0PSish1iK9F
MUSteIjv5j6vnswGRliID1vNVQpLfv7XQ4+H/QA0esynKbOK9gMtB41uRJ887vDE
IeO0Pv6F84MN77nLOioKst9Ync6cEYS4pxQQjavj18sDoEhbup3tYH7kJXj6oqJq
+xUKQqiDli6dOvEFWw51OAf1UouOF/iQz67JU06iJmsQRlXNGuGMygda5eF9GZuP
P3aKRRcjgFU+xFABMmjusVByjK5Ul+bu2sO0R8FydI1SBrDpkVQTVx5E5PbPt+Uo
X5urLNoQv4UhBQ17uKmH3cURJoaDisRgRDhxQHZeEewg6fY/BywRYe5Z1BFDh1r8
a6qycHmkuTkV0IC7E9Q+rvy2Z5TOb8BYCi9Q9dJa2+tXUMX6ix2JrXGDRA/hDm/c
1VnyYA1RQKRjKrzQuk1edvN9AoS/3FXRNdeJs1afWyUFDeuOyGv2FrgUFBmoSnx4
SLx1gOHwLbPBg0s3nipaLGWUxokTMjTMOhUGfSpBeY2wSuAdFlfK5lKPSmvPF8td
zIFYePdAMHaEkuNpcxDgMF+6XV9VIPuIVDTepbxSGlgijxc+F+tSs7MJwtKL9g0W
ObtO03JeFQlkqdoz/uhQ9Z9IulMrDvAZnJw83/eWfOgZc82TQsUwM/MkO0dGnqHu
72+2q/MuZds3BsC+oCwTDZGS7ltfbjCJ8cCib+SXn3kRQjmbJ4ovkrxUAil+hfLJ
gH63k5Sy6UrbxvcW1Ym8KoT5Ih4pNlhljsie/7PXlLUGTsk5tLYtHrFZrR+jblZq
30gdiVOKjx3Czzz7DInmxfXG7Zp5v2+EmB5+yMFrmpb/zDfOXysphpMzhhavjLqy
fcKEeYddQCgCKdBSvxFciBBHM0lD22JcyPAtjVXgsBD5pjIsZ5C5zirWYAm411Nr
fgrW/xSbwFD2sqU6GvPGwYvCNkI37cRVHQRBZhb7m9eCA0n1V9yBXhg9irnwq+nA
eYtzYxUsKIYS+aXX/MQuSYmkaGZpSWAeij2Lc87nqHHumWCxHxwwZIuXIGIpauQD
V7/9v1Lx3yhe7QunGfCPG98eQWuqykB/gN3CZYJywApn6uDjdtq5BgC9MzEnBO1z
vQ8oyefxRqu00+yc7UmXTW2GhEeLGNuXue4YKRgLml8Ww7V+XQ0bdyDJuPVdQGSv
Vpu9N6Yep1fh9k0wGA3VOZb5/hKjc/sETbSnl43Bi4HsS1Wy3bjVOX14ynQiG9Ea
33dscXHpy7at7eUvesUhGukv+RRL64g973Olk5mhp7je2NVLTS2WG9NIMWw9u/Dz
vkHVIC9MIiIS+2PXVrJNOCDswodBaSjJwT7XUbBZN+PDal3ux8vy64o9Hu43M08J
nM3TzSg2FNi43vvNmiPXr9M8uiYbf3wRCS4l/Bj3DJFMhU8HWxPRJ5hnBNZNeD8Z
jOMFBK2A5dwwXPzgCUyQvusLr7FWSqBvJOxp7mYf4fziwyBcRfQeOyrX5tWhrzYQ
b4sESZYB6ardiEtD7DAyfdO94OfSgW94bqR8C4NGOxVJyWvmRXhUF7UNUEwjqsA7
Zw9lYRuujVs9swIb1BePJoJR1VHkdqVoXeuuiZ5JwIJ+xPi5Z3+4K39SFKgYD/+5
4iSrMXzzDl2Wok7BvRjczGN3LcByvao5RD4jhGQVjqUXsN63GEduBUNsfPfHB30X
/p/wZmP+OjBolNUsx/WQFDZe14G8STdFxvLie/lJHpvE3ovY9KAzVmgQ67GWgBj+
rXu91EI+L+dayQ2pTQz54yWnftHFdj2Qe5rhbNYrTdSfiCM6tWvvaWCXnxpmz+5k
pRmGrKZhkZWtmj4jSZ546f08sklVATMFBvCUuY+9zmwK9P+/uJYY65BDBYqWjcIu
YQYKjJa3+SMp28d+3fk8HALXxoPbTj0RPFUKZplYRRtZfYpcPPxwGRIW8XKHmLxI
gXduq0LrQzhFJ7m2p310CtFexNh+AH4jASL70z6uvysopByPwd8727Kxnm4uYg50
yQyLgSqcoPP7ZgmKemizmTXs9d7jUZQSTZojTZNO9tSORyREtk+HQdGqdYB01BKJ
qF06tGSWtv52LSkxJBsqpaIYTfFVcJGaZ0SYoOP9k/WloDLoK4cWIAX/TBvMzxth
D/grXTvlFAnKyVa9WB7SMpsQRrt68SrL2yXoqMv8eU9jS0h5qEZCkpMzipS949M1
gxU2/adP/cEhZXOtVguVdqwdhpj4s8LKnHPgwnNb8gyGn0qWNQ916QuwEIexjPcV
DpCXq0LOS8yUeemvyMWIBUAIm/pxyMsIQuOJGj1JsqM/SOtdWcHuH9EVRs58F7WY
iH5ZFPrTurWH+cvj5XL3d/Tkfs4AiWN5JGaQGQpnGKcZaib5uuX+KszD36Ykbmvp
3Rzyia55l20cBzJC2VgWoVAoWNqIaKFWQMkHz5xFZDAw6GSQD/VLqqmpL+nw7aV+
6gjvF8ZbZDD0PGc/a4wM19YDlUyDfUYFVHRKALw0J2eTabYM1jU5fF3UH1EMjZJO
i0kJU4073QC1TXTuOfKvgytUmqGL8HC2HiKl/AacXZRP39eR0LreD2lMrtlrn1Wa
wrzQY6h/Cys9CR0PD8O4RZKStnyPb1W5i0g5/xddBWpRjbRKl6Np+Wdjyzh91zgr
aODFW1tvXrjUPUXBlD7ZGNH+dtJgdFoBuYyM0qKUdRih+v7XcC3VmH6ZTHmjHLHm
AGzhdl5bsiJyfQt2aAkqhJp90zI3p0i3MDoY76XettrRe9MQrGWHKPJ/8aHB38rI
VtC618/0wdoGD2SOjLQz1bEjHj4w0sJ2jNgHrWIIszkLv2cfNHQWMPmt8rDwIE83
LSkVwIkEeF2NM+qg+7oBzlW60n8G41XuuvSxa+D9anuk2igM2k4zIXyFWX7MbhSL
QULdY8JDYq33yXHXCloQrjfvhcRwuOjHLQ6L6zvuwxM2yGYhduFu+f9Qy8BTWsZO
BFpC4nnYgH5QMoYXNFLAQBMNftqHhtd6pYv966VGiAMZaL0DJDmaudqMBuuAhoJQ
5+MLv1b6R7rjVIoeey0nogJeZqQR3AY9XSsMSuBLDj+8jlx8Lppfiwd91V6b0HhO
gO7ipKvkC1/zqScP88ShWykM2UrAPn/7yHykd120yArA8rmUM/3RcY82PX58Gm6M
2FDvVL0Vd6usPMC8wSZgZLAY/5zYV2ExceMIyZHaA5AxMl6SMiSpVb16Oixep0Tn
xevBH54tR2CZAcfFwC7cGKNhb3OhcZ6eR42G109uyXnwXLRTULUlFrKAlbw3Tn23
+IWBJwZZC4uu1Dfgw26KC7sLd8Him0Gt29uTkS72nLpZlmXaiutTSDTLzRx6CcIu
nsCoYp1SEDroSBX6mP86kSeKwVSEdVD6FoMOaEs+BnK6iH4dTc2l7uLnJGByRSGX
mn5CyATiJ9Xr1pGkcieHtMbqkfgYlbhbY8uB4il56ZyC4a+KxV60SXj0caheJfQv
/bOa7EIItFr/XZ9aEEJymXcUSpJLs/sb/pqxY8DwSUp5bcFtE6BQwGxI16PWW8BR
ACTIXwTUKPfFQyztOnzeYEpReOEjKEtKYrq/Zy0JdmqCi1bDBAQB3JeUV1NANunf
rQuTTENgjOBynIREtQaeJ6wd4bIHUOjWQYMxPACqhaSYRsZjQWpbE1v3Z/Uujg1J
WX19PAzDW011iHChAfyoK2cY/ArODhpzd5xfTU+qO3vwo0pq0tkOhVlES3CUPO/F
KLX1/NiWL8nGwSGrP7BrV6jhPtOQc+bUWdAQiWFzZQvB3CxzBLGojAu9CeLVcYBK
xjopJ91DEdbzKv0AR98IeDCG2ALAJ5UENkKpQUnlaUtoaYAWwwqAWfbjO6e1Ic/G
vVBSTU3IhEaVOHUvO9gHJ/dFDI27CFSMtULy5644ho2x0ZbphktFEFx8PLshSWfC
k2+NRmVVxWx3NpoIo2wUNRXwqtQ6ior8ABg6GJ7wQGVOOmuZq7rE7iARhrgPwXYK
DrADCwd5mqertEbUJ8BnwlqsOJAbj1GHr3ZhAKEIVjWPkXR1cD7Fekw+oVmxK2Ug
GV3joOSyuXuhQ/Q7C4L3zM7kDZDZNc1YmXixXvztzXfFKr4VzOTx+ZGJ2OzlL5+f
BWRuaR83NxW+T7Z80w7SKIxyEO5fURrODl+k2wtk6U4Qr6wy3xfx8LfKSrLl+Ccg
gCasmp+mxUYh0pdM5DyoYA9tanUr6ePxZ/i9birF0VDi9rwDhlQIgmbWBltBcN/D
zn4L1gFqd4Ch+Uf6uglKPpG6lEdIwGroaQj2gLKyVoBnOxtmMnPvGjZ9iwvM1UQx
t46KvMi9qsl1Vri4frXVeG4Joqff5k4p+EaN5gGI6Hk0pVd/6RjEn3yiodgQl0uU
QKd91AoOKZxOpCRFfCw8jeb6FINSm2PhRCpswi+aecVOZ5YIaIDOaG8BEs4hBu4R
HuB65aOeU9nko40o3Oh046f2x62z/+8JXD77zKyoqsFUSu6lr4LKFUcsK/Pdu8hn
71ikhHc3t0SQP/4xz4uMP0t8pl+A/w+BCzjx8cdmiu5pm3VwzcroYOBSKHVSgz6G
F0YlulxwmVLmOgKYruaYq4gHt0nSlmGIUZ33It4nwzxdTyEWqXGz0yeHktqUYWoI
9dbMMx713okRDm0CxfjEv+g4HlPy3w+jWF7+AbW309C51mj0xXzICIAuE2f1ySCG
XkGthpf4plnRhn27tqzHF7yIddyU8tJRJji3j6Ot9H99fACGBknBpmCpJgsRpEiP
OTw14K7sTo8ZbsT6cNV42rVzTBfqVEtFCyG64oJAjKOX0We0UknGvLNA7A8fBIKg
nlj2i/JXaxt8WtsewE0arimpRYskp7AQNsYvijqTvv+62+h6L1Gveb4xJmUObDzd
pifxexjVzGbboZWS5gcctCQ2uRBhSvlfs5u0OX6LNSjbr8p6tcqXWeZdGqI4ak7x
Bse+Jy0Rwpi/IlwM3rjcOF9juJicwNP/J3KstvIbJ1uYHLdKQunNYAi0ZoFeL1bC
nmVyk9+0RZGpPRL317ehxJL6Lkh0M0dsb88GNKTgmeBoZGelDCiDm6nOzFb6/hfX
iNNxZ/V+UNLtbe+mQqn+TaF42P4NljOil5/ARgXM6COpU8yvFBNp9TLtdd+TtpvS
4An4bBtNFUPpFLpR0SwkTKqwAywiH6x8r6NsxV4gYLTzvzzQOaqN4C3VK8Pa9hBj
2oY77YM/jFbyXMVZfYEgHziogDZl+gaB4+zz0sm9RLY3EZumzNOixO89sXcaiivP
ZCPAwP1JbTo9lp+8eO1Jce+dTgEyux517LuclDNVaiL4+3dD4gmjPxbcpm28dqPA
Wo5zAh0DbqyktN0VLk/UFNti3ez83NQjONQ4QBRp90yIk3xGpzMnHfoJGzdEhmby
UkpOZSdY0jl+rT/2H27NnQThnt9Jju1U2lyMCmaw2r6rt7+8fXZI33XzUJiksA4Z
XjY1emOv/a7+BjUMGxCyd8zH0KBJFi1eWCzpfQ1RKvPZmDn3x9rhHhTO7PkJjxpy
eNwioD52uoLOUkOI6LbdbuyAjxjXGDjNHr6b+3cKJ5kVGwtcqBKfNDZ4ipFNS+9z
dQ0d3N69fnPJI5mfIHdTsEBOprgOYobTaIy4DT1cBSvJ4P/R/81vo9KNw7ZwCBwX
hn/6Xaxm5YJchKhgaoty6qlysalxsWxQ9XPxUYAa1dH45GSKLng6mBXZJ2f8r+rB
dVlkEXNQI4GGBIAF5pDXepH/2pp5epPZnsVypWgeP2AxzVeUH3EcAv07/+Mkhh5B
PAPh+qDd68Gtg7o1ovKmeojITX0ePe57oqz9VTwFf+qd7c3J9MQGuHdTyQSsJlqK
FbIg2w3FOeCWlAqVe9sqHbW9VEQMkyr/Cb7osaUQKjd46qK7DbPyUImuHrhbqmO4
47EKxszJpjJlxPchOMCNtsvD5qyH+ecZ+/f1tV31YqO/idyrn8xorOPVOONabMWM
wuUrGW9qKOHVv5LrmYQKnayVCVidmZ6m+QGovmNyKqgW0i6v5+khNgOpZ03/u/aX
ITW97Ra9vvExhtInIhn4YA7AWXkcsLAxDGUowGtpaKTaDVFDtfQjGqwyapTdyj4Y
XCkQ2QVwrm0JQaVxr5B+qHBJsOH663wmXhsjHgDil4WCXaFAVzmWjToKVJ9Vxz61
gDpgaJUyPd8djz70xegm3FfUeIcX5ZCArHlqGrapfs6vuj9pKWqSlOt6nHMU3yXo
O7M5Jnw0AmTqi0qB8tm1wm9T/76XyQ12FFoYuBuq6skfghcCuUYI+9i7ku8CLNXm
l+8xXgngicn63/nngzKCPYi9ZKJapOYEsN/uyC6gJLnI6uo16YrwOiI4IHIGP2em
JvOD8eqM1Wz6MOiuV07DrfKEUJFNGKVK9HBM8gDR1cvjkapZhnfx1hkIhSLskp9l
Fy9w94GZMzaZfDrl2XLce+FPWaaRPAq3gjw1+VQBrS6RRNPZ1es4qfEi1VE0OhH0
wgTgY8vhtnvfZZ0X3FnEhMl3/+2Kvm8dM18oDYSnpMXYm/0tbYCrmf4QE2RpTy9J
DxCkT+/TB37ugw2V1scRcMWTcBj/sgUwhom/oMnXNMGOAM0/JzGtjo2VWltC5GKG
1lBK4VSKW1nHG0vJicbp0mX6oBYBybjLno+MY5XsyMyrbjK/TJhJtqIrAnOd+UFZ
LN/VEgsltOega+HHwXVu116QBaTQGun3+/2lLHpLkg2cdjaYA91UWcH44fEg24dY
ScXsCYFhvgginlt7PSAaRhT3l9GsKeyVb85uC3PYhtaK9Kd39XxviHVJaSKRxH2O
KWDEO7KvDoOkXk+hgSWcmeFIK5BwJLeTFs2+fHnqS8cU7xGyl4gkQSGSwJEmmlQe
/y1fsLO+ddNNf8mdY4nJlXwxl5HyHPGBCJwMqxBAoIvqiamIfh7QukhExfeHObI0
Zta4iLk0DGsGH+uOLjxNf/K7jLhiUiZ4heZwxssyy8z0j5f0EXs0KTospnORJdVT
i4lj6Zssb96TZKYofyPAnuqMPrBpHtsBtFiP5DmFPVS7wy4KfPZUJ5iLuZYbLfYI
RY9EUgMMMPq8tRFcomT63OKAjrUNCm55mrhurRwwXYGLgTCfDeiksBTXqr+u+R6v
BlS9EjIsT7ydxv+7VCOB7K6xhNs+zOCpTixN+PsQ+XfHDHTVv9Z7VQDaXmbKsQQF
04scunQsk/hniP9cZ4yN3lLziqELgkPLj1AeiNorjYtBv5VQX9uepeVE1x/lBi5q
v7AyqzRGuqcMZ5s3nxNJR07HWqOOh2cxo4uWRyZ6/+GsbzBbNA6z2wYGcZ9E4jm2
uAWTAlIY9xfHWQE/TOmrvGhv63YDz+/UJSFvCqXIeP63C5ydMSZqHqdAqpZ/Uc6i
Z3+EN1HuN5sR8e45HfdWg8bFy4Z098Wq0kTrkDZj4H3EypuImc/Lorf1Kiu6SzW2
1NmHR+q8KFsEHf56Oa82sW3mfK/1lYrHYM51UbgFjd/izkPRBTnQgBViidQa3Z7L
VQkqgw5V13X7jWvIufxIge7q9eHPOpYL77uDjcOrOignlykttWQVCnL3ZY/5H0Rs
nMOrxUU7j7Rfo4RFJSsJpNCz1Qnz3PjGl5+0TUFowt8FiEG23r8ff8C8Ye/BqQzT
ahXWcxeQUYUtNdhaihYCI8knRi12XQL5dg6jsuHc5EhVvhYFkVwuLlGizBUffiL0
Iqntxx9ulX1fJvZCu8pbGl+7+/NmXBr+YZxbbNSYdBn/KjN8GdacmE/zowEaMWl+
YJAnA8lyw579AtAP+xoyav1rJtDKybhLc1ZDzUNTuumpTLaY8KcVTxR9v709FC6V
rtEihE7szAeFyh7AR/Ih51ontDsGEwTAut8z4eMqqVnndIsB1mKEAXvG82saI2AZ
hBwOy5jAFqo/XwmFoKmRiPnAGxyWfNDzebkz58rV4aQDCTnSBLAnBzY4UR/TljWG
Lk3lNbkD0wybOXvZm6/tYA74tC/LFeE0URNmGpMh0YgIRwcj0iqE7+cRWnVyWm4r
0DEiWfYV+nsskOjJm/o0W3dyj7QKsVaV1FnH8cY9/AIfbtZWlkApwz7QTzjBS4+7
DxVUlrGqgPpViB+gJ9G+MrOuwsMehA33+T+8zJOG12LhS3RYA259TqFL/ejGcNNC
8AlW9oh/8r2WsiJj8AffASZ9dUAqmTuCen0m17QaQJBMvRXy48ScPKlNRqUu0sLh
3R2WFUF4LK5Spiz9QYCuOkKS1rpfmX3Iey2oWI/AWTssMSN9xZobwVFhFdjOSWqK
uWkqoy1UQ2bYdA8JdPNUOwi2LztF3vnIDNuW5uCard0UeF3NkmT46YTCqCv0fiQ2
7NFKo6vaGYB2R/otxEmfs0zrj1mcKrNifZpsYY03ORx4ClTJJFhaSjxAsUP7htuf
/VESiuehwonCJr1O2WyiZmlGAdfZDYxeja3BRWc9tvUEZi6qhd0i34kd85trjB+5
PtyH6yiPD5riRW0+uXrYWrdoe8Zhvt7voy9mUVxLm4lsuC9Kej72O+9b7b7qw1Ep
FgcCZ51AEar6kP/gYf5cF0sDQkK27VutJpWwAsi1+03MPdRa+/luqvcP0pDYawM8
rO0135RzYmbOpNHu5UE3pdFbFV0C6relwg7+8V1lQPMENy3xE8LXTNAgIzbGGKpd
mYYmq1PCYLArE221eli8fMZRJq/fcNzW7B8ER2KAE05yzmS59/aj5FYRYHb0L8Sk
REbAfg/y6EaG8SmZ+jvqz3zEs3WbwdNOCZzgcmuN3JhM5S1KPuH4O8adFkcMwYaE
4yHYBM064wf3/h496qH9WdNMYRD/Ku5/muP4IlhWFt+vPg08TRuwxu6xdgjWjXQD
5InxY7UNAwe3fymFqqfk6Jh8NvzTzBn6/xf0tmCTua6dkpwW1IG94r+gg+cvqTiL
Zcv9CQoxuae9iOPfsa/UUbjFptNhrvoG2AYgJgHEcanW8QBraWx+0c4rEdfKyLm9
FhnY789+s7DG9QE9nKxfBfQOZZGCMWI807GK2Tc/HL3NIk+S5e+1W+9CVMd1JCXl
2ljMTnT+KdWZfC8fRZyi/6+IOxbKKEJLXk+CNXyJjlPEczpgbg95rQupMvV/njY7
PhMxlYFk6IiBkN5ppJK3tWTZ/B1i8e8pMKhlepP6BRztd0gcoVGvNNT3/EoAUuJj
+lhp6Gs9Ry6lGyLf3j5fDAOAlzKkBbVo8xbYpKWdBTanldzgalixH3LsO5Cv2HEg
kH81FHC62sxOr7UnpYb8Ja1cst0J0GaOHjmCJiLnYTuFmtIOpHPKyuoWhIODFp2L
c+Hm4oaLkfv7Ues2L65qvIROk9rZxOAadRL3X6g/er6nthMfc7C4cATtot3xxcVL
YA6PwR7Jojb7xY8RbhCcn0VLfrnvVLnO1iZDyUoRzO7ZhqH/YC6Ikhom5wQX4WCU
Iv9LMepBn2zQj+X6wVnhIZy8CcO8Hi3I2JNvtqGxTVeOchX88YSH5AzMfnC9Z56F
Z0D7CiyMrnrhMrjCQDfIr6aaJOrxulpxxGlZLsnX7rb2j17El0hikWXvAXXb16y9
PVW76SnOML6edDEZgvXDoafEbcBf+XWT59Wy/nUDbi2kYz6nLSN7pitxwUzF8Yso
fZh+nYqygT2tmCN3OPOVPnPOWKk3ZVpGkb44MGaWRqYJ/QudJJodwC/CXW+l9fLk
P0sBZmuhYQGbwhuwAaUeE//vN7XRmnbSNIoPx14k/murierdeNvtDmKa4acBV+qb
WqyPWutrFFz4PvX8XOJhXV0ItuwifuLLoN8xrEkVKubl1rBBjfTnbCCjej8AgTUf
QgzUoY166h7QjH7FOLdOqs/fY4Dw0rFCxoJZPTgIz0qUVUOJ3KqD1aGu64C+Mp43
nBLCnx+odwr39SJfYyO2UCvgMv+1+32oTel3uL5Vv7jWa5V3MPpgRyUIb0COVFI8
DD/io6TljQzdqqqYUt1DJe+Z8ba2QVIYqbdOCWX7yh9/OyqV/DIVKNQK1O5IU39d
9FmFXxEdZoxKHsCYsBiAnxBi0xN88uVvajSP7gqlIyRSYcBCmyiEvx+syinOzuVZ
7c0Gttwu2lpiR6pJDccW5d8F7+O0TqZdtbbk+v141ZxjbV5euFuOBYMDLE7vGbw6
7ovi4k3QtyH29mRGMWwnMYcCPV9linzDd5lK+Kj+ls1/nmEGasgRxKA+Saf6GxCb
hvsfCTz96ML4iqpx8NTK7HnHCzGzPlcArPMkbPM0J+062/NRpcoJIgI56V8YIzKF
SuEz7v3AXQeC/D1W17VgmSqSf/ErXyR3Q/py4UasdOyZZKwLgX9zts43AL+Q759M
J/6f7rNtpoAdPasqMJUSFMki711zegSvTy6J5YvCgH33L0vLg+MqYya63apavMoe
FFlzIiiikiAGoeJVacpfu6o/ANaVFOWB+++kvOe+Ejxh8p2cnbkQvSEGm63NWXgW
KN3pZwg5sh1dcwd8OKvYLH5LOIbaStwDOqw6/yf67MCE8fUzfSr5h93z8svtSfih
+7SQ5R0QISw/ETyjUwtOX0GuhlZ4Tp53CyEsvGrT9VFePjBRMFCzXQfzDR3lxK8+
O5DAPfcwbY0sl7XBkeDjH+Sqm23wdUwBDTPBYSLEMZyPiYLXB5fPxudooXF47pL7
WbHwOVnleIlKVMJaDkr3O2rdUxC1IxQPcEGsHNexvcLFvpTsBAY3gVwEWc4l9DJ5
qJBuShAQjXVEJFBSk3/sAPRS3FTNB754Rl/aKweMHC8Teber9unqkBYurGiv8rl2
cIAUOsBmbz/0N1PJ9sgV/bC5aqOfMaBl/hefyr5yTk4niNYRr7+1lVsROREmgCUW
1puHN0r8IIE8P9NZvsTBTWobyzdMfFWlGqKF4SkKJu+6C5UaI5l0Tloza7xBfrRs
D8iEfPqcucln7tlXAPSQ1xHQaV/n8lyiKzNUMsBLUKPEQUvGgBaquAlBhchTYv39
A0Sg3FzHSTaWOmw7XdqvnmXCnDtlOXlg9qOgWUJWgqwzYktGpSoP49O2fXM/8jJ4
Ku5mKDSuVZPqUCXX5id14tkXCdfFjP/RP/7+fkzYNzWflJR0nLFwGed0OoPYD0Df
Rf9Ez9FH6B6asEFmIykuGSzgqzmWlzHDXzdnRQ2B/patidyZLocMKkvM+PX2aW2O
QmSW9uBhWcrJpILG09up/eXYQpSJPd/xRPCRwyiSlyAjy+NCqEsRe7YnjEpizLKb
MHRaMUXtb2orusL+f9xeYmZpoww7g13LrsLPtPaWW/MJ2IkZD/XycQ3HtyTKMSoT
fITIpq0W75YR5q3dVP1lY6wop5N3lmYX1kmjkE9Jp7NovcABr8IP8YejEPadoZWW
blXMWXC+HbgehLOisrSssTP4EOYXVvOXB0b6e9QefBMykySfBbBVW5bensW20SGh
JsY9lkFfCmWZQrI5BIJKYBtxqCfsAWkYBpVujBBvLkYdH8PwxuwsBiQwRkSvjVdC
mG3S4qhEupKAy1kPzA6FOrELoRMwp04pzXHqzOatxwkn5X+UXB/BomxmUZ3YCooU
XY1E+72kCh7QJ6PVCnJLxnNTbHCGcMsH/yb4TTQgpinWEE/F3j3klCgaXdBYnw6t
cUGOASJAkuLB3u+5ofRarzOBJwU03Fr/FFi1knssJHI0CR8jq1wI6Zit44/8gkbl
DvkFfqYBqX60X2HcIY6fYLTJ1BdpYSkZXaHXNair60YOsLOJfpzXFm1iTwtPQWS6
b/uAJOCyx5tOgHT0qcE/bkoylH0MRW9cohNMW3QErm6F1Ew8MiQpLTxBwG36VoS3
vy2X++AjLlh8tzaiicU3/ITokImiLw/plKulaMdXCc7PeN5PIi0tW/etwqWwcI+Q
caLsIDZ1VqvajceHG/Mni6pwr4KoEnGRSRdmstmNV5aPguBRK2vt5H96BIHfUJWj
JyChEfa3B9bdfc5D14kZTJcH3SZQVmMClh2GtdkDvBoY3BkmixJM19i+Z4iZ7EbX
o9FbTLEBr8GAp9UjxulhStWOv4JuVQij14HSUYBmr+zP4W6Nd2MuCFgRQU61ef+5
R7nkIduCyM0NELJQtBEjdQXoWPIk6123353qy6qOulSVgB87Zz1qlwAZ5THSTF2J
vWlPyviIMxTeiEfHz8cpcokPF/FDu/yZIGkIyWTo03pq83SnRheRTJbXtCRQamfm
oG4EmsQvKZHnGRS5dUKZaeTGOf/aEQFpNzzSG1759AMOOILFzOVXFg2eU8X+RfVF
a39sXiz9F11D2tGdUGeEI5wOUcKNhElkpsxbwupEC7pDIKAvEBuMr0fWyglQPr0s
lKxqryrnM3hA6W0vQ1zSpJkn/0ErdFV+iPCAwj7rWlTvt+gcR1GbYvAF/ByukhxC
sk2pVgEYkO4nzkqFTNk6oHC255UuqkZK6s2oVswSq1IPz4UjvKSZRUEp7cW91rcJ
12v0mMo955tnypCPrVu83CoOuFxG9L7YsBmEgvvmYTYS8cYZ6eS5iDl5LE0rGgBY
D7imFNCD4GY/tQG1P7ZhclWF1ecqIreOLbCaW3HfN3WqwXyDGhxbvS+Fr5Cy30wz
UfxCXBhaCHHtcg2VQsnIz5UT4kEVu/Mtf/8VDYR1KMF8elfMSm0X1/LbDzRsp+ey
ckrAw1KW3COjNrn3OihZ+LmNhsDfhroLhaN5rRdkl4J7wTd+wfWxXrIuYBHh9v/s
dMqGOIzqCGkcYSzvIhMr5I0fJI1ORdKcnYkflSUDBknVpTT5RDNl7Vxe/EGZo2y8
mIMBosJcus9Mxvy7NtlEab7yq/dTfPKjdncLeExl7Wd+R49Gage4Qc90D/0dJRmW
dgHKa77J7wBapczwrqvtbF0FuKQ/CJxSHambzSU/2q/mnJaIVDtGujlv/kG9Whgo
47AWmPzA8utFRrfsV8E8Exl6b4jCcFEL/oVQgUpVvJxL6pNTcObx+NSJ5cxNZuT0
wEMbEBcENxSEBbnVNvkdP8v53jfxDoh6CP9Ni+YG/qFykJafZBsGTEEu4fRG43Zd
zlqIuviVAdo98lw0m2zMEXHAwT5YkBjQSkyJlf30s5nqM42qjR0gNyUBVdjsyvjA
o+u6rbQEQmuMWle9/GzfL99DwXPdSoIG/vNmmN7WHrpe5+2knczLxAYda969QsMa
wnT6nCnVOZoUaJc+pYBotq0WBPEJCX9wCOu1W6pTxkY6q1uswsbOeU6LBO1yMkzK
ca2/AQXBU1zSl+DzpLlAuAi79TpO7Vl4qZ5YRCnHJAeUF4IfLYg4tI++Z85urOoY
zpzyMTy+dooTbOldz/GvDCJu+SYMrioHbaB+XIFsunkwFoVtdwT4EA3oMWQTQsbD
aYOwuZL4lqXmLzLlKF+3ZbPExJ8t9JnTmevICUkYk1+eflNtUzIb5NK2CSNc2HVP
pThOMND8UU1WAJnpGjtk/35RW3pm88Sas8HjrHVo3DaMM9G56mD5KUQWcsuYa/0k
fAO0Z0mrMg/sEzhkhBdxf7xsk+19wJcSGBS7o33L0c3B9pptVphpvp4QiWEMEkho
V39KzEtYKYPCLTZ3wMb7GMcTmFSCYKP9GBCcGKAKBjE1UTVJB1JKVmbD9rmTsEiu
9LeVtEUE90qruN+wncTc4VAdo7G+dTcJj53vndUeIO0QI8y0rHrQH6OOEsw8UXz8
vu07XvGunMIImx9XrtqCmhh1OkDVKyZAWwyhFgmRZjwzrsk5MZB2dS2YT5zsQ5Pa
KD72gw4b4V4Y2e/wAE9upGMExqkE1G2uKqv0LDA9DkhoOmTG/xXv43lQ75qpk77I
HNehMSLeX6C9tBNWHYXmaMhvH2hs/QdDbxGT2UddrKHbaTQivMz8rVIQKXHsYI1l
ySHt0qB4zOlKxBo3sn8yWe0xbIlVWz6f3XhPvwanMPt1VDu6PPKFMUowANt65G89
ZI9n9PJfOsLDZ9dG8CbQWbtDE76UbmFzpydI13B5atbuUSeqoq4YQybBQZ+F2TPu
vtkiydHk42PefWAUpAoFaD+7nKb+jMIMe1QBa6oLJW4ciFVfeH/GAfnsCUeC+GpR
MQVxIKbI6Jyd5qTFM9KdVkIVh57kssELCzmEckhJX+K8/pPs4SmICB43PJ+eXpjS
zEOGGOyA6ozRKpUP7hF1eKKDfAbkSy3FbZX9ug1o8QO2vamHCj48miQ1/F6KJO+j
ayM5zUkckx5XZ3JkUjzENzhpnSLCInxXRsOjTuc+dh/4hG/E5ciLoXiDvZz2aIQ6
3v3hBBSWt42O/e4e6ihvb6UTdUO1v2rco6kLGRXO49fQOX7D1sBMi+U1QnApcQdi
/wRh3XwDAYzfZtNw0yoJpOusS0YC/xjryDL1cUMzPrOncoXTc+PtteXUTPzRW6E0
YtiCUYavMTs5pDxrdK7VRCOfNWCWkQ1MAkdipVCvr+zuhfHIOkWOU4LnHNUypGIM
1g3e4VPKhjpRo7RyvmO7C0x7pBmjYvNqVAH5aqj5lohh1MQS7WVQLTVSvoZhYmWC
Se+sKsEtwNN4SSEc5tJY5Q3SmtBEPq+FONyJEUOEnva6BI3e51m4MlxHILxLVUWQ
UHnbW58s4n+bByYz06l88M3qh0Tf5JO5jk13bDUn0TNJiay0anzdsN9tn0eMzn2L
uzBKbUkiVhUOZMCAfwqZMTYs91KlKapi4Lgklx4ZQlYll9oA04emoDVA+FQXjtqi
ekvC2zXc0H0O56B6+BjpKmWYab1JKhMguTh1ojpZ4cJTw/XJ0h85WK3bsMoysbYo
62uMJ4lLEqMtwQQ8XJsrqptnHrdWYMTqMwWm0cEtV0UofKth3ZvRgtFx35F1R31l
M7mM3WANXEihVKbWL/vNI7U8tbTguz7z29iQNWgdzDIQhm9tVphIpqYfCo3FtRBz
veu7wWDqU8P040QHX3nZLy9Y6DH0kHAJqt6zjqGO9DLiBmFk+TX94UekSqLTTCPE
TN5XdIdN2BZX5V1PVNJviI3gBFYIL2rmgh3eMpczQIlqL/26hhhQ8bxec5wCUCqq
C4e6mYUYIAYV1Od6XmHK0xtgtDop//9sBI3u/49MVtWfQlIaJ5GX40ou6nQshfpc
Zwdhg5dCjfWIe0rYA2KOnZusH8A8/DrXgiilbW03pyWnb0HdBWmML9t8tenUM8uV
G5MaNWTe77n9kGZ1rvWE2PPJofKjdTXw/3PNMKtKxU0EukN+04fd55kIaMe1ovAK
1+Urw2VNjnDIjvl+psh5TPdX+jvwuw0/4ka8NRio0UCufqZ5Amu06lcPDPlEcuSY
2eM7uLjM8TpgUAy7F5a/vq4ndfSh6q542m0VCWNn8oj4aIpb3VPcmJ4tZANjLuZH
hkduP0I5HWb/2fI9H5UEjNbQypCHQV3PAOYTO2N+3YLeL7R8ucSGJqBhMyZw1BXX
AoOOBqEgFeuGoyicUMwhnC842zg5887xAXxHJTM6N3+h0CNalQ3Gx69vrc9IWqWK
BW6wuf6XykCbf0EgNTCmhXo5WB52R9LBAdVs+KiaQPcAkfggnK5MEq61cF3I8Aud
Xk28ZNd9KGByCZ0/s2c9vD9iJEhBPLJTD5BhCX/jMS3eZVcw+TlhCCy3zP16043E
cnyOQEch8p3NcQ2P7Fsx4uOclCUi+5lH/QCc38ya+HEiqGiojA/U8t7KPp+VepWn
rvnarldf0kDPtXmzw8ifvZkATAgQk9NxAt38ADFAkKfU3wWnKf5DtfnSgBQ6CCP0
pfsW8zZaOhIml9zXuEYrzgZ9l12DC12SwxVFqagpsd7w3Rj0FzB6RTKXQrK91hvZ
ax8Mt7yl7NOEMktiLUrefHg2wpeM0iu2cKX1vuQjNYhDYnWuTD14UFxuEOI4lMqG
MBThNBB9qklDDQx5WNOjzobzyMZ0n8OUZoHyQcizq8wZZWxKLFP8zPkuEhpaucC5
K7j3HUntAJWESAo8Nrv2Eby3iJdotJM32Mkn+Dk5lAD2Pwcxix12qPtBr6h3ftlE
OXmOUN4uq88tH+JZjjgXmhnRRw60y+IsLMLFHGQkLv1AZVlIbEq5dYNFfvRhU/ii
71YRZ9AKrRhXvqlwGi534n62oPMLVAX8WDmJldkw8KmdtESTNx0JytKKJ2nKbuhP
3x3nwcnCMyOHXUI90hz+FKN+Qv+En1Krk6DVe9sTIYIzsvbjhj5VgVqS2/etNW0T
/gbt47m8XOQ0VQRxItbvo13ijcIyd1QmgM2mo5WbN7S+aq1UgrZvfVTv6aPJPjDE
g8Zm4OOo6Zq728uixwSFz3FKiIsm/FnoI0Ny18MbnNrdTaHhPM11q0VvtwNo1wAl
4RdIj1eVztIr88T8V5ezgCIF+1dyWlrJPRCbqoSrL3bT8U5lcA2Qi9BhkfEXY8DM
+dafDyVO1SK8at8SU7Tvnl4ORLexEw3GVsVCZHbKqBTISTZODZW/vbwrG8KHPJK7
MH1dZj8PsR825IXlD2O77au0aE/kLahb/fWB2tKnEKZnVAR06a2lJ/qYIkEiv7zK
XHlGcyORbATh39Ld6lIEsEMtXcsnSFpLd7/WXhAEkFgEulfIQhAVZoFPtT2qqOej
5K8R1USHV8lZZZLaCwt9vknEgnmOAEdMfiU9Kj55JtJ2VRhe3Hn/rPgzXT/wuP3S
70ztMJ6DV4GvrzDHieTm0HzuPKdyvCLiB9vPRQIde/vueDlu0+WzpG6npFI57Eyf
ckLQzPM8EseK51epX/IVuIwml1+AdzSCPvNyGXkIYo+YZ18pR6patYx0IrE6v2MC
YlkeY+7gv0zSouD4MKLnYuhphgKeHyXf7WusPAeRjqFPL7uAsV3CB/gYvtHjubsF
tiqAM+S6fWCrmyv7wiccKP6EXUVL/jZtH48mEQRpWDRMbORwqXZPltgFh/1zWGhr
UlgegmUQNdcFYYa6qPTViry6f6XXt5X17JmuHkVNW1/XbzLWihhWbxssOglO26eh
THGZmSToXKfjX5OHu5uzbkl8tmjjaskpjIccWeMLol2cs14z461b3/xVF8Q0WmC/
O4dSAeL2TV1AFdcDGOTZl0wXUD5TYAPQuT+20cSK2+i4qRf7hdrxqaCAeElpKyko
f+jUH6KIgsyPLqL9NhpbGOzXzHXDBBXh1CuBUKMVsT5/Wb/OWewIEHzn5TZV5KpT
gLuZIOQ0YwIyLQ3OsVTdYAOCTMVjdFjYdeYltc/+FDj4ZCsvH9Z72m/Qplo5EPRL
zW64zbT40OYoUrd6K/OGXkTM3eL5YKsxl7V2pwT8CJsK/hYsbWYvvzV6aMPT90Aq
63YfGge7WXipLJx9kkk8tH+gB0/yLN9lE0IiQvihBP6+//ruKBIC45Q78MokwI5M
2Gtf4elFiHPfEYw1ZK9Zjhn13BBK3Usm5GsEf9tVYP0JOY+NBL3iyvLkK0xz9YgP
yn1CNT8Ug0SJKvKy+A98Iicx41sjV3h/OYFmMvB5WnARBosTPuhMkduIZ9xmvDhQ
93zgHScoidOTFbfhv76lYIUS1PxWm5S8kuuP2Ml85AGulq3SJqwAAksqpsZq+vah
EjI3j+Gr2dPEBhPmMi+Z+xIJEHJ7NajJmAMZPSmjcVdRW9sdvOekfymd91kOtoZn
v9d+Tu4ksyvyuCdjPSryDVdyv1OJ3DIcIUlDoYzoHsUv7swMY0qgdtJzBAoMNwoj
PxQMwK+G519nxHOYIkb/SEEqlin2y+F7yqlzx/l0CVN9c0H5qWoiYGUtT3stiUAb
WkazHu2aE/YvZtrDnPySzmEHiO0SHvGs+HBLkwQ7AShVTQTzKtpCIQVsZWow8CH7
8NfX1Ix+ZjOGrBIma1/eo9UvyZafW9PLTbWY/30AXe4/ilA61p9Ax97MZ6r71HqW
anLZWMKJ38gXyh+VTnJAAklizp3pwgkC3esJWkaliqWsST0jzOcorPoiua835nbL
jnZ2W5FS7Fgo6wbBzJLSTHWBNRFVVic0VAQeKnoe1lXnJN/7n3OTEge+MXH2dgIP
4xB73L7hUeRiztfbPGGYi9/O3Ano+7JQaB+gKIfzG55RL81P5jOMZ9zVUzVv28tw
YdNwy0D1iGcJ1sMg3xbFqnZShph8jau3kXTG/ZYVVh4M4K9dh2PIvPGAkP2LfpMZ
V7Pe+0sEHHrM93IgupjRvfogk4vieISu3ZvoUyCjd2MBRibuk/R3GGK+9WM22u5S
acKvFddbRRvKTikCUnO7ryzGfsn0im7TMRwh5OTMwIsbGDclkGHz96z8jTjVAAW1
kxT1F/SulQ+YdQOJ9l7hG6DLxlHU6GGzbgTPEqyP0FICsqUWGnodFtTszWx6W8Do
bDpOxxexq2pZc8G/erGD1JvRT0iyNa+qsNEEA5PcMJXNfedDtj3c0qBiwktoz5gP
oX+4Jkkf2zflla9t4rjzkQm+1NWIjyK2MVWlLbK3HLHaHI82M74RTHnUH8KWnSyO
YE0GTkrqmfGuGnLk2NNLMjr6yYvF/152qyhhcVwtDtzfUFVtacMeTwcfgo+xZxpk
HnrRxVzqEXrxImsUTXJHThkbqp8QwOaYP/Af63x9jsVFu3GP/+IF8Bj0lpD1DR7N
0DqRJ9380W2ZsE0M/REQd32IjzHH8KBtI7Q/EKjXphAMCWfyXKCWYLmfsyGjgDAI
T098+OXcTY+SsUtySQYIijqft0hGn1koOKCQlsp9Ho0Lijcc58zWgoTlVdqZTMEt
L7D91oRGpxfbSJd+EFquDcTbpwo5kVK6q6GJrvlY43CfHUFkufFpP0o2pCjwP9rN
7qh1LJtmA1FXcjGDayto+ZKYa4i8i2xVjx+LcHG+35uWAweGC+PcnQqCsm11vpZY
8S20MBYpRERfGpOPlVpTqJkpUMOHW12N6PcqtOBRiTxqJ5tBZ6l9nEqJlITha0ph
56Ahnxn2LErt7qFtFSfSnh14HDlBVUHF2L66lBifCyG8PZV8dC5sXRp9mdrSKxmY
ysZ25jpPjxKfHBWH/InMU82KAL4tWiU/hEy4SZRqOUmjgJVrcJmrJiXdfXTQp2C4
S2NsJVihMnPLSveBYpzqVHrQAIYBKv23Z438I6VDtcQZtYfEnniX5omUqUuKLQWW
6JFnTk0ESMMKTjhTVbPUt3wq17LakNDy+0V0oBr67f6ULRu4C45Mypbqg8OAymgG
tWq44HkUt0UhNHFUtQ5AiOtTtWJeSJInSsLaN8TMV6i+lleZcdMh41xkKfWaHeRr
VXRRnEwZTUY1oMTdRN/BSr7PpQKF53FWYyRXZ6bzCVzgsxuXyiLTKlBLRovEsyU1
y3zcUF0AkIvs3/Z1KAUufHLh7cXzcRSZbiF1sHAEzHSWgXg0aOsrLMV9IcoIGFmi
NQlR1Uf9ERdECfayjID1hoMvgk4lru1Er9ydTiphnno350fjwt+BAKdpankpLnP8
J+ZSww4NODnt5fn7eD7WQcYmEebtpbDkW5ZjI9yfPf/0qiNS+bFMBJyoIXocmpr/
fURNhzrjCC0z+f535uparjR5+/T212gw7xpLmZh6+qC3GLPYfQfD7wKpBXKBQIhx
3wb/zB6JswjZp9sTjHlZEM33tmodPdEgZGhHT/r756Sg24RIGb+rHubTugftRJu+
byejS+WSOYY2i9l/U5gWgX14pQ1EpLZBSLmR0M31ZFD4hQILeT7pSY/1tqRjmUTs
ajEBkRj4MusKgPEZI8WMCtTQcaOn+8zU4yPtTvWBt+Q1RzF7eN+I7Y3hCu5k1PoI
/HxBri/Un0DCuHnFOLYmvgHUT+jAk9fUpzZMX0PZ/6A89JuvVuOhYUQqUKJk2mGS
/+J+SXIIb68v8zOq0kIn+vrheUHCFFSownWRBlAftboGlr4reI5RxhxCFQIHLSgZ
yMwGK3toQy5o9koWDNYT/M99+8CCjg3vtpX3pUNIY9J5fktv5bfztESJoVxUSmce
AR4B5vlcK+A4q9fe2NakveWmqv9cZK5uHjaBLo7+VX08wBwBy0vd3xCwLSi3CTOP
ufuO2YR5b5yrs0YkUoHW+40BQXzrRlnGhUDdyHg1ZJfD/EX25AXMyZt9EUGa8rSQ
35750Zg2E1Q/XYlNE12VieahrzWG+Y7KG0H2Q1VfaL47tJhg3XN/DnD/QjWvUgAJ
Rj3Web5dQVET/wcUguDzeUWSZxp8gav7/p+KnAYpo1OW4NI4GgjId8UP2dMZMZyE
DkYE+VYkF0EtXbc+BJI1LcOJm03xr9FaX8WNJup6eWNdd/wwPV0Fmgh0SlUtVu6i
8kqnwhhcfHI1O4hYYBSd//6X5SeK2RKn8r8B6wbWi8NvkvdRKKgTpkjmp1GVumHw
e1dsu8IXv63y0ZyLnW6wO2MTRvdZN2bfOpIdSNK1Hp0kR/ZxPsGff6FayhoLKhuZ
bFFmrrAe7d8kPJYBe/H6pLIXIgb9z+pdagyGh2MmgCPMRbcTH5PSk6SS5gi6ldMp
xuj5N0kAjvYehgXGP4uAi8muI+DqM2KtOde7fS4zOg0JvDRqcEKm17ZqhpVplDDV
CrBuQP329gccvNGJH070R5kSR03WgtgYBYIp1eYm6Th6QQJuTt/zECwW5tuSop6v
Hnk5jqoD6pXx8yWgJpV8+dKGES2xO5lY7Y3kJV1cX1bqNVPukGfT6c5Ldujews1T
rMWGmKBWpTdu6q+JiXlzbCzh5a4wXZ+SPX9IDAxO8z7lBlbvKxg1/JNrT39r3DHK
Xarn+Bi6Qy6TE1T8wAPiInMMzNRC/9txpcWmtveFdJOWlb03NpwkNDcoVWhjbb3d
iQ+3tddqBmHBxw3FQdT7k/QWvEEUBQwXlA75x9y+yiO0y+QRlfprxQvlfNk3hvJP
pqwXDoqL/2Xgo+Mg7r1rZvIIHWUDNUWRDYCX4l+LJIAnBoRXfeoNX5c8IS2vg61/
XthAZaz48M7l7iHV1qjw0GyD9jHAcyR0usSe6Svr/DGsVBveNT9kGKvnSZjJvPxc
Qsf8QjtJiL0OFmOuefIYgYs3h40hDZYsOH5Vf8xwUF/NmJrxFklkHh8Yd49eQE2w
GoERb63rcLW+WkZiOQXccjYZJutgkjOeVcuqpcODMrg2Z1PR5yWmvAqh2A4AeDlg
v/8t0JjYT7OGFmiK2cUfpvt2+U9WvdsiU6yBiETWwlOXb7LRbyfQiM5HqFf3Eo08
DBZyghiArZuWUTLL6yYHRf+7GwoIQ00skWOgGMj9HPcQFAKZgn04izgNM0YI/x0p
TXLcvODEXalSU69PAzofaYcFYHlBPj24zWPsXdtQuy/5Z7e0s39oQGAL0V6Y4gbP
EsMcF+8+QPuP5/wLLqowk60qL6meiohlfG92EKe95FTZel7P3/2q7aBE1fTLzEbm
xPuXA2v+GvNV/LUJatqBUrciypShY55J0BCg5c9uvBFuZ86cKBMPpBrz7Kp7mRBL
AaKuV0eorB3LMyBEA+4Uy8xJZXHFENwLoq2K3iSVKUY7MdSJwY2sq84IirkyI0uA
/+l/++2U/k9h5W5rD/5sqWwSBXGcsGVUUXqJxCWMFPr6uLPttAyth/qxEii1rbj4
h1Mk1vG0xc/Cj1d8zd10xJgYVujN+Yv/koomV+8OPwuoV1WnqNsnQXPnBWUK20bU
lV4miaPwg3xqLbq6jid3f4aJiWkpe/PiC7eGISjvWRD5Oct+Vja7diRivE2Ask1q
Elkm0i97/UOLqDPf2w/cVzc+jkuY5JRHJlAeTQoxuAuZGEA3knEjaHMEtFUGSZHj
0Fy8oeCjwS9X0W1qLxtTJoECzUZ/y6o3zr9nbHFTmMMQbtJTOfConoKoARjLft0v
Uh/gEFytoc7cEXB88pzjlC4kTEqfIGjGw6bYRIWwrAWALuRUjnMo8BauKHnctRFI
WJEi0Ovuh5FZL86AoBy7MB5Gm66x7E6KDID3nv4kuOxOvaQYybPobL5i7375msoh
LcQ3PMzfUCdUrySl8HUm7i6+Qgiepv6V5OMAo16hL6gyh94rgi0NEIsu08rswi9V
yQW9bk6TCv2NP7nYECIBnRIMJLQ45h7Vc/B4cwoMOC8WXumKKIO+Amfz47/4S3jL
xYJvnuYvWbS+vbYAtrDetZ3py2J31gYNoXhXzuuja1uGGfqfBc24Z8sjFRYhk9cK
eXdJDea9BtavxrzfSMPNLHDtIXZ5FF4a4eSiYuEL3+VhiTIpWqWAsl4px9OvNugX
mTUKiRT/dJCSwbg9ukVGace3mWykpJ1b1TlI7arseHUbAuc9S+4jnZWzOqRA3gri
bhguKDN+LG6sOtFXK/mq7PbYE0EYO1Oxag4XYZOYhRH1Zsa4GbQd/G6Mw5IxXbr+
6zshHuKbl59FdIivewaoY596JG0GAgVwdVbNzMSrjBjp6WaXGJRQKaUo+VQK+0cS
GR+A8Y5Evb0CzsGlhiif5ifcKkq0wXAEPIYyjWjlu1BB7ZyuYGpTWz4VL0Xr/Wu/
GeU77k8dqSRkaEv9LOWqx4OcOpSytGymVsRYVeXpeUkGX43uCTVNkV62YQ7mQ3QE
vike6m1Ljmgw9a8hNfN7mO8CS7L+slFajM61DTwpOvRMZEwn+z2ETi8HwodzQMVG
D4x6F/dHU64evd2bhOscFHxNfquemlZ5KZhVLnuVFV4NWq0U1C41hUN1pX4If7rK
ZZSwyoOg5r7iGAv1vs2uiJhsY6fSNHLcMNnvvI9HoMSgXRsot9XRwHobsz6qcGYX
bzK0V5vPuXzzHNshyzkIRr2AM9c0nVGct8PVE9P3AHellBQcHFk1h6z0lURumBYH
z3PuBqEn6AoUkp6E+kGxj/QyNLe8InbKZUSE3pIZySYZEixSUS9FY5t10mSiI20k
pgjDyis/k5IAHCJDX5mnEoKKxmEu2/zDnlw7zdOgznxQAHdk0xRVid9GAc3tA5bu
goHbbGe35uWItQg4JhXEbJ/p0S0OKlKBcE+xIlpgqI/836IkQUpH52GpfzrNhwJG
WLlKPhcWORS0YJVMmXLkPOEVwCQHycGccWCC0Y7tJW/2Zzkb4O0trRVz178sttfO
cqGftQag/rLZ10vGNMq/uZwG7LBjDUqZaOqkAlM9rb4kP0gLFdYKZI/g2knxolsq
eDKb7hYvFZZL/VQk6C69nYX5dvEUWjPUtyIyMh8FyF9dejpKGH5TbGX8IYP5OFQW
esuIJV9F+EQeZnpZP1Re5Ui8gijRxzFJeKRf8isSCyQNEc2PyeX3grOwIFvLsdRw
EBTwJU9potxZuSLMMVAWDb4tOk964NYo95vC2/pt1zhVcWZT/hL012h40zqw5PNX
Xm6DjAonH+AL0UNplT/idX0bj0hvmYIVoBExnHxqS2LhXgcqlxAlMTr2Bwe8TZg4
+4BZIRNbMJSrfKGO+zf0Mvlr2wYmO/c45X2zyxteqoVXRaXYHXsGsil61cZUabkX
0chgGiW6W4NNXMblvy06uGRVyOh0itcJs59m2GIfNVJIf4cyhciuMpC0G02SxF1l
89ku+Y8xJ4la/Mur/FZeoVcQKnAZp8QCIHyBd5JnFNxnNKjcR4xWWZpSovJVuYz0
j3EMpxiKGVp3kiaJPUHesP/L964DCytZvnXob38fVQXtvvQlULdICxjC0REbWoUc
79gOFGAyCKxdE00S4EfwbLo9E2EBAK/DvcjRjk/aFUssgbLt3hhLTe02DOsFktqP
aUOOkiIoIh/KM/k7WghYcSdlLe5b1Su9L7AFfSd3H3Czvm6rxZUGG+8+UxGck2hx
Dfgu+7oXCTRD3pjk1K//OcOIe3FqZmCD2Rw863eyzDZuLeHMwXqWQfg2lbWx3tyx
r89gxxYu5ozrxCbk/oscVTZhSPP9PoZ8TJHXjclW/Iv7k8ZDvJZrKEC85mvD5HNt
g4Vl0bYsVzBJaQs4YgLRenw1vHA9Na+wzOSomxmq7y6ifPLwrOrSE4XEfaKH9Iwg
QK6DYi73+MAlvTuG+ZSKgoGnMoCpdal/otPD5HC1wfUG90Y3P0G0DvJfJ3ilsLZk
iEBAsutzSqsb3Pw5F6PzpKZ+30gSNY8uuf1rKAXQKg8VLwquX/GIso3sZwX85Go+
UXOQGnep/gJWg4fkJSWNa7jta9agxl6OfiA7ACgcg0NpSz24xOepzC9kdjTyriWy
KGakSPpnj9qFEhUXD2aIqIFRS/uP31NwXTDVmkiNFejpu1AsnPDcStL4bSwdU7uZ
82i5qr8vwVkNwJhrjy3yPF3ve4fL4Ccf7lGrqdfAzu5UknnysUJZ/xdrdy84oRTn
jY8n73HxYxujERkUMgruTFD58qOm7XSc3t0JpKRuUVZDPoQqvs5MJlifz9lGpNY6
nVlwFpN2iXKJP5Bzo82lBdFezxwgQU7Wv0x8moqZkep/8/8ODL2YqHCyJSGPrCwl
aIb5hFLhoOcuTmBsk5X/ZqB1goeNH1R6tclWglnEBvLjU82qB8Cb8HcSExAvVSze
yVXUccMAn+I3WuYuLlG5GhEiM3rQINIg+Ej9G27mIcZ30Sd7RF0zk36UZSflOnO8
CG1sE5hJg2vIgUMqqk2bx7H3ucEaoMRUgpmDMMOIRi4YY5QBUxYKMWjtZd90Czbp
d9Vx1ClnO8rKwKhiWXaYu+cM9vSDPbLMTY4EGQNUM9sofKZ3IO9/4wAt/ukz+Zxm
LTBSwe/lhaY01rhtoLQ1cOXOVUYT0K+KIMMwTomirAwCFBaff0lu7RVBl8t0fDlJ
rv1UZNqVyb2JVq3962O4Os+jjYPxe9ZWZqo/prNr4b5n9tjmyq4ppSK1sRSkrNOR
ZDQybxqprNM+dZGxFE8N4w/cquoJ6vpUxqTmaAFTQ3CN2ZXLyX28arYaNEnAlRhw
ln/Z9h4j1PUHJ5hv8m8EJS38M+ntk3B1ImTmN7ie2Jy20IEJiuiEmFxhVXzh3Dss
WuoLgvopzN9WRQpp9RIiBYti2T4NPrzdQATYZxzXjQclOodWSWPhi+D/f+D+zek3
+vDHaR52BYUFRsfzHz0U6jk482nUvm3GMgc8d7z6PiZ9NVYJzN18X3N6t9wQRL3E
sws92ZIF0fPM+gxUAZ3xeez3TzHttCo0Fif2ZVVuFv8RdPNW+IvDanhLFvwTZoig
N+dGx8htbTp3W9p3HmPDVdE9QVUEGY8QrI15gE63EPU1tSnU5kFH9LUEVUT4DkuM
Ozx/HyV0+EjrbpdyOxz5l390uy0vFFExUB2v9yn/XSkc2tuhcjQVhoMuOwEfFK++
v4jnc+qOJmScVNF6xX/9mDIHHzRxMpjN4NWTmLyJwuhqL+6XDfUCkgem07h2d1Kq
hljv+IDihdRVIlHqvkQYxwF6AIBZIeSZ2yaLCNQ5CokBY3il1K8cyMk49AKBL2xC
CFy4PuPwMhpb/242FPxSjXZ98sFdAKwNtCxftYVF7EzkuAkAQRs4q9w29EApn5Cx
053f1QYyDUsRF9w68yS9rzTie+irc99ML4Pk0ZFCz7ZtPt1/qO6Nsx9CpdBBdSgf
AQXf8Egdr2VK2bjC7Vzc4gWG51yvHcxB7ljSTD5HjeYDtCZmz8c4JWD9szzFnWs1
R5yeUvKT1iWMl34VwUDmzy262S4bIMqwRMP43YGmRtnft1att/oDhT+qOkQkW/SB
zp4xPdvi45mYpQ9xV1uVf1pzyzj+/CbIFf+GNumYoLE6BrjJacyKaTR3MV4om00/
+N52ye001METNmHdZkyA/Rf7ckgkvopTNq8aG3bTfc1X/Z/mTiwiNk9FmWOu2e3A
j+uA2udv8tu1GqG9KtZjaJENVPg4tb1/UUrThljlxPmWz2YPwLWQ0EuUFEqh1t/C
xYnLSshzgoMuPxrBrgYjP2CC+X/wCFt126e5CGRkkoAfkRcM0nvhwKisT1wru8Rk
OPanB669uoNjBdYiRcQR3bfzeJFGQiqtiz8CnufBLBR7dHkq4IvwRUK5YqFNuh2w
1upg5ExHIddsm6ITqQ/G9hJCQS2pGJ5XiAlpNigDMGBtkCXihx9tmuCaD65+bt2t
1RpSTnMTT/4rU4S3nA0bLipNhpTqfHXkYsUJc4KMsSTbm67L36fNN4SGM+wJsId8
aXzCmPIRbiSeEv2/11AOfipcnCSxzN9nx8yfZy+gepu1y4rAhzBii2Zyx36hG9af
ZZvi/2c+Z5PapUAighwyOIGFvHhqEqPSjuvfjUNguX/8TzUzGv/N8M5CQQ7P9+UU
QpE43cLDGXDYqPq3w4k7mJEoSPn/U8GFUcURDD4HHzgJgCM/bjrYXFtnGVcXhkGt
C4nWnDfp7Ca2HPeo/DVIOYVJd+B7RC1V9U5ew4RDEvP+JalhcjDmvFmmD8RaUTNs
zeQeUg7+yHOAbztZ4yo6lHYcon4cdJ0lvp5AYAGoLM1VAZqkJvpQC1OBuToAx3ig
tYpt1jvyZYLbSc1trR/uxtkEZSx+IOPvKGinhg6yDyKxyZypK34lRpCOE7nQbSRE
BpYeOtNce55ihhASYeJTR5kVX31kvP/18ulL0luANnhKOcNhPglZo2wigmKx9M3J
rO+Fu2XDAEmKtdPxSZGg1ZlJ/Rf7XqhK8U6nrW5NFDpPV9rbOAESfaX8J99VwA3J
dfaJcUhksCA7JnQzuMXAVCYVbwCztFYZcDKM/rehS4uXI4ESXZpDpCa4MxvvgV9g
FlUsgYJ5fLpPUxdCVeAZ4V8w7aWZ2AH4oAVPjxOrwo9CQ6HX9vuwVtcDMQeP8/X3
rp4p8H6fFY9ZdUsIzSGT8UIqhb70liRQUlS2lbjq9rdDinCVHF5MWRLCtW4AhZ86
RVykZg0/iCGCU0PWK+GhMWDsXIKLsDFqslu/d7hGSZUl5Cv8DmgUGRELi2Yt9SHV
6xGIZFIT4g4IeZWQKQFK9hMT9AfFl8uXYh8S1i/Dw1QYrIY+iyUt3RhaNR/0e+d2
DnKSu5XKA3cJ7JBwAfOBl3yy2cKNc6ptw/D6DC5Qx1HMMsqcmQfJMY425tWdpZaQ
VJHorrwY8du1wmtkECoM0NccqLfUnzJI5RhJJfL9AG6rIxGYeazeIr5dq2qJywY8
fV/6I1UtA32Z0RsUG1ftsxNCGLR4+qtYl8mHNBfqRZKNKvBc0eNPJHE5jPEkKIOn
6CW7DhhVdaEmDKtUjEAMlfrQ3o8G9x5BiR6WbZPFmx+ZGGHXiW3Jjh2jMhTBD3h4
N2siSJ7/05ET+BTP6oCC3HOnzg1aLlmwkYJaE8q2a/JH5NLO1dcOhFWCQC3vKK71
at6mqblm+221fYklPZ0hvmpPG8W9YlHv6YvRyF0tz5Tg0ch3pkLYtITvdSkp4B7/
g+3OdRk9/bsFRvlzogZSAwKzk02wN1lAdQD+ZLDOO0qwJLc2hTK4M8KiQI5U1+wo
4vHsyXevZ3pgpjGUIymWw/DHczoPdmkM8L4b0JUZ4b6F0LwGUyZDjVhPHu9bwkpE
GghWEYYv0yf+MDS+yTxPZp/FT8a4z1fMkKOah9Jqlzpb+PjYaKQG1VaEmA2k4gB5
PC7ddMrH61TqYMLS28wMGu3bZ2dj/k2SWw5eZExrNuXPkpybqWkBN2iYmgn1gri0
fDlNlpfjoj6KNdhVmmwTWUarlV3VjoKjP7WTW7OIOzd4Zi0PDh8yRisFLSSD7N7i
Ixn/WtuP4xJY7/jV6QFiVCKeslzxekpkBA2E60Z8gjeOIrmy5ronPxJ//9Y0uzty
6F7axgXBE6SFrrWtAnWnXvxgE0uvV+IzHcPkxmSHEfaQyxTQ7l91Z0CaM+jvEcRS
6PSuB+dJaqsRHyIbKGeHEM1KTats479fCMJCKg/ttoXoQO+58SWcLJ4V/J2GX9JI
LCwaNfdLKGc2YHSzMIbTxpTHyl9/Nqo/NdwE18443GvdjcG70ruCtS10ft7xhCrw
2TfIgs2ouaQ+zxHdlWdV9+znehCCI5jyyP3ljkurSjKJuj7di1RT+nF+mdFqi5t8
K4LPoQfFntCxq3oAk3D3fFjIBjM9lAKEzwm3u3enxGWrxIfiUovWtNT3JP7HQf5z
4s6oW1asmzFdNv3VhZL6YhB8y1NbYQNxEgeHN4QeVGVRg9FnDtI/GQ2YUliU0esP
kVRpfqVceEdgkiEgVd17Omdq94icF/KCvXE3+D5r1rXKbP0z5AwvTubD8uspe65y
sY1JwHU9/p6jpf35LdnYxwJgVQmnxvckP4jqvBNuYh3yBehHWecoN2KWx8ARhdm2
hB8gvykIvefEO2SbJOShQM4ht6IXGc8KSsq4KVyhFTThQxXe5AEQp7Gl/5j3bwsm
3ruO7OFkDqGlD9RosXdJhExDCoXpYOVRRg/4EYQijYmSAN4ww9qwhKZCRMF7zRLG
iCGw849UGJDkAynI0pBSW1MpoDEfgeyV18gG1AzCOehIeJhTGgJxqsYBZI5AVIuD
MDQ5as0VOq9hPWwtKN/G32dfux8enrmPSx+Gi7iQ5nC9jVCspxwdjkqNkx2HGDzt
NU+z3/D1+x4ggaCg47KbKC3Xry+Wh9hGJYhWvxbT/YxolokDZP9eyqyLEo3eU870
9dPRACB4/L/rNofy0kwZqkZcVHaySxT4nsJJfp4x3LmKxcE7b6ZMVDx32W4sMVQn
607VEr0ekYkkV7mgxg0k7Obyh+QS/9MN4RjtJ0A2e6FTNEE6Dbu2aUuAhmZ5IWOQ
3UoY0JF8wTZEf/p21eiFzStUk5DH92SCAIigT0Dq+2roBXLak3TH4B2i/hrefWzp
RwLZrutCILfG5bgu+qP4I3pmlLI2/Hl7pb2i/ZqDVv3Kb7+f6Qn70iuCufDbS3d8
iJ4Yg0pJMnoz9QVRiMaAP4YyuiPD246OmxlJxEY373q9PbSv0nI64o1k7SsKPDiB
HsB1RhHvc29Mns+CDY3LE/PxXCLHpFDZSykqVShDbMaFr6U4EJz06KOn1B9fNR3x
hhNrm9fo/vWHAF8UqCSRI16gkL2oU7rs8DL5bnGX7QiwPlZznyqEOaw9QAv7Wf2y
hYZHyszGUpgDqHZCWDkgwhR2yWLtg7jMHDwIMeayjzsVm6VJBohF1JskZm0lfXD+
TGtADUl1ROjGrpVH1BSjUxXZIGxXt5F1k0VrZzXFTDpnAWin7g+JPPx8GL5c7IVj
omqmx4+0FMYhbpwLZShMoCmlhKH7aQEflk0tbCLCiSqgkHlKHezsqL30EK1BSeev
6WXegzdip41eTH67DpG+hdcdedctSv4kqcdPwCep2CBwDwSA94g4jtOkS7BIj8Mh
kIw8WrTYN3joPX7aW3BCTmbrbhrQchFLP6mOgU/uKxY8raQw8y2XsP/jiC+C7DhM
ATj2udp+hvjQgl2vFci1JU42KVjye3jZhSkjjN6vNiRH2ETok1961ZnKk0pbIRgr
HZU5dHdoGme/2+M1T1E4QWlPPIsPxlLePaqFyr9QMYI+OiIFKXw1IoZkrtav5ppq
bf5U+8IgKzjOI0Kn/n4VUdVd9KFQWZ/zK2dgKuuMHehAddAUYElUMJGIJdIz1UWY
qkpZAH1AAH9xvuXEsTU+SSdO5Dei2KKBxQGK7aPPvByu2zj6vzlJJdcO+ojLbKoN
0aPob7Ocguykskl5b5TrqP5hPzDiYKqewk5Du6W9SPVda1FUiyt/8XtaBVNv4Qgc
8iedIqe6gRysBNREQ5k3iXZzQlhkZckjF3MAVoQo37e2sfX4rccQvrY4Vzal58c+
RySa1PrsajWYX3WHiwknsKjS/3CSnH7pIi1zIbDbbvs1ofBiJRzNgTyUmfiJGwsd
e3cNxkSBHhhn5O5BUJhUjUfaMGd5YrVtLk2wPJNdRje7k/wNUVVGBQhUfg2FF55D
Fyw06dR5zRYIQRYmdjPlY7LWMkcTtkro7m96tGkB1an3QHyC0FYKdUek8pdcL44K
Bb3jhJeahjY64lXCRlpJ/zl6I71MiEPGqHUPs6+WAkhg1KRAWzsC1RIq/krVYmF6
65xVZsQ60FBbfZTkgt2eERUwK16niYHLdOb9gFTsinLhONCp+LXASV60Dn0eLgPa
aE6qO1EPoffFzec+z0Mr1feHZNoInLTsGOdC2wFwmbkUz8kHCbMr3IBgGCCelzVq
KKMXcijDCp+nqDgtSKMQz9bK/T3lnzrQs3Qrdp8uL3+H2bUNudBuxeVTmK99Ih60
p6vnLr1FuBlilYR2OfkcWgYLNK2VLku5QdFqtrl9NQ+S2CfyRAGY9jK9MvnsFbXj
n2lLDgtyRzZpohm3QaLxmdbOC6JpKCh4V1odY56i7dn2WCHkiBCQwt3GDvZxllJW
qwaeG55Enliwx3gTaIlamwY8v1NipYOyn1ID5/NNBd+7H94HFM/clJOnbMzlJPDh
vFI9Mf33oQLYcbftpg7monbiyAW63bd2xAHGr/D8xnh9BvcCDY1ZKeXhCiM4KnX8
CJFlUXDuNjRLu1S69ku8WNKGaNpGCjFZ3CJtTc5f0Xjlp0OZAzADfwvZ8iDqT4a6
4wZgPyAld7PuhzwO3Cp5l3oLI49V/zZYOha2ubuIpWLf4X2otKAJrpJUFoTGgUOO
seW4oXoZ1ElQc6y9Fqfsya4KV/VMzbJNggL0VzJrxpimaq4rrPrWuSdn6ESAWogc
sauVcDvrWnb4TbeVJ9xkgsikl123f0S6FF3Sx5YUXdM/1tkEG5dAYd9gDoVIGTOQ
vJkndFc44gBJmAh1Ar1FBco6uqbx7oj7s+r5OHOiOkizypr0DJlPUUIlvmJn74p4
bJs6cjMqF8pJO0NuM4VMS9V32kGsAczdLgxUn6xmRRJ8KeHKPXDCq07aFCA4NRMC
rF+B3D8BGY9Bb4Ofd9Gb27XmNxebIhbmlOh5DkumQhH9KLl+xoST0HA/kWuZuObX
BX61ZPleToAMd+h8Adfrel9baKvk4jk0m1bh7tukYOJw71iSfrKupt2VNMClRBuh
8NqQ22/Sr/9zbWh7eAgOm2P5nXrC9+SwvoOlGW1lROfIOyey+nphxcc7IOmpuL+m
ViXQVPCeic/TG8TZ6RkBGnfT8ah4y49gbBYKtLK3wsst+Yr0c9XUqf3MGcz88otK
qFD/U0S0r19/wbtuOK+TLu3Q/V2lZacy1v0ybLnCqChWeiBnSapCAHeBl3kICMgK
Wc2T/Gn0mQ/7gY85xOokp7NAF5frhhxtlhiSx1p9gDeS4Lt/R4QFL0BVFaXwIe/R
kRbL4zq/7Ps7lFQOMiSEMdK5Xs+EnG5aEZ6Mn84Clv7ptusnSAF6mwyBPJkqDe1+
OMKJ5HIAUg22LDnPFBr9qhGNxx4H6uVFWyYPoMFm7r8gZPT6DtbwIR4X+xwZnSyj
ZnK7cHhoFtIM7OV48SSkDSbfIiu0a0zYvpY/bZia+2GAFpBk9EvSn5/TBeEWhJEj
d+vUu2oqCOM/r5k7XJgrMX6IMPJ7IUckKrMMOzUNEFtHsQATkSZsT6U4cU42fsaZ
tbtenRCczGCjeS5QtP7pAHKDwu8cphIMVeLybbtTxRwTYa0GMSM6ttwlUNaVuLak
IwDLlTT5zbx8j23V1qAv2ZDIPob+xU4STTPrz8V5ZDLJYyDwJ/OOPglzYPwzXY75
sCX6xrlTKFKSm22H3swwLNrwTFKJ9P1llxyh+ogICUL1JD+RqQEn3/qfSBbD0Jk9
EXaHqUu1/IPJU8ezvnZnNcT/cw/qJHsQQ3fZfujpuZezRLaxWS6zvNoxiekt5HYi
mBBwI9pQtYbLW+vdb2L7zuY3Gq2r2ce8FD133WAPJP8IXHBrHOa9/vTgrCFBzhxh
39Q48YYLx1BqwAOm0/Jbr2TRPcNmTXSEp3+9acwAHj3IrsDgNN0WtFyJ/ppV0lLR
V38+uPXm8jClhxQWGkC/rH/RuBJ4p0mIpCBF2+Ply47am1gyGaRNmWrlcnmhA1pN
jXwDTzPwwY1/CnCbdrUpbxz9JI9V/udAli2wOBs21RcxDgvE1eIWlnfE+t7FuM86
3UiqIyB6Z7WCQAjhJI8Tv2Z06diADrVrGcTYzEODGcuqIHm2N7ipYsjIJH/59q1Q
kkdVrrqWw3dACIZ6cJOP6ttxunW4ey3L0I2sQBsyAJcwqjsmklwC3tY83WZXjynR
BXaJIe8oElx0bbtLZjnzcoRk7vWuQVho8NX9vsNp95fIkbepfY79lJd+VemgtwGr
2eEuD2rBUCz0tgYwrFtU4T+GFtGu1bT5ghIzQzy5N9d6fIMV2p67OYFH0Nlg5EZP
S4GhF32HLolXV1kukuceEkBx2nI5hmjZuO8KQDwz2jqR0nS3LYJXvRvefuAGomqT
DXGLEgtj1s+9KFSq3c8tgYmcY2XBehAJt/Kyw3Tev69tfSU5RYSbeOOFYZj8zaU8
u0ZAvUigYVUWLfxc3+NfUFL9U1DkOTRMFRgRX4B6f7n3PpBuiOKq3e41AKctf0ep
t+2LQJuhqLvQXu9T/u1m8dsaj7MkgQIWT9EOCg2OJCMkYxn5CWjaX33NtHjnsGFj
PKRg9H7MqZTHTW97FAnlmDRsJg0EW6n3efVrEfhxfKEIfVpmggoz3vfXWK/EACQ5
vFNzfUQ/O+kZLda4gwN289xPiMNhBg1Ji5jbXrfQAZW1JgahqjsbnMcJu0zE5UhC
a9EAQhG1DwXskT4bi1QQWUbcDOcC9sIJAmWZbX0/yLgIlWqlAMC6QmItgZrACLKh
Bxr6IOTgVYf0Gd+N2Xz64YalfdjXm3UIuw1eNYKKW0Y9JzP5bHldYwGy0IQ4arfF
Jc4xApmq8LBDL8yU94NldN3Lb91HSzY9EvCjElx1ySH4qYOm5jraaX0awlgPxbhq
XLb7qVeTqLV8aH2PBWYGlUFdUaDeZLmRd3gGyT1yw1RFK1GDH3pNlMjntg4TsLLe
+XVxQqtI5L9+PudYI9yBedfAvpkNyh4oJ7POXqNHKiDJ5h0/sKWW2nKT/QDq4yZo
mlnmaQx4VSLcrZdA0saYy767YTEEETAfAJC7HQjkpmPzYyrnydRszz7AGfN9vS2Q
Oaoh+90o76ksmH/VCXUqrQLDo6zje+WF5yfRVvyp7mZre6I1BGvjInHJWjNG8sgp
1e8Z+y/K7omBnV2Q6wH/BG1QZB2RRZSEt9KLg1Cuiz6CobjGyY3OWWm+lgal6jNd
1FLvHKonDGCGv3a8ZmtxQ7SmopMuAWzlwdjCPi2pOuFMu8ApYGX0Cye29t19vPUr
OdU0bRB701O8oN8XcqWdJ+OBRYTfW4l+tBBnov++AQPR5rJF9pEtg/z0ueTJKXRb
djo7ud74n5Tb/YjdlfPUYloJ/Ydl05GK1lLi6vMb5P9hRVlsCjeFQmNcO6sR8eiB
b/yXQRQAGkQAF6EFBkb/f7qh7aK6iIj/pmPapLG9O1M+AVKEBntjVmMAekN2x/xZ
DskQGfwE4zOOnz3hHhC9KBVnFs4L0vIP5SP51PeoxAkDtdHImDRvkRMQLQ9o1EvI
+Se/WI9gWWuqrT/J9q7ZW8287o6xk1CZWC+Epx0EQYnu1vYXsHPH2ru3pqrK7g81
hJpLqPxJnLHddb7geE4LkxT1+e9953uBc58Zm/IjtOUuwK+eOYfK7/JFw2TbtX6o
VtU+kd8zgspUyr6kYUOYMtS7Giu4fCJIpyAfRn3k6ya2mkEcLc0gII0982yQMZX3
49YK8RQwLArVyEl1viyCfyWntjy0J+MwMtfrnES4UNjLoty010iJnruKdXwvxCNO
fKhWiCi7X7fMLvFmIHkkgCuhQNF/9Z74FEVGr8qagyUtYa1/XCKtd0y758IK+0Jt
j5gnrHvFg1MYTcsC7vNg140peJEiBUgCYNsgqYjINQK8s3Ks6QNB5ZC/ASNZ9CO6
4PcAjSQtLmYR4LD83Vj0HXK8UOSlAkLfmdX28ERLyXia+wEZ48dJtI09vC+GqVm/
hYwXLlrpJ+8zjX+Ez46FNYZfv2VS6Rh7C4u1Ak49rAVs2OAsBJnplAZufMUktRmI
u4nIzACVYTS/5SGQF5v3pUm2cj5HyA/sNpXLYNnqvYmNGPMNMdJDvNFQSaYf8FRA
daSwlKz3EjGXG4gv7DT9Vx6sinaq1bNZ+sINOA4o+R2/ggVqCDoR6XB9BDQGe2gg
VivdSkC+hmWS3Ep6L6k0NhLW7VjUskbwKTmH0JhyZwfslMy+tiqWIGG25hHzok3d
fCTQ/fnjeSob8ZGu3m6j94tgjLt34JjkfK+E2sv1Epg6ld8cgUe8aD70WJ4B+MR1
3sBPmggczNBpWLM4oDo9TJyYGU/+JyZpzbPApOoWj94Z+QI0rKJ7yMIB3o1aLSAJ
POVKqKHFIMYPSPABM3rFWcsGuU/48DCD/tUOf4tF0bTacJ+XVw3ebX4x9Vf4uFVX
regT/NOjhBUsNHLO0PYfOHE33rKrHBBdXcz6G+sCeBWvXinR9rTq8fNPOe64/kWy
Ik8JvN72LEC6CrqAK1JOJqSVRxM4j2g+Vijv5M4I1kTJ8Q3D4E2l/6d7WQylIvLQ
8ySZ9NIj0CbclMy/ARNadyrtPL9ZH7VJaP7iuoJSJ+k+vxdVPpg5E1bBM60IbVVn
zjOk4ncl2JMIS/sEiq/x270F1eREmMrodIy7EOAJcU3CvK2oiwLz0vz6aCRvh5ol
ViZyP0qSGfDT7gBlj+jNUneR8sYrmXSdQsVWDrSC80gj17m/Q2ILdpsM1eclTgmp
erJH2r7KI2OBixdIBXeLU9si1GMn4tHeSRjyUn/yFH6uLVmCPxDepoOFEEjRRX5w
iK7SnY59BWY4v4hqJoHP/X54HMZS11e7km+whl7FfsQ0/5dtQoixJNFwGaTSnd54
5SyIpinfw810HZoVAQa32wD4a5bXiT09Ql/do9RFJrp747dRkyF3u8FwUNK3FdWr
gEJ8MK9yV1XzN1bcTDmoCIpjCtxEtLTqwt6O5gxcbIRDiNgngDVKoGJ+xjAl9NFm
T01V7wQYB/ghRwTkuKUmSToeyRfnX9+IbNXrN7RdxQr5B0Y3mmnBCx5qklXIq7OZ
2EvwyWtet/4J7ic+9gyakeAJ6QOQ+IGc2uKC0aDnsO6CsaqQ1CpPEMJH1LLOJMU6
3JIBfOM1McoLICXFp8fGOfNuO07eQR8GJLessdNWzyRablfNrWy1eK5VG2Um6twu
qHMsli9kSx7uOLThNmJXyaN3NNkt+zdN8PMiozsc7USLQyKxhjeTacI/Otdy0aHj
Jvtzd9xSvppx2sGohDY94FDcfPJk2sfZjEvAIp0GFgbWvF8CBS3+ZHPfXO1oLeNO
zTHpxOPDZXz1kr7zXDjjhOUD+P/134/j9GC+L9u28iOdMxw07yR/QZLVp9blEANz
//14s8kpzlqBsXNUOr+XZZy78/E3t5iMSr35smNcKlPhGoNicgl3SR43V67Lb5MX
p1kWagO/gbrjJW4lKXvBTATSilKTTtGhNZWf7QUGKg8gUD5PuffLChnU48lZTyBY
AFDp0X6ADlsTlWFEVPDGU3ZPBjMT81XaSNfQnNPcv90agt49vhCLBta0ZQENkyte
9f1BYINIk4aha21XN0BxMwUig4KPQEwQWpAadzUlEX0xKxL6Fwmgpzem4S2lu84s
UgXNgXi73Q7dHp0UrJK45YnhOhZe/K5O4rIsOh84TGCenBZjksyvYOGpZLfpLFO1
Qx1ysN0bOF0LOvIHNGK9yqv5LprjiK0/yNozch6aHv/IsgYHRE5ICJXgLW7xMtcz
VRWGd4UIPvtiX2DmM9aY6CtfoGQzPXfxje0CCZbRvX9bif6fuiMu2147+xvLpfD5
6PsFe82ILf2u2bizJPZtmWjSu7C+ZR/xAfmOXqPpqksbRaxbq+jE5SDL4BT/sMj4
WfWxb43tlokMn6frAx78SK9erDANG5h0/b9g7xeCc3Qnt4kcr2i7uqmDkiy2FOTm
3FM9JpRdeMFfpt7vXgs7B4Z9b4EcR3hWSJg4poYKmznUET1ed3EPISCFNfsXeIyk
8NlNXoEGx92MmI2VPbTNPQnfP0Qgelw1vSAt0pD1dAJOOjayAZfCJ9rnttq//WNU
fFhpfjSvtu1atSk/0awAUaJdOLZRxQVW8EUFqihDNrukNAUbQYULS7IrKmKxJmc7
66xFwxFXvO0HrMPQChtZqqRL1P66EshPxir9gzY8V6xynqqexrhjBSe5IW0Jd2Wq
4PxUfBXJ5Y6xhHiY3UM71I8jNuESSwAXfgSBjlntD0h44+UXiZQWsIPObI2rhPUl
foQFMeWett16wIMSzpzSHA6qQDkxvhcCqgViLchYbSx5PbkrZpa3ByPbsmKF0YSs
f6Q0PXmdFm3dThfty56XgIraxwUDXG/iO2tLuAJxneHVO/NFmBalZbZlEEScNhmi
yBEpPYrSfU7iCFIxBeMsDuCT3Pu7xhHkndCw90rcIF3UW9pzheEA528QEpsUhqnz
G/0g2oxWu8u4G2EhCptYzhVQk4LfxUF+W3d9FWa5QGLzEUk8IE+WfEh7jdqAvXP+
MyEH3OZoaq4YAKfP72iYVZ3njhQEyzfradV+okSYo2FS9RqXDDMHMISOJZQQlnFY
tqvJvy7aEaMTR8RXorlMUpLL3yUYcMIRpd2TdPdhN7IhSzs7Ab1S90esCjMN52fC
UGIVjYw+wAfWqBSEJyaN6tHwLVlDNQ5eLFoHDvOroBHNTQ9Q60RHbERlzu2r0O9F
FAbeUXzTtMREz2Iil88fYCKYJwXVFroRYSpzF366QX+udtA45hkvOpePZuv6PgYk
C2H510MQc9oEul9cyCCJb3x8TUqxFeBN2OTuuv/Iy+pPjRvkGPPbZ9/yMz1TLwlj
Z7IbPe/51C6ocuZL8sLJvecrHPA1wYLIh5mKlRjsZxmmWZMQiQewvCttN5HMe3JC
21PDEXXkAWvtZUXRPh6OhpcXS6l4CF0s112fPzyhwj0zRs5SeuwXQKGR/e+a5hJa
HPP4oW+1s6umBbFNrE+2tfsSVVv4LMyTAj3kK90sHYRKwNOeSKhTiUTp5Ennj2gD
EL+Up+lTeK4vpjqHtEDReDp19jOuHVVEerxQcL5FfsWq42OAXy6tav4Wv1pCY2XH
dZqhcWfbbq/quA3ub/Zl4AXLKpi+hVV0zzvKq0tx30pL8U15FTwdnPgq2WIPkxmZ
u4OWh/JUs9bXzeMHiTmwXWEt1BJROIQpuLxBK5LaPZKBdR22mjr3teYEWjaDjK10
02s+KQz6Oyuf8y7/Co4ei9BIyLwzBBLGTETQ8Gadj+zQy6iouG+mxKrXFUYAfzMG
/mO96xo6Jmqbj07YiBVNVoAW84mun42wY4CdEHY8P2t6ZrZWoMi7aznUnefH8Llb
TogiUNg/N+ETm3Okh/AAmR0Qwkv3pDBNe/tAuKmGs0mWdDQGgmWxw7SlW67vnl/s
2/Luu8MMI1J1WzEG6lE32F0dcaNxP8y5Sl22FURo6Qh2eAQGEjZ6AkKqnpvN09I+
s1zMiuJhLpvSaScOXJXgZrErXVeeWRL/NF28s9iFN8VgWsjgsvk+TNsEEDFBjxtr
n6v6EXwyD3MnXaAyNpsF9VoZHHzfZH1OpEwdwAJqV9WYUJheen1VTjE1ELXQVsne
3T8yptXwRPpR2SfY6bkbjrpvHIasTKFyz+JBpHf10nb5T3wRz40D9pSyFqPxw+Io
DZGj3jFmAB7FxoGMp7r3IxY9sKu32Pmojuy3UHVUApTFK5JKRXaRLx202zWpvDWz
OOC43X3U6WNeohHApmdXXLB6AN6RxirpT9QM9qoPqQoUHeG01c0Ny78K+O8sCGS4
xjqvKKTbCkIQEtvyJXb8k/91FN23b6K76eURbQ8nlibAtjcdSJP1sALd/qkZ66VZ
Om67stOzxehvS80sO2SeGHSpXOPR4/9WKz7LG/ouGJv2QZ6947fOxK4IOldcd3Vv
46I1DDBpbU1Qh4RqJUJxPJz1bxTrjRpQi/aJ74LfItp2Bp3nbMVEG8htE97v8ndW
MGyregPLHPTzCCs7EqSilDFJfBslwB5w3vvs2jeGPeadMGvchYb0A8DHEd+WqqYx
KuImQ2FA2IkUDa7TqBo0UcUoiL8bKOp6/c0MNMcvjAC/blkm31R6SX43BxbEWYke
Bb+QLtyGNqInRp6W7V8U8fWIdQjCT/b5xM1PmNEDfhZIpktsfC4pB1sncFirSuJ6
Z2vjFjTEraCvMCIF5/rbJMMPeGKBElZXEytzxgZtvcKgsdQbeyGJ/oPsmJRaHzT1
Mu4Q8cKmWpEra3ktWLa96+TpS1iOKl3bh//qk95ke2LBkVBokT2csrMWY9UuXjiZ
pzgI1muLfYDbzrWwIdSn3MHBQKPTnMAVsnopAFw395bpDOhC0r7SRKRspAoqJJUw
1k6Cxo48H3QmbPk6loRV/zOzftZQHYjdo5d2EePbhdEu5PHNv/sf580QZwLyQVfd
pfipzQGrGF5VqJDd9kSMJgfno07BFHZrm4NVE2e6fvcb8GMnhj8Mr1wphfdQTLnl
7mQfcNBEH8+gmY7K4pv6Is/zz3WYLnds6s9EaIqv1wsMet0hnHVgHC9oiNUkg/B8
8t9I5m5vlL8EfLmlGO2FWQXnBWmXZbrUag4sBc1z3gtwpt/KpzfEUM3UnPKf5/Ez
SkhtqP7rlD/6cBMIryfkgUVRBFlQA92fJL+noClpvi8vrW/C/lldBKfYr67mV1iN
5dQvfZnfbou0Z1gwVNobg4DX3MQLv4nl9B69hIRtzUHpmgITM5q1rsEDmZLiO7/c
OajQtRddHBF7fRH4lBNGLj5V6/A6cvbh1bYiSKAcjY7G3rtYyY6fdQLoHmxBzKYg
8V3ejs9ap3N7+vDcg2MWyBGeUoJMnRbH2kWI2J3tyStk8AwFHxYDGVNsREA1hyXP
DHZEaxAVkZaR3TNRwbEUWFKZ5+wSLLtaFJaS31we97TjpumIquTGgGvbVQN2G7+l
lumBMdALynkdyo4cGvHtRNrWkB9DMhVWM9l56PNLU8o/nKEJp4OenYnLdjDcfSUH
xphRo4fsJAlNd1h/9edd1F41CShsWj0gJkSKIex2UZ0IgItDl9BjexuqjhrSIAaL
3tpKCH89CrJvkmWfmSe5z8yQfVLNNTCgrcYTPrrEa+cHYEz5b0qtvvvoJDwU0IfF
CR1f1Bzbqa0mw/Jrgffr1qe31oS29ZA82BaxzTS4ATDZ01zfm0V2+hy75InlwxDE
BQRgMjqxQn33NC3+H9jRyV5FQ9oSl6QMAOg56ToRJp2mnCBk65uQzXoknzpzYKzr
fEd+oxTVjAhEWKETn3ost/NMdl4q4WfI3QFmcLOyX9DWX+UXAv2jh20Zy/FfPTrv
9qdeOo3gZ3fW1FbL0RyYCVIt0YqHQ13sKjZgkgvaqR8bprqEjxuex0Mt5IRwzrKM
iZW7+teOi3+XWvaJA4q1bttrINC3WJSyDjN9VjsKKL7GtPJitSk3nvG4EjFUnMZg
dL6R23N2pbaiCXVLVPnDmchoHh69yxOwZt24v48Vm39pspKX7aVH9pZemDsOVvHw
7+rQhHDtYHQutUogZh3Pe3KK4ypi3a81HNRvV3/huu2WSmLap16GrGJCGKnbDRXZ
4DUXfl58pWYL1lU90doTesgOe+jtOHxVf28orRNscsE0QOwIkzbUwAIzHNi165ji
/7okovDP2sg+rG4UZCShH9ewURZycqSOgCBUdv7J9R9dDvrcsjWmn75H5pDGL4Z4
gBnFlGTEg5jBuRi94KkkxugwjypGk5HlTZfbyd7CuzO/OhnbDDWmbv9RJL4F77QK
i56kYCgGpmPC4OW7hPmSCbkkTXJtoHYM6PPUVPt4qvQWdFCNv+ArJzkyvaHRPXyw
cUm4BGk5m666WyNSMH6sPdAc8dwsAfdnkgjiN5nwJj5R09jNNozuqUoZAGcSfNgz
WxDEt80ic+4zy1R4YqO8HYJynO8wAqDtePpeCkEL1yHMDTaV1PzhCXDTxiAwWlbM
IPW6YDfS7101XLR5H9i/VX6/k7bIniyH+JFaUUMjEl0wnkF+71X4iTD1cq2ladYr
Xk9joWw51z5JXVxyV5/YhUmjFykU1AGPfYO5o5ia69YkH1OjB7eHO53WHzZxkpr3
wMUOa+1DrB4wUohpR3oY2qSNAXe/qijMDl3slmM63hhJK43JYnB+MaLIOUJ45bIp
A4wwB0w0IzxfJgf/1nn/mo0X/dy9P1M0ZzW/gbaeshsrKkoqEInh1+t0kEC/3uex
D+bHA/iFEwGuI/zHj+smWlvfCZZZAvTH9U1Y8A6z2NzJGnDK7NkOAh+SfgD/JeOh
1ieN0cLeqWm3dVA1dvcTTt1YqMNCXGAUPxt9I0E21xYmKDvQ+GNWFdOX1OHGdHmS
VqpeNe/YTDYDPngYRDLttE/PChWUP4+JnY6j62tMoH9F6hidC0Wuhb45MMwMWP4l
cTgYtBmplD/p9fz3AcF8DkrQ5LHxYfLheEB21iCzXSe25fZJQVHF6Gvn34XTWOSq
4eGJG3uTSIcOILo1mdwoG6gf+eXkkYm4ahJTk5fn0T8nPVCgO5+n7YjBiWXNmVsq
Xsf5sgZOB+g6Y3j8NRA1bk7t/CcJH7MpbTEyrQ0t6j6Hm4epXe71gQY2TM9hO/ez
/EurfUY+CIcr1vYtZGsb6/aybgP+MphaHHopgjzte1Y5npyTUoGVR9ZrL/i/2sYa
LHOsAog5QlNvpIvtiwcTqPVrIJRrRUZMdcumJepK02lRTBocllymIBCFY5heercj
+jE4y3526JgRyvFZiV2Z5eyS9+ECH3Tj/xlOb9iwT0TcKSU0Vl+WAoEU/GNfsChy
BTt50sae+mcG+yZn12zgtoGP5opxRSl5oaYij0NK7r3ugWmzdOHQDU+X9Hp/x1lN
UZN8gyjR/3ugw/B6XkUN52uo0pZWDWT4l8jsBIBdEzRtfv/0su5szDU51efe5UEh
ZRevlvhbMwZTMImADKXNSII5h9AlY+IspVcQQsHMFNibqUvXrP+fCaHozoQF051b
vLNs1BZDfs1WVFQlXqWGW4i399f0HOggtt3US3wOBpZHF0bq6DpC5zz6WDUSrqKS
Qv6KEfruv6y2Nh8U26b7MTvAmfz8u023bbFWYw7B1Neddda6kjoIPiCA+hWiLTby
QNrkdcAYhg1JneTd+mdC4nQumvxN2zcwpbN2urCGEMFBlJ/WrBpn/yRh1fBSbLWJ
OSOKSdQCp2RuuQnBEZVC5LoWLrPzqWY9HLf3EUttGE94vlARYnB+1enyYPh+s3RB
6EXBBD7CAX/PuAY0R9XjO8nRIt0DxreZuA86G+uJEKo3PUdPxqR96pXyBBNdt4W/
WKFluq4uTgZtei3Xn20M4H914vjCvmrI+wNlXOkRQWqgqzGDLvzE5+SlakpVgyPY
UGbhWd6W5PfLStBbNeN3Q02kaxlXM39FUiWPZUe/VBgLpizrd8E6osv4OvOMzXBZ
xI5qC39FJqyN1Ohz+DkTdY864WNizqevSnMBDKJfW7tvgJbDgIUJkdBg2z5VA8sY
LLHnakR+U9MLxNL+r2i8yTiRLYrGPVYf2Xqs869nOJ3RPh4xDKByh2uo1DMv+3yT
5Dfmt+Y4/qLxsi0V9yOC25sqlOmUQdCYGlNP4TwNyyPIi/y38udePw/jAwii2sRI
KiiwX1smH4TGvWct7YQTtBISjz0uJR11iWbdaMt+VdlcqGkrWzsM8J1oMYLXMs/b
Zqqo4k2+z1eA2tPaQQzNNinZ7KIGoEzAqJIUDqVzrz5MVZi+cRMg2wpOYKwD4xIk
Z4hGZ5gYISPyicpTujVikICl9de/omnh5msOqwTTyGirb/BasHtcQ8NVjcaeragy
wjPn5LKn25frzsThxCUjYan+UXn5HsY0j9hcHR4SOQPh24ZwERICwAfM+5eDP54L
N59ix4/k/6bu7lMjbceQzdjKe1ktd+m6YbYJeGs9Ti0YFTSaywyGCulDmUiMwOaE
xkbq0Nf+ag3k2JTNquGsxpwnk31i3NB2tTHHwMIiIx8wj8tJtfaAnw634liUN3lk
9h4c2Nf3SQ2LOmsnHUhbzkw6Hr7tRp83w6N5NRO3S0D/wbAUG3Rzk20UI20jnkdN
TvOhLWxlS0U2LUs+kwkER7bmrD74iEsHFJdXHtm4u/oS0rNiDdxVzauRRTBaEkD+
rjEErqjoReNF91q0Za8KcJKlsgpVNY/D53Uwj6dLTYJMSK90Ia1BOhTWBiqznttU
cStwJ8QonVHCLQmnkz+B4HDbUiKIsPN/TV1maIDXycEZQZyq/A7O8PRt6gx5Fe8U
9elzZZ/3NzUgQHPw9YePj9ElRIFkfLuhx8vddFFcP3MtfU7+Xz6EsVtqtKMXJYTy
2oJVBm9UkeDHZJWpLIIA8inWH9kDdxSofHdnTOe/DNMUQVtG3hVVHohUF91sqFTn
yBtCj44DNtWOxxzd38XyCzZgU+EEAt7PeBLxfWzDBU3K0PWZ9A+PjyyUJAMgbUTg
AmhzeSUZcodeXvDWFDB2M10NbLEW4DydORyQfT4dul9iLVYw4d0lptopgQ7ztTg+
M1JMAdxJ+Ac3rtNJPDF5X6P/90BapRlT0Jy7n60AHWJJ63JlPDm7PyGSLYxVDs+A
33qFBB4zEmUK3W0xiwsG4rPBZhqhMn+wv0eZ3HnXPdFoVQtxXgN9V0B3I8KQcTPe
QYCiORZKg83d8lBmAcMyVawBjuSo+K4HSDN7/+PzodJy3vcvUKJgSAVjOonLq7bI
FBQ7xrs+7mo80IGi5mSTBQIBx13Z5V+Qkgsfcsv/ZeK2sLb86LDXtNOohLVmnhrZ
gAdgMVfVmEWhGw1IfPKEoC06LJfF+SKCB4sQqF+w8Q34+zrJhbFNkyHWskw6X/2Q
Wl9Yc4UaXwhf4qDgZ69xbpqlyjJ1rbQyEfPCpNzTasJountFGZlrG3nrAHwHtvdR
gAJSEwLX0RxHmiH8LBOzpglt6ZdeZDEGWJP1aENWmoDKQ1YV0oBgn276nhgUrjnc
ZqxX2tufbN/uhUOIN18RElQ82suzN2+U2LrOcuV6a6w2eBgnYxHur9zQf7Tz6XYG
S/ad4K1j24+4Apnrjw0d0jXMBmsITqf8NUTcJTQzL15KP/VLMstN502dSd5qY6CO
p2tnHKKUddNkBkKABsxE8f4WxFkQsChuuETRTFrvB1kvxceLa8bcXkyXTo+LnqA+
YkHvRyHY1kwlpHg33Z30anptNSf63ZCHYCPKwYPo5zFMu1GxHoFlsHKgRN7qjXS3
Qu/PwYFU0gaUHQwzUR+Nv5SKibajSR7oqGh/AZKSmIAtUAfOCPhv41LkMohoni/c
sEh6f3sHlLNv2nvnBx027z66REHwvjVG4bDlOjpzwbmSGU2zIaWiACtHskyR6AT4
5ln+zjJ5KgXFwwew7s7fCIB0C6xwe9WG4n93AEn2g8QnPDW5y75ExyNLODsuAT1v
nwURyXBa0EMcyAAI7YE08xehAMgYAZym1FyXHAawbtIfNGLHbLzzMYgB+uKK3Ppa
ppUrPEnl/TXlDiUzIhf/7kkDYx9UDTQyaVX2VSGgtRH17QaDptK2VlNnCzBv/Ud/
FRp5HZYu7LJPaRrOhTBrNhGO0M4I4SwTdLSl2lo972wJ6FvILdxgKXsdD5TkOb60
MrpB8S80D5ssFM2uuEiRzoWepkihWMRl+szx2LhprDv0JX0kOE7/jEfeHMfdnnSD
SSiiyJsE77bmqxaGvKU42o+8a/xJT6w44MADgBOsNr9eofYxsjmk/fYd33ngIgRU
0vUEjRVLn9+Aj3L7hPmyRs5SMBeVtHtfBQtHaFcySGmHhvD0mMJSECAkenfIO1Ej
6/JtbOo4kg3IT075Q0aq8zFaY5M0KXhSRMPCWc04Ha2roCFV+HnV6R6w+nQ2vhkV
RZogvezvYpnjhk2pnePLE6arY6StpNkJg1IiZC7ULaz06JQ6nHFnbzhypIJh6kJF
ZZYdWhUemSoIUarinCttbn6i2x5sJJybE6ZcM07SRxOll9WbgsYMmDfG2S0JqCoB
6VcousPDuYcgOFeJWLbiW8SeeAySPWtbEEG7Litk8oI4+I91ydDK8awVmIQ/OEPu
X6RxbVUTMqOh5cUAMlY/khNkrzr9qNEnZ8aCZ+uB3nt9Z815Fr+WJ1mJk9H17DxH
m0o5CBGeKN04PPuUDoP4J0OvqL89iso1AocKhptxgoC+lsp6ZxJuLHHksEkgj9A3
j4THPeEEvAiZh8Ydfg9X4UzkmRQU6MTjREMq2j1Am4oO88lNQRup59Te+gWAVKiz
vufAjGSRrFuiH3BQStBJ9GrCOXQviyrlvWPojBPrbUYehIFPCXYj17ucjdKqEBxF
pKS4IddE0chHPHWMST4tnhIC4UQm6+bJvrx8TRshgb2SOyASvrcc/HQ0z5u9aO70
CYIn6JgPk0yIPAXxrFPffS8HWUtxS8QBsfpZ4MF+b06AoQgA8V4q8I1Q09Jvi0eX
bK60agmSyX0LzHkGfnYzJS15RzMpAfCMtP/cDz8KqipTSak+K1jrk3CuRQs+LYeu
Zdi3bncjDecSbdNQQwwSdgRa8Bw17TBzTdf1kvJFzCaMsUFQWTVE8LZ8w2F2vwZX
T5bO+TLBdqalWeqdbolmdquiaktyDf8GnRFBuK0ncS1ttHIEpSi6fWeIupXE5OAn
Au5qaWJL3xuwbdKwfHhdDVJbyWIa5lFecJ6crYMW7nPEhMi8DfFm3niMOf8/yLmN
RybvIMunEUVJftmrfbsYySrhF7bGyiOI+zwLvqAY0jQrD0qwWpdv63REGr8WqXI7
bxiJcQBaK/BRwuRT7TC/wbp2eQVP9X3Qe9sgVlfcBiRqmfjqYABT6N3YtygOXU9j
f2xdysJo8StTVid2aQkDEJANCHV6ocHSPuL18mj+n+4VDnkn2SeOnYV4b+tNKFG3
ITM3FFtvcrpWiyCmg6c4xjhVMXhLsTM/TwY4hjGV0ZTicRKI36wKypTyoy2+8Uj/
gxNEnEg8iRSMzfPZbgxaJYipfdx8Ofnr4M6Gg2ubD+WwiUqBXtvqiAFkUcL7CAh/
wqQoeXSvbRaSVmgJt2t692EnCSrcGl+5Cil/JyZDF1DSu6xLWP6Hb2AgKM33prQ9
D25IfzD5SETIgpBDy7UN9hQEfY+o1KfBFQp8nolToswM3f7aethWpP4eQ52YIi2E
em79Bd0s0kr5bcrkwVPMYnwawG+osO8q93lh8BACUSCOJcB8ZEz9KCpBKWqRyAVM
ppIccp1ul3qf5jod7EzYsOIFirgJVZVhPceYYW07ZAFqCFc016s0ievrf1ysL9dQ
hzq/003FNEHjPhRM65lQ2g58EOnNUXf6hkoRgBMvBdhRy2e1+wKUJt9OBQKfIn7r
lybUMihr0C97iFhXxsqF3iuI26BHnKX3Mn1USHLTDxR0XeMIolOmrqjH6nEz4meF
4vVeFMJgLzMjv6lgBnoZR8wGy5e2v1VHuUoY01yDV5w+6DAR9Nmiw+JGhYEx1NFu
UYBe6F5WgnFwIwR9CDKZs6sEplDpsQq7evtkFKuFz6k0e4OIcm1u5oeUbMtDak+M
3SeCX5tDoThWYdboBpH9GVjcnekmmUXRtMnNI1vJ9QwTZhzpbPRdn1WQQr0fyXo/
kDafvPRePfX6c3Lfg2cEFURYYKOyCydUSOMcaqGHzOx5sRBFORiQ81Axa2VRAFwk
WnKAWlzm/uQJQJZs8wpZVZO91NftgarlRVA+8rO+CgogxfrR+JMWKcqZQ5Zk2g7s
WfAYkv5B+CyRvk3/h0Blt+BdPvyPJKHe0utlJUuQPGETsakmczXkVu1xvs2GEwmf
Oy276bQgFqs60qifNJ7WRSILuoW08JounWmpJtt3Y/tyuHsMj9muNJiKeKO//45l
MGL4zuuXVes30P1HjcpYu9jMVp0lD04kupHdeaPso8etYTwn80/RqM6/Bb01kHQP
ABBjGmo9am814FDqsPD3aAVWR+NLVsrAKPbGACOMa30bgr3PiCGs+MJPLHZcyRwa
P9xPClAuj1kRdzThblXFfWA9wFzFQsrbTEawY1FivEHaTNkPhD/4xRLX9yzfAfXh
81UQkWHLH3D+yHJ+E1PxONqpMmQCXfHzcI81uHgbSx0VCjbdkfX5Nk/c42gzSWHJ
XDBQTxIlF2XuX0AEwePK4VMj91gFb+Vs812iviLdZpOH7Z4hGwS8Y7CNQHeG5VKa
L/zG8SSbvY69SiVZWPihmAK5ktN/VkX6x8itlONKBsSrpCBw3pd+VoDUET/o85Nw
FEk/LgKBpbgIKU28RaAKIuHyDq7oCCkAGMA+sG6/Ri1sKVBQppz/Dkqh16x0dkcZ
3bRFtwrSdSDY2wkofa//jfWSla6PBYen/vS21dAitbpWc30o9QVfPdloA0rjKkWF
wMTKSOEs34hGqfZvyXIDhccmT3QEL2lnC6xf5rQeA86LAjp2eBcY+kzcMP8GBx0y
nucCMINMbdZAQwKGxfBCFAhVoYjYihZPu9qy3Wc/vZLovSswC1xMY3yl6gh9lZCm
g1vWzlk6m1w7NydtU5LvCPyL343GxIiTHCqZgDNMbAD4GpRHJGh4k6jWGyRlI9AH
LI6xG+Rf4f+Fa3SwY/X/sn1Axh8td0MmGs0eZCSNqDdJLV8VnZehfdgqEmD4Kvqz
aGckyFJcREUOQ78aR/aDMSVEuh9qfdpT7dvsp1D0ps/tjivsn45FqpzzHuJtef2M
zW3PxLwVJ5/Eft4eE/rlpA8kxYqHltmMf8eNklx/SZL/zD5OZkDaX2w/QVYabL6G
Py8E7zUSfmCf7cswwY+IjJf1ZFp/9Z5091DG8UHhlPFZ1Cy6xywaxuheqCIPOMXK
xQz+M2aUV7T3+FNIftDtd593RTnppxMCH6gv3fLgTcPM5CZIN6hGmlNL5O7KWMAR
1GYvAykQE4jKf73CeRPjUP0tL4nKregM0pi1x0i4XJmhNqab06BhhAh5D3ytbi0c
T3do1i36EQZTtPbltGpgKf7jrthSGIo6qRd6/MjpMV3fLMaz9nRV4Ha9M1EzncOM
TZyTR2cfCivzKWNuXVr1egntw3NdWnje3m67YLv2yerXPL9Oo4FcciJNgCe1sUWt
WjKZn2dOlOWwdGiENyrggZ2fOAYwdjUyRGzILtPQFi8j2jI9nVFFuZT4RxhLStvr
1gqPesd7aJb3eC22OU3H/M/jomO0q+d7vQAd85oZKL6U6DNKxrgjG7hl70xWsYnD
mj1WDc1y/H+yzcLIt0JmhbWeFVxRYE1hJZ4l9fNPSfVgiULVCqvD+FXpEAbaOoGF
gGUfRiHW6gvfFcInvxZ+EvRV1HhScEiaWe5/JGc9jwQ8lTgV4Z5lJJdMNFGVu5h7
B9ditr/gvwW+rGS/EorDQIQsgYCyA3n6IXkp1l/eyCFYdaRm0TwtMyjkuNvfLScR
gN0IqOW/pW+NorqvDfdeAOKF86tgJkj9v1uSLd8D3bjB2HXi2y45Xe2KBUChKnBt
MmLoc40d3dRd/pVnEzpMPcWmEm/I4Uc5rMFb+ErnZoQ7O8kg5ImfqaT9SYCkeSai
LJ5KvU12EVTp3NyHbxGM7xFVs7lu+r5j0OAwnVofl+fcxDXARy6w4hzlMhFpRDE+
x7Ikbcu6UKZIJwKmKQNnD46m+VrdZd8ElYKZQELSVOExBYrb7abBA3M5C96NBC93
xSK4dhsANK/8xskNxpmtLFvObDo5pQx3OgK+lumbdPScrCvAfYmt63KJe6szJJni
edDoY68q0+axJyciR/CYi4OPezQyOFcotlnGaIiezqaCFnMZsVmUxx/WQw3xbhds
syITIOyiKlDch8B0Ilq6zI5fqyxXINYoeYeJzbFyeLaLoWC0BLTGJ6iN2h3Mw+eC
quPY6b9FxP1oE5CUq5DyoGR61PigLE8ME2whTmschBXHdrFhCXs+B23unpawK6EC
Jj5ULPShi6uhc1+b4eH1j6zo5oXJYpkBuYcgKVsW/mUM+KOLa85RW+6SlV5SvHd1
7hqyX07NR9kgIW4KokAcoQvUVrxKIsoKOGcb3hnkAL27o35/fRV7SUxB8448AGMq
8cCa8YijtsXnUEr6AYBzVELXudr2rWLMoiIqXCcGVkF7tMFVGgLsDskcx1DfSQR4
37+P8VBuFsVj19IXneXq6myRrvibpylp2fHkgAU1YTkqEFKSEitmjZT0sPeLfpGR
f2FyVX8yHQBEh//EbaAWAu0r5aEnuropnp4KP/LJji+IGtwwLgjTstPtbSD6U0WY
k319UaHsoNZsEil92J4NXFsPQeOhTHeSOotXS5zaPVb3Td2Eikouk3V+csbgWn/q
jVM6mst9gskLW84TeOuVU3cJlGsN/uUgHfWfQ8Fbu6hN6o2VSPU+jmL/7PvB7eGy
v+cJm9T02ip0pvKO7GksDKSuSeN7G44gK1fGPG5amIwpo+F1mroY15SEK6y8ZLdd
BMJRYHj3jTc6O93b7S9EbqMCVIixNa9RVumCSPIE1rulCRmFk97zRJWi/Opoi+Ho
AZnNwrvrEuoCFJw/wCeiB6bpK4DbFrudl9PbmyfIQynzSUc/nCCIadKglUccWeS9
xoePZxFOIZ9XENi+6u31cINLxD3AzbD4fd8GITURmWT8uMwncGD5xUIr5pBNauBu
bQlZAf7q/w/D50GxugezA/oUXF9t6i620m6Rhv4L1BMHcRx9yCM+uwO1mAtm89x2
CLRtLUoxX+nHrdzrM/+GwJAcwPYTTehVOSztrZg4CdtuHhv3XDGoDtxd6Ouj47L2
OdCVZgbQuZnuRkgAhE/ZnPElyaKpkM6YAVZHqIUDwhHzdgIekPv4557TjGT+LaIz
LQ0UeKYPsRG+Mebo0elNCV6Ql1MRW/pgGyc9aZXhBVjUnuJErHKffJFKOZTFMCkU
vDcI9vn4e0KwiJ1pAYLJtd7ojKi3VXmkE3rP/3oNt1s/6of4Cltj4FCMEsv/8jq4
5HsiIO2VE2FvC9gvmtfUfo2eRGb9e+OGAUJKg4FTBfcvE3KxgOhMoz0S7dUtusD7
WVv9Sdikg3EGQrJ/e3mux38W9KdzoScm90+Eb5LRFfhJq+3u322wQEdFf2PsgovZ
Spx41JurcG7zb6swf+4Zo+2uGB4AXFvKV1IkwzXNTBVxzAbl76yV4bDnPFgi4gN/
033u43iEgoEF8K1iW+NRV78eXox/L5peYY//4V/7PHdABa24XtNjvxT/etEgWh49
Al0Py1wRYjEJfmg6bVfSiHzbU1gJIixvIPaZPuBAxUK6WmLvdnMxFicDSRNFqQim
9vqdxpEvtp2mnxX7aTU7RrcAOiuEo5J+KpM238WaSOWqP5itAHC71oCr14iYckj1
N5f7MQa9vXjh1WZ4kXXY9oeHVYTPXv91UXt1aHguZewNbLq6CmiMZvOTB5M29Iur
Dnp1c4vBXr2QUTIQ2emb8rB/I7viW3Cxe2ZMlXpcY6RCWPCxoyd/XeBimKH13KGA
D9l25CIQE3tizlMllHwcom7XuCSWDo0XTsA9e0NXTfg+MzueH9xk/5QgOZu6d/Of
8Ifa0ZJWHeVwxVwsDIeoww7VseN7VH9r3Vm6sNPnHwaEFSAOZOujLHfQreVBgT9D
zaYA0zgZQbCuECOztasS87AockLiHkEfs+BKaIHNNRYkWJDxVyseBhwz0704hWBq
bEpsmxvjOcF4We1KxPuYP83Ffe9pLCfcRGH6c+ihFqOF5xH4bgsWP2Xec32HeGQq
m+63GxPgBZqehcimCprUrR2XNMpNd0+0pWpEnC0BDM6ypl7z7mX45vWqFDpmkKTL
/V0U9JniRiqKwvlT16voPpEfAa/rHjZPb/oOG4VMvDtgz3FePUkL0rxfQBZ2e3NJ
4rMU5+FutkhkcywlGNkaviJawz6DuosbXtPhe5pCZMec73/rIebGgfn2Bbsiz1cz
fWlWD0A4dxF2OkfWPhk7edC4o6vVSFLk5kgaIfVEe5C1oTK/N+E7KzTVj3hckeva
rBaWWIKe1nBbOHqhBZu6p4k5ZymJJpJtUy5iCIfvdg45sIb2sWhKxH87Jg96XVwc
ttcVRpMkTEdamQDHco31k8YDuQG+aSfSWOBqv3B4syEuJ7tUj5HdEjlCAmrssRx7
pkaPdK8oFkSkJuMf3Kt5j48ZDqMI9YFoALSQ4mCfkhynNEK/juPskdkSKQfoAI29
3WCSt6q3+VCkjRlZK4UzrjP09INRpGjFJ2FjE4a1FmhNLQSDDor/g8n8BlCqbAtz
qM6cSJupb3oh42z0vMBHVeVsxDvg1PMF8y5zSh8vusV8ELy4jaZzBHJ3pO8aqQL5
lYpl53AoDnjxN1poCG0n3nJKBNYDE5sHnyrk/lZMBPSunBKKUs31MC7Y/LiHT2fm
XSC3+ZnW6HW61uV9zcIHtilaEEq99E33m+9JRYny2ptpYhB2+KekFUv/x0nMAdh8
mFIZ427ew4mc1TDTOJhvQh0ozYEEauEjYG7VH/vB9gzr9lSYTejv3RDbJHV91np9
IWwlMEkko+pwuf/xgFDkVLrmgu0+r7yuuCTJ75slNk1/7xasbWB5tTBZ4KRsKtLZ
Uwz4jvw8y114uDf1wFv9EgtEGk3XJ12Yzbs4/5YBJf1ZZZPlCEuibV7J1ngP1tQR
bYUmMN2wzVb1q7b6fNYMHZp+EEIjTtYIrqwuWlVefZsQRAqN1PsHnyCh/MCzUqaH
dOdu/vEpR7gqFPqJQa1HAvQ35XW1ZaCBPke3rXnSQholMR5LMHd8GZYCbmzkfLB9
h0p8UTnRBYhk1M9d7DRboTKTJAhNS1BFI9gy+tHIsnegNCn4LnRS4FfLZdxiflRw
8dI6wWYhXqYEYS+RjZB+Hs7xebxwe93pZ1h0hwfCtgvPM4cEuupsXk6lz+wUI/tO
dNGyB1dA5yzPgbka8W9edF5fKIber+/pNcBqbh0Bvs8CrYhmK2qd7s5RYbwcSz4a
r+4nFYosmXHBh/HkOTlKd9jfnefNmWViwnjaPHZidTULgtjnHoxWSiJ/IqPSa4Xm
3UnNI1yjvLnC30nWFyx3fpxUJ8gn/RDZYxvMJTsy0cr8rgunOCg1f7Q7ZsJ5QaEk
JsiM+TqCgLQ/+TtW+ODpndKVxXJHALdxo4XLwGupmWNJdD4Vy+bi/wWmIvSpiAG+
PMjOH17voW89urqcePpxUL+Pq2k5HZIUFQAVXjZRhffbtJ6HDOjF63MmYrDZJdbR
IU5cSpwi8kUNFemXp0XuslHnvQJvzQEbpmD4Yp5SOllB1gKN7vpvLP3F0IMO7ScU
9uh8L4z8zLPMFFnWIeJ34uS4I2O5sK6lTmA8/OV9VwtLQbkD2ErwGEeqwvncC37w
QkqesjcIA5Lq3LYaFOCgGMTtmIhSliB7L5YpqaeQmlWcLbXmnS0IgkOcoaq44mk9
RM4fX1bejkc1t0uQVGr9rrRHgI94APzBkp9Wkkt4PVsjnnGW8q5rrpNwMWir503a
uM/KZl7O0EGOvyFvUFlS5gDnakIdLEnH8sAEqKdTwmucDGkhlQ0t+MLAmW/PpfhH
PiMvaDCvCdvqp/Ce77QtOX3Mj7SzZLZGm8fhojzRIKl8BagvDcE3Avrx72imV4cs
r+w1v0+TEOHndjMgCXYwlHGgzk4vtf2CbS7u7tsjxi6lnBLnqUmTNEivTTq5x6Fd
WTwo8GuvKUnbap8fScbFt1YSEI5Q7UYS/WWczCiAXQPmvcRT104HVJxBQUVoARqO
z2ghzG2cpMPX/uRSt27mWgQ5vBMrSoMmfxs6eVf6RqDko2MRDkdmuKKG9wRQGdat
ruIqiNQPA6CIc0rd/eSJZKEDjIQnN0ZCJm00PpeNMAx6P/2CscWFsn1aJLKc72JW
yQxw7L0U6jgbCbVZmTeY4A/zwgMdjEMoGl2ZZMMchoJLZsLbGLUtEHaTMj2SieZr
EAiwATM8tLLlKnw6s18JkGZkfPBh498wJPjKn/fHotxSv2ea4Fx/UfS77MyuAxZD
1sxjhDPoCQFL14tQsMn4E6e2pnZVMrdf87HWqu+3K18mHU6uY/chQGb7JNkcUbvm
LbbjH1YjOgLj0nmtlFv6CYyvTrvQI/GTS5emdTCUjNwh1OnpFKmTcnpScl17mo3J
DFdVxxRPOA5+y7XLCUTjVzsAD0jmQ+nAYaAGwfU/ogsE+GObk5RF2fs1KDbnDmf4
fe/pIg6Sd33VbX38BOn7fYGBNjxW1dkIgevEaqtUA6VpTBzvDEmK2N64qk8U9+tF
2UZ177QP+u3/6zXb3fHxk5x6kOPV8E1FfYGcHH2/6gfyfxRJz9QdvqJJCAN+ap8H
Ab/3dS+dAPGd0DZWD88KmwVjExDgkEuRiH4BGc88X/Mv+vOa0C77DcHWU2JLxjBB
dJYzBCRshJ8ORNJIvC3ek+dzsUQ+PlfNeyRl4dI9npHsoiPFQNcB3kBMQPfVG5dB
dgkapb4baGvof+Q+sGzqwMLog3PcC8aevinXanqDofuT7tULgZc/2zrAVlzOk7GU
3+9EJu3Ab5y6RD1QKvdGxENlnrqb+5KcLv7MJNPgPkNzSSaPQPgA1reQgOqnxyyt
EkgT5UxqJtGFJ4ak5F0Ki9mxfCs1AFp36D4U8i72EwXUf39YMqlLcKNulDzgZQo/
T44ekolF0usu85dj1NpaLDssNV9ZTTcl1DDL23KQEEVi0YszhyYthso6WezThEXd
EbPwYU50JsKAgHRhAPk14HuDJRvx3xgmaNizw9iyog5s8La9pkFH1qLw8pdv9pCC
V/oPiZ+ciHBI/Tf2cfCm5qSkaiA/dWaHZZdTfKxn+uY/VnuJj4gHZgv6/Uicf00q
wNoCZkUz86JpATen3F1g+US9L/zv772Lcwfzb3foJUdUj0v19vaZJxhc0SfhvbMt
k+ICG5SuU0AQsQ8Fl7Xa5ainG6p+uRCuzhd2XTU65ncRcoV6ukndYSGlYcXq0K8p
V2H8amZmQz163Gj8A1zAMD5uCCjLZhqs4fseqjvrCVJXBgetU+S0vzJ1ujZYcpO5
hOccKpg7IVLFdzrpll6m2gRpe/ZZxXg5A3qXLn6nLF4qi2+KjffSzIdt+y7vr4Yy
qnXxIO1b5Qc0rIqMosqBF/NLc2AybtCqTDjSdWfOqpGUbNmPWSkh2+rqfaWyyt9u
e1g2U6GvZISesMCh/rT7GRhKdr2DHMzdG3X+23cA6qajBWVf2IqXuMFGS29DIyhy
9Ah4XGIfXNKaJBywuOvo0xI2drpyptm67gxfC9vk741qowWzT+yEI7JnCJY+hMtt
H+JcGefD5AS1sDB8hto/QBaNJNwQl8CIEA90MUWMkQDMCg/sNBNwLa5EqyzkKa8m
dnOMLoNSDJy4JEp4YyesrID5IT9BisLwaUj56rNx6lqnC5J08N6RG5hnyathP0f8
U9zve+e47+qJxee9egLAA0PojAXU8N4u3UwJ9syIRwATyCU0NU1aB5OJTRkaWsch
gUetMGd8oWemnW7kUqr1xkNPTNO8WjsGFDNzJrdR4DNfTKBy5JFacUiYDr9UAMZw
uAoeUFhPa3fojptfItyezBJxO6P/k2nAupCJKfHHbaTl4AT9EtZDbzJyPiq7i7PO
4n5mHMrZq1fPgiFoJQi6f+tPa5PSyYFeEkTVq9fGiYfsYqnaEd39P4r1P+tv2d95
a//CA5X1/M7nox6nUFYeM+jOcdel47LDSP73SfZ+OlgbEWh03sBZ8KCsmXoEmTRb
wBaeELI6NTQtt8j0xaAvo0wtKt4+RwJPAQdk0QR7kvdPduMAVIZpd5wmFoQsz/4t
GT9qBy2sW64RqLsXxF4f6oRSeRktS3kSFuylc7RxM40JEkFvKa+W+uPFYUhMhknO
1AbJUWF3gTS5yicG++0VKrZgu0b63dRllE2m4Gn+gxBm8pd01b3SFoVroiy5IncK
N+fhxBknkr0EMv+Gh6vZW67sUpt7RQmMNTcFMJ/tZDNVNaOl0dU/5P98WOoJoSWE
qSkfGn2iEM5f/arOpyDBvVVvHIUnlbEmE4OfhZFjrawQQQ9RsrIa/85wzvN6mDZO
CRZ9DLQ3rhJmHdJ+gXCAUDwSTgw1AMKB2UA+JGruEEaFZO220WeFdp2PGhAZL630
UcqAW4D5HF5Z5iy6oECiji+ZyKQZ13duLyGODbBhQmU2ZVFJypfgI9wjT6x8xpDU
B2M5xeQtbzBhv0qDTVvbNk71ict8bHVppha49hyx6ts9lZeK+/Z0hCW1RfjrRzCy
O8XE4zJMZK600o1/Qo95C52R1ar1YbeDh5BZaLNz4efH36QU149yBDTsuEwqS6Cp
NdEtRE1iL7IxYkTtfNvo9qFLnw7UpRV7ivtb7HmcAcWoI4XKFzi9uDIQN12dxGY2
AbQJ3bweF9iFLTjIlg2OGzYy4edBk7eCxNeIAAfsJLYfeWeJDBBvz/iOhZtL5nk+
MSkQnmSU8pA/pnmc0+WsW9n5kHgyX2dcp6deb+m821PttKHsnmV5jT/9Aab2/WY0
zM87sjRbzRBBLc3ucyqjGaT3Jvh5DXSo2Uz0jKeksqCTPRgxBW6Y+c0D2zLNbWmh
7Xz/FLURc0N0qZAR7ZlxLHhVtp1p2uilM3qwdrPjCxxF2q0cow8GMRxTxYYk92BN
SakraeSRh8cFuXraiMfHzU5LK6rpNb849+cLwyckaqnz06MJIFp793Qx+c/QguLk
jj1zQ3j3NKc9+rm93EYFf67WTPqyL8RRhmj+BFm6aItbLBn2ncZWKfVz8Mh+pUFM
2vdw5TwJmXiykvKovhxt+QcFj3B9ksW6muxN5cQK0KZD7p2vU1pznnWFqwjXX4uz
oS+8BqwIsSlrdWOVQwKMZbQFgztuVcpeDZLrQUc1hkh0DVamqZ7uze6EE11FwYWS
zfd4A6ofGbQkCYSnACze56YL5R02L/tuNCDrkfXLiDPV35/X6nkKk8Ji/7K/qF94
N4PgjOtImqniYUMa23QCymLGLOHiO8Vj2RJ7HXcveAlFzsf9sToS7L1ALs8am+AL
ZpF/C78tg/AWomg+w7diJZww5/7PrXLxHngWhodWw57EF9/e1ztm8ToxyRGO4UXd
faeYCdmVzEwobdjcD+NvN2ckauNohCMXvfRHU+itEqHWB2L/+aUWLmyQ+4ZmqHUj
OCGRhx0u/0ap0XRLHMWx7AtLqKeSZZGF/GNCR7iGaN9i5gYaQCmDntNE/z7cIfdG
1EiKLOuQSceSy81cKFgkL1UJ0RnDR4dYJXSup2dG2OMZaXVeyGRepzC1Bk2XYHl1
CR8XqiU7SZT1IDTORFs+fDkoGYP9Gxw88P66wIgDIVV4oqBpsbUFmkgRGYj+53KD
kZIRd6GkF2XdW7yFt8bNu79BYGoi+K5aiK1W4kFzlnsMs9tJHW6d25rjJSN4scnT
CV7LGbvr6GKgHNjZZ+5ufULi5cYRduWDcun5yfDjwpaYApSLUNiKgl/+gDbX/dc0
c3v2A1iz5bLhZt3IcffUydLq/Fbn3/kL0yxM3Ml2jKrhuh4pRJjHJdCu51BYNJbn
t/gMnEmES+DFVFFnobRuuXYP1kYb2jpVGShFtoPvkT4BNeYv+8u4vn1yzT6J+a2j
wa2XZgjwOZh8e8jFRWeYhQoe84L90QfMNvtvHGrXpJ7V3syBRBnb5EvvSZLp04YM
eourPN5VoRDSmDjXBMEotrtvkgABO2iMO9bJlbLl4WqkZS2nFTtvLr6Ctkm3PUSR
DEFuCMF2joFVHR4bbU/+jaVMW1RlfR7X5hnR1ek37Fqg90QSJ1/5SmYbdagAIboB
n3Cb3NY+RHfnPEacit56wdYdJLNa2yQvXgilEfmVK3M9yPQ1496R5JpAvY5I8ac3
0a2yYEn67ydsaGZhL5YM8rhaToYWvtMMoBMj2rJTcQomF7RLUsvZp7xJcMb406UT
pey8eesoYzIU7HQ6jvs8BotUkizTJwi0DOqBOYTPsColB3AudY/qImMXnsMbSIuQ
isrbO+MOy6F4RMVGLVGd0ltNLxO9fC/txgw7m7/df9I3AbYiR0n6SrBSYI0kdX/x
XUYTQiDU14G/hQqDALZRih70IS39d3LlmWgjsJgpinAu+XxRpwxMJJvD9W9aGQWO
jG9Ap/OkEVjohPuHvF8Hx3ZwnX4dY7O8Inc7zwwtUW0x7osTBXWt0SkHTMgf6kUh
J+tceT1u0kgVLMF42z3uzZEiFJgXZ7kx2qW7gT2estckj1z7kbev4Wt6xmJC8qZs
IkD7veinyRJsg1va+kLon4pflqS8MpICv2CL6XabB+yihWDoC7ZP/71Za4zE32y/
tU0qoYzUXL9/geyOpAiiXU1O4riC2Qm/7JNdkGc0jZ+RywTUJ7MqyYhtogQxVMhU
xhs3wLeswrdMhlPW3KAe8G7wQjiFFHEL975v4NARO5+jy8Z0qLH6uhPJ5daScv4N
51llBEl8IZlbIRiDz6yacKmuhpQ586eC8v8b8W5slurpxmuPd2LM1vM0v8tuLmZq
MdZaJBFyRbj3eDGf+9nyVWxQPt7yUtBzF6F4NZ6pV+NK7UQ27AEdHzyefS8oEkEO
Lo9a0CqIVbuvgGfu6PscLwDRQEAMA4mMpc0OTewMl62M0iO6iq/JY5psXZjEHptp
krAASCnEZiptaO3Em2ruR01QUSSIuMoC+a5UabONk7cSnIy8Ad7MAIc8pzOHtBiG
PFJZgMZsX2Zph82G3pCkaMMyGZAizSFLU8W+k6v6G5gtuvjVVMB2pnG2whONalm2
eGcDWCX+dBfW49qcXccamuGCWl3dlU6yTtCn8KyW0HyhHRS2ZPi6blG8nCJaaVMY
q+Yb2HwPyu97n8EhADh8NcB7mYEAIUHqq9k7k8lGGXIrNTQgPArOHvCrL/MpNocN
H1kA82eh+Zfugy1F8ct37EUNnDsKJNE7HH70p8ujxoLyr4UH0iZEIeIj0V47+++x
JWVIIC4v1sA88/g2NKPqRuw8fNbCoAr/U8GoW0c0qpXtv9e9aL0BWHoyA7+MiIF2
OEbz6k7SZQJSnMtQFYp7jTz1bXcKygGKcQ7uuUx+hxv/lKVZw5X6O92U9AJOzSlr
7SRQoTIryFY4Alwxew4A8jygmCj0SYhyXGWkKgmd+kyUFTad+dR1w/rhGsqh9BZ2
miHWme5Vb+PkeEx8TEN2gdLhTVnVne23y9skRO9RQD1hS2o9EKNfs2zDkDSc3r6v
8ZRzNSjR1zeXIXR1JZSqjSPENY7tqejwufMvAUr0/Yda4XbLM/KLes9g5IvZv++r
DKtrWvN1eMImmYy9PdsrgvcajVK5JcSCl/+3AOvT5IUgcSHuJuLhZCPYUzpKyTpU
zGcxTyeMFDxM+Z9iQECoGve59MwgEj72gLiyidRebRW1gD4DGdsB/Q/SJg9vwHQR
1jDYD0v+8mV61MjrQHd6wQGNd/kPubeYw8C5a1DCgusIWgh0ycOD/s6RXmLKBscj
dqXo9y0xkRbNLvYbZgmHVh+qCbSxvA7ybP7rjha+zIS76nhY/cUHnhDQjPmSQQ2J
UdEBc34MAU4Op3zjfpznk2u6S1MWXfU3OkiNaAhczkpgJH7DnKKDQHNsS7m4n+b7
GD5auKUcNmgC01MR4DbyS8fFCpFejvpbHPWijW0nsuHfw/LoYcX6KiR9WqBm6ziL
qIL5sLmcXinQu7E28+m+P8M+UcMPk8DMGtIvLT/ScAcxsFpSp3YVfzGhgL2SG4+W
7YNC8BuubwIUAsMh7W4vtGLOeeiARwzgQhTxYrK/KkCJ6PaimfdWd0govKfGwGch
lLrh8yoWNBmwCWNQf3U6DTr1+pOHH7nB/xoNh2T+YOSShVsEWkmnDzyoMOJ5J53Y
mm0gsEfBWX0zKzf50WKBvps6v/HWEERx8Eb33T9csg+nfgPuK8wTtPAZJPoYTHJZ
BaHWGdxxvTBhLbYkdtHdUT6wtmxm23YLXbDYXGXttUYNYTFxo31F9MjhM9O+BYJg
+C1GiBUnhUWEBwbCsSA9TbsQBOmoA9a42kouwA2uKJ3WGutN9S4BFGYbnUhGMEtM
0MPDJMufwCiba2gVN6yUVTGe67QEOx0dVuCRVuuHXSTKvZoXZ8G2xYc/GGvkupTJ
ptF4P5aYTvosRraNQFYMc+ZJdYeaZimjoxtEhl7XRUiD7uqTEVNuYBevbB++lxc3
d6/NtWI61nK5v65m+fytTY/mZNJ8MY78tmbuAIoZYf5nd5HOZuy8yHNnZCz5WVWX
Ga4BqJNJFyAdCxe2TKweB6i963obswfEmQQ/mO8p+xyBPiAtXY10Mi+I9BGlul0W
iSrhkcfSXhyL5adyRoNylqLJ6353Hz1PZQZbENb/0Tt/7q3+XPxG74HsGTMl775I
JZqfUa4JTKaJcoUDDvdPIhMLmXVTWDMVqrorWQh5z+f9axmKJdl7z2eW2AkmIzBz
WNMkdrSbk79DG2wCdPar7yJFgC3E+9uTQ1/H/ujTbJkYy8KQ42k8ZKS0aQtyu6lm
rJGpGE+ZMtIeezvBYETeXc0jZYwG9nVPMV3ihpCmsND/PmNjz4kKRGCS0L2Lbm8F
5UVotNc6ROD/lBMC0KCeeMwVYNnqKnf++C00Am8G6GLznuH9icqVnI0wb2yqGLk0
00IwGPc+MHiI11HXGL88+9DyxNGjgwBpeNY/rOnF/HoFwOEP3YS7dacoaMwN7Ob8
tjWSZMBU8tJmOyRgF8ondTBqTWJd/nc8dc/l4QUp4//10V/tg/QIXvcelAlPGVgK
E5/40MC9gG4+KDIvVEqIGwacdEXOKZv8RLl8zMJ6ZJEh2ivU6GAYiKafaC7JsFe8
iG2N00Ehq1HuAStk8guRXoCw3ccAapuHo5JMpiJGcuj7kg5QqN2LqtjfawNwRJtw
yK0wX/5bJdinQRGIV92TfOuezCAZcWErCtZtBZklB+A301jkNdY+q+/PSMSN1cBV
OGzv2QGfRREZE7gUqWsogEUKb4+GLIBPNwGeLL/zp8JWaL+gw5fMSxAeaIDO92eL
wRk7pVbzpgm//f6vgyhteD0SGHvJjJkwwwYIb1aLpdMK5J1A9i9OgY9jOiWDg8Jm
xtH167/68U6PeNGeN4tBkPb75I69xNvJiu7fx/xWOF74II7o64fYiCcDi2uSYTL4
1eYyVNpPO9bMMXhaPPsU6BiuSm1RXaw0k6K9Cdn+VZF4jJz1Gh4LO6h2t2xIqGaa
+cybyMtGn3o3b7MSPMit2DzQWSGZRHUzrvxaFa56MTpkWVXd/UM4/lokpaaBOjnv
kokD6NiJcE+ClzH4tfZKQLDr9cxqCQuK/wePEw1BrFyhrQ+zFxsOqlSKj7jpI2pU
GiFxJrR++hSa0LJUPSUl/8lTVedx1sm6aFIiH9E+ob2bwM5Yclntow3ZC1w4sbrE
nOEI36CUNwNFNHhDksl3mtUUflLSTSmUqYfzX1xYtR3NQ6K3tIJqYErOFa70A7ut
Lu2liaHfYm4n5ovwvb8VpGpRgO9WQzybP3H8LC2KVCCvQEw/kL4xAUYAZBhxzf8B
Vbpu4rZK+PwpOEArbehxL2b7Z7FLNsmqA1ZO0rD8xl6wZDIiYmTZKaMTOGgKK04h
qAs7VWIucP3I38dHv+Y0ybQ6vkIkaxcnpQ2lepKyQHW11CgnchHSUm4SXV+/U4rE
oJKK2pyQDaYFoDgNsHCTWGA3KRwYNu5wz4VhQy5hYlWVMg/9y2quXeEoQKNitLos
czzhM+/EzVZskbp8Ulbb7OMA5Pn9zGbFiRAiiIeqFG9NSpPBgPyBe1+TuQcoX3f1
h79z+pZBXSxyQZnSWaAlejvoiABsKiPvSbmLFtqydp5CC6LQ+GgUTQ54i66DL4x+
r0z947Rq7LqpQK0wi3NJXglHIfbQtMYmyTWMcEL7iL4G9pxo67z585PHgZHpVPD7
mr/gH7TMXdUED4hiC486UfL/e9AAQqSTIGQFSq0MLeusxr6GVPeyPC4oywEjTmF1
F7bx4suZOwDr7DYqQwF8qM5Lm4A93+VeAZ3vJwoy10724omD7VVroykPLoQ7LR52
2ES5v6Fdii2iNSTOpS7J7YeCXyfHZKtbIsm7tWTmbk9Se/9W3sO60dPxKK18dKm+
PO2IlgaqzDkOGdRd/bOSEYqhQxPxcJgQm6zZl0huQGw/QWjEQFu+AFAxvMhgFxxd
GQmDBtkH14m6WVyNEIc4BELOybw0KqrC+dsM78XRcJHfblXQLr/v9Zf+E1x4NSXx
0n9Y9qlLdxIPpE9W8+EXfL0ta7UHJxw4ytkIZ5iHyk2DGj+jaC0WvqYIXtmMhPSy
oDtbv8Bdh2MJcBTSK/fHAJuWjpHlXQ/bXB0g6frmETgbxAFAnzBsx5gz+soDDPhh
jUsEADLG/mqteO4UCn/k5EB5+oGz7dlhnwruL7adUbFhjmpEptreJjyJG+nvK930
JefnkBKw7A80SW1oSLafpftEBs4eVots1E72prtotkR9da7EKD1pPakRpOamHKnu
oTy6PzjGYNFGtRbYSjYR3EBVKkoRsYmQjpJ55X991Jz0r0zblopxc5Ynt4nxg2kL
MezPOfwU/z0lp7B+ngzxX7Z6RxIeuSdP6yfUWCqusQ0Iq+O2s9Fu4sl+h0nlTzQP
2keLi8eaxdrN4KXJsUtLG2usas1VxFRDMUQsKLm2fp2EgXPOB3rLU6Zd27LJSa3F
W42Hzh1JA+EkzwNU36PM7gAfJPNGFyHiEI2ZjJys16MeQJtgmp5WZV/QVl4c8kSY
4VdllQPpw9msjf10M71790yWx7JGwoHJ+Lq33C37JxqWLt0bbRxTweA/4Lu5Sbyv
+NOAyagQhWqQGO8XDyZXXGy8WuqoUykOs23GAdK37ijAfbKaGQrSSKlArcylr+Cm
GXZj51ngelGnafiiQk4SLCmR558j60duvtSjQCLN9k71vi95+19Efo4ZI1wQkHhJ
H3HxBxExw/IwAklyfIMaDmU/7/xpavJ+ygat36ixBcc2+auBTCg8jvrMpLPRQAzU
LPQsMue3HzTSrF+g9EpLm2X6TjWTL1TTQJ2K3EmZ5iCNInS9pU5PrK4jZz1EeSte
+eHr9SoUO2e6fc0HxeC6rvrXSrQC/D0yCRL1eR52LEUPWIRoaa64p1vHv9iIfAsP
kmvteUV1YoixM2vLE3MNViG4jXU1dAVvjM6CMGsbUVlMSFM3GwFa/5VUW5bSV4Vn
/T07pOaGjvNoGXcV//14Gu1nX/9g4JgExPSjcvSHBoEcAyt663n3O6dCcvSqzJ11
vUjtUF3z9CMteqKxaV9a+V8suM1SlHUXAeh0pkuo4BgVtbEtP8Fyw3tw/eyGfu6g
rZd19RzEhUgO9nuisDZ0qultoClHMCcCP7eCMrBZDbCqdhWpqPnEm0q6uBVect+Z
v6RKxQtJmk+7xgMkD//KWwy4hHHcv1PSyx9sQEjZKq/A0+PSTmul/0x+36XS2Mwl
wOy/Zy7nn4f0opMt478w/usFvz75z+uj3npLx+xJ+FvphRh1cpVvnqTy58+kJtSh
aq+XkHAjyqaCxaEZQtoVhCFz8BZ3WYGpYcjTltJIIW9azomIsGCJnx4S1uz5H1XK
yJuADQo2resY1VlIEGCHNOCz67FYo8UKMumAkAX5NNQy1r5RRu6DgYDmXtV7ki/3
+G4Yldl49jOUN+1mqDD4zbEhsbnakO4AdUbgxADyXLMXWVogLVfdxKaTgf0kuZCa
Lzgowmaxpi/7u0QbV/p1YJy4XlRvNFnTrO/quK9EVs4MwXmvnxsl2qsFtwkoycef
xm1AY5YfJPqXdmAqL8ohjkexMXxK0sRocHa8T9MCrI10Trvs3p0fSmGwggGralgv
rXzU9V3O7Pgmd3ohwY5SlYQYe+T/MjNtNLVZ8YSzNtDqd0ZsKYvOalddL5+aofV2
3Hv4o6b5IuLyjbZn8ZaGdF3jVVS05zAceDU4h82KfWq4U8Rjoed7BGxoGNp/lg5Q
ZkUerccuWYyzdzdIROM8TU0h48ZZqP+uWNclZwOglOC4Zbh7FsCb9TXbM1sl4Arr
qfrhCmh6JCCNhTEfGitEiuInZeQO/DG27LRYpVPPssvoEcc+T6D3b0QVdDl7eBg9
bUE3G4gViv+kp1bcAfhvYSbIRzejw7Xkx0ctRRloSlvjSPW3R6b70qgSVTuyUo85
eFsGmJ6f9/DK1fApBUuZwxEVF7BmTcZdnXapVoHc3lFfwuUluRcrS9FQFOuzmbUo
0JyX2TUr/DNBl5L42GcSNzlBB1CEgG0WCClJ2OKXTCgOXu4xeuymwYYSOgIvtn72
ZhLK0yUsbnTjIquEfrHgYc5GMplZu2PX3tqf4ADbtz0iFA/7tWONlTNhUij+6GcI
QL3lN2cR/+qC7KijwYq3sN+kVcNNluldO0HAx4SZOznUuSLgLxCqw4R6/DP5R69L
0TnQEJROo23LY4/0N0dBg5XBd5a8sA2Umio2gof4MVmm7uyOXproqp0XITCZzDP2
554PschfQwb8d+Bg1tS4es8k0QonwPIksAxFFYdtrB3pqMhhxdZsQqpeKlpiR5Bv
7ovDnd76R6NuPM27M8O2Ss378PZ/ZoSkSgESKjeFgimlFzcjcxxobvz37BATZX3T
XFTtLEnICC8YeDPPzPStebLyeOelRnX/VICTkmLlkRXb9NELelt+5kKzCTa4wyfx
3a5RUEZStZDkzjp5dAD2xp3GPOMNxSzWYW3FWj/jbHktkztQBukXMWaWK6N8BZJa
KyOspNKDVPTDwAZG70CZSKnVNvB/IHAVG6wo5CDv3d7ZQNHpVgJwfOZXbRakmvoj
1DSy9OGa2Lixb2HLflch0FdHGev4Je8qd2q0gdJXTbegBlpImKnZRn+x0n2cXuYI
cGdi0doyUVZT/Bowax/0PHLpRu2Vv4e0MPs208VRa5KS4zqmVXL5TCTPlN5OnnwD
1BJXdjtcUG1MKaoZMtF5purNZwSmLai9hxA8XdHchCH3pPwG28IdsutfOPzb3EFs
nrftartzkQs2in1mgbV/FYALeftKHSVruH89rShlKPcWSVJy/fudUwojP4DulPEQ
WweM3jpXTky2+lGoylue/jpEcBjFJ+fIww6uQBg4l4vBo+835E9b2BrAmUljD/VH
bUM1B+6M8/V9dkVJ5/6ZBSRgMR1x+uicbG0CN/qUpi/eBZoEi7ma+1zOdBTj4pUP
9722e+CrBALh3crmc2Y35JjF6Tn0ZMS500ob4TRHhgBWv/AgoeZSdaFd121qq/GF
qlKk8mY++ypFNbOj/v/Vq7iGxH+5MuUY2wW0HsTHqbp4rIoiJSms47sTIbfPnhOR
ypeyul6WF99hAivAfBshLY7HVX4wt9HNnToOj+BXCp43kbgl3fWY2TUvKPpYg/rq
YZ12wMeMX9LjXWBPM61B5tKsuZQcULav3hqeWPXruSLYyRRy1nO4FIq2jL/8G9T3
gjjB+bHwrTryS+yHVQrUolXIuq9wyJ7so/9DBzyP+4uzGzkAKPhkeAd1jvs+yXzR
dOWs6KrLYYBGFWaC2LAk21g0F8hpv25CJgWW6MQn91PkjVkiAR2PF/k+kfOgUfmL
nzkyk04BszeQ6Ao+fLLnW+xP2wIgY6EXYHvlz62BXKZNQ/ytQi+iAGs0Zwg0mgPm
b3rcuS8zeTj63NBYcc8NFNen2d4cjb/XGVbHjGf4BAOIeVTzIHKau6qgEN4icH16
x7EBrgIxMfgcT7xmi4yJH1IOQECWe5KHiZU5ATaStohZbbRXCVb/dNGklBdzFYqH
8VYMbD07b+vUyp4lkTwdLv40Z4ndx7F23v8C8MIk6NbDkWPoJNRklS6pHQQhggPr
9ZrBsOF9VrfB9BF24qkBpGqDHc7nm4WNer5Bf3NZzV/3l6jNSR73/rpNhuRuwMjM
3Bxq657Hf0CyvTyRCXqHS61u7WdSJ3AGiWG4Px4qsFUNr7AxgRMVrhh7r9q4wttX
lUd6jtDNrNaU+69EeiPLVW0XiDpgliDP6sK2puf24S8GpAEKWCbZs/9xLs4ovajC
rnqaNb7gECoVfG3qKcT6iDelWiRrLfLLfTpvqCtR+64NXs2k5KVSxi5y420K048U
3T/XcFBMfSFVTvypx+64WUyoHzLfgtXC2GOQCmsFPg2qw4CGhfxbTNfb6mvwK4EG
+exIlHncAKYwv+AWQgjqrSny0N0OZWQG1qk0ks38YQLlhBS7bylknT39K4YApoUZ
A9UBRk1VgddG9WbvUBLLGCD4qQHlIKVrQr+d/3rb7i3zkWC4qRjquijxXuCpszwF
5mQ1/Zsv1PfwefJ10sexiPUhe0xsjEYmtZl8Ya6Q6UB2RJbJ96z53iIDMIIMk9Eh
OKAB9Rv4dUUWK+fW0X1Nqgg/EMC/0DUcW8OPH/P7Sm2bIQOi/gMA81wvyxRKeTEx
8I/EqR4UJ7PL7tPAXsjp9fG8RghtFyNdiMq1HFzygbCilytBLBD6WkmHS/w1tPQn
5ESZ+zg7wz6UU+MW4hokuQd3DLctRuk4/3XOLzx2bYeSGLzfDjMV5rh5754vl1a1
ghVUyLa6eoSCk5D1dLFCe7OVsV8ccbceKXcQqWg/6SPm4OL4M8p5VwBNeIJkQ5sU
YK/3cKMJJqWkzNshWTIPpatMosptpagzNkMr+mMbyuj0LKL0/6MVdkoY73cfGQHE
e8cRuNTfFFlh9rxCEYviojGOT85irU5/wpQGwnvFgKUziZowitlbZaq/6iaoijOz
lyn/Pj4BVT3QOLkyDX41HQIxn04OFwCP1548jWE+tPurta/cCYpPrz3uVs1eSw43
/wcKCAsv936XVgSRlC4sqp11IhLz/4glBgMi/q6iW4/eYZJj+nFV8+youf4ItvuX
O8r2hFcbm/p5SLtqcJKGbYR2MH1AE810pjMLEL0PGclrd37RbK2HQCVvy6Jp0hFs
zqhbDdsKLS1lE6GxydZ9L08tqZmHdWo8L6qqykqHeaEZOHPtoFmlcseFA6ndTIdl
uzADUDdXqO96JIBfmv3l3OxUbos5+pQBo9l1y6zmqwBldjGU1RaUh69qrOl1XTrT
wEhclq3E+Z5/YemCBSeG3oOrl5px3vQdsZ71g4lu5KkSlSiKzfvs65YH7SifxGEe
yfviBWtkh51Gf5BTaPUNGpeyoHzGEUbuhQRZELDl720VmTctRxs2TzqGXVINyNPn
OzTSfhAuyfB4b0E22yfSYXtkYIZN/19k5GUnXtEnFMY5+SBYO+YeZytzVNhUUjbR
EqyQHpl+jRsURKmcZT+uUjcDFnZEk1rWn+LEOZSXfXizTP5lvvXBgJZvxeskSpZj
JfbffddrHx/kbrynJJ2ilV+HDvMZDK2Tgg28GvaUGsCAPkK6AuaItESrGcqWpvOK
VdNhdeQ26jONZ3Q9VaqklBj0zdCX/Ue1osg1tIY6jkxgIc7KRvz8UNdHZ9QbWZhu
RF33r4pb1cX5zT8Yjl7VIxsrZEEVaEUrztRUzeXbYN7qdZfT20K+YDSUj+6Sqot0
rjev4gXi3oPTLVsjNOTWhVyBonfSHtNTh08J82cX65qCC/EFsO0Ts6hQPIQX3sb2
6bpfIgwgA2rydcUbtjty/8OQcQ95AFB+rJFsP40flX2Cvx/gcyJ2CA7Tp23plRNV
Q+VUG4tIeLVP2ZoeE/pL1mpns+1xZHh/m1/BA8uiAJqPHPR16C2pyi+czYJjEJPm
RT8LUdHq8/eGKGdYpEMr9Wt5hxcKeFnE354dSCqBZFW6vMa0Hf2v1ylz9mTLll78
c0aL/RI9C2jsEMjR6sa4huxzUzruHvYpSdHxbVLklOcMIH1Om6KO6ycvDc3YFl/9
ubGlyhJFLyM9WrA+CAXZOMx2lU4A/cUvTSa+GjGfHvZ7Z65+mLnqamkOVsnGkweQ
az1Huzt/YAHWI0fwqC54xPGN3wAzZY8B1jGVcyE0I4xOlVMhrN7nunAJQuw7qOnx
PxdN/xbf4Ao0BahQsER/z4kP09o2U4CVvq6LMYqIZrdKH54hFj319v+Uoexb77Fr
40DHIQq1Ii3HzsTc/xeIzQhturopkoeN+iBNK1P2+a+pJ2I7vHeIQq2yH3PbOoWL
E6fJLzysyEYo6JAo9YKpi2WJ/URVIwIHb6bY/5DIZS+rfBs966tGxYksOKGueSKI
4oi/uiIRAp4C8rbz7ou+Uj0IKDnKcK0pVMmr7ZNwjd7iEo/fFSKcQD0ioyv/nou3
E6KgNk1VIOzbDeFRo0B/bGXL0FQ693kAXUuLAa/q10didCXyyHVkQNt6yTu68wvd
c5QT6532yRO/jGvmzZ2N3kzjY30glOShS8gxOkq2mGRoTRKgxfcbGXHrued71VDM
xz3gzxLNVzq0T82YkKCXsbmWHyrQOBxo5pglNe+corESpeSqXldYmDVp9O9sptW3
tQLv5aSvq0Nj0VBxSGIoIumS/5GGH4CLqiJYhYPonpSH6ZIoB2wz+A8bww89cMc7
0vfiTv1smR8tfs7lAzAJltsG+HN/SWKfeRLgfhGy2LnuSJ56bCjiDelW5tkhLlF9
b40jBylk4tgF+jA2obJZ1BknGT/3qVDQsIbYUJiVCe5vUPdB8ruEnmKtJHRrSvYX
4Kq6bOhjRcifA3f8yCNu1LboC5IKyw2rsgZOUpIIyG6Cx0YE/tcrpHj3wNRkMnfb
XOkj/XwEoFlnzabvCmyz538N+vLXlSwiRUFcZHC3ABO0eZORHTYH7ujLxVJOSwO7
StuPhnOU0MmHKEraxKCobtYIn1lecFn8pm/TJyH/vmQTXjhbvjaNYskRHFeag3qd
/hTaru6WSbxBLsgewigJEZvNfRdfNoil3WpUFNdUB96pakOEFC/yuUqcBYhSKabe
cAOVYFoe5A45qA223Zm4NvLaV6mwLWsZq5axJ+gZoRAEgvP7lblv2zfSWrdZ7cZz
Up8HHzk6m9fM+SoM8EDP0cyZPdFKvPR76lUKpo/d7Iyk+WivTO4BSWm/937xIBHa
HrU3APSSeYAIQoHHra3UAxTbIsc0MQNvsa4qKecTk4uViryRpHklTlJONc6/O2el
FzGRO+fuaDzp2RvQJYtzF2GePKiMsMvEAC++r1YqLATaTR7ohsLvdL66YAHI5FJf
YVSMxu54dQq1p0U1W/hz+ufE71PbDjtrPNnMHxVLCvNL1BlxjuRdTwXfZDC87deW
5YlGvRwTRBkEoycpoS463dqjm4VrXLqzX8qhpMA/nhVIW1SzxOkjesKp+vaeWidt
mdzlUaqQkFERRtxe71yzN/rKRkjhQPTst+aSQKIGt2EYt9p3gYoFnmjE9+xyJMTj
AIqv3fgXZnJ1YmxYO5IvNEFjEgnitPGGlp05Im/tse2lx530VBEmx7v8t4S6lfHh
0Ecz/ArMEoaANArYiSBUockV8PWnJngXo/GPPk+llt5zdf1Z3uMxTjilCpKmQKO7
Kd1wSK79CcadREMXTvzB7PitS7g3CPA6ZumXIdmmU4Usig3k4WncXwvGYZbMl11u
Jykhtah+b9MAJffszXTVPqV8Q8q0cT8uthaI+ID0XPUsfKAASYr3ZmCbD9Y8I6wb
EX8Mjl2gqdGwFGYKe/PKJJNoLk2rCxDathKb4bo8UUYLk04rVSA0jg7L1gT+o8Dt
NlG3NBfS31NkleAgeROPfstgxkZ/gr0z8fG6RqpFETZ2+HycaI+D+ysSfgtXVNpc
4sy0Wje5MYfmooEhtaieEH13XRdQERIyT5Z9RtT/LuWNE2RncHGTqXX83qM0bwJb
7QU5xyrm59qd73GifUXSE9Oz2FG+hEYBMhXSmZu59X2VV5PO/cRo3isX+0IMVXj1
S9r9cEBFZ19svmL51Te81mp1jozlXVIkc+uT+tB++wkj0jpPSoId0Vx0CnrEARo/
f9NqOXvGl7uvr5Cm3HfNdR4ax3wnvwYjs5OWB0m0mGnTA2XbhGcpkRQbI3UvWeJj
RDZ5t+oAitL3flya871lrjzlzvVtSXqeK5Vzn+8ljeOJX/nfM3PnR+kVswPyy9AB
bN2hIk6n7DeSo/9rF95KXNh3585YcGV6rUY+F5DrSHH3/mSjdxlPf/CgBh2shbjN
MXRZLXJNbLOvE5QSLHpwQNByIA2VRr6J+ItlUkGvIKIFMwnmwJoLh1VjfwowuB1w
duWNCGWw5Yx3hvPPDjNC5tCJHFaKBI14AbUrsW0GVdclo4w2CEhG2B4COm/3N4fi
6zvTr/fQOG5TWsCG1T0QWu8J/Ql8N5uwvVYYeS1EZWmPe+Q2bpZEKF9i/cUYDEgp
oOaPjBbOiJZhIktYN0vy+ooH8npUVeFsSBXbDAl64LmBw2ptnVwL8HDpCv2oiE85
qNKGUrPj1Lu0xB7zUcDsXDTUPmM//6Z87EbA2A/XbeFBVShUTSXG397T7IRgOKMB
OloqnMN9LI1Y1A0xrI+cI4z26o7sbUKf6FRARIM48XOxxN5Ej+7xNGREviC/eVZc
WUdpi0nny3/RZ3MqMl1LnRzUujd/OStJwxYkF02F7Y3ha24XrjOI8LzTfY7xMefq
JAZDEwZxQ0e+jZtmR25B76gSxgcD3jJ+k9k4zw9eUXPl1K7ZjwMWWQYpTiFTPFiz
Pmz0sbb9sF/1BU+J6nikX+rSMJI3b83H6C/qQ/Kj7loFNg3r5Iz9Ok7xyBIyHkQ9
RVKCcbZfs4MqaJZGTvoo2cJ3aslWHDAXdhZWegFfWWCSeFIUBT3eGKR+AC4EMqyw
1ReUqGUTktlhKydHdo/p4XDgp2wdRXW5beI6Mz4W7SUp6KF1gsYE8ZVrNrXEWFqo
w435fMtIXpdcfRQadF7kvtY01Bv8RFZtfuLWnyQ2KS/cwXffwzkh5jPrUGtIX/YL
NVRmYPBVxyZ4LBL5rLXLF8/5GfUXUDnXi82QwPVW8CrUTymf/Kk3nofMIp2SXjWS
dJx5f5wAA7+lb75G4rdESX+Agt+aYM3CjQBdeM3vBD0HfUTEuUjX0l1PPww36MSZ
QCcF1EihmstjRRhiRk0sw28tfHLfJTW3T1+pt//bEV2mO6TyHFIQMeTsh3I8uH6t
ZqRyZ4J1FG1lySl7sg7GWO7043wxQI+AgM5dP5oRWJgM+owLjEnDHBLiS61vFidh
XCQ1/glGsF1tpjl6jqZJc/DSl7T6V2NBt5DAEunS8l810aAeFB8viKX5RRVmQFO+
LHGqo2QL2fisz9MZDOnUCtxpDLD4AT+wyFWq1XTCEkRO2d+abDOGwrggnCnPGL24
k7KJKbDjBh/UtK8RnMq4UbRWQjMRSbjBdndlyGt9uhC2hi/XgUPINyE6sqDaoI8r
obamgG2oHR6OCebKzYAguFWzQ5le0XGBkIUOJpiFTaHEodZXygnZY/WnP+A7HJP/
qmnIfKun8LLF5IdGM430uYuOeDw8iOx5SlMHPfpWSdB43ZGU5ETo25WL3vxx+3xw
6/rJZimBKxcMREkfFufNKayr6zJA5S0X9cUWGgOG3oFPmL4IgnDG8+SW/hlkkYND
2n1JvaeV0Rrupyg9X/M1uJ96CsH+B6kgyqDROsbd9wSw9go0PQE/7PzrW3aaR1E9
V9BCiR3l+gfaatAU6iQ7H3+VMCwvmwv5zBRbnuW+7V8iLdXLD+jttTIGglQ5TJ3S
OnZlzCIc9MJEg31WRN9hurHVu1+GvqUfccuvT0ZsQI4iWU8XU5+ukEuc414k2vxl
0qSUhR/L8sFlUVLnQ0IM3TQgl1F1cYpnuRX6qmt3G9wfgyn8qVrKViAAuOV5FjMg
t/G89SIYN6ZNRMUruXX31DKpxEWYYigeYE8sVVb/yQpLauHbI1XrQhVfX5qDYnWI
vhP6ifl5HWzocAdKEkOkUus1Iij4C48Gn+kcxVdvehrRyflhLhHVFH8lME9C50ZO
rPgC3ICTS8R6wlxEc0DkwIudXGHRBZF0FWU73JBBFk9xPQ/bKgEv6Oj3o+9T+g7k
JJ5ytET8HLdIlZyDR+Xfs9+g5MrQnnhGKPP7yfc+osCwgh5HGxNi51+y53jaPCuQ
p5q9fR7TYi1U4/+Y6PsCr4KwcY2ypYfm0iNFMs0aZ9UCbNzjZWPcSn5kXllqsoUU
Cor8F8xjFVwQJk5dxb4i0USDg8OSSmJjXK5Rg0BK8l4yz1yoNXOzemnITlXuOfxg
pFGidRhM7p4C5E/6J4O/AB+LssFb5oku7DpLaKPxhutpp4ZdgDp/HXcLrmLoCjy5
iy3I93TdCnBMIkxYp4yqq5oAUhOvQ2ijLbsK14ztH7MaHHZvzOkhmWLhDvBwTP3J
Nd7ort7APiwaGz/NYnYGbLX4czQAMqL1GBoV1xmAX3NmVGwowbg9fzcpygcONF3n
/PieucO6CfN9A1PJD2U7jgZqjBIlrI0xBNnauC7bVKatRN9TtZVVtBRirA2DCw5o
7ngqOx5N7ZI+IeJbmKqrD04VEHvDUCbwIPJyuMIZ5JUFd61WYywZQV3ZunSglK6j
CCfKmzIIZhBEK6nVUye4j/1C5WqRAkz9Dl4FtcdREq4rEE85PCPgZmapbWOodxeT
M9ToMP64TPHv+9zpL/FiyK3Nc+I15dExkvnaOGCORTzvi6OA2a7dbnDhGxUkP8XT
ch4ycbZn3R7CrPZLrJncDmuJbEY1SkEBpi5a1WDIiu1x4YTAhgdfYQ0Db9clvBpj
thSBWQnZqhuPXz/U2S+2cZVJd+FEonOYiMiDvpOCJ2koOn/O+qT0x0NkpfYiPMmB
7UXuy7fxamjDWG91H+V0oQ85IEgVIOwtW+xhGQtNYYr/bC3wjwbecl6S4uB3iTzF
aJk0sHj8pVPZzx4w6F0iSeiql8PsFU78ANYibLYiHLK8yjL20obxVEi9IcwY0KpX
G5lzhser/L4yXFXuQ9iRSuy+fFvYFQgVeS1kzidF+on26KUf5UjgDaQTLkKYMejX
fMCPjeyq0tSD2LEKxq526tQ0zulxDNEZZDzOGCHMGccBsOsccdEmXGtwUdX1I4Qn
ZhMzp+2EK9HVXheYTZ/48VC4mTHMbFnB/4aF/Wo+GH20RV2LPSO8pIR1iOcJ2KcC
nTkp8mJv7ccH1qptmALyMrnZmDEyXGjnJ8YzYJE7YJIRRsuelqQjSA1EH/lb+snU
DjNYbpOoWsiOeVCMhNJHNh9gb83fT89pEmGvxYeAj2t96CHCuQnwubCjMZ/6vCaM
OJNfkS8jUFtn1QI6nM8K8hZlX8riF8MFY2ExvUBuGJC4hpk1VcEAQdi7OmgIVYhq
2KsTSoetlYPw76f87ga9yeMhefXDO5vHm+TYdbH3xmFT5rUTMXKmxiis0qjoNpcy
a3hZWzCLNCLbuCNlAp8Y0YfLogQsnxLJf7xP2H8SnW85lGJiqp984rpcuzxBq8gf
EzGdk0Ij38c6aFPdvYj4okru/tTnHMkHgDWl6wZ9FPL+fF1M2aju+4T4XNNcpCEb
ZDJKlsduwqkvnGBKuUTNsFFhn08Ts4MuB3fH6hv/hjCCJG2yMx92NnXD6V6tyRox
a9TDxpLioW7dfh5E1UkZjzwTFQUrKvknw1U8w8aNB0dWRl5mVPNVQhpDHAoChjYO
QTAHRooCvnG0UAJQDoV2W+F5910J48VFE1yIrYtx57Tkv9s18n4VmUHD/ud9vjEE
J8Y4WrMgvaT2zsXA4D2Sf7g0h0Awh1YLe1OEOE1bfIzuRvYsfS2LIb5C0pn8CHZE
fYyh9PScErDUGsmg4MedIFqD2ygIu79ZqUrovWVMc/af4pnmvVH3e6Q2hGVRYOFM
wQeYU0l7wyKG5giZZU4ogxqkaGpd0CftByXPr+y6Icyie1K6yWndstF4dSiA0H/9
wfwjWQOPrKXnSZ+Qc/AIt6mcfGRgclDDPZgmcA93KD4Z6DhsXq+OUTVwbEAXfcdN
8mXCyCR9dnDm5IYWAV68HzbxL8m59qVUBoWZ2BNe8zfRmkHlAqKUG0J/4Lif6Ytw
NrciJkB+C/18BD14Nu2X8E5qMQWX+NASdil9XcrGoH2D/U5ADCeCqqNKprChy+kF
eiFsaQZ71ev5+jsrhFcMerpRA2uZaEJ6SaQkZ0xt0HlIU8ofKrRMzk2k64qY+RId
EOVEVYIxE/xiyfOR+euGnBsISmLVhEQWK76hdFnEXibRQFqNuhnrTL+3owk2QVh9
HohzsLjUSY6bW0BwyXmToU2Xw1cHEWnEsoBk37+C8BPlCTwtR1JthpjavFaAFU69
3RMGa+b1AbXsugKqaFK0vi/f/Ek9igP5b1UV5jYz4Pi7eJcpmjFkodOcAx4PtQFa
T6It4TSJV7dZziwpXVmYCpfVX/L3WcIbhb14Ggzbw5Y4Du6tiqJa2i9yFl71CRxb
Gu9YaLrNy5mgTWAwXlUq8bwzWZjvGIYouD7ePSQyv1pgQRg/en9MIDwnu7DQ9qud
ReFtCp5Kv7DeL7bwpF0N0aQpmFVzVvLpUaZcZv4V9aB7/ONPmfy0SvcCBn/+dW0G
SIOh21TY8rzSPsk8JdKZB+GatLsMEk7aQyG3OBc0drazRnroBghdC8YzloxfIzQo
5u4B9l1NDvoilBRUrJ4ggJue46Uo+qDVgjLJJ7rAGKGbMzUZOu+p78NhgCIINoSP
uHa/UpaeLAjGSyd/D3svAHE0eprrcZ35dzsvWoCFiSnY/EZJZpEp4o257C+KrNcc
In351onHVkfmd2Oa80snUZh8RM1OzGrsH4qszLKUAzPasji8tJpxx2LMIdiOJVtO
zG6/PWxDqHvXXm1hIoqcAoCi4iUujQzaArxU0RaCfFjf8EkrwsHyGJ+KsnU+DAyu
BLzJf2OIkqsvj6o2DZYA/oaSG6nbezsa4rdhcVC0k2PBneL6JzMAofSfFsNuWhHl
yjX5NdjsCszkXOZP8dVOG/YKAUyCOo2ZmoEZ1qJlevIcV+x5Lc/uNS0bfdG8d3EZ
N8hNjxsORGnMmiP2ONq5bWpUCoP7ehN6H1pVlzHeOmmXB+66/c8gDWBchgnCTLNY
Lcy2JX/d54apeRNvlH3extWE8S9Bb4QLhM1+Fl2mW4nVXrCKNOC7sF6UKssmaYT6
d3YDRjk751bIpCenaJREy9CPMCnfzhjOGeHLX7wyHF+grAeExnUOxEu4aFLm4/L1
dbStQKM6LaYDN+WtyDDDyZwjyHZI/Gwp+Q7hT0N4xl3qsQ/+IBBDWOIrdBhVQbGn
gCWrxfRvqE9p0R93CybKMJGds6np3mktW5H2CWs/CKw8jvLDH02RQ+8J/26g6OtE
9fwhTIbl42pRqkQwH5TinceXzZpggm4Fwj0tPWTT/KZgMemhsAzNK5nbmCvpOl+V
MoHUDHQf5p5yB6zbn+QM24j1kk6GGNeSgJZLAygAfdEkwQy6VyA5QeJLAyEG70h7
JLtSek+bN6QUn0UFlD1LwDaBRLVkrfkimilmJcBIb3a6hZRHTTFh4JKlr7dPf6hE
k7dyAMdZdzwCEPXXxqaKYa9PtZy5J34VZN2bfqv07qAwpbaz3XQrqqVtPsK3F49L
+279GcJV0a7NnbNM5csYuNut0ljvD1nOThDbbii63XnmdFNuJD2FBrdVrIxJM04I
+sbGloSKSkpRaRU7yhNxjbeex4et7tnanMsK/O7rr+4DeA21+52ZDPk8d23Hb6aj
s8AGwIIH9RO6DNajNl5RTHYwD8N5g3nP1YMWVCnG/jaQhi7QLw54fUWy9h+HKjAI
fTYm1m+mRfaDBY3fM5LRyvNKBiU2MtML6Bvgi0j35O2XUakeQo2gRd07l+23u+Yn
QED58GLSFyeLzkWrBMfgGQeAqybaTeb8XDU4vsF8T98ToyUMMK/MzSUKl5BJADbe
5QiMceQXUJ8VNMpLXI9F4gvDL77ltDDrTWLmHJE6uBd9HlrIb8poUeZhaJUu6pt7
fCV/CEnz7N4f6nOgbq7gbt7UW0bW+sePvymK7CAQWymsH+HPFvwow6Xjf3zRaniv
+pl1c5AYb090JGGvYMsm23EkddHxTB9wCERfk9k3mmuKbjNA578sOIE1lq37Ckmh
vmJVqW2q6aHPBn6ObVBDxVknNLgh3qoFOT2III/Yv9Ao6HEOM8ZfzROey1oBm2K2
iGvHplrTT6E7N29N0PushFZNtMxeB9pMw79caKAEJvmwUKi/tPZWQtEd5RiLZndu
IIFEEAaiA0/kwCaKC9IgGb7gDy3onj1H+/AN51Kve2UtpvKU2bw3KHm4Xr6Jl88O
EboY5rC/Grs0cyZllPaXj5Sx3LFv3j3M0Ob0LmDQLyDXruinmzhFNbCJzWe65f1v
/2/Som9MJZkVETUMO4tFoD2D51pFDGX0l2djCrdGKlkB2YPgijVjrycsYwnimUmq
OXxzh5MeOpXnU4uSOx632oOQKzrQbgYoexplnP7FS78UFXrrSbqAoc/Ryu61Sn7t
fEETZ/Jz5QZq9QgVdfXYG8Vn1kbL4EbaZWwN6PjhgBOvXbbCZ9YdIDefMYsDPl0/
hz3eqXQkTw/6MW/fuieBPz0D4apcs2zO5d7TcffmZKwjI+FTBF4GJwO6B3TTA9Hz
DJ49TbmJw0qlSoP374ZGWvq8z6BzuC4EpzZMMpgpsgeanrhculmKH6gq8/eVtBY8
/URYg6VknDYHz5UHXoTsN7DxXbXC3aGAST5YmNfznCOYYAdB9n9M4q4C3hdgIXTv
U76hWxaPGJnO+TWFMNCMeTcIGiCmIiOfCQPnfA9+incXNPk3V89So7N+M9Hf5+jU
9DBU87fqmufuJXv/qs52Iius428JifUnn/2OqYKAP++Uxt/lcJ0Qzvnwnb7fVGFV
cllMZVXOd/kUXtmmJq66zvkD/rhey3eyoEJvDgBsifSOsl/wN7p/4rTXLdjWufaV
AyBFD+YoNGgtkQ+TcdqUGPRmdUO63iYhRfE7EMeD2W/pmtE8ydfzSQjj0jz5ZBuw
XQ5/dFqB0k9zCFY54V6cMT5y24+5BbtnBWeOiWpPFebPiCsDpJWJyefXm9zCq3Hq
pVlVyELPC1htQmkdTCHoCC18F4CMmxJZQOqEMQS2hZX3sSe7dUA8W4knIeHJqd+v
MQlgjuT4IXyxqsEHatVTIjbTZafdNnYy1OuTHoVmkCs2fb7pYhxD6ERpnzOPeT5S
wL6OPeOJyuv3VYoix2Cr0omLpGwsyhJy/ua70xRdaO6g939gxGGAGUfk2x8Fnpxk
cvx5vBU/tEnbdfeS5VRolaEzWCulqW2dXuBnuDTTALwYovzzsj/ybDphX61vJB4v
ZwvPH5yAJyAjdEt38vlS4VAhKjGS0p3mpHYy6CIWI3eUcpdFusJPP/N3BZZRjuG8
KnHzTj7JGd5anjuuAT45gpItXEOUq8hS9YUDLlm8YrtnPTm9ElEeHB3VVNlmDWV0
cgSqQQ/SVFwDzdQRrUxAMeXGZy/Mb6DkQIGnlGLV+JXfQrPv/tO4LSUyuiqvDlvY
pnrN81d885vT/czOVHn6H2KrX7oR9iXaLo8z4gcQUOHzd1p1UDDnSb5zN1R3SXei
Z+gXkOVOoc7x27pJCINlMHOjtAyMB/ABeuo9v9UTCGg1XQ6QGAFFs3R/QHFNyBF8
0kx/KIxjO/ANSR5Zf3X9YXcroyoOC8jqX7d1x2u/MHizsCxUP9qaV1s8cq//Ztms
yOdmrRu/0+5zSWH6bjoWNGH2B4YQXQ0czECJqo/1Fi0+bGYasAT7Ul5by2NfzZFG
j5L73MvLc6sBJDHmffcDCj1an9uCsW3eIXSqnGvFDZYiPspjwK4gXV5Q1PO4DBsT
wIze2CmxWQAey30vWMZ64rbeQ1gHsegrBZ0dzAAtsI2hmAjLkpAMgQHhsz94cdof
uYv+jf5stID1xIm4Z32NCOhbA/MxJGRqI6D04pR9qiVOPdAw45GdQoDPDzaD43pF
nm1HUFNQS/DcpX2oloNpCEntgP8J4xFXb+3x5XyepvfTBYkjWjb7UzzUJ5t8HDaL
uWP0t4CIOZXyd2fhz25WyTDMRsZyisE8QN5ulMSJZC8fKXP0jwSF4Ne4Cn1f26XR
AB7G3HesodnJSHYJvOe8DgzO6Gzgz1DIInBeVH8KLYalWiJh/LS36ncYYDetkvpr
8U1BXxRDmLzCX5NtoM7072lCmEcdSJiUVBUTcOYOVrKAOgLgkbl8PcN3CrabPdA7
ukgRfLSkBKes+8d9FIflPOmpQTmVF0sU6uCd2hIyAoACI/UfWLyVMNeixdIZ1Rfy
wu82zvdsZJElvPSKsSxM/6Qr3MjnUUQDAw0TqXvTFtp5aX97tiCFIEd3i1McOqy3
X02bAfb/LfBeuu4oEq2DzY8ddr6TTG6nxv+cGIqnCGdXbpm1iUEVUOWEpT8sfTAl
jduoKATQ2BdJpIQftMKCiEn5k3dPGiUJJWA4lMhpFRuajDRY/sufOTqTpMGUH7Hs
1fPEIFUXB6Oqc285OFPGLGzlwpKDuiXB+0AE9mctazxfepd91+0gtBnECO5yPkiS
TxP0MQSLalP5MIIM3AIqVCitPGzZQ/2HJkYgPL9XimRFDYXYf0Gs+o2RVf2zTUSM
WS/0M/XpQIl3vH3HCJu94/k5F5nciOIhyouC8goqhTAJVjWK3CjYPuD05LvPbRkp
x4dlJx1cO61B5VSBEOai+wAFNsc1a2NlxZkMFdWj8lUy1c9joy47VvT731TdwCs8
7Ppd+Bh4KR20QKJzgLxaLwgBoCyE/bx2kMpLcF0n948dDYMKDd5fRb1ojQ8jmg1c
b6Ghn7ogzWThUXymrWe8wPcv8k7JD0waF3xfEoJfp9MXhCqJg/aHCngfMpoZUYcP
jVyC1d+vwk8+LZFVGmnoVcA4wgsEmplEASgTYi/hNb9ccXEeBpd3Xjp8N8KA0DPl
IBpA/tja+vl5EYLxxcTxwBAzAI3llpZSZ1N7uupnd4l8r1M5VCe7s06er6AnVTEO
z4bXCFucPvxEr1DGdAfExo/OoXbap6MFyAMVUuzFCPG6dT1xE1Bfs1aLhzv/ZSzA
qgo8Rbn47aog7AxWa+NpOhzKq/1o9oTfTJ8A+WLJEDGZSrNrPiQBq0Z2u0BLGwPL
WIQXa/5daz/T9PJEH64b+yqViYhLuVBLjQkRa56Ai7AGgS9dE2bfdF3+Coe5Ybm/
4DPzY/OoYba/kYthja8CMQP1JMFy8x+pc5kay9zdgkwc5VT/bKT31QvWHppLk9ow
cZ2eqd1Urolu/yeiOS0jM4JdPq04XWnWGqXT1ZOyuaUXmk6GeZmxuB5b401qNKj/
PdoFMpYRWNCZNmDggi63pe70h3bK3cdRKvJdZ/3zumtxNDPqfrBigQXcciI02w08
rokh6m4KewgTLzlzkOwYO7Ai1FhWEdCWtBv3/NZH5Zh//gsKDJduRWlD3oW3G39F
CN+9kdHAZMtzmCIr682zIEmLXeSRPoqm4rFNKC92at4WRJLmAx8lOwI74trYcysD
5vLfuppKJMdlXsBZnHndRXlbZeAf4AJ5eVGMFCeA5CRpZLjZ0uXL/mzXn81EutiV
ZnfXub0fKidHYC9/N8z59ExmmZc8uOLNA0h9vi7OfOwP39qU9e9fZj9ybkg8nJf3
uW7ixeCc/GODTKmNp6aAKuwIXcoq53srJUZThJaNUzS0+ExIbUOZdio/lFc4aKOA
1jCRRv+cxfnduIZMezsvRccYFCJNO0oiTgGeGu5yfrWuhLjiJWJQoLZO3IRz6nBO
kZJx+5+iDRTMchApKJRV1wdvYU2xKigOetKiIvR/R0NJ2Og3fNy8LYqo7aLr+nDg
JikyWa63kUSnsgBO6Mz+fCsbUDu/d7TBqNzT+qYuE6RRzf3+0zrs3gWiVyq11k5n
8RI445d/tHevla7/SCugK01E3UojUWGNLniKVyC5fn67Z/Ba9tDs61zgQLsHGpuk
mlEtMJs8fvMTh40x+5YlDyJiWgM9sY8KINwgXMoK3b/SN/K62Cn/SeCJcxoLBgZL
UW8fxfIFBT1UR4MxPbkY1Ne01EdY9wDtlhmesYyMCtXFJ/KhNa84WKBEZQaEXVP7
Vrf2Ug/koVXJ6/+lykfz+qiM/Fcl3oYOInTkocmleYN9JNDn2w1NG5Dxb6iQzPSJ
YfoLfI+1bKMZujqU1VA4gKv0VttVlBHdABQxrfunAElzE6ZpF4TU4P29P0Y7G+FB
RY5jYji9c8fpEfjEQfmJ7r5An0Wy+DDjD09pFib7umx/NpmH1qw1lehOClZqYpfv
SoyZVOYijlv5oNn/BvJqVZNfldzd1Anod8yD6cgUywlhRp6slJ5quYLGKWmZB/JW
WGlQziwkjoMdPi1sMXDpKOlRJvUpBfwJpdclquAdCBRSXki5ewJzPtFaMmamnlDy
rc0hC++x6SpDVjtMfujGo5grShS8V6dWk57IL6ITKU5o6kNvrohiRnbASPr7bKI7
OctFauxhTLraZSzPvtQTxuBnuxLGfDwzkm6ukdTlt8mhRU92cYnw5hB19zWTmSra
7EIASzjFLGGtu6RNSfMlIkyNUoDo1fpQbf24T3CNSIdbz+DYgJKilXAAlJhgvcug
6PtqCgI86QJDnQ6etSuwKecBZjC/ZScBou2IRSW+0Ihk0Ns6wnfSQGb8zs1zIiBE
0nLXzII7FxKk/Z5uQFe3VZB3u34b2TXsTiccr8YNLMKHv4wkDY+vFBWk/1uf/RVW
F5gWJ9/Z/08smEzhSegUijON6Km/WsjmvuABU7oRKMxugLZimfIWQNlL5fG4+fIP
eJXuR+gGJPd0Bak3TFZSCc3n1sI0Nw9h9oLSvCzV9Ky8LX3VAYsgGaFH5dZLrEGS
jzKHRFZswlINi7F3T5Rnr4oIybcDFwS05Mq+kVyFndLsaTlUYSpNUOFCw2F8AOHI
+FHPoyFntlviTjoIlDXBG3dw+4m+f6mCnhNhKfTpMbmtQ0a0/uTtpkvk3+hM8HUa
Q9jUxwEdl6jCCILWQ+NGx5I8WZ9tIlqD4FayawHFEl3N8q2/LOhfLG3DbSyqxs9c
mTH0G/3Bq5Ro/vEt4SegozczT8M4ReVYVkRogPC1iN9vRefpbXV3vu18L+7aoSQM
oNYKU3Gac/eENe9kggVEeq5a+9cJxEr9TaXS0rbmdp+L4cDAObZOxdCr0cogEpCw
mU+8lCWO8B8EBSBmTK6yO3X43WrBD6WphlYcRVSdJDHX9YSdBAja2m0KV9JYkcIV
h6W9NrX5RxwjDAfs7vpOR32f7e+8Ay3PmBtqX8Z/cv4AgLeV0KM/GUjBjMeRvmGZ
MZpXHpwf2vutheBP+qlUW1l+Ax4QRilWjfkkUL0Tv+PTKt5gUcf71+jP54GUiVp1
sY4s6597rP2O+e8mkXuilAHg6OZhXZVYfjBbrYExkuKG5dJyKwH3dyL4+VDxfCOT
v5ZFKNeR2mV+CBL321pLP1+K17I11sV/r1EB/IgVpOvFpC66xc8IBBtnKYaGeNWW
ZRfwA4IiHSDTqTG3I9ZwF+Mxl2B70+ZaWN7ikhDn85C3cHvrbs58KJa1cTopjy+v
fAcu6/Y1kM41j7UWKCD/IKpoKQZeKLaJX94q1Hd8Ajf8o4yAKwtz7f7clmzI4WR+
+kX50CMBL4qCWzGpuEexNdSnmiK2dQzmJ8g7umrS3ie7OPCfPia6akgnGJrvbysL
jyTDbYovENC3La0uUou372WTkcshx0PQiP91MCyQ3OP0zlMrWZ6DZRJMv97hOwaq
yvr/XuKaN4LagYVm2KRRbc3HHySFQ881k2JShA4cwnxMqPMZTC1mpoBfe6/q/vff
Pn1bfCCN3EsmOi9f9Prqq3VvZDZp1ZJmQ8u4UWxWZp5aOH5CUL5DZ53odaC9OcqV
b1fORlsf3Z3oeplAHzv9mbacPqdwKE1SXFv4/aKp7h7qSt/joI6ofDrSAG6hxewg
l7UWqsDSlOkLef1tCss519Y0qcrz1NG98gb9r+5mmt+QoTURbnjPIw9XIbe56c8T
ckTdE+nMymubthjWowiCs01I+wChE/Qcnz30v8h1GKP4hMBIbcu+wJJr4O58jOgf
BMhgtzaa8g7fQsMyicis7M7xONv/9OgdLVIYqUPN2+bYTgUsMLsJUUCYB3wWZ9xK
X8TUMOaUMdwvrQt8db8qiRHEX/ysben/51BLvS5wUi0iU9dZZH/XZhaMcZ3S2le+
3wLrGkhh/rTLibxM3c6Ba1aYsO4cNtfyhNVP0jBQgj3Dg42qdIF6sbelQxSNsFhx
1KWT2E47zHnCORBdJsqc86frhRquIeFNHLw4EfdcZHoAwpIZDV7GykqXhwbMJZs/
aAL7iCosZoFsnyUUzvJE/zcDqN+vJ64JBE12pyrEl0k9f6ID5+JsoZWjC41CPQWk
012/iYuJppDj5fNT5HHlS/951V3V0JloMvGNG62KvNU67IWK//arv7XXnuP4Wbtb
AmFGWwvFSu+RVX2R9fL4RJr4M6pmv1St4/6mVbB9GtwAAIcEl4pgtedyxgpPArm+
8X4kMCQ1Ud/dl3JrTBdfXMHhJn2GBDl2ThVaWsEIr54WFt+2yaJncDjUMx2fZG37
UyEC8nqQSVGSGgNZpaVJcNCef9XYpSOXVfkgzbIKXin0BcJvuI2Doanc2Lc+f+zy
kZCFMLCNl4QtCnsyJGxxoJ6cWCLh3QjCuw7ousebwxiO20/r0YUbgaDMDpLxn2YO
TT2I9VXFMRv/i8YgN/BYLnuK19X81xyrmcHRCQCZTzTDbRcqOZN9pLrTJOAA113U
2ySxpLfyI3BdyyNGLZc48jgRVyVZtWGoDcjOT91Qqo9tjequ/nlV0zagVMhPQIII
H4sd3w/hA+HyECLR7XZ+JjIQrYLH/VU+t0AKCZWnl3ukVVkETSJsErxJMMQ6C6wG
KzrIU1EUDLcgaXgsPyGLVGaEy8MH/wXFuSVdPL/uJALOlrK3UnEshDRCoeTCXgd4
MCnh/Edkekz3fDkAgouww6PJIXfutCN83djRZEb8q48QeHqaF4F6pinMQepx7Mx9
/RLwCEHMRohuzKHmGxrQGxRpNOMD7TVKGCipiaregJSLNQVDZy1A3WYg55hLNvFq
p04RkGkI8oGkIg6qky8c1GyAAi8qTTP9mPTkl8h3G0OR5/Qw/XZOFUq79Xs6IYtr
c4zWziI1VzJPO55F7NQu4IFpkMH8ucnmkI3359fYUkt4IbAbHiu5+vujxWguhbwY
mlIncrx9V/AR8ahi+3/XeqIn9gIBPviMJwOtxExj+Vp4RudcPimRVMyztpR6HATN
RRkN8+iLQKmrTTEes0ZBNvovzBzyI/KmyLdLFYyOUS7ehnyeqq+PDrz2jd1TerBM
EWgy9lAA7xhPQfPVwPNvWbKRWNGhWgn0PS1dTL5EwxDsvwtIsu6NX6+f49DibSTC
zPHx0u8wrxY+RIFeG7+0ZnrRSKk6GWjn9EWFbCdHMNhraL0IiDVSofUDXThwXSfk
SnGLPrxOh3QPheYLEOBEpzCwCiiNS/BNC8/SqY1PTCwbk3kqspheNp8ZhoTs4IYl
gi20NO/17kU/wzdubYw1ITQq/aswoYt01LKS68Gp4ZTnrZXXYxg+D19JMhrGkRSe
D06SyY5zhQBbJXCA3tHW5on4VBYjqskqeJ+YnaCHKcYBYb9NN02sogTySzm36W4X
1aOOYXgnbol+V4rjv6f2vxe4VGLGih3Kz7flWjUk/cKH0Mlg7u4pUT67xBXweNxg
VkmPEoe4equja4Bp+jLbOZ2bui5nfoiLr43K9ABJyBIH7EEXXdDAIZxfNm1ieFKo
ZGU+ecRq6LAvWgWG2aSSUbAdDjhQYCgJFApKFqRrvymPA0cgDC9vt6aRn2NddLBD
R706LjBUkPiW/Acz9w7jSxzQ/oRfTiiemjMk3zB2/abrUY+RpHOCpgn0SeosRJFK
GQGW+tOEzMBPHYcKrMoS3WPA1VsAriNH+StgVxCiXOZSwF4Z7IjdP3n9djr/FYyh
PTyqNVCNLWFW9tZBC0zE6zf+SpdKXeM9ERiTz57PCbNVLPTWJ1N6LGT34fpEWFK5
jyxWzLAJOZe+LaB+rmluS6oM/nbFxo5rGeQtr8UPv1Vau8FuI+72E+u0zA+tNcTc
9nUda4PkH26/K7atkn3g7yx674M/L9ZPXWISyt2BRuSKHH6OUTsL/lQGNFptCMEZ
R1Gh6CtFhg/yMg/lb78ZVr+KtEgjed4RCofqk6sSNcTvdpMOtp4sNf89BXtAcWZZ
lBGUYDQKMCD1E13UV8KXhfTtker7Eyb3pquEG8POxfdHj47rNfzAPn7J5x6gc3SH
d4t1QbtGgXX6NtlTfUwWjyCBphLNqgnksx0Wv4h7o4KKmC3GpDyH6EfnzRvJ7XON
jdEmFySPzi98MZv7wUZTTa5MaBX0kuaa4NJiSCDoMUzLhzwtop0CdsoeQzvvFD81
p9cR5WIu0+1W4HVfdNn67S8w0L8cpb6OxiO8zpr9nH10fe9Z0u3zSXCziHjg806z
u+48WR61867QMz3MhKbPKhK3n4Z3W0loPhvlg2zFzDAG/lvdWFkzVokdRLRjBfBc
7GJfNstk8cS0it6NbPuKdP5cYRiLFfyug08G3moyoeV1LLHztgvg0SiS2qbxs29U
44nvuDZJr4OAniN+iD5oLwAq536bF0BUWtoiGsMSDIY1DDPTpHTOaxYgNmek+MGZ
Kmi3NIzKx/MyDsxFOeansn63HfjTzNXS/BmzU0N48Kyees3k0KREEwJK7GdafZ2Z
wlIVX6Zfg6ojy5pjEAnFuutrkDavJjlIkCzFSYGFTWlVblkPmJ6fxlwxcgqoOLv5
VR7l8k7770t7reZbGxGk4XLgaSZy+L87zCcdBl/KLjgWS+AOHmX5D4FexbPmkxbC
0qHIXCFsysXQ3oILhQo3YSJKhEeTHMTR8IN/e1cspAN9V8ZozXSjmX7kRz7dsOcJ
+JkqN+aWWkliQO7fakuoCVj+xqFPg0Vh7uvwAK5gjWHZ6L3T1sirKI2gyQAkg1yV
fgr9lRr99E+I/R+aPHB+sb5CnUkfypL4LamEBoo7qGBUeh6n74hKzfyhK6DwU9S+
7arSfmht7OZQiiDYzPr88xx/kP3XkZDLyjs7+OQElZarMrH4v3vLg2CwNNTJrL7Z
VFyJAFGUCrBxjQ1Wq1jKSj+sxbU4bDRrLbVCb1NvH14VN+YYujFujSrVpxw9QQYc
q7FKSKOl/RIcl2kHJMpbIvbFGze617Jor7M1oKQ7SBIgms7o9Nf/j3hbHGHXlO5y
CWMgvIDGNtfJbFr6PvVjS/fN2BQwejLgqACqqmMC/yaKcsI99xtc9jFKj9WWpGqS
5SYQzZFhfRAAUzEG8ze4Gxnq7fSWhW15K4pEJIKpefcw0NuaaXvN7NssDFgWOhsW
IRcKkZZWMo5hIfHXH3MBOz2dbm8jSNYenxA7TtEzcJxUFhOj4JvzDI1ff/kr3cFe
4YmpWve0Q41nJT5zeVYAxXb1mHVS62KQ/WpfVKZVqqgCZIx1sgPyWZSgX9GOrush
W96RxHun3B5tIhUPcL5hw+nrauIoAgAyQyGHenXxu/Ow7NNYwqyIT7WWRqvEelGM
FBXs+9a8szeHL2OFfwrn42LK/vHgnV3m2Zw+sBC5Zgp/MtajRihpDHVZ03sL/bxp
mqenh2izKpni4WFZmtPqL2JgBHaBrn3r0CRMKk78CMa6+v2bAuIcyxApXlDDByi6
JLtbokBHT627antxWflpia41PcMEe+eyBzHYtclvlhPyqwd98T223z+HsLq1Ry1W
VoXUjFOp1HWt84UzF6bvsFZqGLus4KVM08iH6p79+2jaTQ+dh+0l1gQaJBiSoD7B
gAdkmltQooeLH0yxpvnIXPZ8/3lQdLBKPBQ9ScZwpQXT2kS/nDliOrRQ71ixbI4H
5oDsYVNcqkCqkeOALTqKOyOab2M5qLDVP6BWXc45felwjIt1sd6oChsiXJFqU4GD
ndMIoU4z+PYb35rjVIYYMxf8g+IsTu92X4GCBJ7p3Eh+2fF9/k2xXUsuA2SL6f99
CDETj7e0VtgaHjPTxqIfpFeT1aKxXQ5Tk0iZKe6J56CZtKvz5qvXh7E6Uf215UFd
8LWQ3Q+pbpq8nq8SAfOfAvGki3kxYoxp3dcqSD7kuWjAgzRPEg4+XokO8GaXop+W
4703gXAt9nszhvVCv8ruReCwEcilrQf1cD50aV/CqHpUZFOfDOilcpspZZ7dZ94U
SGDG9f/O2/iyeNLI98a3QkT8nUninDTJSo2sE6adfeNQtk7icg7wEBZ0gq3fNyN1
FoIdA/QPoP7evzs5QRmPyVnHEYq9ykTgGEjKhpU6O/So7yfvYRSu9vjjY7whDBLa
yJgQOIfD+EblSLPjUL9vpIFZq1NiK8RiPcmKjFH+QjFsFf7WiJLIlGFaO3UvIDaR
9euLTT6Vpdk/s6qmpwKG4nKq7Od04U+Vf/CFcI+b9O6mA+FNh/8lU7aLIV8Yu79U
awXSBo6FlcjB1u+jHR5n1weQ6w5lQdSuPTqQ2e6U8ZSJluNfBNu8QiSW2yz/vXBA
CiawaEvFV/9puXoYEOWQZKPrf27Xx4XF909aaa7oUpPSjc8GtW2ubOG2w9lWMFMa
e3p7XcRip6lU5Fb8FYFOP2zA0vpEJr4i6zt5LtFlVOBxg6pslfbftxeQwnFBz66U
ZMlc0mtRa7LhJukGHKTLPrREiN8lUeKYlgLQ7i5eMHRQRuuMOHv+NlOYToz0rhAR
bAY/5J5TnZbvEiUyXNnyiKZIfFMDR9FHSTB+W6Qlho3BIe4B5MhDZ1Nlq34k81vG
hqvtF3eSocviTcqEfOlPIQ7sbxuGaLjZ9zSqleM6d1r76Ru2mBFzzNpv6M7DoeM/
/H3fvCvAZ7mNUFxOltSTgcd6rCNClzOtFe9qM97/MM8Yz4zT+VYCG0EDp9Dbn5Gf
GFvNBSJZm4vyNJIKPoEklKmTmcXBc3t9/VCiY0ZeMsq+IW02Q5EgPTPbwAR6KvA6
hX2Zqb6kmNcWgGouociABgH3af046B/2QN3BA02tTQ7Fn9lWbT31H1oSxD0Zg9SF
ROqkqdIA2BP0wE+GJaOpE8Sfv+qSKt9/vsudjJgCNRZ5dEghsYc6LaeSzpEfSigM
kL1O1mLYdochufK/QYcXLpxQzuLIIt5izaERhSYGsZu1k4+GkSRUGo4zOgi62MPo
vrEQKtt3Y53sAMujGzn5kN6BrM0DJT6jzetAutjyIyISSP1Jwje37j120wEaXzkR
FfFFf6ulL7GbOUCnvPKPWN8ehERrg88QLe3DL32ZUzrREtxMAOf5iDA0dlEvnyvJ
m6d5m1R0Jn7GOOKjrgEAgfh4YzVXfQRhghgszEFun9cwLpMWhwyTY3itIqXeveZM
4oHeoImADxycbMLbSJiRz9BbZ8xmtP4ZSK05lF/VNvnhzed2y1R1hFwOt+Icstow
TfRa0nqnboq32S6cfXauJGsZDtyag8YPuP6RpnSrDt9uGmquX3hywpzfsv30q4oD
vHGN+AqdTMNlIIj9vX3UGEXSgPnTSCRHjcZMSn4aEs4svIDJLZEqOUK7r5Ggz3ct
1q7sBuGb/ZH8rWU0QnCR7u6hev/mvPLsryj2C8NiuUylr1L0UJBivSlOaeNY5DOT
ZL/HuAdvqKwxRnSUPGckBx+H+rfgnun2Z82EqwyaBUf/neKsxziGotK2SwLGMlvM
ZY9AtlJVpCQhkcwCDL/oOE7euSuuSVhEyGPbxv/u1v23nGKrhfcZkSYGew6Qdeoa
l9hC7xehOK095QMRgUngrgguWSGxWP1Zkg/8uhVP0WvUx4Q1V4knjmEki1LLgM+k
0lm7bpR11PqGzvx8LPxB2Ppsk4F4p4kyoGoWrMnDeI9v6X9+xngOF1MWmBX1FjG5
0SU0QGlUeZEC5AvO8uptuG8XNBeLQULHu5jHrvz2Ky+RN0et83E11ZBBZZEuxDEf
P6wpxpjVVtiEZjUmDBpYcmfeotCa3zhO1cFSOGd6wQ5lo4zOhNqm/MK8M4fBBTe6
jNnFtSZl6GKNGOMhVwdl0fBP5Qw9V/rYRKgBjvPCBr76DWYlmFiAYJy6FbvG9A1N
Gwp6gABlZ5UVoQAyV/d+O+cT/UtNYm5GAMKhmdr2FctIFOJ33H2AMkmrNaz5tg62
ExFz3o0QIuD4/mx0TzDDN1tgUawMNB2LvLwJyuVRX28zJN6fPRqJY7bnKwndZQHA
ab+D961VHmbN8cat8R3MyEQUV7Ujrcl5dQtsKfb2Xz8JvYdCRbyOc7/xAqU5YaIU
DlUjr1jQBcp4rcituuYwWl9bzhrSsmHY8xLEDBnxsVi7B2AILA5K5dUDVPpUvXl2
HINALKo3YEYcttr2wMTcIXKAMMGVyHSzkufChDHdiidmXgAalkNU9AXlcd7iJqt2
EQN7LUU77ObrKx06bwfkTcs+dPPMPl7AZdN70Wm9EaVIIvgu4++pUzoFwBlXLKNp
pXcYKBlwL1vkpTRXmg8Uiwu17RO1ImTiUhsjJtb7BX//9CyKcmi/snyG/Ho4eHR/
aE1N7YxiAEOj+/1pO/7sVjt1qiLBqoiS2+kEP8CTjs3OA0jnAv7ewc2n4H6lwZcj
aaySoZ8Fqq79dvvcDHgzb9ExELD5j1ePx/eizkSlEAJ5LoMPM/fesVnbcR1QgSTE
WTK2r2U1VQ3EDkNW20dvJ/UBlglCh75Sm2+zLgY3FEghGjME/cPfUSPaRhBnoeiQ
RQijTRabejP2Nu7cNqaLokNgsN4nyt+12z3zG9fX0litWm8ngEkSh8FuJHiu97h1
RgBo9nvpZKgmU3UtX54cy35PvelGZuuzFJEC5aJkNNs0MjTOuoaZ/Fhn84EgSF7E
N6chVZ+0fIhTuaoin6Me3fWKBenwGptsrBLaE1FFaQzALSKpWh7k8aF/SaGeIans
EbsZvpveRszpz1n0k7RpDL0afUsl8fIss3m43X4FRU8P5SGMIc7wnPuI8ZFn6fW6
UfKFTVC/RWbJFOFJN31UEaE0gxGbOwKRlsxBAMXz29iphPSy5HIZhmpG2EEuJFxn
CDTj5befcJSno1d+7qC/znyY2ir+2AEHPqEZWGhjxtizyhfP2I1UiP+VG1XXEsaK
Io5ceeaJDChkrcXISAHHkZ/c/5zA2jKeInACjffL3m+nrv60DQYUMOXZ3PfWwxhA
sD2EI5dxrlkIFyTR7VSvXLG3HwCZHQ8S+CT0Smm3XfubN/UcpKkvheUtD059iz8P
vY3tCxkiagKko1EON2THVZxdofaIKBEfOIA8NjY7clTvbzkGIexWwRYScXyR3DF/
mL5yRnTpgAKt9Aog2rKfpLaL63FmutJ1ge5guFxCBS0kPbYDKEptHTVGET1/wr2l
nTKb09UloV5GbebEuf840pSgZk4DUU0Gg9cUfclRp8kV6sazPIa9JDvmpxzVUg0b
DIeY6K45sAZCr8p9ygPr+Q+Dgmy2T2oSs49XISJFI2DJIW5I/dVPHKgyZ6b7uc08
LOFe7tr0LVz2yYQb4crS/kTwn7OzqjnFXfe64flBA3V1ZV7bFExUXsOTF7dAbuop
AzwL60+xrLJ5upobBdsu91K0P/bFE+pi3GOsMzOZh6IkV4DCgHFv0ZreF5T9KSEH
opMKhyydt1ejkLelRJQ6KYnZpuE8K62fcpS2MsQ/nwY5vGL2sZoSOQqqyTrpIkF6
r1aqJFY1TlRiqOD4zFL2+aug88qfrNx+vPXvSPhN7/Z/QDuRONtPu/7ygnnKKk8h
VnzDcl+5ZXVwtXAhvRsEPDxYjhgN7ZrDerT+0tb66/gQhHE5HbDIwd4cavrrwyHb
HPcr7q3Cye9Qj/qczm+jsaK0TR+HzsuGd2MRW6CyPmBNljUGwwQXjvfbk+dcRxYG
mBgqA6+5z/6nUgsibv72dAybYGsq5EGCZUB+E45hPHCttV+799Rr0Wpr6pdmywRC
K2DkmTIE29uNfbk2N1S7X/NoPAYdTyitqvX6njAMz+BsZmBIIZlcev9FpXkVRxbJ
++JAmTo+puhGmCQH1bZ1kOhNlU0V1mgAxl6+7tiHZpPuqREpHnKqKsutxVGojYwf
zYZ0AlmNoinInWPIeBBT2FNvCsYkszk3AxbmnqlU+s/k2whFduoMoAnrzVVP2uhP
SzfdbOL5vhkKPc04ZsafnZGTag3d95fdZmnKt5nhOEe1vOGfq653rnLZG1vKIiHf
j7DdK+2Ui+39zQHHZdQMpTVVqvOnRty0z5tY9C86Cnl0Z6ZWgi/ZOeBli4vuct95
eqxLruGA9/zFxBXJUI88cpjp2/q3JGX+Rqq7FpwdpvXvS8LC//A2Ad3maou1CcS3
C+D8PA7rZ1RhudFZvzlJ0T7qVnwBHLPbEsr525MEpRM0er7uqdJ53PRp1qiwz9eG
2MxZ5uOZA5cSTbEpR1Vh3NjqVGKXlE5wYdjsm+dnAxSHxw6qGFtL/XRnESaF1yj+
d2EmHCg6nPGufFNj1EsDEcZuyCj3yAnjxDvxYy8+ksVl4KOC53Yp+bu9c8lxV4YC
Gf61tnzsb4FHG0Oiw6nNw0v7+6i+UhlbEi3BwDd8LesN7g+ZSxQ3tIWbTmWbLyAb
vQ7e7twSTUOOfAt3JY9YIYWx21XTRem9cWPQFbDuLa/UnCZaDQi9qFAkxCohOGYL
ZAiTDcieoRm+FkM/hu9EEA6NcWR6/0faPaPTFohycothhp9lsssra8Tvvgwz2QFH
fCs5aXVRvUBGUpw7wyMDKF8vT8l1yTZjjjhAj1LfJRAcMx3XHk+VFy5XNMDH982d
NB0kOr3gNSB/YBCcs5uZeksxgl548oEUjW4Q2wMwjnUMDo+RgWN3JdAJ2nzpFtKg
Wlp/Q3ejKSsu5UKbeXNDIX0mBeyov/qRVbxGv+UWW3NUajULK4c+4Pgm+JQTWqZc
AgX5Yk6mnzcpQPSO+c+rSJ0kM2FKtfA8tJcTU//gnd+fjPgeb252wDP6nJJX1R0+
cM45Oo+ksEQxA42ctXIoytvDYQMMcbmCvRwZy2k9dnpDUMN62EPfc7pAuObgdmn8
avc4ZztWtpm2yA4QhD1+bdo7Pg1R47bNkvb7jBi0ygnVx0PIGQXbezAgDIjTuw2Y
HIgUGS+n/xWJLUqaGBPcPLjOlvc5QM2xipa8Y/IlzYDBcPour1DKDN3QhBXnp6ws
qysgjug0vqgfBzj1mbAqUTf2RhLvPofvyyKjC0StuAeSFA2sA/yNUXhQhUcKTWD1
lwNmMYBtQvw4lrvo/fetuYuCP7Iy8/lOe292jS6achP7/1QS597RRveXZLJ/pBcE
PENh9X+8YKZMfccjg4OCa4YVr43TQONZwItQQgKZ/Ys24VPJdaDZIce8GgLW5HDB
QA6HGlG74a1yHLchKx8asNXdy4D+2l6TyIMFmhUFFVPTiukJnkSx8HHajRlAxjCi
q24xWV3ThIl73/fWfr/LuJvLeHVQsw+qTaMo2lhxkNDsfKcLuYWaryEXRCf7OBU5
90biobdvTATsqpJx3lhezFTB25DoD1w71wvkfaNemHxf+9Tzc7xetpug5nqRq9z5
5xmATWnIubgpuiHLsAxLZADZOSrUckyDPSaAld4gwxEKmHqmPHOlYPWj++5II8X2
Nkn8ElLyFVRwPR2rY2ySdZuWjoJ8ENxF7RQkaRFS45mAf4TwD4/j1FPVP5uj/Ddo
+/0HOhJ2ikFkmAknSN5Qx+bxojqnoyMmNuXnPi/OY4qC9snv1Wp7JcUx6pd4PDmt
S3yYJirIIKFlbKcndRHS4eIuRYz23w/MJxrlraZAjiqetEINmo8e+qryf2Bhmd9h
ZopLRtUoevCi5U8X5iBcVBLbaLsSVH0BVRro2UpQq5F9hA3OkjFSoLcaICC7UDqk
gSCMtzBfvYBgMEfbvfLSAmAWgemLBjkNjtxbPM/3rdm2RG5voc2zbx2dk0R/kOP/
ir7JMWU+Be0MiuzjNhqZjJ54zVeolIDGvE0yNEtef3cUG1A5JEJ4qjIVpIlB2AQR
nrM/U8mtczkJMmfRVlJYUDsZdVTHhzgYBiaM4tkrm3Y84y9QFzLpYR4oyCZU7E9O
Hv+B0itmBKeZGqJqVZVFF0WxKjau+47je/aJOTeZ3jlBD9k9k6/lqJ+M/bd6TWKA
2cTBMLBDTtFF4U22g+ievDmMNGaDuwq+kaeexQPbuyz2Ac+1dREolHaRVOh3LjCR
WVAr7RtCP9B/WEZsvzFY7jUcIog576DWN0osnKtIUEIPUHMAjDomm2Eu0hpLuu6b
UnuiVcX2G4omBrf+TZ2wImBJ04b2Pumw0+5XmNbsDYZCN8EgcEJWTAyMP+/DMcWB
N6ZNISDEr4zxm8ZvO8NqDPrtJ7ZlMWTKslRWTQuAGWx0uBCzFTJ4MzcGBAte7Yky
XH7nJVX46rph5eZimeuhnFLAE/M2DNegnHZ2daY6qzuyMjgBFlO0m9X6xmj+cL5s
lj36LyVDFTAfSNvvULKsy21uVYKEzCp/pYoGjmHL3PyuRwmvrFKnthdPjF7Kmfi0
zyBYj6DRQEBtoJ54Txr6a/VnTodGqQHg8sstkSrUY5de9cP9WcYjttRlQlXyBOgD
Y/M34WbfUq+cpNoYO+cBqzfZVNq1rdr628lAkFZGeODggy0BpNkItqtkClDxBjwY
/DUYzFxE/ljqXFBsHd2ptq2Asf2jNsCpI/6ZPvjwcjomsxHKYHsKtPQkHOc8Se19
8BCz9xd/s+M1X9yOYclVGYVNbLvRk2gjFxaoc8OjY8lKyl4dgjoAheT7bgvoDFRI
MSwM5zct5nvEQ6qnJDZUnXOC/bZFSNhQ4PTyyReULnCKEXNjbMPjaFPUsG+/lpe/
5WpV2CR4KLNaAKLZMnLwtJdOp4GnL7Uy6fJlmZsPjWYb1HNGemgcTpn7Wy3pr0z2
KsqpkAPtK84mmzx5xbjjdXSthrwPABaOujLbozaZLJ3Hh2OablproFRZZ2UrVGR2
ujNU/qPW8Gi3TbnWIdpZTxpWhwder286bIU5xZ59sTOBfIJGsYdaoJH/DOINUk49
1v9EnThlbWV4Y8zMmNm8BZqlEkINvMU13Si6qXd2rze0/qTxpDv1cFDJasY9eGSg
3FWvXHuvUTS6SZVqa8K7c9BjBgDBfzbBeeuSkeA6gHpP/0s0aqjhOke7BG1/rFoh
lGfIS46iqCGxssZ48badMV1CTvaAyFdTaDlylFIp1oL+9Vgp2ccXUNN+j4hjcyh2
Tg5KU8+Ca34lldy79izucn1pB5j5s26SzTK48bl1ljzSs8I513wWnYoP4U4Q/IhD
iW+NmiwKFc1iiulM6IrqNqIcvxpoa3tAJ32Mu7/kQAyd1Ee7f5mQ4LuQYsviYYSv
u7XSBAzIaJdzwTg+d6IycVvlCT8JetHsUp35NiDLXiGy1F45dSp2nb9YuhTdnk1D
mVCuIAzCBwCYY6AxilHgqo9NmSzQcVj1ixR0HmyvMxBh7ScfXEn9owEEN2uvKCGI
VVeta59XGKTKX2zdh59z+n5MtqA/hJePNEbXhoVDALgpp61uh1Lfei01B1qi8aBP
26nz7Df8Vj0T9XvfH+wnNT1TWhk9H5InguWKEKT9h4Ms3qRKs1zF5Hecn501dEll
fdZE0LM0ZMfr7+9x+zFG0XSzg/9Y2y4ueiYz3HuyExdOevdxGxsHpJUI6dp/6kBh
4Ut5uX42zrOXG2BT+lLYBI7LKbfZR1ZO9QPosOK7SOq37MMzWrKRaF8LR/c6kdk3
7jPzg4mKRSD4CIm2qqwAKuCINCmihpiEQYfPp3snYZ2NGZ56pRnUESsNO35lL4k/
55VJTFLz0rD9nUWCrn/4/6jo//1KrCbGBGurxuwb254Q0vWtu2uOOfN4N7kPAvQn
lYEwMpUvoo/FgQRe7MlMHvWcZHDXMVzWbhaIHKhDVdGH4jwu++Y7fNqDxY36YEHr
QBWIHMt3eGN064aLUmab6k3S01gD0A8rZtVK+mody4gLLEyKWzh1M1cU3/LdIpRZ
DnEqY1EMZo/UTFbfvDH3tPp4F30gakyDEbVjaXKaKAbItxZirS65ZUb7BCbaFrhL
jxoXIz2fcDqJ9gcWz370ZU+MW75/qdFCvTr0WFWR9QCOZjzkASvvWjm3quDmRppr
DcEMiC8Egxr3pVdGE0TfJOqQDXGAZNXEVO5fAodx/8f3avIwrwBaOrMs/ZHTt1J1
6cEHJpLWNO4ZbxJN1Su2eSw3cN03y7Yhf+bQ6IUQwrwVFP5gfgaeqhorRM4VZFze
IywXbaB5w1ALHDWdDzradqGFWi7HDMKl3n4wAZkMbKJp15ZFrV2z4RQE3QTjJrh6
RpxR6t09X170Myjs4Qx7YoUqk2/WswgdxK8Grsv1R8fU2ZabQjrDUhOHuiK/jUlh
BTqgP8K+m62d2kOtlmDyJbjx7zM62W4KuViP8pF6I91JLRkrO71mx4H11AZSTLJ2
+NR8aleExeJYr3wJq7BxuyFOspLKmSJt5JL9Mww1RSNth3eXayGnqx9OGcfaba5Y
0to8mPZbNT467ezcXYbZdffd2E28WPc0TuC5pgL31qQpbc1UWP4N7gVSpDXzVOWn
apySR/r7PAMato/Hl5PejjYBXPQtRd9P4zlcSOsJyIXPY2pzR3OPsYDVH0ngYPYx
UVdXLZnYInVigid3XVN9F2AoPXPNPG1BQphygnx49iNtnomADs23PNxGqZ+GD9fc
tl+So3yBTYUnVGOBocw6zr7gi6bfKEKclwQBHG/KW4IQayEyRp4Z2Cl0IXP3iVBu
Imf91VH2QS6OrTwVnl458o3EILywqpOg7oHPpg/1rMjRPLzJo4+nB8EphD7X6mPo
XLkFkqAYwsVx8Uf1wVvqESQRiGuPFoJ1cennmItRq82YkU2mUyQWbnUePR7e9JBV
YU3+mG2z3JOyW2q/l2F5NyVJz1j6qMjNlxOq8ETOPeFNNPVax8hbqPGnmWjhoJcX
/dO+oVsS0dkDOySecX38LCzEf4/MeDu3z29ZKjeF2mt1SZCHqpw9qaHiV/Mtz0r1
dYFyZ8ycluYftyW8nEBs7fVqq+H5ugCa7dm9RyEKtcyd/Y0RIAFFgeRhz3nTBkmu
nmt9iMxJd1sCW3ubkIUS+XstY8393VK8gZ/1HTddre0tmizVPBqNDiNzS1iyYXxs
pKbH1g9ugW3RcAWBAQ7zFNESSqMAa1MsO+gAZkkS9ilT8w1MkQYDZzl8sXInHN8b
OykhAN6mjpal3/Jt2en3W9KmWIrs33vv58GpkCefRfQSVdam8mFM/aaUr40XnLA3
UWDskqVcuXax5Hhz5Rv76j7ro6rzFZPa/qRyZiuipiGnXjUsNjFYYXylMwoWHoVm
qiC6s7IKsgp2+6bIDJesn+wMlo595f8HiZqDk+1XImwkYYyeU08NP2OS1Bw7mbua
vxcF5xKPX+to/gG45jNoHCg966Xs5z5lVR1kg87uhlT2pKd8zM1GzTtGurVnE5nf
gskD72s42XdTZ8W2NciNzTrnxO/j7NfprTin+ZfFkcHeMu2KUCSZpHB8UnOjDphD
kn3hdTSonLPWBChrWntWVxVW9lRk+BNuFLY8faHjXZnH8bqfsp/FdSIHPUkDuNhC
WJfpg7YugAVDRy4TGO+2hMNVkBZLlTUUIT3df+Iu97xlFsOhLbnEQXxnmA3emwkN
062YIPQWKpo/4JQckIF8jppEAzvXI2MupaHlF+dOMuOv9CIyO5z90B5e7FNqivu5
n219KvHQHnjeXx9wfSHbsaBldbQ1qHJuH2RlNzVT03vBmcxP8nqUbQvAeUYKOl/I
S+ps8FDiCJSM75YHv742KE0oqv2mjasWIBAwmuKx7rKGChyHwsjRYKfu+3KtQqfw
UJrWpTXPlaC6gyKF8N68gytiaJLe3zv/JfPweGxgLWbXYX66hXmIygA7ZS7LCXjf
9fLvdnfMhzFodi22EoEE16cA4n3gRPhsY7IT0huqgcI1Bxio9xkcUdUYVzl2Ay2D
0YHJr9uROU2iUfXovrEslIZ5Lg6AuVic3U7eXGImt5rUVyK3x7AdMRusyxFmBz5m
v7ttG3pfO9EDUagOJ1zYiLGaRcwOwsweO8dMqCmOwTUUSCvW6pNs87PL0+zuZOte
xfG+fore9+nnqIiZnkoA13Ico5JzWNKp/GpLDMmTi62pKa+dBC8fJ1hQXAQGlSHa
3T95myWKP0Or3dTZ9ZvAMvFIBhKywM3NUq4GuDmb8OehT50BoHfY+r2YIbkK/RFo
7+rOs4E4Vt1jXvWS7dS2UhQQxjAxy1aNZJar+g9YG4eUXB8xMUBlTHN8I8PthOoF
3iwctj97EB3uAem+x8Z0VnEk+BYLnOWnX3QVMlVdzMuLwb2/R0hf8+KvIsihUl4/
uJeXMLBNnvOwCoG8bzM+hp+nzDsWNTl84oMenB3U+Ip732hlW6psEtLlBXGncdS1
m6jW/QWBNKgpMLtRhpC4oInaJpBLRoFdWPqOXul9B+9qj3D4pDCVBFJu8BMkaprS
oQ0PQVQ8M/CgffADxSxLvmhIsVIRY5eoPW7K9sjtR0gTdI6rt9htyQ2CqYl+DlDq
vuR4Y78otwJZwN5ZBOY65f9wA/vyGhFATaoY8ENLD3NbKb0lDBzXfHhIkicllc4p
u3eEWlgSgrGrLm/UfYGdNrsRBuvqq2Il1NYR/d83N2tHPAFzy9nXozCK6gkLcgJb
U4AHZnZXoXzP7QiqozgZMXAb+CEtptO6FDWaAF/oK7DrOnzKAKGMWgYv8Mkxw+OA
AJYxVcLCB1ArrfQSVMn/e6eBsWoWMtXSwZWJ5RVEQnCHdNMlns01dy/aeGdQiSLu
znbpBUOocNLkcaPXgU1rU3H2qKvR1OwSuOzMuVoXnygzdQxSj4Nt7jQzmJ0fl+PV
TxxPyFB/UBC0MnpqNqWTktMmPA2+SqN0cZzpPJwMEbZdngcs3XZfJ8/XBScfrQ2X
tSHlEM7z1BPkihU0aLSzeEwKt9DXYCPKE3F/OzACCz5XWZ+OmhquY7c660hSUcGo
0bCRUCsZMvet8kxqNibAGstWYgralfARbaThaHDCit+5QtMp/xL8oUuqzT/Bx0Nm
L4nfELmMLaclA4vVQOQtsWB3Ork/2eZvU3EYO4UjL8sD6kJ6K1BhR9Jovb98TTET
aQ+VMbF2+MfTvxWzAkROA3xr+a8Rr8GGuKXLcxeTi7WWsam5auxsRW8yh0GzlotF
kgafpg7IlNS4ElAmlyKww4Go6igu5LrvXMK8WUoYpTkCmkg6HN12LgCf/2KU0mmA
0AMB3uB+w9sbpFZRs7U+C/r+ufpYtZpeRNv8c/JV+AR/iUIqe4ujz7iqKyPXMQBs
lF6YidenKZ6XApYCAu995oQjskbuwZTqYWm9euxPgJV+ax0nmYy5F9WfoloQ+99D
37DMmjNRW4oI+S70D9Vh6DSNJmHey2YOudKWqGtO/gZ81oEW/Gw+VAO2J+HwF4II
rhfaShFgCv98//f2GnyWRchNV2lVJopYUdd3S16yQucAOExDMidH9wBYZZPWdN4f
mEm6ETYByVnPsgIwRuFbqRI/sPWT2j/M55jww9/HBWA/VflztFWbilu4eNpoUN3H
9mVaf04DSfCp6IHYyAkL7PalzMf7JkvZrlTwkEEq4m7FjM7R3YVydwM6sl67aTIk
Yws9FTmlPbOWefcTallNH/ozT+w4mU3VOamrcn+sR1Ry2OYVFDCd5LCETnyJaIuu
T95nxLgmZp5NFMXKfcJpSC8oxJrsF4gZZIrxC40YV02Bmll574p/f2tOVT/lvbbl
LtjtPx2uDH78ulsm8nn07ROpl5WdXFbB2V4xuYjHFfy7XBx/zRXznMfB0wIia/19
Lduqm9IH722uGJBpkU/DN14CUBab5PeWKR2Qn6g7JcEItGki11WwZEsc6ApJvIVl
O4W5Jm919+AOfkUSOSHQ65eivuD5zPU7kBGnyv34DgDOFh8A89dx8mq4jwflvGXA
ybVzgz0iGQh4LYNhDKdA+L6WCkhXX1aMqxCNoBzkmYKHq107GXHUvldlaNG/U/Hg
g5RjSaKFPEz92hybPi4G8A5/yMYIjed6fkfhKTZQfMpi/LEfAmtjoopoguhy4iAE
6KQLY6mTQSZ+Jp4tduHsb6vdEHmSlQ0N/s1micvDNDwhBaOmF2LHsFjBWEPFzlPC
2Kh2EzAE5N+np8RAfKmDmhy7Fm/c1QROF3iwhfoWEz6cnPXm2S5dcITxRHn6/sNl
xGurEub1IdyvEpiIHqw3soxiHhtEk3FMVB5Evnd9zXhfaDlYEWl8XMD1OCg9Pu9K
pvahZ1ZTRvUYhaPM2/N0LlNAicBjxhafjJ0/HKqJNgVa625DTM5Lw5xHwddnyZ9s
tTnEXjZzlLkFZXhoIDkYzEvJ9eG9CujElaQxXNpE+G3IJNJ3aqGFIaSufpNpJNSd
bsrddJ5MZySaceIZkhau7+2yKB8so5F/E50hMbiJ5iT5hzT+1XlQH1HKu5pIGoUP
U7oUn5Em/e1O+CPeOcivJnadhMGMXyKI+iKhHD7W2ihPAmP87Cxi8Q7FYLzz8WJC
2jQhqQ7tKLaBXGj3gddWfQ3bzWwrvdcDIomHsdB6H4kJNvIS3CZb1h6PQF8P9AhC
nTaSZYC5FREDLrIke8Q0P76plMKXUtGiIfP5nJKUQeC4a5UuGI4SA6i1MMIV1juO
SJ+BnL+t8mksNpnvVP0J+wNEflkMEHMw2LYv3qnRjhjHIvqSVQRi4QtJh/ByiCHC
T5m16xRRbpU9Q176BvCjkKhbseEo2fDuHZpk6GRpAtA8DdCTRt8tPtB0Sk7IyPOe
1NrLI7cRDZJtUswgX4PIORRZ4GXpQRRUx8cHk3+qpcYo6SbKZqOyS5hh+9Fk9J/S
44WEsM0Osbvn7apoGTw4LvN8wTRl1xAxCsr64lrEjhari/0+IqwG5mSuPfv9i02v
ha3zVsomF0dbjZ3tVqig1jEa4O8lZJCmWv4VFlYO+QnCjy6R/Vr16FAUWjkdP+OG
0adsTF5La/GRFA03JAZzrRID0U6Vy+CYx/pjZ+0ntThELrKGnl+F1N4V00y6+yk0
shBej+uJ7qYa+qN7h8iHmupdzeLDkZCWUDX7fZkPfRr2ljlqVUwE2bhYtiLnYDi6
DV3PZ083ymWaNnk3O96s+RA4qCKt7TkNoTtMPDdqglZQn/tHR+sUUvponWnY7scW
HySbaBVxLT9pIa5TN0IzvpmeW7g/WXsLI0ghwh6UB1dfsmeAShrZp/Rs3QjCuwGJ
j117TfBbHxR9Xz1KOGwMVyTd+YgeL3rNe0bbvRhTrf++RjfZB1XPDzWCIzOuYm1t
ZbjdflpnMma6vjowZ798sDchQ6Q5wMwTyMYHYvjPLuad+Zt/BSZl9APrL/8ISQ54
RVgHGMrwfRqmvex537EpFeYKxl3t5PO4BjMVMp8HtDF0CSzSgvNtaZQAU+o3gd8i
TvRQRXVVINP81mPm+Kmd5y/fmOCODjCvgUaQgELBkUeo4ZFSJaNosr3MYP9lidaP
t/WxrfQIjbW8SIa/8UxGr5EpL6Jh2C1pftwTv2av59mZn7zwDveZlEgAGm1lg3Qw
k4RrOqlrn5JLdah0nRDzt2cvFlq9BN0VOAdbfQWs1xfcvd+wBJeUx3tIi5BL8xsm
ugnHc/7ZS68ZZV/WKHrKTT0f/PKI55cZILaRWEcc/erzKyeZT+5k323r06DUz9ms
e3rawIjaWIYHeN2muV2Gy1EYh8E7jygHRxhoreCi8lUaxvN44lecIzN07SFZwFWd
vJqDqdRznCTbTAVYZaULdnHjS8vAFBbD7Ebefw9qViBY50l0hbv3ooMbhgWl65bd
JZeYupO8j+uVUJ8mKM3v7vwrCVB43KHctJgysElHGu4nkr/a8+WkdCKAxBZv/nbs
PVdgrrvOlNxAD1NxShaYBl5ynYe8htorpREfMnKgViNWNQu743ou5iuQ0LftbtGk
KykU7xrqx5NbuWJnph+3srvmu7dys7GKIN9Ta4JygnpjSzDTTDboF1XtuyyNXlYO
beR0tlqDLcWu/72Rx1PfXA9NHqOcz1ZsKqv8fIvODidpAZatDuKMMi6geXGEg/sR
idlTVfWrjJ/PAO6cqgVjzw0Dyvx9QVr5qL3MTDYi+G90XNRGTaFrw4iK96+rZ199
t3LnIJ/mgrXtGQmHT+2xTYxCfGK+w6CfX28xJh9AUkznYmAW1lBGfzuh2V6bSpVy
QQFEgQPVr7zNJbuoqKamJUmwoHlRRgPl/sbY8Kj0jW140yf1PX97QUO/2qvf+08T
EVcLp7qLRg+PR0nzx9pajVIjfNicUgrSAC89Pdw3HR9OUsYuGxjiVGIEiWO08Z3p
R2e2GUhfvGiHpoYSPSJ1xkFbCAZJIFeE5912Xhk3t4ho5WmnHzdFteYiXF2dS9RJ
Zv7zKgNXVHVkN6JQvnuET96ZgQFSJrBVQpo2sfLH0p3fiW/+HmcYcsT/NVoxMJf8
UEItFVQcfWC9KDc9LtuMgBwMyEVDK7mnHXcb2Et1wqFbltrNoKnuiuUXuXhOUs79
8gNZOlP+mojT+OAXzNRr4bf+SEVTNRti14jgGbaVPLPmNvGh8FRhranFKt8M8EIR
LHHlBtDjQ9/yhwgvzWQc/uOKp+fQcY71ZOtxe9GJ69oYXOoeuMFfuWiAPvHFdA1v
BXwxpm9POiRHUJz0S/vWxzt6s/rHBwrDxgwPQiiEethUpYk+vULOEDAydKjeMX31
5rlkmYDTqkWFM1U7DsINCZTKAKv39xIuHow3HVrac2ov9b3+rvQYDaBAe9w0FpTr
ddQjBplQ6tpDm7lMem9buDdFyqsyohLLwq+RaweNRg83B3Z3xlsuXEoPATe5OZ6y
GRzH8aLKTifqu3TYq+qeMUZT64LNshMXe5qYttVwogNzAPC5wT2DLSCOeUPBGPwK
zk5VXaQX+lvup1HPAlwXmKGZ+Pt8d5EW9zInUI4haHxK+FO1+I9A4BMuma7MLQoN
sMIEwmL8B3hjwZiJwjhYlRQfEoZ/U97aTalUBe7XkQEeAgYLZUVR0WCHpMgQCnfs
38XkXCq3FV8qxaRs8F6xCYC6NQ0Hmfyn43/Cy5ulP5WeF//dVm0YE4ypdUqX2VFJ
S8DHCVha5wFgb0T27eSzxsjpy4jDdlhssc8Xpcmp5r2NClTYPgT6pIdaQM48LYrS
rZVAPwZXkWUWzjHu2AvaY6p7pVjgH+IQ8oqJ0raH8Y/oMFnRcY1MhdJMYtz1nqE5
VFowE7e42io7rB1M1GSWHo8Pzbo+aUTUh+KJoUDsum/pyTd7gbgrWmwc1zpOcnuo
/8PYTLkXmHGmYVxkjw2vEcSgc2NYYAPQYB1f4ququdC+bUREa36jrgSHsui9R8Rw
gaDdnfGetwjTdpYbAD3yi5ZWujiaFpFV6SOBm6cXYfxxtZPz+DBIOnztevfNCMIg
yU9NzNpIhYh5XU7RarmYVtMHb+mqykBWkSC+5ghLSkFUPpJmRiLtu6oJ4C2O/vII
x0ZORc2O1zJf8t6S+WcV9gjAc6SGxYXx2Mif6IQ0UNb2q23ywUXUIFloUSdQh1wC
pTWeX5xXd/sEAkbhU3qG4K41JTbYDBl8qyYUA6wBj1muNilfoF3W358Oq0jfzR8P
lcDC97yFb4bPyC3bA6KA5OKEEzRxet+6ifaxVhgcfP7Wmz6iUVGgmZyP5mzK8d1x
VY7Qx3AcEVU4O/Pf6mHetiF8DwzYwaYlWTcuVsfjLaqeOITukhIPJy3xy2B1EtLC
MudWeEcYSdwoff4d9VE24nWz4LDajlUXkZMVv1tZz3je4YGB/v6I3qEmpmq6jmg/
RPQQeeR7xKIh1ABA4lBgQE2HsyJehiLSOCa5bYfw2Bkjn+qP48HY9/uw7cY3Wk7/
UDNBM5GT8rqBlvGf3X7sEs5Dp6DKgANkkWDYRJj8Zf9b4aWEdbsnOfobSn6DfNid
OZZcjqDtjduQ0VderyI0ierhHiPF451T5vbFQyv9WYCXbamYNHITBIfB7v6Bzdvo
aNr73eRZbR54GFLYwtVNVRdEPIhw/e2QWuUMOjpPMTAu15mhZSbwi3NP582eow6o
h8dh5j2XLVGrkdDDNEmH8SxgNT2z/JoRA54UXwZoFQM39zXDyZyd/TpcKi0V7/Jb
5XU7fJpuykKU5+oJHX7bzHbBQTxIOMRoNdoJloljhowiwp4N6DazUYSwMhMSvDfF
pfOHjtvQoGnlo83TM2pFNheD3MEbNtCkqufRyC1P2KXjd2TLJJEj5VZGxckcmxXC
kP748gDGvyiUZBcjqoSg3O/HhHs4OBMLTa7UuRDBR8WpA+X7ZoX6NzhNwJgTJQhR
fBHknKEU/+3Q/ty5MJ4xzKp0ldyh0bkkD4r1xk1lGydnijsgdFkMYZhP6zoIckpm
2oq8L0JvcRQUtFQkUgOkQ5+aWhUdsK6VQYlu6e9VjleYTXWbJPw+KlZQswd57ihA
APd/ckurbE3ELTDN7vwTcxy+zZyoDom1zbtqRJ5aug9sXcz5ZahDlBC+2rBgOFzg
iJlbDpoM/8ycmMFGK8I5ZP0dtiBZQ06KQBsHUG5IYUpbwA5o6YsuwvZR7yDXwt3v
NuadcTdsimInSWpbyxXt2eYXkLjyXyalL8fp2NPwQhh9zg2ATNcxvqfotyqK88TO
4GONYX4/36P5Mc4tf7Tc7YGs2X7rwqSnwcSCIBhFoTODjyJqU1OG3BCFaZt6Obh+
fglf5LIijCDi0f4V9f+ibkCFyWZYLAzrc/WNaCk0eExPciVBx9FBD223EP4oOAQf
lFwK+Dq0Ym6aq0dINLlYTSTGbehNEO9f+MqnfrFeNo0osI/Z5Jz+e4px2jzJ+WED
PMZPTGvNFVItJN9TXzX3C2hb5gAgilJPn7W1feh9am1RvDog1ricBR8EXsv7vHFN
7wlxgaaNuz5awrRy+SFKzHVm47orjnSTVvNu2bHNjcnPgZt3UbSjRpOeb6U93nCg
xhFXYGUh2HcQ+hRF1zDy2z29MpveC/qGVrPnjiqQBwUZfiswTtjiOacEHgUkTw59
eVSJnCMaQdAmxXKffVLgHZzMXINOLojkzrfDQnIKBkUsY0YYpL9sybtMxawrLbaK
vaSNx1dArUnxqYmx+ocWzmb4ciAxkEG+A/mFZHAfkpL7tom1bjG1aTYwjsnKDERt
QjZqigWHO7OzHmL1w456ozyiNFxbvFi0eNrg3T0Cr7YgBjmeArY2WlR8SNvvINnf
DlkcoK4T00Ney0HMKg02Lzp3eOcvA3HbQYoY4D0m7frwpR8F3/LMtZnZltxnRdCb
CTgSruaOnUnr9tK4pksH7HeOAbh8zp9zA5SGEMvMrwRBHPSuQZ3zf9ffflDD167g
+gPRmMq9k+KWFrGyuwvXJCW+lo2GfdyNJwKPXumlXXvk+5LZRiL4e/1Uku1ZONQU
ZQfgUBI2vRoV93NEqzwd8N75Vtx+7zMj48nT/eDDnxID4Quf3fn6y7zAnZ4NAaQn
5ztcwtvYpo+CT8bk/giSC+zIL+9LGhyhhnFMZ4lbuW9IE8cIYruHsTfdTzkrlC3V
uDha+Rd5e8hDFTAoe7bv9yaV56s3DFoFJmxSxQY8+92RMjOwsL+g2UCK4/lGUkaz
m4tvK09Zu8pqp1h/iEUakhBXAsXtvlUIAMQCJGEpOu6gYTHoyTP6N8MD35y2Stxg
Ml8gxVb1WQRoVRUnQZmqAN9o3vMV3dKaE4TTEdmzoVCg9wWzQ4WHeLj/WmnDQViL
p/BIqTOrPf72b+45PWfjw9RQ7d7iaGc9p+R/zOxaA+xAKy512CMuzUAZ4fFhI8x5
dmIV+uE4m8TFnWwMRyaTtGH981QgDWeWXXz8rtzGBa7iuPlChMvSrJISOI3y7rBl
5+Tr8oPoNaExP7DTAMD03bQFkbuvv/BYsreacyleo7lgCacNoea3OBC6LUMIjT48
uX/uPgkNyeCBPhUsot02g0I+DB1QH2zbvCqWEi/fO5CcEjyMSeVbTPJtZGvwm8kf
VNBffDno+zVCEiMsyc2SB1th0vpxypoYR07VcVWUBjGdnf9DlphovPCICff7qePM
t1uwUwyfYUr9v2Cs+ogwAlTMpg7OLVeMgBvCls/Wy8rQs/aYt0I1ENb78Kbxqvd8
3EsfwuCzJIQLtWxePN6PJoXtYtKTOSLMtshComgGa0rjbsHsuu7QqltUXqHmjlYt
IQvmW6PArlWLPlIlQIODsHZMqz5htHuM92bjdG5OduqQSnsZHYTODR+srBSTxlS4
g/bfCRniKjoR1Mtjlw0RfSkWSWUgWS6RWap6i1jIwVFdubFg26aW+vZYKIAsjFQu
DDZdLoDEwSS0004c/Giv5tz2tAVbqtWSpWDkoXUEX9YljcTTDm3fenS5JO27sBxb
Gw5Akjdih1sb6oGR6hYxus6oVzo6GOtBYyFHNLYmMCYnYdm08U6FfKqtXG4yeTBg
jEa86IFz+KFRbLFPMJ7xePppeS/hHDdeeSvu2qX0dxFkZdkLbOmqWCLVVrsKH+He
6Bw0mYNa9t0TVdcYmJHL33kicQXB45nVkv+jlTKRwEkf1IGeJ1jW7S+cCd4TytpU
kFM1gBRsMpoD/KNGL/o3c+YoWCZ9eYOicxFsyWEegPc38n+HFIvsGSlVAV9Nu9OJ
AF08karH77IfMjbp6Bg+Y2J11AbukPwf6jCg6/pTdiH+0ta06SDBYFeBkwmAijWm
Lk99L8LYj79behirDe+tGbJCLh7HnWkn9gAcI2eh9PeJ+B3t70r+IqYtKkxRXwvE
h8UtZrJGc9vWXyj8Wt4lgvYtvQ/3JxAH+XqqmHudkOehAtORnLb2liUf6CPr11tw
+mcTdAeGxy9fGg0OmQgBaPS+JIA/hrOUHVSFuAxVl8VSmEf+bA/3HhJYXXgngnJ7
pVzQ2sqYYIjKBRc4CuYC76qse5rVlhgmeVoZ8Xgatc8RTffIYqLvnSRtO0vlP+PE
YEg7kJFYafnjoFPavhMu+fKw4vbWM0crkjIkpTT/g4tBbP+YbJEgQd14oe75RwUR
Q7LXcEupaoqR7V2dXuPA+OAzmdNqd9Xaozr4GxsviRIkxL1TaTRwdkCIkELD+mFB
majKOIWAkh6Mh9rw5h6WBy1C35z01XOWdez6bzOyzbb1MzUkXFnNDPXOl7BXyyzc
ej9rpGuoGSM9FsjElCgSa4uuSz2D8sL7U1xmldpM9JfgcgDxymsNYm4B/TPEEPWg
IxHUNjHj3HB1rmFHck5lwuQmnIBduy8neyj9hcsvPDgmm4bHIJB+LfaEJnN7MXKE
G36g0UOdH2SXbEpTGVd9PGXQQLOXpnegptTOYsKXM9PCLoWvSwurGyOjTrO2t8ut
RUsBd8xnEpTLVowT5uHmcMVQJ1ls3QdQVRLdujLC5PxQ01ss4V4lrUCQscWIsg+i
BNAZiJuKDsGoGYAzuZsiWCQZmSoHirs9IlRNfHTiqSkXs/E+NZGZYmcdMnjmCWlH
RzlLFPv+14CquF6vwMBefeQMKwJpSqBrwyl2oBN8DsCzjLEAsly7fmp2GE7Cld8Y
dsN3wNiVmr24xnsNeqpMFO5TA63GrIBC1i0AP7hkuM63vED9K42jBgjWz5oUi5I9
hOeN4rL82Xif6AyduyCLAvYn2vlfBAtLRfHmdCzaOG21N/3GLzZz6vUksj/isG8L
ihoTjooOHbqJLwMaJ7WA9cKHjsQhM5W1Hg9QsgGv0JHMFc5Sz2DTzW+h2cKRfPA9
9KI6gZ/VQHvUpdNR49V0FaRbUDLFvKpfJGUL3p61emT519HBWbwIL1iAjx0RWQ1w
mMxcX4M7wCnFB7Rn3VkLj47Pz+UIaC670wDSJj1Ph/MgX6eQnpvDYmMDH4A4F9UQ
ytIX+wLwC8MS7ieH8bh8qozaJYRSZOcfaUfHM+im8K8SPRihz0/QnDD3wUMEHkiK
umg+oyivO6tudnwdfpFt9flMmAF07h7JneIGq5aMLoTqgn5FT4pJRbylpP18dmsV
rpFtX8e+sKRyOFMk+k2WYnGaka1qTN+Po8LZhHClM7GJFA6hDvRrTf4yqbn9avFJ
3Bo5KqMGzxaLvTBhoHZXSF4lUQOx/6x2+DPVtCE2VNUWC5NehGh/Sme1EhV5DyUM
isQEn6aIsJduqm+Ds+XMYRv51i0EiXtBRWZU1jcrSZdEkheOd/rz0vRoaxhhb48k
w8nbotygifVZ6KXvDdFwPab17C1nnffn0YOjcyDSoRJSwO3MIweqp7+HyNI/5Ed/
X+Rh12NLssrO6prTcvRpePHRcJJNXWOwKAwqhRMM0r5LtOqRjbnNFva801nNUOj5
zh2dUwaa2xpCimsoMU1enePJW4dQjbWJ4UGtGPjD+du8kIbKIbRTkQCxwP+KInd1
PXeRs2GHCqbixocqn2rFu7mzSg3sN+uH+5etU94FRaqoTEu3GED+/EvEqc1F/rvY
2LMp2V/FDG1JQJYBJbLagfQBLMjwIjXsykYToHzMZyCJWhygRRwcteLLdcWIvkL/
Zv5JzMUeZHbO0vjShDT8h1MZBbhd/OEiwABGLJCP0LC4Ahsc2PcaagHeV4l4xgT4
IyRK91z4jUXhVRiAq3VP8vp5lYe39ATXjpVomYikv/So3pVrwb7pSf8M4ao8zmsD
1EMY8Nq+o8Q8JC4zJuma57MsU7EsvtZ5+voGcZbg4j+Vt5DdHHZnjxmJGF9oLPNS
pd3ecb16t6YtyUk5yQNKnrFkT2Nn12XWxgw2I0n3ICUY4eqH1RFYABSnJogQdBtW
t0J0cf3h+2QOPDWXlpzS58E9B1VqiSkXp0fL7gTh4O3t0bTFjdyn0yQwAXzXYxTw
5elrolVn105GSQENgyLiPbrYhUbvdmlSE2UO8tW0Hj429SGabaW9Yuse0PFp6Syt
NT7LPkLeH9QOyC9tfXFP7LRPJTwmQQ1UftdojJSRbJyulj/Sk+BvxdGWbC/mwDkV
3S4Hgvv7J58gi9R3mnCKTlovUi4IooOVKQuu/pfXDHDQnskJrFc9aCTxoD5QSdW2
CDqVkAR+LVnV5fCN3t5RH3FGGTT4bFhQ74C6LTbhnCsBVHnxNia0x8ure7ZhA4iF
rk6qE6pxeLTaVy1wOL/xiwHuuV6JfBZyHTmnPeH1hhMyIEOjaMCX+z+CV6XBUH1B
jjAMhLN2qmZCzaG0Xh9bRFN647JLeHxp/EZ8pO7Ih3GKGvUyFFt4WNjVVK17Udg8
3dyje3VzcUZceoZ5Lc0d/DoxtQ7zpFUGP8NInuGMe84kYUGNMyV0sexuR6TvyD2t
CPqK9iTg91V45aQNw3G++OJNJHuXtsuMAkIT1agfyroeOrC6YbIztwJlknE0TDct
6aMMBXftBoDJ/WRjGgPpTjjv/A2RafPhmHuOMF8U/UmAshpgiuRB7CbFW4CuF1HO
qZH6MRTHoxEg6SQG8pUW7vj5CYTVEy1LXn+iy384Ua64k+guA4XqmsNnLIkpXaCm
tbG6Ek4rSN8BzCUavqZljE9Dq69wudWCqCI+gDM09WVbLt9XTS+n87d4XD+sW0OA
qEqNbGzAJTeFbGtr4BFElk2MFzutP8K5RjOGx/ZXsH67F0VaFwAomOKPwfxmxEOD
plsfU47N6A4IxiZ8PqVz37gAJYqZuxioRNrNgEJRAFQT/kvD1Ht1zzKrT3MQza3T
ZOdKRu7jkDPdqTYWedB01G279TbU/weS9k2bkmpn8NJ/v/oMbkytTJBG9e1UUVa6
EoSjC/gCIdBdyTIwe59lVLL4MjAnoocdAO4uexZlrXNx3wZ2xkEEJVjgD6p0k97U
uHrFHLKh1xCIMjzaIbwX51AXhJb/rYz2S2/522GGjS/iEYf/SwoalfEFPbEbix8y
XMOvhDZy3oSeYr6vmkm2PV8fwHliwv7dZsCC99GJmXiGdoKIi0T8NoTpHOiAwbE8
+/pzKvhxRT4eqW10jGn/EhGqRlTdQdjJjyHRuvra0A9CpcjX3O+rJdST4+wCxxMn
7dguyFvrtNCJgCa4udeIH/U8kail7BgMMlabYf1/J88S2EULIhEXxKWtSi1aC02H
pBaHuny1BsLmQkKuS4muD9T3IiL/HgSpG5SGN/9CjsNNyYtuGXTqZ+RQF5+xBAnP
+JTt+yav5LOcf+x70HQoUn97EzkqXcH2BJq7+I4aek/kay6sT9sjacRoR4r5fNdI
Ie2YCZ2s2KQWotgKP41/7ml78m2qAPpSjbqcnqS4o+9hbEZaC0YMiKBT+1dd0H1i
rRYy1byLDLHGGHdlZQOpaShyjM83QPiq1JDRWBJeQtqgUibXdUrWClyyMxmFJuyY
+6n/tQc8xJU7pYbvKRbRO0/CQLYHW1m3F0w3j7RmPNLG8kkaaS3anBAoDYkb5VDx
Y2WgUpOPA9f5JOBfNkDtja1K+ZE8xQaHflmbfA/jbcegfty2eR6eds6U2CaGejtt
gQ63PMiFN1YvBiZxzFLIq1IdDKyi0nCja5iAlZmECgFQX/IZXW0Sk8nmB47rxKkv
Zy4zo5nY3ryAnxMKtcz30CRnKGen1TYbH2+ZN9eAEwPOolf04Mva4P+RBBLsGDV1
nfEJqsMf5j1dqHrbKHuwoyrBN0lJvg1CPgFlhvxZe0LRvOh810hDQrlBiQwDQUrA
URW38fz8g99Fonhf3m6GZ1oIOSeaxmPBXcJ6am7iRxv0A1YA4FGhMwWCRiG2ZMFZ
AK8z/tW772A9WwuIKV3oDSodith+N753Jg9QMKULCD+D058xUqU9azK/ldflBvkU
2fmUZv5qnEciP8G1oMDwmMWdYnI0ENJC40u44WtMU298IobrApPHPWhgkOF9w7sb
m+i+SiHKc+CPbkH6/Y6Or248y3tn+z68XVwEm19BbfA1pA3ANmEaN8KVgLSbQG/D
thF2q/tURWz1AXseaSSm4GIGYyQfetS/E49rqw9wmFGYSqeZU/Ji3sjxZp4IEE8S
9MDji+FuJ4iQU4Awp+DZE2aLpxuUy3GK3b4wfhRJYhKnViHh3aVH3kNi09FxnLm7
mgMAOqZB25ZK2KruHuweu0V08U5RkeWfg4EVG9LSNiU2QrvJYpmqgdTnkxalNfXm
Gitg+9ggyPkdxaBjlqJUEwyruqMRESa6LEyOv0zJw8vsalcJjHwJnydVaccE056g
oqlUOlF+utuU9reYzzpM94RsrGSl+6pA//zVlTFVBIFbxcDXLvUUSCN1H50SS6or
Lk9ISJTv4MRcCFA+mSmqHBQ/AVH+hxYVQfOHy0WUYqLz8LFOsGJM4T4a1AN3N1CW
wM7wj3yk/8mzi3Z+hG1F3sBChJrFPRSMbFgms1wi4pepyuZ9tUGk6uWNUUIsKQFB
r1XyNdf3X+Y/weuli7ZcwjyQNvMrBT69sEZejV0INJTL9d8uhkwoHN5A5u89oGTO
wyZBQCz9dJAmA92rCKdkyQEG/4AsApGO+kgDnRZoeiqYNevCGvsKdss11ASVe1m8
onsk2lfj3lFuQq3zTrRvQ85ZFqHJdUesR3k5B5nfXiJychM/d/pzPUL/kgXTuEBc
y1XQ7to0+hvaOaQCxDeVjUY8lXTmkgZHypp5aFWTVIzpJ2sDQ5ywPsvZK400TVwe
mmL1jJBD4iw9ksHk3CAtA2qZ+YmNfOB5imWqov0SElkmmupLPVR5Irmfz8RwVNTP
9GwGvwnsXc+hIOVTRTxeq3mvMB6vfIiwXo5i3lg6v9pkDMEwrbBEZv5WBpR5Yjz6
UcfITXCtX0Wd9PeJTKvKbFaCGJi0fVtuulji3geuAxXa0ZVUDVjSA5QAsADFcjaB
AwNc09YNBJQ91wxypTWFyhlXWZtQaIzE7C2p4UG50Iuv2HaFSve38+bp782hfidq
6vXjlcxPFT98RbIOKLKBuw2iCH/ZlzLcytVTIgfjBq3LLZDnjuG91YpMF3o4TF9g
HTvHhRbFPb8i3VPf18ZwZosYAe5U8Nmef76DWgzyuIjCX0yP8wovQQ2JKGAJjMgm
dthk5PbUT25mKFeWdNsubekm+ZEkxrJSEgyL+y5QKDlmEkSJ8qIxWRaXdDDRKqxK
HzdiRQU5oHTK8Z1iZZ05Q6KNvlDw2T2YiI7MSBvk4ma5XqS4s4vX8B/YVAJdmhB6
tza+kBE7p+AI/Eo8lN5afXuLKJ+TtBOMn+aL8qKrQiBzaR+JP2/HpzOTXuxZOBHZ
nE8WqDf0FKHT8Kr7CSc/0mH8b/3gS9J+v2VLJtUjl/Iq9dQA4xYTUOrCmLcAs4Ey
BPD2kLuv9xzhp3aYWin37hz1Fd8ePQZP95XGbW3lxxIABNQz0wqCZXLG7gwSvuh3
7YtDZIyklxjFxJjpehYHzzx9z/oFU/hSSLecjEuT4o2wJOQiUaLmECyFZIPIrjoA
Zm7BZeZi5layQW1CHoCx39KoH+aXPoQeEDdx62C+mrtq6MvFLe/otraQOZ1mznnJ
H98Dkga0+/zEA/Y6eoGk5DdveNoeBrerYeq4TlcLuyF7JMV9jJ2KpH5S54fTAli4
sAMrnhfuFwISHArjun64RaNbsCXU8V/U6M7+b08vDjAlifEuYQioy9i+bbnamWI4
sZzJNqG5g/FzeLJ33ovV22guNCgrI9jsQ33DHhDmnm4fjhk4UrWbX6hm3qKdIw8U
NGv6cbdIom6Cpig/tzxieT6PGFlMrQkY+E3pg2d2cS8jYWf4/5nPO3k6P96QtN0F
de08sjiAhz5r8vk5jXwi3UKMKZi/CT7nPBqtFktKZGMmiQ1CkKGlwDeBMg0Y3ctk
133nf4aLhrLeNGKbJ7uC7VqU5Te/SLiNE4MjXEbHNzUTbZQA7At4E/NvlPw7mzVy
1TiUUa2q18z2q+krM+K19ZJMEI9e9PhxHJCfYYgJKwlNnwZAwsus4iY8L8AuS+Az
EFy1W0l1wC0xvjMkSNEctoYYrYAIPwO43HGS65ErsSIBb4NOgaVN2TcZLTQDv3r7
Hkdy8vPdMCeDksvkne6cBZ4TfWHQypZuOS64kUnLTbnSQdkUaqFF5eq0GIa+X3YJ
Oac14auHRN7cKsz1Rt3r1X5CRZIcBGsoGEWxw+pRCFHvsqmNlid3XTXyE8aY0/bu
eJmxkCJ1ysn0EYt0yUKLt4i061Qib3T3UCzLmJ9Ey4VRO9bXtCQcn6k6vPh2ZOk5
kPsXiguGOZ6FEx7jYkL9yRlwkEj0C/V3JHzRRmpBbxUkniMrLde8lPdLiZfxxp8v
WS2EA5NZiNp1f5OGEc2IdX2XrlTshaGIqOju/MzHouIJjxrnchg+Ec2LXzKMREVH
Be8l9BeHw4phHysRz7j33tJXgHa+xV+SCNgAGFml8/Ilqb7Uyf3wHRQSDV8xByCd
nhk9o4PV0A3KDVHcE6YGtS4zAaRpFY/czxPvj6ac9vu6vyvZB2Z1zEZ33nVotKBP
KNVNNYeW1ooOqpys62OhdStY97QTgEmSsVXFDzbMZHBow8kTWAFFxgwT8CX1uFac
8j+mfrYp0uKLGXaFP+EPxFfxYyUxJ9OjuRERVupmScgQgJnoYHYIK7hQkvlWMsul
lsXECaZWti9pgeHViDl59Lkf2buXIVLOPBeIWPWTuZryxW77xsWre9qGHUpX/BtS
qHK7CORuobH+4z323CL/1dt35Qh3IEQuaehW8sgq7rk63D7IaWnYXA9K99S8wozn
g5IHJE0v93RFDxWz13p+itzB6j2ovkcWyjQFYlTk7qIExLpDIZXGQH9NkjS9wiaP
HXI5cHpUfwEoL5Li0PAaQbtf1Aah0h6b64Hz1MsS6fk4BOaQXcNpy2Gs17aTZaVo
l4Po3bUmbK7j5zD3ktlSU5UA7kvvGQrdvXJudyl0tI3qibLim9Q37clML0mqimik
L5aNc3RE9z5nRbtHoqGebz834SeNGySCYdNPHGCYZTEjk9aKHAh1nPqGl8eE/u0W
8n33Vz7Pf/lnp6EUeqnFd7Ux7gBVi9EHUm6fS7HoRxnt9gVAGPqMeMAQfYKDprIM
RtwLCIOxrgYAzejor5gS5pT2kGkADYZV5dNfjYcM4/B+pMknL7S0NBAHqOcoKWxv
rQi+d0Nhakc79nBsRfz+F/mgKjBUFaYkGezHHbQNR4La0dX94Iy9W4R3Demv7/3g
HY3mCTSfWWS3cumHnHSr8lZvJdnae9ej/mdLj6HPGXtMpd5zvitu2GhfLbRWJoTB
VcmyClcWJ6FLmOJzEezRu131N8D9XAKfSplP1Btdtla57pfCQjiqHUqpqeexE4MP
RA6Ilnhs2fRUMHGIM5JFd3QAw5ffgpdMz/GsdoY1dT3c7iJXPqMHHQuoArmyrG0s
S4IzbALFvD7dnpeDg3l6BrPv0asR3k54QCBiW7VJKoq6dRDPylzHZvtp9valEZKw
eF7RXN3N6IG1zgyIClci4YoN+Zcl2ARZs+NXSyT4QzRU6/Si5KVpsIZDN4hJLGsp
q29JQnHPe0LUGhANL2Zx4EyYhPlmDY7Xg0FVAcDp9DyMesa44+3BDRgdWW0vnP8g
voIv7BuvcSBJnsUrWPtrISk7QaaY/aRf23arOdnQrZM54nkDLcOEzDAr6QBNP+sD
1D7Is+OnuIdVGywhod4r1ZLYT+hCr95rC3hTlT8qwQMoEfkG9SdCr4b8Eq4h9RHN
uE+WvhhUUEaleHtEiVGGIbnyqwTWr+c2uGF6X1nOoCK2ZquEIf+slIw5uws2Strl
dVM+/1yNe+8Li2M8L1RK+RfSB0+kCqLw2bIuDBBLD6vzyB/Ni8vQO5x0YHKsJN1E
DJl7nq8DEcpo8glQwyY/l9Bf1aFeewnzcWwdeImbE4iZVzPJtKopC4wZrTEOwZty
KzOlQPgYB5Kxo6VzY5OaHXhICt1yarclLVq3qNyhecV1dt3nr0lnVklteAMGV0FM
je7qcE1K1SGoIBTXSr25UUcIZaEyRbaCP7dJpR0dQZUz8VVHPMmDJ3WD4HtrQS8j
2VVMwgTxwwFgQ1Na4OMD+99znC8UNXMRYBHi7ulFGozV+3wo0+FOyKzl2QAQP6dF
4Y32sc53j3vPpsiA5APqLqmfkgMcF5zWUoDtF2o5dqdRovMF5Xt2l2jsGc7iPKrk
f3Fm8WLz73aZR9xCqDypZCDZz7i+HN/lhu4tBBaak+QmUWTMJipN5dfHiNUTc6Dt
E42SmoQRb9LTtg6Cr2mux4rmsIkIVHfsOF3EuY+jXSXtWGcPhx/s5nCzqXP+J/aj
9jgH9LMylywc6NIl1jo+VaDSlpCiFhm/O0/BflHGvG58xFJtqRRn5kYmwDqLGAXu
6Hb9pwS+YR123Ju/0gfjkdO6CNf0djFJtNsGIcrA7o/M+eoQ1G42g6KEYxTZs5TS
iWghBVXHP0Stmg2xXOFsD9qZzi/7i8gNwL8kJVvem65T14vWAe9Mn5XMpCfzMxLs
x6DSojt+M4DSh+KAJtgNXx/w6iRSHTKgnT3cXN9s3ktrAMmPPpEXZxedTABoRZsr
9w+uBxmvFAxlg6XrgAIbymqsLJDmGbQd/O5JNi9sZRR/y0o9CT9Xlzslf2fojZ1+
JYaXg/4WYFvnm1ShXUQu28EeglRdzXBtSYrJn3DeaH7sZzyo7EUIm52FyijWQLT3
YiyqeCKeJNYBXfX9KEbhO0pOXiEJsWz2B3S/k7qoructAvAi9CviYLDepr3P1nDk
Az22PrMHUxxs2vzRFfsihXmqpNmvd4sUA/ka3ayyr3QjHFRQlzDAVGP3hFwnBvAt
n2jjYBDcWf/uZ2iO5x4xHWx0WJm9sD/gmVivx6VSpigYKxdPqnlM2MlUTk0QTNWq
QIOtrbPySevMvfAVX2HtZWCZ0627bdOGfU8kn0eqex8jcnEHAaQVY+mq/TX+qLDi
HV5HrzQlwNpbD+/c5j0Bgi+7R8qA/Q1W/zUZksUsWDZkDr/uMTsfqmShanivOGTp
6u450c+OtvcooN7Wrfo5VvEhjQiFncZBhxInIsu9x4Angnccp7/uwApbrmA/8uvl
ys2TgIZxv+241GQMxJN88am7n14xoQtkMiLtH7LqgbQtgbGwir5HMgitv4t7Z5PG
sUXeEGFCRBRKwl+K9CmTlcULimD9cNuXbc4Hy/gRWrQceEhjAsUozxfFruBCxg9z
/JYxZWx8HFH/3aFP2YUH56SfUllHreHovfy3IUeZF96JoYH9ztJNNhPGDurj/1Bh
b6ILdbSqlCYMQvcbY4EnnTjIf+2WUiDGtk/LlcQE2kOvMbX28K3eWBC0xOVWgzHz
v22BbbAJe5e80pzHarq/cR0H0DpVXS4JRV3Iw1ATx0fvRns++RYDNTk3dMvUM5ov
+NCpDj2qkMhZk9mF27T69wxKsQP6Fyj5qJPB9bRGZppdyjq+Hvtx/4pPSP6Rb0oN
qmeP4eM1r1H8pPfqIqI4d+Dg8v1+9N/4VuYGTRUAHiL9RpzC0y3WISqjHpdngfaN
yt7jc1C81vlcE0obIggTLSwv9gBe9gKl2UnASMuDFSHBrojJuX08VmDqDgz8uL6o
TzL2IgcF9GnCRCXOvMmOAKgxOFcNL5DUtQ8JP4cQg19avGxZ0jSDKPVrzXW+6Nfm
m4kFgBAk/vM0KxuR8H+mkuJDzxeHyxCJGhD2j8fpKzKg1ud8y1LdgfYa8nkW82ot
PUHm4THyeu98S/qy0fHS0XmX2c69v34yOWAk13BUUUXC2lrngqpFArsxmY/ZGac8
IzfPwBp8h/YviiaqoUemLvIpOs+EN0MuXYVR2BX5n67hGPzIbHqWoAQYsQ97Vafo
8C4x1a9dfN5KDmUAJUKp9ZkezMkqw0DZl2xTXtzHnTZNvmaC+RscX1yGGCdBfdya
eescBjehivdhPYU50Uk1sWp2tqsA6uS/goeyLulJlRq3ZICEh3/efp2Up1ABqCFl
OannGgeQcf3OZZqxtmtY/dTbFCWEqVm3UGaTNRWMmwQZK3RWo86AygL5xt0dPAfG
ap1ZrmjUGmo8PAs2ieX/mJqJfxcgJmAP/JtzgEFsF9FoebfZSmCRE5YaWS66glqR
LAH3CmO464aP8EOi0XyiawK92omquEhW+rG0OxeBkWSZdAMK/chPe3gs5i7wcpgz
RfAzpa75ggDlt2SVDrnNMuioRh41b4pXytP69OVGJmlC96BCG6COIWIpPO6DqS0x
/x1fgaRVY4dSqZq19V7DuWSsbd1qM3d3jpgr68okRkGvS7tto5uMrp5yNo8X+COM
wd2EfukMuBnShj1Wg6FPBxt53xSSU6YhOMJ893zr/+s2Z6YYsJsSCU7djG1+1MiB
SQR299/ZlBsgaoWWepcJtDe9VQo0Id7uJoTuQs8Sz2QLAY8rDzp4ae3eR2vxYbDv
ABs9nJZuPWXeuhh5yI6sZ/sLhx/SmlUrdDgWe13p+02UVZ6LPRkl85lvpSCryBLf
XXfMHCJl8X6+WXGT0cObWQmN+Acn76KC3zF3zpR02BdEFRbR6EmEaWIwWb5mmpzZ
yvtb3aUG6LBFtNWZ9UrvV3XnIEJr2nGqWhr4zwGZaUS3nJax4ZCRFz0+V1kyNFWB
qMj94wu025iH9Z3TJnGvATWSesqszus1WUAstv8fVAYK9gQoDa+CqYBy6Ir4fJtG
k7MrairyCBKzL7oClKn7g/0LWvC0twRe74sCduvbqvsd+kqAW+lvTCjAwh7pO/13
DyqohStp0cnJWbliNqM9iDBAIyPa3zwVXtfQjiQoNp34ct39Az+EaiFOsjSlpvUV
/OxeM0uZJBE+DaZZ7o9dtr4YH7yoCf+CGybqtTgOgUqThwcTr2j4POSpR0acsleI
lokvaoeUYGgrZBq8UkhUXujT8jlVoz9Qg3ynEzhojQ0wBDsTGrnnAdi5uuq1ss77
ZVLLcrUvrNQxIpErPTyI79c3/c0vRwH8Zhm6PDXrewZ7DNMEn95kILA7xTPwgrQF
JfRMdaxSSg2s3E8NDpEQ5B2CouH11QmBebZHAzjVxU1b38CqNSYROKNVDoiCRXP0
UU2X7wS4FfYM37SIKdqSuwTiBA9uAzSkY2esOcqCtoCvieZFld/4J1+iKvTyftx5
1OyMsjW433j+Mf9Aqz20yq9Np+wr5nBJwDg4Her507KqamZ/KofisMn01FPhrawg
e2lmEF8RDc5RQwMZEoURShDCi9KT3xbMVzKy8E/GFKcGT4hrKqq9lKB4oz0nD+S+
u1L2MpHavYbO/HbuGuwdwdbaXnoZ8GiJImFPKt1iYJg//fBfHsjig6tfU0WGpQUa
i2ooiV9a4MfgbEJIGNMNcv9WZsCnJZ3OZwEnThENd1aYXlsgA335W3RpGFikq3eD
ZgIM5bHVZslBQ/GqFaP/btIJ7P2OA14VUos/Ab1gjCG8JNss3Es6teYsqeOPfRAY
qC3CY89cwXbIgSUO7r4rLl62dsHr44qt3XPIM89uYwnRqOelIwr7kWegdwUWOVIz
jdktUpp1XP5pSiyj84lGr9raDIkaMIDBlXAxKa/lyM1MQZoGq4GL3cW/4HMcnYmM
pucZxWGxGaAugBIysngyQDIs8pjuQhjyZtSi2EKZqPmdVc2xLxN4idMMvOoaGVRG
8ioADSleTo/HRvqeUbSp6wQ+zKX90kyc5socBOz8TkSXHl2HdjG3TrEIyzrqBTXK
l/qSNKwO8Ey0O3m8/AS9ju5MMU19q3+8w+MQK6iMLeXnwmONCOCkkckmTEyNfYv7
zfvgkvNtz0NjVYjtVTer0AKACPu3xo+clkI90c3AF5T0cmBM5n9PR8uCKdIfxwht
OUD7HAGikNM7ZiYQ5V/0eVkp8dCFds3Z43KXIFHKDqxJGK1oTk+m8llc4zEFN3vf
6i94cn9OAzaFl1Ktb5g3jiyYeQf3CA99+Zp7HVmhie1+XbFhjFp27ppYudfdZMZc
PWbe4kmU/BZCI9zG770SYokbohST6/wc410rv8glDiNq5/F2hSP1ahGZSSQQJZP+
5yxb0bK/BjNeiORhkYx6K7kEDhEbTVgSMg/yKWvzLisHQQK/aN6D1zUf06LCV4hZ
yR41UgAeMhTF8tPCXBOuqGvFULz0aNhBBLyMFTxZ0qXcXUBwSKv4+tc5fEepgMYk
avA4z7uHQtwhKWZftMwfX4KldNyp/T6Tfh8K3g/mAygtpb69jXwo90z07B4ftfn3
HO0QH54g/B8ExYHDO+80cfsdvpZ4D+JNJxHqK1/h+/2JiNIx7Dos12U2p3VRz+jt
aleSIUuJYSRAul7ADkEGey8MFmHaGSR1CkOypjGGrMLgBiuyEDFSaNKaZqguURYj
kHRcjaAEyspUoo+PvNsNZqiBlUdg8oSavNkGDuUbG1EXkEDO+eMBreH7on4xz2X7
aeAxRSx0k1rnemplX6X8SC2mBnzefxiRJRD28UgcAOZzmYIHpDJ/wVfrp0xO6WzC
M7CCpmYd3t77LqzkTGK2yd/uSrYYu11BobhoBxdWrrxnboKICln6y8IhO9vEOAy9
pBnKQO3pgMgcVZVNpsPueMmId43ht9PLi8SCiKR0BfaP7LCviRE7KaDXbE3m4VfP
Dm1fi4GRIz3mlmdqdAUTGjNeo2erjpfo+P9XtrQdlQI7Y+Mbr/iJS4fyZEzVR9Eh
qmJi2g793iiww2uOp7ExduI3ke26LqZ9biR4v/dznyzNoDWEyXvqnjvZjobPaKFV
DLRRI7KYW93L002DO8gFreodP/hfFNzDaMoIIrU0c25l3uqdJFyRxRoj0MpWi4Ff
bZqELDrEEPwdMlty1YJhaAxk07GHNhfMWfuFuAtF6dkGz94UzrFUlX77gA9LUB1F
V79Btt15T0750p9adXoPu0j9jne1Bt4XKYV19bRif8GF51j9ADKg6dmIWujlSUYw
gqj3O/cL2AqGHBXzAAnZIu3GyJNuPhERL1FEbuirfKeL8P0eucmRUwWGCpt4yHif
KLK6bL7f0mRI6V+rWK/jA+oFKoCli0vP4DjvPEW+iUWCR1lSdkoitTNIVvPv4txs
/Byvj5+bw3iQFurEJKjna3bQETFivALegf7KHNgOjHzkDvg/k9IGXVjMAhmX+vma
0E1W+wIjD1opT9xJIMj9RIO8HVTN1lqSSrHTpb89M6MnGtTsK+K286/PSGBsQ1AL
w7G5XMHp18PZMyaw2MNXuqiYeWUbkuBxcPfUiNymrTCM9ZwfsUR4LQcNOs8x7paG
NlOTMx8kacC27MDooorDZ/tatxk8qCHNG2QjStZfByYGwE9uaUpCpaGD/HinKjDq
tRc140SyyA6tX7Hypm6r3Pdvgr+cTGwcPIDkCqPJTTCOQrpCKV7y8liyfiKZmbLG
bxuBBL4tqvo/Luy2EPfQEwdoYST1ktM+XIcHfzdGGChrI6N9mBRarKcaoIf43Ae+
pfhVQrSWhh/KWV6HkDOe13NMsNOq6MkS0k6R8QucJ2D+tsOlkAG3zmDsNqoC2Cc7
zydg9FmvxGMAeGU0E3gffHYYTU6dywU/88ck27E8OwJTw6IFYZC9OSKulSbVEgs0
EsGzVyU7dzUbAmnsKffjSy29oxahspFO7zATJRPnRogRVK+qmsHr7E77a+X4doAK
/Z01n+WPHq4Y2hNALYq9UZefe+aT4YMOAgMn4f/K8rHXcMMcNwEjVKTdmv8h4yRH
dRi8OZi7O1oqwTNPddDouuLwHargnITYYAEdtMw9pRHyTqTtSbzWZwrzzfqo31aW
R+fX1AcEF0KvT/PSuMchOGsmqTe0VPjzSdFnOGmjGwqidqMUrPn+zFW9Z+uceFn1
z6FPrF9u6XgE1suCchKgUUF0TghlC9FRJxEnK/d+vCaUkCZ3twhOiYJJMqLvcpaK
Q4u1U2lRG05FmZVLPV/bmBS9/iQDZYpsqPAODd3014VTmwssW1ERDzEYsoD4ezdD
uxfo1ZFfYZNMDjBt+12VC3o5bC0rAZCobEw604ZS5+mF3cqEiwYr4pCytMcmIPhR
F35egFd+t3ULyJF4BaaWznmosLMZKuVa1ZhXa8DcFWFJZ8AV8nTHrSs/I4P1QZPm
+GvNzWgXk/oMA9X+dAt9rkQ1UBj8iNybakKPH6S4/C9Cx3+TxQjq3eZXWodxp6/r
g+ZY20+kc+wFLKA2EkkuWWxNfvFlu9H4/dl16kxgiU/vqRebMicACsh3tK+FmdSL
0qhz8af4Pe3nATd3c50/O276apMrZsLkJ1clmsQ6kMnESYSIe5PCSRG2aQEGEglp
8Zn7tYpeRr7iqB3xHi/oHXD714w0PfL0mbPtiG8Y2u8osqB+bK4kO/0Gob/yaloE
i7Kttm+hr2LDmNvxxm8EVEX/kPYs0ONNaOVeL/jpFecConva+Os/T2FmieurHLeb
NzFrfrw45Rb02ypCLpZV3MBR55Vin6iMal9La/QkP3n1uPJUQVsMG3cVKesEOzlL
VWQopOWoiyGjaCFXcpR0bUQogWBQtX+u74XvNSkZtA6ZxzcxRcsP5rxgsfDWjmAZ
5+UlY1ix3BwBNTinp4Xque4x7pMKWH1iY+tkVZvOh0v9+9mltYVeyQSsuw248bkq
6RcjfIbRsgbDwtUURxW+kV+/Qy636Z2MJUztShMnlJHUnCEtYfyQiC1qmM2M8R2C
0RUkgiypiJBlDnUgtjeO1C9Ar23wCBbGBuk83K1/ecKmtAGHcfIcsF1REFnlbwpb
C/fYDsSHhk9N8vAezOZUS38skmilKJ3yAPSrJzt9xVFOj3PdrmDGHKoPFI6EG4cN
RQ56UJ1lZgph6RmFyHMh7+hFM/gspgHmQ0iZBiGvhb/RJXSnqk9ZArxIlfkhX6v7
MQRsLkpkH9vbCdmmf6FD1xYJHqT2d37K1qfh7dml0uFL/NOm6RqYsKUZefDyeq5N
+Sl52GXaHNJKg9Fi6DzyVUst/f+ti4Jq0BCFGHdS4rZ7oxrr2FHZqz1uPXvEO0AE
edQas6AgPHv01xWIwSG0OWtkWcrsQLLQYuzWycG7DnN2JGWkdsDMWOPZbJ19oOTM
Es82yVjEOS2yNcXxO/0EkoSdb3dgYOYocfF/t7kuBY8TWm6JGyKaQ/Hpx42ikZPu
oOwVmWe9XFOeQpWfTHv9idSSj1LMHwl0xol+DjdMZdsvADSisl7/kMqkmSJIktt3
G6FzGhyxA622LlFG5mpJrz8RufGY6JBaT+H/Zwu62gg4ZDCrsw1ayl2679lAklu3
XZdVU6lOrPzXG3CIElxLf4q4DPryB/Uur9Zz8BUBvy+MomtwLqOw0I7/AyBgmjMx
4HVsE4LUQ1KlXfCnFGVzJ9KnQLvdhkqjEBQTbtsZOo2HWDgWzfnp4Ez3f670C3Sj
+xOhpudHKxtVT0dP5wdLwevONuNsn9Lv8dky1Y5/SKQm0m80gEl40ORhZ0NAqh9D
o3lVsMk0IVEoKU1xssGETuY8wfTBYPW4n5HccHQss/d1rnVOR9eBxLhS8RtRnhUf
MJk+oj8NyA9+Qi6Yrd34hPXHH5mXvnxUGcoMRWe98NGAF/jm7GK6F8qhg6Je1SSD
aBhbVb4qcDS4GPr0nSiSfep8MmM7WnHkfMah4PZWofegjOJrkeCIg3jwVC4NwBbU
+8FCEm4jZIK6jv9czb5UVrfKsX4zrd8eYO74bbj89fvgeJaAkWgylM7rKTdS6Fnn
2FbSKtzZqoxRoaeiOsL/2iaOwZbIwpdJH0cgf3D91TqtgZAd2rI1JuM4ig6jyv3Y
L7D799kH0g9xCLi4tJFJAb6FTmrG+xPQhKWxRcY7yjxs/YIjqlVpozBXHxaQQ8fW
1qnOOAhdQH2+cEqqD2qj8s1w+sJ1DDmiAz7aoUTVLryI1utRIcFV4bNqo7z4s4jK
Y8G8H5dwYdyj5/urpGR6YjseFkghAbJSNA73GMjHB6n3xWo/2oVCgJs+Snak1e0J
K709tTCY/eTQ6ablzdw48O1ptEUfJU3RpjJGkO7WcbBWQC39pqhkX0fMtGZE8J3m
r1HbD4VtBOCrw5VqwHxtk/sFLrcT6hnKt/t34afiJ9vNYOX+ugmB+7Ms8/ebDIJE
gGWCHMgBaWepCBLE/aA9scF1ED7Z+qsQUmfQW6MJCpn+ozgRuebex+F1NYUqOO4x
OGA0GWg/GUSdgNsr2NsUCpU4zSnBZiABYSSU5GLWbWiEzWgJTG2dp9h4JOuvNBHP
qJEWONr/e8xwavxv07xUlo0mJGZ9MSSlq+5CoijzP+9mF0/Q6/AU2ZmpuVmfUU5A
O+WP1CavkOLfFGytxl0gIN6bz7B8nNqUXadB5LozpM+/vhQNsudYPNlweDjQ5sr7
HtVngMIxNlCCx8NTIxD8UFQUKwr5zOGn/31cHKzUHDAwfZCWRtKimzpZi7zXYShE
HMcD31d+Yun0vMPgGdDqKRBYSHIcI+pPkHLDJ1RYeW4GlaU9YIt8hg0oNmbTf9d/
hOljfilJY0ODAevtUikVUuyo+vbcjuFu5PfANCRWXj0KOOkvKDuTWt46Wn3imfrn
c1VWK+Rxs25MFIYBi00/NHBsbyRZ5iJGgaOJLRgFeq9WPVfY3vD2syeYuexDhfkl
VThPrE+4j4SPEIhNIcVrovZPmOjIIdEvdkXODauX7BnwKhCLAEmFlUgvXvDhBspW
bG5+SDT8FfGpyPXnVstgZ8EG25UxwhBxMIr4xGfeSIJcgkedZVe+jFjoovAngfW3
IUMJeSk55RRXJGzk8lVNzx7nqKhp/u7olRnqG3JDzmNJFroxPAmA4gt8g3GuYmb9
wr8WMQsVk7GYt0krilKOP63B/bkJIt7uZqbuBnqnqz7209V6WoHZS0ET0nR81YLQ
JtSVTuj1EFN2cpLOCbSAISqyfcUmfRnISC+ikPGVB4OV1Di+E/QCGG5CUs+jO6af
qN0jWujT6wqkpW0uwXcJXTCXn+JGjzMX3hxFq+CiJZ9jOdufYV5zyPJWtiF1ieoz
3Mp6yWlTjhjNovxXF2dpL8h3bLnnDo/jP3Seyl99B/wBp+mPzSxRcLaAjf+4GUov
NWPXLNIsSYe+oPPT3TnwH4IjZ+cFgtYkr3+3M+cdqjXoS71V/DS0AtyqZmdKW6Vs
x5npJQFJmncqMGaKbC7Fj6h939sb6Q7byHLpP+1lSsZHTm4cynXxaFYp08vHbTIg
Gg1D18N5kndVmYC+A4rBFC4jW1RM3gWyuIPQCqm1e9tm05UQxAnWEneDAxraFkkK
of4lqPsF7BsF749rrtJDXDjF6pBPGirhfqVVT6qX/FEAOl8z0tFSG6AgH1/QCHua
vhxduHA9StbBrYRjYyYA/u+MLeuYlHfhagVTUnMOFBGcsqYFiauvn9TPTeqOpDf+
MutYAIZ9qBI6yoHI5x+vOPW+0MiKR2SsCMpciNNBui7kWOfMuSddCtIaLG+PgrC8
F9AhZKy/SjnwTlONJN4ULVWlGys9bxDG5TF4H1FYPhkfR4jqOqKy3Vy1P9gcNY0/
vNwOeo6TR0eQelE8LWmSB/Qh0/A69XwQ4zweTeJoJRPxIX6CScSzxeVV9ljpHxVR
WT1S+K04DrILe+QG5NGfGf4VViNUAWHbAwUx08+AWcUoHZV5AVZeD822FOgFw7pG
kXgkBUicYCI0D/rDvp6rFdjF+6H9eZ7uZlGp3+IfvmLBXZue4RPnABiEjEAo7afa
wJQkeY57+/QNXdO2iTdDfftuD9oRtERttc7tqVB1uut3QUwS8/OSXTvDa+0HYyrp
6oqgM4oXhqFplSuBaeyG2ovzCRemsIlaTytbMp+IxKnRz+mJESZYY8ET0IPxFAkn
12ZJU/MQxiMOKg979nDmr+jGL4mciwV690tL5eBC9+lEXC5f9saxGaNNW9W7gYdO
AUGaYBA3F3+0nV38CsQZmSPK2xpTE+l2An5b4vg+I8W9TrxIqBtXvXACJ0dStXBy
guXCyJeemR1B5KljSW+XMqM3oOyYD/cF/6SYVh1HZjxU+iKJhf8+SBBY1Ejledvb
FlyTSL+ze3N2M7ROcXkMN979XuieRWO7oLmpaKsTNkx6PibAPazDYsHHLaxlAuC1
J4CRfT1Cwjwk3LDku7qAa/Y0mRemRfnqKPearNSnFVg8taZ2UKbmNt8x3NteM5GL
EGjo/RnED5pYpZcSYHZDFcZB/x6LhcOASaNdXt2ISd9kQYzW79E4iOOqfMPS6rGi
BPH8INHN+YAIfW+kbJaPZDNKHQX1TwiwnvtU0sXcCF9F6f71y5b2HH0fdOBoKWLd
qYaOdr+vbBChJeTis6jRO0A4Guuz68BUZz0PBkfZ6kLtqPjhrWZYJTaApftr+Q8X
zpRxIukSwDYPsOoiq0I4HEIoI/SvXCOa3nOd+MbiNh+01FLaHAXg5KjkrORugVRy
Cq1osiBr4SMuUn3Swusniot+Y82wB0SsP4IhN01MqXrHaMX91TcQ6zbCUl9B/bEn
PEjGI5WuA6UhqhSVl3PpUTvCSUHCkeIh58hAfOYU35BADPuFkyfcYqL67Y5lDrn4
vX5DFKy2pN2h6dZ1Ta7jpNXnPVJlsNhpSs+THg5MnRe6x+ybWXqPH4IIf7bZICkX
mTtc6d1MqNAp5Ogilr+tTG9t1y5SBjVdx+hVfYH5kyn9L/mA3YOa2SXp4ks0E0eR
h1AF9xEq4QPUtEe7JUhkP751P24Ctg1znwGBQ0KQ3SzdTFUpGt43VzhH2Iw+tE1O
nw/eY6W/QFS4siznqAjKMHCAvP7pGh0Zz8M9eG20mg6XqV0qP5uf4n0UusOs75dc
C6DyETkb1k8DsvI8x/vtBdb6zBY2izRrXFWk1bpsnYazR5jfuR7wbzbLF+sojpCQ
5Kik92Vy4Q2jRfbC734G20pWZsbzMIWXIPQAMawUSsNdVFO61taUe92ld+8RYpnU
SUWyvjP9MLMQIMD44HLI88dOsTG6slgyJ8WSIwgurwtn4dUttHDijRpp3Nkx70K3
6a6mWkqUd/m/8xAQlh8KtR2UPSfZ8N5AupaH8IzT8+Flc04YrXPg69HWbJQn/0oz
VGPDry63ZgfbYmxUhNRPRGvCwJqVGSjGbC5P6kE9RjCoq+Q7E17KpqcgRqI13iGc
g339um91athlmldQpcdF4Vkx7ixnu7tgn/9K15AYi7h1NAkj906cr0rV6UKKOzBM
W+WDv0f4m0J+EmoSl4u9qqjiNJ7+76usSemrnK3YMtXItsv9vTmUwF0bn3GFb2MH
hLHQGkRxi3kZqJWeoNxhPMAE6VMua9S9HvtwcdjPWkm3tdQUw/GjHZrIfv8y3EJw
pNb0DMes+PtuRwttibOcx4LDIsD9BerdU1R4Y3lWjXvtKOCA/LmRiFH6pQ3iXycS
buLx6VYqBLXf/oRhhp7ig1YgtMEMmxf+lxV6QuUmhkYO46fYPeI1kAUAEWIzqxOk
s8eO/wB31mySvBLxyc5kTNCE/6M/CCdbrl3hRvfLBQ1dhn2tuTrreIa/nc0TyVzl
rPBHsFCprFUJykw66NZP/uSHCQ2QLwhGy1yy8RGV086bz5WFGiH0DHzWJ4IAYuv/
NPzZRHIOVvqncm5hev7ewPcRB2oY5RMj9XI04Mr0c1rkgGnK6iGirOdfBf2RdR7m
RcIJMHuAGCNUCNlGV3jiXzo1+XzReXV1mW2gktqdVS91kZtVYkS5xeZhgDxcaFsn
y46QRqUMKf6oufqVa85A7d1ANcEEAizETuqHv0tWP7H8+SZdtse3vhYf9reUr8Rz
IK+za9RTAvxOkl5aNCV1j+A6Oc0mk9wkKIfRjfc8Vzcyh/wDWPH5WYhCMJnkJSHd
Nn4YxFIBdeTys3mAkNw4R6bdFe7qhyJY/fTgdQntEKxpK3bCXss/2ZKk/xo9sOFN
95jgOIpzSROcx7PhsdJRtm7cPVAz0NPW3UeIaJtbiukupyRfJmfisEKgwFKo7ZTp
USfQXgG8Dt4Og8RRegnSqOP7JyRCLo5O7Frh41Lnm4QhGOe6NShcDhWtFwLlakJe
yEyGACSkgEKABUVN1T1Z4PjX4R5B02/tjyxem2gWF62aWDUhyh6Q4MuxaeD363dd
TKxoGjtLvMvsH7sz2O8fAFsFysqXxfVFccRPbDAaySmkry7s9PMkw7r0/Z2P7hdX
mjEOA8hHhuM2BTV7uT1VelMPiycZ7a5rElz+3TLBhAQESwsK96W2GdQT/h3ggCUV
fIAZplmnjJkTZ9qrZREy/rJAcC/wgEJagQePv7jwFUyifl2eCrpsTEAJfCnq9bFs
F92H58S1SjRHR39dKct7gHQvNmnBIE3RxEsszTWO8FikS2sYksRUUwATx9MD239c
MZ1Puuaic/dbi3G5M+N/sSrItxtB7KDOf9YcsQdC3v84IFw+JYDsvfWRT4s7gflk
ZZqpHh5k3BebE1ldlwlOA9yA6JTPTBR0/6Hjyh0uzSiDlVxro2Bc3kJMlB5yKw2j
Nf8f+XfJEB/OJUfy8zAONXaVLFPSCa3Oa4N4kNGvQmjaab8aiKjRB1PYnLYAkcpH
2ryFib6XOctRcF4XhDckcMN13evKeoHPnsJxIcco3wQqp0b83I1PjRtGSWKZC+Le
ltjdQ/OtqX51D7s94YoWWesBAdGv2/u5GmecLhv2/H/uSO69iM74uvLc0ns36ErQ
7Xzye+6B43SOp8buxGkEE2HFSkBeG+wDTv6XdKaUxbA/0961yqmstESnsdnXKk97
SXCIAXpDVlvkBlvTKVXGI7OHWvw4Cj+N9qW+sAAd9LLzVlnjHc5gqUmaErRBdel1
PIsRcOnww1llZsJZDGQCXvT3CQK1Y8KmcWLfH/HvD58brJsC8JSCchOgV6WG4ooN
1Ha9e+krgeIUzVl9TzyRmGRRgH3RY3e15iouqtIw0fEHlZnLJ5HieP7W9VDrs7MJ
MAqut+dKI7eBgjUYIArMM3UjF+3xj4zL9trFTbYfahrKvRTR8fycteJpCl4WCSOS
aaGBd4tdNGOTEFHzvTulHZTbXc+YgDRlA9hjur3F2hJ9zWbiFiB7piwkcJ0sBkSK
2v1hc+8elPsP4QiI0StW9tlHvIQyUdue15OooZOlRK0IpEAmC0ByYfzrQxgGp7jq
1cL4hNicukwxxApt3oCTgrYc2MYzpozblrGje1PXlOv5q9X0EhYGDLupobLP3/mv
e/M+HcP2GtWrYE2F0o35zxqzo58m0tb/IrkbKagiA4KN1uQ/ovaq9Iy8up/WuuRr
vnNy0bP6sxh0C8mhkH4annMcPfKeqJYkk856A9PHFWfpHADYd08OMEv2giZJAJyJ
x669uFEZIpHVeA3xm2Nr9pk7mZ00BgVZZZ/KDB7M1djWQRhQbfo7ns3MO52ddka0
afSW9jYTCfoG6x0ot2vYF4Pyyt2z4pBuubwNaWc7sYeWjngt4T6SnRD6z1UBiTGU
OsAQQNNEZK40AVRF3JZaMCHaCbE/honjEmyMeLf+mhuUHwRhVYcqbJVKQ519eNpU
IqSYs1JTXPKegK57DRYbKu/RrRxIey5PP1oE+DK9HlllDPj+cCZ4Nz1xWuqegc6T
SUuxebe0HBt/naoZ/XcLj6+0I8XdtP5jgiIDBCC2gCt3cLrPxf8m8sYXi9bawbPv
2+GDQ1Lz8eYm/Nat0ErTg5Ltea49tC60J+4zeImiW5jZLMNmCe40MgfGUX+525Co
+my/705oD1GAU3N+1tOOnodKrXT+p5elmmNIzDIS7P9kBhn3h1bRt8D3yOllOIV3
1GBQCeYd/fqkegX2a60CvbcoBm1aJZoyci/AqNRhG3146iLJbBDVZ6wmWDF3KokQ
5GMUTnL++gKZ+Ap86XvN8yLo8SUhPrPuTYq5UUuCUwVSlM8bRkXWajtN46+t8eks
NsgNU0a6amHQ23rM5uYuMxJfIEKlGLXuAqU6+eJ9BjsWxb/dMKjl7QHocjZeZCUw
RR1QfaeL57KbLbPkmzhX+moJ85vUlZQHBkwas73kTpOt3lJoJCbkMK5136CbbgAT
L6oTOynek/45jDzuMDT2o5GSdc94/oL8wbRViryebIWtB+digUTUgx+ca7Mmqsuf
1GUY76AYQ984w8DEvgXMNuGrTvWiqRLg4cROrdl2Klb990x6CGZqu4g5MHycDl95
/UJ2XdUkthgqYeygBwBb/Q71zgLoqn1sWmBWkJsrmDBLb3T8REQwQTI1kOhjHwIh
/Gsft5zcxJaeLshlrV9NWB0xoMlOSnvfKXd4PPsqo2KeZYXIm3vXkAydMTM5MB5n
UfbY0QLDgrbWTuky2xZCgVaK89mdlOqmxTXy9wxuIzhGc0mA/l3yCVRNdJTDQazJ
aYA4geCUboH5m6CvkESxRqqwa9wXlFCFWq0ZLRtYWn3I1sCD56bZhoZqI3ayXnp9
XetTg71AUK/bDfISffqRN7r5nVRoOi2y/d8jyTHAeycd0BiOlj7fuy9g56RbTjbu
CSXJrK5Oj4Xrz/B9fp2Nc851g7crNK6Kj0b5cLTUoo1dsOAF5iOezgR+p8jRFO/A
66F5spf7sh/UczrxUXqKCc9vLIhOsut7HEUeed33kdK71hqBWXi1L9Di4/hmkA5h
azDKRQ+40Z5ddy0OtYsgCra38LbJQIPdA8XcYZ1JWMYcMuL/pM7dRqL0UBiWRNjm
Dem3f3d+ceEVmPHCfutDhtj5JdMZfVOcjCsnHJAZtRQImkNeCillpHD2JOZBrQbV
tzZCzsZbsvHYbi3zYg1ZvLOHLtjUdiKhsmlzPxKixCsTNrxeF8SETTH0cTpyhmV2
Qwg5x+24GIVcQiKiAlvdkoyqI0H9I1+pDIgK2Wzlyin67YvKf+tMQf96PaUUdMrd
KgJKNO9X+gbc/B9eHkIjKTuQG2l/OjTOYyHWUUYkWSy7KG3Iu5pi4S4D8PFIndiC
sDtIO79c91LfyeFMmPB83t1Q09IFWdUGB5QDfM/bLKhjaSoZBR1qD0XjZmOydyQ1
xb+E+VDab0JYhfeXzwIj+HxuHzdY3syP/vuMq2MJeanHmw0qfPN3URDBDljZ++Kh
j1tOpd0zMXkKgMK+iEEAqGMi/YyFCJ3xGRU0CVFDWaRPal5DdqwHa9KiR1vJ94aI
1n5dC0fwNe3WHWcmMeyyRnq/LTRn1VW78p9ygqIr1VXoIX17E9qMvglJ9AonR+lj
wRilEUaW7/wOM3xAurZ8Pkjy5uqJXx9RtTLuEAFIBXBgdXmWmv0rgU83yto33lhO
KAy0gTamWaEsFAQBS3KUBGNCztim4nNETlGF7eV2pr5ttoSk1OStllRwiMrwVWBI
SS4Ej+MIhtV9hcQUUBzP9ugoBdj+k3kTNzWvTEqMQnXScJ6EVbDKyTAtfa9H7/LG
+CD4lJ//b1ALl+rU1/4iCwDHsdJRKDKXvxEe7B3GIJ0gOf9HOgFklpM+1S9NDgjt
5SrmtG5uNtYvenmh0l04pjFWwUeVHm5NvTpoyvullMgTuC1YCjubLOWA026irU0T
8YFxV5JqplHoKNCMSj4qQMLsjrsql3GuFy2rlpYrFZjSK+pJJKqaSfJXWWsjVRH4
bPcMxPxtiblytFmTGcnbER1T4LZ3B1CQuKAPUqVudHuIs+RbnADd+YE9iDPXvZY4
iktXMdfwXkRN5hy5Cw8FSXALHbkvuCBcKKzMWA/8FSqd3UdYc8S4Ow/vsFJVyx/r
mi/4I3na6stpFnCyhxLob70Y95+xf59gxfcboMRz3Ur47GxDOM85yFEvUsWpIAcN
RRNWOJ3qxc+Q8XRLY5D5xBqNzlp1WZN+8TsXlJebFE+Hv5Oi2XHLmIii9ODJL3E5
4L8Syd499vE5ISfXouEstejn6yEyUesI8t/yjXWmcXz27+UK7JvwF98Emp1z1S+M
8ezR+gra5ON6N8DMlAa//kxYJD7kJx9U9rppYUviNMwJTeBRnKPkTsoL4BtTFBWQ
h3E14vRKAo0p8PhsNB4k5vQfalLHzV4AGY+Y3eu4monKDvhQCaXKLQ7MypjXE/S1
slpfefvdeUm7P3FkeivLWoeEUgR3RAf3NJxjcM9bOE05c6UrcyvUKTDd//au1lHS
mhGzg/9ZXsjgB8O2hGnpOy8EOwIOBx9XXnw1eIT9J1y7h3rawOVXasjttqJPF4cM
ohtV6onVIXAfvQEB8+q5ViuKorM9mvMZX6+cvaBQTMLlcw3OySfELOkpd708w+cx
oumjZ3Q1HFa+7TA6MNICg2M3j5GCCXjvnfmj6UbcPgroGcTMnSRTGPW36zFJ078B
ZXoQS1f2AF8S5UuFc1M0U+Os7JXMSaiEcFQWzSW42nzlnphUA7jhQoCP1Ha604Lq
53vSNhqKLebY3Bg118x8YQ6UApAi0uIc9b4myuEUJQElIe9Nq0rmN/sgAHgnNBBx
lmtzuTlsBdyvf1Gls9tXb+JOpZ7H5sB23knOpGxsHoB8njW51k2OXcEoTTCi9nGy
5Z/g9J0hIsX1r1o3yji+uFYRF6asVgyOO/p+sWLicei3ERO4XyKkscFFd9uISLuG
W2KNWyH5NemHuvFcFzYGTi7H9xYYQ6G4aqRwl/IzBNir0DEmkTBAC2yENkky+/Lb
bbPVkl7TEpHg6sr/+7AR/+uJ2Xz1miin50ShNNtKWoUjmMLj49tAIxynwIf34GBL
9IAF6x3M7ZlzCRiNMEZozgOUI7f0LayqezOHmmJryQGRoGwojnVjQO+nezH/4A4J
Fsggc6Nz6IOXwBsBWB3Jaz23dCsn5wiZ6XitPMefn4FXi0CbnGTkJOtkNYJzs9Vk
jFiasxwvdrmvCJE7Gw05w7Aw/a6bPzgzmiFCh0TMj7W8k/+Wq6Fg75Em+xIRAfWc
KmHsXb1+oNp30xqCWuEWouoQiXRMvlErPJLCZbzUHdbvvkXQmKujc24ZkVbEU8S/
khsguyYPajMaPLDGi7SODsBnfUlURy1PojMuMGu5nYPCEOjXDl2I4NM2SEpHXxdt
oEj26rWsYQJTomV+mBck+x0MTTO9JATjJhnwYofTrGGWvvVzuYX8C4MyaShjiu6i
w9DuRbn9kyzw5LyYU+1wiPazua2vvD45xsq6rHBMoApZZP/VygkJujCzf/uOjihJ
Ko7Or1aDiVai11tU7o4ePBXi6L3cPgwTA98j4kl0jMI01Ek5DZ3WvufNG1Y6FxbS
w+Wv0fRmkS1yKX+U81xb4Vi1mmAQEiBAo03c6jczmujYzN63MD+EQ6x1CJMjYo6T
HEdUbwVidQblBEz4NN3CgjwZkRnQGcQOWDCP7ubzgUuGX3iaK0O1NrXyfnuC/4b8
vWpws7JlBo6xBZ4qOtOhZZTt7bw0K0yVwXf0BdqAROtdCzhJC2AuSZbHcmsiMxCO
22Y2Dky7CxUntIL/LmlqfBo34WacHPp6bK9sAhPbIClnrnZ3Eop7Qe54775sfTpy
3VlB1VzflLGebSpzpcZkqB7QVl1tBce/+CjUcReKrhUMmk0M7B+V/GquTCuYSAVd
Iqz6TIlIJOtF1q3GKgLB0l/PUsGED6vJDfmbYg5kj5EjIVnS/s716uDvmTiX34y+
pzv/DbQq40w35BJAhO/dgi5MYi8rYP9kUqC/O8hVzLFz2mB/lCdO1XDOmciYZn4+
iL03pjbYzTUv4G5Zn81HAIKz3IkUIKbXjwWc3CET/2iOX+ol0cSeyT8n43fXa9qT
OyagSavOn1fC1h/dN62zrD3INPrODdA22DGCFWNr2PZe9wbc9CiJ8wTJKglAtIRJ
h9C5fYV0ntZ1y2ioNfi3vspoOvGargrTUW9oZeIboX/BJKSFEQyqEAovGTWPy/MP
8x30DlqBP8oy5WaCg2tgkykujXy5bBVlCi3Oa9UiYKJQDXX1B5gA9RXWTW201Vwb
UG6k7/bUsiXCzHS4VSf+xcFzyQ8Gy/hOggAkT3qR3YIbRY5SKQ4UBLcg9+Ji/4kz
eL400GhxnSywnyKJfRD2IEvUuxuOIvz7DaXv8g+9k72obIz+DbdktKdUgro1F6ji
IRsTn8kglnawXgSQsFjMgreUjDphGp0LZ5GLnO2APceuRv7fjPhHIKFfU9D5SgGZ
cW2hI4y2YJCGHPRZGi18E8gKHoGA3qgxL5461fSxLBf7Nw/UT07BgEEXsj9mLqms
xkxLq04L0aPdASp4zu1HCQyWhYLE/Uwv1v1DWECtF2GldsyYEywpgMFI5SpqhSJ4
Ut4S7i5nHc5NnzsUrs1EuzDxMot/plT4Eabz5zVrVy8wQTq3H6da7gHBHL4+oLzL
oxCLvXSKj9tajvuylhMyQONU2C69cHqEG5kzRJTk+FnKlnoQlUvldmEkP9iWr1LV
gHMb5L3AAOsIF17jl+WUizyn8v6yjMndnmcoSHVa/zJC6Y9zkKw2jMjM/Wyel1gP
Gj0MzX9NWo8Rdy4nmbsnI/Q5J7YpM/7XAOSY8g8gL+lg3xP7VjecgFs4+IObBcOU
8263xHeVEfg9Mk2udaioHG15EfLRrCti2Ea50/oVSyqnMhH5Djw92FjXcRF6Gr8h
H2Wi05E1gIXwpcAOWfBTXef2oosccHPttBDlY/r5E2MT3baZ1152PobFt1cO2aGg
si2qG455Rm+zaigRYEcLsAlXgyCy4AIMUGa6jj9pPj+47HvFE+/XZ1ZU6JrbgiiG
Ql8PPva2FyeuhE4v9TjRN935XaZo+dEtKb21R5BjOB8OoDFHr05j3lsJ4xg6G9L8
AVONAJXLAhZ0dfBEew8eZFizD/IMNIGytvuh62QkdqHUMKJwUq2qkC8RIx1T2PmN
53GWn8ndhrs4KIGVlpohMAUOjx9Jbn/UAIFX48ka2Qxw/jU1cQ61edq+J8eIIiJx
T9yfu1kDjXlasrfYzhvS40orb8OzMD8iOZQuqg+UmBGZUhNT/TT81R+9gdL/vUgh
SdwHqwLtEbjxrUNVpf9Elp8ZG+IIFQm8R17U476/P04g5eb1GjxuU8zGJB5RHLR1
5/+C/9Tm1LMM4lZDNKx9rf+ncXUqj5oL/vvNV0Y+Re1mSRUYu+J67Yo6eckYv1ZU
SYZLoUESaNeL2L5LCJWQI/OJ/Qo7C6HwN5nZWyiVEAv5V8QIouUtPGnZtpr/5HKl
f7TPqFlwGIpwBUFWRAg20S+/rIXeqiDUSyP6NQH91xejqSHmmSTRqgLKoQ/sNulU
ys0POWQjmgJlyPftLtWwT591i3OykXllf25Umo0zak5cw/qgr6vPQgWsPbIQ266Y
XdSTnxeRf7uUSg+/MSt2egyu5kfB21EsOfwGfCyW3CjMai35XPZ2uSLXZTlL3/yK
q1IgZ/glaBn7engA2Px9HbVPOEHJSoFgTgJ/REyW5/eAJNMVX7nB40WV7gpTBKam
UUrfpyoWMM5xOAKxQAY/zgR3ujpPbhtUdT3BGkkP+zt7JPPjGc3bAWT5chWG3bnZ
/iHhSuZdBG+qx2pHCHVE8yNmltqnTxbDIjnC+R1hlWX2493q0xL1Aqehf+dlZ5bd
BCSnrAZQz3Y/rcHsD1cBTAZz30JZj8mfyb5CC70xrJ4GRSjGcQiQ0mVwlJmE07/8
88nfhW8gBz5m5gzwFO8o4xqEfL53q7u3aYH/KuhthTF8ZEIm5grFpxSz8oadCRDH
/RA+Zruab1eKyk9vGSzNmw778NvWtS8Ie5QHJ584E/6Nbnh93DzQcRN8MsHbcgKQ
050d12/RInP6yp0dgfxOJ9oCYeSHdq+l+kxWNiP+FIxT43HctNUamXrKlNhJB0gC
4+G8HR0P19d0TisxU1rD+WxmL1/jL0LUCu/Z5JwCD8X+sgAzNubcb8NUQn8UfDTK
tn9JZrkABNtfISMmobEsm+nKO4xVw/5DPJ513F9JhivpxfaRUnV8enNXQx3rLdhn
mLuJAvrla/fIgTOubHS9BZoTAMbhJKO2GFXAsfv6cL0Aic/bMhD6TluXBCYF8s+z
6TbYDqPnnXdXdBH+njUwhtyFxNnbZbfKSHbn4cKh87d6uqq2+in7s0+cXdNiY/Dy
Tc3bIc/CmIjhN7IgXvcb0xDTASEO7EcJwabXJO9NC1Y01JmO1k2YFbL7AP0vLK2P
Zoxbo4umZwUZte8IfLJ1kfWp6hOjUfvku17TjOrojL52glcrs6OhNniBrCZPgCR2
JTisKCTCyBefEHwi2XOK+blo189S0uTgOygNYDxovhBcHpx2Ef22uyd8W5Pho2qD
1D82HldQilcExWjjgrDB3gaoOLihBTEZ5yCcIOHkbdSDYsLCIzqMykqWRT1pl3m8
7Jq82FKdJRTGeql/f8g0r036bdnA6LDTxmgl+ePfMn9rvnNEANQy2SBJx2RyLNUF
ZuoJQwM//xEeKD2Fey3Fsvtmd9GZ8IDXysbScMklLM4nRXrdX8hLKBs2N/jaxywB
X8kMIajxFZKDBVgGtW6M2jPmeUvGhhgiyu7TCzhwVuYUGC1B2xfKoOnLM/0HH0LY
0v9Emv17y9bhXggyiDyEXx9c3aLMx48LXUnGRXaHH8kld2r9HTWi+0XHxUxwiBYP
7NFUbbFKkPDJpcyJpiLElRwlmhb1lidVKERiWpGdE/MMQnQRnfGOySUtHBvEZErX
1pNr/H4TBfs6dClq04PaplJZGES4Oc1qPByGEis7wKDEN5GpLuYSXlCWG+nBPjjm
fnwe3ygUpEO5r1NJRGhpyoF9FKhQ+nKWUrhSeAwoYQAvWaBkVBnJjoqDe4Dgtwz+
+5N6aV4sXaquW6lPZ2SgBVVdUTtlots9MY9t4wsDJWpVWRoIH+LfEEpouTcRG0mw
hfAEKlI3JuZ/b/e5y7I9cVDyrujZTJ3iYm17tkSxyJYJ+LdgwxjrdQfDXxRXnabK
7mcYuwRoibUi0+V0+8/Hl+N2/V9+x0+MQm+sySayvQemjJhIccrdM64RVVVhrBoN
9MeMT3pRrZO7uLcJfeUtKhL1NLZKhR9f9dB9ClSmgzbuJXSU61OjNcGZDSwNjDSI
sHZa360tQQhWe/hg/O3OY6kmpZ/pTnVts3c1ajm84U48NaITskUJrtBkQnT7fpzc
/HQCKTGyS3TyMmkbTevPwTBkFJ0Eb8+Sdchpk+sUbEAtVixK+GWojbp9St6HpXC6
JIxg3QyoMtdu/y2DXgdWB/Y6ZyiR/Mbd4Akc8NlMT5CfwTjOoCOdL//Oe2VpCoAz
bYtQjNSfz0M+5H8enjxbQ9wtWLfPZrlEJJ8GyDo4AKA8ObhKACK1+73Ton98hO5X
5U2EconyMYB5aTkHPpYb7ChQGJRpjFdJk9Hg70AhRgYlmsIU5kKm5A9rgYJ8oHXj
tW6wPoBKvOePBIIY2RXJjI35TDeGjsso2wJHzIVlwjOFP4ixRVHiBFKkTKtvWvzY
4i3AtiTqIeWbjT3LfKIQ/aeQtvx1ndDX3fU0HQJAc3JApxxXCqJG2EHnrzN2+bm5
eJmLjRkoDih/xUhy9rGHapIFnAJdL8GVNU9kC05g+GPfLZqxrzrHglxfKPpOzst9
8mNKBUl9g9C92jyaV+m0B72u/1Z5zK7wqrjj2quQ5fJaXWLfHAju4rxXYkXz67je
tIrEMUH7PSbEYB9JajgdfqevgAocF8xazz5B6sdpOHs3v9Nje+KBeIvisCsGK+3N
n9X0qP2ddfU6RbP+fM5U+8GNqI2yOa8dbZ2eg3pRn9J9MumdOe3AmFArMR/52Ytw
D4zPjSFtsew9sXhLey690kSbZJsRdHDpKypC381X74GCv76g9UHMKwF/NzN9wNvM
2y6Q7zkaLkD/4JSdAIplW6vCf8jpzOD/+9AGrsrkPhHeGWPPAMZuSywsZpCv/JX9
aZFFk0NgzhzVnRwFEYlX3k6PGCwGC0BduY8JOCny1hPdpgGyGRGGefB21U0x2oxM
REYPSg31IifjGQGFmdUAXSbzkOfW1I54+gX10gAqR+VSbEfjLN+fFiacaNPjNJDd
tKnOKEcvge7qxws962RaXumLJbhIZWJvu/hZpIQMf5L2ZlQJq5c/VFsRqX2VC3bB
iFCeHlzwjmw/TnJOfCOTVxy9hL8M/PtpAzb55cR8wHXLqFfyAy6ScEUBTdIlrjCN
xA08hf12ENPcOngKCKf+iEsX1LEXKlT4KLYFajHJ0S5d5u9Redh8nSxm3BFgMMNV
ORQFS34dCswl5FWE0cBi44jflcFiqrRbXf3U4bpEFsWHY7z613oToTsaDsYz1Kb3
H3BJ9Sl8yZUoxazFPHxlpy+YPhg88deHsbuaEE+XA50Dn+PJwOK5thZHYA2TaOpe
Fd5GkdaEP30vAZUn38iWBBJVMuxiCXWJ2xUhr0Q7IYnabqXxmCTJFsTEZPlf80oI
wbBRiMcFEGwPl7oTrpPkc68Cx44FSonB2YHKT/A2C+5QV/qRPrrf1gX/nSnqo7/p
wzaPK2YVMGo6N8m/GKv2egNo3XdMFHRCVjE3/YLR1T0Tq9KrGWhQ702NbKQuNAYD
g0qgxGw2uCDHTslB4NGQ05UtB3+O28KuMmllHZB9MpLlbqVx25pGn4Vf6pzA1jQp
lg/sDlr4w/bgd50ISqlgzWMKKX+xqj2W4PevXyixHNGnLeFWrE8OSOFAg6CU/YmA
Bs/iYXagsX47mcUzqGxKw0nFmnKdYVLseYvHKTLsppoMdsWCRGSWYmOTRgv2jO5d
9meJkkxCcbbTAGpmc4Z3h1cw0hB+4RxeApR5jPmgNqb5acx2pV8ptNXzBdf2+NIn
Vq6wr6PBwKdNGHDlfSijRMumYV0O9wC+TIgV1QvVhWxWJt+NR0uyaisJXnZDy2Jc
HZpq5X9kwD00Z3AOoHRsd1P4KW7TrX3LmtjbNYzKqaW74KpZ7RBLGZcvcHSntw/q
5jSqM1oWCJyprM60vnMpHlhUt7jC5H86LHrld6Z4+qe4scWyNJQ+YF/SqSfcUwX6
v7sB0eCA+PuqJsY4yjVoNHmb1QBJFyGYe6TzDkrH11lc9QoItfNAxeAbuANDz2lo
3NUfW2pH7p4Q7etuAPwP0AdYKeBL+gmuEUZiZii3P9OUY1dA5oURiCbswm5oyrhR
SGgFAdsFfVYTUvA2u/r9aV5zuasOH33fHGT3vJSfGUur1lUdmvSuCWF7HDLkh6Rg
56s7kxqeKbnGVl2yd1K567kBZoDj1l8yJ07vzal9svZ8rCooFiLx8owUp2n4jHM1
xRBMstuq0sVlbcvnLU25wjHOGmgStlETz0bqoqisDbEFSGnHAgpLcQFqcP5LDjDu
vryOsAJAbuV/roMdKT0BGHb3ZBdHCkL9PYKIz8aYXdMs2BcQS9JE3SO4/DNzli70
JcbMAnAbtPBSzPAzjx00bMh8C+t+gCsvG1nQvbxKlwI6cYLXiBmYLWFjaJmNLRYl
YdQ8kXmaiCAOig7ENHtWeIovW4EP/JdCSeJOftaEwgahuRMFu26PmJRkaOYJlp39
zuJv/VugtQP4DmXaRJjzEUlC+yWM802TAk76kKLS5qUOB21ZFMsp+oao/Yz0WoMP
8gQ4b6gEg5EohkhvchnEmlsnTkpDPFBBQ/Ha0zB5BHogbR2x45+LE/jl75gH+CWR
bdR4UWtdUwtwE9+7ip9umgYTEz/Q48RiKHW7i2ct4GBjpFO+DuNgI080wlgEKc9M
v7fZtn8wU2kvh1dWjajMk340xfb8W4wgzGctxLj24hsXdKJaWlEX6yNDycUcKoVX
6GNGsLxLOaiEnxDx5IMXgmQ26JKThhgo6J6aupUc7+NPygI+WmdYOLfKGJorAIy6
zOnAA/NRKxcWs8rFikneMsac88m4LkRttByhFPUTfGfsZaWwQl9JyB9wMJB8WwXS
RdijK2LlTt4pfdqgxSXQnANgnp0ae76QZinfgwmWo7gz4tB/3P55F1F+l5vdQB9K
mWHDCy+lZj3R9s3mAGTAQZ2N1tdRrVX03nvzZtzpyJJNK1fOtVtiwp3zA4SN7QyM
raQJKco4r0ztLF/oQjsTYITqBoMGs+I1sZeycvDXFIrCjiTt9EnzdVdsGcVsn1on
8aTAJESPTjxvG4/B0cBnHv733kD3trSbYlp1KNp4hzWKujud2czNTcBXjzf2MUbw
0Adeu1hxnVShdDNOrh5DPNcpl/DMp919O2liYDvEdDyHpBZIVoGh3Y+Qr1fr9Ood
RXvIoHFk5K0TkaN44TFEpXjM8Tx6H6xtTw29KZnuQT1H25pU6dkh98Yt1W9x5BIZ
UCesXQJo7aTUiX6MANNH2tJTwbLuM7V/51boX+BzKjMLdO9KR8iR5XzX0TnHEhmu
hA/c37VdUxc5fQ4JOFdUHXKRBr3AZaTmaRQ6uR22wW8Ucy4xFJfz5rZVze9RZOxC
Tn+MsuAKR/MTcY2wxDeAoV7G73vy1PkTJgV0gTyQbQO89+0dmEFmFZEm+LVgq9zy
deDuI63Jhu2jg0tiPTixB208CotD7TDFYwSJmFJ/2CBfhveB14Sawin+pC928+mL
QvWfR31pdi5KMP7YeTBM4gVkwQ5dA8MK1FjFUeolAGmjT8yEnAPRp6uIPQU+4weH
jNW2QzjN7y6SlbHrqMm0uvA3KYzMkqngsF8YygzEQZAOtJtFC01xCNfgQ5fNY8I0
QKvYu2wnwxvYCJbIDQ+vPGSTEz/WJUwnUekrsaoW8pFG3Ov6lY+Bs/AFpegJiT8v
7wxf77nq2KCrR2Kc20EKtcUz6snbFwdGW4S1vtUiZ7C7/4KH5YWlh8tdvdmKpY2c
4iBdTlGdd8vFSILL9qF/VV51UR/2d/ULkTEMWmujzgs9ieazEZL8LWKgZrcIp2V2
p+RCUXQ1eXAA1K+moAQWJKLOrqfZqEmasVJXkNWg8MHY+dPHpJu2fYCXJVfLkB8H
euWGjCzBr/lV5eBXVvGNXKNdkh3aLMYANlTZWVIarIQ4DE58m4YbMVU8wRTfP9CB
9/23aS99rNea/7Zj/2/YoXonUml85uTgYYiwFCpCJs2LtgTW71BYaiEeWyb63u0I
jiv5Tzm14COgYIZcYZmPEsW9FdO+7t8Qbv1DGcW7A4rA2yj23/wciby8pG7WqnsN
LTu3ROXhTY+0tP56zGQmkimzOUFUiLSvLGC+JHbIREdY1qS/HvbdhT2ha2MpqeLo
KqrT0Mr5dekV87xu7xF6zpq1IVVknDKLxBcJNSKqhw1MlF58DFKXzmS0m0tIFRQg
JyMGzNbhrVVf0iZ2sronkQV5oCGiyrDcHw8ZpDzQ2abuoqA41aTXR3KCp+pbUEUa
UszaFqO6Nv1VBJA8yX6z0yHGeaB2loUXBsqt/1aicgpJPhrmEZhKwU1HNo+rqYTE
kxYLgEzFYg8ktcV6gnRA/aSKjnQYjq+CwJcosenFTJQdNWi7apFbSHLP5Kz8rUOE
m/LDP85U3hh4F7QxtDnvIbK8ApLPq1xi8vdN9rBC3oN52k0fsNCESF3wlrAssZ97
TABSXAu5u9YIOKI4GdeEc6Fy4mr4OfjRFYzA2dLEJZmJ7KQN8DJzwDqCvkMzN55w
vQQ6dD1L/8EfneBJDI2e3i4+3cJifGrhlh9Do4kFwsN5+9MxGlecG6X+fXvCb2VB
2EjSwYDORujVzJA3hzDn0H+o8HaaOWTWQkGVc7XFR6wnI3DA/kNUxaK2chQ/YbD8
+i6pOk9tPvgXCUfHFIgKVa9vb9Tl2TA4Wx7jkY54niaq8Qss1kdZKLDaUUMbuDpg
fGgHw1DhLo1Of/Ayxuchzi4dWq87lQGpIHGwrvwdh6DTpbbFDrhq5ci97dr9dXPH
GLShpnBiH3ZsSd4JVVolamA4FC649FIhlz/Hso6px8tSw+r6eQOXRQbEeX4NsXkS
o1GwuP8GDa+QVpIJUN7EoGhtYTzZ5A80rTmQa3f3l1IvLhiw4ZuYX0V4xOgPk/g5
KUyPCryFW7Z0Ul0S11cppnIYc3KsH8So0weGdKR8Oi+uA0N68nTwW8uRqLhofY9x
AjbxqK9RQYQw8SG9M6kvahsvwbX66fb8PPoBHMDmMK6bcjCfxLx9fljs0ZyHD5ST
aRRoBN/8zT9B7EOpR+aSRFCMlVgyMoDnw14a1xdKoa5GZoaPxXG9IZA5FuvxZmCT
Etj6Jg3fp7Hd1Z/R8QPLCb1wdvNn3eV68v5pejLQlqfuyCa6nsTQIeJrNuKtl9rZ
hBsrfM7/rSrUOBaB7XA2ui6+c3dMcbgGJRLRhUyzSYPbJ7IsIh8O1V/L+K4YTLhP
SLYhf04x2bEF1gwYcz0qAfPyKjfDSbGLxsXc5Nzo7EjPKit/Y6ySUsvcd3Ojk8rb
hFPv/Juf8ZckeZsC8CbMSKs+PfUUHQwGndG52Ju9CqFbjf7OD7KW7Z/TOE+sx57h
pky0fwCIiT9MDSdTlIeskMmICktUbqP3XFmJiil40h8/syN7Iwoa+BD1bBZs4nnv
ERNcLDVUpiLdfXM0EEeW9/dtNmuElZTuCCyEg+ufl2LtCZ5dcy+28zcnZ5BFrG93
sjb1Wrrs7bC2x4qi9dc4b2+2rb7FsmzhZXW7U6idC665D5bNm1y4d+g3bB6vze7t
K31hy5D/O3TIRRXYHxhSNs+rRJ3mPwTv+bp32CVL5Skm3pAdCcH1q2r1WVoZ0G7H
J1LhDhCE2E4P0CmveVF/J4ztG+pCJTNcbIkDjCnsgN9Bt2ZUJX1l8k0NGkpsH4Cc
fXZQ/WUx3UwVsE6ZdKcQSaYbH4oRpvXZxI7JjsDGo94bmS4dMUTppzDIfHWpoXMU
cBjRY2GTh8EjuUWXh9uQgZyI7p7Wb/oo9iM7uTRtnZYo+cxg2VjsOtUl9b4RnHQs
3zFL9chZjBHjv4vDQyxB/Te4nZjmZu5wPc/zKJU5jVenzhMejNAgkcN/i6O8v2Rf
TyqfKnwg9He9PaOUaMnJiz0722x+E0NGjBymZj1yYqtxbbpx3iGUz5LOCFHvqKZX
JZEMNY1OoxMzPRO0NL+lI67Lt2s4iHUdxVUAFKLPIckuQ1/+4R+Lg4naJjcUZLIk
Zzlkf4osbJTG23s3Ap9embgKvIRvT3tDGQsr7k7MvuJynDw2IwQ3ccW3DUG8ThX0
LwFsSELSSQVz9Hyek1ZSNA8y8gHh7ZT+nBuzKa7Jy2+oo7oTtUc9P9usSG28BWnJ
PwTmNwD6uPYTNYcSEsthhwrWl7XjdfCME5UafJaiZDtXMhJswoSfVaSEPx8Asbt0
1M9UAdD9frc4AZc9YGI1IYeU5ycTQLtAgHqfzz4X859u2i2Rc4DeTXvIMAhzEcoV
G7bFhtvABU0y/Yjmk1F8Er66bp6eTXqNTA7QVASNeKoRB+mDAsh8U5e8JHheo6eC
NDT289nyyJLEBqooR4uZHFTi7o88GDhG4kHzC84OapgcPBJI5p7qkVzQYYYK+m0z
1srA9wzhFmXCbcQassgvt4F4aRdtbDlnzfhAX+7CVmtj4vWFeAJcvhpgm6DLBcxF
pnuKHVuUgVIXhQwnbomDzdpF8pk7jA/2V7jGM3ASKIgcuOEKgkgpGJ+1a3PfW1QR
3/fVyfBOx7mmdvzRagc6yoPAPAiF+jgICsgyXlGR1GQ2bbrgJ7/NCE/b2zkBidO6
yDkEqxxLqBW3L+uWUqFsGJxABm+v6oj97Zm+JpmkhFQFGZmkvSpedrgsuVxXuzwo
qr5RqK/HKTH5czR0/ASLN8/Efsdf5B1zHJbF2wl3iWvlJdPtp4hIBTC6FXGcWb8b
kuSxzFwVbkAOijIC9gpSxPgO6xYTDU6mIorhndcgTMTkhk3rhLTMswge9/17O03v
6fFTVSNrym02y+08C7wp9rTxXff6IXADRGWWpWHw7mZYTqPGbuhI0n1wuJKWAWq9
gpf334gvWWlddcgaGOr+QJtt9V7/4M0N2+apeAJ1LMfLCnFQ+SXKD/dpv3XI2RjM
Yl5YvCw1tqdzNIFIrV+9jFQ1yn3mf4a6itDvfe5TlIkoI8/157Ctr0p7OdoJywn+
TygN1GQ0c6Qmn1q76m5fyUfJw9mBKtDH5e/oHhKyi36up2ENciKKTK28mFsOX92A
8Ag4gsogHCM2rf6vdDDDw/FLWO8LP/Xv8Eo48rf2TkZ68NeMdjK99yZq07iJrPV9
Cwu+9TtFrJdY+6UYwGksrwb1u1WZQxoR+7A4Fo9h4CXQBDZJtxIqAcE1qgp2XMun
LZVumNxaygshpBRBTWK6/WpSW1uKowGqsyJnN0VMU/2vEAAh+qB4lJ/jM3c7sKOQ
OnY8J686QU4iUk8ALIkvbpdlginhJADr51f6lxKOZj2CngfXWJE8ivyRy+ZvzGC5
2owbk8tEUVkF8N1KWLEf+EiyQ0/q+O07QqgWWagjXUYwVXfpnkZ6FJI9YIgoc0+P
Ja+HqLu2TKQfAq00Riy39sGA6iUMe9Zj0Y60t/Hol9TEonxB5icgbplrrEo9Cmq+
pZ+sxOlbx+ye6QllKnG04i05zRlMXfxIIYB19oItVR0Ns1QVkeLr8dF5cWvW2LPb
DcwWtuDwPZRAN3XypFAmgGhRFh0uAZ8yCJ2TJfdB9zKv6z7GocrCGQF8iSkzJJAl
jS0HgB24RVG1LY+qB3eL+sd3Z1+JeVeHerEsb8MkGOebXlSlJv0l0ALuzXLD051f
d6kFBJSac+UtZrFr9C4oHO8RY1lSQYyGx6+zjcoHrBG0Zke5s+G3ZnIxAtQI5CKd
pp4ntEF5q9fRSGUU4B9X9+FGQda2tWN4o7BT3a9qRd13sof8tAz89JrZh1I2HSU4
x0FwASYfdfP5tw412n3etL6uB/L3xZVksy79+GMfMFDF/pj3PJ67hVsTKvkCITkt
UZdyajqoud8VY2bB1MwDKOYoxWfABuYJqnKdRD1bv9WOUoMJv2Ie+di0nAzhWmvq
kgkgBJ4CDYRATSFqoiLEdPwzmtGFJPWOpeA+s6BOLC89PjRB/Xm97SVsbtd0VGhJ
U2Kdzl7Hoa6PJg3hotbDijO5pa3ktz0xNeSIFmVklLKxHHxrZEAV6Iabl2cy1DOZ
fhqahcVYO0o/cPVBYDvTcKjQcki+K2CwGbZ+9MZxnLfLdIYmn0+v1X2jQlOQpmaV
MVAEyVemWnyYTrvbyK1SgdJSJYq6d5hZk0z1TvTsNbYH1PxIRXdo5uaYcuuv80lN
stF19IxK9HDDJt0tIOkCPlXWPaK28lUHNhk5uMgriuqR0cS3B3niDpsO3Stvt6LW
/tzedTRNe+GkF50TLaN8/Vs19xg0nginDYLm6ETcRczSlFAgANwg+tSKOf07Er+6
NnQzk8jX8yu2Be0XrUTo3eVq+6ZbMvqKPbN5klnBpyRYbsqX3TqkbR118Nq52RWt
+O2pm4B9ovebi7XPT0qFCIpNJeVfzMAJYRrmspyxGUrFEefes29yAPe1c6XypSie
h/l7xJDDvzhoJodRBlnfGCDGsY9Sd26xrWGxoTRfqnze9dYjKuk3fqt2QIR3NY8p
8v+V0QlWdvP8G0eKMEIrlcjY6Gkd88Z/Ve0Y6InBpn/ntv5gbpDcoKe2+iqVtk7y
cTHWQWQKv7oMET3BIIKgEobsBIXrlEj7aDaZaMyMrBoleSlbVyQCsAtloo/gm7Wf
caqJhNivnMN3CQRiNKMuU+nXjKJzyc294uTzSVXVjUiwRc70injlaWZQknu3K2QR
nnc0WjOak5+Pvw8RoWuO6WuMNA9+Uj10nyX+TPar3TNwh/xOJz16s94awJO2WA8l
QBr7lMXUpqJDAZskwl/QFunN1s6anM7Gi8IO2h9cm+7dsHoaoKqlQ41AJUoPnfO2
TTXFdcDjaY/RCB3cka/4VC5AR3Hzom8tXs6bQsv9UX0zrlQhAnYUy2R+dbmnTdo5
jGuMRuhUYQ42DqKToOqhCdzv6FpEyliaTGsUvrU08y5xWAvo0j1g7Ig6e0f7BhmD
nI7d2pxEkm1dT19mj0T71QsXLTDWwYmxsYbeAFiY/CS6UW/zNngsd99jt/Sf5onH
eIUtQhFzl4C1MTlRqM9lgCF/aTTIiLn2wkMprUh6PNzdtaCAiwrE+w7nXn/S+YYq
YfR2jQ5b+VvcoxV8UR3MjzIWGOilBOxpGSZf1FPCaW/fxxcLGjMLBnnrG0PEO/dj
DCVOPfZDPc/DDhGSl3Lj1NqyaXORW4P2AgZ0XjVSclgE8xHv7iuc1f6N2iep7dEz
UjIkPv2pU9CKgI1iG8N4fHfZcvaRrJRanqktP4AZpBi41aKWgJ1P+sIfyyZRYI7B
IS70aBOJuyKqDUbHZgTzKaFH+S6gBykBviKgzL0XV0wT0XmCmK4QsEM0/+zVT6Sc
DtbbYPVJU5Jd+2UfOfESLetE8rnbMJTKhfDrEc6x3rCqXoNy4f3sBgxg5UKkAjka
lKWzXTT/BUYG678Hcy8kZMsaTjxSoTTICj6I3pctujbvYnCgtlPQdtQCbQpSuM/R
wgLr2VithYg/ur/5525lPuFfj0357RaQVbQRJ7fK/1K5WRPC3CrHck3cP4k0cIRa
gH/Vrud20x6e98qOSJiEYFr1vqrUhgP6Jm0Vdt+j16jXNupwf/9EtHCMBjJRWPUR
5/+T3FH22S7GJemmKoX4lxHxItdz6xWD6R7f5gPVEIZs7s0tLtB2PXlMtsytDeiH
uMV1xFkhucT+4WoJCCqsFlMOxvFAtFchl20F70KcFPw4JOxw0InIhsQ5cq96qKez
fw3R48gVOfzwSoXm6LRpaDiNkxBkZM50WH/XDu/I6A8ArWqH+5/tVt4BjlvR/rV+
OViuAPYIp7bizJsRutrqiN94gN17R97Na3gRUnQaj6GDbprKY7MuTeQMUrsVxxYF
AK/F2vz4ZxEgEZralXhbrXZ5tZqsDdZUs59RwbtyXIMQZDgdPfD4xfwWoI7eAL4A
+CtsLF5R2rppxA59glwiyeitWj3F58uGy1wyEN7jeT0+QSQUICUjqweHApwpfp3V
ap5/MMlcOwKsxByKKCIiIiTzR5ksVzz45+J8hXE92ny6VP6U7K+kCSDE8Yasbg9Q
yEqFnE8yBCYL44dTaYoODq7ClrSFNS8psRQlM38iKqGwpu/yeb5V4T4o7j4OcxoM
cWtOR3132dZF35d0J7lEa/WHgksaSmsqh0J4EFV3J5LjEh4wIDAbV+FrSQTmOqDZ
MB2+DFgR0fOTS8TJY3RzicgMWSy5TTK+s0OPz+GvpXxB99U2OV1UWp5OAcOCV1CS
TzPzoQ2JeD/MbN1wtlETpYpdb5JtG2I3Vr8Hdq6crtnqNyzzLUwQ1fI7uFUFFvDm
BcRqwFI55hYn1fBle2vtjyduEnsceYECwJDchpIWdcbKs3wYRugF0XgMeciUr2Zv
A3xjsNabfU3MfgkFV33m6vKkFi74mQWNOQcasaKB4K1wMtzYoqWsAlNTLFiVeP+R
n4NSOFuX48dfRIaFdEG5663KwNDEVMk6pFikmg7mQ3CR/9y/l3QmL8xJsIvmKcKl
2DCtOxa8Ni3CiyOKUTpNdarmHiIWfCjwBBbiro/f7im//ZfANetw0QXuMY2RWgqt
vP2WnIsDj0gb2cMStGW3t0ZEifiv7pslk0LM7FfPS+Qw+onMfXVuZM5QJtJYalgm
dqtXQkluuxnvaPDexamRPIHSsGZK+OLH2vkcpuGB/jlWixxuRaP2f4R8ivsZxfj7
eREk7BY7T2XEsBiAQirlSvchPu00op5kivLGIqu4UVVhq90/ygMWhM+Fbe6Dly5q
ZqfdTOjabLRSuntYSGIt4G6wgPkkpTnrTkbnxWN6DZvMdHmt0MrDoJzruOZDQ3Ug
VF+NSrCtlZzR+xV0YQkL80w+axHGWafrxrVAYxM3dMOWSCW+1z0E+Xvsf9WyrXRk
Jdd50WETSnXgH4xik48TAQziJnmvx1A/D9RnkgaxyKe8/IDdIWqN1NWUM+PHP6pq
/Wh09DnbyWf11S6P8EJ4gXum177UxT5lAPMsir31qQaaw+pNIDNWJiHlEinbKh7g
LrsLxjUIvfhIHcxCZHDZPo9vmYNhqXuvVFh92H5B4enNR94MJvYvRvInP7gNaLOh
lUSjCTW/D8pgGQhmpYBLHWL9WPNtdv3Z801nS1fr7HesI/dLZNMsylN47lW/FFiZ
j5yJXSmlLSgNU1vfZs3gItOb25Of+RI9Vd1XdXda79Ydv5rC0xzLkTe4kV3bcYi4
vzQWDib7uL9iPcErjnrbVK0DIcFW/5M4a5s4VZxJO7uBvF0rmsEMspq1ggirN0qW
T+Dd/FskDOTzvwktprwr1nNSUL8yhcHlNVCcEisNVGhtnACFYyDJvCG6Np7ruBpK
tMM3AXbSPYBrlJa1vwDKxexh6eBCsXpXZhtokbpdIaCRqdhlA7dyirdf+obij0M4
PH/0s5obxtWm7a/FQUYGZEOWYc0w5FqPr07A5tP5OFJc1yupgpLPLCFSJ75qWG8O
woGmPr6lhyiedFjZPaIiNdhTlX8hmqkMtKIUeEirRLiQWcGtkLLPiEIdPdBdRDUI
jbURqqayAT5kJQrPXJoVONpRTg2I6fT6vp41MBPnXaxbgaV2Hq02euq1mlAhrdAr
PZLQCLSQTYiKXaDLRPLtjKUaC4TIaGsWXpk0TFMgxEOWN+PczvGUbAJDqN1SLql/
DBzKznQDoiEzoAMGeyueCjAjUwazw4Yo1bvuV44F/cV/uRmP9jivOweyk7L5z0t+
UXd8zNTfBkkahm2WYMa7H/SGfNcXTM2uaYq3eu1/Xi2s7HMy2vw0HZS9kGXBtsbB
1GvB6LVDrqrPrlwpoF8SdiS23OxYECB7xteGZ0lqGhySgyzOXVGcn4VGTYY0AkCX
an/m41ymuova82ZRiBTBr2bzL++U6OMfgXYxi+wustVtnsfnWckIajetQAkw3YR7
H9GZ6A3nN7WQd9zmSLBUSnS1PSkGr2dWlLvZUp3e9xAyrDRY3uNKS41xe8qXKbaF
appk9mq1X9RXohaKPkotSaKMjQoQvCCN/7uXKeyrziCjvITQMIVgOO3FZvx3nTS4
gDHqX3GRnDDdRwMoX4mKNlJx6+uWT0Rl/igBO0+Vxyi9bGemQPwYUF3uyN0nPpb8
A8tf5RpBk4MC6Y2kJaBxeEo6Oeyl+SOGFmaCBoVF3inf6LeK2lAoQC0m01tDJqDH
fFYiA9OmHi8CWAMAOCeT4V+NXPkeA5qZ+lR2Ad6FXQT5HWFO90qnSpN52I/TnTzw
Kgw3sYQIKo61TknTmbrPh2Pyh0xpNDBIK/nLgDoBz/ot2CUdY95FvB9MtwUrLtJM
fD3tjX6vmPQ0V6fVC3LofclM4nFB6efaNKeHCnnoEHeVqVGCaNIw46370H6/CBc3
7YxsOXCNuGDoQb7NhRwSeD+K1Illc+juwPh43fImYC3xFpqb10Y2E55hwlUvY3Zm
1GbUkPWI9hiAR41Q58+mOUCEePd0g21D4TGAtoesQTJZ9URFaLIR8PxYD5jDL+36
hduELGCUPdrup9goVOq1ozSyzAWO66kgq7EnWl+htrYIypss8pSMPnkTLq14LfFe
iLnoH73HxOBaGFhGZM9gBipJmgCm9gjnB7MLnTBe0Hbipvy6xR7n7SkCYWa9S9Y7
gLM5Td3QFrh89pHgD1/ioaRlzU78TUr78uaQ+Lk0AcCAHR9SXmDcwn8z5HuHuPIK
3s5ygEpCu3p4+7jXr22q5mRxs7yIZnpaFcq3IR/JXi+LCs6lqAZ2VPsTijYUKkp3
45ENkQJpzOyg8AVhjiMCas3/W341qzBytmFBnZBfuuGy/whmT5H9SKvichohuQ1b
5dRdJeO9t6mZwIvRSq6K5L9Gu9fgcLxY6+GUIaTBg92QXQiZ9ShPx9emNemlBg/0
ZbKPTIxc0Z8oa26KgvlqhA0ygCH44CgdlITo7HTt3a6lqBoPwHuQIMe5xD/3MHQm
XT/sU3pybR3qg9gtMXjrOGtNenSA/hx61Z+czAQ/xWnI8bYeM5NkdeNmA3ycUXcW
N0wX6+8FJUlT6j8QeBDokkBTsIPM82t089nnHyaLL3/m0DR+rbmOPKkv7jcy6m3+
aOoq7MeYTQSTxATd0MJdh4o014WW6Jdoc/nVKhPiqC6EA2EgdlJmVlOOFf6sCBIC
rx/pDWKec0PrpXHKIJiwrToKVDXPt4adKLio+B5qyUZvtSa6Z/esz1UoGOuyRnkE
AGJdEHMwIPUF5/ws53gIGbG51cQ5ElJCTwncELrVqu1C8ciWrpIqRT1ANZCHxsfC
KXvDftAWCPgTJvVnM2Mou63126fAa/GTMom407+5AxSyhRu4g9cmQ5A1AiV/4epJ
Jm7AJCWg9y1VFEFSSDv/WZE5RVMqZGnMZ0PLA6DeAk8GF7eq6CVjZbT9L0NWzr0H
Z7a+EQJ/3dGuFjvMExBAcZqa7rftxmLkU8bSICnzjA3hN87hwH+GBfyCueULZRSl
LycCXKb2bWMLoE+Nfk58nCjDTRNllBExhIrrH9s6cx+YV/5XVGO+LmD7XDe7dn+L
UrUDRY7dhi/QXIaK9ReSNWn7fjzCXS5a+apuJzzB9b2JySihoWv3Tb0ASTgzodJ2
c4KdXGh/i3WFFodmfgovGgl24N+18PnPzE1t3qrIHuD4+suelKHgZVXfmvlcyzo+
ta92Wpq/f1kN7+Qi/vrwRFKFIMDKvcNtegTV8XZ+FPiaFx0RcEgKBwDYKesktGPx
7+DuKWvN+gJD94x1bv55jCSlWksB4Egh1Y6SnWdw44RfQkWz7fhRQvB6cJ+TWyEG
j0KIriYOME145q2Tf39UbZElpMcQeNESZVoHBCHRd08b+XVJfrTuNK8cFrQc74EG
/jfqBkoGIJX26ASrJ4pCq6Q/fkauBTkvn+LTJiP5vH5ThGLE0RVVgo3G9U29NGbA
G+lhSh2e79LSWfL52qnG08+A/ol5Ox1ZYE6p0ZLzHyJva3R0M9h5oSngCQKVHbck
UkG1tn/3xMkwngAYqR0UpPtSkHU0ltGDRNbtRYIRuaexRGAZWjaUXTl3NsdNGGLU
fCAcJU5fLxHfcjvQvbN7LT1NTpOV4Hn4yey8uWVn/py6A5i6hs1bsMAlmiyzFXjG
gEFoqWpe/zK+yX+9veGOu9AIzVMzV8UkE7/J6MfAL6Rf3KdZAkZSLmXC9wtnYwVg
NRFJHxE1IrSaC1ehqzVB5I3g9J+fo0ocqwwB1hxfdfS1sOqcdXROliPIGjciInBP
EpMNf3esg64w9phndi/KmmxQsXrTJ8Q+79Wmvf2DDfBzIpMUzO8El3Hj7K3R4l3Z
IKLhfZxD8y3heAinFuIPqxjOQydd576zvF/8RfdxPcpV1eCKHLu2IJKlbtl7chrH
/olq5dtnst3M3b1eFsWAb+FwyjeNEiyzbRpnJKWz1WrvG67kcskf+tgFtUE/kYHb
3LjAY0mmeapLeaSsjxGdbiVOEMvVbyefZKwRTut4J60zFOAfysEbrrPADC+Q00yR
BOnA4Flw1TZ2WufNlf2My+L2RxIGQP0c7Wbp+iHY16OBk16bTP/imxA3n6LyWJye
b3SRLh7Zn4MoRnOZHNMiGQDotZnWwV37Wv0hBwggYgr0PC3t1tIuBDX8yErfIEsx
qlZRQZg6J1tJZxT9sp6Vr1NgAQS4rnIMebaIHcDH6NlCwCD6cULfO98VEmkNamsH
10iSa9OA+3KphOhlrC6wcyBqr3Sp5nN0+o4cvNtYlTLq6jnWKWsXhU0EyAnVbsic
3HDiauffzCc8XrHhmEzq+i5Za1CmABYCFfpH/e81h5GXo3i5c1G7CpjM/LRNhC6o
TUQXwP3u15vN+cu9yYBQP03coX3NBSku73ij+ZMVMybI7wqxREIBvBmNcftY83x/
MYZx/fT1ju2bxs+xob7CMy4OkdK+XX0DOmNqVUYc4/XGXfFRzJGVJWuRHynGj//8
whOzk9srY1Iu+enAq6iyMOl4R+fPKX1EGuub7liE3t3yGrm82YCMLNLxBKJ4YhT5
ZazOyGUKccJtRsE6+zvrl9WGOJEA5r+nc7QG+1Cihm538o8MbhL1LHWZm5wA6iHH
yGBvQGUpxIMg8nfwps4/YoYCGxeWAf5AAaS8uG7VylFfE+vExUL3wbSw4v7gEL4J
rHWEF+jVv6g6UaA0E4BhwtRkqFMZMaijF2OLAKKod6B38qX27k6YmXz6fDsX/qBM
91VLtQAgjWFEOV28s/opMg/+B8IwuBfBFD40QiNFo101YCc04WtTWbojVDwIPW8i
xRaEpUbPwPTHPhG0P/8cCirWozEGsXDSkPY7XztsgNEpr6Xd5McHi6/neKvnG0Ix
FfSsIuM9h8g3OvfCD4AZhlAOBW/UyLC2khfxbDsbh0SjWwlIepbenyPEUBmJh0fD
PtAqRoH5nDNFL6D2nu4nZ5sin1H0m0Bdcc/TYSxld3CWnoT0BD9K4Aoy1lOMRVvU
yD5avrAvQ+Gbg211etDfU56a3jXuYIpR0oTyuqDmJp/5kbN27VAW3K0MIx7qjXWc
IH316zgRb5I9eXqZ7MfZFcobWBbKOIBcQGgNBwVmbBewxi+TNH9dRBXQ7klHY2bP
9XJg6gASYTR6FKkDmWfHRyWU2JoFewv+iC0bDwlDTWKInsGSu/vrSRIU6/VJkjCy
Vul3t5vntypnlfTzP36C3dhcn0UrcuSgjOEFi3mfrO6CfK19mBlFl/1K6FwYW5rA
2ff1vfZa3IjgoTV3OqiwLWHG2pOpgQ83cm0WJAthK+/4N3ek9jZMiWYqg2j4Epxr
I6ERCdNtrQqMPoTi9vhszTxs0R77dhkcBe/9gcKW6M5TK9PqL3NdOeWmKM87GfKK
5KObT39sAjY6vrnawdsgaGYcZ+mDnrFUXJpiBxrfYUfd7EepI5CKMxDvEqLOvihC
ue730QsQjj8WdwfPZJYMzEbXKIK6W/AJyx4d1jWvlsVXV5DZr9zRDAOloLDfQMbw
t/ha4e6fVF3EFxB72OypvuAW2GpxxR4qOOPE3muTF7fkZsb8teG5W7dHMVNQHCob
pk+UnCnZbrNamEjJITdpPVlDnAi9MZutlLhQtsH2cjBTvB1YcaYYOGFwdGIdtp6l
j4QZBufOgLeeAQFIi7ESkDTiWa8hzS88/0MiAe3FGFYDEPDID6OseA5493QKjlN6
DfZlfPi+yj7+YImNBklk+V8NrqV4J5iu6j2f0kWToCKY6CjxOBihp8Wvt/TjDwms
IOlDUTdO7rasetDEQcSzLkK6dcOMxE9KG/W73xVHbcuMSNl7J07RGNBvsUGR1+36
uaQGcdM5OLk6WGp6Frwe5e0L6HOOkX28Glwp0J6Uyhg3jwS2n4Ia/9kToTaG3D8u
eLOPVAWUB0d6Se3kMY18hMxy5wadDboe6XrDak0HdEp5xBGiKyRLDOaONd4lws8J
d+GdANXOSp116jfLE1rsFxL7nAJo5FcuYInWz6z5Xr2WvdpJaRbCbUwTWqIG/bJC
CKLBP84+q+hijnKM9O/DhNv2TsAJthhu3oXIWiOtLg35Z/5oVX928iPSk4iA3P3S
Mo6E8E2qtNRM1v7L9avWs0lgGuV3x8QbuO5hr6AZrtVjhNdR0SFVOI0ZLRvOV8zb
c9isnKHHNepzO6W30vfEo4f4Hv+DRERtzBUj3uwCqbucC8vU8B6pJjQXQS72jhUG
NVGX72Dck05XiN6ZzZnOkW48OaAswwkZtqXOqu2QU3K17bIF1U3+7RC5F5Q1qg2N
0wGXvjpjSYovTrhqg+QzKKqC+RRwwXNUyhVsHHifI9qo1Xgnj6J31ns0MWTLyir1
JtRSOKyEyru0pUGPuCx7kZFDbmlLJQS9iEk/VPjyDjAZuycY4ud/UipejDPJENY1
92cm6klVLh54elW/GFQK8TUT9X9az35DSmFEFRed5fwRKk1KRz4sYUW0K/ET7YkT
nNv13iwx3bk9td0r5P4Pi11yq9uNEHIzpN7o8TYRKzFF6WOkYJwFh9MOtuzd2Ayc
P/Z15u6vqlYbFhCGCOdbylE8elm3M01B6KfyjKymrfCPnRit16iVUZ1bzwj6eFls
BQ6IHnP/DM2CZbc58WtIBkWcR1ppKffDQs6gCYS3c6qcH6GIIFqOOvEmucK5hXp/
1Qftr8VPiUI72Sdkwl6z5Weu8F6VkGfhP9EX9czPhqGnlAkXg/BwywFM8nPzqfqn
nxmUMF6lPkbz843gMIN3BeiJ+CQ0Gsd8d/iIE0Z535JNHEGuIdFU+Ri/33LQyyH8
ySukVGyx4Irtb8C6S9jj60hWz20q5A5KnNSSJUjpBjP9MJsh/nL/elCXZvRkuxxP
WFgDq9EsIy7+GJ7rp89dEcya4VZtmUT7DHHh7ruWvy/0tpWCBiu4QSMkIctafWtd
x6/dnp5lGwTpJbb7a1bY9twNuFIHoq/Le9sEa6fT9U8/qpISe/5DztbaHU8t6RPX
JBAvdnAOQMro2ZypFIdVx8LgQulHUCfb6nqeGMH4fCmiuWHLwhL0MEwbYTYIrSSE
pKm1whRDJu9A0oSG87XZKNM+o/WxZ2B8o9Vtqr4LgVPTRFbNkWaJIsucgaUWHHsn
kmEIfcDvLRoJZ2EMQroMuLJJb3RqFJs9XCTHeJ3aBhKOiN6HSKAB+Qhvw277j+Sm
e1zae8ijAQUmgNjx1+ELQiWI6UiBffdJvUQEcc9TMeUlt4j7ZRuI1Y7+Q6V+M3SR
jlZFd6nQ7bXczfiHaABupdUysqE/HO8EsZYKpkOZQ1pd/VP26X0guGBH2cp3vKBb
k7lioffI8LuCqusRW25IHsNDKLU+sCVDMpV0c1fxeHDn1V/u2+h0XZBS9oz4VJbI
B4Ve3eTElXsNa7Uy7jaNDi3QTssGmsCg6q/iLdBITh7uIls3pZxGgpmjgekF6QEQ
mnoFUpeVTO1SFgIG6YqFB7pAfwj8F0vsqaXTzYPli2fJOgDVm9eIY7qZhxj5C3eS
PFpgIN6Pol4TwxLLL0OD7ZyZRsbBwtq78j16D21faoasSr7Xxzf4uUADBcpFbeXR
Xhzk9sMrKNLlBhMKBdOXN1GE35/aWr6X+EaUz7CPT8WCHjrF8+O7S1qbvMvigGLX
4YL53dV0CYPVE+8q1LMXtJCePCUSN4/5UwpNbxxvEdrXdbkVVlQDHwmY6U9/zx7V
sn1DE5E+CBXRaFanZHVTXRNh0cwIKHABnFl5uDpAsnmWpE4Ur8MENW7T14Qrb0hU
ojqOH4c2+0CjHPmEkDMojzvaNjSgfV2Ta1H7/SjU0NunjHsZmiLBLqRd5jbW8sGE
gfAiZ8kYg66TYOYgHLfc1yr5NCRDagQnijNE2NlMAwKvK3c9bTsk889uCbOliRgl
ZGMb8XRkT2URyN3D80fwGVqheCXO9alstWZ7vujUlvqEWoKn5YjR9wNNpghSisfG
E891iqGz50CmZq7w41cpk5wDOYqg3xxb+rvFxl8vHI/9765pZbGWJfbu9UYRCey+
uSqf15LWZOlvH1f2a7tj6YMScW35S13uRROejbUByDg//lvZqMy3JheB8AkvFbK8
9mdrsh/tvINuNzEsMuQcZvfIUiih4A9hX/IdlWthnZNLsOssJwHQvMuXqC68QHuY
eXd4WbqFsLo32NrYVSIArMWFLpd9+2bDiR+HxYGBp3FSbbUwlpTpGL81FtWch9VZ
VgmcshLgfLGfU5E5XkhvQZK2c58X0n5lespgDAbVJbbmkGUKhxrTmCT/Awv4Q/L3
xXzlCpdM0MePYhiTmdw7iWSyQcnW1GiGoSRLdACIxbuVYPJ5jZcpGU4FRZpkSVRN
DDMwxlyoHYycTs6+KTc40Tk7A4/EmDVpY2F46PKTJ3Ri6iicm9k9rgdgN8q8nqsZ
UUZPex3OCiplW6fTlTj5cjwFp7QkWHPGY6Sayx64hOJsYzHUuPJWp3KkBbYS2gwD
1lGVQRZuIi1fERbX3tSgnO43069eDs47U8ox3MoR8O8cX9kMOznm+WFDDjnlx2Lx
8NJBz+uGO9XpjujQ7bcLFubBxaKorFNiibpbh8H0gMZm5aRHpwRgF7OeiFNjk0PE
Sxr92WJ5Jfm6Mgd5D8ttZqgzlk3PFs1yidwFQdI819WBpkohAFy5Q1qw92JDmc3g
LNXO8xUGR6RuF6+6vnnY5IE1G5c1Wfq7h8nTuYMkKMmZ++jYv1vlNpCUuQPSRXmW
LvUJypfPhvEmEezyT9KuzPLQXD+kmpQsTpa+riQkQt5x/2KSVngMxqKPUqX0tOae
4nM8eZ391LNdNJEFj1HKBIJjdPjGUA89kuLGSN80ZqQol5eEH1s01dRtThDc6vdo
P9IVQIqdlwGg02f9dXuWQF4eozmh7Yax3ayE7qgpzLVEuuYT+m/NHZ+ooiUqUofw
xfDu14rQZ5tZRWVoF/vY7H4WQv+2ejViv5FxjkU3CwOUDlYoeaOowbxn0cM4AwVf
o/s6A9zKIAUzSGR8UETAXBaZ+ANEX6eDDP+cbiBvUM9h5L7xQuEQCUAWlzgeqm2Z
LkRQaPUVW2ENWiOOhK4hVxb+miHGFC6FvaJOFWh9o4JWqrM/ACFwKOqap30cwgaA
OsCgtoQKpgOtDDH5B4W1o2gWnsvyqG+5RSHZo2eygx+87XAKUFM2sntYzYrvwJxE
ncbtNENZ75NicxPbLRRtY/0/MCmRsOb9JewofnQQRLy/BSgj7o06bDZf33+tz5vg
BpUrmnuUpYtCd8Oq8pVllCeQ2ycAApIfD1O672/EFo3Lg9sN5ooQoKas/OEhfPmF
vRMxoOQGT9r2n1PD+0i95WfUHmYJ9bg7lrkUU6ckLPZxc7v6qy2Dnl6avNTHrKMr
wMRD/5pv76IMpis3ZY2kJZYRvV39G1CbtFvobrLEJaQCGPZOLJ4rGREzJFOlq1l+
IWWynVzlt7qhM8UEo16iZbL1Q8CtU8TUWVNYoPh6K4iUsxrnMKMHDToX2IQz5o+9
9wGzpTZCVjocrmNkc9Eu8f9mn8KsgTTs775aDQKzy8BhumHiRjqjpFm9CvBGMx2D
YrDbWb/F8uspR6uVUEyt7ztDF9eVTkBiRIVeVdEAI+Hst4tkivoiUQ+oi5gutyV6
I7jC/i7yCqSD/72xVnsdghSP/bVnkDX/2tgliy+sIYbcrOJpKqq9K8KSC+mYAlST
6XG3Ah8Rb2wOPCSWUns/vsHmbz7Q9AJb9XVISu+z+qM67XmpF1KG+IVeqNZFvFUH
m4viGe3hkwrt3UhiN7LRoJXE5Y5ZVRh3AqTezX101tvs6ABPRkEGwy2lMT+HrflR
6o/ckbw6B1Vl1XBkkFfDWYS58KZLWKLIYcsTIiGXBiDsWFyKn2voGLwXNIuV9W3f
Ohl79hdRKYh3/f3OZQWNLU7ZLQqpL4ASWvHrDytBUIsU2obS/vUjTmZv3XHokNI8
0yQEpWlE2TG4DRbpFd8EhVyxkkIocgB+t4A92Z5+LglXwXBWoAkwJI7/fi8Qjrbu
q5XPN9SmxBcl15BPWVC/pFb1aX/XeEPedtNG08CuXkRZ89w898/+QaJ+74D2APt9
KMfY4LiK62Oa8MQ5SeMiO+I9BDA+8QqewCvxLgZ6OBl3r8nArw0BK9e4/YtxXjcp
Ne8mbSdfkLQpRNm8Z4Xqf03Kv6MR8qPDi7lbY9dBMmcqpQahcTl3OqU6OLcCDCke
yjOldkzHZ7JEDnB1F0uWFCcaf5kE025M//UiY11OcX1I0eZPto/ar1pR0Y5BpvqC
GQciC5o5UxJbyfZk+B3c8yQ3WOfK8DA/acpo9UlyXT6k7BulsPJz1AIhv7m3ce3Y
HN9dOzpA3+1u9FnmJi9x2oef1HbiTwySk04xo8xhvR3pFMZ0m1hNyr9wlIO0N7fi
DpNdSRW5pJSoKki/CEy9zC9TWjGqvDnbi3O6mSX4H9AdaoOTRpjYHOt3SEEulllo
wq9q1Iu/XmkdyYbxuMbjB12FAN9Nnmvh0P0j6A086noCvvPGD2WfsvuhuwIL0Xkb
uHWwyIC7KusnldL8uW203mZY8VtNt8hbIUBdshNwzhZ53kftvGKhB1ZTlxzWNxqK
pE0iDadbDGSjdL5qVEpE0IzS6uJzfolYzXfviKzkaLmRwOfZBMYV5dQDalrNRmmk
5zYIEivzZtZSuh/oQYFozw8WE+Fzm22RSsAJGrOXdf35sb58Hqr3dn8+3r5ET9MS
TAuSIvLUvBVpRt5wH4s3VTMYJeo63tlWQzd83f8awBSPvOX8Qn259t4x589/MkEg
xANrVUswreVGdWsHC2zE1pRsNfPRDykYm2Q5hiyGSQdJ+PWXUDVtapnaLZBDoNN/
FEBKUapIMoDc+j4wrFdFye2eNkKUbLSLJzSeNTMcTTmFcpeM58zwQVp62YATkxJS
Zzv2hseG8A26/Qvmxoc18HrdY4mFKE15fS/xlHgqCOd/XwYQ+01FQFjFhN8R/RKa
+3SaVcbMb+pOv4SMEsGDO4PyRGQBAZkCv8meu79suo4e92zuyw/dr7JJpQIsbveu
/h8BDeG31utnzol2nLfD0TPGnr1pan5mAuT847w3VR8/WCGnsSotROP7QMgzIpIg
XhFEPTw1pi4daCL2RTetpq6erzqajpS7vrqfUUHCYRB/u0YuCjsc+YXcDNqZWgSP
qONxkiwwLRL3bygc4ISMXxKWuqRC6npFLLezRKn/LN3g+Wbz2DtfkRZ2+bFYvGMF
wsmWKSKBImAVA82C2ROIdszaXTTHOPl6Hg8Zq26MxqSWZyZaduBOBf9M0RkrzKdA
VxUzxPNB5WwUCFzSM1GFkDJvJpzpsZbJqgAuoABYIQAmq8zTauwQdGh6fh7OCICl
qzrBJUHRFrEtrAzC6y4JAusnI8K9MtmRE3A8lj46VAL+bBQMlNCauRMKH9qxoEMd
thjruKIh2SQkNwFnI9ApANWPDgGt/xrKIUWDBci5bh9fH0ZSCQByGmZQZNZVY5im
/LOP6QmV5gFy/OhuFW7GUhbvXjz7ZtbQfJCp91+tMyCXMg/e7/UQYLV9nU1/Z02N
o+3bWLnLcT0ehH48WscT2zeoDFMofkbr530hFanomehAC2PkEHiJ0PmByfPndCR3
JQx/r0dyTr7WwnzyQPqDuARCpK7MdMY4+3FbiI0sqMqtQr6dYTJeXikzKPfAjAkR
MYQg3NV7IXE53oZrpyznUghBOO9NlKgul4ELo1+QO5aaCEZF9xmJ3HD0xEO357af
WXsgWncmH6MzfCHD2IFkXLtIO0WI/mRWqMLnOKoXJxla7qj37dufMfwHB+JJczk9
cezupqj412cAVQXDIkWixA4Fe47dMK+T9gyI9mbiTekYihwJ819H6DEqO91fO2TR
+0PLbLtxCUWvtW5KW8pj3MJrE59JMVmoCrwkQBfPjH5elT7mx+5O2/+35OfNcy+Q
eBEsc9uFzS//f0Hs9SOPqYkGYT4YIPvpaE9WUz8uOrE/ev08ZgXPXnS/X/F4u0C3
R6nuhcBDex0T9rePjDw213xZiJOsogKLsqLL3JhTpTUlYIUe+9V+ueiv1yfrzf7p
4Z7g+lS/QhNE/N4TR3vHqAOhXt8OS1wLFmPNnUXyAtdxqv+IlhTOJgPgnKzPN86s
Ovy0aCJHCOsEh2hIviCWvdSvVv8xwmf/ypqF0f1RSWtgBloRLqK5ymu8ejg8oKvx
ouG/QzQw2uCAE07PRO0Z2043ldKPlUf4JugSUxXVNpJDqenF6qaUIxrhEVpL2Ekz
sfEkDiSs8EMhgXnKt4sWOEtWj7d3ArUYQaRTIKd+oAoPX8X5nAP+pux32/KHBdAj
fx6dKETMIzmSn2Clg85OanswinqHtW3OOObpO4BAGWs5vtGENJav7qfSB+gIdYG6
k0aSxxHYDs74GPkbFJBaG7oKDSK6KmawlNwDf6xwYkmsHOS3LZBbx8JTajq/S4AI
ou2+sU+t2HG4/uGKJhyORDunLdsXP8oF4Fi/CpWMihIN+GC0tPbSgpM6pM1HKaKP
oZu3Vhpj6QS/UdFkEJLk05StF35S7VFh6b+UGiHhU1ifRD5JS/7oXwiQH3zbKOEn
wiFe4+m0dD3it8/86ZBGqqAM4xVOD7ZGlYR+6YT67KeDmeuP8mH1I8iT4t3/Nrcl
2hctJ3sR29P2HJS2V4/R/ZNB5hYdTXOClXZEMk/FjskSCQSB9/RmE/7ZBciB+BHa
atESg9cZXVmf5lC+kuOJSFdR8FGi5ugFoIzhkgWoqtf55jVImCVEYNPUyovdDzRG
AkzpvP179CY6DZ+QpMJJnKKrXHa/Zoyp7RijPjbWrZHYmKuZOZL5JU/Kt1/wXI27
n2PGyoGexl+8QqooYdQ1/rNbk6LZo+pyDKGy/Y9ooiSkFl8QlkWQuZU6LKXgzLmy
0TOjTGm+gQZZ3Za4T48fOI4oG3/ZhKBsgP2IJ48KjSCOlBf7k4pR1iNUg7JnSDOW
dPKftQpPrGpGO4gQRp+1kEbNziuzEeBMBiVDSY0aWMue2J+OHdeAJU4tDa4Hx0M8
DASZyAM09kHkjCfP895uryLkI0vAGN/mBuO9gARRIb2/TGJsgXDw43ZmXIadLaed
QGTur7S5xYxfALIzvo8MdbnWgNExairpkDLI6ySeWkikSmYW+y76OwjHRtr2VmtG
4AmLyyBDGbEKZVfZGC9jYYr5G8EEfKR9gLp+YJ7x87BSFh6Y4rFiI2YqG0myLkHI
V+V/WCTGtELHeHSpLvt5Kqn2xTJqKp5dYNnQsF1q4grhLFOhwA93rpNeI2/ODmMp
/w+IqpUdVQdiCwjld1h7t7CfJKt1jL5h45VBOStvztFGv0Oh71sMx8vKPSAWqRU/
jzB1/cYSl7Re/g7ANFVUqaSZLiGpLXtOcUUU7XAnkbDd607tRXdxWvdAjihA4Hck
WUFFBVJ5zJd/veuLXy17XDjf5krs7yKfbuFd/MAeCebJtkRx0+Z5LYxBfYkFC47c
AdvKFC1xgKQxFQMglIpdltfgJS+Xv1chUbml0zR8aYfkawN5BXQxIuBcWzAn2mi+
iRycbdZWkS9Di01mCwLnpX1LiXu9b1UJnrjfn2lL0VruWxzej6XAh8qY1w6e39mB
8t/lcfYzaUa3ZjaUSVojBoVAofc0OzZRhXdx8UuJxR8zsTSTXDnVf/trux/4KEoS
cXwzmEJxaJlg50yYg2VyJETgdj7P0JFWJNoby56d84v7lrDsCtr+8TBXq+EejlPo
uSYqYZGYNKi44h9KozinYZQsDi+Do6OONP69nd4ICW4pOuWDxPLrzpSsVRxsoKW8
r4gV4SXu7acXZyYUImOIB3wzY8qi6+S8tiIHtZqsM5WpGxls2SL6FiWh97wMgmxz
329rWhOlkrfZEl1DTleuffzOkeDzESEPZkUi+bJAZNBjgVNwBZHZalkKEmaWetlO
n/7ofw0bp3lzAd5fJ3w8I9y+DW6IFtSKPVXp7Ub1qE4db5VXUwU0Mop30lSO5JwV
Hxb7aIBnJ4B+94R/sWFjE5jCfFRUN18kyci/46wDZKrXJq4/kOEfiCmcntbj7lBz
7H6Db/vPUQ0wVh1Zii5OZOd2/xhcT11zQADdDg1jIhCUd2zzW29ctD4PvlhmAANs
Z4AX0l4xNXpgqp3k5gPHKSXql7RuWG2AyqmIzvgp676Ff+EmoMRylKJw2JLjAg5y
llEgavGfTPwQKP541glBuv5Vlxjqlsc4jXmychSFOym2xEcAVQk/XPNcwQJKydC1
Strq6WT0FuOfnwEynqCEgTBaLNpTpKSgU2PG8Cpr0uwPdFNEKwsmpY4iDGNuzr9r
7p1fUO3nrRhkwCBt/UsSE1XlC1Tj3e/6baA/K5ur62WQz6F2DCPRFyDCu61YM7T6
OmmZcYwPYN2joyQ7KLcLT9fst9in4rZAyjXD1s/2qZKKUY81DZWzIXC4JN0jPdMZ
vw/Vl1jwNxKVGnwJeM2XPXbW7O1AF9ISsxNFeFm5qTEQF6Jhuf2c9cSvmkElS/Vo
Rew6B+qIEIiHo/vKEn3+vZCkNmawTB6xVSt7sOFJBbV8advZ3xNqQ1Ahlj612M7I
bK1XBvA8EA3kOvwaaYts5SVSvIH5Fhm0d/ICSMA38xQYU9kmdpGMICtZLZl40cvk
a1JG+PZE6081AmDTrQL8bd3qqCVOkgGTCWZp7i6Uvk0iQdfhB1FXWI/RDXZXhzy8
TLl8UDaP7ESGagTZSHsKgacE3DuHlVvMCWcD6ZfWSnLkuqknH50PRn8Dy69GtRDM
uAqQFKYDwJlu/J3jJh5d9DiZ0ouhDCkoa+9+i+UdzRJeiAuIaByKhYqGjKCnRptc
eWYipb+tHaykfYjmYmpe3yHODz5rxSbyhNLtOjrU0d8PnbrqwEtya7YGvoZdgXYC
Q4Zd139nhUeuZY5XJ1yesE+j7yGwD/Yqyj0HRnXRQ8JRzfisGeHjYtwcHFv7+jiW
wczS+jBi8pieZxJR9orkxnnAOWD4w4ooxWtu+6LNqY9bMhDLEb4F0lHirpFrjfEX
+Q30sOyANt+ZofTFqu4ZwjLGQdemmMY5EtpYQrtJ+3YAsVZaQAp2CZU+R/jCwO03
QevwmH82IGOVAYRojXr4WWP9KN7ss8QnKYtsbhTYUlHiLAhYKpQ58xj/dXFZ8mMc
nJ41nlJtC6lqsXLxaVipBn8YxHRhlKo9hxe3opVc93k0F/20MqsvHpBBeSuwyH9v
Xp5skAjZwx5HkUIntvPC5oGEbvi8kIPkB7dZdUHEACyUzlXQ9MP058ixrB9D3QxC
5rHqHxG5f6tt8+XzbHfZbm9fMvSv8ddlnfEejFBzDJMcbJ4NYKaPzL1X5zb6FrWw
51FLCwsVFXx4RKmsm6ZfXYDPbNCIgTZcSQHuCNvYdJBJcWQyEo64dikAnyfWNVbs
FwyDNOJMf7btQgXAb0gwbI9LASoNKNKxBYsUmnpbv7xfmSgBdyy0X+wLIMZNCVTG
8H3kQPZ8XpSu0pVotcL+1e0uYeCtXO14MqUKxPm9X5pfmeogzt8af3VqbQxnCZI9
OpUrMjZi7hY6QPNTMC3YOorIWMJ8maU3YuTIANkLs1/n4Nqsh+JD0GSdTLmZ4qWi
D2MaU3UiGm9Ggn/JwcRfKOYQiR8lKOz8ybestAIxnKD6uvoICBB6QCNIGOJevhdQ
9ySvGucntxDzi2HqjIUXcXjcTn2QUouiCpJ9w8yazaLHverOR/+b66rbVKHIf+u6
G7rBgfL/P1sjLgZpnoNzOg0kBAfAf4P8KibLEuHDz9i/jo4nfoKPjMYXVl1g5tJR
el7r+JPlwPpKEtjCH+kIfvfTIEYIJNWLIZSg9lQGxGskr1tpVEbidjlvZs6w3RfB
0p35Dn5+F/vM5CR0A/UlSL1JHdy0XtOFGr3cxrdESD2kLG0gH2dDh3cV90NO18gp
JbQwR9q7rvHTEkpdJ7TaWPddwyFEAp/3VYw+1ER6uWjQYYaIi0QkkSOkxDD4+9uU
K+9inWfavu+bmwjB9QCRrMMrXaQTwAvbbQiBAdIFqiOreiquRVDUFllpbpO8v7Rv
2qiyJkJWhFbr8YpRhx+UMsJ7rlbhD1DMC6BnOjBgOYrB+Y2Oi3o/ERPh4zR9QJ0t
s/WtZxXz782NJBzrraRDoEtXWs1KUQcH32A4+qCSdW4TdU0o95YKdElfp/ibapcK
n8OSqhQFEBD9tlpmSGiNXf2EOItBzaSV6+8/9CkWMWD7NFAPQY9Ocx23xR8UmgF1
KSn30Jft33RowOU3oZA9bnhyyb1qDIkrTtPGN3wIs/ogiyz1v8XThYvejb0Z4vWw
flxIbVKNe5MrQag+AOk43Caasn+bp+Dye2ja+B/+wrQkDoCfEPm7YiuDgBZYqFHQ
1WyBytDi2cvbWkFr+mxxiT8ycRn0EXvBkaCPCQ4BcOc3u+vQC0+lHkS+8iLmcmmV
M4CA42mK+VAygDS66Dec9eMcbfWLhm8i4FY6jFEM200ejI/0UKxJAuNVxL2Y8+8B
hinak/uKj0pcT8PScPHseb+dBzl1KN1prDdFw9pzPGkmgonwYcvcGBLvenxJqU74
RJGw4nOyjU5+9sIPPcP6/dciUP7GF+5qnZVPxkFf+nxpvewgBTm+pK6WX7eJqtar
71k4edP86eWGvFEAvz+bzWAA1FkxyKJY/J9U4retfosvVysdoHqfxUbcx/OGr3l/
8tlB6EUdkw3jwPxNDr5bCM0Wwyr0Dt1GjI/lkL5miIVPEYRa70imygYSesh8X1l+
b1zLsb7oB4qim/0jMj6rKi2tCWJcXIF8G/jW/Ph3XznAcPMVaR49QhUreThhSkCI
SqCcYdRJt5GT4yXPgnTTOP0krxQtOC3eQ83tbhyKgzWmMSQj0Lr0Ks7ukphzzfK2
I5x6uoiLI+kQugEMTSUj99FpRZ0Fp4l3IeHE/gtxJtys8qDUPG3jc1jT9NrvPZVd
dYK/3YuL/rSkUT+NjSLdEJA/IntypWGJC3HE9xCLb/aLA1e+a4ADJ/GuEQl5LfqB
43ftMt5yP/Psyj4NEwtcePw/M8NUNTnAMC7yCkZiP2S64vwfP4NHTJCRG4xTA6C6
FHF+PJYSds7i1edWJEP/Lp0F/5yjQHurZ3IGZVesySwDfEsBJk63xtzRVlFubO6p
6dZSjFEjvAGlNDIK2s/neUgLVFKfEi216m3kP5oF/JHNbhMLdTi/oZO0URLZE3G7
aJqGrWOHYgPWmd/+KciFkxN2H5tkIEUeZgHIcJHfaTt7FSF60pgvGsiNZpKLi/60
yu3wl4bmUHnJ9YGrjt7qM/rjD220i2ETsDXjPcv9+AGhf7+6cF2IGpQBHDJnCvNc
MAFfp9DFeh+RaGYqZfyTkPoqEIHeI5q3ZDush+wtKK6pZ40CPKPdt574AqWkZrDC
RKOqas9jAQtBvk//G/YMlP7lmUqI4em9knIJj/CgtktRulmN+34RTpz4pFYqaFxB
V8N0qCzVKOJzbucO2P6fyOLbA3QShcyaEvTY2k7393JHzE7xnsQCPojp0SD+3GJR
Mz8+vPEeC6e9Pyk2pgFa++5oPfP7RxG0c8t5g9vTJUGQkMwI360zsf06uLOe+Gix
zvtWOk5ZVhr5pxJcR8O5yTgxCPgQu8c7mMc9ENpkevge9TMaoDD1rBs1bUYv59tf
DdVQqFYVf48MwJ37eExBLJIfQXhQ64L+hUJEeS12R7fmxluGhCjM6ANFath3b5S5
rhGxI3C+YkmC3GIpSD5JNT0xIqwPBptDmUaq0aNe8+/l5bFB3P90bWW5tweOqk5O
zkDen8jlL66568GrX3POsxdsq9AosgA3XAzSH7h+E964pxpH3xNQAdbTzxf6Pox2
jCh3jawoHXxfpszmo6SprFxMsuqHQqEz+n0Y2kBVSn488BqHSzb1L4k4y+EA4ygp
fOM01ar9HDW521ZCNVWCZeLBiyUzMnWPMvVsF/CGidTreoZeKfuyAVQzAJfDmXK7
Z8hCuALnokvTBx3NwujIdyRUgaAS6YzOL/qLYzzrd5kkuEs8P0PYAApaNN0tlHbk
uaHNJohRfvTRxZ+jKEFqM/kNDcdgVumUuCxFLiyefa+bomcrUus84JAzsJj9Wo8q
h86Y5t6n9A/UVnOuhlZwRVmswfa7UysBwCyIcISYrpgkSFKhOhNjn/W5epsJzZJn
Qx2abqZK7pw88n+/nhu4X2nVn12IiFNJRnrr1F0NSWJSRjpqPvdUf5OK7+7J73xJ
6w+wrDtaGRp9j5+RtuJlEkhRLcsnUaxGK/2v2vg1PlWD3TXIjQ41IdmkDijyovYP
KvQriZPMEs7ZI1MW1UDm6OsurfKs8wNajeTtL7YUdwx9wI4Ij2u9u6Eax3myYRqJ
xfdcIOdz3165a/CJDMghk78YFOwHmF6Rd514oZz8ZzUpnnhCgqL0J76OLFu3Q2EZ
4/uSZ7/7q6mHQQFe7JeZBnf+NTGNBPHoTY/YM6DrfE/nTIbFKZPhLqzJovG2jUlc
IJyQutvownqrc0LPLbHc9E/QxFLbNYWh4vAePiQ9pvN+txqrCPZfIousPxPrPjUw
zalC5MbEgc0lHjwbXe45whVkUIRwrieqi8GHB+2IVvt0vEcV/wxuy/JrFlCyPzpj
jQET71dak5dGVHkOb1TNRmzs4tHT3AcJzQiUrB0TNjpU+rWDZWt4JcXd0OLX5KrA
9CcwhO8J+cNlyCrBAcchUTr8rfBiyKfAkwlu+pArFAtIJCwg4Hmuc/gy4iNpkwAb
R12t4xkcWF+tDFAkn6ho8LRph+HGiPZ9rGoIiaGBB5eimm7bTssB5Z9vdycLdCpl
muCmRw9lA8ezbSdfBOwQyIT3c5+7J39KJ4keHWw7EL1YKjhaspYfcPQERxGrfrWC
JdI1bQ6EnPy/Uyq5rbDvJVkzS0BafiDa++LuYoTBO51NgHPC6f05YA7pkdKbWxBE
ODuIkQB3j7efhBX96F7thrv63E/vcmJxjw0szEP4jar7rftkf4CAh66LcLTUJO+i
UK8pvXkCLaR8VnzhhjsYxI3Lav2blLPOnoKIux3dgW1Ri1yFduCm2RFzySrDKlYm
pttN1fRiVAM3XSKSG74TlEP+OoPpy70idq/Y5+rptYDBHPZl0/h+iYLzTQ8kp+XW
79obONk7zDOLbjWG0DUaiT7veADOmD3pvpP7UbPuUCHFm4mpOZCOHfGahFvR8wBc
9YI3KSlSukuJILuMNeJt4k7gaO7fW3n8FqN3U4RfmQ40Nky2q3r3C/xdu5HlH1Ui
NVRpHhHyOj1GggTPX0BT7du1AqJ2Mw6Hdsim930R855K/ZVVvh0snxwbvzNlpNKL
PpNUdSH50KW7X0w3KyjLtfUqZOc28GGmYUpgPbU1Ym+4pB6L5kSfyR2iQLZK/sb5
6iUQUcQfxKD61nE94rv2b9BhdtOmV6QSMbAJsxgbJKFuBEKeJN681DFZEHCpbDbo
mcR84swUdLeWz5BvJojtEzdryG8yrCZqieOsWpCNZ86NzGmyDGsGQv0gEUUGF89F
RqTEJloUELmeiDvJlnFegxVJXOEZxier4vWrJXL2g9RZqKj57uYxPyhy4MIyEVNq
Uc3+3GbBT3KBaQEHFj/PlCPZbB+xA+IernEMzrHdUZJyLJFNe7ehlLDTQKocdt8i
u7w0XUGMBHFMS8VYqmIzdFiJYicsq+BgT9u7xgI1I6QaZPxH7Qq5CmoxwpnjgHgy
OgWCRbcEsK+Pzm4jMw+9e5RfZkW44UE0Qmh6Zsf3WYJFUKIxJkcq+JbOWqxQ5EOZ
in8S8liZm3rdVKiosYA78YTMiEfxpCvW+oiIPsIyNe6mfgu5Bkqng1JSIB3d4T19
Z3vDSKqQu2TelxfOmlfVm5WGHZRLEKm0BweGJh8LorM6Dc54+IwJFJQZ6dELqWPU
EStB+cm+FbdtXOwK4cz8g76tase3LIMDRz6o/JBlmBIaBLR8MF9hOHlCAEJgEhNL
71i0lxLv7HKLwfsX2EYbOq3z9X0nqTybTmb7jprb1AxsIbGveMebvLQF026P2xio
RNONHZHphZC7fceEhP/fmg449ayGR51v4Nbq8AF0zUR8tHy47Tpvyouz4zF9L1Lk
SMJ3TdPx3Ga4JlFBsJBpETuDJalhOJYgGSyZOxgzdaO1gUImthO/wmMonSX7Lw05
704LN6Z2PdWkMCg0G523N3UFfJMZT7vC+Uaax6N+5GqyEq99D623fh9J6Gme/xhe
WIAuEOhqSrSHCjF7goG7JgsOL3X9pVGjzfjmV2bcG/Dd3HU+cwtBsYPeoLmQbk4V
TE5T1mhHYil2b6QzcHqnL+LGKR+/f+hEN/i6kdDezxDZCCArkgqa+OFrxU9QL2NU
WONJ9woCugQHWqLnbJW4rk5W+bdzJlyYrI6rYC/fVgsF8wfadu9lkmZKU06uxViY
XNb7S9kqAS9f1GCzXhXCQMt2K1nxuMir2vAJgBezsD8FNSAHPGdG45qutPeRX6Dm
1fU+d7DO9mycIB2a1Og7FySn1kpqAFQF4fx09VA2VeUuTt5nBdd1CJm3/XY5Yen7
+OYE4BNAHs3hYeSv5WsqhOyYvxh5Fb/ZvnW2XMMMpCxpMYUcElXv09KeqWZjP6Ji
wwSCoJ52UDvH0qv5H31dNV57dcbtIIAbbqx8MKcQbJxjN6PFi+Gq5YH4aZ7hH74q
dsjWkE5B+vSsgFQNZ9uVItIGCTqf9HiJii5UwPoAoPM+4loVX5krdKMj8LivNKIA
KyOLb+OjxTmDWEVKTRJ2oFxwMetDnIIjyakASd2e8XwZxSv87iY8NTw/1wyQRMqw
n+KR3V6Zhe1L0Re9oaGGI+gBEDqnmZomjvcUdZXHdyE98rfnEVv+v0siY/TZl5/L
vokrI7+SKxZNk//22hK5C8JfOh0gDZJX5Te/VP6Exc7510fe13R42t8AtOTC7cUW
UVvceudiyGBO40GRCWqOs03t0ebNi23XsC3At3yeQ7LJwcZXm80IX2VaMGeK9Vjc
/5pIGAs/PSBHhX+UTUDbyOy69kinq8Q6SbwrY/F0S6/EY2CNx4AIWTjwt5+K1FlW
IVPeRjMCEibtygBbZWh+mDL/w2XE1JlV3/uervF5zAhlC5q6S+Q+1yRIZnQRax7s
P0RvsLBsDrVk6veU+82w3VFib2kOSzAZkwP86GU9w52JeRT4L/uiwg+CfEfAzwO6
S/7IAw/THJQLB8xJ0reHO+6IcvoEg1IDUn8h4xkdPzEgTgtRxIp34kfzo/wQMQ+3
7ymG2cvO8K4ZQWZBUB7CykXkXFS+7W7mCEzeZRWEmu6dGI8dr1ucHxoSLIbyhClp
fQnJOsQqevZAviWL6VwObr4ZaQL4EZ8/fZnVO8eeLvTvcgX46RvoA2CeZe+yd/qD
F5jgWiuRL994uhNWDAFoY9IufrN4JV9LdjvCqmDF+prCae29QQkdMdW525BgvOPC
7CE0xrQNHiee4l4n9r7b5hpTSQr5N8y21w9oO57MTrq7oa8V2zH3zHc9TCz/vNr/
NjYQJDgKhvBSny747ZhoDtTl3v2uB4fR6CLHSW9wnazXWvKcpUcqFTrjSLb+I4Q8
PKEg/7UnqquGZF7i7N0VCGYJwSMes+zreQWepClNc4u8pM7DJcNMMCsPojqKT6Xd
2Lok2ss7w6dzkdrMQxUpSgzvrS5kDGD3pDF7wmRI/OoZm42vrLknSI9Ix4ZNgVpS
yCIu1Vw5afNUuE5zy585pYbY1pOoRldH+LHoSTFiYxX4AQaC3pHWRnbB18rFZiH7
nqkEqx0bW6ubecL8egtJPmd6JPwc8+/38iCjZ0P0McAAZ1UQeEw3dHhSVQd68utx
djlviAsJasq4UtdCwKVJ7pjrdcF5LdHQS6NpaaO9nWAiKiJqgZuYVCXzuMMKoV2+
Vgo9xe5qYOFBLVXu8Oml7VenqBkwIa2rhCWmBLgHf7FOxNfLQ60quiUGxwuvh4r/
K85iiCbSKF+mMLWj85HQAmPQ9BKmwx2G9oOWRvndVGUQANmg4ks9Sk7C0l8T1/5m
iM7X4xknFa4z5DP9OFQK/sYMgVDugA9kz9K3j5OasGIgIk2twSIhP8p7qP8UjkJB
gl3G2MbuqcCR9RPPKrkCmWCnwLtTh5wf1vfg0FcanD7oSqw3lT5239u6ZMo9UIAF
TodeHPfQQ16N/uxMsT1zcbXqNHwA5LauNi5Fqu+ZzZPZcc0cDIbiuTdfia3U/iIY
FKsEjm5afwte/r1tCwjJ02Ae/yL/KpSFyJQQ6BhBW4HZdg45ZALpPWxIkpbAS6TL
wk9xcK+hRd+rSdub9Us412JCoM7Ge3UsIIztp3JtkqV7iwZ6K4+cy+6bj4QuqYYC
qDJtJswbgPhSVoYarTFjaqDwUpyCZ2ngahDtmkKmj2u0TK0Eb956jgmAbx9pdYw8
+Eg99XFRdPqfiuvuug4sQ8sk4rusaeuVCn6S8M4q27jcaVvrHs3wJlXZaDeCDS59
9gKMnciXMtHRrSZMYwxsP7cYavJUa4z1H7WOSjGjvnnmXXY3q+GXWxU5JRgv3qvB
tgRON7U3URFHQZCwGSC5i0gNE1NxZv2kB/cyJpWdmlxapZRCRlV9fDfjZgEzqOCK
U+l/evWyi15ELYOje72u+2JezZmeztVhOlbr88arAEXbufvP30saNeVa6/EsPWgW
qV+7VrOw9XEqdA26JJd1WPdvqwUgBrba0PhzTq7wyH81m1++ki8lIPr6n3WzgFLV
HnZYsefxqUDy3W7HbFBNCqnkRzQ/yWqREAZsqcjZ3JJv5tvNfebxlH3swOv+4bGu
m7rYjm927zuFCG0fYdukL5W+suxB+pkRNRh8TCp0d2oSxBasgMJBLOJutvzkH6Rq
a1D5v3oBzoSxSk2VYArGrX0a/wDtwDsMXTsl1dFpsZDox1NmYes3hWHcLn/T+O59
k/lGwSSXDdYvb5upUhC0WzELypnZArYf8sN4Pdh7tMl01ggB/XRYysHyxmI5jL2D
J7gNLZJLlW55LdsTBH8jQlMp6jZjyECTxb1UdbBfxYQjj552yRMgwE9Xc3zFt+nA
iM5G4hWW4VD1wxrxei/57cSxc16GLC1TZDR/XO3R//CdOQvD5UvmKusiYetVQjkB
8t8tM+AZUePP8Ixudl/DafdG+LJpO7hmc1du0uhp04jwSrdo9W7D+rHnB3DrQYen
cPcgh34b6p3irqxjhNL9KvFIinO498YWSioT4tQ0EXMY0LmuQPQDZYs/66qf80LK
aDclT3LeruqFzwoxmlxth5dCk+Kejc+3zorYEqPN6QDJclD1Tf8R2wBBbxpgDyv1
ry9UvwO3F7r1vaFgO16A1CpN++EZdD7g8DAXY+R+F3tlNpmf08fiBFXR9k+Xe63p
Lehxej69YSunIzTuLGW40L/ML2QeI0qA/hUx+KS5Fm1yC+HCBaYAzU2U3P5vhziO
mwdGNATMhLTORNuq7hYUliTbNBDkmKmI38eOkOV29b1pjU5tuLGWPrkU8rW7nYhI
WykM9910zZWMvxV3/aS9w03xCnFEgWhmZYwkF3pD36D7y0jOFya4717hfNuLvTz5
VUepWvgyDHD7RUuf8qYZBZFih4WGlodLgobLoj2Ngwf/2SpehNzJchVbdeJXV3sS
QbbFCKDqSMj8Mew5I6SmrtQxosVdCLtKakqI/6lJfk1PKzGpPWUEtA3c6ZzcVi5l
pwH0YR1UjXK8/YDeu56+F4tgrELknt5TGP8oryvVK+fZOE7NVJSjbF2z13AyUV39
E7KNfMVtw+W61JM+pTexRW4PUo9y9xYkN3RJEVj48u6NjhYzhx2pUC+tXEH/flQ5
J2EvPObem+QnCacrOxdUMh63oPhdWB8F9Zk0v21pd9GqfiAumICLVcP1I8wQwXMR
JZgPTj7G3ODgbAaWoq3YF4yOdEm30K2UWFJGMxxYeOXWHMpM7b6hy8fI/s/WguxT
7bFCcctUblzJ8Uy488O8cdFuoRkgqxj86WQWW57sO/pJnYxkQI1XJVS9R6y83+b5
PnVw025q8Dwtj2ZdBKEn1VVfLsRMnOaSVv7462bU0bvcYvsJ+yUuxwwGawJOLuVX
tLJjI4AVo34kjjWI0VFZJ0Gdli+EpnHFy8pF8GCnj+k/iAEkPNH8lVonmLq2TwBi
+E3JrEDR9UbsRn3Edjd9GE+xI3Em0pFsjyQMGgKIJFYF01Ny3EbSeZMhanwYnMea
WCFOoqhAv1b3NROlkKrrH98J3avVo6neJli2LhkJtx4TbogRPZ9u927gUE3gej62
vnuu7VABNDKe7/sC6iOG47KB6KfYPzaVFTHeNmpUOWalvpZAD8EcvwIlHZ4HLDT3
xk+4tMflmqpPg4EPZprAFIuxy3qlntJZg/Zocbe13FuI9iCArjlnRyS0IWb+nhs8
WjfvIpZAuUk958fbuIIQLEq2FkFvs4RE1U1fHGDgC4YcFrHxgxe5jaJLLC5sOiEj
hooWhekojsK0el4eaB749yTm2Ikyq73O+i2haL7QF0JLQaDbdTIig4yJrhx5K9l9
NEAk580nACLt1Y35dx03doqy6F2OYfUTnmyz0+U74qXLvmua3zF+PJXSw34J1ThF
kz7idlUz24PeVOiJPWEAxHeLxvODTmK7w86L9LJCw220z6frex7ZWcdBvUlM3yQK
Yewn8qp1YG6fXPCPBfdo/4pJ9RubQTbLNYgpNPV3hP/yxj066JRsA0Pz6Hi3iubn
1GNuKDW1GBZN3QHhi8ezJR7pKaWZAkqbk0oMD+7yKvVqFvDcT3Lg69yfJRTmfXq1
BOKpqqfzIXz5VHw5f0fEPAnZFhzK31YTn8fcbRbyZeZDVU5wCHzVUrV0kXmc84lc
k/XqRz8UCm96TdcZkHgDXz4762V/Bovxv11sWq7HJZfobadZxsIgTCSOzIsZ3BIO
geJIAWC6dQo8xjw+eBw5MF+aM3H+L8qaAuHOKmWvZZ9aTTSAftuWNgdffejGLq3C
uUm3umtDUqkLF+P94uIGPjBWucfEMMp89ITjAXXyueTIm6M86q33lYMxtSwNPCqt
N0DZtpRYTGA7B7Acuo789kRl8ipe7SJZMoo1EuKuNsRVEu1zJ991Hkenpol918YL
+GsdJ8iTR+9UwYZVUXzBctLlDH+hJjWQFGI7wnbxXlPpwa57RmKSLugtuIgPK6bA
p5zefYUtWLx908IvaD92+rDwQLTYqSxmG+4KxPG0XEcUQtu7PenY8nrmDdwGUutJ
RqDu9Hz9y5/lgXbd2+nlDTcUUE9mQDQsLZ4k4LBdq+OMjD010L4zPSFoKOpF16ge
t/2+nqx0ZDLyjDxav/zAwcsXyCWVuq/x6vWOQbMBa9ExStDYn2vf9WJpqD2I1siZ
B22VqGOCKIG+oUa8R04UNRJdM4KR96rOTulnQN8A8csoWUztbv0fDuNiwgHrAY5E
ooYibRpWMLeBhmYMBXHjEvIsr6vRhoH48bb3qTH9PhiVV4wckTGWcQTJqX69MeRa
0djrY2wMVjHC4evZJZs8TLunbUi0gS+E7kHC/asiKUsbLrIw28/gsgz8BSj8PFri
RPKjve3qyLlFFedbLiad1Vo5tcdpnH/cIx/lY/4z7IAWUccmLpYuN9jfoVacD9eV
qMYBK3vO8aljbPKwYbTVWTxYwoT3n1ItRpAQ0+WfCGDSiR4GbZDe2qF90liWWZsU
FeADLiHt/2Qv+NlDNiUsw7nPM6LMZOC/Ia8Iiy1eCiT8BOTlKz4/kGLTQkbe+q3C
iOKx6aP+7oSBEruwjpaW8oAL8E6GCpGl+uVEpdd5q4aX8lRQw+nPhzkRdWWi9f8R
8Qxr7ERS+qtaEoAXCo1Mkg3g2yovfzu7S03kGyVqXhzkvoNnL9xa1zb80mzsoIc0
aCuW5WnwdD3PpSUhFpPuRuclfgzyMwYIp4wwbpHdtcqBiElqegNMDobAk2Z80o6i
0/AMCLCnurnF0aSapkaUT7/JRHozRtMqhAuj/a7SKsgu8dF114jowuy5/oPA8nwW
U+nnbPAUParc15driwKGqbYQ/kY2XinfE6JR9FrMoX2d/+fQjxfTw9J2Rol+vppn
syjdSqHMt+fL7o9C6ouNM+OuPWMHCpbnAgx5C2VjFG4zREC0TUUkmbIzQ0x4ycyN
CeDhz4eFptjGNOMw2IzLatpqnWD0xt3abUqI/z6x+OkcVDi7Nax/6ge8J9pDmBs3
Xj89INaX5Lldx2dNvMxR2siuNg5LzhY9SzkQarQX0sP5C+nYfdyn98NDF2sLlwBy
ndNaLD7xX0KrLt6uLlZfhh+tpMfMt/2UO6VmRxNX9/QIJjfpj92g4pJWGnU5SuYM
9d6NPOEiIU742Toej7VWsJUOoiLmnIZlgJyNIyduN5vD5PJft+lelJ2rlb0EUBuI
aYMworRR03Zy/9Q/ztTqG74sDyscmlkqY6nsgahRoDzAqckE1rywLVy8dAi9MI2J
z3rkRwl14gQkAw2Yf/T+RNbZhXIvFKo24lAz+KM98+n1fabI4BfWCUfXjbK6nWlf
vwyUB7jnAwSu9gNEnvYZw+w4Jejz3MAPNHvuHI/GiMKlqLFRrDD32vbMOeqSa59F
YsOcyHBRKVcOsTEcEVEItdWlghDNGHe8vyYr9N9VCnZzk2eRUackJBEN0Tt1wRGl
T9KRVPjBLhW7wCksmra7Eat0N3ab4bN+QbNx5yvLGrg5DF0Ug64LbLwXTMmqXBEN
rmE8HZT67O7AApa/6qYpxa3VOdvjnwDwOxDUfPRV/hoLQUZalUvQky7F8aUj8yAm
dq6gUWkYEHYCTVOzkfyaRe51hcfyWN8JIYoNYkDROvuogURllFWEQgFvJQdv9QvF
C92FLCeiAz0cY49+71r38acfZdahASux3/ERrL6YdcSxObhVC9vzqAzn6eM5xWTb
GhyjRlKoSVkZxVN+L+eHb4Ri096dTKeMMUji8gC1y1kYd8r0X31IgqSX3V1SDvej
xcH07ixyNWOapXqMgG5x+CAXG3DEQk4z5T10iq5Nldm206OGLnnBiiHdnqaKtj4p
QZelUhF69J05olQMbnnWPajawwRthzh2tijZSHr5IB/sSbefMFi3lEf+YJVKBLUx
+05cWCDB+8Y/AKNihE4uvYK/jVG7kJyzfYgFy2wOBwq2dtRJf+IJeNMvy/na3BTZ
WBhv4SWgf4IQfmf0NHrZXw0ln95hq03Ra56N32+CGh3i4hTV9ztW7lY1CdvnCEeZ
25h/iOSiif357Dmr26f1dkOkZg3s8rRVrs8ppfD2Anl1O825bs0LR2YV0TgSANNx
h5uDlr+9ezCDhS4HN3eeDATDfHuR0JbJcsGuzBc7yavaH2GrM+fPHZZEQserNi4P
uYMEuX71abmGqkWFGEDZP8U1aHYeFv1LA3vXGnYzXvHXINnd+rddm2pxIW+hApMC
c3FMif6gPDrHgd2E5XL1IdzLZ+5kuQpv6VixOQY0XHbLCM3lK/9fmCQmjNVjY5qf
vHe5b0PwzGwHihhSYpK30f3QwS/tKrxDQz7e4nYq5xsi+zxOZBaJ4IyXY2E7wYe3
MTqJZJWPzt5PcIs/QBd7U6tBP7GwQMCXZL16S63mXwbp+Ma+1hPaA1/naiEJlxN+
RYFYbfAWCGgzPW5prMhrtdsO1aVZ7rf6gla06HZ0nep4wjvlG121z9S0x53jj9tc
PkjvVnY0F6KZplsqS3jPDAGmuD4cHyoZ/mYhQY1h+Jas1RY1uEv/1JpuqpkBYtzc
M1eAzwp8Jvzk34Sd4k6gsdSs5JwFUY9FliOaJTUB/qsU+PU9IqAVEFZCW4KwaZCG
cNodZmZ/WT2o4vOfEhKpTiBsib49SWOjHU5gZ7g8VXS3dE6YV4kprxx0HZxtMxOx
DGkf90TtFzMi7to5nmwLpViwhugt2hBd8g2nHdrgO1Lxb5iVlKxtN2Jmj8B3HSXH
ZHeprrgbKCMEStLRt7IzHxMN5ektWxQj3BYORmTSQR94hMNAGsEuuF+FVZBkVo2X
odolm8iIUq5gf0C9huR29UpIN5BSErs41A6wQdf8TUt3R8kEV8+93xkl3wvemjRA
hnLD3L9+2UwkJmKxMIWClTgd+Zif4TFb3lYmtPwZ2gDS175fQuATid+sZQ62qmwu
ezeFyhGMqtjS4fcLBl/vqSzn4RfAUkrTKV+4ciR+aTHXzHCS7kqL/bf/Bd1Xjhmj
schWrE22oA2lHHJSPO28p7XuFxJNNsLtMmgoqen1p6A40UwrQGuI/oNTOmlkYmRn
QXad31bjyKjnNICb0UW4mTM0cED/mESLW5ddqSXOBLBhEBd0beUKuye87/YswbGo
d9OYrMroSL8Kuqp0qp8+rYu8p1dxFdaHM9X313VkXDaXVaLA8dtwetKf+Sr+JbjS
+F4XS2DlN4ALYhnZBvQ0szPrxOQxEwQWXzfajJx0F1xztlcwGkgSDAmVNbUeII/D
1SRqjGlaxNI6jJ93Q+ub/wWfZtnegzagPXuQx3YH+t+nEF0aFqi7ptf+CLBaTt7g
7QsGocFjAVKJQusNqzcNA/+m5v1uncq2EKZw4OSWzn3zheYbMAtPrLSb5+JvrO8e
SPDML2FqR7zjnmhg5lFiRDAO0wfRNW4V2gBKDY4Y/CWhXvBsMq5CqF8pvs/XE72R
dt8b6SUX+cANve+Mptf7OfRoEJympYKtUSmLMb2QMEzS3N2lKFEUUR7Zy9YJ3ZDa
xfANuHpk4kOBpS8i3THFYdrv4iEcePrjYCby7yUDS7LjcBFVIcAq8Cw8URNvAPVw
FdV2QK+88XR1yYEs81xIUKhO3uxGj4ItIZdWYWGVfJKDD7wuHRVjoetv0lda9Y05
FMy7qQJG6U5jtasoqc6a+wOdgPsNLXosCHXPbNoXsuvuZJ5dBqJYV0WzodNI3Klt
jkHO7Pb2GHESRNu+8W5bSvSlJOABzG8GV4S7qcyGExcjpxT06v5i5cQ4DmNZySVB
6p4ln4hsdNKcbZBVfS4XMF3d+X1y9L6LVDN5Y03LQVSGTVrJdw+7bfyAvfT3tPeC
RRKsA3169/xgF+70uvuPRPjJMyhS4hCUcgj+YdhXscjxB8Zqbbx8JoqiSz7h7a3V
hsUuRRqgr+4Hx5cVk6uNIiWb52APDpyprimCJRMX9ktNVSAFXz/cDhyTyETQFKQ1
iytebW5Tze+yphbNTbVSKtDWRQHwcbq0ltxxJeFQ0Q4SeWgEEoh3JiBjgI6JeLi6
RL6YuCsC4nXK24K2x/MK6S+uPzeyaETXHDiaQq2pPJlEf/jlYg/5Qod+mv+Qldtm
mmX4k7OdOLMDIdawUsAqpAmxBdMjgPs20Ymf2rMwT0uWJ4TmEEqIv4h9mRFdKrO4
SeGcPvSle+RYhUXuNDcbK7GT0sGwq1lmkIMyCo7mBsqoYsh6dmdCu8SQX/V7PN0j
sB6kplpfI+Hx0DHA2kY6F9/aCouGAtaaWJjJYk1frxSerAeMHiNB5xzPOaA2jfAP
J6S/DHQqJ05N4QPreXTK+bH/08Lbr5MEtNUcik7KQZybUhMMKTf57INHruPyYObr
HNo2ujwCUEA9jzeyIjxgnJ2ynj88H3KbglJOV3DcrQ8e4RNL7rbE09eQgL+UdUpQ
67wGciV34a7yZS+1X7L/ukgmSa70Ocd/zzSHNxWSwSjZKVDuQ07cmL4fYBBeLfDT
YO47As+eALE7mg5rIXm8kfOJnFFUbKj8osSIMn1Jp0+CEd7s2RnjLyGCG9JmFPXi
mIMdfMhhAgoLC7y/Dzv+e1PMZby2g76VdLhh0JJJipmIJ0Jx3Fffq+3WDUwl7FHi
bt8RyJiuVUK6f+OEPR7RRkMN86C0353DUL7YRlKb50acpjIf7PMiAayU5mh5Xihv
X73VFSMD5qVjRxXp9M/DBmCt/BPGia4VxhHlc3ykh0ZKSsjYHLkHBANcZEfFW5BG
PP5FA8Ar7j6fAg9HHR/xxIsW1NX+gTlQNkSF/RR+wNl6vT8CebJVUvFoVi/SMTdK
OdFsSOTFIsNJtf/T8oQJOYBvkR3nNSo51hka9xqHZ4Ocn2SvqjRV9iNZzRBcbOO6
/KyBEp1x7snyR7/rMRIZuIpvR0zCITUoMrpcBBHVoXW4o5J0Wi2E+MXIOCGhayla
TjVyLyMpa9GIFU2Y4f8Ls02qOclb9SHuROHDcNRFM+KIAYTY+ZJ+i87C0bHX8+aM
n99Ka57KPuvZ+zulYUi4Yk6F/WObHI/RVhEVtDowLCMmtfnujdJr3aKd8/kciHPl
0+4fX/Kc7iUnyorxG4aoNoWJlfQZXzPTyNc9zka/JivJAM2uJ8uurJZHSkLK9jPc
DY48dUTPu+9YJStTdrHNFoMAx1sHfJG56dHZQ4anAnCTNiJSGf7FcncfHIgShcjl
ktie52OBBddUE7lOEwl3aemg5apFROqgeDgUANHusqv3zzceEAsup9MjFdz8o6V4
NPfv/gdkv6bbVK9yCwiw3iAoUScAdsR1uwwfeiRDTJOUTNY2WZYCaFTELBS8LZSW
ACSVIgLvEZR6lnG0iY+CYotd0cV7ZN0ngtk/5puNyxX1yuZGaw1Gdsw+95wCelcg
lU4bFUEvN36WS2njMn8drmqjZVzyRA6Fgu6SJDqFEA+guBA6caZvffia7gQEeh04
etSFmrJQIb4ICL+FRD0vgGqwfJk3pk3K5VDYIkJjyC2oAUsLif/Tzn0GfKNFXqPG
5TR0zmcYzqAj0DW3b3DY0u07KoEntM42RPWa5jzdMkxQMsw8mupqBh45yMavCi3J
yI6H4cXy1qsrOOZMKMyKz4Nhd24+P62YZFYCdSOTWMy+ssjENHir4fSXVXOxYtoG
MoPYeZGEDxlZCw3VuB6WZACtSK1ryoVAFxD7/9WlniBoqntgfGxXZGHedMlTveai
3OVIHcMgArBEjov0dB8f2eNtXZDXilFaNkDYkc243YYkZeWrO6eZF1ZvZ1yO6PGi
aLB+kcw9aYqkUS55aOKJmyajMjVK+sQ+UyxTEBrB2cxzI3VWrOn/bYg5aG0iq6lX
mqSUh7hRtsupEf4HFRMbd3Agyqzy5914Lri0UsV87p6R43hY9Qthn+yaBDOAg4u/
TAmGm9jxT3YQLJl0hVxsVSeWpNJwFGR/kn/KNLCSJSP6bKEA8bY2RuCsOuY6o9Sc
ECjikhECcZrgry1TY8i7MAaMh10peYpCopfnNw937iAWKN54N5NF5S+U2noYwNp/
Ia/h0RWFJCsuvJcJy7eQDD0uQUHoB1U+XjtWJKAtAIXYA2ySQGowZGh6DqNl38Fj
IIInfMXWuW/eLkU092ViZN/XJ1GltklB62VkYgDQA9eHOEh8GkboXCBcwYRQwD9s
o1VJWHzxXB7B9FKCUMpB/FpKKiYcEFVp+YplEDrVAFwQEg5l74UtITABcLqcioar
GUtjZCu6t7N/BjS9/dPXPO/kbZrDdqIzQYWnxIVXC/yqRX0hQ3/I8VbxARGfPKYg
XVKIZGMfWhXXFyVBCzX38xCRm9nEKsOrG6rZp72WEI2JhdTBDsItorYHgZHhb2a7
+FO96dLtjPO/1NxdzOukNFe+EhIrDXpX1ssEUCJYx7t+IdPhhvB7+OZJgxU2Ld6L
TzARd3P/wDvfFSAUQtFwPwCn6D/15q49US1CgvD6qJwaAj6lZy1flB76FxiDrfkX
kroOk5q/B5pMCy4ouZdiE0EXbXBBbANV1kRqP5ZPz3I1ktLSPMTHG0YZkHpHfQMx
4w9NwWWhwUNIEMVzg7XwiZJCNOwDAmG5f6qLtDIslQV2Jl/Rx3ArM49Cz4svjCWB
Cnje/YBcvTTEefwy+dg+Rgsi+blNnKR/snKt7Pqykz7jnRt806yc7WdqZXy4JC3l
5Ldz9YAbzWyZX9FCf3J92Q+HIy7cY2Z1JKxvb/TR+OtMVXjl19BnE9+DPWtIE8Nl
6VugXXopUePYHF8fuXmV7gv05c4mD65Tm5SC/ylMCWrzsi5edXMHzfjtktdrFxM0
BFWEGOP9MviVFXwLXmCJ/4ZUdPaREOofDH99qrIKTDNxZtPER722eDgJndjLpEdX
yN2MXboLOmv01mJ8PCURr+pLe2rFgHUTkuDZ7/MoR4gwLTJOSqPToMfI7ATLrBfQ
S/qJNN2Z1yCTqkhiIKHxESI2xPsqaBQOLIcKu2J9Wk+n3wW7K6X2+tFuK2ZbjRVN
L5uLN8oaN7eTVLu8qGZ5s5XLN/SzHkutofu7H59QdFcBVrp3zXxGY7QWKA5nR8FC
O/Pk+i7bVJrXon0n9S1cNpkVAL9uzJ67DU8Z/fTJOkzriQ1voe102tKQ1DKxv2UM
C3wTg14bmOgQIRYCmvnwbfuguc5vmRl2jWxLkzR89nt/8bh+M0LxdlwAk1/Vj6jb
sOqA0Xdrk8KhCnr3PLjfKKeRs4SNSSzfi5/o5BBYQgWUyk5YrzyRP4xR8pT+4HNW
GEOT23iEAg8zQNKItUc4+GQA+A/p9kpH3QyNihAYwOO7IdpPVPdI5suTldgeA4BH
tlrF2QuL85hGUu2JOFd5q0THm0vDo8W5Ef02/dhRv/Eo4JENvm8nCzJ1y9I7FpgS
RfiY0wydRXGsZ+R2B838KRNPgnrXiEjNGPFQI6HImZCx2y7ArpKqanUSwXJEm8uM
rbiBPcp0X7MSKc8kgQYoNC75GimrCD1y71tooJe1vNEu+0LstQrRDerDmQlMnqlq
ZbZ7QF9t68A9TyqePwrHC9It9Av7Wh+0OqcGaWJXZgAFIgc7DYZI0wxnQ5QLjG8D
zeIhEtEa474eEMAmkX/cIxZkT6rHFHqedoMf9lIzxUBM0hr3wqtAC8wE2qJ8Yf70
rRsHYVRV8huKCEeXM9kX0tWbp7VxjZHixsFFm9NryxOwJwbs0E1HoPonEO8v8+N0
ZQVAIPeBa/x8xv9Fm6RIJcofP9pRvc3ifwVXN6WKjAgqYFh4k8Baww7K1rkBd6gt
ygGHxssfRRh0e8Zc/TCcxQ0n86N85xwIHGdfBOqa5SGwYtBazQaKT50YN74GaGMl
CSQzx7rZEMf1E/Jz3eLTndJIagSBPmShRFXTVDRqW1LolVNml5cvZ9fI6lIF/j0Q
CYecLtEmwYNOnibSZxVsJOtV51lv/EWrF8/LGkqvEILXQKuT8d9OM1IjDeW/uVRg
toNIu5+2MLuApUFQgc0A27jCJ7q3TDC3ss/EYDLayjWgJtKzzJI0uju1lTqU9f55
gsOG6dEIKmBcmd5BMbVpBEsnEHCL4ugiYi9XcH0oog2l/6NvcRIU8KGxPBhGx6Km
QT1VjWJl4azFlop8OWyQq/WrrFePWtK7JkHJLqrxrKwC7n5uU22mkTvQthwReHuI
Aer72CHUT5ZPcz1vF18tDm3kLIOwfSZ1Jj4loHDHgBUBId5FxJnY1rR3I0Tq3/4Y
rNUuIUiI8yfmBPjfeOGyOlm3vK4xB/mw2PtSvee2VJLPvl2793Sk3TwKjOt5e0Rn
nlI2Ep4goMGXuzMxpsgkyw1HLj9rK4TbdKoLgvP+1XkShwntepIlaFdgiZ5CoSsh
P/p9fQuOamLeTmoTmiXKbS0TrHbakX7MxNsXhvuR228gqV4qM26Mi7k5+XpFuYSN
gkWOBx3LH81f72CWD35Tv+BiPCVH37v4r7bFHN5OeSkXiWdI5w2rgUJs9rMfiwWF
9h5//R/j6BuzBRE01XgGwBkZkjTpc2KrRROVuY4CebTXOZgPoqtwUK08JN+rjFnz
bnbPVHVF/2hwGTRJcSdREJoqWifEA8iwjcfRDSC1DCK3Z1IFm552VgDtw7imgrGV
TWBQAQY7bJH31cy48PTuuW1UBStR4IlgAC0/qlFSxD+0T/qntSQMc+Xtm+D7op8W
69+Y9+FslSsO/VQ2Ve2jgX3NjBpI/lY8Q/D8k5kxLQBay2Nh5RNExmyMOl2q4cs7
HhcE5IzpmoNvisHeE+KX2wPTX+aD9+UX9/vhBaIcpDGggsqa2aDudIE4r4rBWJtx
FDydbFeyldhvjX3jOHwsl7EbahzY/mQyWFT8iTLMv42fuJ5kODDb+P+jfea4yn2x
BNTLp4LdoAPZIRdCJJtNJQxQseVEauLTtQr0YKNYiObcSFN9b9GNhpwVgVwzAqTZ
KpCn7JDBIdK9dMjlPV8Xe6yna4taJaOLf47lQEvenvqPHZz5YW7VkAWsUnpxAIzG
wPB2JN/9FEFMJtL7yxbYUU4svdSdmnUFDSeYChQmdYtGr8l+BVJn8GpNTPg842JF
Wdhtyb455GAsfA/od3MQyAqX7djXaDk69kLWARKh//Ne+KqmpOB/UBe0ZTtymX9j
u2LC0uzjn8Y0+rOxHG+hn6bNToZebsXERWDiwS3Vw0CjDu4JCOSy1NRPz2VvdpTE
5EL5vuNbr9jGxnHnf1f/9yC7umc2I5F5XC0usOzjTGu8HElffftwLfwn0Rh5bCpk
xMNS+M6pN2Bxg1FRO8YX6qAgwgwIjAZHKDhS5g79Jh7h1iMVrYnN8HsPRHWlkyOE
56PytR3Q/C2iqn5Xar6adLkg1Hk9qG7Arg1T3act8mk0JYkAsJTfGGWXPBdulG1J
PT/3daTZPr7G+mOEMly4CggMUI3fAVP6IzPuzw2LNYMlPGUdS9E0Rf6iziiFtC56
IE7eB3XO0uQSFA5gbmTQtXtHQhfgWHb75dbUM1BeyNBbzgJLMGNf4IZj1t8zwdk7
rBan4hAC4An6OtZfKgcYvzve+nlV/QLtIoSzMWTJk3NyfAGrLG+yVIhpLi7QhpTo
zWN8EEGBt+bpSox38o5056iDCOjTa1VUp1+70IHd/KdgSIhEKY+EM/JEY9h4GN/z
w7eICYW2PdZUh4kAYKX4Y7Df5wtjFeSwXj6h7Ac5XgfAn6TKiR2fL2I1c8UBnFo5
ADSSMicPGNrwpJANmTR9tCDVPr2gWjz44aJkomPAThB/u7NXmITB8+/jHpgS1uUK
/7IBkc+iz4E3ujKCdBE5gYWR/Hwm00mtE+saMkp6Aqg/Hznjm/2warZqtmHmp2+0
M0xZDCRNkBeSnktWT3jbP2UdccuTtU2TzP/CZsLS5oEi1p4LSymyXTCDKjZ2d+4x
Mo4SHGUgyGkY4IC9WJnqafoHKzNNVnDxR/s7B0dpHn3DNAO3+MHAiCYV4+UsUDiA
sidTpDr+IxixVIGzF5qmZuX5yKAtbMr3rEFZggcAGSBm/HrBmom/Y00Px0eWw/wa
itzn/HIG7C+za5Ueu8QW5vxxoPIdFby5kKIOSlo/ezUh1PDB2IrFSDwA3KBpJ8UV
6zI3lTZT2A6UWuEtI5R9GXoDq3X0bYOe8qqSom0q6VsZlEHOpAO7R+bWCt8ptAdE
T+3lxxN/DfvShEaCFC8SYlackBXwoypu7fVRiaoGmWz3KCmCJmU5MaTYUkZe79xT
d/b4q29qJ6AmyrnIEhrP+7fdT9Ns0+Bk++UQ/Ye/MqKrrrAEkIqJUsoQkI2tRV5I
h3vI0UMd7u24ECfG33/pKCf1DyVPdutd38X76rx65fox0YG9vpG2dP/JcwF7BKIE
54cunuNWEP4bAy9SfSuLzBkAh7QSrXWenQQwmnmfM5GLY5kpH10Eqy/hqiUhI2C6
B9DC5JgaEsISZdS/qMuFvUEiOIo3BbMlp3NmM1HY6sn3jQIUqWfHA2njWkac9hQZ
v2z9XRNUmfdMzv/BbGCiX2VOoXyYMan4wyvie4c6mfKYW2lF1eNMstcEmuPaMha8
wKA1g5zaQSfwUSoxWb9zy1A9XJwi820+U91r0pOlcAI0H+nlpF8coZeuJU2zevYx
SaKj57vxg9h0jxdSh777IZ/gQLulj5WjKYNWCwP5ikMzunAK9Guq3EkTG/DEApQs
P8UnVlukS9uMW17S4gWUJPR6iPeyc/WhB2kgVBxDntK3l9K9JhbdRLdZHg9oKK/W
tux0tadxuh3o+PH2MEgIa2MOdPE8IpMK6e9CtNz2obXTLi6+2iS/ytoJ21Dj9cWU
Y0nOpevHbZtGY0kBVmwydpXcvCEoTnU3HVJSEj8jies93AEwRdnDBtFSXmhXSkCK
MS9rwZHk9zU/Vvd8QQgdL/qYCnmquWhB/6wIThf151EuamyDy8WRQQvDgNCvp5Vu
UzEY2pSsFOgop7BhD7lkmgUOfnbXFbbS1MgZ6VVzWuXhxI2uZHCp28v4rlFbRFyp
BfQLpgCNH6gNcrQrPAmyr8Akx7/YevaiirMj+kB2VbdGBP8RfcaNBnYOV/8daL/q
ZFBDKcYXGJxFjn+Zd/AZ/A+UBplk48uM0nkwgdEhVT+LSwDDY5DsQ1i7Cu9SWlbz
5eu9efYsvvyJV79tPFn7MVRPfob3qSeoKMVQUfN8QPGQ4eXu52pVDjf/O3XdTf6I
0+gOGKBXZZJDwhAlKZp1t01Ht72fKpPPOh1ARTCg9jhHMK04brYc1lPOyWzhV4KV
veU7CH5D803pV2sl7cMCI7PQXUt04wdL+QPvArQ7ZJ30v/zBSquVdd987zRv89Jf
IvcQmuw6GJKnb/SRIeZ3yhxqWrPdXNhtMsxYVW2xoWKdYxcpv9tBKt/vGrEUDGf+
ThEXITrju0tJgONHqqplAXZNeIuT2g8aN2z2CH57e1b1DTb6NA6yYXpedsR9ZzhG
iNbv41jKEHuV0uUcuBtYxK11ibDEI3rjs+MaUNON3lX+zNk9K9Vw3PE58vrh+xz6
L8Qs0D+EusnKi+aZv7dFMArgbJ3aUjpsX4eJVnr+EC0AUKneUjb/SthT+ZCaqdZs
6C33J1lJU/t0GkT5NigreUSE4q2uHHP3NlaWsh9RkKpLemktYkqYF8+U+7jIg+uD
Sa0c8bsfDgj0A6Wu2sbd2eYpjoPGqCZ1MQL/t9P1cmuM4cIdOawXDkDzggLDEiC+
4XACVgjOvKczn8oxgYX06fIp8aLeZREUGPz2OU/0kwqxFuZVur4ojPmT/6xHda5N
LWN2oWRvRguJZhY19PKhh/oXOUCfqO9/CRxrWjqjKuqxoqZAOwsSjUYmmQxvLwTH
1GesihwwwtDQ7gxFwnqHdTOQkcg+JMvbjyCbGvLStuKYVEBJmxlBl6HQ33uMKsUc
MQPy+vuIQvB380yJldNNtRFwe1nA7mwM7V6R5P95aJqVV+WeWcXglsPxCpj7sS9C
a1fuBRHQ1qZShucr4LrgCWWRyQAbXVcNPY2FluG27EXJmjA3Zvr5j2rH+MWNXQ2K
EUwx+mauY5oqYgjECR1R8OIVe/7JqCYtmf3pnUjp7tz+FdLyCyXTR886GTs4DG9o
dI6ktXb5S+6oxCTOfIE1AJKsOuefljUwyCQ1hmH7RXbTW0P1GHcUAtp1WgnMqOjL
j0C0A7h9Z6Yxixt/pF0FpzTKRqUZb8avQhNosxqutRUinIVmj5ZJub9ud+dCK7jL
XG0ZAozlvlpKY0N0hy8a0F/5ycrVzWWHwdc+3TbQYHhdewOuu4xWhjA+yDtV+Um9
1MwEcH5vwB6/x11CbNIldwzAO4ZQFZcUZWasam1U10DO8Sw27h+p+sgopIiBcMpQ
hk3PA0kmDXjcZCFtsYbjRX1/YciEswZzbSGHg/QUAmOPCAdxgDIsahnWE22sH6gg
PwSd1jbhDfEdr+mauR6tGagvDbD11mYK5/2l81dhoc4x/wMiu/OheTn/5S2CLSI5
JtoECCMp4yLL9zewGFIx9NVCHgT6iAdKGR6J2ek0YyBnAQVjfAuUidZpg8r1RHXy
SuCtC5yfzBmfhkicrrFdkcCie70HsWPKH7ikiAS8RlILohAuRdGCaGNIgXMox+IP
PqvlNvWElcW2cfTRJhL95vFW8XFg2D3GDqq76vLpoUiL/RZmXuGT4twFQZAM62pf
hxn17T8EJNEGg0Y9Lckln5PGDrha+hg9MsSBGgyu0gBxe+oom1U8kL5209yuIwWB
d1LAxh/7F4QNNnfRCTaWSn5JYqyVBWFtWPSYaoxaw4KwkCQgMFEVmR95rruYiMl6
WsuWwj0njBn/A52iZLAyC8gHW6Tb17dMtpHRvToyFl4gOuzizUOsj3GIH5wGp+D2
D94DOM5KYE4bDX77QBuR2tfGAzq6m4OKXv5W1mMjmef3ul28egs+kRELxuS8ED/T
HtkKSi05E/TpJH93BcIxUIDqXUTJHTBrEYdQhUUwmHJvV8qTUUAaanCUkkMAaWIy
iJ6AlcMjAy4sS9G7RwowDDKckMp2gpEF8UhLoL1Olfv06stbGz4fLOr1fXT7dDQg
Hu7hQAsknvt/Ve8QA4WJC4lxpQoKbg0pGh13xHxVVoICcJWZBidPzyve+O9Ko/an
2tOAK7UGp8G+5VSRR1ULcyJnPXDLYyDK3s9oKd38TT9jJh2tbH/XPNEstZgAog63
WlQpUNosNaPw8phmM0cKVM670wLVmtUhAA+ijrWVlQLYH+LoxCumOIAhkJQkQIXP
lQ6bgAO1JxVCyW9VmleUPA4Jk3gnDwTlNDUjQyA4WEq2REiPgEdn+XfCFgkLiomG
gVDCyG5lu4tdqGYUYoFapRPExWD55Bc4ecvnDwWB8R+RFIIzt9zpizbLuG3T/r05
NSj4cBqPXxcy5lhIkLrA8dy7DhoaiX1W/hdT1RsbU1+nfee126kuZtIva2SG7tXC
vfSTur9TutKU6MXmCq8XlU3Y+vXJ2XexAAHnBFmlViUsTO5yOSLoZ8g6I0zKhgvu
zSoTrc6xjlo/KvOTVpoDmGtlS21u11s7MDsckYRDt6zlOqj/whWlFym+TzyzTzCD
h54sWdgVdx3YD3tj3dDlPiJIduqTq20kgcX/mjRHiIyd/uH/0rsLhvlo6WsZKl4E
RxbUfZwvelCtDkUB0pCU9U7+3ZxFR8NfYTeA7VYy9K1qVc+EuFfb+ifuGNAHZJ/j
u8z3/y+/crBsmU/Wpvhcs6TdQTOIcQJiu9AvOcvnYE+l+tG1LHFJeMuvWh5uuUzt
2xQZ9FExynwcLJu2dZAExM6QIQT2Vev2mDMeddN9027W5XYYg/SZ1UPfxh3XyOc3
pK1s3LJx2CJNZoC9m1vMwqq7VlTHXH6LdPqmQjivCdxVLRxCpi4mDPWqeM+0Lx91
+/T0rQxb0nzu3QzSihjMDZgOx27zFAKJf7cAI2lhJL5lZ22luM45HEcTf9GHewP3
EnMV2D/RJ0+qjqeZDuc2nqfvAquVx+WswFBove+NaCWLrrgl+IkVvyKDVfISIl46
MblJ11XZSqhH8uv+gSJs5/qaBPLnEfAhIepzYdZEPQA/CX11C4mu/8y3hCB8dWIW
xFXbW+g6NAok5GDmEjS3qPKy603VBN3+Mts4VRtdZjue6waj0ttsa36ATfUxLzTM
a82az+CERY8tmz2/f2d18aEJ0rCWqqMmoIT5ZusrWq7yMBmcmD+C/KmxZHt1w2sM
77S8SXq66utSElzZwLg6+iqji23IMXdvXFVJwRK7epfXiOTSII4DPmFABRXE8uYm
Wr3i1nQj+KnMa3T0EHXpw4oAUsaJg8Sp1EFbShAwU5CY8qrjwUslY5POLnqvZ+aJ
6eVR+dkLim7jfUAB9OQD4vPZgbvriuv6xIa4a3PITAZC+pkackmai+nYg+4Zy+dB
odwvA/2mvjzCYY2ZY8DSbhLtMHSnSD1kM3ttdc6C2XTSOrYnbeUGzH8+4gxzZciA
Pw12139G5NsSIN8lLKTdkn0Ng65dtxva361k0M6c2VOnSIbkvDToVgbOS4mPt2sR
HjgiTh6gYimBmt/BzJCCEPZgr+lmpTOBBVROMgAkTOUenvVY/P7Ph6YaGP1pVMn+
T6rzYmsTIJ3zE2Bn/jnZ5Phw+ljOBU8wl5oGGAi+dklwh3+EO9LYsZWyKz/Qm9iS
PNkGhG8+GPLq8UCmrvmv6Z4mE/4Nkq9M9VKyziDey39496kqPYwyP16kXVq4IsyF
RTTpkp4i3OJNWxthPeEhY4WGycb+TtW/VflRkuG0OiJ6zKcZalhVfUY/bRXwLbwQ
foCsuuYZY9/rrNl1CpAGr0v58X0ErbKZNrXM/S5e3rbd0i/4q6CuBn8nM3mzxREU
adOtTL4bLjUZ6GKoI+XmBR+GpK4j+FW0zCA7z4zLxy4FehjCzIYgnH/TO7r1pmXQ
/nYzFyuBjxnuxap4S2tp9ugWpS2S2vUa2olDmxEKZqC70iyWBgMFYKMoUh57pk5K
u4Oo4+QGSVBJ7dEy64QgZnBY1K2vsq5FLN/i8/tH0QtDn7CAgGytpG4OPWnlKDED
73DEHICp0ikEc/1BsW3v5/L4R9r4aK24+ANpU9BpRHs14GEN7k+J7UHbRDPrjb3y
g4rQc3R/Z6sNNLF0HoirZFu4XHSsE7TtGWXT5x0uZ0P9d2SX6NxAvuI8rd/Zb/Cq
tg2ho3VpkusV7huNu8NMI0Y5NA5Ozpz9rvb8QqKwkS06qQbb1Sh2OCyF/IBXraBw
/U1cNT5CzpPzEpB8a+Hjxn4fYqyMziiLHgDRuGmsUfEchDxczSSP9tUuJqvP5vcf
2MrZdSVzlm3klnX9WiGWWgeTaES2kCOlSbgvPCEi9BypqmFi/QfcwtYl5m/Dq0+r
J2+m1AhnnLa9Pke4uoKHwrAZ6jyOeRwMA5U4F6QTOo5el99mb0R4yGoI2bSDIRpM
JxbaCVznW9W69hBFePo3P2dlQpKmEiFDBUmPIHkKFlzmYxbZJglke82ECLczpNtQ
HuuLo+CXgDYq71N4HuUkBgThYQTlyj4WqtsgUjjdpSM3qWDjAvlC13wrLpCliKt/
whux5YFL9Mf+o22VlFR+w59D5ONl4rDsHUshT2YXcew1bN7R4T+UIY5UJSZuOInb
TfCih7Lxf9vYv77qLYcccB8bAVtP9CyoBQ3ZC59k13MrqWo22mITP3fbo9jnvQ8c
Xr7mR5eQRsjgIVf1e0p0Se+fJwEP2ZyGxfcHNz6x/qTxEuqFtzkw4vldrcP/yX7p
iSU/czGO5TzbhGj0sGaRWtY+tfageTlr/+TBzY8G4t5ZMLGGj9orZp5eF1BYf7MS
SftbrBS86MbyO/vGPLtucMQ/B5WdN2bT8jxrQ4xQWVmCP4zlAS9GDJr0HY2krgl+
rPn7ju78VumUALkJQGCU/x1fvMGjPbsqivo/5I0b9SSGjzgznlBWYudWMqO8qmqE
jQq5rgl6kbzn05ksRH7B5RSB3iR9kPKb7GnQs+rkR1KBem751OUOJgGvkUe/Tcor
HlANplNIA83qI/v1YEyVq2adJ55l42WUQiv7ydxmXLmTzq6e7L1+gets/9nYQwpr
USrd57nVu4qBQjeut0OlwGMqMBocR3Pqlu4BqX+b7hcQRtpNnu/4p6LBYvEPRjc4
mrCHVKdoonwHu1X2uKLczRgBsC87lgNScpLsdvxoKULk+q3fmLqCkut78Pmt+1S6
qQnWfo5/ngl51CpjC5lTi+Lo5lyf5AHjkvlnSWYCVDLX/AIx2mTqY0NLOLwFEw2U
1aUj8l32dmpvKQQapSDwbCgIehnmwNylD8042nnjQ4BAgA9lVmBW35VC14F5vBJS
bFLYLR/Pxh6FeKUDNIn05eDAHytDGMgdT7qLDp0j/MNKfOgBfiFIwj0gPHqul4Sg
4Ekb4aSTFeny/NHEP/YmmUIlYPJfZbGI90tjwuE8x4781gB9qylwlYvBm9UdsmUf
ZNItUJ5519zYEOGpX5iKQvtCUV0mHaHqDHPZ6uV9YdV69XVd8X33xvMXevbTfLGW
Xc8cjQG/AYIIKVS3xhfZGUFcm+WI2plz2WyCVROxKGsvvG0/txr+/Cp+ISyoOl+0
RnBp7w+qyeKcGkr9WHIqvEtzpFzhlSIXOXyIiBrHrOoJlEbIn0a9GpuRLxT0I5LI
043ut4gYaeNeVjFLx8+cY4EwAoM9xMwnORJOTuOW1EeUpE14oihNIHEN554GQhQ5
wSTIyC/V7d7qolqR1YkWE29JTzSZAHIAOO9xzzTrE66VM/b8lekDfA9jJLS/D9I5
fePkGbUcYN4tc3VH+kUGq7h/FuexcpHLoZRYAodjHiYDIqXkyXVl8v3Kn7+6Zcke
4RswwtFWj5YlTJeUW7sBwPoZpttpNP/+sg+hiutLD9bxRqPQ5AX8fBiH2E52a2xQ
sY86RblkfsUBHiSXE8aN8b+yq+2vclgGwk4uL4y8cM/5VoCYGkwi/BLdB1WtbtUv
YuSUSZZzTa+MhoLpODtoTwhmeJUNotk3Ghr1fa2uQ2W1SXvb87jthKAAmWKq0rES
6NgpKd+EMzAe9yE6XcG2Y6BT2PoOneNIt/kyNY2CiOaw33FbYSa/rEzN/sQnmvgO
iPDKCG5Y39uNXsmzHu/LqnaP2dC/SqfWPpII154Z+19zddWp5bW8pwDJ9mBRpNyu
X73xd4Mg+vXx/YM3aC/8/qkNgExjOQTT4qo2wuI7BcgFG8I8VBwAF9/8pVsmNO+f
V80KHYjgFBcXaBZGtow6qtWSUdBsT4hWQrLe+UT+U6n2Rg7X/t2vUC0AguSnaUua
nYMVk3QR4ZKgZfWlwiPWPWCLPzYocZlYrImgaodEKxtRbGKesDcvK2ioQDEf/17n
ryndVQUouwJeq5bUDOlGcdZKLMAsIVHaeQ47yG13Vf+EN7/da3jNVRreVmC3dVhD
dSo9LpP/rkd81JTTfHVfQnjWPX0ImYNUVBJnL0QWQbph61fNHhm+5N5s8H1Jwd+Y
CpHxXYoHaGgm6DZmbrlj473QIpdrrp0QnJfz7ncFvIoTpAi1fSWVlpU0+W7UjRua
beerNmx8xNqKXE7bRKySWUl0Kkfyw130pbXukfI75eH2rTIalNJXNfYO7Tfn4QCP
j0OQrb9BL2O47ishcf/GprWNpRo9jZ6r/t53ZSK22vbPO7dGhYdNQPVs31AKwMSz
H40JtLAxdVpd3BDmrqvF5N70Yjyy6+pZjvYDo+byiAmy+bOy8ysQzwW6aU4SpZlD
g/cWIt7DWV5gZriJ/xvPd8baBDYOCUM2TuWBOmsCzOf4ZGjkBoHn3Z/BTlFlUv0U
rdjqXm0pa6KLfrc6nj1P+eULZc1nBFmJlchAWg16+aJ6191Gf4tf/CEPOhCUtvF3
4a+6WxqdHcq6qdxusM0Ki63ivqjNYC+QEPlXybPnyv1vF+BSavHT9eW+wysqRzKg
7VtBvhRoaXccTt4sumujofYggbMKKzCvVVpH4bENZs4GHVDY0VMwFDe1BpFfEcVP
On+zMGxCBMo+ZGfSrJcwQnzb76m9UiaWl7eNTRwlKV/D++vI0+fM40BXo6zmjD0/
rTWrMfcOxlMBxMtVdrijcQMAShsvyXx3YUjamLbTOMhuwy7Bk5tKAR8i6sLGC0y3
2cpZkuvqAb9SeYJ0W046Oy7ZNEA7RPqZQK8aitoJQPG9FMXIVi9spiCCL47KoQ9B
6TM7KysuWp+2Cxmnyv7zyU3b1yGmgcF6BdeY2PA+BkkJ1dX77A+Wf8V2IkOqVthN
c2o2C+seLlA7cEWJAxh5GP1ZdqGQQaTB68ArEDFeZHCf4qTLa5u3MlLm7ySigWjU
vL8gK9/RasQD97p+mOfcyLuIK4GLurUniPMlmKzQEyJ57DaO6nckRrd0HNOB+NB8
S1khljLRyfUbTAPqO//sd2NpjsR54S1O1kYNocVRn7Gfof0b1r5VdYCDBLexjzuH
e9QCorESav4Ri4tvCfHDH9zFehoyKTKpuxDgbOl6r8Cxh8a89stRyZfdohhxS38e
5PjWa2KZLuP+WmzdjrUKHRtKPf0TSymLQbU5d777T/VbHgNTxMe/HIfA3MGRTg/W
8QyGswR7gIqi2uQjg2I2pSGfSCaK1BCgenflExBNOCTMaLQfnvsLD9ScFcj01jHg
U8/NGC8H6RzMAOLwHIwY/Ld7oxewRYMiXzSpFtiMKi7Ye2jDTfZpGlV2+23Qyz4Y
uxbCCAK2Zl0b4935n9RYOzIEHK7Jq7Px0rSaydmpCa17wNAgqSNyDlaf08KDPaur
8uwFTIFTznUvQ7GHR/wGV57y1/cxhOV/gpQ/QQ3kt9cSGcGewby9A0kLP9yfn5Bk
s5BQtlkgF0I8q/Mcfsk9Zc8lIeKwen1seAi3xuczBHipKhyeWwPzq0sGDrluxB7O
I/HIZVkNPbB1aXuls75SH8aaM9bW3NB9WlZqdiLoD3qS5Ia31x2i41DZhWUcxKTE
c5im8cwFWi57sBTTcywzBWWQhXoDuGMBDn+o6MB3sMRuKWk3prZhzUC6mPfvNIwG
uAuQvnRgbFjKj6FSDAKbfeiIpUSVIrb7Ss4zYZf5R3d23Cpp0xJ4ABodP2zv6J4k
M1HxkIRwDR7oq+3gzH+ZjBnbtFfIAHVHHWySy5moWjZJvMQjsI77dD0SR1kL8nAF
slhKmZ2VFrdzjv+iz/v5em319R+HpbZReqPItQlnb9xXwmLOF8Jbhz5OYMyjffV3
xJ+iXuNL+ia8wCGHio5OaMngUdIChFzgXxQAHBkeS0Ni5cKoQ4nRURPnJIgOyGV2
yx9IIf12PX57lplSz2HWkPaDvoNsOErmoZfpiz3zjAW6nn7raSFr+G40muzRt3yy
c8BPssZYm5Y93ldVXnXJo7v73sFMLH5r+zF9d3FlCHiR1dEkfVhVvPUdPT9rmY+t
uZwZ6Zb/sKBiFfQVA8ALneg0p92rhkvXSI7DdgqxsxeGakopRYK+RQ+sDiDQh1rF
QE+F53h8qKRao/VqoHC/MhfGCk2SIA5grTOD6x/EXCmIJKd3raWFP+1cfVzOE6l1
pD1TnRAw0fkmewZfmOh900D7LBzn4iPmd23OVDnIhtpId1gkYyQVHVMrJxmvkkHW
viZ+boNUi4SANAEkvT/ccOVv8PWqSsRsd39y29qmGlIYH+18CfncpW5o+mAY1Faq
rxNFmUcMr/7igWTvLZoBlD4bdlLA+Az4ZmgzA6XOIxVx5Ran5WqW76+vaAdC/YeP
0Ct4fKZVOFrdpZeEcWBwQWVS2fiOh8EmigODTT7peeMWRNUMEndpt7t9es9iLqAF
2b6x4H2qC5iRlArhMqwWCxXzRbgKSEpXtc3vpPS8g1ftRuueWL1fdNupCvflACFZ
JeMiA/jD4owOZRX9eC/jj8PtBF52ePZAbxLorbQY8wwcMFKJtjhRTbsf4PdFRpwu
wEjVtJXjC1LEw6Od5+D+/aU3/OA2ejfPtv48GYcK0IfitwgJt8uhW+Ve8yNjhsa4
SmxaIH+Y2Ra6sFX/e2+tImnH0XEujSDkVhdvnYRnswsHVAlct0tUj8Av0tCSxIEs
lchhbaFDs9g3qKrku9ZAyHruNc+Zq2VNSwAJYFkt6u0fgPBMWJX0QWlk+gSlnGPE
+ikg3ov8GTKspryfaAVEt5aJPprX8aIwbcYbh5o4NwXAsLKOmnFbVomr4bWKfRVW
7+Xw0HxNQPj6jTMG8fOroUk0mCXdhbAnnL/PQOJYVQ/vYk5F0rHOXoRBEgVpVOBE
RXml3Wso5tRxrfU/avH17Tz9PwZXhE8aXhTeIm4drmXGzu6jQVDzUvd6RuYEK/BZ
4QQsJWYluExk5C+R0dkuW++PA2VhyJvGwhtss7Ykc5RWzDz90YXpm3txMYogZGu8
qPNXMpd9wEk8Tt2WQp2Hi2VyA9tqvqL3+S7CcKYVM1m+lYXxoQNtnnNMbOh4LDlr
zhaLt3PPW2K5ORtsaKmsVwHZf42DMbHNF7jPJD41lzAC/ICEh8KyO2PbQu8gl/Bp
5Smfe7sT123jn5oAqXE4S/jsNBemcgoZODccAUX8SQ2YStcy03xmtpbvIVx+n0Gq
x/67eNrj+fQMAp/S/oS8nvRSr/E8LuOwYmkB/kAViVN98UCD+7auQbGR864rKmSM
j28s5rcDfDa2ua7qe85KK4JcXies/eRcn7z06xF/QADwQSIDk/19JAngrYVCrSgZ
utouePLMKR0XFRm6+8mrMUMa2Rv+Atd2L1dohPpz5I/jrQtvEVMrP0BuLI76fuTd
Gyx2H1dNfywUJT/wT8gK3yBad1Md56ThwYxf7mLubqilU3Q1Ly+4L9MbcBsXj3Sk
hmFNo+B2z0X1HvdzTprWtlvGJp0vy0V4oe0zTg45GW5z3D4gSnjDhXtXYu2S4D4k
VTgEEvIKh/iuY1YNdTgyrxUEVrPZ2FFRfw2mgIY8OX2LuGcY2uGEg0sRQ4ZEIBvc
+eHLxMXZdHuStAW99bO/ljK+cxkMJOSOSwzF+ccs+abVUgP9YTANcYhxE2eQYbNK
xd2rDSjdkLUeqbwtf5TV/ISFQ2O/LHTyZuBP8EbzWg/wQB/QcHHANwmro/bLNc56
BV9X0J5iwFDtosvXpLnk6ZMI4nW9Aw7qMX975XkaMjxk5xUvu56QjHg0j0mSYqdK
GLYAMOkCOQWjad1AbI2LZc/miS7eHPSQLWYLg8VtFzsrXdP1duSW31G43QVXG8wZ
0vYmRQeyJURZnRdrwW1EJ0et7VCygmthlxLp6qpdZKXRMecIG/rYIAEAFIGupUGM
CKddzmf5QLYY3L5Riy8fmVe0wjTYwkEomenvvTPjt0qb+xvvNY4Sm5VVqPE6yTou
PqyfWQeAAtsz6XbxDjuIHV/MCqIKj2i3ffXTzwg1D778tG86GZDODd0osbmPYCwG
JIiRdyI77lwW5JNBE0XYR4s6g5nvmVlDCkz/sFPY4MUWhsY96CqBOeRxyk0Pw4N7
07YkpLJwlDgG4mK1lqueW0oCNSmwBPnXmU/MeDzvXxqyJiNbWRZ1C9Db2MSZQmTg
QdRJZVdE7MDYrbqPX5TrGXynM9hFdQx4ITQbEPuLB8XmDq1prGBoA5WRZjFAMfpa
KomFXWi3w28ssHeBrxYECwEe5F1X6zUB3Yn9FJvURwRKkkRVG7ftrX1jxVf3v7jr
WeZxcqiDL4RHRL+sfqeIUQPCeAsj69UC+0ahYflzwASytYYegqqvBAIstR86zdVm
XiCL5OBCP1RqaCzef7tPKG0ZLK+zYg6ta2xidlcZLPN67UV1ZJ86vLqubMbU+/P7
jcA6CLdNDCS9Am7UWS1mf/5TY8GuqhTy48eVgxuMHV0nwqYal1BDQIDUAQkInXnT
f2WPnBuexaENuENYZ//pmgIeHxKDC3Kn9nYHMVHdCxonIHJsDSh3DJeJjUdTR2BR
nENqlKZ0AENG4R3g9E2Rsjft2pCAhpItPCofngzKfkG6CDZuE6+PLZy7wmdzuvIM
KYi9VWSlmwgz/yJXNDlzmAWbfipIJablDOCEDtASF47IB4PqsWHCGqhpotT+dn1W
uuvdw0mh6LiKoKSnYTPPd/L6asoPBhU1Hfks+WHdBoANmBohhrPUBVYdvqZIkQRd
1E0KJ5uxQg6XO+lse0gnoSasBKRloivbhgqD8VhQjSrHD+9flNW+zIxLlHwClyWp
oX6tT5yoRXKpt93GNKA0jF7fM2J6aQRfx5IF4HoazZE6DwBcamPdH3ahRav/TXq+
AgqjX4dmJwyobeGa4pEL5eQe7urdV4sIkHbeKuv6A8sJdlnAZRnsIXFTTtG+Yf8A
epfz39R9/p4WrICEeOKMXVzvDcDz4lavPt90BDsrFeS+5SeepvKoko/gqcknTbFD
z1SSj2kznU699lEfmOhxVvxKbTfMkyBoEGj5HgOBCLD2RmVRT7cOEMTcote77lp+
d5J/789QF1DFnrV81w7gXrr3TQHN/83JMOOzOBC3aXzzlQUzlnRQk1DCQnGv+15T
ScVyIDuXJKVt38NUnd1hnkUgtFgHEqnRfxeaDNMzK7L1BnH85BJHpLvn3J1Y2D4h
rMuSbCXG1GI9zEvVgcrUwhpmzYEW537ERiF7SK8rTKmhc3miOkCx0p6J4oBgcnds
elBTAHOb7CacbymwGtrY80lqpXPKPHIbTar+ssofOZ1LDcNvVxv5a5NEqPr7PLSI
EHGEsS0OjWA3q74u5h3moZpvYq3b6Dv4UKiM2JcindpeZCYlds9fSqEK5N7IPNuP
GmEQ+VBRMGXDbgmKCFEU1g4L0d4nU2nMPmqKjfFkTV4udg0CFlS6dI2d31O0P90L
N/vSY3R1EOT+hFejlAi1tUMHTbRn1I73C6AyqeA/iTkt4ylQw8ihPMx66LCWPP+R
LOJx1+r5tpR7Jl/uuPD6wj5HNE1+5ul64JTvXKW6sVZFfARBtTcRc2yX5Bz3K3Gb
SpgRTix83ASCLyyi8UI21/VmrAys01xf+wIByERcgc9vXr30JeotKwaxlgRbRpkv
FWyzBRlqMNQvujuLeNgKc0VBeK3nxLxM5MvManWHn1L0dOYGDGSVlka9fPNYlSVx
UG1MruQiLtkLQglItkZed7CHtiEr+0M/jxnx+enOVQvjowdlas5jpi5GgO8QOto3
QXlUrS1alBApQ0W6EUalEHkkHZsuLrE6CwFaE2O2S2E8e/kPvaAO1hbMm1iYOq4+
xu14fppdcbUnhs4SuI6qCAhC1FAjkcGiuxTILa1iEJUaq2cpF+UHLgnxkzJ4oD0g
a6H1b015FIlQYfAitXwulBOxLJcjUR+a8W+R9rvHY9VO4nN133sP3ucemSuCzrU4
Jw7O0fagaKmgV+GBXem8r77HTZS7s7nTyNiGKXMs4k+L71RYtf7SMZvPZKJt1f++
KNN9BAXhvReItsa4+HVKzjwkDhAwtZalyKJSuzGehELAQ73yt7Fa3PLf9k6LL8M+
eY4zHiwegeno95vN516/kRTj4Dm6Nr08cUZqHzUxY/58/QgSBkKZmp6MU3W20jeT
NxioBtHSrwgdOdl4wTBMzLFOi7BpHPousZzP/xhliaCYKAG3/h2MqDSqiXIBv7gc
o9dJO2YbLcRe2A5BTKmRXmEGkwpfucdq8F0T6wJX+H16LDlwA38k8Le7wBwjK/Kq
p1rypBr5tKnCCQZ73zsJDynLlq5L+Gix6V6vFCmw42Y83pn5kJLelIRaPHEaOfOs
uvQpheUCQC6mSzoDxOv3NjuC+X4uRce8lcQdKa49jK/nPuuPEOsckZX1jXrrxHeg
RbvK9guUG66Miy5bI0gWjTxMmO34c+bQcnO9aykHfQafihCf/WrhKMWC/sHs+wzJ
EjVF31DaeZmMSIZtANFYDKg0fcDyNYfJ1sucVLGvRvtdh0oSfE4Ikqo/ybT9Qhdr
yT+M4A2V1fyJECX4aMIM15TiFz//y5VV1Lo7O83RtyEhzMNOKxx+wucpceM6oO8+
9bP36RsPyhn+6oVBB5NQUvhoStOq6F4WU9+02yvPCxcnnn0A5M4zUr4jV/C5ktHS
nTnbeJMCPYxuySr7+ZaucD7pdxnoaOETaWzV7BTCmBOVNu0hZp1Mf+DQNohYpbag
HeYgUjuymSvcNKbPN83k6w4O3zRh0uXK5esqlJAI3dvDksiFXdOHJEpOSh9698Yx
2FwBP1IGm6Uz/JhIQ62d67yyMgQqL1ByNlbtLcgOFSn7Q9W0tivk4paMgz9Aer3V
G1bu55o4hAeVHQTqUfZMchbyAhWLqKh8qT8icPD+9pdzwz1pHfuZiV1kjomrPgFh
0r59Q322JX8vg7a4XU5Zg1gZA5sa/xSaQUBAbBKM+5nh6Wx9bO2T64ZNYVt9X9h1
vgThXD8g11UVu4NRuBf3sOMlOd/SCQlOX4DPIc1SYQ7NsCqjpaTxSaTnRqoZXHm/
vYUijE+Cq8E4DeA1EjP+8x2R0lyztCnXZgZh9QPUCz82aUXLIrc1EmElepxErRLe
g282/gf2YskrJEv1jlwtnoRY0RmADxJVTw3cXYiTqo9Yz/n9wXdFELLYD1457feN
7Jyw5mbjMMfOU7i3fm39q+qcuE22jLFc/SYSIoQ+4IkS9s2RzOVR5CZI589YRPkz
hNoETK9CaMLZ8Ghco7+7sdRLMjOcQiJeWv8hxQRmB5dBoT2g1f6PM5lfI1hTrOty
fht3gIPbiqaXuDv+6RnSklD1291hJ/RR1YTRctNMRM0z00HYD1FHSJJN5XfHsWsO
4hiWMKrrp9qZ3jBdVIt8+oceulleSF7nv+FED9zmaeCsPssxAoHKhYHU/7WWnShG
6cn9BDxdPzalu3dRiL0mG/0NfZ8+lQuBk/nliApGvL0DJ9BNeUGKcgLFzCfKpfbm
CazVlZ6glB88YXpVye/2RUK57hHyQ9T37ioQ3be4iyfSgVHh3mLnz7kuysvCcxMP
Mylrror3D40sggVrCjntjCg5OpIXmuQ++PSeLAW+pcBYV+N0Dg8uY6lYp55UPAbO
mSTst2hmBnY/2LlWsffTU8+FgK+NeImJSDpNexJRsvLnv61yyp4LCku0MTlpfyJH
7cbe7zB66xWPB16iwdrtpVFmLk8uf4sNCYRybrtkzWzDI4LW3h6xTscl3PlCy7hj
oFL3dhxPRN0AP9vwntdVWeCgAEX+KFbZmVtFzndgC9QNNDEG7lrDNxKUwkxKMRCP
4mxpgZNrozKPwf/8ZH/IbvFk0/LvKJtAUgODrvTYbKSqXdKPDoz3KKBCE8f2KwLD
Nke/Ajc4GTkmBZ7fHFJnsst3xjgoQ6NR2NWAElj0HvE+S2FiUoFRylzSFLDFcR6r
ytuDMhb29TdmKX8AUmvo6bPRHXcfa3h5tUf88eMvQRxIgYkpCv0vbpbgn6lGaeL1
Awa/SSPPanDsY3ypfZTL7WIBIUMGocKgkncuAHMmiZZxwhAigD/DepT3W1lIHsxT
yYJIKWMOK+OJFQMpfI+Htrga+lOBZBYD5l6Dbxa2PM6UlztRPkDXwfZ6tA1siG8O
7LUqL0XHt2+K3ALF/BgsXW097y80cE36wAiKVru0siVXU1V9aYXHHF+E4umJuRjy
aGurpuyfDdsAiDOiu67zMvGeNPiG3GYcDbM78XIy2tJSZeyd5dhc6GBJZ0j4vEKU
CUJ8kWsKx1DzC/YDoWmlSQA9fn2UgcG96BVUrGifazaRa3WyOh/QPCU+38qwPJq3
6ri7yGATUQPrUJwijdyQ1V2A9EBFEl94aytarK4stBmjZ8KGO7J/6XINy2o98yU/
s1NjY1SZjHBX4aMtayEzAB8/B4iAoGplYnzhAVtzV8GXtmZm4gyPSVg3hCm7OT1f
Y0iIZDQ106Cc8KtKVHfwmjvc502BsuiErX3BMHvAvi6LRUcMSU1RRm+sZDh3tnE1
iwUaOlKxKi2N9BPetOvh/ReQLVqExQYGnDB06UakLBz7v/mEWU45kzJozxfb7CW6
zcbXxbCDqoKVMvmzUYy9GTNfMRxxrzmg+XodlbY4PySvU7HFLUc+CeDa64/4HE1u
DF1GWwjnzja9buJSGYeQrd3GvwhSKgnysWR+vtT/ptCDVH94Uv9Lh96l/CDvSgC+
wnCaf/pskL3ZsI01oqdYAWPIRtnywHU0FsYVE5nR0gFi5uUaPoeirXRyuiUxJhlS
h73ukG79dT41DjnocpYgKrJKPWUeLF+c/U4IIUmxT7n8gR7f0XI4LoWy1fE0IHEQ
byLrhtuhQDmeN3jivd24ku9A1JvAHnFdnlV37GXV5BzRQCFbfXFIrt5vPVpfdLLg
ily9Vn1S5brDaaHICR4VWdXb7uyrazyz3n173NPjaExgBHuD4QjZtKnuYn2TPgX+
+sBtcuoxJDBpaIhrLiBQnJkuesAwXrxED3JReSOXvLdExaAy7fVJkCr3jDBJcRyB
Ry+qZfnp/044/eyj/jVOblYbV8jroPCvLnHMRyW18kuie0pY03SjRPrzWvR9/hsL
fcVk5c8F6NqvZREnKdUaOnDSpuoM4ZaQAvS551w3uzv+dA3GdKfAzvCkxYNV5k/w
JyZlVd0x7m05ek4AXSxi6pHZYePSZvrqpm2U/q8B1+sPzfyvp9zHBqYQYBFdDsw7
lXqiFxtkgXl21WpJVT9+q9obI86sxXTYIbhByXVlhiw28TULPMC3BGSy9nulviiN
tmEeZebtjc6M2v2Nkn1U/n3K3BSo7YV6IBqy6cEPNt9znZ4yZbMGXd9jrqXShaJp
D3eP/B/RiLBnk/N+H5L2HALgKebEAPA+cWCaf76rI+IdJ0mrsVp6cIlpWpIh7Y2y
vbWvhibFhoAn16Z2tF21NEJJf+w9cQNPNglguQGPzbLfmQQXVPuTbidLkEqoJOC3
Gs0T9zzIPfjzWdo4H2qONAxO03GLk3rgJHLmXYlkNrJGs/NRkrT0WQBa4L43kSF6
ZkUydAgAvZhBu1LTPfswaLUmlAJD5z7qUSqIoNZfBD3BknoMsRFCV9bb6ng5MqUX
8suQCdTNHDdUfaeWJkvPviPwbOJGez4o4OZ1UL6LoFLoQ+hZWiiErT5okqW7b1tm
rkPRACj4PqxyHGEE5XH85AW245RbRekfhsYjD0NEsZmbK5WEZNMNCxcxNFNCzzya
mGw+2fVcEgWVCmZON1gAfzFEFRVtvWFsVP3QyDBOcfbH/YlSZPSflhUasBO+kDQg
B3HPg+26A2RiVpUXL20whPpwU635jucbumn/yJWXJ4v8OJ7nxtWiAj1fY6cGbmgs
pmTzeGo/FDrE55szEVTsgnl6YQCrAtK9T2IGg3/tCQHgNRFllbZ7SgeVnlf7jgaJ
z5tLpW/VAS26kERVf01mBaPt3mfSpadb9RLnPPQFATCEaBSAMusIpbPpFBw3UISD
78ffGhTCGIBrqPRum4L9BbKNq24Ofe0UG45NeccSFPlC+sav5NWQ49FihPCd/oKH
Npc+Vb6C1dhCizaK4YjOfTLBaIruntNqOIqjJlfHDBKVJJz7zYtDUDy8z8yeR3Kb
r6ZXLuGEzF5yywq2uhf9UPIXLulldoT/ehN1pFkhyWDka7KAZ9fhgmAel0yR7QPI
ZFY6QOreV1DvVOhINAHGmmcyu93EFtGChBKy1zT72A7eLCowFXeo4Xi5lHAXKwEj
j7t1Be9tsLoM/nX/Wi3DxeId9zsc61hZTpomngKm6+mcpAvJaQDTseGrkPbHBMg3
kG5ZRfvAs1y/FAz6oPohrlem9YgANzAgjgPVfwPRfbaMbVlTcOIvoCCQFb84Wpx8
tQZs+q6r195eqCiAXcxptXm79WUDenLPrT26+MIc8VMUUUPtcMCBRruCSuRqodXL
2CyxeDiOO2QQ38V2pc280b5vW2b/KWYzJ7ikjH20FW0z0BiWcYq1Uu1CDi0gEZ7v
i60iPVD+Eg8mmtkg5GJxavpdzZFbn4OpE4hYSzQRaM0f/e61TdzSgPGw/9qthUt8
C8wix7nPMTaaDsIBMkfxFmyZgJtRXgDzBSsVLj8WbFDRc/vU8W1rlE2i5A4bIhvo
BlxRoxeQcXfy5Q3oSwUfiplvu6UKaK9dubfd3UBYvoLkfc+htnClnU2dLS0peSXr
Tak23qzpMiy7ULCM4Wg9VnN20uuxg7LvlDtVrHZyQFfKj+pVD6fjq8GOYSPC88dF
mcBINfujCwHk7AfaUEYtPnn5pogN16Ht/u4yiauit1QLdT1UqTxAHtIJpmtg0mBs
Wd6poh4livZQD0QjMIdugdTknllWJaUGcftjaGg0RwY7FstSadq7bKYIA7TZ5ZeO
+IOAH2k7HD9DckJdHNUI+8xcYux4m2mJDY4CwuvSa8BO/UdcHXcw4V+bD6KNpWoi
p1FulKjTBbS+jcCpIEvPEJBDkse1Lnw5Eh2Sc9gB1sTnnPTA9xBJ8ODJv7nqGjEA
MeXZSy/d/X4rodHkOpq12j/7KtxCiPKxAhm5fTcCOAS/w2X66xj4n84fnj3PvAqI
8eBl4JMpfbHwBHBoK2A0BT3KE3KzaAKcEKhzqhKnuZ3yuD3lHaYv/MwgPXE0Fnko
rNASCWUkqfLPiGL6THCUgQSwUC0u+L0BtNXn+naW1kxzBZKyqk2qkXkpIxmM0Cr3
vEfaz7WYlC/82SsTVwI34yxKlB8D6YmdsbrzlNOsb/+y7nu22I7oRhOjyxnML5QN
OnSChdtsFT63JIZlbpalwAbChVOusdkxz119lbatcxb945YpFYrz7lXeHdDjo/2U
jHNMA6QeSY8EMIJZWmmsJIbHK6SA3AM8K9yddQ0iQBKDggH7wQH03HoMuEIVno4N
P1o4f2UUQoMnWjuig1Yic4E476lkfzXKhOwA6VjXdWHQGQM3cOvu7a5TdeUa66GA
iq5pwoBYc+0nQ3aXBVlFeWKCEThtULTCMmw3zP50DrfYDF1vkETkMAAsVj19Omwh
W0RXGagZkrrlZyuyjjx8kp1jd3lf/Y+JCy5P4bUuzSYjbOuN9nNLhNtsoVaE+YLQ
EASGNnWcgNunmeaqguKpkX6g64KU4ue0d2sOg8bC2xbqaen1iIy3yudhtpeUbR7x
tO+KBBk0lzVfvOS9dPczXbq4LPzlIRDm+5Fg99wBAS8cmT0XvZFa3gMjQjevSX+v
5axrmJz9EmPj2pt+kcNQK0IyCOpANBpebJnzrk8BtYPHrmnU4OyvDQJUEroWjHJ8
OjXPDjwUWtnlHmUOH8fum4hgJeeFLDw/M7HiqxP3/yoLdhAOeyMYArdJEWx7HEDE
3RyORHmvXPT+aTrZceZSmNOYBPAurrme4k8xo027h+iTvjEgqFXNtq0IhOrauSJU
3MRh1EG3Z/13JM3eUZ21NAWjzz+r6U3sD/oeafsitTqX2pZ3oEIXvHRWoct4kyHU
lEeFgcaD3wR9cwPpKp6pJnseUfSpfhQTWlla+ExkGEYHYOJsLoaZfQtybqez+EM2
q032U8ALfMrIv4FmnQjRVLMoEP8B/nxypU2ttULUVVvbpAVt4p6LLo9PLJlvEMFf
kjS+dw/oby0QoFLKUGQPVDWTofjYctksuscz23vN7QB52WEQpinOvLBNOW26/bCf
II/hBVXayHIEq823wTRziYmndESUe+zP9iCaSFw9BEFDbk4kUtRdivOQqK05IOPv
gZO1635d4TZN4PAAncR++qa9EltvuB4So23QglgnhIM6Ryws06blLnu0ehkmtEYE
gxXAsj6KsgFRfzXhDglZqoviyAXV2oS1qXnQ8nHtlbi2RazzGawLBA2R22jGegKY
wXZn5EcfoxnW5p+sOaF1sez5SDegy/7Nel5rPIE9Fnsx1Ojq8ohLQu3/74CY9FpB
+xkkOuiPF4L3o2b9Q3U6NjJL0UUi93cNwMuzpLfsagvNCj0FQ6QPgICO0ooJQo84
YNNC0xxRye09s/LkOXVBqmi1euPvjSshtem5WtaeDejZZR+Vy+XdNFuq2RbV3V6z
rFZRSY77NEnyWPhHRmt32d+iIplAvImVytJS/BAdMHx60/KAEJlEewp3tOGVELxj
E8VlhEizALzd6POIeFw217oVcTFY8xgs11MxDe1LE1s0T2dXeE8GIKcEUljFNZhk
QNET4ueiwX65KNQHX+mbyRJROr64/ldUZI82mfLllTnkScFzxeL8Th6fmlRSkFhJ
iuanUtWW00kJkHxRolT34jRXcD4VSeQ873dDKa/MDrG1wgfAXae+oTNO/WMkfMTn
MQWwgDmp3TzQ/grCRxlRwt0a/19Xs2MWJhlhFMbUik9aev6iCdBtvjx6k8XGNOEE
AXpBH7NG4bmmIVTHoIWLz39uhpjT7vXi8BrnogCy9t/PLfincyOVge5v9Ngxv6qU
M2mtau4lDVWJd9c8fISRZMwvIfiD3OZ0myfOqefdY3ZjBAaphpe0AX0TRKKpHkA3
BuqhFwDv3ugVh+6FoYxX0MCcw9SNgjKBfhdgRQx7bfM0TRYfSrVZRae3mpdteViJ
WX/YegDjVGWr4yPpErcJVmVYlELcFMWXTNbqm34zFl2/6RxMejF9ADUE3fYWtD9X
dKVVQw2PM35x7T6WkUAfSxYvjR1dGBnCzRyhmHfVFxUK+ZPpbiISU1q/FyYCE/MX
NwZ6V+UNf2jqxIkzGkc43L7giaNfDARk042wdbOhFJ0wYFMJZjHxEU0d59enzRVL
JKD1tJGSw62BemLwVZPvyKHJDYcDbGVx8+uye5QobTd7zv7OHsn3WhWAv/BD0e2J
vGf/4xDKL+HkjxOGeW3rm5bEnGVAzwAHeZa135IcWmK8scGcndc7XivO90/vw/GT
X600hRoX2jQ9w/xRqwcDGOQxPPKIdTT+oo7S/v+b23chUUsvkm9eDI/6VFrel0Yd
f9BnVtgDxNv9JlIFgxolwGMVnADBjV+1bXVyEuJDn+IhFeq+mHWowoQYFoDeArj0
4QOrm34JVE1ye9GrwJgOAgmmGoRdh3Pnrpnm+iUIDkCQfVwY+8m595YCYPJGtwui
jzsVH3OxuvOJabCTcuDlbqVdRnFcv3CFSYnf8wSjim95/3VVHv6zJVyKXWx6QlzG
QuTObFYXNiC4i4w9xnfl6nOl2pDrJbRYypHrMjV0gVC8E3ZvrpLddejwnU//FOeg
yiEPSIJCkONXNLp+f9T4HJoAwNAO3ynuU/gFFvM5m53AbQ+BfFIRgZ2zJ/du3BHe
OXIeRG1uy/G7R6gjN9pvwNqImV/mgeWZTSRwOXj38PGGXuGQj/snJYl7cMLblq8V
dJ+kqMR5ho/r+iTR8KOqAVqzJAzcUL4Iepko9kbKfqzHevjki24E9oQcDiCgfE4D
jEI97EoG+4qRBgnIcxeAoQcZynyWsUoon2AVy9VujlUOWitzKviDuKq1qr9B61zN
ezt266PxYJCjszrwhZ5mu7FWFhJ2hBuwoblfUgrpEOzWshEsIDr2XCwM57mKXmHd
+rDfMIXSFjVKqhzG77BURkbKFyGMB5fI6v4tc5ODzV6/UP7frBGzw6GE3sMBjdxd
zVJfI5XkqIUY8in4Nwrj1CkuQayWwYMrAYgCgh8wDQyu/zKtG+DyO0i2TK2AXZtD
5nIkPVYYp88FgIy/cb1ne0wJkl7exifiWBwg6B4zfhFc9K1ALdsJWEsjER3hH6zi
qPMyGam7LmnCPC06J0hlvCvFbTBj+wByJ265Tw6X3JoTS0sJVo5N6rsyYWCV1IqP
+vv+N+4Pvw98C6R3BwAj/HxpRskOGUEy7Q9s9qD6TiMKLgR7xVsBLR9ECqG1eC3q
CG/VgSGanRt0epuI70AKuQj4BNrxC55ix53rMwqM63Qs0HlUb6hMdwM+OT02ewle
drSsqjmdc7olD0A2ADBs4fTKVsIzE6rCNxcGxXqQcXzGeKGAP1OP4ui//u00aL8r
wK4rU/kQLCh2SWd2T0ogSRS/RARcAkA0EqnygHl38WNHPzu2Akw1pne7G9PG4IqI
+ETkLavo/UrI0uWOcQKK8MB/8p2uW6K9JaNchzVViZ2fYUx/LJBGllZXbvEnV10h
QF786YinuJByOck0wCumbtTYFFiRmzyaqKRNnblbfDJaxHy3zAmWwGONtmlYdDTl
aUWXkLGIILQQEm82ka+29jpnxgXoQ1bVcLJTjOhFC8ZeR8kolJT6otMDj2CxQgy9
9USElNYZrVVYb3r3+5rZgBXBzKDSYCDVwJlcGVGoWdpK7GlY3jVCZ9Wn9FfpoMR6
g02hYUN0kGTErHATiUTvEU8H96toq9N4maY7ZXY2gYXorjZtejbctPkhSG735Tj6
4lWM/PkJW5SpL1x05he4M61FB3Ggnu0TFCrrqVsmyICuPVr2tWbNfy00l8rzWWja
0h0vPxiHQnmOoF8IS79v2+ruPRr2Pw1QN+/2yZPrcM96Z+qQNVIHUJeLbP+Fjj5o
U4aMKwbNHscJjKTTtUWsWEA972GJ76zWnRLRpmEI0gkWLt166YqBtWfWFGgHTBlj
bsmFh2EwX/ywfScWtdxX2CXXR37D6hTX3g62fdvV6C4WYCcnussvoXGJLLAvkJvd
vjwngp8nc5qFeF8BXgFoSnIGv4BBpRbaD3cAWzu+zkWUol8pslIj459D7voOXMt5
uj6cXCVlvIu5dPnDog7e3qjfJjW4jBN507c0NAMiu1ChjgPTvIiGruBmdT7uFM51
7LUODhhJNc0OyshZV7Aul+xPl80DbnJ2p8ZWF7y8MEWsisGuskf3L4QKXl/KJG4W
BJ9sq+AEuhZP0xxTV6+n0Z2I5zIt5/9Pm15cIHOLEPWzfUMHXYdf7zxFtr7fTXuk
lKUcFIwi52Wgt5Kfn4NIPEM6G1ASMz6KPeJqb/UIlyMa7jpRLwqxRlkcrBcG2snM
fuDOrbGkW8/biO4ldwSO69DnHFkqKUsPyMRjvMf0WCjORAJnNXk/dDU04XA31V4n
TSDK0ZK4jqRNe3vrDXiYMynunDRbLGWiFeEiUZ7D0JUK9Y4IHhE4nSc+4a29qjze
yJcnEsBMigzPKkdVhoUflbJPvV5vZXb+HWb5gC5tvrs4c7sxT9eAL9kxALcKcC0Z
g0oBMzFR7LlKdTB2yFTex85drFlv8i7waIAbRRC93E7hLUcF5W8oKDyzTrPK+tN6
N4E/ZaEjBJ8nV4OJmTQhqXr9jUogXvByH7ufUFsQQtbay5LlXsByqLs8bpcy0V4V
iIFBDefYhQmyoEphJwGgjNCeuCAkklB+F3yrT2drVQELKdU0Ez0drGO1in/PeU7b
TZk3Jy+nszO57yWK0coz6gZQ0O5jzJvo6YsXNwePLQEaqd9ZvqVgurw+zkgSuXOw
vKn1UyFFzt6Yj2kTxjK0suRZ+uysJ6uDpeFsklQP9wvytgLAkop4EsR73C8muPq8
uC3Okp/OJBgSHopv1He8/9kM4C8MGc3oIOk99Y5v1jDqBqAk5OfmK821Esq41UFf
iBUe2kU5bYIeClWiC/nBvN1rZnqS60wGFDaFXJzS21mt3r0WbFhdGbkeUtVRAs1x
VmSQi8qod6AWsE7UFYviYPTnOh93b/WreQhkCT2LMfdVRmdupvkWicDHSBXonMZj
ofS2yAJvpb8sEmgbVEmbV3Tr5OcWyBwdwC70sBe7RP2KwbDvVG+kOYxO3JvjXvll
jWN7r2qKg4orYi81TLxJuau12N3j0uYE1BLbh1We/o9kU9Zms/0mpre6iq5fzLYc
b1jr0w9uz6NlYKrEjdTA7asY7Gj6ogrVRTqRGyEeZhBZTSZNrvvMCMRh0E+MLrWN
cjDM+O3mif/5h0Xr5S1kVpI7gZIy1rSR9vbS0WgSn+RIWixvGbrBlLHtB51KFYOP
o0poDlXFXSn8McAltHseK1L5+NmNM3GX98jUIx5STu84Z6PgxN54SZ1IrZlz6TuY
coaVw+kfyrTpx5zLt/Sxc46ZGlfrmm/UH8WakaygZUB5APz6ssrYyaNEpPNXY1a5
No3qVPrB4NfDqfSpgjDDP4bKKhvBqwgdkmVPVqi/GWqQN24JApT/iS45T0jP5VAi
4QQvjr7iPRhD75yIR9wWuXNRjk1NNYGsaPC9YYPTXMEHX2PKKGUCTA9a7wEbazDj
wQSV2vcRhUG8iCYICi5BEe9op6pL2wphKCEo5fQg3UnIPKWFxBD0MsD6wIofHDh2
OW8K0Tlb/5b3kAoYFf+qq1taHOAzpTfUt/ycW/a4SzMkT1vaMjlTnVe5xT7soXfH
JoK3OCbzQIXDaLwTAMaTUdgam+LEfT4zlQwmeFf7/xoZyD4F6g6cLrBtLEibAZfm
nsZ8rqKpPd/EIJw3egLv4qJyir5aiT+VjgJTzjijRYcLJviDVnhM5OLAaIPUgYe2
RwYcqCbjBZT4+FyepLWJlBoFmW3dunKIqERjih6HvHVUOf8SYBhNy2HNE4W3Sjrn
GQ7eQD6/cDicp0BfFIG8qdCIL6G8RfVphwrelT/P63UgeiAYSE4eFaKb/+stC2Lx
lT8Ftrd9OKWz2mt4cM7Rnjrd8CNrBqWgffqB/i47XSRFFh9D7P6RvKP3n9LEkjBb
dsJqFlHqm3MAyjTYhDDZjMfS39ERfuJtY7T6TIIvIe4kSgYfvh1jU3Xl7wa/S2zc
VwR61WoPzVtl+bgCySJIop5smGwWcJr0ntW/TUghrRFUkOzZBeJDCxOkOsd4bIKv
tdFUeFxMJAO/6qAvvnEMzoLPJFnEKJtsUS8OOKz9bX2h4IHoPHH0/ztrHoJBQYJv
RR/TiOXalSHLFk6BLSa6Zf22Jj2RVrMCMIl2Ic7WlO4viIgUDCVfq/yoR4ZnZdc2
kYgff6vIFgVwkdFYg7GNZdd4xN6HGnrgBxuymcbrOX2HLtrVXh3kFbTv6CWOS/m5
O08njKMUmjhzCdnNPPWUgZ/vk/R15eNL1NovB0Npjx3LNawzj29RoiVMZsOsspEf
Tp3eOwZLQmmCGjzwdA9cFPR8yNC06tseABjnpCi4mazDXh8cEAh+j5Wd8+N6VcQi
aXPh6wm4WExw6JcqELck9y7OSH00BGmQXSniJe/GWAzKjIXLrbfnl0HKOp9i2A2l
zuMhxtd6q2uk5yk3JDtDuKIowQ6/uy5CnDiYAlxjhRd2ZKwetJzYtJiZ4equ0DW5
goS/zE9WtEJ+/RzwMuZFTzZyO0lcC86bln/e9aIKNWBiBHQMBbaLisiNSW69UO9/
fxw2b7hCYxkuxKDZsZTCsxGZhPWhcAPosacgsiMYYxnLsXSZhvd+8xovPRCnzYqA
70pIAh5BypPQGvy1WBgD/3GJE3mm0kwFc8P9Chxt9zdYx2XAa9xqSAcia8cNu3+D
KnV6bStat3MpTcAr5h8meA9gUaTyAf63h29FBzi5LTJihGscA71PTUaJ+CnznMYq
31hANtf3BZFicGJ23sd99791rrHEVaewgrC+pRFMyfoAaKl0ZgmxaM8NdXxTvxlq
S/IAxf4IIxqXF8Rlcrgv7EvVDD38R42zgDOa3aQDmwr4C4Q1D5qlezJZ0z31byeS
sEhWrorM3oaFUgCXhMT9hyjNwYzoyYITBe5MEpbAtOwJk6ap2jtJFaPSxFvr3Iwv
zuo8eHpnXfIErbIiRtAMf2tuMzchv59Oh17Fe97/GPJBXHAmeTE0RMUM5lmYhssE
21+PHC+hSPOHaoq9pgLmS8NjFtHyw38DNBsYcEjzf3XIfq0IEWev/+ZX2ykSEJK8
NkFAvaOfwNE2SFZ4UrCV/yQ0vuzvSjRIfOZhbNB2WvpeDLMAxZmX7yEGcviPeK87
/yLpN2w/f66+FbZxoGN8crt2jtd/+yebNbZ0sUKoho3xP9HQ7BI/ICwnZBH1M2JJ
jLDqMLIQDpKS6Q++/ge3QPtdJMHh0llJGdGFfay0FdSJ3ARWe1dLG1wsnykTyIm/
h0FTcNJ0bYoUwPHr+fl1p4oXCnw/5adiAgDf7+KEIUVwFCw1fvYSXImzYxqBoov5
LXJF1rYudn1yRnX8XShdZRVbbt5ChdEExMHrqU03xZ2//vfAv2DzP5cMNCWC2/08
4a/FD2e9Gbwx9jlwH4ShkDc98/9ruxdy2ce+oZZjdmqw8llj4kmqYn8BBOfQgNIy
zt+LXUaWIuphn2CxxBh/T7zVP2W6f4kXHVrIno60TWFSUEX0EuvHk5Eoe6WOsBEo
t6F0TSHgDrX2WwHtJdtywaLTP2EyFJ3mjOhYNZKkXpNBLzyjR6XYCmkbGKAOCLtB
BncV6JzCsxBsoW2TQKAtQDafqjx9FuQvBk/XTekJW4P+vnf/NfU+CpNKGIokfB+g
thhJv5ootQHtn4toeQaysPHFSc4/wiZsydAb6HWOnBAIUOE+XwJspGkKf8lY5yZZ
6LZ45yUK6A1eeg55bbQfYTWL8iuy8cb6BJfg30bvoMoYFSxBZWZeYP+jKg9H/JXo
VKI0OP9lCuFP0YU74H/uc/P2B2xXxAJAOXIdr3lX5OWPZh0va1uBgeozru1FjlB6
f4Vg5J4VTLlJULScuumz4kEjc/oVRuRsScU3xziQbZTH+HAH3ozLivGJ366KqOri
EdfPDpA4zeSQOWn2ZX85SNiH/ZrhlX1Sl1XQSxhZVux37eMoU3y4eMPGkjcNNI7q
uuEjT7q7aKNP4yJv+fNKF+AJn0BjV4L90ToRFrwHGYWZvnfAlby8l07tAewNKoun
aeLj/4A7BXO13/OJBwsARZTG2G252l5UNA+vvJQg5qMsHtj756ZEun7zQqzl61GW
OIkfEisz9xONJLyZZP3jjU0yhFhdnouDzQAxXLLef3t85/Rfk8XfJUtNLuss9T2H
Gd68MCPdL8uTBN5H4QtryrnufuFNW7L9N5DoojEzLpz6dWj8ZPRWNNj65lX/5xWy
2gU5MS/uOS6loonjUtDeHcroXxOe6ZWfVt93ryLKvJ3m6HW0k/QBpM5Khu4UXcAW
FfKJ9pXQOk/zzZHq+lDEcu8mLD1kjhxsnQKjHy3oqcKCytHZJpA62Bcg5eV5JSV7
gieCwtwoT4Vuy1zkxIcx+kkYfLlZAE9Mvxo/NijSCW7fwAukeuYktzskGxXuDaBN
7ePg23gfyqQcVK6qk/EIsDFUI1K768C1n0AYyHCDKjNDjEzkvhhxt7ywhMLe9APH
T06lst5XV5rvBuyjZ/UWS3XuSlnMLBmy+OaICsXIx0mpATy/ZRCUf3+Cnexghgue
I3Pdb0dBB2o9AZTm758hxv7glhP9X/A0U0C/Npo7nsREzNhijFO5RuaV7JGRI/Vo
3GlO0v4OFTvUfajiIWPxewYqVUKWybpTjJKqukkPYZMFqwotuetG1IqaeUrwsfHN
O+KFiqp7SeGt2C6moZ/hH9ssXGPG9FeLG8Q96KkrciNuf1gcKGcBSNi6tdT4RGx/
AOvnaGQFMPt25EsMy1gZQhTaAaeldCX4Xe/uBtsX8y7zZyTa/aw8fgx/PsiSubWb
SpX8bPM7ewPhfbQPOtHcUkLLFBcHobXMO0gMBTfymn5sAkEqEmcLMsA3O2UuH8rM
zOFKrT9FsGVKZ4vaLx8G4EY3CRK0gxLYk3ry5UKFmrq2uU7OsTSFSjaEp//8kcRY
jelswpmOnHHlpsS3ts6wvi/9W83lvxJSmt9oMmno84n7cFIMH4bEML+jz9CvUp9i
bqxHoPiZQYDUe5iqmW5KqC34TDstgv3YALXRnGf7QMoCKiDOD5fkBiqVaG0nTnKr
JGnbbC0Pl2iy+GdrWWwFqhOro5IDBx+Ol52qITGAxOiTi3qUK0WgIfEQo4lkK6zk
qk9lV6jyMCSv8cBEunKlwmlCReCLQWMFdTpHynHOm5vJpc/qnqzHTPqtYSyhurrm
6Jra8jdsUoLFU3nXlT+2J+77/HPsmjhHitL1m2EWQMSqNXZ5yXuEZheCXrzHiDcp
u3AbTs3RF/lK5zB07F4k+kXFK0PM03VtNsgB9cWPvk253O7A1ZIOQLZfoTaDq1kV
fIVIQjPj80aIuDLxEzZs2zNxgEYigq7o9ZmZqJLbdnARbutNPQAnBziBpH/IN/qR
iE8qafAkNby1w1XqyCaybo0rVWNg1Q9yggbB/sfddny++UHgmpydxa4zhbJ9b28f
3Fo8jRcuLpnPGWM2EQepB6Q1susNHFVUchzBwHcyH05hkSOoIk6fht1XonSpBdRn
Zm/43XW3LfYf5QW0+XAuSGSnRUpuCM33NXoAvnnJJxXMn7V+1MjgTI+9ALBkkEd7
L+lll+a8TVLSSzpymBdPAQm+CUcA63PcKrzdwamxuGoJKWNVdQ0/otDO87VIv9+D
DtX6TYdZEAqh9a6b67P9AnRHvB82W9G9DqWMRDotPM3T/1coHL4zuDmcmdvE1dNW
1sOMsmhj4HREvgHvnIGWOyA2fyLXvEwE0UTb6XwvoDdgUOaibw8T28AiOHWVvUFQ
WtmfPtJhWoA9VlcpCEhjj5LS3BjWA+LCKKnCPl5/1bEdAjqd1lSI7hu4aQLRu35G
32pz/6gIwXkNp9UsJ1G7h/kYKd4KBFL87c67DZtfbr4vRPWxGDdqPrP/BpTbtM1f
Mq1Mbak7l6cM1HsDLUvln++QoW1lsvQ6QGR2EGORqSC4BAeYQWtQ4H0QmhgOyQNc
g6hxaNYUBysx6jj0wmVLZ92NrX+wGpLRE59tMZlEyaRy+6rmqoliBP0upeE7E7bW
84HPXB7Im66Z/gXNZtJnTjCBqiVNJ3WNAAnsQcKJl+etxnQduVYNp7ObjBB78/fb
FUxkTXMJbgUfNFcWhiUmUCPBS/R0f2yLpK2TbEpLnf6e23zNnsyuO+hVDk1v6QMp
wF2n+C1TpXryoD1VshGWaOpMGcbIkUp637sFp9C8RPvmWDAaClAnMLsJSe+4/z8O
+WWJcHjN0hdZZzklLd3Ppd8+oR5KrqP70JE9SJWIZHSF1Hiewc+tYwA1Fo6nnfb3
hJfRM7zSJg2cRAVc/VCAL3jOvnDphw7gd90x21/nSCUqs0gnGPNoRDJemXNKdCVx
MYuvqhieiDpNUFa6SpLjGmZ3f+ahsUAMaHgTbPvhC95/rQ9xCwBwmG1Ch9b3d88j
9YB7H1BH6PGi8e/cTFvN3jV0+hbx17V7ng8YiIVUsNmmyCHaYTrglw14OPGxv9NP
jniKMzHE2IkFDuI1t4wq233HNnH/fSVkOnlYgpFFT3BnP37Mn+FwpnGvuad2gDQ0
y9bRZJ9fjLWZn5l44+zvDQoruZEXp5bqgL7cFzUVnvl067tRniqBMvRiLgBpAaZC
7NCJ3+iTdFDRIYrLcudpDrrhnT+6iwgcv/xqLnWnmJCJiVc7wiDAXnL9KkceoERd
olkkZkjUx6HY49a+uVsvkl02fYfMRdgkxaOrJkWrW4NjHHVHPqBetjjyUyfys/QU
COWpu1/D8FObgvHzrIHvLdl5hshQDmHiOsafc+Gv7brCNcvYYFOhcKDEqRizLsYw
E4UVMmPQ9tWzL3BpatdEAxDegFNqDRkn1qtLn7WX5MJr1d/TLaFxvshjR4zUkeyG
vyXDiXM7acCof1svCjuvNeSIeQUwDrkPw5mUGtkoXR2LnNLr4Yo4L5bScfyT8V9l
8jAzXDPifw6jYxwcEYo5Ib3aL5S+6seQBh5SX6zYhRiSOcUx1Vju2Co2JeW+hPDR
JIna4pIisCt55qpUOyqafWREJVHDFGKrZ7Dyaw1O8QQ7oamVcA7OlZHNpHKy0977
y9cxZ+owRC5vpjvs2FCHVt/j6ofRu1M3FxDtWrusYtIptYUoqXKrq7EWRBeAiNL8
TD6dYn2q8htcSDrVwJv6ehMetHLYNjDdFsqO4LZ7VUJpHA85FoIIEgoDPNUsN5RT
m330AIcJ7FY84y7Wi18GLRgwp3PePl+Gas4pqOHDxKABTYHgr54XxbWCwqba3zvm
i3svJoyfOfIBF4lfagXhMANU+JPRoBqDxpmmI7KqqJbkQBPx+EljWqpS8yZ8Pori
4+m9q08hVk9UThAAkiQnDqewkYjmH9UUsEPPDWXoaczy2DGTj7XiJDDxg924o8vT
+TvSBXmppMD0tD1R39st7hPGeeyhKzcPQ55nvmCa+PZAigusGY/n3+QLaaZYTFst
moT6lpQeX41I7dsybozZ4B2dXRCyKrPQGTy78mzlZyT2zIKNCS1CupapjrQ5QSPt
kZSHiP+TTx+lR1rgCt1mmrKXlH1ZS9g30pMo1faPfkN5DJqbNmrlR7w/fRGsRX8M
QWOowskcgKoUhxG8dwqZkUoeb2GTr1SI+EAuXlz6geDhCdoDBiQRZcfqcohWUgPl
40QN/NvSOy8SU2hYGe6hqpxiXM6h7eQm5gBTcZtgSH0ktct/jPtkv1Oadb8NuhCa
8BIOfqZ6Iqzd9o6t9v/xpxsUAKi2QczAK8REx3ZAhuxgSwmq0ZSJ+zUZn+Th3Pit
lIOAq6672g62wosCQsDZz7UdBR0sF6+ROonrHNOlHXyHTvJewQtG2KkOnLkZ+Ubm
3RkYeKEQpBAu75zWVdHab0A+CNatgKMOLTYBHavYJnoF7dEzP7zqfabhpkqCYo+e
ySPRq4+zgbiaCDrT2iqqGsPQVyvA5XCOmvtmE0l+YEQkGgx+mQ1nFbVZoFYIP7Xn
Ouebb55ez12X4OKSsH6SDro0Xpf8R7ulpm+InfD6u/SNBejzoqovC4VfrtXQlYUW
b/c+DbLx/l8FpUmZZEFxNyvavUKL+v0vWEKYaOMbYqlUGfzop3XiFtXQP26hcGgz
BIYPuw9zIpjnULCLyGqBMDLGkHs6IWoKoq11ZfpN6x/AuLf70cB8ao6muVCettdM
k+LL9kQ7Bji2xNqZEgw5W3YeVOmIXLIPhVCMtsCSHe331H9p+A/doKbWC/CwYmWN
9jLLvWZOMqBgJWpzaazjcFr4drDlG5hCmqYuZceJjGCU4obnz+Xgr1+eUUycyoq7
FbA+RnmVWPj9ZhEtpNZKcs/QTDjZczZUXjYnV5oKolLI469KCifY+ERpHxSdN7Fi
iD/ys+T6LOuNE18jz/0JzqqsxOefk3mubt0nXgjAf2neeMMlRlPcsBpEMxbz4L9W
pb+FfcPyxkUQ4yzN6GoP/cxrXxDKx+GWvksLg80mHz2/uXMcUei8CJknpL0losjT
FhCbnVmDSxI35Wibh5/uUDyuJYQ4NVfvq3ZN8j7MBvKYTP6aRwojygAuQgkVh8In
7qgwLpK0Mwgp9z47f2FrBKV6IbwL4s7PKCcwiWtLjemP0GhNczY+Ba30hnwdqj8j
MNI779a+crVlPRhkaDiVxcfaP7Te0A1y1DsB3KA8/rrY2fO4euZU+iyfKcB1MTrB
MM5KxVew3d5xPGyUuP9b0jtfx14uPRdiF+I5vyOLF8pld0vxbMbiKoKff3+U3UId
zJoeKTZTWtBJnzWbq3ls7C2XDeza0Va0UEbQ1FnoRa0nf1Lkoa+sI1rbvyEdcZUh
75b0i4BlBvNQ3NK10vmGZhXFaNZtbScigep7oD5jpMgEOyVd19beCGRtoWJTUy9k
18wwXCOMWS3DayaRXka+uZc3pT0L2PStJiXCirTBpOMMaggD8mC1+i9yG31bA97c
dAo6yrBkbvGcahHcIQEnfHm9G+Ndw3OGmrzXaG2VqFFTUjBLIMsb3LcHFnTBqARs
xVAGmKSES4Js1iWnNF2/hzhDoPU54gauPPl/5YYq7Bz//WgNV7ifxGROGxe57YFh
KQDpylU9p5JfL7cITjeIti3a7fQa6pu3dDMyf6GA0PdM05jpZjZ5d9TeznKjX+of
WZEw2eAwFOl08k3z7uDyjg6/a2lSj/ME4m8/jzV3hwNgV1rBsoS9a0aP0EuvK5uv
ne1IsHGdpiKYnvIVs8Ew7fWG154f4JpwMt/Ds3y7Z6SbXi4wKs2O9dxPwgiJGCEl
X/ydSUs8WmEijilovscSv/TF9XWFJQrNdeWVOhMzno3tQnPbRY3FqSAhwspQVrF0
5s8/IaCLc5VGRHCgI2dAm4UnAzWPNLjQrD2CGstfNjoRUm+UxMLun4SGZAVE6Xrb
OVcc8bnpUkH4bsAfN0TmtPggDlAz4xCcYQpkeVxr/1ts+jU9B5gcxTK9cM73ngLD
7oUjLk8KaJZfWvAmkAfLEahqapVGxxD72dS7tkXpSNOvy1bkKBx8S9ZZmKxG7yOU
ORoEUGR0f23kufxmeUP3shsfH9Z6+LCX6HdU4Q1gvCmJC8OyYjGkmCZwmL+EiaII
24NokiT4V7KLw5uFOmTGAZj3j+dR7Pk5qJGWrdgj4iaGya7w/MliSeqJ//q2W9DM
PmLTCnJwjz8FHGUSW1q9cEjKJBHXtV/ze4JJ8j+zbUCbZteueblDBaSPGTBMMQNt
dn6JJwIfW0qwXtnvaPIcQgVuTdIoslVgRdddYAzCwiUJ+zzib1BisKYUbiK5+Jud
MjOo3wpxD8NEBrKy2OCxhCOlb6Rgyz7gRRzus0KmOQnZdzSTvE2RvwE0gtXh4Eu/
D8Lp20KwQwQNAvrFW70o7/9jOKz3/Pe2GIpKdv9qc2jFIm7yV8tPvVLR1XZbCkfx
kBny3TRwWu6+3ay1vp1V//q30ggSoGRopzDQcs17wkFpI313WxM4CV2x032WGLQh
EPUXSyAkue+LjQRkDCKP4Q1+iYc8NClE8R0TwGpFyoIA9qg4hsaVSSRRxyGc5wTH
O/JF033hogkCWUabxeOqZUvhX5DWxuGeK7PbNqJq67xIma2kq1PxG6+YhzR+tZaV
Tpev/EO6RQTElt5O97mEBfq3jcSrVvFP4JHcOMYe5XW13GB8tzUglNtCdAiKI4Uy
Im2zX25wrUybN1CIR7XMfgZMwvTlGhl52amY2CfH0W1g+VkzSriZG5JsMOQxQ40o
ZrZc3uQOYqbQvUQRwait9kzPG1j6FEkOYy09VLYB+Ile+E76pzFURx5EhAfBeFWt
2tGe+bYQwbmZE0sydUwUo6JeMnbcGZp3EnP/2XlDwHQEtOw80d9jsYmSfH75seaO
a5KnXzxLf1QHB9c+YhvcDRtwv8UbKbrtBYRudxfXnNa/cU7zzZbLiFWzFoqZ0qSG
nJKZOtBIjvjXMruGHvfICqpr+oq2gVUBfsWeV3qay+ZEDb2OMj4VNeqYwC+9qhHj
TGjVPEZLk0BTPfsRxDwik8KHYshIMJzde/aeIa7xDLVi0NckpqVcJlATQGvKQu1Q
zT7rZsOVxy3pLUpdPvaPo/ojyYmcOavDzne0F4xaJX83qDO8YG0nVPWmqJeXRGQB
vXn4FkjKae9gTghfhBQIr+OB9z2H/1qUyrfBT5eMap9eCbMK0u7qWqUwow0Elhyj
zUMlSx4iIkxALbdnBhjOg7Bqe/LqzK3SpXGbUTe4KoSSo1RS+sBQ9sFkPuSrQnXe
NMEldXJ0JXdxMRwBPDEQ+5T/TcBTbSgLkGdg50lzi/r4/trZfg/0loSpfW4zO1Jc
9CxVvqRyeU2ayGfWYb6K6Tuksmnr4NO5ZmqVRMsJYTb2cnHm4HyKMjjgSLVZzSyB
zWpOgr1ip67VVL0suiPcxabwUeSQliC1LiBqnZB+H2KTM7H4Z5BwyFzcr633hbEd
/6N2YEQ3PU058u95WiwMf/mhCIzp503hDUM5ugg2Fb9uvSq8XYU8Vfg4M33zLLBV
9AJHCnwISeg+ikWpY49ZzrUahIm/jBueWQ/i7QPkwgGt9dBYPLCn/OCF9dQ/QCLs
zQbZ5XraFNatbkw+kZL//4HnYNg/aBPDowedHRhCGwKVU/tnogwoji7J8NyJy2Ui
2p1jSsuWyufkRZRwHW7ifeJHozfYlcICISgA9pMJOOnCBV55IJYtyZF3iaNxYT+z
7v+0uiJNPC5kwhy1nMzvpWQ8thU8IHQG1/D2Mc/EoLtYBTtg36S4EtJI5g+cBUWF
PYgjTO8Pf2hSPegiyUW8sf9aG33fJlDHR/yhoiemzpZsmH0x9UhCoMszIgd/dZp1
y9pygXbkW91Zmcl24kBvTGKcdbYhH2dY2eH7Kt73YGTv9n9FIr6V1RhxNWnfWBot
Ric9hRmarhFJZg1WGjG6sgRSI5aRMUNe/h7ADlTwdmfZ786ZSjcH0a3/yqRL/kPb
Hgmd7dPr1Wl3wG8Mbq0WsJKxI3qSswDP/OxC6tlF6qm5yt8LtmpT1SJVevWFjR5w
8tCldPxxEe+Ir+iBzqeR7mYa0slICXodv9HSvVufOCO1SUntz4+VFbjpTrVOwTUF
SUWJdq3wn5rgLG/640wXq1+ej2+CcZgn+6lYAqdFjXKQ9qC5Fp12InQme9hGKycX
14b8x9J87JngxFtvIUxsOqaAB2Im/7sRNO3VJPjlyi9cp2DUGC2uF+JoIOmbGCcy
rLY4o4z5pt9lNnM5geo1O8JTUE0RCTpuzlHmKbe4RhqV0Dcn46M+OQyaxcdDYlRO
jEWWA5YNDG5dsA3PmGbdsHmKRt/yP2HlHsj5Pz6kqwDojIuu9/XGAhNLcOc1uEUf
oxFHeFk+OiCFx3BvII1PQ44B6ZcwC4dQ/X1r+NipkagxNsam0ER+pYZcXPMgN8+G
X8jJD+Dwzh9U5h9hXShZNZifJwQLFJyInKtddX8dmPKecyf7SMtcoQC37nbw4muA
ckuaXKiWAM1GcUCf8EjTJjYB5EaD1hyDb06qvy5A4Jmbmnfebs/y5qQRGi3hmw3N
rqDoQDvzez8BS6rwuiB7qUPTFsR9e1b2MZz7kAvwoxU+j4/Kxy5NIy2DS3WDH9k6
oc3PT2fwTe9PP/SrAs7DQq/MFy0JV/xwWVKgSDxj1/rAdBdjrpwdfrgeETviXBOV
d7PYTT/TN+iNQ4QG1Ob0V/feEJoO8dMcC+SzjRaL+xLMO2jvjLyx5qjgmBM+JcX6
CgOfSRoPAzlEimNhba0Sk+Skwge5OLBmF2uCEbvtkNADoSbxjsJyWsrPzeuxFcSs
xDrKK5nsbAZfwAj1F+WzoT+bdu9DJIm7LU4sIUeNsvccouXat+5nUPnjdB+3JDFi
5mmdDrsTzbMS60IzhkjJ0SY3Hdq2BVNwmpNm+PWGYbOTGo1L8yAUINoRvFLeYd+L
S2VTlu6/4w2Y6Vp0YRSooKwZFWeUg7eegi7L0YjHiGj4z1fME0LizB11mxuC/4v1
4hhn9ZfU7AEp1jfiP1P9+EVC7KVTgWLRO8CG8U6dMqwPTF1zl2+kWHrMELH5jV2C
7ptdIOW9PROLVWhfYtWTzWKIrE6PMxFUJViigDxiXU/iI5ZlkToFDFhzb8Kz+Y+C
JLD5tK4mo5VkGyM5M2CFDGfbQi9fZLWvrX1dp2lFFAAO668FZQFX4cFDDGtVAxnT
3zlicIBcWWiCVpdJeNvBcVG+IEUkJinoltUgL6frbUmpJXc8en2gfLstx/Gm6TuX
4q4TbMvoX5uE9k4ZknBMJcosAf+BIQ7YEuN2VWpkiH/CL5S668rY01nw0bmYvL60
kAIag+N0nbWc01wIJYpBMJkG7et6twb+9ZfHdaWQPiIct21ydLvh7wkssMIDst48
T8choQmNXEY9duuUlwLw47eIsAlmDNFFRrxKxhgFkCqXnw9zM0FsyELtFwBD+hgE
eY8u/fcTLpZdOXar4fnLcqcYakAlc1LMqli1hJmU8ZIfo2FPowCf5XWyYAJ9wxzW
QZ56BO+BrPd0RZUMZXC4jbHWgpr/TwitjRwFRh6JexN/BVYJxtf3In+/M2KD59gr
AppLLeUD4xkvDi1h0Ba1n5NnmE7+JbsT4CZqX/qzn9DqWks8Z32yPoEQN7VCZicK
A1ulUHJ+F5dlLeLQ+TgPC2r3Fm4sJ5HZkmdQlNnG3GR9hcjM2Oa5GerDArW0ASLR
kjFgNGVh9vX/c164YEeaALcTGfHRL4qcWpzgIfbZ/mII/asxQKWhMjqdFxN9Q2Be
VM1edB7lTRw4EXPfTSgY83iXPsoIRAEcIQ1W8ATgkoGV+1y2uadXV/40/BVcpgcf
KYbyYGrI7HRb4F+W+wCrSEveEwhwkkDd3iSMgbJ4Uxe6IEiVavpANVxYZ3yTCci+
+orKKiBzBI8F3akgWQW9lbUYAHyhoa5mL9zIo2Z92ptbA79e2Q5J55vdGeKAKbgz
BxZCoDiOEspgMbxNJaGzcA0J9Wz0DEYHSe6k+gUhV4bA3mH3uNXimwKypmbnMt+q
FZ659KJiYEvzcPK5TDJwMr4EtkI7jBNCOeWpDGxevF2Qol5wDj2ATS8LlaMPhVFK
JivXXWuoKtgUf1a64Nfps3V39/D0by9M9a+Px0RU6x+/CaZbQ/udsENQwtOJAQLA
1t/dxW8KQO5nVN/ZPRJLxJgWKfdYAjjHJCgG4VZ6vuynRUbgxvvv0t6Ufg84DQ+6
lgn8YZpdgnNMjLEhwElCImiPTt8g9dnRE/V5Cq0oBdOxryrfSQsQts3j5eCed9QU
uycWYZL+neIGirPH2ccV8BjdPDifsbnAHRc0rN6jbey039+gVx0ASgj7o0g7nvkm
4sydbJH3DUO/iAKVvvSPTq7LmkziMPqyDDx++x7LhI/zyZV6byli4OOqNR8ngC4/
OoQfxt4G8P6XgMNOH8KrLI9qVuRhPx2BluBrF4sGILw34GpcsknuZZBs3g6Nd7P2
KAjPqEomf3MwZYw4V3QhlqLx6fN223mk903JmHf6NwwIMgbCdXA8FdrhaeEbZRsD
YyPSHR/lnVWNFDxGAn4KlOZxFSPnwLPIBCMx4mrGX113A/m3lcItab4uNhqhzZz/
q78VLUQ85qH0LRDc9Mq0iTXCbLqpSXanc3r7+HaKOKxiT9c7LibG3+cHRuD3A/RC
sJh9UuwYfaijpkIZng1A9cFTws/pXs7AHONgJiYmt9DiKwlXhagZ7Oq1bOspkMp5
6IcM/KK9/tn1+21IY0HmXf4RIzmWL858jRAal8GedL0ldoHEK5fbPqCc8kOiaqeF
Ia8zbb7IPbn2UQJlP3Ty4LkGkECPCVI/piPPDuOvOTNij/yn4Y/ryRXyJ1tbu9GK
9FKS4Q+rzhyBv8qMixG3SXLPwDQC6p3yZ6E+/q11Vb6Mw7isrXeaqxGESCzfg8ux
roXBZR9zY0KZsHsBVjrhhF4vu5YwrutV/kB88WCqOZBAuQuiPP1QFoEIvu7msEkV
OGxaKf2Ew4LSPL5Vb3SDjaVHGG6L/On1caB32IjEPHj4FPAb2TV/uE5t800i0UIy
PXGI5+1HuOK+1Zp86tv+AJC9KKN3MC4WOg58TyAp4i5rk/dnDR96c0XlC7Tp1X5H
YSosC8cRDaQK1Z/cnCZd2JVSp4++GHixK17P3xRnTnQWUEuOoQmvy1tSVjeEk7OZ
XaOixcpBMmA0hLu3PFaiaOtzAtsNQzlP7fayoCk+e3goUHYqRdM/n8/dbaD8ErOx
pEDA/o1dtbXTzmUXM49lwVPMJoVmYsxdhgXtnU04RQXAPXprpg/wjcwdviyrobIZ
xpu39MkgqqZgs8+f8ja8C6PIO0/oCgW7uuEHzYEz8iPpyPNSqnYELmb/YGfRSiSQ
39X4xUbqs55KEAUSab7ORNv5jUinHFgPh5eaXjWzdxYcelguMCcLWQZNjmnkDDTB
HpxO6hol9zaYKnXZnG7e61XZHDSqHFeT/nP+sxB2EmgM8LcNWiJ0rjnn0Q6jXXzL
4c2YPgr2wEC0CgzcLo4R5xbgbm/v92NZ6XueBA06VmQSAFKOWZpxaZsGeRvoBfF1
fgGCjl7DUsACM09DlAXjO/E8xJvNJpYmMDHBKCrokKOj0jBPdIpuFdlTGblSxRmT
AvZHslzSluW1xrxng4novxIpqNYfqruWOeXjlC6Ycni1J15Zs5iXRvUYI5p23vX9
6bmRy7LrZMGV+Z6C6boBFt8an0Cw69tNnKx+M4JP0j5drTcd+3ExYmwcDS0zhYHA
SPUP4B56CSP/IRy/QpNG1BPaGsuXYUTgCMIgrodn5XRqEowt9CC4B/9knig+wNtn
nOkWaE6DaHD4u9GyBR/7mW7SpYX2z8EyFJgUmx7QH9+Ih7rkHp8CFXecveEXZbwu
b6APJGMLoZYS10liGX0I/PZ7cLakLqlt3Fu2x6yViIgFlxe5iyBPttJUo0yoNr3Z
rarsj7DEysnek7DdMaZ3pr/E1/AOuqTsBM9pdjY9Y++8ThIMTgvfx1JYAKz9LCoL
FUkMdn+YoLIWCyEm2cQI/RsMQeECPkbOA1/xpaAZ/QPOxD7wnRP+CG/prWqz8AeY
bdqyDqcVRUVRuI8RAxvIUgdQbtOHSAXR7P6e8nsemGOz/Pz3EX4f/qSi6FV1lv7r
bOyyWf7zlejbYM+sTtZENuQx+HYJfhUvMMGrKIj1a0vv44gIwMMAtLwO3cpqOm/H
Tr1C2R+rg3Wn+esUSLnRPjMf3W7ip0IPLJjd2noCGdanUVEO+HTnrD1bDEyB5byP
jPElTWZ2m/VLVEHi2O2rJ5vLTqubVkP0WOllyM5rWkQ+Jr5Zio//MSkBY/w2x4GE
8q7aL/cu1jwjVq/coLWCVpq+I2FeQPTC/vEEnGfpFsCWQ0jxkllRgpBnr94/QMGC
Py0Nfmetfm+zdsnn7TMV7R87DPjN4nY0oQaYhtYG9jxIRWrTxaroKij2YDsrA4En
uPU3tTOG39qy+jaZntA0Eh/KT4hwV57hR0UIlG1ONRvqk+X/BbEPGbgnUKe2wjFM
7lV1h4h3l8be+RTLW4WJ8iq/N3QDOjTytyh+aKOvlTpgGvJ4YQPt6v2hpDzbrzX3
NgRe6qDFaPhJx+0UuPB6F4AfarrWtI07g4mDqnC548WeOkTyUVovsAJde6+tew6Q
0Lma+KHZ2K5Xwy9+qV1ZBp7D7hot0kAduCNWAltstvtV6Iar5WfIld5cQ5H2oBsI
VvW7TpmxKhP1GkpFHOnJYkLL7l412q7tvD26R3UtqTVT9RZSp3Pykn31u5TLQj0e
iVa2i/8iYS+q8DHIAE7900u9zq7g7uiWeaCq5Y0Yg8D8L957MGcL+Rnsi6iiMCYJ
AMtnBa8tql73o2mCC+sIEFX6yzpbmZOCMkZIgch7IDlpggQXsuyV8ig4R5w/dAVT
W1T6ijQykuUghPCpdDCGCcdus/PM1EQ/ox5cdtviSkUlgInyg+AsmrW4XssDfSAL
G8EBcahzvQDJHu45TCg/zxZ2bOLiCJ4NJ+tHPSIt5Dwo4DMQ8ldsU9CUHZ5vU0eI
F0NyemLTtVkGMiiEhPfjg/P2msTwTj49xCHqgoHVnI4kztp8N0j6jZ8djC/rtzdp
45YRw0LXkzQFdcmb3E0Pq7eJ/AXZlOuijbDCskNp6gxPhIIyqafs0yMj4V+KKVIf
2tp0yeJ45Wn0hUpzGUasp5gUKpGBhIZ4TrHlSgIq3vewAgdiTQHiUm23r1SgVhPp
Q4Q1r02qNh4+VFe/5Z8DeM7CP/OzCvWgFRFeWzGIv57YBiNUL4DRbvbRWy/njIP4
Sbn+kXuuMF5Edk2GKvr23CwsV/PrktHEccmn5pPo3sUlhXULME/bvPLUZVY0Uyu3
xeIq3SPOeCA4UFC8QcbsI89zknRcT/IyLEiMYARG/ErFs+uC0YenFPhmmxcnqkUR
hrvkrq9glwQKv9DYOH3GI0Ifga22AYbfYhHhmezXrlFAWJXs13Op3KMpLkoVCLlb
LZtGUO/3SSKAaQf2DL+VXlI2DhGnEvFmyB3Kio1Cm80AmLNlQmlAIplSbbaO6tUx
W5MZnPwCpKl+IgtyhN1IpEQW2W+voLLsLTwHKjp9vJ2XSQN+hVvSvYg53XC3DWNA
0MnvmZMmUmdeUelsCyR7h0vNUFLED4Ub6CHWc0KWi9asrgrtU0scCs4MdNR5cUy1
koyl/o4k9nZhCTCNENiO1zMp+u+4febbrFK8Zb4ScY7y6qbOMhW5z4Ljl/0ruOm7
L5NFDD2gizd3FAXb8Osli3p2VPXEif32v0QJnIFleP+Yf2EaO318CTzRD8y1l0Zb
c8BN1++ECFkbxeapEFEpAo32sa9WvdJvynm98L2QtdzeCuKdbJ3zcPuBZTvLqy/w
IJN0crA7iiIKxU4HXWO/LbvpRakpULgh+tqtYVDJDXJcveAKIYuEwzczteFgPm8o
XmAiIuJT8SMvcpOdX5Dvn4uNRhArfu0Hjjl1lH7eaV5epkgAMBOkdDv1/1tVuq5h
dbHbaGCxM4UMaNDj5VJA+tFfP628DWosPbqPzuyzAdQj3K2tlpcKrN5ATsbKfNLO
0piklO6N4kqpHtTuf+6sqca1kYLTfud0OAf0WC0GbeNTBlndLTifIi+18zK/wUsJ
slukO2A/ar/Bo3yleys2lXsV/1ZhDxKoE3AP7Z+wyQSqu4OMCp7MvIe8jkuRwPhX
SGuyuXcDAnFoQmZLGu8SDzEu6RBiO8hwjjGSoZDNBgERiTKuZqeydrenygXHGF+T
DgnpyY1e3xS0SKNcBb6BOEG+HKNJswE9O43uwdyzeKv/PDNkzkjS0pxPJA/+O4kA
2CBuGe+8pSb8v0BxYrjS5wvrt08jm3vbMnF7HESi7WoGlnb+ERgQg1PhcXshvZoG
geAfPfJGuU3Ema0b0PT+ec0sYpgY7AkPGZI0etyAWu5waGCh4CzTqBDP0WluEKKY
KhCBnvYSBEfokzyCkOyQJvrFCu391HpckL7jqeeJeI+oaN0HfSm5gYNzPTU8srDo
zljmbN16EpZckLN3fahtdYi40qNXltkw3FiFwdIKDPbQGtdfkcZodtlVR/eDh9nG
gQI/hg3BSwYZoBXE1BqOjryAH9b/gV6Vq/DBAoARlM69I0SFAz9LbUmCyZgbOlmr
f455VSV2QxJhYUqjOAm4D23eO9j2QXpBc0z2UUZgF9tj7fBXNlVG5nT0yl75yPOi
pNKk3IocQ49N6tff3oYYv/0Bf9l73aSkQAeggyXSLLU1viZeMJhlFCv+WozOtNPP
hcI9AeldLQA2xYLW00rYDe79+x76nvx3v8C8s1CatMJ0n2+DFDl+fy49n7pSyA7n
4ZpEkCT+28i2oe5I8vK3LsajoizFn6c4Qzs9FDKl4gah6a/vefoY7iy0TL3T/O85
VFn1m+x/NfQE4klqerljFzy8kmNYcRcvuwPFkoOcRWn5GNrNLNKRHlikY5aaDw7U
gw/LukpKZT2ASJGPY4KVS2g1YQJ5lv0MOvPW0AyuV+ac1cDHPGbv0yAnyga3M8tK
bKvxmOuQFe1yxvkjx7SFcbQAwfuNnVf5pN7Uyh/ZXtHxGc5gpbJUU4LkgYLbNtFP
GrzkVoSH91D6r3iXP3dqsBo3feT22crOdpGpMpWy7NyNKmeG3QvAfhPsRFqCpnAm
hKaC0KFr9al+8u2bNuy6A9PEArXxurGzBx1vFfF+7uE7gH7XmRLvMlMRANZNfCno
N0DteX85axEwn2V+5Pt3QP9fpGkmIB5JQ8Axjl7hdN22Cmax9f4aeJ9bWnFlo3zH
wZSNRxkAk393u3SADuTfq4Ihl3U8pE0WF2T1FPC+sdGYm5wM3bCpEpl0nl+/5G0Q
ah2/QkoXtfv2DcWSfqDIhKWz5vtgkGaIHEByicDu6pbLxAvwKgsbTPe7tAdRnuR1
rchvzzBLrGfBnl2idmrZgBcR7mcn9cQHyMVns1o0bYgTQ9CZP7005wZ/LJuzeE1N
JeYQUrcH/gJsj55No8qRpD/cMehbxFcl5MmQ7tQYOwCuAJZO0cKThWIVPu1JHMt9
mxhgZ7Axq4wePZXtRq7mmEZDzcTV5AnKrkwniS1gqsKg5yQlwNbNhQvp4xMQqN9K
JSFUDOYCy+6cA5lcpizhAqeu57AyrWdYHlG4YNq2ThJbzaTW1NqAztVJXyPKfflg
el4yOWnOFppjyrYqzu07cOf6mmBGv5/pds2sdUiKG6gSQkd+2mAVFwlzKWxdjf1z
1EGK1sdI6RHr125G6TDyhMqB+j7lboF2rFPjL7Loj5v1wXeTmHrx8J6MPS3RL6vs
yTYmro9mu473fo2MR8rlb2rO7LqoC+WbZ4s/1lA95B3EspqgVqu9ehBMqFVJCZcg
ImE6e2aZU+wKA72cqBHzlG6YGV9FM9ODG+9gysMAmsbY6wM5xSjFoom25Gmf5wSW
4XIlz/+S1is5cugtwc86bWY+L9xIy5jDiVoMTqW67tTstnhT5Siz/VLHgYLl2EZ6
01TzYgmqKveOMIfpAt5bqdGhvHwLXpE+1At3kGf+Y2Mz9/o5mfLCJ2SOoTBRMhT7
Kg03zS6DlyH8aJI12eLvHlDt3xhkQZ59h03m8Uik12I8q3nU1GM7cUyOLguKVzRX
TWhS5brbCrzq/HI8ArDUOEsRB/QopCp9T4zwjNBzOEFImcsGNlEGi4a82vuVJ2eF
njrYgXPzIQY/rT14TVixR+csJnYTXm7E3/hatJfiq19uA3TzzGJxh3XR33T1d/Ts
gSh92H2ZGRoAy5QqjyrnSHdgpkjSUahyCvsVj5w2SjQrIBfckBUzo3Xg9bdl8nd6
h5cK+dbWCFx+t2Xl62LDuhxSVyL+7aihO1VBrT6k9nPNCEG4TCDU1adVpjDs7NOi
oBevsleI6KBPGwVdCqBf58+QogLGRfbDLUhazm+tTMgNMx9c7kTmuX1Etx+7HTm6
8BSW9dQhxbFei3X1qaib3jSnjv6+eYgyBV8KoylkSSvg8AbPvyRUol520c1DBAVe
0XSxOuSKNaUkZAQbShHdGkqTSaa5NnNg+luN5TBlQyi+qsklelFt9vAA8mYXA4ue
4M579pnZhPF3tv6pEeZGQFSm8zJBEj76YMZTpEN37lJV5OLMp4hnGa9nutCGJQNP
Gas3+cmfOhxixgnO7NaKzQ1d+Rg016dU07EInLGF86vLxlkq8iFuZAKNZPs6bwoZ
Zc+0V/1KXfiTTrLvEWKyUm8uRypDkWASXMj9Yk1lU855CnqaWtRqdH8iETYPpBQE
Gy+5nBfEjHoq4rtbIisOj315Zi5VKCcng+NImfTxE1U3gomlpFkl0hZ/I2Ez8zSC
ompSYMxN6S7RLDRuMme+gM//Okfy5rgvRNEYPEB4HafvNnd/bh4gPTl7bfdWrNTG
ogL98N/0B8Dk/s5aZD6jwMjoRZJjdQFh9UR/D3XIPIeT9x8N4kO6lGTASW1xZTTj
9EOLi9fNRA/Z2xZeHkmo63mnoV+EvpSla1SDFNBRkajxdXTAFiZQk1z0IR2SFSOx
GiMJR3ZlVBpCGsL+uIbXognYIaJKfwMhcZjkwFHE2DorEfvO3116vqp5/g9hf8yu
7uCPL2jYL7tmilZdX1taHvhEWP3wO9ZIZTHcM622C7FZH1Iu6CsxrU5pzQShZ0wb
AYRBIgg500H7WR2as0sVr3lqo2aysIiZghK8Un3lrYkafhEKht/6VMY+LIZiiBWq
5q8QMC/41ts4t4VdSpk6wlRr4exOf2JVXPGgpYlMwjLWc4yKSAGnMN2vdqT+FuPj
gPYYgqrOT6nWRI2tnj7PpRZW1CO3Ev4CZRab0kdj6taxab4k6G+70TA2o8ainaie
FisncPiVpDHKZsjogB2JYvd0NfjM7Uk0znv2o+nKVpCWm2/xbDkmg05590EsQbNt
wesVA7H3T3lsPo5o6UReFPetJ/8mhFTy/ZqJOKVtvXLo9/c3c7Rf1XyoG2lJN+FP
JzPN8FWKYIVfl9sri1AB7yduBf6IT7j05zwCzdV8x9vV2ZmdUWKQebRqewdkmfh0
aRIFluoxIi6fp+1oJ3kaqYCyylTmkgLeMkTZoYtIvMUBJ+QHEqxju+yQVIzlFRLW
mZ/cIdpDwxLwOUdQI9Htw/U7OU9kWYC8mh/DpR6scJGSRnEqysE30DfpcJ+D/X1L
QEfIRZxWj0CH/6uHmvuXBXgQA0E49bkiKob0fxHXh3wr7/sC9iBd/VWrV8/L4ZjF
j+JM+Okoo9NGWQPBNx9IgyRGS73eOB6KgMDH0e3UF4JevaCHmci4efntoFBIMbuc
KfkSSNzaMjkTUEYsLmGUPR8SyyAqwbl2p1+YD9ga8xfZyORGexqEhW6K39KoAGOv
LuDVb4IJICSbWSr8vN/YfY8Uu0Qa5ZjMqYlMfzo091QwlyEJLAD5Ij0O6s4QpUgf
CGEtnY1eBV+l5kD0rz/zp1/bE6WUC1YpoG3T03dmG1QhLuDsm4kc73ptTe534F6C
YpviGSMScgruWUabKwQ27p5xFJv+8MKs1K73XP8a+XM5iGJCTKCmWifsruWrlsBb
tYe94qD6G5zieox5uwTOPDUkXaHm6/NJFGNR5zvb2CAsZzXjLRZhqSC8Jpjl8K4g
6tdTtWU894JUkz9zE+lA3QfcUBU61cVTLzEoZ4vgAUxshL4KVJHF38d0gu+4tE1H
onImJLeaeqnNjjuR5Px0V/Pc7sf5w8nibBFek9Y2TSLRK6eGQmist9ixrvftuVnW
1zRbiBts7Mg7FghE31TQHUINnqpByHzKWS6JxnPQrndHORC6h7wnQ7LZVxGcGe0d
shFkMoGbI0GaosB2veeHgCL/849RIeUCe2zQq5OQixy0VzXk66lSf++FQ1d4vjwb
0dlrN7alJYNeTHZS62LROTeAaOm4ba1UEY5CdKrXSkgJm53yLD3WVsXEe7Wuk02w
bnrR7WxWP86lt+1+sORSMLWD6T7pjWcMem/DRjDQcwQqpB6JbGAM9dhMIxzYVKLT
iwpWctXO8WJMKSiVfUs9N7DmEv6UhxlvwqMfiPtASnQYwyfP+iQw7V3Y+ZQXy3/w
BmO5KMhtYKW8NBd52COHqhgu8ebXJd1GQYgrqE77/bHGxgy3GHk5zcr7sp5KUrY6
b8H3G7d1twKCKmubRwrcyKPdJ0b3SjRhARC55mVqNH0DMzWaLs93eEENnx9NYCg6
9d3z6OUx3XvmQrb7bIuyVmox/c0811OvRGDugiOv6zdfDjuwABUUWmv140C2SuOH
IsrzITk+/JxhtL1aCt11pRWEfDKjHCHiI2JNMepwpeRFhoejvqGYdBrK6cBIIJF5
P+qs3ShchIswT32wPBmWbM9ukqxtCH58hINvkgEghVjOVoKjrr1ThwjRn67xgmCZ
jNtQXRkcDKW777ORDgU2CXrKEPYXWKh+PRxWLncS6pzzZRJTmcY5gx9ma7P9psMW
7B+OxPrnV2Rkp/QhdE0yPD6iRmO8q7Zavqhx/oOEzcyCFW5DO2jzL71Z6Xo5HGWw
R/DB/izVXucx777gu4BGZe4yVgU0iVpclF1t+1xhZrIJ+Jgl0C4arbZnULz9R6Mu
LGNPzFymSSXErZqUQJ7yCK8MttGvgFWizl5ipYpG1WAvjqQ5rWKa5yzDtqf1RyfN
bXLiLgsjJay8rZ1EwU7833sRjCna59TCOYwtANWx14+8W8auM+Ow4F6zFl3mMLqm
86Mtfnix85beQHmkEVKl9jUsU7e+4Jdg0f3VBOzAcM17/SY/4jh90jzyB00yUPxs
D1OO2Nu8xvKu0cfqJTXO2fDXnSAwV75dqM1M2w6Ay99t0WMqfHINq2Ocv2o+8Wka
S5wRrgJIo1vcesncUm+J9iOTLR9LNMhHwbPVXMSRqW9yLBtvicUac4adLwaGiYji
fjV/PQ7hywKHUpZXR1Y8H5n0eWwp89QEdFiJklIRhtvX721cFMD62FoUFXsmF4gB
nLPnSJq0cqCdvgBoGAf66q1pFENq6zcabwRo+7jVa9iyZwzBsHFvp7w93ebFrVnZ
r8wIl/oazF5nqD8AvrSLX4A4gxM2OuzPohg4M3uy8f0E95t9QFzBu/qkdMs9TTKV
lh+1sXzHw3LmqoRMZQBQMEcfRCrdWNLb1inObC1Rk46eTscPWZ0kyItCqMxCk8E1
cDPCTzyklyicAyjfB0LFHtRXNAsBu3Ncl5tx4eseMm+89QhiHNURWRdHRLsPEtME
Qgun4DbggBUcFOndHrLmCxHV8IVbHgUFlKdpajeaYrOx3ik6SSwoBX1oPCdD7Sns
NA/rTAh8w9y/QaMVp70fiv0ShL/6sfyrtV3GSpprQWsfg3gzLBasMknDj9TFEwZA
WeWSa4wwpJruaY0Z30Io9kyN/VrbBi3YELao5WkH+vRGkwbFGvr9OGc8CTbGhb6B
1+dCywzdG0X4h6C7b1078V7Jr85fFXpU2A05+86Ru7glV4eo3klnGYxvwMwTUDCX
d0uNJKXnm4VJHMWzhVoGtdr2qm5fL5MmyRU//GQK1b0jccvTZneTB97qurqkdeSm
8M7h8lv+cGf7oo4R6D4gnvLynuuMEE2+KHjAJSqy+A4W7Bp9dfFFofqtbIn1i3G7
r+wjS92BNQtfPzm3utG24goZx5Tw8TzFv2jOpgessXXCtTvT1a916Wtzc0WmgUYY
hQK2rwxtHKypVL23SRduWN5959tMeg3ECeKvE2N66XaAU7AnqkG9/hbCR5QJlw0a
70qfsN8FDIS1YcSCOzIATrwQjxSdtNDFuNtFWfYZi7gLuogfNws3XEHSr8kU+woK
24FxDHWJGGvimEpFt69q7TEToPdvi/ZS/qg0BrkHGrYjCI6LI6pf+9GpjxO0tt1G
f9Fo3l29K+Fk0Z0SxCJokNKsutEyyUwR9yRa5SR09a77Dp8tB9jz5JXYmM7aXSGA
fLpp6uTpJBrIlaI08waW3XX6UdLvUoBmHOp9xA252SpL9B2oDVLEwPDQMIVqeQ4Q
QdFIXDkZRfy4qnn/sJ32sfmx+l0LNRA4YiWpWpkMuWuSLZAyBkEELZVxWfx7nOQw
SFsViO1DPb6eqGDbUm5G/h2OleytT6PoX8esPEJz92E7qwz3SzkRJ0ypxBUCLb48
Jk3jRlT0uQoMRWchCIMm4N9SEsPx7z/gWasPFWspopKXoNAq2sdNeBt6uh6zVmd+
fw32te48C3RRn6IlpfxHQ6YlFhV99auoILIMDGs3YcjLGYd9SO4HcfYaDMpgEEjc
g+ZHyIEF26xXDxke0tHoG3AF0rItJhf20WEISbKQF98Fl6NOs4D9kDAp7m0UUIXc
41i3aurYwG6ryWRMfmN8FEWFYYuC2Kuf+oM99uhZjSQVO4rpIwwbQSwnJfLPuMDx
Nc1os4jGOg84Z6xy+xZ0FInLJ6rpw1vGFwbH408+cQ0mnYqN5hVyFJIdrvR4J1+B
gYRopLokNg3fGCn60lTzW/7uNIwnaEz1XNTnm6BHw62n8q+vJQzX4O6v+21hhPlQ
C6nDJJ7lwKrsExoHawa+59O71hqD2sO65jU55+cxm8P6j/ZIa4z/0gB/dQAJucPd
S6RhUvZCOePpN0DS444CpqZixdI/RU/Q0ZomSLe3G6VY0nP2l5vYym6dmv4zYi+5
IoB5P6dX0DE/oG3Wi96y1QghOGvb1WUx5P4g2xrx8cP2uXDLdk46qU9CrGPAfBrC
AMgfZ0wcy6rzSUZtpHPRWkVbA9XoFtS+oq/bQx8xOK5z8MEA3OcYoa40xDHhPNuv
gH+Xusi/sVdTP//WPcCfNsajA5ww5nuEoAgU5Q9DATBwbNG7V6lwyl+XGO21v1tV
a5r7mYYF658Rb/pCQrlyXbDNgAtDRCNxLhSXzriDXq5oHVsymk5zeVPRvVKGgJ+8
Kk80xNQ3Grrgo43jkhhsacROousYxu+HEhIt/oy1jlAaglf/neEGKTEex7ZP9yek
eSvW6XCzpEir+S+l19KcSjkHSF/ASXimvOSCnFyNjAneHa10EYc4BXlwu5jLP5Tk
66ho0ygVrB2VQLmepLmKPMbuVkjxcGcdcCgBSfWJWHgdqbhT1NDEfjvHgnIa199W
WW6b0qU4nFe/+cBHXkukEi4IBFYfDU9GW8RQqTxaqdWoOXah3GByHKROkUgUWAaG
JHSIljFQ01PvkTEwifmgTASN0mzaTzvrQvA9lIUY4yNcyAx58Bv4pgkzDBzLyYWy
oF+9z3Agof01nsXR97xHkx0wabe8HuQzJLSKXgX8vbabO/iNAIQjsVicdnrWFSoR
t1NMugZgtV3H8U9akpfOm342nP5GRZdUVwWOJCo/8R/A84EbKMPUkl8G3Yr9Z/4R
eh6zFvP5DCp7xkePBhO2tI9RegxsYska7iO4LxNi8WYDtRaeaA+ZBH1m8XhNCPLm
Tk3pCW2c/3r3nSXITiadNTCUsCiq47byv/QmaPvsH+jui+gwyf3Q8ywJaWWIS5zw
1Glyw7AQdN79ZdazkJW4GlfI4/p0xO3k9v2v3mHDVedUJr7t8ANiowZ4wCJeyypI
stDnu6Mhi1upJRVu7OvRmWzhwNZMEEBK3j9uKiauhxtw1yTvbvHagjvmtLS/51qp
3HIodrSfgfLwN4rCdcsr3oXfgnAu9prCZvuhuR+GEGsB2xm7fYu0ob9+EPZgIzeg
XBjazoRkXOq6af4rx6QQ61GrV9a7GhFrmT4gVOQ081X9RoaAzX8Abv+xdVHj7IgL
Wd2vEqaQwAO5FQqfksnK+2NdSyeCzXSl2f6CJbTZuday8LtKyc9hube2VPWtnQzZ
Jf1Er/F4XqFIv77tf2MyfM5atgQRzO+ziZb8JZi4mLcQjxUVR9xbluGoMe+1XLdA
P6sxdIqZaALJ0L2fs90IPEPXSZEjzqyxTROcRZiLP+d3qeQ5xi55RRqHq6fiSaYu
zLY6IkIo5vO+UsdjIgSEew7vEHgbDWRsBE86+pjm2F8CmOOgv/X2b4/s5UpxCul+
3pCUHOid9AkS++EyVrxT4wc1dSvi6mMoO7KF2/QwWjWpLUyHhcla+dhDHcWAns6l
8/Po9kPTFnKFwRUwlV4Fe4FPWUm6urzbaX8hTHKkncQylr13CIbfUGEGTaUoMz2W
CAVwJM8LwLMVsM60g+9Lm8dKfzAGJTqCzwv+LKq5KJgrqyH2hCjOP2Y7Vvodm8g9
lwvXs2HXuMzYpw2aRApRsDyEX9zVmDqmS+aIg6QzewYXiRyb5BnHbZOY+d+xOxHt
3naonZOywFD11gzMca6vhl5uLADYNTY+EjZ8u9k8DEpFg+Fg4DDsJjvLIBwdk7vN
VjfPF9U40LvmsHmkCTQInN8G45EwRTSvcwhp4YpmujEHOhqXVJmNWkVlUij/sKVV
JNf9LvH5bJzoZXEBfqWKTLpYkUKG4JsF2biPccGrsGceRAqQoHZ5zsy07XyHT0be
87MbhCTMdF3jsc/C2hp7z8CO/mMINtH3GPy7+rNA2iDBxJrvaF4jeOwnx1WzGrVU
sY9Y9klMcgAiw23AgwDt9++0CPtUuBYaCvgGdR8P1Fnvc4GpCBUxxLBCz7dUatXD
0FMUz1kojKyTr7l9KNFZXKXvVD8AfwkdnC32RoxuK0OIwCRKOTn3296gZPQWkea9
WMqEKiBQJoWqvfQQ0yQI5i2vujKoNLlmwBGkHWi1T2cVewmOnrHHJkFPAmeWjCcq
bIx/NDF5BjlIcA0dWjBlsxmQemfgnwhxf/w7dvBpRrhDNv97mZ/6FPpXRKH5eYP5
nDvWb/lqhfWje+B+6e5twAWY2WvCzYRy38tIWfWnRDlvYuK7EZg0GB+lhWC6Ahtb
uxkLZlmdXRZ18h2ssU5ap5Aprhw8xHe7pSLiUxRdyYp+7Ioja+dQSDGgkS6zZWIB
2bkM7L/wxspOLCOXNWi/yRB0FVkqI66spK7MZX9G26TEhh2C3IDl5P1DtWmk0R7U
0h7Gya0dEbhgvEtnfNi/NXW9FMaswLaJMqKAPoauv6RLl2ZxlbmTGLhL5SHO9UGs
6hjZ43JeXPBooDFm52yNuNWD9OFsxK4TiMIjw52s/dJru4pRQLj2i03nXGCIsFIv
YprbVPVRdiqQPjFxXdCMikox6brAQDTaafK1V/fnsEgK/ZQ+t4vFGM0q72Ce8CcN
XAMqHJuifmXDg3689K1JViQYplNZNw5IcUBCEvjQ3cElcc5Mhv+iIwuR5UJUIGar
VsrK6AXbC3rhZ+5D2zgqluWr7kGhDw61otmm6GxNVx0pYx32jEEtEY4SxbiH6fy1
IGVeoDHryL3U/cCctW5Tt8bw6PjNgGMPWKVu7mNPFEW4WIROpKYbdqY3hJXrMkI2
feMdxm1TeKx0OC0Yn+Xu6ExCtk1O7CNXJAazYRza5twp12tULZggBtzkYB3G9Da9
J/B+6hvf0bVU0MzvL4KCiUfor8C3Ybmi81Jd1ylXAJ4I21Js6t3gy0cH6yQvCSQo
qSbxI0IInqRFHinx/zFQHZVpJemDKpBTkYJ3aWyEC/UKJaWcz9AV975dkwUxlxJs
iy65VzYDGzm+hivzovaICehzoPKJuI0EIIod3EgL4pUmTEv6ICSgCDNosJ3LgIbm
5RzG8KdaVn0fYKhxCSZB8tR2GsgDYwYzXxX5RpdYZPH2WevsoTn0kBidYilUGv7I
KGoTmMK62u+ja6qQnh0ST8d2yOU/jSW7lBmkFqnCsAYUXgvP1v5sPsAURyaHVADy
IvV1kK8hcOgiYcgiPJ6frGeuS5kiP66tMb/DUSQ6DTL56SYz/eMdpEwwRBsspw7M
Oda3lKWxVND6VqU86aMrMYYwxvPA1V20pTVqNivEV3M31FDAHhvoyEQ6wiFXF9W4
MOmX5d+bBEZMi4Fsjn54sMw9Sev0oRYAHdwLKDcKJUYssp8+52OoFqLsf5mBi2NW
cIS0xx4Ddosu1MCaynm64WyjkVleocfG+4kxxOiA3pv8dEWVc6WAvY4Y8wfZg6fg
jHiVze75jPivHYRI227AoY1oHdMvpZU3tKupDMGKjXaeKaRQc4nGhMXPIsti0j7P
UNsjdJ3IAQU2cwHHZL54pvW9xAaeP9OjYiZ9M0m8FxTsg2VZZDUszdJFoJrbdDhH
TREIwix9lmdqs3w9KpojaObCLxGxTF7DFO4DuHFWH18ifPolk+DfCKW7Hhu0eGS5
AlwBJKuqxDOIKr4KLP53KoHC02+IPFy5QIo015INmwOatxPhLjwjqCuvfreOH+yt
6pPlAJZPV+HauWu1wr78m3l7jA9bF4h0IDsIdFL7aih/BPi25s/WgFirsp5S3e4r
5OBImyHC4MtU3FCNRSpQ+hQHDWK9v1OwurzaZ9oMD2kkcuLoJTFM+kSVhaFujfvO
1FAwAbJdC5N1y9HFOAJd3+TCZKgVT22sZ6VTEYNqTLhYfaOHMGv2PTUQ4Tmz0IWH
OJp69HVBn4dpNNZRQ5ehLIYlvIuYQ2X002NOQHtSiXeV1NL2YAl1evpUZjJA1uMn
oq7hA/QdYnY+C6DP05pTyU5914iT6kG8tO8jf0lkkSYvKsqZmTpZ7LWalkPmQ1vT
f8n2WkdzGU+jEgNhRPDdCm2hdGNnJOyaNkcyhqr8n9pP75C5hRSWX242Pj1Mo3KK
0eFLkpJsok+Nz2LP1ZKRHqD45ArvUMHWFBKg//cHcAZbTj38awwHKS7fYzhVqLJg
6ly+IjKHIFQUinr59uZfjL71Ay5PwXoYojJAhoKmRWUdVnAsLLLSwRgeRA6gZ8uP
aoblUoDK4y9q1aGU58wgx2KHHAhTCGUcD6pIc+5qX9cnjlmUWRNHbp7CuDEPAEpI
QuiqnysaNBx5vKIzWNXWCy0EkHA/kWpNHbTGuO/EIywpUNQFlor05RFOzKtfSSoV
N3DNtkherV+ecpWbxeR9g9oD2lTUYlL7GIeirYvTggzNGgoChIsPHM+gvIZB58bc
Z7cavfbQZR4sPEURtJB0crEqC396dzKk8oGG6bma730h7A7IuXxEyL7z09o4nU17
hSp+Np1twLwrk5VGCeHcs/aewrPn8j/LUXqkht4icILGZRXt4BPc51i2BcHLg55d
omXZmCH652/VCZtJ7XXKLxri4Dr4yfNPVSMsoyiHq5rgVNck9YBCkkRpj9Z++sWr
8WboadvcPFSGAIXip+7wmYKO6EulNNrRhDo41qNzsOAnccIRcZsHt6g8ERI7T/on
YPr8+0VMSBXLjBqIZLR0W2QxrLtbR6vM1d+hCMaGa70APswhkyOXIle4oPv9BOuI
lHNPsy3MuC8jreeh5mUO4c+157gAfjQLc1/lPbSdlIjeWVldl/Kj69cn33EiOZ79
B16n/GjVE1EjTqego7LHEs0oHncLU6CChNwp+d/XEx9zGbNGxbQlAwMbaoLZqTu0
8kkIeD86sg7zGgphVTjb2YfkS9zaogCamXp6eweXvf8tF8FIDJwMsXpbhTCgrElA
PhsT0ZTw2uv1sDsrEKUMudp2zSFm24q7fmblLfUTazu1LB6SOhhqgdUnymvbMQWo
OeiwgqpD8sFOntiqIXtyGg/AUdac9cATTKS/Mu8lnfq2RmINQ48zi3VQQZyOlL/q
jOiRFJE4yD01nI/bt38cVJ8Abdtr1aMtS8ldIltOM/3SfOyRHKuCnncZz+yTX3hB
jPItrbjcHq6Jb/vsBMV2tasWwY9UOgavV5vvbp6KzCPUKOVaRjnOtQBPMZI7A35L
CKVMcUmteXDCtwEHnm5izpVZ9QaG+ZhCy3hzMt9QuICPMHhgdpbZJlLWsbps2Cnq
+aFG9sAkAaC0Zlz1BDTELG4MnMizdW89RznyvvOwdM1VY/o2qi7s8nHWeZvJH7Su
ztej9HI6Dh9vRrhuG7Y5szQN8+or/dimbET5QzGnQAwWMAFsTk5H2mmT/4NreeCi
2cEUCxqn223Hp+J3r75NbiJAwEtW5Pf3N1hgWb+sRU2ooOj7sorAS5eWhrb0zKh9
JzHGH1Tvz6yNoBI8ipNRSTlSqN5j4FACE2UUx/CaZ9gt/svZuEAMPek/xTZcrAhq
+MlQFnOFaDuh5Dy4Rt014Pwj1P8X/lURiNJklDeEABn1L0OPMKoVACbmLDpuGk5i
8LwcBDn9K7OCKBN9dWaQrcuclLUB+Do3VtSrcIovGu6TZlZ1Mqc4foF5GbdxdKW9
/vSNQ8lDTmOotSXzsRZfXO/HEHZMVJloLWe1ORE4jKZemDn6enFB4iniE9DfK9QP
7JUZwK0HgL7pqKOcBUIlHMVYqIDoK+7kJ263ICPGX8IWH17fY01MYcyWbiD2rP5c
42ICJg9M820IPi1IHlXrgY2/WHiPXPOiAoJbukKnnNTYcBRTpGPtT4c6tdNDRNoa
bU4RG+6fBOsHOytIjRLquj/7EbmXq76tG64mUW7YWyFIsgNmdn1r1OtXdbjOuX7s
aJ9v+wugt8cRwvej0ENjmBVmwwrXBtwG1TcL3aWdKC05IzTn5ulFtqh/BJ5dHXJd
H1XR493YHbRgnCjvztqrVMJTViLKLH90ai96hYKTa1OI5/dCfLC5NvNhrk+FLQDL
LMyi9UuMw9VbyElAS8fWFibbDnUll+5VahI9/j4lwky5PpGcA2chJ1DwWioQJ1xR
olhSFvFgaDGQE/KUtk64PCNdywhsDGEO7rDkWCE5LK+oDEZMk+WXHGegg6ux/gfj
jdIKcgpUW/l9F8QvaYchxSl0WfYgQj2JxVLJNIdCS/R3IiRDamFh7rZmb5IOI3AA
PkYYvx2C/ooVSG8O24LAVlB8z4SseRokbFUFsMXkSitfOaDQGTf8AaA7tzMg+Wp3
oSUT2axgNkmbkYjVsi1HLfr6iUrCxFqUV3MGoaoSOCLBwy/BnR/z9kvmMKqzp3dL
/xIDUmLiwUapZEXtTc8Yong8ZVNO9QnU7Bi+ZWvBAC/BAHoHxKZuVlb+LiRw7K8K
5oXOTN7Sqhf63PLVjw6HLHEMrc/5z0lVpTDX+qGepoty45aFLnVFdPQLW2EnTHJu
n11HLrbsSKdGzyVdoQXlMhl5IFn/rek5klYM6y7ZxMAYtBfUAjQE7FEyMotFx5St
YlJ9+JZNM7JAMopgvwWxTJ7/LX8RB3Ix3BQYNJEG9+bpH/6rkRKRId8GRnU+n0qW
FlHp9tpcrsSETlW/cICMDRscdEDGW4uC4xTm2vmGFzMT9dt+76QYvuCMNiqFKgZ1
cFcatAgcx24bjImr7l/G9n+EgXoj2G+E6i9YTtURsZ+8t3EbQbWFR3HnLXVuRxrU
P6BIj8Jc4y45fvKq/4msydxrqJXiexa/GVO2iqgJgTn6Bi0alj1NGtq8QimN1U82
x1Rn9l4wScJHL5RNRXDIyucOeAWBlfhomlpfuS9Xo0zfw2bY5pQ2eKPlQg/YRR8O
D9tp8050dsvpOba0NMGrhUK5s+EkngYOcfDvdikD7Sz4ZgWHGjPg2NMIsxZv7/tg
x9wBG/uvhyfgSUK5slkVwu2kxaWU66Bch84OMddZOTaiLxQ+gUS410CEInJX12ah
3p/DiHGBObPPLcEUgE5Nf12YEEwuAw4t62OUd5/C/WmnXn8Hom3c3Tv9IC5eLDLG
eHQ3XvTYACpwaNG8sSsUPrEJYYDOCnyTd/LDJrAQFqRgpkfWRU6Ut2RAHecx/DKX
pZmv+SlN1YqwNl+qdZ35R+O8lBHFpjHPeGfxW5s+yNU6jMpb1CvYB6nAznNm6zQx
cny2tMqLTyxKrPkHV/Zf3CHH5CztCvD4Itqppijess7clHJfn+XFOxtFxWSte0At
F6wRZnLCsV76QbLNTAJ2PTZV7BQL92qkIkvr9pIU90TvLxdLVBCLhau7HRVz2Pq6
a/JbOhafMEPOtvLwMYwLSV0qwFpPBDfAgCmmg6jQTAsbNICk3t0Tf+TOAFT876G1
jO5Og3rfFsaREBoWDDE/1VNAEMzy+iz1eMImArayjd7IrhTuaCF1jKU3ieveCX6r
M615Cati8Va0pEsupNH7QWdfjDWv/akW1Bz7ARs8yILP1fjwrHFmPbZi84A1Pbgr
isWZMbRdd6VUuhSCHYTU4UFVwMPO10EC/7U/3rejOivj2vIJhF9PRGTJ67iCXLj7
wYVikmXzETbLrjm38ZK1C2WxqYUAZmKK/iMMXHZUfvutauV4M3eH7rf/DMgFtIx1
D5eb/9GSI/9LjXGS+kNB4DjmIEZpsThDnEQm8qzcuk5lZtI13Gdn0F61afOyRQiX
ULoSj6XDZ+tuj7O0saTxeeO2JAhq8cxaiuG3jYp4JTq/u+W6GGUmh2kFIpw9+sKB
ogBjgD1jHx+smDp05u6wGb+4d9HxtbBZ3xxNTnEdmmxyT5Y0ZYEf1fN1twWnRkgi
dqJ2wwzK6NcHjfEwZfd90Jw/O3ogz+S2x30/+n2QMRNCR5qmP5VJU6nQL/IEsgbd
RZ+LUUn4/XbmwRtiPQODWhJEORNK7+yh9cDiK/HxiE3+7mCzqnFLx5ThqrCtqmd0
NEsrOJems1ZEVwz/b7WGcl6HwymcrJMKmg9J3K/Flg2BZWFbZD8o8RV+DO2VmBwP
lGPrdFvyX8C4BsrtV2JDSnup9Q+cvtR6ivx4efLCV1Pl8vQ/zu7ekpf6rLh3TEX/
++C/kQeNq/IWaB+2eqxw5MFBqOo4am+UiykFVBZSI0pQALHlQyc8PbUI9f6l1zaW
WyYHXAKtEqgAFYsSrw2AiFnXQFaMQfu7voeU5GJ0jCqm53vylZL0g7t4Y+1QIvjT
oISBMvUWgk+dvDQT81BJ7N/4bLvbh36305tMtr8psG/V8VDHurV6fsOpbk9ndQI/
S5oDtrLGul5LX+/0KocFnvLBWA3LWHS29jo6yCQ3M1t3AvbbOT5aO0Iqm8JeEqZT
J9+tH7TYCrqUvikZiizlba2GZWQbJUfzPzCUnQzlktsVc3z/YeM+dVJXdRCXZNdx
zGGRoc2gBX/9TM0otbRAlPta5Tkgg1fn8dViOT7c5rWWNj1X3VmWAu3FPma4oB3/
pCqMyfVpg0IAfslB9ZaTJu3abgsGofXxy39g5R1NzEfxHzOkRnUY3XPAx4KmDP23
EYf1bienBjdjWDjokZ2T95cW/uYDSOsGl6OhX3E1iRACwspO+YvxQ9fJ7QVgIppd
2loFXAK88apUlG44We33ZhtMfhhVs4wDDyiH94KM0poMjBcj0nyBpVkOgHEq1n4d
+KB92kTLRS/vsZdu47keRt6oWAG6SmEkckr3JUOjsUTJuh18rMtGOSrgAAdtomMh
enkGo+B08T6OUnm1IqOMov58+OwoKz5bZMc3jY4uUVLLguzzme21zvqPpxJSpex3
Y4WJ67If73cy86q61YJTBKxFQO8gttrTecP0wo0F1aM1mQqtO8e2PPglXAguPmmh
Vhw1h4Tw2VM4qka3YQBGyRO0iKepYQotFoh7GIxtSWJL/FazQKi6vctJNbXp4arK
eLW3ua/IXuCneY8Tg82qeUqpHPPU8wOPS4aYLEMzVMQhVU6yjGS/9fsJ2CQYXdzZ
6gV8LL8eZyTHMwzTMUGLNm+q56EUrRDVV6Ng/oOcK+eNG+oiUT1BkbHdkW7A8JP+
ZBg9k/6Kz+qL57uTweM9PldTRqD+Mf60ZnuCdBT36GwU+I8gxUdTn6UVtgU02R3J
2WJxtDShk7Lg0l4ZNMUv6t5Mji9nsXPDPvQoUqNyIxzpfA95mACNMwOTWkqXxVna
myrMY+klyav4tChaTLno678Xb+HeHni2E3H0Xc7Ti1PL1dX9WeB/vcOneMkNstEF
P2A1O9mRdVXQhBRTrgfZeK9zGNPp4jDmGm1346w0RT7BDyijwXy26KmGG2aL1sit
2QFG/DHO/PJVtCqS88iA7wC/aFDnIhyb2uHCGAweFeY+WfcSZWl2D4PoWJfYS1wX
qu/SR013MZn8TbTqzpZfckgUK/Kbph+07GunGfM3Or15lgxe1x7+8FRVB969MOjT
O2artvDjpPYpS4xXQ2v5emS5BjjgUJqSk8SGy1Q9eV+BkgmZRSbK20xyPW5/6Zjc
TmZuY38aXzUP9X/uGRm/ppQ9546MIaP+CR06F9NfWLIizK4Qxi+vqOZHDjLwCevT
waWp0Mzp+6FXHXzXxxtg0W+GpZLrMpppJIkTsPS2gymdKR8zmtrV+7C5pZi7rJ9r
qUpTmnbh6ZkM0R3EVrtcD1SUaYswofuKXg8U8cmIrMCYOaOYQmftzQi6+hy5gAUp
YabhMCxKZieuTyLKa0kN1698TqjS2kMF87Gn+lzEpyBvWzv+du62kWEL+IIyt5s/
sWJ9YPcMWwE7BmVl9ZcIfP/OhWK1ikDpczjM/BwOxmmonpmCU7ZcoopVhJ38Grha
6plIMf3U6eejhyYZOCUV038F0mybIOx+PlpyPrbA819W6NqHGTxVs77WoaBsEkA3
N6LRt7zOjqg5+/2zg4zNbPpk+zsZWOa28n8u0KBTm74c0oB1CLUWFjyYM0vY/qW2
L1HD27sWLkoYZGCSe6qNuzEEBl+xqVip+YigWGhT2nTi1ABNusIUUxHKwGydnzQw
tdUqvx/IjaSaTDHma2XczHqLXqf96+hrJB1ShP9tuEPQQTizBX9ExzjyPF1IjoES
y+MxRzvq8OG7AuL+PDDXRk8SlX95GZzswnuxuhlUeXkq9CDeDKqJgh7dC5sxJIVK
yKzifcYfL+FlO+QKFNRjKsIabAI1BE3h+94hIOrOVt4wXFtDbvSkpSEVjR9eZ75Z
x2c06Xr/BUavtwiuYaDLXUNm6qcI8+DF0Nsj3rYBA091Vc+hKFJZjPxRZN6BxLcg
Cik/kn69bUYMXxCHh4a/eLMbm5O46dIBrjcfjdZk9VZsUNzy+gaOcvq+MK4MDsiz
GQ8HDwO+QBYS7M27/g0R9k1oGRuxPPctjqQ/Lc6StENyoZV/oGkVvJXG16ZqyJ+g
E7jIQ0iF1KfON4MH6yCxvijOk2J50VJHf15qLcqgwkJuWM/0hHAgXaS7jR6pC7T1
85Omq4TCVKsHPwtISUuL3iFqdYYO9ztmw0S5LtId5LPXL7/dR5YfL/B3X+oUp3BS
NgS1YwdEU5nX7SwGgFoXWldeE4Ycb22KqIWZgfdjuy+ZeCfJMIo3jwqbWMrkjro6
gfOy1lhZAVG3FOR4YIQ+UQtlC1EiyMAaPOUaSDa9yEyPzPYsSo6fgiHXkg0qYwtf
A09Ov7syUCEH+iBD2Mu1S2Br1eNcQ16shASDATldpBiZlSg8vHQ+cwp2IHIx63+c
91Hv49oH+xD5iiOXgVjXbo8GErwDiW92+sAoENPJKtPm+qGeIH4Y4weZtNcdNmCb
FIzu+nbEMrIANe7sGMUdoHH2GxapdEkws1HUQg+x7Lf+Im3CSUDvrd6kse3+mBZ3
yt3wZCQnuAJG1PQsPvYHXQjy4go1aBLbrW5SRe+tR4qnFfLUnzEpUE5qqquYYxMD
xElUxnYECxjNBZUaiYU07pFBL2PPJDoF0CTZ2akxb9uq9snpSqN9kGSfXiOtOb0a
89mBcdRWbNDxC8Wswr6zS5svQlbeEn7QL2zKqgvcHGDJ+5QV39NZUfSQyq99wBEp
QmjYbnMOaGBO4U/leEe9+n8w+3o3NEk4/b3KjCC/VVPKocsXMmib1f5//c7gxSj2
9EPV8H+qZVNu56sRxNHgzcgoWh2yQV1vVS7FzALQeixIEplQGTRx3PP3yETwp3c/
048LskyWSQxRVR2ri37jQNNXYvJXDMEd/sj7+LfIHogo7XALNcfTI5xAgJU9qXwY
vQnZVA7TIrtYIeJAyfPiNcqE1FErDbXRoEotHB/6mp99I4YTjwtvcaesEXQChIVk
4juU5kkZbPAfHQGv/SjC4NOlgwoEJZPKGHrtMCcF9Nr4fSuuofjsSouk5EJ0KTTT
/q4T+AUC5ogDBH8OXQ62cXRzda4mfWbRDH+cdqJbB16K+A2lQINXE2t3eUPjR6VB
bVtRiWu33yEzJh+zsD/kqEbt6esaqEuAQKFlAMyLjOFXbAUQKk6rGCTz+IhH04Tz
J2SjaHu5Ybb1CgwEALGZEzHtOkpS6r1FbGFaWO73Ksc9AG+VSZg4P6tKvNJYom1k
IheIIhuEl/3NTKRHl2xGXLIwNEP4TVBnyOqPQ29D3v0VO1PRrAx1i1JShp3eJH0J
luiD5t3ZstX9Rgbbxq+luWTKW3ttdUUqjP9aTSIBySZ+9jqBm2uV1Dicq/nNLmS0
XGhj0RFAhAdH87BCwlfNKfNO0wWJ3ojVNq6CQzC3uFwemyWn7of6n2nkg2YGZC+C
pp7mm4ToOjCeKTwFy/nK7GuM4JIAhlkxrVxmoDshadg3w4FxoaSk7INsHKCPTY+k
8GVCOD7ewe0sTEi7ghsTT8ZhnasFp0JL/BUtPdWWL2nd+KHC/YnJAvRCnL4kTwO0
VEd9ZEqfrC+GLI4aMHidtbMENgZbnCM2Fl4Z73hBz16bMcdm/HbFBmPcB/xbQr+q
3MNkcr8CZsRtzapdHnBwDb7RnljdDrUuEaaWhDusxt9tvSKoQ8fQXcfJnKOAHO7a
S8btZxrOhrtLTjld/AyP6/XExFizP+Xkd/umasLYZ0pz/gF40rKqND3PRiHrhzbb
91DpTeC53ME7Nj9Bx5/BsbQZ1BDVqIJwpwf1Kmd/lwBD2MB1kTcecYZVXiHQdsUr
yYyZO02t39kkJQOdIkIOZejcDk1cRCVoUAkXrw1FsSS1fe5qo4vhUc958dstlKfj
nifj2dv30S/cxmMst2Ee+bbvxepMBs8E+dvk6rI2JFd3sLInRBSfOYO72H2XJlOY
0LR8baUPrzENbs3HEr4fD+gRRIfGMp9VF5n7KWir2q2kgv7rN/2BlFGIRxnROH5k
p0igXhoIJhYN2E7NMjs8X+vvNkLUtlpwRQDWNBAyKm9zMpzBlKHxr3DYuC+mdi99
8bEzeq8PKqy25aqHMBqCA+SyFb1IGubgFP0Ywl2ddkWoSoXfoQqIId/azIKkwFFm
1frnN4bnB5KgeRH/7X5jj+sHYcEe3ry6SNcCkFXXO9ZxsCu0b7WgwRlOvmMuxwHD
UFfnKlJqCxZQH7M7WVEMzZy5TEAeF7FVb1Cs9NINW412jPVYkeb9hjj9pvjGJ+kv
p+bdoHPMyE7Hh0SqqfP9Y5xrJO5kxNqcyYk9TFihzIXeZ0ugjHYvpOr+195E7MDy
yLxGzbZF4eBRcmwmGLDwWoLruRJp702azaAZi0yzeP1QMsvh86EaF8tY8x1QxFvZ
AowABcAqhR8vGX5z4cnr/9xvv9r8LMilRvgNPkqo4QMbkRXUHQoe1hXLZPkSq6QZ
JmE1ZZtSO1dLMBRs2GtpuOE90/0m7PMP6AC5cIAfgujP5MMY5IJbiHlaAfp4eIl1
WibFclX7S5WsSKls3HaB3MOb672VpsOgra3zN7/ArSZ7qp1mngUdJoHRbJKqtKjI
2a3OBqyixQp7WyGJep+snjBctt6R9avkLi2jK4/Dn6ysNrLmg96zWEeEb1Ps5JMc
WJQGjzrwPJZu+MspXbrsuk67jJJZ0Vk9zan69AK9L3fJe8jBUH0NkSZjQ08A+V62
407wsGezPAvv22Jk/4gBSyjCrcOFT/slv8sHKZbkqnjtY/3ePsNNcUFO/SNg3/5l
UZomsl8kbj4oSsyRHeiIlXlvsVk2Vi+nmTBH3Y/c3ii8cfPp4n8Q/WGd0eWUhGim
0grwz5sA6Ut9mH6w0xZAyQkpY+w2v2pNlcCKkqniPOoz/fR/Y8+cmVeyk7evFTCu
FFle91keI08EArXgcgnwbDenv+m13NkToitDV4gAHOKj/pqJT9V8BR6FdVaz6szC
a27uNsLV3U5qWjKc+hLYPjwoIU5qa2KTIPW5bYsxTk9RTdWIEwJD1zPPzViQhqJe
InYaCCVZK8p+cFX+GdDPmWZH1Fm2RtVo6rgyTgMjmZ2+3TSjZ9mNr4h4N3fJWn+j
uRm9FyHnqLeOneHaJCGZXQR4AflMG9bviwRUPwhksRcMqPpm+CYNBvr6cl6S4Ptv
H4gA12+PSGeJha6NnQ2a4vPLXvgXy7yn/d1yiQBqzzTV/mBk4G6z62QoXJfLKhaO
mEJsWSrKYmI8e0clKbhWHSXdUdn9FKxE4xohx+Mz4AYN9WHSoi34tggtSrUNWhhR
1VNocykev7uqKoPIFy7Gs5W8uHvBjUhW0Lv+GZy1LD+c1M+OxdBn+/kXBR8bvpYx
NBgfIp9vuCCT1gcJMuFnkU1+FPgqPHDm0TnWO5jGsKjPnROqPfp6mlDCYYFYOznm
d9Eie22iiFXq9kIs6hjvizORolE8V+6GJzuaqQYprvg9ALjCjP72r9R6QE+V48Wu
a8IwpwHx1zopOibt3wjs+r+KGHpnb6kFnGBVafR2sFcAQMs3zIydi7EFq5BXSO8z
lfAScTG9KTlcQhZYfVvSRHCFR3P1eDQZHncrOv3Wksug+ptWPNfqgmmnoTrqhYeZ
uAXNBAMpKwPJAibtdduyf+QOZq7ti5Pp4Rxb3SprWo+XM4D3mkne3nzgbdNQ8MWf
7P66dbayYHxQfOmPYSIf/JTUuwJQYB1G+a4lGcWEZClU657RVYR6MvrlQpdKs3zm
NR99fNpwUN52ME3Hm0NavUstZTUuUS6NWchIXRMYh1JrPtx5nVzM0FlTO1VkbbAu
7Y//y2O/7+pNh7V+/wuuPQkKqsIDi4EHagxMzq3jsvIpe858H16NJXLB+/ZOtzE/
YH4nQVenmoJnjanIyr8lFiw3zHCnHBR39jieOB9OQyrfqdFjoFoBvIGWzJJDQSYj
dJEzs99SamS01jm32jN3ACSrUejcM+NYd2//c6aH3qqPUkIARF6buT3ZXVkIiNDj
NXObM+5B3sRDRFkeMAROG3oI3vLen76go2r7xyvkq4Hh1Sm3Jhd4bpoFpu1uhoc2
slZUtG9kKweIKMXj7QLmkTDNZJogqKzDFp4leYzeRilQXYpIiRtqa2UyDbWEljaj
CibmEOTPT3YKdAN8VwyofIvOk+yBAVzShCp2aKMlLu9/hlsypy9zq6psyH/ews/U
0CoFKgPxOtTN3G2e403tldLRq8GK4pDmaPiBKJivZ206apT4emGbxwEUnVn3omxl
Mvgt3ZCgMzQ+F0czAZSfnGxRSC0IDsYM1coiqAUIC5+fLoz7S0iUSJCH4FBRvqYL
OVrY14mm10fVO6Nbkt7PwtKZJwW0EowIapg1IqSgA7BaFSumDhk3fnkpp0bAQz/s
2Y7JCL5K0DKOMu7WJcns3wtX5lXZikZMYLSQwMoPTYWvAlGVkwG0ZW/KUTrJXAhQ
ow772P+6/LEktO1ON/Tzm4RTfjQE5W1STH3J5VzYeoSMPad0l+m0+AUj4YYkTe7u
JwC+WAdJk5wPXlTkKL/Wae7Kp1e/UUaSxPTYQmVwXB5rPC8sX4T7+XtQzJt8PsAY
e3FWSs0WZYALGH+knBWiNgSWuj6wO/EZ887w+jG3nL/MBk01YM3ZOeFSasP+hv3A
6vPYd7bOOj3WhJagp40Gq/D/SkXcEjAWsbAZK4eixSee1j19e13JParPo3yoPuBv
fVnYxK9PIvjWIJoh6p/CKvOcfJAytz8ZXJzlTWqW3C99zEhP9dajL8hPXKO3Zdqm
ke3FzY1NayenTj6bvPiqJYOFP3OkEQx5u2EBuCF0zLjtRnvGb2kXKBR2G1HDxQRv
XL5eke1w1PAjxtktU//Iqe9vhVYLgjWJBLjdAheJP0g9KI0cRhqQ8GC2/3wfsEy4
kajBemjobNAj4lJkfmY5cjVetTuo0UcJMs57kXyltiM02LCDV7NldpTBWQG7MhCh
7BUiMQF5b4KdYVwovLWVnp2fPUqWaDVbCtwAU5zNNr28J6HmZd8nQH1VcsnWEwT+
yJFWPO3jVO5ZU/gZ6kK/hEK/kkzpQKWlI5Vd06s5n2614SNphr4nHZ3sSm/hjSBm
S6sHmCBQIfdhmMVHpvrfszhsceFnaoQFqx86zTo/evC3jCGIIDzmA3lzIQrYxJh7
F/yMycqlPZ8sZFRCulAieoGWu9LPwtjA6xmYRvLU1f8HL79W9yvtc+4fJsAP9J5Q
Tl/9GXpxqkHN1MGn1hXKeLTW4492cRFKeC85wx51+wnlJty2bGeWK1C+R8zi/SHy
3IAp5cCqq2ZzFcKeJdHjNXPOPcHo9ioZzpFKQavkWttXICaqMB5Go9LyXV9uRNxH
TvV6zq2IRMNohoqqhtOT4LgikuP8l1R5952DfnqQE2ZurTA/Yc5b9JuqgbufKVKa
tMQQvqNg/uyLLoidl8AftHxXF0NHsUq2lirdZshY/hVPmtY1+QziOq0DhC+BwlTZ
ANoFu9T5H2p4Hg0Gmzin4YYB8ur61gfdSrtcQUltompl/v0GjigDXgG7nAHgpVPy
W82Y75hajqgU9MGiLxyUOuF9EeWxRd6OFqWuzUCjYSOy0s5b92B6rOZ/zj8+Er/J
tntHDghcWfdnA6bNi7Pi6uYLkz8iXl0iYOAgur1M+OJReXExlwlJHcFDSIJc0+b5
27cNiNzEu+XtQ3peOa64VPNh6uh7pnuVK4ER8RNjeAG2p78g2sWGT1gxmLN9Isyh
6a9qPC8cazy2/Mtjjk4gBPP0rSJj+XAgIFckQom4n9RcnoOhkwCn51Kp3NKt+hmX
DqSr07qV6oupqJ/AK6P9MypnRfmxolvHGwH4CRv2xq7bTxQajKFKlHIfdg/PTbV1
ZqHZhxvr6++KUYOZ2VZBCN9zd3lrWnWZW34ueKROr/bpbHYNxdMkzXFOnU70H0if
3OXTuK6fov6pErts1iUSPn8FZAWF+QnAIuExyJktj6wjw+3B1hlmm46wub4Dwr1f
lvXrX8503TtyRXJJ+1VhXNweRNnPBNr8XPnqHD4qJaypOzaR8UQl+Dc1hIGz55kA
ky1nWWPb3zwRzFzLPepFYDK9wNmKdUysTO3iQ7xNABvl6QzELA8BSWqaD7WicZZ4
YQNwGYszB+in4sXKJL23jKoMUkfukoHTs0qEN1/eQc7dKnBS8uJuqsUSSexVzX4u
hio1QtSu4ILbWSvHBUYx2Y1G7SQ64rT1TU/1GyweuyY817+p0zsIlnqeJC7bYoRr
EwkJMMiLbkMbOMc/Z+9KVFvnIbYvIsvjJoS15BnEljxY3pRP8gj5OKf/EAsolr9U
Qh8uuR9EsWdblDKx5pGoAB3Tp/s25l1apTj8ap974ZhcNMy6drkCMOXgrQglO5mN
70InjizOW33c9v3SYm6OpojVltdZL/h/D6qm2WK2qtu12od1+dnwq2xkgEdygFyb
y/PlYkgwCXeLBzvKR2brCheE5k8ylinMO6KAKbqH4dxjVvxrP5JuRUVNwHj6vuBu
3z9Q6k9b6ZzhQY2fmuOVp8vgypNJ0OkTQURN0c+zGHMpFMIgUAimuPe8+Wd+I/Ae
Lg/TTsdXk7hPk0CwPysoHjrFpgeNz9w6maKlMp9+sD0QnWcOm3700TvQu/jFAQDo
uCpGqksRzKw0qFlasRajIQN5mQ+EGpp7ggEi3fKWHxlbUgMOlSUeVRIEv4ei62vz
D2VW3yPNm+0Nx7KFCo6cpylh8r/udsYpFtxarqFsRN9IIAZVP0RFbsDzjzMwjNIJ
lby3lN0TTUoE+r/Hj5ZVe0lDHVqi/mNFOYwpOB+7U1pdhfRSKsAyppXFze7Idpxe
zIGTLsBh4bflg0eOqzmSRZz1xvhcLmNEYl9YdUUgAmDKugHVRoLO79JG+GgGv87Y
ybJ0t8RiLdrF39cV7UR/qGigmXcIQjbf/rhM8xCb06LHkAIORwZKLbr44eRUax78
Zi3D9dcXSAM2LrhZ262cZXzTHMfXa3VzUXafo5mVtBAIshBKgxk+zO6RjJYZ7Zk8
ho7A3EH25vEj0aCEAWLCZXQRvy0XRB6hej3tWfMmK6d4muXuxmYS+RbWOZjIzGCJ
pPwN+mDXrvwDvhRxWlbgPDPIDs5b3QY6To+SgqahJwAGQMn5zgcyIpl7rtykXAI5
HaKBBvAKINJldg6nXYSxCZz/agzMWv+Wb0bX9jOqO3CyLP3s9WVMpWReawtbtaAN
OhF9UNhasktLgnEXlQMKjtgi6b9PYaIzfOPDoaDVBTFB+5FVVwHatpNjbRdouCZS
yK/qhf65byRkmwC/KtwWU+chBKXBvnIBaMUbdTkc85l5iKNa4XyuAqX1JanoK/jq
mkArfdX/mLv6VmkPQKhjXn1Z59hu/aDicgqz1UBIt4eM5CCCWc4f1YxgPVCxrrGL
Rfl3bm2KaiAUWeuFrE3cDsA5rWbZtQur/qWeuj3U8QfZwRYWKUNDCew37dmw23op
aljH0lJ71YIFmxpczcIBkUwF7EdTd0ODX6qzIhQE3YkOnixry2M7J5dco3Ck4jcL
os1OmOBw2ytJzHkHxnWVCiP8hkxJMqH65xMBgqfBOJK0qQ8hFNgFPeqnIgunQAcg
D6+zjVmdJ7N8/MZfNlB9GiN/zfAsN1VBfgvk/CN9TPlxtMH38MziftuhKYGHVnFm
05tBxt6U6nxv/+biP+gReBC9gzC2LOlyhUdIUem9Rukf03Whko0B7CA8Qf6AzN9o
TfvWrQ43vS6dLJBh7pIRoEZLZJvtrjHVGaxWOVNck4McSAlK21ve8zMJAujJ8cnq
CSft0Gfg+1CZ3msO7il0AXydf0OrzeB42WuI/UGkDmfIUg+o+c4Vg5Q+IT0KLUPk
ckOW7C1H7pvyAyEUxCrQfUAOG0eR1ZhEkek/PxeJ6gde+oTA0LBtoJeY7f1jOtVu
aBP25oB2FLw0eYcWunwArR3xTjGGeLK6kxPtCoN+LJnTn3VVTI95x+5OVlhr/6/h
MY84ckhIWz+5ZLgR2x24BepJOzfvh8EWNIlL+p8bCSXOiXlLiYjcoYVAwhLa79tC
dfW5t4K5uKZupGt4ZiuezIhacXSmIRO3PlaXa8chC03OaR7L9IiTHZi/CdX8GKdV
LehboxARu4plXWFfjJRklM++0AhmD3J8qVfqTzOBI6YyWCf5N2fXVdyBoX+BBmdr
5B639qlJ3t0W4fFdItVlMUIuPzX8Zr5ddJHVLogkyynsu1+b+U51/vCM+tt5mWmM
mWvr/ON3RurGC9N6GGsld3VCpCOUElWtYh5molTr1ntsDfmMY5ritH2C0OYhK/zS
mu8OwxXPllcf0pXM8AgI+EtZxSKa2MnWuoWs1iTDPZj45ZL9oS9LYo1sS2ffzO5i
XiVQ2sQVK9tKHMhrRhyBndEiPViRd9nZY9gCp9j1J06fo2yTiMrjhT3A8KkkPvqe
/WAO4YxdL/0fNekLEeb+OvhwDK80QfeiIBMKM8MSQtPqih6S3KLMc5s/EcRxBOnB
cnDofgHo7Au49Dp73mLuOYt3Tn4hh1QZU2XoBNfy5SxqPPNFcNQadTooqjoJ+SZS
UmdX+/Uv/jkhvJALQGSFbzRbXz9zObvnSpmck7EbBxBxTvrzE3Htfc6OmambmJ9r
aKzWFNt4b7J6chO0mcQrWuJ7l3JrXvIAgmqnLs62GBRtePPiLw7Rk4e1K8gXhJyE
7arQ6Bx4cvxBi5jBHEim+09eukISJBIxTGcyCDWYE8nT7Wtp/PH/JwS6uh8C60kJ
jseeXX2rKoST0XKO/Y4g3MQoI26/u9s0yZIxLkhhlzH3suPrglEcx7Iq6LBT67QE
bSfGynZPSK0CebTeEbnwap+zJSGN+kPgJT8fvXg/251dgigYKnCjQqEf+KIju1l6
9qTzB9TM1eMqEk3VZYQcr5etQonJtXW4aZIGLnQYwBgNku5SeNgqK72LdCSZsEgx
ZOqmJLFc9L35vdLPE45idDembOx9hum5igw9YyW/1L3g3H3qXgNxtrFJKfK9oWEg
U8A/nmfO5gk5nb8f0fxiA3Pa3O70VM2P0GeM+oOExc1iRumicNKAclvQluIBS15q
erv7BegFg1Jja2t4hGnT70WEipi111zXzWQ7xKexa4LKB7vVEXCxFxlHp3w0ldGb
qk7s0iA9FX7WQ5gR+rykJUssDmNJH7lbecidnqaA3H/bBz1fA0V1h6zbM19kO32t
gaJtknVL9rbljgc7e5ozfx/zioZ+tuo4RkOc6tTGUW03rRJu5aFxavNFpfmVltY/
vSiMgaU3P05uqhxmwdYliw8dMej7R1K+UVtuDEeOHIFazx0j2cznU0EV6eviqFNK
ZUQL4epmge/QywBUncVfb8t1tVoBg5DsHFDSkgYwOFiettScut82BGUUQqGzMhGf
UltW4rkVbfPwCiqSlIxrNtmthOQ2Cgeq76P4mWEvD2oq2/F1UWwS2yb4j5X10lOz
AHY2xcd3+LXQyxiN6acTI2qo3ekqoCoC29KUDCcD0F13gM3XO9l1a+szU5CCYNMd
nlmJcH5uzW8fG0HQH8g+NxSW5n8lA8uanVECpM2iAPbdjBqrhqeB6dh7xNPM4ssE
gtrh1stDkWlds3yqJWxJ9TX4rLRGH1KmfBxuZqOERNbbVsjY3fLMZLNJk52OPqZe
zSLMKYcQDTTEbNU1HnJ+wl9Hlt41Y2jfu80WNATzJgwPm3nTPB5boBVdN9To83PU
QM/KXCWKuSPrkOyrrndzw/NJ2kt8dtkVhrgGTBCAJNonUSxH2skrh8px59QLJZMp
byCZKTwsXOCMD7uahO/SyW4bQNy6GlbgBg0Xirv78eNUBAsocsF1G7m7ZQ+giGqP
++RSceZ6DMrEFbmGBTMD4KSEnNwIKDFYqwL+aRq17lQwUN67T4DF02NWH5onnNS0
sJkxsovhAo9gm4kHoKiA6hqm94gQx/HSo2Q4GTLzubgyssaKPCNwGA2oAriFjwR9
vLadFeQ5mC4iN1aA/bbP7mxVJsJYY6Fk+PYePt6nYvijhkDsi6ddfgsY7kBHJBaj
qsh8KEffqVC1qXprSjG4BTd0p/MdtaNky7HSHesT+/bedosquGYVrU9/bPT2y2CI
ouJpOQFN0IYrl6OAimufV8yf2B5Di22RLIkHPBFXi3VbNqw+KAlU9P3M7SEhqJ6P
TL+b3DmCz9nTFtTRtLZGluxZGmwUCqTfs7RGNjFSPTitH5Eqk7uVLZ9oV0B0f1Nd
b69lXgkbNQGuJLUQTn+a/nDwk9OXJt7jCmXJ0x/GV2HT+KvoD7Py6UTEdtCiHqg/
Jk7ZeymX6ocYcAAa7C3CBFsvfYoUuH9VzVOcXDyDLoizSXHs/0h+fMELKd/i39ix
wxNbtFJ+gdMmG4pKejj/7j8VleTqLBTXyZuT1AhQQbilW8Y1kuXdz2Z9l9kWHfDt
DZ2yNC5zfnhnYLISDVVzqZ1nbykXKo9SQ65zwjDiv3vSWyeLLA5830e6NAthp03b
sV0XVkSrAMLX1i2nzqEwLApY0GVChzGDux+NfFe5tL2/7frszlC9eFYQ/7PxQ2Nr
cBjcQDx1Ks5dxAV7tkyqBxquPKsu/qcvHetofNQKJTuO15W1w7EF6w6luyhZYDk/
PP82D6p/8vv1zisEZKU3bifp1dMBhtlO/t9b0/guUCIfOvHe4JlCWqiCixRc47yB
230YxG5AoXVqlzi5jPYh8e7fyEe1vjg7T2LqfsVH8AePXbO0LjsRZsR1LPvAUMU0
+Z5QCfVgMKdOPT/AUFuGLX4ICi0B6BQHIv756c48Co++7Zx2eEUbFOMM40NGR4Ua
fGAaUj0FMK4IfxLryCQojw80bajJcd6Vz9t3IrTxy3eod4TrFLOYp9T5fMRSNEzg
jPegc+DgsWMUsTni2AGEpaqRsg/AeFifHaJjsZluzufULfQd93khTk+21dppTpqY
JXrA/SrE2T/x/zpl9Sns9+QdNhoYNRumRfj67Sd4zAW6/t9j75aY+bcCYj4WWMY4
M+kxK9V3VCE7XnGb+d3iB2SwjBN7fKQ5izzEDczyRsWbeCAOw+S8X+bkrH5TS9Zv
5V7n0x0NiYteBgbnwHb6S2pdGM1qg1VIZoz1hWuzPHAOmsu3dIB7jN9chAuKiKnY
Q3EjVVlG6WUQPGP/5VyQ2P7nhFU7NcF0ZVQs7u855yxCONH6mH2jDIX2Wtzcj84x
SWfP+kPfuuAHIByC/rPLhxsbfquaxDtspDJsWGQ2xsskssmoehDqJNJ3u+oVaeX6
qOW/4SyIbWppuOroXgr1GEKRs0bAb6s71E2HwFtX4weo2JxCfQWydPiiIDgAQIMx
MyIUb4oZi8akeDkOdzCvBMlQ6Pi/ujgRgXM6grDuymhamAyYXWxy7HutdmmExkxK
giXeksfm/tKzlfnj2f8oCadz+gdk+DtQQCnq1P1OoGRnMTaxivuPotCcqors0uQg
8Yo1Hk5aD4BdE9ByQ9UWFFjDyeP0I1UQTbI27EVuSh1siQo9Ei5di8y3obWYk+Yv
h6P3bGfwsbsvC/J1PG7u+IHXKZKmvWNw+qPX6yTUfdKgIPkNxqeEZ+puO7MI1vUf
jiHe1JvYRsCPzJWkGV6KBInsERvWRvXtIP1RkNZDNK7hwr/5nPRu9wZ4BSf693dw
ax591jl/t780vve3ckn7QTmXkBa84M34PYhjoKTQOQV/DevmOvvUqic0s6VeD3Lw
ayYvkwvVimjq0TMEiosWnTq9sC7+98iqXy8SQ3wq+BFxRDTscAyGMiiDgv8OhFGw
/0CbVVkvJzOjE8FAiDdA7oDO09avCS4C5HEEbEjKixbZEwCPoAD6jea50fb5/fTb
83OktOGmm7ZEzN8E3P7mkpsUyyeSFVJUV5iLz9+E6hBO2b3cssX2RTwh3yXBlRy4
Nvx3d9/j/SBkYPwGuZi7dqa4YGtgxPcmrizmlUnsLC/4YLERZNPK/hB5b0OSJbrz
KWz2md5Penffuj0NX6tOwT6DtoNzUYZbyk0ukY/podq40gv+6kMNeq/xVvTSvIZt
slv2AuK5xmmY4SO7yQdZYlOTSDesdEFkBwvv/p1/psqT90eQYFlbJDyaivH70i5b
RepL8yIdcnG82EtbBbayKMxONmoovJ104c9IyXgpU+N1hB7rxWQl+/PS9xWeZOYE
MsUIq3ZLLBHIvw8mbVTc6zsHi2CB2rICOjxumQ9MQPb0zej4AA5mN4ZBTjKMTyXl
QtusjCuEMTCEYZXiTd85fCN6FwajDzx7ysVBd6BJCLJAmWlWE6/wonmFBg+y6hyD
rNUSZ0xtOXyzPinjktS+yl2IyWo+cAWIRi9DNoaCBClBipAkOvyr5U6EVxpVsheq
PfIgXpzmsfendS0lohme9Pk9MT2ftYPMj6YEgCrSybUZLmv1g7V+33jl94NGcimH
ky1Rj1haf3j2RI4SIV5ywpwh8JfX866QuM2g/kF2pXIwidCKz7S5BdBFLGV0BeP2
fHgdm/NyVwbyS5RCBg2kWmyQaEgLv0ssqZPmIL3x+ApD4sjMI1S12vT8TusM9hG2
Br/htrUDUfPp02CPfxNRyPC8mqB7TrOSsUugHwtyLnHIzzFGA/dhNoQiN3GA52JZ
18xzuuK1vyjTs20+QdOcH8jvksRtbJbvENfVQKA6Lg13IJEKSrt+go73bCzdpPDN
lLJHJilHIrEhMFW1N7CsdJJMBIEoAWse6d3085pXy/0DAbRiOuwQB5R+Ehoh1tK9
XXQiYFSootPxx3Kpv0QqABbyPS2sMxZowGioaqsyxv3l9C4efE/7C6sDcehIttu/
GJtdu2/Ald+26RmMfRIzZJMvj6svURdEpJTgPhuL+3ehpxYoZUOSWbf+d3RYodYj
c69QS/jayPNynwcaJR9c5KKF0oPycPF1/5pHZBw0mY4yGnRM1nk+QsKOKJavQs6j
exCdHQW0d2P0eRDw8tmijxOxxhUT2aX2bLrGjHHih7MS785rOHwOYssquRT8CryE
twSZR6XT3NZwz6b+oWDpz0C2KXEYIcHCyxlSa91sGuJSN9WlmQVljiUzmmVQC4gJ
I8FFvBOnN3gDYKFCgw9mUHPNNXAnmF9dQI8g1yawk7uR2jZLWuXUkKNK/HgXcJzr
0V1GvFdMhC0d3WEhD0MIfpXe+fV0Fqnad4KdVtoAxL1MhMLtdaROpccQG7zIS6yc
F1EehTw/7COZ0EDKeTBwdkLT2IkYFct1hC+DJMtBSCx32uM9FfyfouZteIxVycfp
k12idrJOeaGiiXYJArens/9ArM4UdJIYQj+xbiZy/GavTRiXLnKDTCf/pFHHIqBt
yuHN4iIgGmzKJYw5DDCkVSI/8qqAfH4ahAhnIu+Wx8QMtTOUm/QnzT26oECuyhve
gsLUsydMRAR+WJzcypwTg/SvfEmus+KlfDMZqMsJ2Evcm/AKcV1v/NGYmn6JYJ3q
YfOBbXhpL7us3ahe/YvEAHIKUYyT3YHs91JW8W6mwj3THBu5qEQ1C2oC7x93mdmg
tG4/yU+Pa3dNm+wecq5EjUrlN6RzTqOX/A3dP0TRmIMvmCBhQkyhzaImFgdxBxM0
7w2wZ9u/qvCzus+7VT86aHooB2XW9MvaJNq5xXTFfXXFNzeG+MlIN5gWpk+K45rJ
vLIudB6O715b1rqGUUIjznxiQdBHxf4ZmdDRvyWvwQRi28LBc4NdkLlJBwD00c4x
nVPiNPpIPzShqAcbEtDKbFkzH+kFEBNeW7Ndln68uiKO2vxa9SQNT0YivH4XHDUl
FeW+x4INQ9cpMukVv0eIa1GnTvayRfoc+F0ej4/CSx5rRcAIGuHXwdatt7h7acRN
FsNul1wPuZj0zw8oAZGmTC0PdrKgKnO4KQg5ittYhvZs0FfOCQEBv/1Rx3MK7T8q
AgEHmt4ASGbQXD/ooNbHVo5NMESASBZaJWe+v5brbvXY9rGQXd/EH0Eqpac05wNR
WvXMcz2CJ6pnYpHtduTSBVD9quUiXV0my6fUaL26bq66mp8QklvVTK7W2iaptgnE
P02CDBarrAyTpvvErfgSuWK86jrxSYlW2s0aU6kuVmNC12u+z9EaDS5tustrPoKd
/mDxDh7VE5CAB5ekwYb5yZrqDOTNojC+jGP4YnixLaY+7rkTLJ2v11Jpm2AYpBcR
t4z+pcilYlv2BKkTRMsHe5/KQ626CjxU75VjpJiogslhVUFqWdMWyPnPyAUijN88
Ci8qG8u7sE1ozQZATfK5/kj+ojMGxWL4DivekBw1S1TFEl0+uSgWke0sR2euWviZ
RR4Z6tI8c/1Q5BIupDsV4On2NvuFucVSZW/Ls991S2Od5DL0hWxE2mIZCGOevfRe
GUxBx80lip6QtzwwS8ue66Iqz//j1wDws6u6bGzSCWJ4+lvuH/pvUn5hTJS26Upf
MHYSz/Q8fQQ/1og2jBZnOoGyTSnIUrK7F3P65LFNfKKHJGJgPjmLMGvUim0UIJo+
qDQnGB178kc6EglieHGHzEskdDDp/jvKSvG/SsWuoJFrXxD6M9wYXYS0tTiO4sSY
sZxCOOvFqS/JPJOUt608tO44ANACujlj/Z1/EWnFe4c/QvLo7VrcKRYyqDqf9FK7
3DWxsjts7wUIVCB6Se7NFwZxq9RQYU3HobGUBMZeeUm9bIRcZXyM1USCMVGYGGVf
pveFxgucl8DYtog2K1r6bYyPtYVqseHUZfuAJYbJzIkoKaoUppngCwfYYu2yhCE8
4b6G6D+/3Zr4+TAAIRpr/UfcWPhFUayWy6YwcHo6e6gecABGDC2jSeBzAIJlbSqw
c3V6bDYY1u5JwlxPRF/+1VU0cEiZLsz2aZs8d1Pj0elhBYeAKacYVenpxWl9eZXu
h1952nMk3epvT8wFr7rDUHpUGrKt1WyXEzIX8zxoRkrm2J9B0ELA+vM4psIVGKRZ
NHAjnsB+oNKfrFDgP2o8IIWcnEecszt5iLMgldqgdpP2nEHBUMq93gEfHm+6qviY
z34LQBy2yNC8+QdZTVb1haU/d3JIuTaCcQxu9j3Sdc9TFOXRBhUVmR0ULmROQVgP
Gip5JrOTlMqpt189X75Eqx2XDgsBQLpF+QMhWbY6G7+JI5vVAvZvJPUn+MwtlXdm
7dop6/19r97wEAqa2EXtT6/B5tenF0qU/vx1IIlc/k4Mrxk8aBv2wtLonMUC3xW5
TOt+U6H/NAiskGRxDRfdycNYqKIwnrZig2fUnFGbl4FP4brHG50qaLJl7836wtKQ
1je7xtEBNlHZh6YEcQdnloTFS2zalKekWHnVEFzCH8zslTROVGfyVKo//YwDvI4e
ewj/FNXzRIwx3jQEczHOlgzY8K3RgkDNaqqyJuW+/GMw/palOjUjpu7VNLZp5f+I
dqfhxMxWbTucc2I20xC8XmuYhyFF445C5LSv6NTCvXK7triK1myUqh3MIEqHwVWf
07PPRSUWGexWWZK9jl6dYDalrZrjaBg023bVxfetfV6haoMt/aNFL+g9OkZNsyCM
quMhL4CVEr0G8MkGxdfRIhDNbjTsCIZ50qX5nxZg/f9H1SSRxZ4owUa0MO4flf76
vY4DWr4et8QI8BDbsxkG7JIZZVyao9Ef1qIIKW8fNld2XjxZGHb1/YJGUU3h6ZZS
9pMfwD/MxusQI0aBrjR6y1F02Lclgfup7i/UmR6u/J3kNAz1p/EKn4h44QSGRv6L
a0rD8/AOaPQNQwPJ7FmEtIcLCZ84N83BSzdeVxJWBzMpHdJkQWJqsLAQFPZAFIbc
aYk0j7PhYKK7+jcAAnwWntLHuQVITb/svtcJX/JvxXuJWGMFYPIFGAZ0PnlIetkr
8zwz5bCRQ7ahcwc4jDTvYC0mvwNo217UQLx3ZtjRI/PclUs50dwvbFS0CA0iyCpl
YiQ/dYKshnahvQ4SZnTHsxOswL5WQPty5Li+y1aaBYuzdBm7YB3px8znjUjD+SJG
fVTtM94/UeKzmLouBe05Q70kvRsObMjgwwtGsZnWUVMhhDbsAViNkF9ynhoy+/8p
0hwmAmf8TGs3t7TPlwWw3wamSLmRAJsr5pUxrsmy0UDRxNJ52WlCHMp9I7ar6ekJ
P5CwY0u9OJDDTB4LOTG4cKtmKzNBcH1+aqk1E3NvF5pWul+0VQoRLKE66Bw0yf+F
gm420/vLIbjr2tvbyxQfMB+T069vXo3fHYEfB8q1M9wWQUz3yjaFmkcK+Bd6QPeU
K7IvsTfOHHpviJDqKrLImaibHmh/rEVenE6m0+bZYCz+Y44lJHKjlVghqXYE7/06
yxERTwBPzYJ/JE6iXGEoVIY7YcWGXOnWtT6idKht2UPoawA8t+5XTonsnnFG8gCt
bqUQ7L+p8f+rpOfuLTN2xwI7EUe93FWBFoC1dB34gt9EjC0aqUnipdSopAbnKg8r
xAc/vqeCN1mncy89HIpjc8ZhUZ9PpbntdP9pIhOQk/MvqFwZifjj/YpLtUb+JILZ
cDHv6CWaFy0qP9Ynetbg71FkAaWODx1/5Fg0458Tyny9iZCl6Hz0rxfcxyAcjjTL
d48hShNbYH6B3Pl2AAg990V0gIiihnID1UqAN1nB4Qoq1iR8LkINaEiVEgLRYaZ0
C8R6WjoD4FM6Rtl/oAtPHFg3fucZ02XL1p1DS83GPg6g3TQ3trKtZWMPCb0g6U6Y
fcKfpOGk7A6We3UdTKLRJziCqT3edKq2LdBU/MvFoKeHE8kD2BJfyQXrZN8q8dFD
nnJOiuxnGDhc1EPQolbo5Wnv1cVGL1/yXQtxQQ0mfL9U2cfbJd4qt5IZNZDZpfOl
qrJodSCLcKCnlvxmF5qXpj9iW2MYZVtr25Rj2SZen6C4bX12KEmNTZAaFZqSlHRR
Tulbj8gq0pPbRHQ4G9NpKouto4xxW9FWb+d1V3oiOTBN9gaDAE41SZdM7U7cThxw
27g0xIFXd2spaIz5Cn06C5MVO7ylpat8qUp9iEpNj1VWEzeVo5XMcES5E+/RBHmP
kLni0O5ETZFdqnSI+N4xAZ+B+HQs0g0Ki2t8WRi4+oRd3E8FNAdJjzvHHKRgnDZw
HCTBGOWm08Da7ERj6TIy5VDmYcYq0001/+cGNaOcjBmgmYPDZAy9x50+vF/jrp4G
ed5OH8h2vF2L7k0Mr4qvZfv+M8cmYljLjZXT8zS3m1Q1Q6Ze1Cg36vUKHJfvgxve
5LVJvoC11ZvYvelvzmuwW6rj9D1QotPgsCHcPLSs82iMizpOatNQ8k2obaCYXVne
RssGG+c/1I9HvWOGZ2hPD8LgZr2IiXPz5hNCAKksmmUlhPg05std58ImeXu2GpxI
SLwm3Y0eJYOJrok2ooyf9ui9Cl7ty8rdUCIaEVlwXI+j+eqFmsMyIEsf3Fm8f1EX
zINbO/4f9gavLtUsUTbQELCz0T6PIbbPP6lukq/HxUYVyrm/Dg+EY2XE07FOHeE/
/kbS++C/2S+87mBp8rACfy4izF1jw7fFlonWukNYltyiaTaPCxF9i4uJoKTXWoad
ua01WnFKtQN0fTbZDJ3fjRom50oHoFLXSH3fXBOoLbkAR3Hb9wRlxBDMgcyR70k9
b+afk5GqnFvbIhrbUmgNvvREi5WelAN1rSGh8lmA052b67poni2pFa7Bk1OTlOCe
MKYn5rXHhq30NPVvothYts5GPWqFZlAw3IWNWVPIlxKxKpKIBuW9Q30tgBgAcZoH
extr6SymE82moNFolQSCwaAb+YxufKILGc08RsUBUzgjLdSazmIqRxqqVdaN3ONA
Er+w55jlY256dRU2Tjdr2GIXvcqfZrioY+wHCpg36t0KE/uXwoG22m/rDOVdSCHT
tJ8YPEP5C/LQYij3n6pur/At6km3dygXP0t3Kf4xOy0yiXCpf8twqKf/MapAJSDp
ROQH0h0o5ae8sqxdm3MoNYOrMDa6uUUEFE40i0wIrJaRWEANZELB2A6M+O0zrCaK
0lniT0ZC4mBhUScjV8ImD5LxOFskM/3Yqns0koEjxQk2q9MXsIkWCuBc81q+isd3
RKAD4foVThLJjGfTVHS4b/YR4E/9/jqwM2cVxzpAmW80jo22upzjK351BRzYfDD6
cFlK8++05qvcbPdPzIlQH9y4i0Py9G43Kn0RqvO7E+2hTdmIVpcr1b9JldukFjsc
Y4DXtR79nRARtIKFegpfB3cQib/hiG/RHCzkJrhJsLgC/WnFMYSOLbHXwWTWwWEw
Hjn3jSN1/IJy+Y8iIjhet6XCLnjBGlg5wuGijkHa62+tvVNeNqVu3YVZRtrlyJ7O
WGrzZjbJyt0ncAH8pYtzUZwnkEtDs90iJe9ne6zTK3RDoaCd5Ap0ukAn3nPt7E8N
rml1SRwLH/0kiYQC0qt1kRnbEBNOt3zHI1ug/zFM/i7zNlYgU+vHnM/3YmjeO3Lc
DyZUSb0g/IIogc9JZFh9ltKkwOH1NjXStYCtsRmuBsBj+/D1p3DGeoQR7t/nr6/x
C3y/d2hEigKloiQw2HmFhhWzdorOOf+GN2V90Txx3KhUn9rT2PRlj9WLIlrOINg+
/Sp+a5gYmdKvKSBv+4Kg9vUFR9CiHzPRVBBO4CPH31eF4yZJIiKNAi83or3qXh6B
lJ6CpH2rQeaL3Gy9S65Q+/9vTg+DY+VlZdef7AacfdCSrXXcQ1CO97oUXhCPKHQo
zl6ybzIAAvxtoc3zwTEzleL93O7/ZpUq9vFiBcFRdfJ4pzNwhY/RclZWuj6LCd7k
UOk9fpG8C28GtWPG+IIcV2cq3EhW0hClLaqCySW0s95oqB9F5UGGcANzBMIDFIhk
pQsnadVpaa7c/Esqe6oam2lo7GpU6dLmuJwZgutjVGKnLkXckRSQYoscnDaZjwXv
U3R8LwDMJsuKA6to5kZq8VirjgBOan/KcXHOf0h7nFKxuBhk5NGWHP9w5AW8UBM9
/Zqrotpi0R9jK7ME5JVBOnDgbLmn/sIZ7ToOR/ejE5Ld+wsZnSqUL7gfoWx84rqx
EdrJSoqmnilaelr4w6SUFVYg4damim5Y5/nxmOfCGJBGJL0tdp7ZIsE8bS+BQ6rX
dJNbhGihicYkVck0ehZJni0CYGjBWl/ka/UqFRxCtAcrXGLV83vE4bqutefzlgmi
+j1QqM1M4jF5lOgRMR6j/TrUmJ/gRJajcSXDUc0HtDHdP1UdIqBkom0QbYExt2Bb
OvRoNEI8zuv9VF2LCEsgf56LGP1KayfctF2YDKH2X1YzxPnDjOa/G5BEsH1eQ+w5
KKqub06eMYEbukK0VZAQ/WKXyfkO6JiA0mbgysy0tNNX7+m3Ib0Jv1kA7+Bo/vHa
ydjAFf2cyEIqRHro1oYOSRB5vU4L39PwNV/vlonOQCUq0Nji8n+tEwXjcLWkuFSo
YKOyGBfwGK7CQ1DnLCsvfzzYY0YxDvcjpZqyjBnQ2NA76vp1+Lzbys9r4AOWZXeW
ZHw3cdETr75m86yHQnfY4FFoFGe/xPQ7miAjVeZpRogeQ7rMEuR77A8aUEP3Kvwj
oK/VhiiwmHslCiTHG/uyx+DOH+RicYItLeFEuwMO6t0Bmisq73+SDNW2z99AkXuV
tANeakgOCU/Z9Hh5x1s87cfFPL88p5I9UxZGLRdgkBIzN95J0HuoAJ+BAITNgGM9
T7CQW0ugy6LSww2scIGy9T55U3WBsGoxxrVxGqoKCiifBLliq0KPs4uG56fGio67
gq67t9tHF81oeFPYLEbkslkP0cFfbsKmulzqIPK7zuD1CQTttLcvcqD4CUyKycdp
zNVJoo8gOa2eXTUKXkfvQpzLi30bDbNcZh10ezpLX8OA8j3TKhNYBN05JtNru2no
o4SBBDdMUIOVcOuC5yqOEaHvNbrP4WiXIgWYkr4XltdS0k3MnpG7chHpPhyU058S
Bd3cjwDd6LCv4+uDRCxCelej6/zyeRmVzWSc3ozw2O9jW8JPGhX7mxM8NC4Fdv7J
nPJd91Of5WYAiu65brEwaQOOavM01PcUIwC2+hgGk2AkLaZlYypuLtyYJnlM+iso
XouDwpUqA3iScRggW878G+JT9Y28k2UKFR4uPr25TNSAZfK4SkTDdRMaATYbAfy4
xHf+nypSBzEfe5iTPI/SEKtV0yyHJASsFf/5SkfKnXAQt/3L/LqDEHfppaf2QNPk
THFSWmmxR61rfF9ql5i5Bx5C1xvv8YNkbEGqbdxKQ766sLKRZffvoSQ3f0KEnKcS
T10u9cXRk9QqBaITCWmvoUHye1EKHc3i8+wjWIYqzYOcRRGpwG9bYJ5ZGYsRVFJH
dAbOeTiO2W5HIxj0v14fS1m7M/BLARfSx14f5bC8fPpaEfXtWJ+gv68C+hqQ6BZi
ftOu6iBZ1PZUMTRIQWIGrfXLSsIBETXBrm5DPMqqlvVIUQxCrejy+9db2boZ8A/5
KzW9zUlOI2zk/NQ5Kfmsk51qOJPv9NwvXq5XZuXtEaLjdhn7TV/SSNqZjD0uO9ed
jYSWrblGfR4h6M7VMrmhMcSefIwy6DiwarMbky7P7Fe7UnVlmBR4SyOPUtbQaknY
rrCmiiS7JeUeUZMyUDEeKE/CFO6c1zIkru/G6/Ow/+EFwrDWYkh3tpxWUhXc2fFF
E+D+hZHbfD1lA5/90mOFto1ZeB6f2Bi+XVnKA/XMG8dURn/hFk1qoHEkELXkjkgS
qo7ipFtgIAzlr6bRD38mWDjMmUJieily4ShkIk4wyNtjALxkuEdio+YTV4XUVT4a
WSxsgrOpdwYVRo56/HTn+OfELG3osBmKlIzFeB5skOFXNzcmiRWVy9mx3blqhiLz
h4fDW/Tik7zhu9PULNZKW/rgbw5hChU6wr1MrDCNozlqPhvtauFPg3trPiO7ZVBq
wA8bvLTsynfaKuJLJCvYjTzky1nbpCtLy/9CWax7PPyCu1j2WDS5QQoXYC3tXUzD
AFiUkpjbJZYMRYrEVlI9AzKAv/Bswiv2LXj1OcpJMbZs9qLQzYKcytv3UaLSvHUm
D1YvAaNu7wJc6xPh58j48/vifawxSy3qlvgut/OZUTqulMyElBd6fxkfpnkIRsyl
tNqbfQR3YOZ/b0Vlmp6+KGZXJq3ViguQW+5CNvsSTUR224gDAIHlllu3hToz9AvH
vH8eSIes7fVneqzkuM27vDrHyweJHsjSizPlz5VI3t6XHfWIeL+jtabqeQODmPD2
9tza4uc6UNe12yvs9lh7jkGfI1rahliQ0Dzyc0YIKoBY5pF3BdfNEmfsaO1dKFUl
Fxaj0fJ1MVSoRHfcyrNmUfgw7OEYlv/EgWnerqDV4tXXn6E2JPxwqO9CVZUKVVTT
wpFlvMlZ3aNwNibH3v7ljR3/bDweTDHrXWOKML9fNUzb9PiIkEP8ChRNWzM1mKCa
tLtIBDzSEY+VKwrMX7wKrG6rk+ArCHxR3afUb4ZCnQu7xULO8jA9rgMZSotsXs4f
IxJ0QWvEeaI+w5/W2QWWl19+UYBRUpL0lAEmIukfYxx/g88tR6B+5qyL/e42qgBV
Yz/vwhxQELqM11eaoWfANRNx/zEVnZ6+q7aFyQgUSpDQdKEkwSB0QTE2hqobRgzW
1pF81nXX9dEfGvX3l02kYY8tMVxqJT+7eLa/5ok+773LdglnxEzSXxs7NCMQZaFO
wgZZoOjTvKPhGalVNp7Iqgjkv43QEMLPXCIJSF2b+i2LnnYDyTA3b1UsoAlfPiNJ
eVjwxtHlQ9PUY/xwPKgCXy1XXEQ//z6EBBv4Tb3Aoh+QLJpPkrqxAU8TDZvDzTwh
xWRrH+uX6hbYgObPdaWhHGSRv4XrukZ2kKK9X/p5Rn3A8Wmph+fZJLESjxax0gD2
tZCJpnpzBXy8VtccpmUufLmmUY1N7+p3jRttz/LyGCMHG/Km9tgzyajwKbup9bpJ
c4irXWTEsqDpawdyUlkKbpeUyWJTekuBlrklz+cjtVEBKih+x1WRr9JrSgBvpk3z
AhUexCaUW15X69z6AcDzUYXILS+wCtYjmMMabQNf4lbGOn+I611+6aPJTSIE2468
HoS6PyJsxk1Rqpo/FrRInxZy0P30heQFJ386B2oROPB7NfwDYiZIIijRIZpk0Qmg
oIPUPqblhSGzGHf9OD6ZtVmIogvHKqVRpz//K0Sv/YdQK0omxfiZsZeZsBq4dl0x
d2ndUXHJXrRsgXi+624DbCOqiGYw3Ielgx8sQXEZA7sH50mL1hR5hfEOffnvyw4u
vjrI49XEDVLkZTNbZ4cnNN2UPj5u+HQldkWb1kRDCDpgAHfgEPI9eOV/kxR9vRUm
c1E6q4IFNS4oPVEFcbcf0IRrX9ycqUIc56hCfMYAJggwStIMP7x81xf8fZbyFNMw
66X5JH7987lNd1HmBwiGqjq/vpx1Bas2DqSZ9rya3CRSs09L8fZR1tFIY5eeut9M
/6IRZKFGut+l+hYTNFHqrkLrX9EufzLugl0TRQFHmnbJ42CCn1++7z96LjVrowP6
mHARMo2fQofngG0O1DA3DwcP4Al6fNbM6lV4M+t3IaKqP/a6cUSfzuKktH3SsDvU
+udEcleTf4ONedzEKgoDLmV2yGa2AskynxNbXj13NOSXm/kd6EClZuZLH1AmXpGX
d4LQkvlH4v+17SRtARu64dgeBgeFDqXVAEG69x++0u7D6LWhu2LEhjoVwf0JVQ9n
aDKewIL0UWY2LsnpNRgRFmReFNa8L3iRsYqS+c9bE7+VBMnuxDwWMmLmuT5aKFhq
OUmK01QlBwOfvSg8+O4U0Vh2PNz44d64DzyYNDNW0YBIRWphM1kBWha/id6v0D7S
B8IIUHtPF7C3Ceur3j1pia4C/hcU860cAXUp4oFytBEV9hU7EB1Sjv4z2Dj0yxXO
hINe7WURNhBJRw/SoIVSg1Wk6LiKf93OBuOcLYDdWagD+5rdEq2Q1LRowC13kzNf
nsQbJUD78SNJSOvruHUO9AuieutMnxT6+YmyRVcCXRIY7d5dJ7EYb6cH0e/gfbhq
PnQ4/pLWiQZ+yEXLLYw2taos6gulltXZQ+Jl97tcaDuH9oGnVvCYXLvRIK6u0l6I
KL3sncBWlVVn46Su8BZoimyGvvwqLtZU8jB+5yjwj6Y2rOXO6MvDGWWSMq4rF1n4
mjVYv/EvPn7o31kuEkCVPDWHAYAydNIdZ6oVnRj/seCjBZQqJxeauVZDT33n/P20
ec4ukc2T+U7gkqOqEXj5G5+r6wNx3UwuF2OM6KXdw9M5i/FcyRxZBxFambvSezRR
u3GL8kY+oVNdU2XK0HKlDTV08QqmpB60++7JwkdQHaY7Y20o0zbZ2JlknBE0zm6C
KPC1Hm4bD+FUKAv0+mlEdNvPfrVpenNRMDgV9HoxPS64HB0Yc0ni95EUBR+2+CXa
2gogBirzWI1HJxfxuOfj0p2KjS2zBP7hZpcVKpJVdC1qDBkuGw9/YQotePja9I/h
Zjxa9i2MGrzoo2Ft4pKB6cAyQ6D3qdgpmo47Kr5OqwQoTNt2VBei/+/jjtfRlZbm
4w7oQVPq/gxrNdHJ6MBqAqKC9ee0LQH4QLHMGPGtjxRMFIGoQBKdEGH/fEd0MjSX
G24uUbTpi/xV/nYZhAB4S0pLnfNi1EpX0kv8wI405Ih19oex56BhjEzfYKq3DBK5
b+rpqCcQ+92Wk8i3WHDbvoLkLM7qiYO5ztm7+Xa1lU51xWPLTNo0dpB76HVGurmE
eEjTcXcPu3hYtPtda9YNuxqTxxK2bcNWArVaqAdozL4e6VQS8tvrfgbSTNMRxLD8
6JK9Wsu7y97JhCk+awE2fkY1hBrYCaXPqNgD25TCysXjlwS3ieGJ0ZESLshWtABK
iDihdiWKC+oyKWd9sfNeS5as+23D4in3XymrjJOuczAhlkje0DPYGKx4E18sAsml
qu9d9el/nflVSK13hIZdG0gX7nEAziH0UComVqnQOHzAgUlhlumemPPimz+//ldf
MZ9j3l6zGX4H8C7ISUtnG9kXfEp85846+u6DbuCCpS32azBb2Qt5aErrUsBG71Of
NPtbNbFyAz9hJ7CZhFOox47RoVktoQeM/ieHXI7vvM/eDYZ9Q4MCjdmRMlvNkC00
5bHraIs6WGhmvWdi/LQrXjGc6axcFYhWSqaKNPLvvVnPoQqc8lKpgh7ohKQtUIxh
UQnG0l7X1l1oXgc7+iHs9jCEonybBhJr7BMTAS/20JvJIdTivWdDLODnBRE4bqb5
xp02aopo8AbDABqbe5X/SsRlNtJjzg12iY9aL3VtbNoP5L9YQB4iRLc9fmzkdKMM
dUr/rWdbJdPGdFBjwM/qzKq+1dZZRIj+OSwua4yhzz+CoqlCfl8XZ0PP0l65dlDR
kmfLzUiTm48dnFUCZJm/ChpO1raU/wxAGUSJRPjjRS/0sQC5yPdvMYw3CpyXTvBQ
I7u9apiAbu+E8eVeecWDzj9HInTnMBoSnOd8uqOnsG0RyImy+4A7DIfsgqcYjN4l
XVOJjCBk4ZZfEEk4pKpNpJLg3cIR/+E30MiQiFOesI2TloT/MuV1khj/lC4K1b/I
T2YpPT4jRFawe+HLWEU2AnyXenMrgNP6gBzK+5hh2+pG+N42cTvy3AIjt9bYHTsJ
X/WlwyHw5UW24aLS6V+Z8lOUi4OWKarPerZgLdwicws2inUVv0zd7LfP6UYofYlI
tad6SdwurYIxfwU+p5C8wAnvbcbvBwX6P1uPmAQhyw45mUCXUAf/5gePj8ZbSxgg
TSZbfAp14xaNZru9BOdH2sw7NkbpQ5YAwL5in7T2ZEB1WtLpH9/MlbioGzQ9x3I7
UH1vGDirHefJJjzG/83IHqOtt5+HsSBMxmu4kPr3APAVeCLYV5HpzPgz4itq2lSY
SvVkjA069ZUPydmyk7Fb+WkVeUCbmUCstmrxSOL+qp7mSH4nr0P9A67zRlQP8J8W
WF778GcFTHe3iJ2AnxQuQ4uIAHqbNAOACGLeAtLZPTl/lo9jTpIqJeoY5dt7ZcQv
Wbhyn4BY4xFEsl/nlQO2xnIkliYGGEogp54f7hNba6Fup586gn2Me8KYXOA7tJuF
UlLFNb5bbS7zcD+TZN13lsnNTo2A744LTqKEHt2Lr/5JWAbeQlTjF9uT9o5fxCMS
KsksPDqd15Yb5EgfJ8DsT0cIevUBx6cviNxIG0WXW3rzW2UITrIAJB9/GZmqsgly
58fXYC6FkBM96BGkWDXMc1UJdMuoduDKuygcGT4gPB6CKTuhQGz50FeZuhJ9xwMi
Xhd6QMfxPzkryX4bLjBQH0Yrr4Gb4Hc10cE7aojv+vnFfvubZKjTTl94TWrzBBxB
Npt2LWRg757a8yEz+Tpgna2X6z4osZ4FeY7XgMT9d21BcW6TMxYeLcVocxrcmIRR
PNSShKSAttDQCcHSde83GC/IfvMu99vcrNniCzieHticAGwtwVjEmsBu7Da0yoZL
C1yZi4kVVPYZrtGfLqy0TazKjle71iEhp9I74UC9t1WkJIHcXxPELvy1IwySunG1
81QAk81NBEeLt6B36p59CpZVSnjK6d0yN9opL3qFYgPa6RNyAB2kVHH2HEKCpjO1
Ls8th0mvpZtRS+/YyIoHX6UC0LhF0vV/XV1odr4TumCbzwaHIvMygEt2PAKqQvW7
FiKDa0c5FOQQm9Vk7choiPnLRdabWaodJ70L0V4du9l69nA1SyOWYkAz9WZudZVE
SnI3BYcEr7z6Kj52M7XOPiS4VKNT5mF+3OW1pc9s3l1EC1Y3LdnbWtkUxMU1f7fj
1brtkZl9cGQdFVKUoF+cPHaj9LKoNG/aBP9U474ZRW9emUZ4MeAuhkIfbvepMMKv
3VM+OVGmUIFWnQTHtJy0dMPaMEPda1SOt1FxIoCiwnTJEgEVHOHVoK6y/ryZviQx
D2atep9LZepbTau4KcpZcHO2k6y/H8rHe9TMdgiihoIGiLySg3bYYE8cpRyxWUOM
FzQ8OIDiySyl9xcY9xrd71WfXacdw5PpLFNStvpOc37ao7MaRdVHM4qYLkKzSilo
gcDCiL+dNZRz54cm8hXbHbLBZ8IRqo3JBwabjBqmP0naYUti0h2N8zoCRJZWG7rO
1xgDyPJE1F3xkFvKptz8aN/cZBqzS3YhIEZ0eBE/ZJQixrOoFnEQSVpLcK7DPvW+
wCqpFAEI6o+dlNxzK4NKV16JuhRT1gg68Ms3GF6XlJJCGmgsT8Ps4puasWVXSEQ+
29pHUojdgDWtu/EPXj1SPfmrGFAFLYZTbLPrHYQhqWVkJjroTzY6v/S7G+wFyXNS
TevTrmElXyHKvUwyOltFNajgYKV7GicKUJOJMgSj4cAWw4Wz6x6Uo+0z5fc163ca
1D0JTPBoCU3sPJgLdxwMhJJVeNgsuJuFu7EzFOcixGG7YMO5phZg/VpeuVirEIH6
NprehfWNoXMrbI9+iBclDo31SwP215dkda/8BRxL+4xBNQbtmcuc1lPGxDXtlrhD
LKOLMvxIpmh8LohHW2U0fONTuyB3BVF0vOMUNbXEDTPRkM4IWDl6EnEkTyoz3V59
3CELdCGOYIVTBrcVk2WZe4Qmg0w0v2brrN4gs+emtpAUt4HPv6lxafF3sFEEZ/Hl
sehWDeeD+AvMP/lntj6+zUTqdksWXUzmDZGrF8Y1kGQcuiJLCOA6Rg9XfljuhMNb
yhb+hlpW3Re/gH4/7xu7+prWF2b4Xxh0Tc9ipCYBbSsga8BdH2d08JG+U3Q3h/E4
DTCw74lc1mXcgeP0522ahURrRAk1nYlubAgJRpZrs3vADWGTs52tRnqTgvsJG61b
PesWizfLKlU4D5s4MbDhvGYvC//liOaVKKCeZxVX9i1EStEDTL7c+Up4JryUXccO
EUZYl7v7hudcd3kZqoFGupyESALzI2Agitxu1ZcolPTLW5bTr2/SDMyn2wIEKVBS
mB0ReR+6hXdTJ/rMMdFTIKuVf91wJ7V27LATe5066fIH4iHvTeQBe2Mr3Xq5UnJF
Yrp33lSkB62o4Yk5VKY3tTTGb8UxOlHMknKgfr3ta8W7w691AAb+67cgbLNHfzSI
Mp9473VVssJkuJc5PpKkIW2nVfriJj2dwy5hsyDt3N1Z44/+7JoxSIcm8K8u3BeG
SR3hDjCLrrw4tm1RkjSLNNkkKl1f8hqgVfYT97AUNOAZ/j4RN/tXmyR1x79s72Wg
CVepwLYhLnmbzVZ4oJmfQerZQT/aqixmoDEl9sEOXsQybgZSKjKVJKCryLw4S+mi
EphiXpFrm15LrTT9XGOD0RfUD+LfQU74JU+KbWvmlFtdHJVc+dFdlXIbYp4qu45d
DF7EPu41r9jA03BqZ9/HRKLl+m0qiLVEITZTV5ILkaL37cZWBBzazxlR113qgtya
P5JLLPa7CaaaCbPe6GDyGszdpPsnGl5nLHd8H96KPy2vWBhYN8guZhtUYD4frOeN
m8kpQluanqEu803NHerRauRRF8Um9yqxBbQbWmnlj4VGj4dJ5XRGGl96rLyOlhS5
++wW0cW52pumW2iy+JsCMXCfOv9cOTswUFxB20gfp3dXt89TwoeHZ/8SBj819E/9
biYkEm8Gt27eV/whCeQ78jvC5DxVsLj3HM/UQkGiHkg6/AeJi9gwwdGYNutrjva1
292fAoSy/WfnrKArn25JGDf37lsEL/jar3vk5g3BtcstbauACIOiT44ZczLEiHxr
wL+qbhVeDzB53mFNTS23RoU5qThy5rOVnNxk2gExQuNisBm8W8QwiGQAjfrJ9QBN
WmpGfD0oO/L2NG0K/dWy0m1ArdUEdUvXA66MhHx6nDrae80qHa6jhroY6yATTCXJ
yZCDtYoqRKy+w+a63spG8VuoEKGdOulIpDWiPxFN12uEJ5ADKekIjv6/KKfVxIgM
zQikq2WzxmBF2yB6j/1Qu1fgr5zqCS9Ovo8jEMeCLIiuOwXfq4Gn6WX1AFqxKSJ6
CviHtDkRY1Z5w9KbLuVkL+DvNExwsrLYzY0ZpeiYBT+MJfdRfjvOyXEZGarkHYhK
aZajzVmuXH4DWW0aHlMl+mRWacqA6p8Vy1n1VbfS4qlhwRobMJvLtDN6AjiQk9QE
jZXY9J7J8mj0ucpLKTbfC1DAkQ/JrwwURw631zlqlnn2CVMl9lKwUkG02oy+KzU0
6IjDavpJZdHD1eKyp+E7JLv/ZKwk1ASroSYbp7dz5KRvChUDLfzepcz5EU69LiHY
8CSG9lDTe6BaLJKf8mzv4VpjkbTJbch1qFGeq6a+k6JqEiGvWZUTkwIEnsPLF5f6
4dzHhwCrT/tInEKznI+J5PqpSxTO4ITAnQcOYqKC29KS/4yK0/c0+Icz8Eo6Lp9e
MYDQ1gedw1l3WBfCYmIByC2Ngw9YZRjKZ0vVTd8uxrP+aF6reSF+1kABjqAC+YnM
AMuUCzK4P2pSEFvfD0BhkIkSq3P148+VYMe2K1yz5O3ifSlGHYe4b2fTsFtevS0i
thEi0QQY64+5udRUittInnfmpEiZCcFfSTFC11NpLdXgP9egTOJOe/pWeObilrWe
+s7Mxml0rxAexGMOQqX4ZWdW/Ju0727YcEtMZLXVjfwKeRiey+iNn0ylEtHx3tOs
X/rmqgebuQ+cI2mUtH3oPY1Q5dN1mvFXVppuB3RXmPYeM3ZuDwK9zdG8eHzVwOkV
+mDwmo1yaxV66ovyUuPrFlLYr6qgxhcM+NU/z5xncFEdOQXEtrKteF7P4536Dgrt
vWh8Nwl7m0zsFSkKz8kkBsw1WQLqnsXhlGeAKzlxDkFHvCD8CWwymVgSeWoIKxMR
HjsbJMbBcYSBHWMOzfiH200lAVknOG3rZuAF6oojkqp7PlQRx4hZfpBTMgYnckz+
KilhkCOeObG32cndCDd5233O0FlOIkSPz1WabEyKxCUcyXALfV0sSnkETGkPqcvk
iK/gUK1PVy+EXWkFIjjAerHjBUfqMzJuzXwM59VAVfjeO5mGyZdbAx5pq4wsefZY
+WAHyjul78StpSw2sXXaXlWsziuRudPSpZE9WVe15adM1xp+AaRJ+s4O+AVDU3aY
n+WjBw7HpEKLrlpFppCuwdmvXzq9rqf0yec+KDPLaLLCMmGj2RcjaC4E2KPugppF
PthnBjMEqYTM4ae1Xxz/wxTI/HbYoqOwCbLPsrv/4Q2L2inwNkGNmmIf+n4ukXJu
JZ7ogGTLDuMhP9ySfr+Zp9BNjW0Ej7IG2mnuPSZjVRXqsaAEA6o/ZxCaGNNTLFAN
0BKAXJG/u0dibSpTe0URcwQVo+8domwjY0ThtPC2d2ya3UNiurkarBLcj4Yix8Si
vcFBT2WnzjYlxrCDPgSOBWZYj7LXG2uD/Zm162UTmOK9RMAbC4pboel+fdmmQM4S
pXU2Khp8vLOwQvlpdF2yWnsHCN0YZDkpC9m2qMyl3kPuZQGkJNB7YmUhyMWXJhwj
Qmd57WO5fGEkHUiwgUJHiF9lpwwByt2bAFQAAV1r5XL+Jona08rWjDZYHMSq/azz
dFk0GZwsNkW/OyETYyN2Hk2m1s3P9vpqGWp9SBolBCjhojm2EZaxoNhWBDSK4Vnc
gglWylL0jwhUxU91lbqXafM8iAIJNbh/0APmRaYlBiFVrwIS2DJ7LwbkXzdXXptQ
UEvVk9tzSqqGtJaqkXDv+h5pkr5gTrA8dsapJou6p00xAqHXJKrFMNV/BFT94xJ9
RRXxPKa08p6pp3TkEmlA666wrivLPG1yNvXc3B3GxZ+LDSoQBvV22pTF5zNDxyUX
4Qp3DbGHgSo/rkrsieindnZZKK8k7c3463MIm3aYVaEJDAxf+xUCWJWZQbN6PVAL
lUFneprkhew4NsBDRsgBLZRGuwto7sIANwjWQBJ8b8dhK8v/xRMHTW6qEkhPcTGh
zfZyErJyI/auX1ee0MZgoQMkxeBxEMaI2+HAE3/ssXgfxSN+CFss6Crsv+dW/dO9
AtyjGsFS8YVgHWNsWIgh8QDITiOfafB1IPtWtBO+P6M79VbwdFqNFAIKYhkcNToY
MnU3xiZlRaODSRaLDO7SW5V9AwrLgbVZuU+GHnSkEO1wnVJE2n/xe4Tj2Ia6vmuf
Rp9S2O3ee5wkb8w1SnNmiOMJquqCtC3oSDwkIFcHURard1TNRl2WW8AxmJBc9w8y
ro+riZUMbT0uLM2IktkmanKvov2JZu7TWHfq9u0DFYQ9tW13/SW0YlTpBchI8Haq
awZa855EFVLpwKgoEGZh0vyO9xgdS1qKseKRYW9TqMH3Et301aQfKOGteHDSKNVi
zI3hONZ9SulZGFBxikcnFA68zJW2vxVAwWVw5WonHYOyD+rPrc+u6NbDGQ73xlvg
SAHhhNS7m+4bTMyX2fXlHcGgkLP9L+gpVo+NCLT+cszaqgtn3Zv/PL2ar/+9PemR
TO61PX0CinHCzvjCtaA+gXDlq5+BtNkVmCG5+4Le0wn3pbfhTv/r0UjYeRQlGjK9
/UuzLfTeAGaxZMcayezIWQSbj5vqSg90iJmxdTFtXRJKdMIQ5YvpSicfRXoCr7po
Fb/wf0WyN3BVoUXEmU9JaIKXd2Ju2DKZYW1A+jkhT5iwN9BUFGRc5N+lYsEuJ5qH
AghCXhISmo/8tAOGRu3M/giOxFKoK3ilC1CYEWP5/6BobiWfdeFSxHKMXqpZnM+x
6Nmyz1b8XCiluz//ug60qMr13V6oy1LOwcKmLi7SnHoFGdluVbjd/ytjfkpgXVFR
dz1MMLD0gCRk4CwYlKdCKqfTc7akfDVcsO/2ZcN99TBDZW7UDUGXXju3jmgjxLRq
WV0AOeUqn5Ymnnll9um9BkwLZwZ8nQ0oD24m55KlY+n+5ZHI7GfIQ2io36wUymaB
lCUTh5z49COaaXS8OPIncz1rZ0njaK5lw8SnXtvqH0ReLkrKmWzO3SKppoLU7yqy
khPb1XxqGYPjLsXOi5c0wNfQS1hGG2WWBgq+m6zdMZdLtUSG7DRJSTCj1hiQILQa
dQiCSaZhFekS4oIftBQ2Ai5Wk3P01iN3WyjIwgvG9GHrpgr3eTzzUAzJ7xwA8syT
rpmxke/PWVEFfX8dBthJOmI+DXz2ek1IkSUb32Ij9sa+socm4E4QbXRoTlfSUZck
BcDohNJTrJDJgJyGy2GeWj+SZIxa+FLntUfAwfngTBa652HynVTL4TNXPr9mmz3B
ANhv0Ji1AQSos2roQwWbbpWTm+HV+JHMii2FoDrZZEefjPcHVCO9GQEtNf+fm5F9
IsXacZAEOSAxQjLGpkYH+kM8cGwpKYUEu36uZkjO52HRjtPkfgIy5VrZI0iXiQtH
8fa/UtjONvcaLkARDpO7N3RnfHCQVRVG7NizYcTHOa/3RmSkXZq3MRG9ZoZjul4u
EgEVEAbsMUgQiHNRsjKvc2hywrQG5DejhDs8bWROa/gXd5jd94asRY71XEQPYpaS
YjSg1kFNWcRyd8nfq610H2o2tkUOEjLM+bPCZDR/+hRdEgrF52//wA9JSb6U3T1V
1rrSJGy26+QxWAx0Iaqwd8iaE3leOy4fn4igm+FmDpjbElWakD8309IUYub1q8GM
JE844F4PllWe/zBVo9k6nyZ6KTXZMv/ObnAFC7u7LoRT8fFeger04tzKeaWinNdx
akaBQwommob5cq0DsUfwRJS6jZcpqd0H80WH1x1f9I6pkRPha66BS+GUkZrpF4Ju
BopQqn/W7tuMlzUUSJAw58fFfec8YN6TpVtP3jU+sK/66lhbqRVQR4tLgNcvxuTz
/Of0NpHuf5Q2uLoBXmt8iGHk01lso77qFRgZr0bznHA9kfB2TD1Es8CHLQ2g/ujr
aa4PLawmou+RIQTF9A2Z3LtziBPwVwCrihKRAVmuI7UYKg4qlQmPS0HfXC/s3mmU
99H3Hdt13WIhKGwkh+SC3JdwQ8Yl0ifH34QRjuXx+0YSMMkYZAmgtnP1D5zMAsCa
+Q1WkZ7VjdaSOpv1ia7T4mffFMIFXmOnD/nt1i37ik86PzIgW9cS3QNwziNdObcM
TOgISDr92TOqVjpvJqUD2B+Vwr99XU+piPAJPnrEzQm8BeLHqxyHklat57f3BLjw
wwKog8RRd4XmNlNQqxFax6/WrL4OX7kG8Hx73oEB88ouLyoaGWSttkIUnM0ENaUy
qSgvClTcqY4P4VkKRL1f8wp3cGzD1Quvj2HP2Rn4iJLBjKbbUFyoGqbVRcKmIdzc
g2eZAIEb7sDN8AjZCz+8GCjkQ7EMZ5p+OqBjJGKKYMmjOd0kaqLdBzkJoTQHUkqv
4xkw/0hOFI2sz+FeZR9xbmho62PUikCkMyTwPZSneAQm6MBUFBKxsJ5BLRFcsDf9
MCB4MT5ACnwlb6sXNDUHRJX3DdI39hifFzTL5K7xN54lP6aaVKKmWk5J+AZvpq8y
wuzIykYM9ODGwKe8q44pPxqcdSbPRxZf35TVFZ/7700QHbWBpG5LxnsT2BWVISoC
2tEQqzJlfr0cXfIrwHuZPMuStiHsJSt6iuZcxkqXj5XP7J+otgnWzpSdAE2F/8ft
KRSgmgKtfLPd5Q/fNZ/y82pjPJQyYmH9Wa9Ou/yCwvD9wvSkbMVQoLha2KrMHy4Q
GR5pZjNoo8ix9ViP5VcD3p+X3aCQ2ev8gMMouB45DhAkUAAJg7KvpD11C+yZhs2a
WAPmOjk+Oq2/EvpNlpA7Yg49fPxahM4WiP9Ri2DVM4HvZXc3n83nHYdTQhRbS5Xv
j615uwojzUVlyoS9D8cGCt6ABwhTC2zFHj4kXfZzaBn9mVIEqCMveY2DV3ERXJhC
neeR4T2kY/wsutzbtgBdgkJ8NA5ZkJCV2/IrnAkK2KKe99ijBdyKIKztmIoMZP6G
ybb+hn/WYnBHuZWFWVd8thvU1Eo6R2VnST4+p8PHZJCMWWEOlY8Zfsl8rNYqfwsB
eMeMjeJKC3tsZb/SR9z5ABFtoaKT2imMASGMh+Mkrf6vQTmxSqEetV52av9NZEij
T7KGiGGCQoVhhc0z9UIq21fzU51ncUEbkE0gFvrc4A+ZEfv0YV6FXitlN/ZBSgss
0gloumprw+pZ6T4wYHUH9Laowd2z4SWsu8VpTcyWBZo3mAka+djTjNN3awcd1YsS
zlY+fu/948YDNSq3xbuuJtdApbMwOoeW717bPFv1V5tmzf/CY0fKiPweWE7hL/iY
/VJiPv5KhbxtOTdlbhuYR0eiAOoS2xIhO4/TJULnR1xxmUKtXiUKK4PyYXiYI1mh
a7sp5RopbbnuIq1EdWbVSXDV1kXdPc+PRetu18+Jh3jmtkP/8l4ONCg3Qpm6Dcfa
FA0er2t7Ix17FiBJ81aMRGermXm+D3SCQtU4G0fPMd/4O6z+SrcL5KrF4cC9Bq8P
lMMU/ZcvaJ4prdopyy+GtOCIl/kUuo/H4tHrf5iWRMKHS5GoS6PreCYSF7yZZMU+
PwKGfkwbqAkyh60tEtUEHYDf4Bdg1bLKWGG4gcvl/oZ6uirLxMfASAQrt3wNQQ9Z
OcqXK7uMKVxwAseDBHGndIVAzUp7/JtaJ3DSaLXng3PUfH5Z0V5HzYqE6XeKdbZ9
25HbHmgM4nC3oU2Yqx65Tom++HWWSHD1A2As1y2bnMljX8dulsIuEvwk4eyztEgI
qbzR/hxbgELOuvfLUxAa+OeoskMhuyf9fdnx20fYkSF0J3cX0CTvPzq20CebHuA9
NB3owr6Kr5Dnz8p5P0c5miEBYtgJsaZo0F+GHHksN7otmYfr3Pk2zeY/Cxv+HAvd
37aKhVJ6vMN1DhhDo8SiiO6K9vHHF7f04r/H1PE9YuMn2TW7nGjGiCqkA1nnk65Z
Co1cuDbrTf3vTY615UP47FXCoICo42IPxkzkKyTl3Ypd5j7a8TqHVs5Q9DPBJW/y
er95D0R47kfEatIX5vpSGREabpeVZCyWNWGM8dT/grataINlW4GA82+yD6fc7ZHi
XYqIJgElOJ9/zUU10DNSvo61FvHZ564Ni5inRgXwSeAtlgsrVt+yYUoGQanuIvdO
hEv/pSysAhTS5YJBT+NehuTpw4uHR4nePpPn4rfY+0oqlDqJ7ipqNK+dx+XzexFC
1Rd2s3tej5uU/l3+trYc7oG74LfHmrJnWRg+n+gMxqwNtwrajdD39x6pyjypMA1M
K26QIFQCorM7jv0a/VxYERWdnUDBWZPcpshl37YPfAEQcxW9V0XzZNwm4QjPf5l4
8m0QGLifqFWRibimRumHP9hxW7E54Oy901fysAJ+S30oztHRU5f2mgjbERu43b6c
iRqd7K9IfAgmI7uaYqMjrss9er97dUcbvNGIghIXxRnGRq3Lb1NU/FuizNxCM1/+
nyLcs9SjDLU9KOFdNRjtO2lhOsImkbcLdNYSoSjSnGCjhnvsR1RVpuGhHkdf1ue+
bgNLgQ0Jhi6Evf2ARVytnfnEEIH7BCOeQxjT2wQV+XA9Cvsgvq7j5mhji/3gvvJ3
S97W4ikhK5TPYyXSGHhT+1BKIc6LPW8bORzAjaJpDvQBLesAEr6UsxvSWA98c1FB
tUK2ecI+WB3MjxpjYdcs+6ILD1dv3jkmVFWFE5MI3/Ykfx20CyeaR0cjrx9lVgki
BJaWTVoiBE2ickZTDh1GVOMryo/Tmev/F3iY4ND65i1b1/MTmwXqtfSm7oP+orjv
gr+FjfyhfysX8GcC2aq+OE+fGxn5rj74MotKXzhzSYaj3j3WTj/7vFSFMnauL/K2
A+nMFKucsTSPmO7wRqxatnbbiC4DU3ZhZ1Ct6AHKGyOts3M8Bz50B7/+J9zO6fKv
puTwaXIZBQgtSKHmpOIPXPd/oryKePJDWqri+4PDFW87S0vInDPn4VccGju+Jl+X
hkgmUp3/ESwVL2N7tO3LarAJCF8Qmpwl1oWgta5L6v1scToKP3SLTBsAkCMwnblT
/LTeGBnK/zHu/uirm/9OD34MUJlM+S8ZtVXUPWS0OHSRvHkiKuMnjGwwYCa3FNL+
o6I8U4Di7emJTHLe6FuRYtditIx+/uSZAMwpwhLdJScvi1bBq8C2Z7JwjZjcEhXm
UogCrzmV3tNT4bDRojt4UMlTT6mXrNjhyvTHGTQ/ywNfG0DImOtLwkJbPAeq+t3m
bsC+HoeaGscXkpoPzieb6srA+/Qq/oMCEV69EW0Z8v+JByRPYeahgW/LYnOBvvpi
VPEnLQBsp1A4633RoN8tyYqukoy5lL4NlDtFmoyjIv+/rRxE1y7QCYnColA6CncA
KRxHmgm0vBb2KaaeD+YKf2ePUNFjmcB4aBr80bPg/KVe4K92edJpfXJ+6lVOlF+j
G9+Yq4nYbIgOa51/8E2UoO7CNviMiD151vhVnwPH5niEsXJEacDDGsSX8ECFqy67
kvsvEx6MJQil9z+NEyqvFICMzVgaMThiMHaVLKA8BfWCfwTqnNFPTB7CXXQvR7Uh
jgnWLAOw4nD2Kqft0scZnPvXOzgJdkbK6aZqLxF0lcePH90yedjDaynDG220EQi2
paEwQ+b6BXPKJOTTlS658mos29Iicimj3zyx3sspXSczkJ6OYMcZzyM6t1ADIbzv
dI9a8M+qQu6QJtHnfRMQje5ys4V3SWZiEcwLBPIpdd05opZVEfLCVa8iyKeNZYL3
pXJKdRdRPMM7Yx/X10yK1wqvEHFeIIOhM/UvLn5zo+BH3FJE8XSvUdu/YexhNXx0
B2ANnr5CDhv5F8JJV2hbJarn36jWHhpn9vFGteGpWYLpp7D7y7MnJzEzwrK31Jtd
rAv/NCTuhyAzw0GapwNaAMlVmKu7MzDrXsdfKOHh0Ak6BjX6iMHYY6h9mTWVBL8L
1ulGWG9iS8oB69/kQ+9w2xkoe3JrrKsszNzPctYrp2TNcfPCB9ZHnURJKAVQHBVS
F5Do9+IWbcjS4di5ThRSHdWaCZOVCEzuEtXDNuhjBrGn+WJynzdi9IvUlxsfgRlt
/szvPc7GGasxEL53NIxHCsRpVrMyagMYiB47L3AntrUOnnLejVofbCQN40NgHVk6
XvVomxvLKH1WCP9bSaFqKjkvt/M9SoIePJHcvjYhXuwYIYCYqHhefE/sxhpydywl
IdeBfFEoEyc3qnKsYUMORo3ILpQTxuGY14J6Yoy3MQ0oo7IDFa260Da14A0arCrS
bcOrWcO+Pt12fx2+sNmWisdVcZ8trWG4409WePjLbpunyNhLYY+EaYAEhnJ+mibG
f2cbp+FssUS5QeoSYkC2OKJsK8IRTngY84bau6mR1SvgKYYafMIf1HGpkp0H2fsO
iTY5WGLiskQCAaVTneGs9Gu2m4CJS8dPuTTlxzOLVncZYDjjrChiEyWdUsHFFJA/
V9l4r3k3hd0PZbT2cMe6OFdluN1tVa5gWs33KigDwsq8nPNKnLS0lys/u+1CoctI
F++Y2uB3Qs2mW9rFlN0Nu4DRWRfX5itHW6VTycScHEJYM/XS+v0kZIIeiFWFZK3+
2Ni4P7ZY1XvaBg5IoEPvW9kSLrVjA/G7/T4v7Q+N+j6S3r8cLyNcborNMxZxp+ky
C1FBgFpYH+dJqCvI+O3BsJZzRxThRWPKSL+U4UrC3wYBlyTNPFetzFgphC06NfBi
kd6DwCWwXrBnGC91I5vobJxYkVJG2aqEiIE/ub1Ja4aGlf82aym4UNBt0Xw4u0Yn
02xsuGiRgaxse9Kbl4k9m7xryBhWT/h9JT0KRmP+LwDL8G6OyL6FaGhSrwppnnsj
8M+9IF9EIBafb5N75VrM4qU9ldlJI6I7AAYgU7DvGOBvx034TK1TxoLXILdlqSjJ
slIFua4/sa58UlhiV2GYYoQE4pq5I28qPLY+7cUJMaIBPBVkn2MMyytA+koMfQAx
9f1LM+0KHXelw4bh5RcZp4a7JVI/4oTA/QlZZfyrGRt4k2fLcVLhQIhoFSepdShs
0ODm52bgR4aEGU82DI1GagBsY6eTj4xbl3u7PnZLirJKeGoacJL4/53GAPc9myAo
0q53qSg7BmLoYj8Q/U7k5Bo02FboZhqzHuU5F0B1jLBqSz0BY6+h47BaF2hnP8cR
XT4HQAVBwn3jBwv9JSJVGB6dd5cF5bMDiGF+TZ+ugklr3aNCOYyX2Kizgy/wqwRg
COMVwiARq9Zb36OKNNXWNxPsxXDrUkPTzGBTr+SJLDmAjubBuCrkrqdetVbrWSqj
9NueserlT61qXIW67nvQ0DRRPyBctGpPJ/qJTuN53rQ6cASmL7AMdzGiQVv8GElA
P6p2KaB/x/7V6wVhDer+O4+oJYGD4wpRCFeXQOA+p4c+oNry2LU1yEBeTQwiN37c
BjrsHLk+YwvgNqE3+C/PS3PnXplkCquDALj6XR60Wl1xiexcvWIIleNvWqCFRlyx
Isi4W2bMIo9eacDQVZsrBb+I4Kx9I1hzpj3QBIi0d/5HvrQ11ljdkhKu61ZEZ5pP
yPT+SKxVz2dRxzzGHQv0tJ7jPXhpaHOR7kVJQYFcnMbvxTQQbKA2JiLxzEi8Ggph
H44taRUp71bgjPdj4Y/PuZTcOLp55b6dQ+RDBHnH1D0m1PU/6I+GWy+LNK2cSQXz
MXVb3e8UHUmsumB5iyhU8ANbzrVrTGAa1d4g5bqRMM8Xr57DY9edSReBw1yT5c+S
33xOqorCNNNZOKBQpXTpSBDtyxEZma48aAZ3iX7oDayYRAGn4XJHXi2LVUGP1Grb
7+f32TKS2PazomREoLw1CIjhuzV+J06ZVoTb3KULA0UP0kR2OEXVW5mkoCKYYPn5
gLiW7qnWscr0HSPYGlBOxVQZuY7XFedoRTME9vvqL6bcBe3Dl2YfQUP04GgGywRH
YICO2yToD9KDMQPsuVkpY8HdS7frYZ1n9t6F5IxtiDI0PngYCTiD6OUKHLEalRJD
bhmzBGKW9L85YV5ubbkNPyzOZVuOpuM52JQxbYBxWDFsVft85na9LZhUQKtE4/uz
YLQVUV5ic10iCbcsUV3eN8FrLGIbCfuyBMT9xiJ6LbKR7izjZNKZv/wwIFosOCGl
ozqMZ+0nUPr4lsQcnuAHQHF4jnoSK9UTK/16bHXEtQxTplJdas3gv+JKQDIHPWuv
Eh2YQ9Y/wgAtXKwHsQJS5dMFpEWTPOvRKhWkgrfkmM9beZ4KidAtsG3LCJd+WEU2
77H8/iJ2ExCK7Apcaj+Pu2qTZFvaVfN9R9US3vNHdnY77ot/LoGD9qByst0+t2qT
B6I48ksfSXZALDB16qlZ1nwvg5F5M2sObN2WAid5rPohDMZPQVhw32kz6jVLu/K8
N1obSU4pSdMW+yP/QcSxUfsSdE57KeWprl2juLyvu3r8JCuRdmnJfrLAQ1gvy8BN
xB+/zpyugG3R1oYo816Q7/KWVVplmZuEEWDgryHBj+wEx/UwqHykWW+fy1S25h7V
YNPuypeScPYVfCD6ErTOIDDqC2iaAM22C/dzTFGml8OhbNiriU+nT8JdPxJQVnCq
mC8FJlVWh5Pp02dz+6/qMWbYusaGgJ5UMFFrRI1cyl9mwBq3C7OWzOVOOEFiseCc
Far5VTaxdzYukjmZlwoYKsW8/OEQvBf3pTKwR7G0LPM7OA6yh4NcWK5fCZRGhTEJ
XU5nOxBZij9Q3IsK/fU2nNdAb/TV/B4rXdq99iS/VeHoE0IvUlZOSuNSRuiblobh
v2X3p1kAY4yAv8tMiW+B7R9Ze+ekeX2rIMKIl+9GUXirpmMAxLilG7KSaBLTR1eD
h7Zj3TGT6ifJdoCepvkYaXctKbzWM1KRGIX2VHa75SxfrxquUHhT0/7Q/mcw78aJ
g2t9PUA+eDbNONAcgiefYVCRxfU18VhUNU8hRGrvgWGkoYrWcnXO7yf5QiqvGBpS
BjIC8Hxmc60r0yPwuiiHjWBaIsiMzJPRTMk5ZwTjet10Gr+5Ob6xmTZSYszvX/uV
bBJWmHTBIVj06EwAs0XCXISWa2d/KJ7dvy9aEs4KNdOJ2K3Zs0NMSvXcbhBCs4mL
w9tLJmlGLNw8UbZWmMyP8epUVipzldb7bjSR0CrmbQEe1r6bQumEuIz4ADitio68
xPBpjxAKsRPr3RiKOwc/ln5QbAABFdK88CbiFPGcCp1ESozg9GsR1qyRPdonU0gE
thCdEQO2hjtAeH7RymP7I+R2u0K4FDV08Aif80MrNTrOuzt47grJkPl5ePHPaBni
Bs31zBPIY1Yj8pJhA89yDdWwVbt/FebgnRG+7H1lGxnSw5J/VaNt7cLVcx4M0tWc
ydoUXlHAtrfZvlMc8bjTDVRvsO29G+EIW7/Qf1YqghbPNZ76rV2ri/Jz0sjQNK18
MjweaYBH1A2fvWhXS1Vcd2WGx+KzQFeokTXzzu4egEiP+Cv8N9rSguwegHOYMen9
J+Dwjci/GMFbJRv09KEnx8O+UUcSH8flDFSB65pK2opMAIm0JBdMYV4Rhpf7XXDC
Xu0BZIkGzySpYG6nkXXNkWdCL8QlInwUL0LIKYTMNE8pc2VdEVrKAPNCmnIMqG1g
bxgV74V1DkXznuRJ2rF1e+FskDqWVLsRkDT67h/dJ413fDE3q7LsNtaGDycE1EMZ
5AHIy8tgoeOpksB8tPLz63iil+nh1m3VDhsVnytivpEVnQvIR/Pjc3hxRcFdj5w6
gOJ9hERpN9+hIIKdxH0U/AzgHjHcibpA8J5o4C/9XtWVNfi33VIL/VKRljZnRfwr
kNrzfLmq5LvdAiqGorxVGN0OrMCRcIOZsUEkDQ6wTUF/M5P21aaAIGyAg3KDNdOt
qS0snC8PDG0y+31GgKm3mLagq9h0XnxmBgVe2WmHdD/zZlP47DwxQ2uUiguX3l12
keHpXQaVO3raFd/aARFDuHqkHXVhWNcbNtvuiTkOcICGE10BZCgZafCP94YPmBJ5
s9G4XHOLGbpRpCddosEGQIWmNaz8uWh19TXtoPz1uNy7s9xhNpL++21EDRuY+En5
rUxlUtn6MlH6IXCw/Fm/FSk2oRaeD2zm1iEH5P57UpfSrv2ALahmhjAJpfogq8OS
3l2+SfB+USNaQXX86wR9clY3BuilJOinh0N3hQl5lCwy+xP2LeO6BFblUX8WGJAm
6OiKj83YqVq6IAM0YJHRUJcdDT4wdUYavzFU/W77kH8KPk3XndBilBpxTYEw1Syg
A2sCI8yLZN/4gFNLESHqu+rH7deU59L9A+NzuIuZj0DSwAJKa0Ctk+o/kMweySH4
b+lWdL0C6Bsq4ktytyVd6kkHPdFS5eQ1Q0RtvglKy7g/USFJbamKQiUiXmth4gkH
JQr7LrSgyxXfZwMzBoqCUh4b+OntiLkilSci1RaoLD3Jn3kfrdrzOf4oQfYOrPdc
jpe1vfnDZacrZOXeH55yewMFGrtZJPBVg7UGuZY3WZhxMaVF/d4SkXaSUZFo4uQS
NkNdjDP9j7PA3YQstomzk+UAbXhIvFnArlbIwy3s8OLZtvnpPICGPr0E/z2dulfi
1xskEy4dVKw1ZKrSZCvd7vjkUneqVeP19th+qNmoFNKLuVitWIfhJI3HZDzts4pB
CguE7zeSfBPphBaoWQ3C378d5j0MRhoTJGmolfartmdYXBqHESjYntUqOXxy/xLj
bTLOPH/3OKpd9w85OX3Obns4rlshRWZbA0aXHwtauYdMDzaQamavA73nzMgPS5LM
KvdY4By4BNWwE/b+/V3Gj3ion2ehwfF1N2OYctQCXQpRPYxI3XzSMnhdepmtQO9U
WcvBTUgyJY8pwD0kjg5crfmbYwgwrKhVhzw7vaINFWEuG9GVHHCycitFjW5I9DGM
9qk+upvKwpTMO7K30OeYOxpnGv/0cNj1t3IH0z3/YBS9+XUp8saOEcNtMWoGac87
iwkkKlXTB37bFiKgqwVdimn5Uz81Xcr1pnjGv1MZ62s7ubKqGSXlG7ZVQxwnAy8j
3TWvB3ec2wDgvq++tEj1O4lY1qaZD/1ZH7uMEOYpFwtqMZxmVkKA53cGZvcAfZRd
opbeVfn15OD1Xw/8eaI/NZNQa775VUEVJwhz4UW8vTSDwDD82V/xqYt6rpfnJ1AQ
qw0Ck8WJQ2nZNeFRrlkdYylRTPFn71s/TLnsbVijq5shNPtdMjEycy35Y6BcOn9p
1tTn1dAMIYgHiqeilDdXNoSkevAERt9rKzVbryW8ESdejajXqmrDBQRc3PP+pHXM
BjZ8lThV81HctACjgsTOJXtWnAC0WqXfDbNmQ7mNdsuaDwRYX748w0nCnb29i4vN
Nu4aqoRfmUV7fdwfcdN6zdZutImepuTccO6mHkG6569oOweQ/DRQlm84LtteQ3o7
an7UQ9agwQyoIivAiaVB7d6oNVC90/iP+eJdKC/JG4X1J4OcWeTsNWm07TK/B/jp
GyPHWT5tNKdf6j8T6uep9VaITcG6p6TIaxl88jQojGtQ8bMqr9hBxJLYIcfTw8fF
XbyHFwiXIw3D0a6GQBnBP+nId/i2vhwHslRfbYxQKqOke6vuH8xvOAA4/DRLGVbK
w3FeP4DtiZhBHAtC/QEfLpMeP2kIkXRmHrPfIRZt+Pu0W7d/+zU9rEJUrL83QY1y
TDlFh2AU4tb+WhGU4Hmg39RDj/6hwJajAe8g9eO2zSUfMfl+FdLqlzM/hKuhYoG/
uRHH3Zovmka5lEc1Y04zZmq6ifCi/X/zAvpfOxxaycSiZVhLEAnfubrOxmVQlyYf
cYSSIKT8d1gcw7ORSTEab6uUCrD2EWnpUZrXwTQVRbWHR0poW+O8xj7vWxqf1iTE
6TTAGLCeRH6UppNuwgtY2nbW8aAPXD8AjONB+7ZRVqRrz6wyhFmUcz02u5lniGOW
TxKtJmNoQi0ws9RSeXU+5BDjdzls7wk+a85AIs31zrlqUaa454FH9iF81OzHFo8W
vMADMr1hTnBo4ofJLBG0URoOH6finn//qQta5zDhCLnO2JbWhuGbQdAhJWbEoIts
tYc27fo8ox6vVhY1MW7sM9HHEVinIkIdS72/hwX5hP+MilCyTgVfBEYKodBrF4jx
78DWOoM3hECmv7h7jAMnU3aYW4AM5sfNMCfBkR9g/eqKcB13fa8y088jpULbMvr4
+KYe/pHfCN7TYCMr3v5ieJtlm80x49nrZokyr0+gst2C/AARUx3CokbfXGBSS5Ys
YgnkIUz+GWx1Fmk5LeyjRRHOKsWXeBTN7GZ9OInJr66CFrA6RGPVqsPPUEH2nwsa
UEfWdMaSs1f24MfmVQBfRzMDFopJl4/LqxyCh9w2q7MHR4TBlg/GR0mkKis76ffA
oJaGNuShNTdxxGgkSxHbNVz58T3sKMmj6StHw+sLchARQGOW2pR6VcjysY2xg1SF
HyrNShCyQ3POMwhL8JFTi3F857StoqEv4Qk7qYljpCVS5HjSQLZShkWoBibXQJUJ
jibZ0WrbpnHxlGkthcjaQJz8ntzwym2hMW44w3gulEsgJMR9v1tgbdf12i0WdB0I
64owOG09ND26bN2TzcNj7AAID6JeBhs8RRk9fCCbzIy5ulMsR3erBx2R8cKcMGNp
5tcW7+KhivcX7zE9HLcs3/32S65P7NLabBNvK9/t60s/xShbw3cC0lr4hSflHqFm
0LtnSb4/Y7l+LenU02KxgP70nNWTThWQmOoXKMOk/naYTZqKzscJfgpUO+yvx8NU
fdslKHXF2TG+QrL+eLbFN5+FkC3LD7WGHSbLrUxM9w2eXkYnXILIqnKXlUbzbZGO
vD5D2CXgYRSawU5Sa1UQjT8C7eLATO//k9B4h/eKyjsXZxHgcAdhyvzKOcu0Kxxk
c7P4vv89RZvEZlRwJhyitvl5grmicSitD88erDhkPQC5zCkIIO2J0SnTtmrbUxHp
d1V/rtoWuKY3/el9oqs1UvEckx3Zl25Lj1onyErC2Yvd5/OI8+oJciTf8CQDK8xi
TK2rwacXvz9p7HBshd3YUq7TQJzH9ni5P9RjMjdcZ1HtFZCpjVUIyEhl2ta25SlN
FVF3CWH9gQNMnDF02TczdJ6Xo5/yNfDbg4tXrpdc/kPSxVwyROpTGFsBx/6h5TKZ
SHmRpeRG6ULhTdEGx+zA7UX+HU1hx3r5Ylf51Mh3jsWFW2fCvsEK00k82XfgxtyY
SDnO0OlPqtcK4czXTE8Fw4Z06+7TFEpT+zvO+PbuOaXvBwi30a7V3SomTwi+/Zt7
Ea8YB0/NW8DTlkcFOaNAz9BS3HH8aFmm6Mwz5+OuWadMpDmadKH+O9M2eyH2la/n
iEALKJuu8ySx2isnhvIvXsKdZ35KJXGThDf+6c6KtcMDv86u8c+xmEpWZqDRihPN
thqfaBIAi53vBc5296dZxN9wme+zBa+UvmjAcpQZP/vxEJa1ZdYXUBhL9Wm2m0fR
8DrBAVGZJd1YQs6QQLsGq6jCoqqgSL+piCkvzhf98Gyav6PZjG1jDWfFKz3dmkhL
3uTAcGKdAHahqweYoFujZr4HoVZf7WK77T52UZJijieCLiu84NfC7AWJwkTE4KNe
wPqEiXn6eZ+J1RHjuNss90afICvxWzhUAmkkLuBZXvj0yP3rF4CKI4RqiBsQM9W3
N9oP/LroEVKLvKkXKOZzozJ5vroCjo1NehzfN+SzO+XDjqCKW243UZ4bHdKifMNB
KZsnSVoeDpeBLU0Vk4d5G7qtGMjp6x0q8JBEj/mYcdo3jHOGj23dlBbk2pM861v4
+8sd3QMlcB4t5kYkjz/E5o2i6btGzOoU3+/zibXmcKD6W/LC7Uj4aR9rTzEHoV0Y
5uTbdPQ3i6XG3rm6AvJdfaC2Ix9DthZHXyScP3KorNzG2aCBDao9u5Afd61cRMJS
VCfg3us3hONvQbgEpG9V4s9jNFpwC1Uqcz1dusgikvELQ5rkEHBksMNsp6VyAgvI
H1OTNxYSyritiaFoU5sbqAzeK3Dv5NtzJbx7QRoEQsET2H2FNc6mDXiA2SrXar17
cjnvxsSgaIt6JwbjtqLcPItOKsNmJ+kDQg/5MZfXfCuNfBlx4PYLLfoK9076918k
GP27PWGfA/LLv5CZtfuCF3rQBv464Czaigi3IINYQMieT5cHZuJXGSLWXT4rC/YT
KjNUFkYk95nTlwPaWYr40U9574rHUbRvun2rffSGfXeltvWLassw7Z4KQImpLhsZ
iFR7R47BIhWc5TVnMfVtRa0WrtLS7lWtIoY0YuE+ioP0WGFXGquWN/X1HWVIRQY6
65IZ81R9HPUHnJV8qNAlim/R271SuDxwrvE+i2qr41PPrDQJBMUXS1B32GQ/Wmfq
TIa84Nu/hn28hxDsceR99g6RHOOabS3Rlhycr8VKDHG3mcZUkpZ0AR422etkNPBW
w3t2ittl4jZFqVU2Qtcjl27Z7f1uBPnXkg/ag1OXsFoDtgBA1xNBO07/eggxnPw3
qxn43Ly8v5zOQNrzP0Nhbhz4iizaS7Wfrf4hQbQ2vk40YbQaZzWmzsbHbi8TWxmY
1V1uIRAFgbAkXbZE3tOX1ECp4l5M4Cb3fH2jmy3UCsgMdGdjPTY3Aeut6okK1Aej
kcOTqgaYWytpXHZbtEXUPu46Kff7UaqyxtfRd3DoBhEh6hLQUPYFsw7UqJRcvY4V
fIyKK5NMvovvAUiLKJPqLTBQduLkiJ8kOkIUW4I87LcSZEZnIfh+hhT5oaCthdJt
aPvZW1PvvgrWDAHBMCrInHaAXEAqA2PDPPfM+pnu3xDgvQuCW1diUgYXG1DGB0ov
3ywABsr+RJFpqdsgengmKcrX/JWzdKfuvCBIdBmXt+N9NlZAmKL7spVsYaN70rJ6
yLm6chOn9CeJq2su7ontpNnaItOUOsgfqLx3U2ilAt8WSEu1QdqGU+O0ZcEMcYRw
K5ffrVBTeutL/cI8a3uMtRQqkbKyLA4NrqBHz3k1B9C0txa59w3A1Q+NGjB8bRGW
SNj4Z5Nb8zefhqKocMi44fKlv8lbBmRoFd5RmZjdsyp4r5e0LkJISBwQixiUQ3gA
yAe+tgIYRzd4yLorCMl+sfpDDMJ9pioco5Shxb8iIfOpnuamqxXfZWuoz6OMuq+Q
/6SLCy61eNHSL3w+yD5ehSPXU24v3PoX5umVQ9k2pXc2pVzaKm+6b5hv2f7znDWs
hJTt5VKmN+oeupkRH9roIB/K6g5G4a2L0ZfVdyYSouyvT3lw8NVTT4DKbHfQjFlN
GAJ63ZpNlQqutkZ3BFke3SqyxcuZ0I+9l0MZbrGzWUDCWG6FMJA2T+QtTw1Dvu5R
11tHCWav17Ih+rp73iPiPMrbKP8qeThi8cbhYJk6hzMbafUimiy88lBH5KXBlhDc
TJ9EkDbnhEDWiniwHLgYPMXYzRT6tIN3JztLol4W3K+cLgC0Y84aTyPxh3VWpYbw
vVYCHCvtd4mlrR4GHLuMQRxm8C5wzp/fRsdGv1mMfxp+S1sp83884CSMSogp/I/f
Hg2aX6KM9l41HbCfxZ4bzeFSzweGAMsScPH+AjtX73T5emtfoZv6zfjnFQQ2U+e/
8+XloU1OmqdLRDCUqzIACr6cM5+N4Pt/+toqwBarsS5fVCzi3mB4PSjTPSybTmgq
nezly/cfJ8Wh/AAy3adDWp+WBobvEnyXwIjF5G5xOmLad+bh87h1051NeKyFtr1h
QT+iRWkzKKMrZrOT1g7PKJ4pJ467383AjAqlj5cVbYHvHgVak+E3xeuXXBtbzNsW
EGa1kdBOUS3Ky59rNO59HxcScWUfDmqxGjqg8qKvDHvzmD6RspjzcIVkhxP4eiiZ
kSv8Qtf++TpHKti/cQ0SUfHWH/+dSsCV4eaNTDQ/ABqkw/sk1ZYA6HUcSLUrGuU5
piQcf/LyVgzqCFuxwKW5IISrXMnEvel5JOGT4JqF+PVMD8/LU/AH8VPci1LSsAfU
EJo9cI6VdSy4zjOyjB6/XHyfz1fzejWz8O7ScbcZCWxQG3TOSYlWkTspbzpDowq2
a/uAZAzWwtXp0h5BNl0PHFExl3/mFYIAE07h/9DgozceR+hecG9wN6OtiinH5aEH
978lGzCnTcvTNkmufsHLl6SvgWnmD8Zb+0IZjLtg1G+JWro6sro6YD0QWeD6mZ9z
8PGhrOMXyDrLByYbFuzSDazd7av8vtdWd9NLt2oFfLM7xKIGqeb61fatgMG5YjDG
3ZMIF0ij9tRPWrsJu/DctBzennNzbDaFD2HZb8f+njNETn0TRVtznwGw/XO/Io7D
z5Chh5XQgFritVoRyUabsT3owjCUY492U5rko7hW+wQb3f6jxLdZ5nRL0iq7dEAr
KDwGP318zchAhLrpe3a2NwBl+MLzMHYGVqW0uw0yBxOmA0kYq1j6e/aylRHsWfIL
ZwkakaOnzZIRF6fuhV/BPtrUdZMabRKgreuJvPr/hlIj7xEojL3WinTYrM2Sy0f5
NX0dkewlsDz1JCmkF0fjPTaAxPicBZlUPmg16tFAAGv1hVdma04JGeoqBShKp929
FaisuiCF/niYn+oOLxw+kCAbuOA/BxZVJvCt++PV8I43ToAbbcMl3ZLgGnY3Kpr7
LjHmhgpJlyItAhlHX/vsWSrWxBj1kO/13PqdRI9v61ciH2wpV2wTn5eR/dZPH2ve
WRu4LsAdJ9XaU1ROyWmbMgrS1GTJyi4RTnveQgTNNnGjdNn/T037nsPjsqm4RDUK
i2AYabwmSJ6NkV3O/OiCvDTIvw1UwgpD3HNLIx0qeaGukKufOib0DyGCoCkyGXh8
HYTNeMWhQ2UNsm+Pbu3CJZ3biLQbbSCRRa9RUJeoKcLzrH6SfZ6+o/NgKVUv0qrB
hOkE0+ggIdBLkzOpYp1/+NAOKZHyJfYCef8uvakz+FCtaHHkWyD5zfgQprBBHKbC
zl5XRYn1CMXqejbO7brsKSQeh0eUO9ROMw/RQAViW7h0HZBhVJ05NxHrw4dNeavU
sikSsYw2hhai9e9ZwQ8sie29jVvD1QzXTes0FdImGS9WS7RVJp65gML/a7+5onGg
yW6ZFkh2bKij46Mcp4hrxsse5mmt2RAeRs8JTvSS7Lr86hSeK1FcMQrR9FvkvVJt
i3j9+tk2xGMz0qrPA/Hb0AfvBuzvgLExQnc6flu14xwo5JBUx5ETYaHErjh/UCVH
AXNDVx0iJ1ExSnuJCmUSBI6CLdwsUvUXMvhQm4kpFiNmoctpAdWkpCdbe0fgpcCz
svp47sU9wvwHSZJaF0HyUc5uqkMVCNgoxysDYIWmAUcHRG2pOKZAcBO4h5+mV4BX
oLr0vxlTkFNfog47i7pqvGLjl4UtHitXqhSwTfivgrhDTRzsIkpAlcWT0Pel1wIl
nKbExZ0qHSrZOy/X8ZUuOwPHQJANLwajEObA4Mv1X7IYUtBjmwr6HTHbsn/ehkYc
DKPUbwpoyADWsXbBHdtrVxHdMIKDIW4EZ56rba7wPMfP/xyy1lLj5WtZgucreZ9i
Q384CrIDfvWBfaDzhFnEIJIBYIb8bt1orHUAzKd/zOmMb8oTuKb1uxVSlm0bHAls
ylW0BMP1bqgSza/VBJX4GgyNkZM5wEKM354DTKslkIza8LwEmWtTAQ5jgoCIRpjW
A8fVU7dd3Sdw+4VkGAsRACx7y6LfkAKVs2l17ZGo8f2RqokvM/mQuUJRHYQ8Gm1J
z3Fc3Uhm5r9xf1HulxYES9DZB/GgJryxwQ1KHxFOS5sEdSmeMB+0Be4Z+kKgl9Xa
2zGCW7n6XtVU6cZ0YgS82HxCPy3LWANjMWUsvgpovf1n9ohIpCt0Jb2uI+2BHMwa
OpQF/0S83FM03hqv9YBJhVAsRCmyy/Xi7ciRrfVtzuvP0bhPLHqMRAB2Y7HmyIzx
V+ZQ9pIqh1ZGxm3Q3dwzU3jCdaKriFn5NLuz/ysouV9mvqIKLCMnvI4XfsRn2iBW
BZgy2NjuxUHcVcJzg6IWsyp0o/s9WJa3g+NBgUUp9whU1+4+PrV4vad/MjnnOur1
MfOaTrnb7hTAyNybIlW/X9hU8I8SqHpGCBVHwNOUrB+uKp5pxDsQTdNEfkhV4t7B
eNGdajT8+HvQfzX6yTuvrCBl3QGoXv/gx8WdiX4gM8TflgWfLdenE5jBsU4yDf3K
/o2XHFvXdDM3RQhsSDyUnjU7qOdtTp1aH6Zxc757jCEhQIxYPhFW6VZZC/ZsQ/wm
VZ+o8AX16goZY1YuBuybZVSWGdJhHoBTd+nHDIP7IfHRCuSIU4FI9w3HMz1QjGVA
tTDXe6VQeIrC/Re9mdPU/01MwEt0KKieg210rpByR1gD1Np2v19GgmL3XM2ygod2
BMCSByXdXMFQ4IPCfgHci53ROTI0P/ahYTiaoEcZVYgxffdSJwUT13YSpnvDCKT4
3S7535hSQcgch+I6eG83eM6klk76vBOoJrLespYTtFwpmTQQloXfDhFgBkpW2ZuX
Xpn/Svlya16Pi4OCuijnATU1Jdazuws0C2UEfkMBDuWwnomZop0vauYpJZzP9DwN
hPphyywmNtXDiPDei/44ye98kotN/1wXBrPjigmtA0wR8Am7g3jMbhyZutgni5pY
BKhnDb1P48EAWhaQ9HhYMwkLbzbE84oCwoN3n7ljA59xDYwJ2zmWqfo8YdYavH/W
oPHuwZTjFDamPiLCLaiIFuU/e0yPaFTF/NWOD6fkPRYmR4682btZeIyca1nF4JSY
1PLf9OM3c9I17dfUlQnjBFXvG22IYLPp2hMJuRTohw57+rvoHCeYYAHhtZVksL6P
8Q23Koc2n2y436aFNrabAyB+HpOCuxA+gOWFi/r7NAstfnLocjQ9+PF9iMYEI2YJ
Ox8/fPCinCUvYMNYnvlihHoERRzrA067OgYbKgrnLEKA1iRrMyIXGO4SNbGkC/pY
x+Ncz+mndCLN6kuPztB7mJMYBMSJR9TDh6cObHhlKAZtduHDfBjkyc8udbefyazz
vwpGyeptjl8Kiwoyj6lFjvC2omJ+9tU8vx3GsJR5n3DDaoCNkTXgAScKEaBUbsH9
gYs3tbCzr2bTtdOYfeHqwuoEGeCVte5eLIiC1D/FVliwTZAWH0UmNudV304UizWS
TK+rWvjmwaSCqgp3EL7LAR34NlGmSNT2cRT82ssSdztpFfWCdE9KxLG0gFbk2vdO
B+QiUUC/ShAKN0jmI4BJHGeNdliADbtIF/Kn5vWpxERUrMQWoWnnp1JwGilY6Uab
itSEswPLn1+CUg8cEAM5B7ehc2Ns03v/uy6S4s7YYa+EHkOhA50APQsWNrbZfvSu
ynYnUUk1pSc3t/eq6hoVgTgUDy0wQzMw1eT4PvjJ7+6fAPkF9bqd91d2pryNg2YT
PTZL4uXjbKtDBITcO+3WErGrKfSo7DKY+ZfxuJB2ERXHNHW1wq6mKLw+mBfycvyv
vYv+Hk5JKMca0qP9Pmmpo1DrtnMbvmfXevXWR9gAWqQnm5pv5/7f/CG9M2puYWL3
ANRH0Dqf0TZsJ6zOLZx31tHz0xV3+/EHnzjIO0YZEMOpTT8Ehp7VCx0sBRCGQpDz
R1bVXrGK0dv31uBiQnsM3YL3vfdQIjGCcBhmq1qE6buNZxBzB8WeXNImSQN6WHlJ
0dwPOY9pUn9GL6VNIMd9yBfqZ/Rm+c4+JXJPc9/VqCEHCq1LBr0TL/E5umm66TEn
3UQ/s73gkhf5QgDuOzZO2J6c03Z0aJy93/zxkeeHrvoV8lMSowxYhB1vxYOQMr4B
acMMLI3W+EINpkDhFnE4bvZwhXIMS4eN+MZQu5ZuYjrk6/vdz2+bKfPBnDjb3Yjk
IGRPzAhdOGZJYl7QOY061kmETQ2GPKDtd8sVPOGTXeEZbyy4BiLxuRMWQSuEDv14
rcy1DY7Y9zZMRdwAGy5DzGXFRrSSIKAA7YgqKndI9wLMRhMO/kH1iv9vVXM6pKk+
UdXFyKy60uQbGvKq7x9npW+ZYBPWq7qahw2IeXgv9t21100FyGfd3/jnqNeTmmyV
ZILvSX7whAIA9q1i11hGTKoVUCoGQwZ+01hGywbF+uyuLqdHK/nK35LWnH+14hS8
TSVgevW3/nrF+t0O5cdJ07QMAwk+4XaTAyX9FxOlPo46MXgnEZDyL7Nv383Baic/
cBVoKTnLLs0AkWelfu9CaukvROrEuDPRhCCWbkOvcofOZTIqM5jVkuM2ddkLEhIf
wY/xvZcnYgeYU9slqKONFHgPkxp2qVEbSnl3eTjLyX/Bdms5i4HKQEu2W2/M+s5t
hHSPOQyx6Fl7ghIK9JRsiO5DVsEEJpmOu0W6FMOgNCGORI35Rle9L4ZuJJzWo4FT
MVd0vk3XXAuE8kc55LcQEuMXMDvwZJcl/nXYEWoi0sWMfDS2qD0xs3UvqLSB7wxH
sgtC3N7kJiiDQlvQwM6o6W2a9TpgJ3qndvmXPmMrRJVBP88qDX/Un4e+1cPUFErO
nFzeelVxmlS2tYXA1SuZAuJlMwJ2LuCpa7u5N+9AhFUrfapnLXHDzW0C3AGNIwin
dbyuW0WocKh9jOPPf7YQxESxMKWVru2hJDesmV0Tr4XvtgrAQFSPGYZFUrPWNZTO
hxbWgiH7CUVTx29WayvF8H7iCZHFADHqQh356lbprlxnLaaRf/bbIumCRHxbf4oI
ryupXUWpm90MlcjwxX5HoYzvVDLpOLgsXU57g2lDLGQ72+R6z6plwrTstwMZSHbl
2cFbztjeKLsFbGAR7EbBeBh7gox55pG5w/g268I54doBZNtJyienP1raCEoeeDYb
ez9SfdPbh7r1pITNQoOxQiuOGxK6Vwv/rqoVG/gDLzQns5ZSySnCNQiSY4WRW832
MmqHf4wn4MmwbtzVQ6jOvdr/MY0KDEyUbDd76FD63TBW3RDBV0wjwHiWlOVnUDhg
JgoNy/Zua2UOo0CTtzIVMYZAxff/Si/is2KEEut8PoeKxb87AwizaJP2Ev46OL2G
4H3PpNirlMOBeaOWrXilA2Td/f5g43w9GXTIMp3JglUinH1tK72O3Yqn4CDTNGdZ
VfgtbZ3BVzPQ3uJ0Dbc+mrHzHfwMuwEAoDxRUDy4Owns5JWRqxerWwTXzuCOiPCd
TcgnT6l4e/uT6qT1kHeSoVWdXPvd8qzt54t7FRZWPeVEltL4/RoNsfMurlcLwM5k
ShHRXtWwm07wQprwkh89MAW4oPz/YtwqEmKVhkvA8k3lfIgA4oVcqDNwiBfl+c4a
0RbKZ8gfacDhNSEw6rlUcy0M+KIbz/gqBiJeyuuESCXYjw5g7FuYrTQ579H8Ger/
dmffkgRlFpDLr4iMnj6xqNvF8fNgvlRqGnQEfCcgHWK+T0iAkt4xcku8ojMJV9n7
gS/aUhVhYoLQ7UzetfbihGFsm+WL9QKzkHZLLW/2yhLKkSAm0gRC0p/p/0sJN8qb
nM9YnJigfvYoXu8IuGtLpcUNGZFqyak2uDU5J/+nXiACFAdHiSVh7mU0ikaA+Qw4
/ZLYVm2SSEv4i2CbWulhrDveuxBdU6+ZWUE7T5A3iOl6+roypgumN2s88yIz2sZb
E7D4jX8G4nA3LUyTELO4gPqxBqicYZ3HTdiw3kcxMSUFw2ULvjOoqtiAeXjmu+M+
gykB/lbZmuZ2uaKjPnhY5Zm37rkLFeFk7pRw2TjENgq335K3ftVaDHvp5b4vdfHR
ZzncLwUzJ3JRFAht0zt0yAY1zb7dGM4shF9xTsssQMdFh3OyHrofKh9A6oEr4TA8
hVjh7A3xgRNwq5fPeOPUF7n9nMACTqUZaJp5G+/DvI1GCmuEyCUBFdhvy++/ZsPt
xDACNyV27l84hnq5tdMp+DgpOWwHqX96HsiZzP3VE26iH17MN3t/sNpP988kSEd6
FMLilH6DYQj8ufJH2Xz0897Q27cHf+D7+hwP+xZXXUs3PcCKs3+WvkyAWwy6Nezs
eDC+IgQrmLB+oteZeIiBekah8sBwVLfvaoPrRABZ++qvUsxk5cJsS56xpNS358aT
K16zWjbV54paZirCD5+2bqngptdvYRJX7AuSNEKsDCn5D2cHY2GjJmOngTvFylNj
DJ1oFm4I3Z8d0yNpd4fBrE1C3UlwlNmpBvJCzGnMc6mq/cQMisYXGYD6noU18wwK
eQDhVBvb+pLLLYKdZ+jhAwulGjaRS0UWa8G9p11mXPXd/xUMNrFYo45FJK+YhQZG
a/s4Gvj0i8HkyT47pNhmYITsH4BfX5pTR0T539u+pOQTC+sE+JwXWjc1M2tP2R++
xoMWTrS/uQhwSCcnkyAJw3benNfaSq0bW2sqZlhzHXNqRP9LUyb2Y02V1rqm530u
JPXHoaE0JBuwQW+TTOIRfHQWzOpdlXNYwGB4wxRA7GxNHGm3VkAZJWjeSdgvxSLG
R2MGIFmxGzR/MfC1vEflui1eMtu7bT4r+brHICRZ561UciSgxxOUYd8+7oeTk5IY
iMnvoRqHwwd6mcBgIpgYkMvZKD0R2tmAREPHjoQCzPoOL53svpkevOii0IBikpuQ
mz4Hcp780BitlBMr5MEnwlDyqJoI2VJCzSlb2iDQztIqe2iurc6tLU0Izp+NZzYK
raMptWyRVruXXy6SPQNQ1fxz90sIFprInfnuPOXACwh65H2TSJ8Xa1Bpeo1QJxY/
u6iMcXp78XftrT9chbWwZWIoFWkvdLPEO3lJKIevXbnmp6c+o49m8nTswJQilveG
bUzSxctB/zv2CdhocjxqI9DAlhbCfGoL9msZGoXXxrKICY7oxPrJ/ypySMmLezoX
551GTHJRzn2i/VKf4/1nUkdxpNNYz5HkgcOtX1PcEupXyL6+cC3F8XkInbsSgYLq
XlwDfPmpamfrTy4vcXo+bEQZhoD8/QhI1Gh/7/hCR1jUdQGuQ9RLGL8op2I6X6cU
R5SVitLtTu0rv4INM3wDn63UNaTsy5A0oxMgjeolXJ9A41k2an1nLsR09U9tuAnr
MHmiLzkXzWLcfbriCixjQ03b0ZSdIDUhe/+gTdn/Q8/6KzTq6vm4rvcIrLXlHLdh
OQ/7o3GZf5jDjnt8qJIsG8Bt45fuliT8IVB+GkiuOzdK7xdTiN/MqGEAeVFlPr1+
fbZ7VPmkkR25FepYrAelMiRTeVNyfdhiHEEXVIXEWdDMhTST9FFV33PBpwkq3H9x
3RpEdYoxoUDhjpAlBjZrrMsoPk9h+lgOHSDGN0UpE2dTaHhzcGXvGmQgBMmTVA/W
2OvMl6tmXB7BRi7fVHO9prk6OJPkvvXWXcJdiTEKkclItZ8oDEU5MA2qVGVp92Kv
EJEUfxkvIW50J6AZu7eo2Xo3+5lQ3lux64SiZIllz98aWD07van8WOD3IggZHmYc
sUA+6BQ420Cqd9lwMouBVPzXCftPKO6RWyrMJiTPgc65DQY+qivo5Lhml6jWFVt2
mvyqLnzbaPsrudoWy4jIXMHLt0KaSsJbA+5rq9d5OA2ELWEu+6Skws9EgvbYgtzh
9In1VDwLXoFjifH87VSZBKfRPqn1qfuamwKrOOPDTnOTOTXEsFhNBIlDlK+/MLWm
/OIQGPmFoXhnjTaHc4/HthYoMo6jBjaQsC8N4ke5uqwdJKReNYqBnA3IBabLZ0AL
P+Ae8ubzkWnvbu8yGbVPZ/B95dFYZCoIK5CH468SZ4ZB4PpkZrZjnZRkJe4MwUjF
uFQ6AgXV9PLUxdQuGhjlHQdj2gu0WgNQkAtqxT0mjVyaRqLNfh32haueShWJWm3K
FxKASqN93bROFcJUuuQyc/W7qknIhN36WUqSI8AcHcc10jyfrCXIKVFho9hCtf0n
V312E6f++lgmgG9XUrWSMfDx0yCeedcBjI2KVaF3FvuoGt+g0VdBjrnshu5x5Qc4
439z3IGdoX2lP6El5AnDUQ7aejIW6iO1K5np2DHcD24ABtIVd+srpYroD4mAi+Tx
SlljQtx7ceKV0SxVl6+teHiUu7j8U9LmVYVwa4sEGVSnri5RVbps3eM8sqFkSopr
KAm4HZqODF+5Ej2UWGUQVYmu56SibcVGf5Dfmx+C+FtczYGOuWiCAl0lkVa9QDIu
TajtikpUo0pMLaZtZkLB5ie64d2BeEWdUcPVY+d540JT0vCruCQ54TX0SejOz687
YgYn3qxVg83V/hZURIGJi4AkYLYoCA/lVBMNU0sVK91uMxunfK4K5Jfdd3dQ1G3i
b25HWPMX/Eb+sPs94TymX/jSOtuiqMYRoFWetCz7wOu3Fb37nOlgr8dBV7I6Vh8K
DbSEV3UbkOJrwPogywb5b+jQUytIHMRwJMhI/aSSCWTx5G1+6dD1ibGnjX1YdzI5
YX9sY5FXucwGx35GyLK8dHzprvMwKWmY9zIj79Yblo98l+6gTwltgwjCg5AHbB12
Ag6XpoQIdou90Zlv/vmRyRnYu/awON6Qfx1qsrB7/UwrRWW6KGVKRVHBe1FbbCih
7lCPnTsx/QfzOqgBwyiXKMbGrrfUBoZPBU+WQ0rN/JSg5ZLLfH5n0NwiKytkoGcL
3oaXAp/cFQsHriPCPpmadEi5H+jQJ35UtJAPzEmYCmiE/2wc53s8HqJuXdzdARV3
p1SCqCUe7MhdSExHnlheq4x9goU/vh1tPqVMBrKCrqKu92qqKmj9oHyPbm8KAm1u
lPmNkJLjXRv4BHLUaa3jrmHuoyQGyhGCFdwJghxUEYatnqtn59uCgDnXUv/GTsbG
BLYr26zp02Ncda427tvfvtL7qpGLwRyHJaxcPnQTOL+DQpNPXf+Pfqp37i+PPBTr
hCITcDOzlCltE/bDn1w7n65S+WDProyV2PRQuz1CrOkw2WRKTq53ooBZ+A48Y4W9
NVdJB5T2kqcr/HKYAXP0ORn9lrOL4m/MMkTlwn0ZPHKUJQe+TY4WrPng0/wI3v3m
CJDasUWXmFXJx0NsaXBOrMXMJifkOix/gA/bEozWKPmK+/lA+zeb+4e0Q5J66kY6
5358cDUAOltw/5Sl6s3+mUweGCEuwP7OoDJUK60jsDGjXh4lfIQ3qCb5TO+dN2QL
QJnT8z2+8Fvzz/Fs3ugZ+mfbIyPoEbS6wJg13G540vJ+rzIjFWUYBpeJvLAj6sjr
GMx3yLOwp1xktQun5V6vHYERYWBQJq6e9ALjQ2YzRzcmUpzfk+qv9j6ZeTSdHYOd
NPEu73Y63dyQhaYw/8yQSiT7Ck6++SHI19ZfE3ELF9l5AsCGS8ozSc26tZiyO1Hu
d+mQ36rJNaB9fQMFSLm8Ap0pgQCTsP3c2w4k0/bPxrbSNgSEJpfEaBndA5s+IxU2
vDZcga2ZUEpnD0y2Fcuq2s5KEba26j087PXW8j9wF5d9y/mijKwD/e9fqGRO9yeN
Qc8fhiQh4pbuccsgOnq5ZJ4AjwsZv6tD40qnHbTgtOUNCaJpLIEM0GJ640ltxYhw
hoOo8AgvKK/99SZbKgYH4QrGBnUuagj5+ZVvMHaTuVAx/GyvpE2RjZzcXyOqoCKM
Tmvk3vwmrCJ7OjkbnZA20tN3navDHlzw0YiYbn+66lsR6egRGzlbJMqx8wtr2D5s
tiMvtpoufKmi01Rk4/eOMWC37E5yW/6pag1Fq2zvbidx1ZLOrpUj9hqxgaHOFFXU
Me7QRUUeGK6KIanfYyxjxshL7RnxHDQZ7KbQjl8PMJfsL03f7eGCPEgYe1BvMbna
IFFy7xLblm8mWP6zzIEBc9B+3Ur46yMyejHVBTs2GEPOdFeuISk9QdFqHFAXHW6U
tiiIbNeqTj9LKa+0QfD7KURVyR1chR0VCpPYP31HPKXv+QqXMxRioxybJSYHzjxr
d8x+JjsEIpRaBfnVm74Afe3AmNXMHdSMCEmVcE8CzGESavkoxSrHblOIBRFXNVL7
4U8i2Uv6szJ3PRFf6DAS1Tq+lBpQ7pLT0kZM9REI3SHiYnPr2NXWIveT5xBbadkf
w7EfWm+nMmEtszNVXxkYM3u9XsEocYFNhHwav2Kf64YkMpbzvNSTa1OzfJn0D6Rc
rOarnIUwfOSvpIIJU6kV83pOqQAyhUP1zw4QUQ0h3ajaWVxUFUz0Yau4Mpy1Wwv+
t4Kd0qa+zf4Js+HzYnZiyT/kJ3v64UfcR7XsTopBzFtb7zdTGc97os+YMDUjj9+O
V+Sj2zn+TCaKPf2UszKQs8obzPJDZ1YQP3U6pl3SgEYteJmT+G1jOnKgSkeUk7HF
hszdkF21hP7nA69bGofgdgFr0xSq5rFUJZUtgsHkN2Q13jRvQxi4uLu2cru3bCXQ
OTvqCCRugXCLm/45IiTaJYG0KCRk9Dd8Qk4ZBPNUCEVZATCYxp3NJNQ/vdvz1YHw
YJquSNdS67g0jfSnNj7RBs+4DGMmOgo61cEfu6Z+RfwBJHNxtMx9malEYPlyh1me
5QzqXT0HWBgddGdMY+fUvMqMsSngmICBB9WMorOHk7dLdO2ny+8SCgpKJytvsNik
EujnWO9zW07Es7gDjU+BwI4eDYe3s/O9gGSET4eUJZKO7KSf16bMNXazixDfcAT8
JrejgVV8V0/fjP0ACpsKwqDAB2BGANUa5zquECIkfPtITUg0WaD6IlOSRYIYRAHf
arH0gOdVvjicX4LE2/fTcuoKwQfctuGEehVw0Qbr+ef8I5bb85nQ44bxDJXy4tA6
5WPUUDyYJiSMOTFPAQFfTnVbWuD0tdx5lUZSw2F0ZX5AuHdZzGkLizjn68Wwc9M4
SW7bXq1x7Jqpjxudy0SFQmgJmKLC4OU9YiGfDSFjDMzQjIKQ1R3yTr58F4Iweuz9
9vaksC0pFGUxP+AIpaO3fzKlSlHvg3vGRot9xwK536Ir8ExoWQb/rtPWAeqPJSAy
oRFh5wnLzQKAPmH3Jow+ef52cKscqeUJgHJyrdMQjm3nJR5WExwR97WTcc6neKhH
UTxyL3XyM71/MmTnSl9cE5yPkL+Qm5MwslAR7nI2rxBy81O0BlCBsV4p8ubvzlU+
kiad5TkrRS9HXsc+hJjSRMr3GEmj4M7izSizT3QJ2fzpUlmR1aF7JkiN8h0bb0K6
hRJC3pTjsb/uVZXqUCE9nKuvdIZrpIZgKxqxcINEC3Ft+gbm77MZ+WVF7NwLTTIg
elYCWQVBrcvrL2GnnFLFDwbNjChmlqcnNHw9heTGQrsXLyQDD6VhqIwY5wupXXp2
MdbynV9uhcGQdNlM/UwT2yn+yUXqgCszKjSxoLB7MVnAQcPs7X3UhVXDV2NsNP2U
P+ubSLqouNN9hyi5x1BLvE6Yfvto8dL9S5W+VjdYzUijNOEbv/hOyAfGhToQI3uW
YrFitA3tIT1vbZ9qv2tD4SAMGcXIrFDosN6MDBUwtvkn7dT30UicuE8Yn0N3zIY4
4575IM9TgfSk2AHjudrY3r1jCoqvsQYok7HrU5CjyA0HbEQvHB/Vx+yn41oXVyhm
PBPK5VJpWDcbAujsU2Ke75yig/Jeld4+TNyWCM+vlQBxf37Gw8XK1sO8ubIMfDZT
ifZWAj3lvPYSSxmJtJT4Rubj142zeLMFgWRnPW6kDAhDe3kJpRsUcxLlrGzaI2gt
Laupm8+NYPwPYxWcs69WJptIPWEx5nFKpm3j6yYfnAVj9NPgfzGp9P+NVRquObKP
ijxlMLGQXctFiPsxbK4QgeEvSde3ZgM7OXB5kWuXsRvqfeJxKGnRrrxLwcomnnRD
vmsPLytaxTt2uhDg/zqGM6k62sH+l6F12+mfxNjiPl0maeMPIBD0eAB5/zC55LN0
QOQhIhgp2LsO4dQK4q3GTAEVNBzP91OQvKzA7LnK0aLpuSXcu6WKCCd/QYC+8avf
wwuFNCMbyJOODdhcMb5QgFWmNB5kDC0tHdPnEeBkoqu7UNdr8Z0Gchu/PM9IhKcB
0goux4J2sj/qKH3ok3vNZJks4VGeEaJE/41B7algVhRTGLeMJentcNTDt++FJD0/
EcbyLPEfsXSzJZZZWU1aVlbk84WJd9JUqmEGbGEn0NJdAevB/nBkGsGIY0pqM9a2
VlfCmoLenpE+vaPioaqgnwftwIRqfRWTmD6avwfsrP3kVHbxFwoceh9GS91mqEcn
G3REkdXeqzVPfb3gIIVWZkV7Z/0jjn5wZO91MtF6veMajY0gxOM2M8RfChr6oTu8
Tn5umWapNP/ZSnQJaWrwg8Th5I3W0RFt7SSy5u/XremtvfndBKdVrrN6P/ycRpN1
WZhpI4GggY7kA8VHZSYvmaPQE09NRsLt8whlZMKL+60btAfvYHMNMfnDeq0XVkXd
hyCkYDhbOM2BAIPA4ist4ilVytQ49YkAFzMlho+GIXcf7xPd5ZqSjNKkD2gQEO7d
5Nno6AdxQ6rFOXkfMRU3x3tmzgSoc+Fnu9+j48fiunrIG9zyiP8JXaCeONEHf3Om
1udWRsns2fkKeQYpQUbnWlAwXU/DG3toTDZ+cuNgFApjIM79IYmzFEO46JSqNcHt
IrymMaVTYhZzfyreyYnzBrMwq3wSMBvFYbwCpa6BED1iLw/pdgtUOONjz7IY7mb+
mVB3Cea8d/dSF5m96bvishoFuu5jrm8os1NTjacpmpxJuhK6dpyztWpLHj0/JYRU
uQvQGi6Qa7g657AnOcSkSEiUByrRiFmt6I36PtL8+jZ5PjpgKCzNU2i25Uc8Xrw/
Ek5ryMsc7RywP1NcogO/ZW8EyLFC2Rl1elcX8eSkzIk8rrpAvJHMkyhU1tI9BSRb
9zMl3i1xWnexQiMc8ojDBLT0NgQ8QR9wmUZzJ7yqTwk8gTqQxcPZ0rH9kZ7usXME
UFPO20Lsnb0txaqRtcZWyCXBtneMMsZNS3p/mau+GOggWow8iYirzS3XfXxfKFlz
y/MjJrywfB44Dk/Cbbu+3Ay23X2k96e2hI9QepML3N2+NYCN/cPG1TjwRtyRs08i
8CBFgpVMXPdWuL5QTZRoiW1MCliM083bEoXqBejlfVlTjR0FiZpOns5klBBfWGEd
7bSR2g77go2vrO2j2f0NL3/Wh/Y8t9qLnY8ABrX3xZ086dd3Pa1/JYfG4eHdxI1j
oyOemD4knB5srV9zBgg+N6Lf5ot9eG3xWARYhQX4HpYmtKdt5Jq3q8DEpkfcFxRb
l/jcjYuN1UEPyRKA1Mk5+DpNnw3ZZLCgjtoQfX7+kfu67xPTGdj4vklQ60biwnBs
aZvj98FkYkGJXgpTLkvJW2beyy/90nWMkHOozXupp5+cdpGqWVcBFI1i7XbWjfp8
vS/eDL7EE2gNUzxXKIVxRPgdvcV1GNlxjR8V8ww1gv2xRBttqIe8LnZEwDLP3SCe
5dYbTjiO7hVbjoMpaZm10wNa6qrXGEttDmM0n8Cnxj8g7HeKubB1x0mLao3VEQ+Y
V3SeZKLlUJbPXRjEHQmcBsm2YHxQ0QhQ02Qhw4f7x7rHWGXlLumYjIuBHwOqaLzM
qHBEfb2FtzjLuLG/GzqkpTLBo56WCHG5tCDLZJK+Wq4s0twpNAfCROwlXD0k4CGO
5WpPZd8Mdly18LWuNMyw/FaFc6Ml0E+D4FSK+XILT+ne+F/lLeEv/B3/1IAKY9p8
vMlAR+nRb2GvTujuAAkr/N7OPp9llYQn6StUNdZ/fUqBX4a9951us7Cjc+mZYiH8
jCDnFKr5HRKFE1hW/SX6JoxYFkefpHmwFoc2m3iKBJGR4WUuuP2s6u79QXNsCk2P
QoVhYbOZ0I6tY/+Cy9SRYCcvjJkLelHydodgp/C0f4qUvc+nZfT6kx992tbzgCvJ
ui+2Mf4ndFu5HiqHjgK8M/FaO1MlNyozJaC3FCz5EjopNj47T6WynW1X1N/ScDn+
R/552vCiqxxk7ArtQokHvnSnFsOUPyKcUpDbXXqDqa3pZW4ihpIUTAm3zv3D4O/C
DggZBKd8HkyFsxbV+479ebaM6XQhtpQZ6uqoYEIausR0c7MJhIcEss0B29SUkaNC
OJIupAUuXEn8dAXrvfG4fCjzxMlUfhbGLq29yc3r9imA07d7/bMkzPI9Kg00ai/+
326UdFb9dmszf5VwoJLd5Jc1lzHIAvQ+g1zIYmdJKZcA5LpusfuRhDdKu8GBYl8/
PMmGrxdXLYD6jhxF9DJCmuC5T/GGXmVMuCZxDTALlMs6HrNR4n6bKGUxq27l+JcW
4eP9lZ+WkisAxcXx4H7jzGspwACckrdtPqJ9qFI2fc5oaoEVxTHwSN8e0FeCcBXS
Od2mb3itmqQKNZxoUxIfOG3StMDjxIiETZNgOOV8qt3jZyo5iWQCvkGx8UwofzmX
JdxSz6WgAqmy4mRNgQLGuTaCETgBnAOBgv7JSUTYiRMfLIvhsfACFIi8Hnkl5NcO
2gu6Km3NaD/auFoGwC7HuXG0aqEqfFu57RFuNj+gJIBYoZdFqk5EHLm5aHC3FJsc
BMTxIoLQKRUbV00odqLtJE0n42cf4aJ4Ngayf6WDK2CQa+KrtcXHOvYFynNaDolj
842WE6tCszqswi7UtGDBG2JscimCZz+Y0sA79LFU+9AODotGMV6TkokQ+Pod2+LV
R7cfbbO8DT4UatIdJhGL0XbUpwM4e6wi/2Hr1kMjaphjq+RrF1hWDdx7pWwWBtLF
ZThqIFSCMjE6BHXw+304PnA7aqH1ZCKKdz1Y0RSipfY7TLxYp/S358j9EwnCSxaW
rbXo1m/2bsmJ77jUJoXGvVl/8Mll1bzoy3dJiB+AMAf9KACTYbik1VHrMBt8+pnF
otGN7qiPA+MIFKLcXmC8RbzyUERuYoyqV/H+iOlBHtWITYqp5Ix/ZVbZ2E6Bprhn
wHxDqRnW8w2XnBYWxF8DJe20bO2l0j3dOtl09Ng6KKthEtXky0bqIolrEAVWdnqF
V8OAYR4i/mRz7tLr2n2V11Zt08yst+k54Kw4ICQgXP8KR6C85k9UhlVib2Tj7Ce+
xoSy2JAuRI3vrBtQourgfYFS0PjL+AUysQqzcobXG71/nk1UMbB31cH7Gr6v5FZx
qUBDQgE5AfQcSyZRlTDRkPRq2W5UG1wKlriwnGmmm2SygUtGNyHnh6FTUqN7zCJB
yXkomBbCtVBfCAX48Mh4veKFZNoV4qCTRDo2JfO4mu+FzQZvkbaRcJokiIycJC/q
xTZPwv6pe2RB0EOEprKreGuK9EHvHaWKfgZTnJdF7SzGAHZ5+WsgYb0C4/NwuLMQ
oucNMKyqoUj5134H4dLET+LiDtEkeukG+OaSbJbOl9l7xHhzkeDezyAA5tBN6vsf
8vSMJMlOFNhW4tsUEjBobHBEg6x9AvWFIMyR7NRMQ5nNAYTTVSYwYEW/qORB3LDO
GOXbKS5MkwLm0ZlOOgU6y+jENHjPg4Gr/Ed+UlIdR3lfG0MzviNxfBhFiV5GoK9y
vSkXP71Ovu8Khg+74K1i4L1Hc8LmME4P8bS5JkSoXHhxSVdjLn/KDJFZ9LMTe6Aw
eLI1lvZajlRuDNug6a+3LbJfVshF+R4SlQ64V2UQGAVUA/h5tQ765kUORIexnBVk
aq34fUvmbNIYEJsOtTzl36/ezKyQ+DDyQgGwS8eAN7oJQowrhXqD75N52D69cvwF
X7K5/IT6yFtfo0E+xiA173JSymw2fPRLAP/hErfG4V4Fkm8nF1c5ZCp8Cvtj0Rt6
Yky8m7GJO0rr6td6wqXdIsjhpqq25MfjisEmUCITXrrb6Jy35SUFbLejzwMCWgCr
12nEGD5BKyORoklwHQuhpPgHuCtdv9bfhGN2SyX6PmqGmmHNGoms8wrfusN/aa2C
ekVc9Z7tjD6FodCgYxQJD82Oi2Xyg+r4bnfJ9HKbgXkdkWA5IKMR3rZU/Zqfz6Am
vY5NcTkYXVddjcQStzDicFfjHn5/XOIck0vqp3sVSUOp0IMNGvafd2S0NJ9GQAH/
6A66X7myMORsAfpFyaz3x34lIjllhERXzNfdL8xcAT52MXomMqqV7vs4+oQB2Big
AMXlEe2yf5WJugb+KvMF7cd8z8VcMVSgsBWTEG6Kpvzfk9EQ/VKt8u0LzBiDu3Wq
ZhXEGswO8ZZLbcLvuxUtYV4D/Np9YwVggOnmgx07MknyaEPIfRzUizXmeXXSdMdK
i/nzd428tY4NodYekniF4D25OEPeMjbrDcr08vOs4KwnssTwCJ4Bu9ekXyPTZg92
sNwPWAf7TRYXDaagljKPnkuO4DaEONjaSFy0R9GZ4wN9OLCBGXH4l7vvCsb0vUc8
TFe4MLj74vL1M96Uj4Y6/wFTtcIPc6PESgLeEm2Js0r0p2JPduAp33pi3YcFlOQn
s1AskTyvFgiAqfcqga7+YjqMZmpYM1CclWeiyoxyDj5au7IlpmMicxuMrvQIW/c5
uK7nkn+PwZL7L4Z+2avEHtouUwx2222iJ0uDj183/4esDFumHKgFXJINqsS92pJ3
w/Ozjo9X1C+ehfxtoIZZAiHs4wqfXriI38b7z5XMSlxi86yrKcUMADC1IgR3DrR0
Bey/9jFTP7V6ujk3PVPyaDVvl5ePZlf1GxV4Y6hvo9Pz/1B7Z7y1ESJEBmYUdb1l
Rfx/xAnWpT4Ny5RkCt5nh2eqW2+7oeIPUbRZVuILDxWX7zap/bGNS0qjsO9b49MZ
X1MG36F4QR8kFrj6NSHPGvrTWTo2Z4btGfualQTcPO6gGT4T4lusb6FTmQBMqLtX
qElrRx1xYnsLoKxob+rGbt5UGUj6mKYtYQeCbf5GXMs1bxox7E/qiVfdkAreRGcf
3GbSx3TszGR8yrL8Yh50ItX0qG+CsS/mMrKvKz63Lqasi5FVbOVi5bRZ8p+ipwSc
vGwtjzrgT+q3El8tbjUE+dEpHwVbZg07EgVbvsTiQrmwFrNWN3w4SdN6zIuCUq81
vL212Fx12cvc7wjAG7CiX2hR6K7ryCgtqqdCTCCC7pHWTnMkcC6GbydAfSKTVWeS
pxMjCOxCgBSk1dgoTLK0i6srLJqxAP9SPpMw9SEgDzFTp0+gSY666lCpK7PlzIgj
1VOqtcQbFScQX+tli4f7C3iFWenTsGBIhcTrN/BbaM3O18loN2GK6tu8sUol63Ht
H5kE8C/Hzdflrpt4hkwGQZ5o0LA1yg5SKOAMcFgV7wrhXdx/1kVjCASvf2yEy+cG
nmHb8lYjYN3m4uMzwv8aQAYGYhlqqpZTuWQSBGY72z0kShuhQJv/XfhIZMtKgjPo
oBmGi7s5JPU64HdEJYDN+BrNAK4+bKenTvohpCqL67aU/vM55CqQyPtMizDoPmsH
6FKfyDx1wqbO7XcpYV6rtGsihQvcoyUmBRuwBdjsgEKe4gov1Pi+aOwQS1CSYhs2
+DqkKX3ittU0Ta5Ex2FIfcdfBk4BgeAuNrKxz6Q3XZAb3saOFZonE/II5Tjco53D
dVerfabzmJrZDlV23GMvgRkEyIDbcushz8orK+m7Q0SCAfu0I2xoO37czFuhmOHD
cJD67klJnmFtFZffsmwFymQsrT+8+VVc2xUkHTnxc3kIKzXkKur8TeHnrPyP50E3
m3Ognc7wCBntNYhc9+YUVtD9p4TUo+wHnbAMQjKm8fTBupXr+VeFD0exy29MJU+v
YGvKxdRaAjFtBXBF6bmcEHcYFd8ApETkzLEeuoDslhlRngcEU28D4CRi9pygCfFx
5srb4ZZ4jsfzhn1wbnC/kO6G9KIE3y08wZKToQC0gSUpcsDTKc7qK2FJPMtMCU+f
aNADDPbJf24RWzkMwS6VJRQKQiTI9PyYT5lIIHQcwtECzyCOc4cig/FCY2AXvn+5
B3vdx4Le7jJSz2+DDFko2FxrTdOhrrbWfLJUgetSzgztQwribbXJmQPY0x+hpknE
pA/ReNZFaCYskwvLCJTmUiSrNyADe9UO7RZDUjIORPlGgxONJuA/Ep6OzG0ihjmY
aauA0k10OX5t1UbeQt+CKeZPKPv3yk+iRuCR3D2j2d4i2VdEOOm29dvTEHPnhEdJ
2ANZnATipp2fqQWLj398GcnwWWkPsKOHRc8V2wCHWor9JGpYD9UOFZEpTEtf9NEb
evpM5s52gsrWbswcxd9w/vbnpKIcqYMvIgaLM9xYoEm/YdD1IjBOK06lchvDzh7X
9uet+D/V6maQHB1mQ/zT0O6NmykXxzcU7mI+mapBk40/pTtCAt+qOw1m/N7oGfKH
lPnK4fGdsW8CsW01zx4+XcFSTnJpi3ru7i+llAb/VEflDZeJ5lMJz77RZGoheuP1
IMd6sD7zmv/OoSYQPSXZ1QPrijXHlcgtNEPJfCcxGlEvG3WSMTXvyOgcSfIYJqIO
DcvfxAvyKuTF6VWsTT9nyzuJ+DY94p+Tf6Yw8a8v7oqnOV1nhC01Oh2uDZ2FZH/J
S2Aza0e8js7DDKOON10akdktfnZlGKCAYDNjhe/sCktriSnED10jaBAzExW5m8BN
MUE0dLyHZK37racQkUltAcvbdtRDXcjKTOOrh5OLz7U0XRFlUPak7T5iwUUhkmAk
5JxLYOqgY4zdj+ASV3CAHirh+jOcRJ67ggAdg6pCEjtpZ8i6Xr/AUvUdgPEFCZlt
9lv2DdjPkGYbEb+ZDobygpKpXWMOJe5CTawawkWSqNguIbOCDH0yt3bMSeEP4xeB
UOryu4n1W+XZN+aesYpGZkrk5kmm0lc9W/kop2lRU9HI+edPaNIdcoHwRvYsYerM
ZJ7Nr833zWdAbxE+lG+Dc0kUH3bKl+yUxbW1ms0yRh41fznkqcJb1du3YwMmvoIA
/St957ZezKOuDlg4FtAoTy15eSFxacPRVKZFC/+dAF/StPGS3CJuSWU0kFxsRfRI
JQ8JQ/4bPSBoS7FrB/YJxHZGPe7DEllZhZFGWqU8upuKXQwhs5XrZ2a6nslTuYrl
joYa9KI79hi9r3c0eOYaKgQd5utrwwUK8V8NEDzxUIGPY7zaVxEQZAyOyJgD+8QE
SuTM29U9v9B8BrhIpTHqjv8Lvh48O+QVNBuIk5SVjP8yakd4m7UcaLbkkLKxsuPj
vKzVwb01EOuzEYSyk5Fzk8uY/CHbo7jpZiwrGXgbIZZm2PBurDD9ePZrSamhML2k
xHS7f40ABcRn0r6C1ph4avMBJPyeaCtks6Vz/GW4RQbaUs0wj1Efjfds0I9F9tLa
npTS4biBgGE3JY7McILCzHPKqf4VQLs8sE8kB/Ep5B0MGNKRA+1gFKRDrxQvioQ1
HnCOmkxGH1pcoVLwQZU1RRzJfKASb4oaxLjYThZzRnhQkyl1p4OOeBmQxBncmUWR
Fq6YFCo27brRQORBGr8HbhLEVdekiLd8j/0/Cp4UNbJtyIeu06Rops3r17PcgzBH
zGl7oP9kcbcsuaQOZebzQOxAKzvP/ccauPb9ELE+U9yOwHUQtYNKC+s8iPeIGVDu
jjcgk7fROgJBT/SHjouaK0TvOGXHCPKHqY3k6ljXKb5NlV5z/quZia/wKTYgz/cL
O7B6JLhbwZbIUfjO68bVjeOFrcmt2PTBfQeEKiIJlvgAyiAxnC5l9mHG9t8O8xDW
zMub9dmmURpwtmHFy2ssVvkQu+x1N75bbPtMYK/DILW1iWoykDO9OFzDqBsZEz+D
D8TNUc5nGCD5Q/zuKRqaZHU2gbvECZwo6/zP3VWiM9et3tt1IWK5m0CthqxWzIaA
6IymmrP7wKnIgi8azr9o08IlJshMqI27sl+LF1KIIpJg/lEjp6MT1JVFk9PvYr2D
aZct422DQ0CV83SYUxQK3owWqe+0XT3LrKyo5Ec1EF7/naKr6wKulz9eX2+SfzfC
UNZIegj6aHvo9PkAZAsVlhozz2DiTcNPiH0GtBDCNs6OZj1H5WFRAfkCvPnaJykc
W3pn+Hr/d9sIEHXpoon2dz6YD5SJTA3NNT0BpjM/DeXPH1yQAqCqLMKYKtNUQ5HK
UBlDqKBGW4/Pp0j/i1uJSiDWM1dmxgcexZOhz2aGcA75IByy28xEblqbkDg99o7X
hJD0rsRB3yiwO5Li0Oy8UgQtFZYZhxEVEWrQIDPnd52JpN0Zir/SPEgnipm9Gtil
sW113ruYHYPfWd669uaWTFQp+CI0/yB/5bzxPw8Lr2wW/Revsiea4Qr0BeqAfdvP
bqOWhRc4CkBo2S5i2kx0l7KURKBlDlmwO/k5s1U2pAI7qji9zKfwe1fj7LQLyW9q
dBpb+0zOuF7tmUlPAGRyMWskrECQbsM5/2XeUPDMpq++vVqa04UZEzM6u5X0qp6G
n/Xu4UXW0TKL2YwxE/q8D+ZUrHcuFwzMNAhXj6VXsmHp7xBzmp1A5FA/5y3wWSRD
VKbbNZu+3OxSQwaQqk9zEyEZ8aGzhEGjrLU7KcTIZojkyQcjb2TCLlJPJk6k/mP0
FtJVKz6TMpksJqwtgp6jkL76aPtBXKnl/hgq2iIz3sMkHbP8MJEIDjMqKCOCqEeD
Jp0VgNmhi738KWHXrjTnTU517QatLeY7D2bLAyGNYPtZFA1LRvKBS3pVriyR2Z+S
jSAs+f8nmW3rL37/LZigoC0hfm8yUgydKk45bpe8z9yfV+8Dva0q8ymep6cls4zP
eyZR8XK5Pq+MCU9tOvnLWVjOAFB7/BfodYp/cqCfZdjYzPr/ONKVberli0m3xNd2
1mwymTlQZID672IXkguExJnv9JiqzacnJfkpeWjSVQAv1X5S0rdgMUC6Dnjblckl
xswvJkzhirQji9ojMdrVw69nMC6LAznW0z8bV47OTnbubSqgO/5EGJqZH/gxSXL/
GtY8GmfIBMXj4iun/TxEjLO7gDE+jWKOE/6qA+o8U1UoMBuLm3KVtemVnve7jEck
S4NLgo0K22l2vipqRC778h9+3M8nBBC9TQicsu10g55nPTWwpR6v97paOX8YBCAA
Yr13BWE2Vr/0czp+BtmAU8RmA10QLXm/ZiY8W6CJSlR+xKfLR3WU4E7PawlLZtyj
nwldtOmh8V1hhujcSZ33y+OdKUt8QDt9kRcEEuPovA0aV9SKpcQc70QlbXk0ws2d
LUuxr3j+60MeaERK7Y1UwN4lDhg4z58GugrgTopP2bu5HRgXxgIPHtwNgnA5LRPo
IXB673Xi3NMQDtqalsu283mQb+9I4ZTtxyMGDnfBsMh12UOaM+168ShRg0zs1yNm
p9I6wcpO/Z+n22VVQ6Gn5mtknYFrZZv5zYtpmV5EGJwwAw3JL7RUJXYzgXmcgpT3
6ljo10MsrL5pZCLqmU6NTqRAcQBxib6/ce46JGsl8SDdWG9TME6TBoqW3MtCkrIN
PJyvPPE01q4qrIwlR/ugbrG++KvrMvsQ22S4ZhEesbGNlWJfx4H1l2l7A0NgFAss
5szYJ8O3e1M4Zu94TfYOabf+ZhDvKtoz59WEuNgcWkz5ik/ksdkW+u1Ji56J9x/7
eVQ1duGxVHScmCI8yZ04PWrPtPA5uFcMGrCDZ/pg+3j9JgOsSm1mJ+iOQtZZUFih
GUNfswJcXELdO/o2rPCCwNROa89BTuhFDIYsbyR+jA/0DfKjv6VgrwN5HdcmWHvt
ndZgh1laMlsp+PPEkW+f3ezhyk7c6eSagrOwQGgKEINr8bkFwl9JkOIa0HgyZmsB
vOV4QZ4QieFeEXe5xU/LhEC9Y7y9ZIUHIZnnAwWxXdQL835jGRWy02b1bIKBDZdj
vyvLXSRe3ZlYUt24dK/w38QFypf+njoiuYgk17gYTPsMQXC3ejBis7xnimoJxVql
nG9gJgRZY67/jfFCKdFgd3F5Q8SGqNuOo4ArI6iJFPJxqHrQ3606/5WMcojeh1zv
4b1bLdHQ/mTVyOA1EkhE2xYSmFbT0bh2Ucz1yTaq72Qh9U5szoXBshV1Nu1lBZNS
K8wtH7slQzHTnSjt1DJzF/zo1ZW+UJmjC+b818+A4ElN32PeLiXSKZ3l9ZMvT9IU
eDyNy9UQjp3k4qvqv4wqMiqhIoMkNSPwe61otcWgP01dvUAGcnNP5FBwiENV4tyf
MQJP0G3U3xVB1u2tPSQhc5renF8C32aGyNyokCMHTxRNAER0YxGJhPj33CgCncbM
RZED2MUWLJCO151sRDkLoWRAE9RyTfwEjIMioaNMkWiRXVsYD+kOhbBoc941zhgJ
afhEQROjrVxf+8j9+zpmXuL3jpcZ4ip6WSSPpxUWT821RG23EBpeoZ4v3eaMIwil
zTQFkFHS93Fw+6onIk9qB7XI8GQQX2QBta34+TeRMfyaysxh0tUe8k1nuKSAY257
QN2Q/L3hcQNmLfMqRBny69WH1l2CkPaKPKZjMJZbw+zMOU6y0RyBX2qElgGCuEZ6
aQZkMRctDE5Rze07buWxZFYY4SD74R1bZORRci5kUBbV9DMNnHl15SBkkJT7xr/J
xRjWRfFooM+Av6iA1IKCAPq2/OzrXJTHGRC8DNK0uaYcFs5Vh/31wnAXKhki4myy
4MDrFg5jVlwZz1KtPxZTgQTtb7ZJc+WAnXpV+IYhhv+drz990rCoJbWNvbZlfj34
6g91NWLEvSr318x5r6rwrQq8p48ol7le9X7gtHAL0IcupgaMMtuTRiEd8rGf88v2
lFpwakEBUH5kqUf99WM/fnEveWWYvnHTfWggS9aF3YypkVXIUz1fyaiJI4Z4HBM/
kZjYN9XZr6hwI/ql05dmgAQPwq6H7wJKbVIaj1cTyVQ5l48fyMVAON3M0WfnhpNG
fbngDxF9skbq42dDCBqw1CEsNfK7PR9ZgFFu69JVDhptI9Xmr70DRn2uHtU9sWsz
lB3cMZlHeWNAFxmloUvjFPzRKQrf9y7sx7b+GcfYBrgcs6C3xHmc4B126Re5QzOY
+JMa79Xs4fKsSoqoKBdNxzZ1eGuJR/+znttaK1O3jdWrHoW6sc8rXn8sl0p/2Mw8
g+e/4sTDsyHsiTHG7fGK9+j+IAfdF6Sex6uehVSkocJLORWSS11LQJNtoAj5g2EC
VBxDpJoVy48u84QKguyqELFfyIdlFx/P+H4m2UFqKVByRCdykr7CcPQujSTCXE65
bm3NzhUyL1o+QfHXo1w7f7MOS9bpEIAYH1IHS+6YjcmnlnBT3zaF+DBLxG1eB70+
vnKnQagXDWnw0o7bFNEhd5nS8TpqEAjJgFQnipjmvfFEruv0PGSO2MeambIvldHA
vd5rrSomvwlTapFx8oBrWpw4Jqa+3wGn5XRQ9HAh5+Fe0g6A8VAm5qILOQ3sVVQ7
YIzk/hVGS8J0bNFtwAUI9/hoxfxmxB2cSIMWAKCIzuzqqDfEK79Fe4hoKMkg8pUF
Ck2johHAcyiOh4Q2/uijB6w6u50eFkqJDHkuB0ZHtaZCxUs1Y2wrsN0RTnuBjMci
g2/jY14S5Vdb8uy49vaYm2ldqsZ/okgUq0uoDoX0yrJvMYq1MApjcBhifiAr+Chm
8ZVg+3eTAxhwyGtWCg1C3LQAFXALUG8qymuAEu38X8zrzvOdi4USxsgD0u7FCe6P
Y695gqQfIaCEkKDDZjGdsLhqpfebUualv6AWxZpy7r6xK7umv0qjQzIIJ1GPko3S
1UBVE97q99pGKV/GfCzbv53jYb+EXu1R44BP2/ob5oePS3Ulwt0ZFRJiwYETTMZp
BnbCqTBqWM8uhekNq/Zr5hVBCo4ubYZz2nbRzfSpdB219TOFWfxVFKWsVyRvhDBN
TcjpyKky6nSU3yx+oRsErUZVJWAu5qtB1TAlwTkzWOL/0kROrZ+KodKUwio31tkR
2lpLDSRFQzmBQajcqBOitPmsZxRf+wmHPNTImDS6+Ha/r0xLMi5DRl6UAuqj+YlR
Bou2ZzKKYSYtL1xE2MMZ5oEb3lvE2S0EfN9H/bpaGjPvY8LLSBu4j3GOl1dtITbV
AC2ovlZBN/ru5ozEV1QP8qTuZQRvyskUSolrtTEUc3rRCH0cftk/pSC8gHzbQP/a
149AUslvEOFXgoNe5OrJe2Hz/CrMfeXUg3a6WvJaOMDT6yn2pB6g+EJTfIsUpsSd
O3LILeSfYIknQYKHyqbEgmOTqVx1Nb5zASJrGfERVKohCZSm3rqUimxPpK0izHFK
i3wLB35SxKfSf7wWaEwVbI1nwBV65k6ZFfVGpJt9XVX/Tix4OYTUs3AgAZ5mGltH
icgq6Z6zOiNzjEpV0J5WMC/umycyMTAQX49JhtXdHtGKl9EfGjIPRr3rzI8CIfrN
jx1h7OX/gbxH7jLN+lLmbtAyyEfWqAoKxv8y6RMaKWuapvaEUmil6Ch/GR/C1Tj9
cX7vD03yjv8L6CydCwoeSirXkS7VMzjDT1VEr8bW/QQYt/RNHOHe36Uhje7VMTXg
WQmpi9R0Bqbtvotb2dVyEFA335Y7IH/nDuUT4efENI0FlouZ5IFtkcbiXIeeXXDQ
XygErNoBYP0y/u2TQolZKGG/gNylVfYe2Hy32rPzCVI7K21PRAd4OVCbH4z9xZnw
H72ozTt5awa+wgk7/57Ki+N7dO+LdhYBA5Ndz/jCNuMQMdmkv9tt2KxyrT0wHN4r
gzpFlm3W9NyuNX40BkPrpMSosXrAtgx3sIASiwvV8mrdjLzWlLVOmPq7aEVV/0xE
95YGelBB4PT3SWWXtt+6QtLt3kyAajYY4V2fudNzVtrUDNXudaQZW0j8jHU2z5bt
SZEe9fDYjuwH5/pAPsqd1S6zfhEwU+xoSj36K2+Q9Ll9lcLbK6wgdrImr0l7d3C7
YDBG1dbtFFeq/a+xYRhbkLqDOdrG9NGvYSWG+6tY+UeICZ2iXQhUtHxzi8aPP0p4
fS/ZNlpwrwBlE8uvqfCKf2iYPvLzYlkWN0G7jz3uaIGfglzB/PUI+L2h4ml1qbgb
yhy4X1x9YJKGTTOEqh1q+1buezR6Yb2Cm9vNrKW9OVEuVELVzWZRve6unT6k0iRy
AL+7x9JOxnrmAxL1/5K0P8sCJhXhwtGYrIhN7lrRNwfW4TC/EQaLmhOKdAVIM6wr
Q9ZK7nPPbtp4YOnzgn1tzggl0NlxJaZpp79Zlv059ukJ2fmB9AnwZbqpTzohOrVs
r2SWW8mmm+2/vGl+pc7+D3IyrrGdaUxyGdYI5AcF5+cDW8zNtUXmslBLhveS6Rgk
zOWvs3QEKdDM9j09e6N1bP14Kt5GRi5rjAxZITI5+9HnzNICtdDJaRGx056N+1GW
vSFhn1BM2spjvrucWZKuR051+gQ75zf55NaSaa6HtTtN+Cy1i9UCataQjJEiiWFB
U8g7ciqt/wP7FmCJZZw6CiITeJpeXImDfTkLluK2H6KnXUnmOFz8jEmmcOOIyz8f
s5sYa9M/ysYpOzk33Cm/z12J7kiCQlhPTK71lymlhMkv/NVJFDndLsz4Fsm0jS3H
b7qKAtwGSH4CVtcClv/JfGWIN4J75LycHS4Zlt+bntTht7zKMFW2AJNo4VL9+1Q5
6PSw2EYKAauKWXdk2OYEqRdTexvTbH7RQ2dyH9PikWy2Oh9/jm3EVYc5j7pdterQ
HsJISOFo1skAxHd4GckTSxemn19sTwqw3icp6kmSh1gilFYIfyVfeUSknDXCxuGE
0jpTIqo0C/U04DJAI3BY9yc3x+pmMZOJnQhBVHdEbnweCMU1JsaUie7dctEtCB2W
6SASl8vcvBAmHje8IsxWpwROf0A3zwwaSWKClMfPu2I131NPzKNLrTqfBhxMpjzk
v9hz+Bir4quBamhftnb+13syoFB+ehCxOiL9MT0P8JiJff98TOjP+FDbK7UVR0Ij
K+TFlmfsCpGdLdvEOT0lJu3/2+mwYOQG7f3avrTJhmVwOqWiGrEy6uslkfS9yaUa
N/i2rzL6nTqIekXwSKJIyaRXSY4cJSsMFmba0YbMj9MTyjFYggoAoO7poXlsibTT
xw2JYJRleJC1Er9PF6PRQHBM/X44BG9MJG3s4u1UZa4Z0JWavTX235tQOw3FmX0s
3VgQlPTBcTzmaUYg2cp8CpIPkuryGRksvqP/Y8I+CO7Y1Z0n0B7juB1EBHh1YGg/
X6NSjwpAq8dunoR4HYCNuhsCsCR1/Rwgeol6iASWCnfXWwNTLD4JRX5qaVqRvt4W
/+o+ASFw8422J7FYpjFY88UmNStEx/9WUUhaPiIXbqjWZzTSjGNgR6mcidhnjpaI
ZPxwL7oqH7NXXwxUZXuodjameFAlBWVmK0cl+wFCkTEsFQAsd6cW71LbXtiFq5dm
lBxSBr8F6yskQCINVf4ulU1dDz/TgqX34h2dr0bsmx2Qv+4qk1vO/LMw4I1F8s5i
FU0UCG16sRXr0SxApU5uGf7UGqLTeQWWrK0FRAEnUWPEMIw3x7Gz22DSNN8QQ1sQ
bEXKEFNzPkrlDQM4bPD7xBqxop77vlP5/w9wmButKlzPEVrC73SJD+pm/W4yzuSo
gRXtsgyL2NYHZhCu4vAivoIp0lVUXpf3jue9ZzNgDcn2B5yFb6baOEKukRUv6/xI
WjayG9q3RIj+a8s8Rma3Ven+U2ikATJKdAr7CvANaqZsHqvzfRKsDYImkoJPXR5A
0zcpObNtNJ8vprLsKr1gH8seLTRfDYWXr6jzjMDzH+MlxMJ+NalIW0xsRWQeRVoi
j1gSmdBmW/52BZyh19bmq3/1mba7J1eJaJDM9egj5JDaw86PZnB34+OClPpStixi
9IAex+pWsvpaMfdHDdUQpgXoMPZTW9OAusW48VBaM/1f5Ptjcinfx+xPeV3MtT2A
HnTYM2QMPdknsJ5NJCJpiVGlbkUwwHxqHCDycnk55OjVaNCdW3cgX8Bl1BzoXh0i
T4U2YUE0//mbm90i2DtsiDgCtMRMYMORXuTNtbdkPgJr4DHAcedYFUE2+nHmUqiw
03sIKjnmaJ4roNEj5xPLw0Z8UL1w+9BLQEBywi3Mq7YfMf/URoIbImY2M9/qxZTa
EAbJyu8wZAAFdCWRVXbWZdrbva3NOK0f1khChrqIPSskgPyucbMYWq/1ovouMdH9
KmBieCVZm5GtoyEFeiaMAuf2KKe5L2dh8qYNd8/YOMbziRL7aOrFcJyTml/moHQR
kiTieV2cVl6e9fGBDjDspfX2mSWnZeLvL5yfe+QG4ZEQt/moY9lwWPZMc5WStdpT
srFlp46G9xly6/hyxKIrESm/de1cDDApHnqAl/PotP5AF6NCW07FiDsrcpew+uKE
3OuktqPjBkD3Tc1Gt4SZb1Mda+8DHT2KGmKrknHwcES1e8mr9ErEgSLrs+kjAj1N
BV6so8VM3G+WIhCa0iaICQWNHxBLAvEWTwtkhrm5YeCEQ8tBVFNuHiQGm1bhHsJy
VR0X7psU35aBYOBjBeYH9Uaa2gA29fwUAA/Kmv/7AH7Gcb1kqrUW4wfTJC/OVybQ
Hackg1CwPOdadvKX6JVA/jlVMNTBAz3P+YfmVhxykdDKrACb9Df+R/n+WHDYiNve
bVik1MhTFtdzjtZWlc/tDhnGMpr0FFPCsRjvWMOnFMLDehLEKA8HuqfxKE5xsmub
ux6nfCJJAdKQHMCkBY27Ltu5r+Y21zdaA+J+q2PiRKucLvFz6RCRL8wIR/h1793A
PbVg1Jan57QwlNFGj36o725zmKfK0DkTRHjkhl6AMLqlgtoPLs2Dg4NKB80Z4az6
ABw3Ad4KX7RhP8PStC9q7kahC38WnDOCIlAfnM5yYW97dhHR8+7PUNeLzf8PDUg7
GL6l3VK+chvrcDqKYV468zufOlOovrC557tQebx+6mzAMuUKqxFHMYdKhrjLQ/CT
/9fGgnu171NgVpykit7HBDUypiDUKvaVQB50XcRyu/WyPTUAQwr6J1066yk4uwP2
xCN130YAoCAf0JT5QThIBL2SZzX4+LzghYktVGj4b0KyzcKCWhTpxAfNW4PYVhyo
5bv2P5YtyGkujuZKb7UlMsF9JR2PNYipqj9ekkblr0XoXeaxO+Q7+Nfa9wGXz8Zt
So2eG3148hUiZ6R9SHnnqo1BF5aFeKDlUPJSuRKDB6JWFXOIg1zRJaI72dEurwNk
MRggAizVhovTEhUxbQinAtUsF2mRpt5wossJE5PsEXyaoZAe+jhkLUSfJX6RhKGd
2sIoQUJUQgUsZiTEXxA+s0tuiJkpralEyvqWFLQs7ooU35gKN+PqELVDl+SK4l4u
SEt3jdnVEWONszQfJpAmBH8PuMSxD3Kalv7lJfspWWuexigDLb0eLi1MFNczH3Sl
fbWnTo4PsOFepYOliDmG3juNqWmY95zUk3LsJo7WlaTGLGavmCNDGbdkclsGaB7m
pgc1wOH88ZSYAbKbC04PMKhvX3ooAmKXWbF+CsS9eklxLixZ4Uxcp3rhNeBglfX0
sUCvKvg3OBcddR+X1ttmVyqYzxwpBXOKOg9A8c+lwJbH2j1R9TgQE3n5XVtIHzAA
OGH8DOTxuKjXGrlBmBV6ilvlddu35c9VrZfAlT0unsxWRrTkPGlJYx1BjYfSXBrT
og5RRsw6TshISfdXjpaHWTkBFyUalb3q5PvtNPVwCbpVAqsmLoN3HwUwd3QMZjd3
m5NLdzHu9X6G13111QNX7LqI7oRxnwpa36ZTrVNwCDiORhUsVOuArQsKywGVHPGs
EwQNyawBbK8RWK6M0P1HGCuoHJ0WaJFuQXxMBbygdYNoe9NK4svGIUrcxQM3CN4L
ZWd/B9zfmR9NffEALUkBFLHe5l/uSaSxeHaqo6g42+hqLH/idl73Tj/E2TC5Z6xy
7lWk7rjzBI4HSf6NYmr4byi6ysiQlxTMACB6rJknF7MteNHrvX9SOd0HvVjnYdhu
CjQ3P+T3ju0VdSRp6Gw7kTXvp30hr3aue1QI7437Dn6uafKJP416FyhlGC9jPU3R
cQ9hvJqg/IrgWWO4KgJcj4JHCeaaEH5KD1jiEGBSnMBef6ebxref1Pvde9ua47ti
+JAlAFwUYJIzygO3IWhTCLL/hJyHG8bHPMqtke42p56zxJuRbc0PsBwqvJ5Xb8FU
YivSGiDhwqZs/1+Q3VUT8WZOrxU0hFZMue2yDEVZIj7H5st5o2/D/ZC2ehvW5bHO
nrKlJsYpMSodgk6xV3//Jcx0WeBujnwbnTdbtXY7vBzC8rftJ1oIoRfe9JXHniIG
/malIjUNYljXGy0qKsvO4UcPMO6kUs2Da9Wen9LDZ4PTbiXmvH0H3mw8CsnRqQZW
1oVPkKmtW8N+Z1tocIn1wV5xzrmiN0QLOC8w3y+PwilOKfUnoNCzjMmWMRm8iAA1
gSWYFh1fgN3zRrUFZH3P1a6QpM4f9dP0aqFN3GX8m0AQe4CDISXbQsq8jCBqqacS
SXv36A+lom53FoxKH0nyhu0o5ApdBE1QsY0ddxq8nO7TpXZt3rLhSyJ8Qk2zgC8Z
8ppV6CFWzn+cDh83TSE/46QGnppD4d8cV4FmxSf6dkyOHh0lrxFaOed4brb2frNs
DAVYOOFnPYJgk7WXNsGvL9KQ/+gz83dPIzR7qEZyJqsW6beDayGOf02YPOWM4dTm
Hxp7vRPXmjlYsn1SStWBU/M8Ph7cxw2De/KaMQ5Vo6IhqcTJUn25qkEQQseO5SNE
XmMWf2S+zx5Wonh6VUra0u1fzf4a9rqN03Ggc0N61fSVDx/+4lyC0f7lmdjohTvg
Sz7GUuqlHZjaZ8icyd6W9ygXQxbGc3WlI5UBoQZIf+YexJSdtL32ipJab05CoPjd
nEpoS0hFwhu3k1T3bgE5EBiPp8nW3VS3kGcdd/9Jd8swdW+E7bpRQwHjewaEaZES
ghJTscUyq4OUXNEym3uBiys/E/7k0SNMSlSnVopfv2ttZyeNMO+2sc6UwdsO92Zt
NTdEF6GPiWn+yftTCGMckZyO6HewJ33sBolzF2cRtV03/M8DGjUzNSXPRYWUMnCW
Bol202nT0/NB2y7vFxCe43rZp+grdHVYM18BuVzCWMMaeH//HFCQ5RQ4B4TGVj9Z
A3FEXp9wNW8/BgqEWE+22IX5pfFQLGe2UGrVOXDe32h3f+PR477CRqHyybIsxHmy
p8uDtfwXG7ELL7/b1ZlggKaSRiBAtz0exjl6Gtut7PFwbgsMiBUzatcGo+6VGR+t
/6oZ86GcNWKbGgF+6X74Jn21/QWDlp+1lIPkRqkNFRDUdyMARMugpUtAOHUc1I58
TcFDgi/1x4To64W2kMUvYZk0EMEjcpB8g+V9GMryTvYcjeVH+g/1RpqnAzbErM4y
H7e0jM+rvnpW6/I9WI6R+n/MN6/ss3Iy78jgTOuwSn1AC+TW7JlBZOVIcWk/4Ap1
7Nz5KAc1fSZ02bms20xLa+K2SmEDdGx0v+nNWLLbtckxrfQURd7mzZD132JHB2dt
yKb3pceegkBXH8HipFOb6XaANVYe/iXemLAweqx/Y/wuFfjl3qEehJWJo33V7j/L
nyyQQ4N85rEuLZCIIIG8PdqeiXnZWS+yyJDscW4vjVC6y3QtOIuNwOkcwC5ht1En
pnjHGGRw+YkN50LHGv0WHG1Xy1vMCNt3LZfuAVwV6h1dxWyaaj4NFHQIws7i+hUY
vFeLEbZU+SJ4O+Q/bVyi/QPytoJqxIhBpQ+6i9/DW2PXTI5MyHc41ywMP6PohESv
biDguglgWPzwyf0Yui5V7vGruBqH+QAdlf3l3cRT+Tc4GKqvL+plHuFtp5oJ6CgE
rwSq2XaN9fcLy5nfr0JymviNJfmKp2FW4IbVb/1J+XKgISlz0Jj8FhD0vzWO8Jp7
UeXTelRkL1PLM+fij8hEeL+6bN8Hiu7YL+8RnCxq647jQsumjEbVaLAyEJAZqX7w
MPdgFB/F+rmnIynWhklvrz3vQe15ga0xNc6yvCrHKFYVDfFU1BPRxzR/vAVYS+yQ
QKWI/n9plvxreAqFRCw0f3bhZmCVQNH2ZGamfQm0Vf7cC0IKyRDpZZhYdUV1VHU/
+zDJL9T1TICqOn2YSauHcr7e/IV3F6lxv7Pl8YUjGJHB/LSXBFZLxUfzBFDBUewv
FxnhpYA9bMXMvgGCBmJNqnhPIR5p1Lz9F2B4xT7gx/ycWxzs4b4TEPiVCPXjLpQ8
0fdCvlR/r29y+3KuostRESrcKS8SP5Qzq5wul+OQ2ZDRh8pC/9mcUb+NPRpAqHnt
6jASLxiGU3W5DS9h+s7UXwGK0Ug4/ljIIg3IAwm2rgS0xaxtQgMaGiUyJfCyQu/O
GJ9+Y/iXiH/p3cXvd0UdI4KU7YovX4+B82KmYAWzC3HrADYLiIO9QA90L9rGHN8k
D3m0+Euh/io3jfebhfN69YVjaK0L57SneNDxBFs1gW2KzSdNuJaOBE0hoRTe6IHf
f6FadGV9/eiov/xxHj29iqRQGkWgoSNSrIFFnVv6aEMRaDdL1qtpqqdhRirSMH8P
5Jn7NB35NCIoMtvYB1j0bJvcudFpGG0wVWgzipHNib7FU5sDLg6zXBZR0QTxcha4
/P8F2ZPi3LDGp1uxCwQVkgp5dhXyTNHT7k/IQJ9mbRLFHfeL2sbL50YCMfV3vDmi
ZFku5/lxqYdUebOuOCqXoLlVoBNVZK1nDKnbQzZEam3gfQBTsaR26+C3SkRr5mD4
Hqhzbkyio1gQ/ac+EjtBvrkFUQkrA1VqMiPFi0b75WONiU3eucT4IP1t6XNTKt+f
GdnTrDVanGSS8jtRynVOKOmdEkMeQXu/AzEqvAKnstbZ7HqKY0XWN1IP932GOJpt
9DB+RcjEO2gDC/Q5BJ3XsIMhTm0dVhSEd+5880AoQ1mZncZ7tLnXZiTJEpdUeR/I
RAxeATpTrMmZm1mz8Z+ZNkI163kOefCqEmr0tXC/hZS2b8AnbCk0h/on3YNvJP+n
opS0z+JXO4Nn9scU+WDEhsKsPNNpG+wzG3IfdhUbKnskVR9+oRHqIY0H47IR/wA5
IC9A5xRZYxNrnFCnuSHQ0xA0QFawfsI3JrZXLAarTNrVFNIT1ICxJkyB8pkMwxHz
4KA3fOjCm8D75pFc6DxOJPuvZ83GVMp1dgzhU2GNTvqMA+HnmPlv7NkBW7nHje+C
55fyQmdrw7Sph1rBzA2qQqT31jCjOTWeMxgIskOtRDrg4aEbvrmpPV46Nq07lJEO
6wnoBFhKKk9SO7rcJkTaQ6OGvcja3yt1NEfOBg9h2tA4bVsJDrmXiafEs9EMponP
3KSw9VKQem1YBoGj6r7eAfy5AIriSyfKW4LAOzeGlml9hOGf68/e7PGVgkEAVb1X
ZZA/38qmBDXOhcgnZUnBxMjj3E6/sh3gwNyYQ5PuivtrPH9b1tv30f13znlvvWNo
OzEdm+9Z88wfDedQc1wtcdWVJbnpTw/OTBgCqnqwpvC8UFDG+3lJxG+Gh95yvxVS
W9W1VebXg1hpLp9UeI7Nn+Bo+e2kl2P5B8tTA91wo2+9KQsoa92e6KbbbEdvgG9t
Sgz8/0R28F1YHFnhY3IkIWKowVTHSjAFFB8MwLfbIPWkHRCcIJvbc3NOrTWsMKOp
bS1FyrocU9wHNc4z9dx6oPjp9lL8KamvcWqqKzrpUnXaLYit6ebPaR/FuvVu95h9
3Cu0T2/uJ+KZ+2LsEVWEv1ZRNfyowEoDNvMdXgcLo1HvQHglGTZuwjFp2ZcwDxHO
12icuFKwie3rZNQobfxsFFjVi6Nm6oh7px8y9t48Lz4CHYnf357G9EUKdJ0mMrzr
1ZIfAAL87Z/qhLWIJpmCz+Kek0TYNwIKaSM6w7cQWlp4N+Nbju7UZTeZQHTvnEbW
dXhqbLykj1/0JyobIYXN9yebg0+rh26YUGssJtyv/caAkn7IzVyDPUODnsW+OkQ7
+C49LFBWVoO40yhwMM2OGpDfsv3t3WcmMa/MqtnmMi6tk0z1MojAIgy2yWTQO9FB
Y74DPBCluOdqOMY2HeQ+MVp1RIMzxFffOp5TP03KGIN01PQnDtuxJN/uSml3gHno
bLmxfE70jkpWZtSCVofApvNH/GNtlrgFeZE5tXghL5lqmz3Jwb9hkn0sjz1QDIS0
0+tlsFqWyGy3GzzKZs3aBznv2oTiOR9bcQUVbKN3k5F91dvlN0ULn3KZLOIItat9
WfShbhbJIreo9bIwCdfQXmiSGCqruUfc3Z6AEQjES3UUIcYXdSW1t13p8Xczfsb2
c92kLGlEQFGExCmxzLFIiQEhIIDD6LtnCZ0b1EBP2uTmmgTGO6NxNUiYYih6S0hl
vYViic/k3FfasLSUv8zv2xixRkfXs3W22XuQzz4tphl3VnV28RX93LZyYtAxlfcP
E1aldW9ElmUEpIxC1txtNK9SZtBGmCuu3AhxGFeGNwiM3xKtY+VlLfa2oavcnGzx
1qkILe/5mWV3oVNwzJm93wtTPMql/fVVBzalSvR/6YcrMgFf2CT545oIcldXMcdn
JumstmXtYKMqAhmCcr72v2Y10vpqLBQG3RuSanhg1SWAB0HJzB0vb0c+/jilu2Dw
XtENVYC8APsAIqLml2pSUjHcxN3L5WLlNUSa4s2z59QEb0Ni3GbnpvUYOXNbQAwj
9l/GFxwhu9P4SxAKKEVWAXMKlU0PADUYWYenx+5WA8mnSHx8NU2ujbSzquVEypDz
/sThrMt0SOWZQbcElSgnOUrMXG2Cd2AzpcfvcdI1G5/piKAQAdQ+iSJb9Tu+Fu3M
qKOiXEmjyVMpfVQjkY8/r9+gX9KaGrTB/33EaFGmGEyw0xRuuOVfSxIDQhKakGh7
qzSE3hHoTN/gHFn/r07AxSQSOk3KBZ3WmEZIPiNOsNAH/jD57xddP/G4Et2glSSU
uqPT6sULbuvJmqqxrL5ce5Nq8F4xfvN19v/sA+P0xSub96O+sFJkhK69aHdqp+4i
F0WaWBmpgndBZGXoO48XSzQ11NtauoBwd/kpGgbCwEp3AmBqYgWMh2u8+od9R3S4
U/sGfX4pp9YgcnA8utcFt2BmwkMQhL7kIbw3HybJYMuhRR7j9nMJGOKTS7fPnIgb
2ZoQgv7arRo0Uwwmwb4ej8Ssi0CWM+lAZxHLpYzT7Gy4YBMjuTK9Cll6LWsyAGgV
Xdjo/jDstBftfDoDKTGlNMrCkMp3maEphmvxbhHZmNzW8ptH1tWp6rRovlZiObes
M21lA7Z7BfobtIFdhub/UNVfP8VNlO+DvpCbl2XRA732gumN4qwCnslyqBCwrqQA
iFdcUaLsFbZfMSRBRSkIKJwUQ4qURQXiOa7z+hs0hfnLYmaxlYp9s0rVuizPEiAW
QtAdp/vBCFbJ1OqSt0RFDvDkO6pJz9Lh8P70xKTP2ECOXneByhMPaPo5pdNrNJZU
MoF7i2g3hkfPUhspu1ShJvI1K+ESb8T3fAViEpufzs6SZ0BUg2Fik8ElwTdX6kUO
7aGcNzeZOkPEdsRdAmZrf5jdhrNqR0dnaZifB0DJuVIXCi/XpWU0GC7gRXcUwr78
1SWM2bowoXGtqT8fH+MhfhJFuST5Gj5R9Wb2r6a4EheIVTxZIksVgiU2gmY0PX9l
nkh5eOUwAfM1D0Wir6nDX1BJ+yh1zS1Kd24isl4v89WjpluOKbIK+lP2PnhYrK0d
oM6bWphHA0U0TvcUPD7fPyzhw6kFyXsc0RRreFURsrDScd1LrE98QStZvyS1z9qc
ME3pDbiujgZC5kxQmOWNcX6XolnMpXkc4KmWoSfHUSVWvhZPpsdB8fikJXbyXJxL
/aG4FunWgQEJoxfZf7zLarzIdTVG4t2tN6ZpcM3TkBQFUuFIVuxfcEqi2G69hd0G
E4t8Nb4YYQ8EynLCNeb7lpXMXfFcUZagXEqX8VuV3DT1gYiwIXPjdXIkzrTG44wj
sJ06TUpF0SIPDB4nfoDdgkKSaJ2mh9k0pTzX91sW07LIKg10rQc1mSnw5pn6TLVV
GeYUgN1U4QcbnZx1imVaqyI6+a7YSyqIJvI+Q1FiAUb0nEgpsN+A9EgmT3Sa7cyr
qiVkcoFoBZAf5Kwgzs9kfOQOmdp+bYme3wEoMNvEYP+xYyITtYXrQKhFuR9+GvPh
c1V81FWSokBUb4RU2uIB87xNaqwrC2bxhaStUpJuVxhBWjPvCXI4KR5kwdGGSxWO
jKVpI3XTNWFgZrW+oFCFpMhox3gUSW0ZChdPC9tpm2/QRITTnRpnlBHL4EJX/UFz
uWKReDAsvRvy59wWSkc4RFw7KxxZmgYkxPOV2L4v1nN8Oyin1iLOj2EsYNHCJXSW
SWlZheNSY4x/frONrbJhanTx6o6Db/PYgZggVsnIvmfrUVQGcdlhC4sXilX0OI5a
C7p+aBCv1I58nt0jV1nRRHNs5HQlEm8IkyarmlGAyracTmrAKROksxNbcDaa23V+
W8qVEzrB7Zu0M5RsToPVWRZrqX5vUcoJjvpMBYEgZI+Pd0pBcPd9913V4N/SRSh3
ypQiPsCMXwKrqQN8hsxSCgZAwe+55O3SWcaKhYfZhmrfYaoTzl2V2jcEaREKKXxt
aedNZYxctURZFdY2xk6/f/ovzBHBRh1pXNNLkis+avo934X82BYnkYn+SlfHDIoD
ajWArRryjZkXvdVJS69Ewdv+KSqSNYpcW2COOEww+2nh/9VsPzQEgYNBoDbHVOS2
P6L1epOu3F7gzKeiRmmt6KaOB9Q6KG2OgG6phHfrQ6VUEV3tYz+cb/spZA07wXUV
V8ueXfqBXK7y2nvJxo4kJRDmn+TIodUwXLtKpzSstebu2X79fxlwp2k3ezvw/GmA
O5kiWZFKuTAFnj1Y7drWQ5mphrGFfUvt5XpA2hKUgMgxF+R2CBJTc5W4HfChW/bX
PzfIMadvNxSobra96hjakG92NPkE91vwUkDdowpxv/Wf5+JPkJOJe5LuGX21STX+
AgSUlMFhTn6zBanhsnTBWSDbl9ANyxoNvcf+wlzR9o4gFFe9sXOpO0cNcrw6XcXV
+pe9vYq/fiXqCL3LUA0FaX+6Flj3mrEy8qbk5PCql96hQI9ZdIRrRJ/up1ss2Yec
QBjvkgzY8aXRB7xNrX4lZRUxIYtpKtPUrY8t0Em9oh7EzPIcuCZpJdc0MqqUpPUE
8HMmThs6uRXeQDwywDM0fr4Y3pJH6+4aA+lnRUH+2N73UJOBiONYemzu9/dZV40e
qfzId2UwzrOE2mfycVOb2WPQ20rlZdFdBoR+4efyWzRJMgikGxPgsCaqSI1XEbY3
SNejzBsV3XqnqQTa6PA8mjHlK48l7nsGzG1iOLWZgU27cXcbMLuCjoc/XdnVppbt
9/eulubir0jbILMQ8Np/P642zUG2hPGF3/qnJ46UWvS3ouMX9fyOwrLs93gplxfe
apRvm4g0BkWh/vChRbJTLlap7t6JFsh+y4Lb3jlV3/Dwm7ChxNQ9UCYzjBx3tDvX
HKRE3FHKAb9uzR6qCNE7bsf/G5HAo1IHJU3+rlMqwAQ52stTGQz0zoURJYgkLAH0
J66XyyIVtJHcwc+b+Xfsg7uFYvhJDLydpz3a9nN4zDHdKRSpp5nJdIEspgEALUBi
mlJ/jhmJY61DfF2zxGbb9CEk5GZOXNJLeLVKxhE6MIFIHJWhTJOOb3A0Pf4tlF7b
rJRFY+QwU7Wd2JKzPrC0s2Bdm9rDM/XWuBayoKqxqcbSXkwoLhyeYDXDoCbHbH2z
VspkCphG6+FoMMcsSa/aA1Sk/Bcv831a8k2+wa9dtYUA829Y6BU7U+1l21TW/LHy
uS0V9Z6grHRfuVzV8IKwPH/IY52Wvll7k2/TmzdxOeQVcaBB4YW/MNlwsuo1EWL7
s208SGvzLM7IkpiyUmCtGj18npeY42b+iXq2SHqNpAVHdeVvrYmTRmDvbByAKXzw
Azl/HHAuji8PPf5VoT10sU++X7KaVg0hHfmOlSfclSoKZLoaJ3Rd3HCXZdenbDy2
1n5bF0BwDxmUcDl5IGxskMnnC8xGxwR7sklkxzBEDdIEwVoRaDwfFf/OTFpAt5Iu
W9zGqG0w1ozzIVqMwmx6PpSSkZ8lVV2ShBRh9/kOnmSMu5dkw4TfIf73FaY+Ms1t
X61c4fNt3kLVOmSX7/kacLLyXsJUXqkL7w04ZxVu2y+aA0vcx0VtTohYF7JN7d/1
2prxZTxOKIqiJHzEOcWqkkmsrQP8IAisbPzhu8P6rOhmxfwEmsozvQdIGggv7K+G
8kGTjsk1UpPRlRSikM9tzZK7tk926jjGd9AD9LFylYaxEsGpCDevGzdKSxnnXWvT
LvfchDV9CyhrXiTqmU8MDGBuD0P+auRXyV4zpP9Px9uev5DqeAlAN35m4buDQK73
FXztG58NN4PAYSdeCdo763qa4M8xBEKI6MSinXAR9aYYzOzrQgqJALyp2yPlp0wO
YyWei+Yqrhr6eGTlSya9pr4m96+CjjzRI59ghs2EPh83NYSflmyF9CsOikSQd1Z0
XSvIJieinqIXswy271aOWlES0C6adXgalG3dCzSmOLtXhWW8eY2/bFU9kwRZNeLi
w8MKCU/1JsaG+G32oil53PeSUa8bnPX2kadE1kAcCovUL5kCHuGC8kFpnTmImcj/
n1/BrmSXHvtrrh0hgAobVPn4tiRfXF5VuqZxzuMtGb0zkWVUNIkXmM6WcAxyukUL
IFFtZ8bh+lN9aZAi1Su+tmuxco2RSJmMJB1eRswcLL+hHhqVaPRHOYgIeJgVg6w/
bzZBgfP2F+zy+GGLuYGbmJZhg+2bg04WyS+ND7d3RqezMId0SM6ptUabRP9F3V+x
hqDrnOLe6hbTwC/F6IE1sNNAHnqZmuy3lP7nr4iX8XoWvkYbdSBGXkV5tVgylJUp
xQHzKyIo7cKYGBYCn0is8nNhFBBq8xddc4jEwhNALuNHl+iTkzuelbNYRMHDU8Wk
MtJjfDtmBZgtPHuJ/XcQNmxZ57PaPtgxlf77KOXnfr0TZwbVMS2KD9fCbYsdGjYS
qkQ4+jLzVxUZA3ETaVfJkVmd9/o5SfEIejAKa5oA8VXxzvz8yJFxRub1Ez2fkmZr
Mrl2Q2iVp2UVLZ25nDC+oMnr75fkNcYIdSTuM/D8M0OQ4+QNEiRrswLJ8ldahUsY
DvG6Pv/7A+q9dAsS4qkZKWuqX1TRYtE/M1g6D/0ybExJLEIUUEwOvPz+UeymAjuk
eaFtUZ1ekqIF7WIExJ/iBoZ/DoVh/bB4TWtemukcTHHvppT062lrF8SYWnEw7xir
8qquEwJdi1G98tGtmhgi1rOfvflAdE/Zf5z4k5EZTXS7IhwxOEuI4ViXBoz0KqJk
DhlXh5gPp+aoyEnZGKD7NpT/zfVNW5Tjo5o+NC+oWXWjSmjDQ82l8neqLAZXvUlZ
Fjk/hIZzySwzJY8+kvul06TzxmWog+xUjbi3IX1VUMEaE5RsbxuJBKsHG8AWjLJ2
VwfQDLoVhhf2wvv+1Hz/gtiMvVZFgnWUDlWkmVi88J0HNeASnoEacR4C28S1qeRB
4E6yjBVlXSKZTwjCYT050ITJ3mmmfj082I3mf9bIADrktMNR57e4nbSYMeH2LEH4
po4fNgOGPlLMMdvtvRy6caVuy56TePV/1ASJv16RCVImSW7d6DcORXocAmvQgaUl
sejK6d0X/Ty4qiXhaSv954UFYu+vDH3VWaVokpkXpyLV4J2AFo84DU4m4yojwk5e
/f0o0NsN+mLl4c0qo6Kfz3LIjI2PMIry3DA2q9tMdyR3pjNvlQFEqbDDlRzOZUhC
dikQZ2OpssszRDYhdPwjBD8i+X68xs79Msu/lWURbuGwttszhMDSJt2e9I1QxaLj
OBTDN8a7g8t8ytuXd+xFmbYKPs4UKh+VSOh+h9DmM+0Y07k1EEgOrEq1BagKw2ux
/DulG4x3FsMqMRzOBwNpdr4tUgZ+ORN86wha+ig2aMURSekD2C+VXhoSagZNz3wL
+oKFmXlUwwmZ2pfQoPI6b/Op+gSt2RFFYi5UqKOaGOnbwaxRYQ7ao2ymnz/RhGkC
c8onmd02sqLhnU4vpso0stA7ftJ4zqzAWrVGbXbzA6dI6xjtEXqoUAI+4JO/wVXi
MLv3cSdxryvhZ21+3XErQ55cKloBdNUn8pqwZl2DXaV4KOR76BRWKLU5W1+PqCGP
pzNGQr1IWPJIYGAic77COAAEj4pY1tULam1saUpVwtfbGVIzNtm14/aH4YdBQO6K
FslkvEijJZD9AZovM/xQIPSGf7gloTk83FnqKcJYs3ttbg6PLa0SVIuc+nLmx/lX
vc+YJWiDc3d0X11pncv9pdmguL4TMneo/T0ud1ymRL0Kqu8vPCrnaJpUZee0BTvl
kONH9N17v5DGT82WF9IHrHjN1iq2Qo47RVqOmu44sHQvYETmWIV97Z2+rJYrkX7r
h4M98pRlhZ82cRTG7j70K25Z+Syd/JIp7iWtn+0K8gWJ8maF/LFDewaRPRxMOaQV
TfMWlVXHWGqpz0O7CqD1MHP4qCl3iWeMQMuwBP+gJvqM+m6AFElKJtouW/tT36lC
omDOvmUfPIWXXUX2IMMFPIKNWBrf+Ko4JGLqESTIfjETJ6/VKcFHxVoTk8D1Nvk/
v86nKcdOW00H32no9AtLFT3+4jy7WD9EzaswDycPA7+tZWGzEv1GoQ3ZJVxxnubL
RIiVFt33cROXFEvLWVhkLa1Iry8QwS2+urtYfaUQP0+aO/2qwC4o3eNd9JRiJUmp
R3riFOFMwgwZNT4jb8dOWTfAJUKxjt01ypjeGlg3pdkmoBoa11lDVG2za+10ncvV
FDUhzhunwuRLIpW1bvPJQWrUtKfwt0/qweHphnWfDcaWzDvv7VcAUtry3ZBo4RWU
ObejUFhLZ1mPUyC7bTEvTGAD6cXvSaivVcHVumocT4kMs+3hwzaSN22pMpZNwk0e
7t06QCOc/7eVv1cYOQMEbQywN4YoxrZa95R18AMG4p1WUzmYCpQyKa36vSp0Eda1
16rqHWfOSojf1rD6f8brljn1ScMNdUw40WtjF6LiischMAk0i3BptoZV4Wt7M7zI
XFigG63hflv9bi1R8ui+jDvHtVfmVN4rNPRWVDid+Xty96mPLGelznxmFwacHCvD
vUb9JKjzm4oQ/LuMv1I/UcSz/l0SOSeD9kDFObJH2hqpGmDsMBdtw3GWMMB5M5CO
zjofFqiSO8G+Jo2UNVtnqKXr49CeDQE7RzGUF0gA3HkHnvIucvU4+y9ukli1r1aM
5sXrocvk5TSnebQhxwTtoqMEN5XAP5QgiY8k4gkH/GJDMD6NOZE5HOBrNO6a0ExK
rPGgqjyAhYruwOB/LmOjfeypItoJcb7s8qTnc9RR47loQNkPFtPsQYivXgHBfunP
E86FOCcPih5ZRqFIVxeiz7KUM3+sBHabKUgIYTqnQFJof8+svh7up+a9SGdfmq/U
ftd4AkvpG1a9W6mjsPxfXO2kHZtV3hLH1eQ1sWDI1XuKzRzIBK0+pKOO482C6tHB
c7FDII/PlD1B9b/t5JaruEPQ5uZt+8rSTnGmrRE0DE/cCXnHSHTCyeUCg10uSC39
zr6ccoF9mL3tWrlK7aEaIDHzyuC8nF4Zkr3tpgHZ6JvK96qMcm77HOzAghv179VF
/C4fvNR/OEtW1k/zR5XVU+571BU7UhEPcd/hdRaZ6SaKVoZghcgLhIas35dwQ7HH
mZWxW+zfiTAPnj/f3ZJgl0VPTUVxTisvsre0UFRWgGC2MDCTMUd1fWkAF00cGQhQ
0+ar8MR3xKsifbacG1SkzBnjpdXweDRWwpbzIHesx5HQMxyBhE+EahjMMIy6Pqeu
IrjN0iB8x2OUjHBmwo0riFl7eanH9wilZwP078R738msoR99DJ9tVwlCddbgZLCF
RdAzhZq7lxd6ZvbeT+L7TMAid/1Qo/cI6ZqaXxff4e4kP6M5Vb4ZJhrN5toEnc/8
oYWqL11tKjnYoiNCFhNwz8bkew9lop+oDEMv1QudG1krwsrsO48JTghAIwLOhk7Y
5Z7l1evKi7TIq+/5Gdfe25i1IO9+opXch0aHWhCh8qW9nZmhAAad3XZOeg3JK7Zz
FBhBJnOt0RkSvUbYU0kg/RqVVHKOHbMW7vCMPBCZAV6lR4gD5Fq42zUUOiwmuncd
X56MDfRtRQlEE4BZhmJmhPpgD6sSk6fSAaETRwkLrU3EcKeZOrypJ5Z1Nm99uKVY
xT9LFYaxpuxbBPsFN4J05QsZLZ5Cyc/haVFFf+WAXGn/ySEmqjgHHqziSisRN5CI
ssmuMEnrYnNEmegbP1TzQERl2BMmR5qbIQiBSZS6Gvjr53ThBjnyGLF6wp0v6Al6
hVRzinskDvCK+tLOlVP5kwQqK40axvnPyxo7lEU20ac81PA4rZ98Gs5QYyhYcbjn
dXa0yqndU6m35ifxt9vINw02++svn+dTBu5QHtKsZWajmDpqS0/pUPFPEwKfL+Bp
oRENFlUP46Am7d4arLTeiV7IeyMEywMTUmjxgdeMW3vACXf2SUpcv5O4Jkgt7KLQ
DLpmssAoxG7inFtEvHxxm0aXrg24tHkbfWbPwR3UNMyQVokZr+8E3nJX7FJtWOtg
JtWrvLn4MsB0sK/d3wBO3iT/oq2vrgg/7UoEIUenuGd3XjRWl7nQKQDmjPUmXxvL
dQawR1ELGOZ0r/9rraFr7IS07eCYNqSiGz0Q/s5wye+VXYKiptneY7BmzjVUvGFu
LYLryI3/31r8RQZTlnsBb8+OfWHduZwR/cGycDZRfGtZO9aeFxik+koU4M1KTgYz
dQlU8lNCGMfBNQp0ifFBaonCpgaewM2zMubxQBtffo2yS1N8Fcui52TKFjM+Tgmv
Q57VYkyBgpiXCWvq8ejYxwOIiVShN8omVJYBG4CS8zdDEV5yahJt8Oqb4c23el4M
YyOb5LjaJ7ffUH9f79ZTbo/BHN9sfMLmAzsyyg1N4aOHKgILZHqwXlMd1JmFAc9K
WwYUMLzsQbxKK23vGLjonrQzRyFhdSotLS2arVRWqGUNX4HOodBevBwgyhpuP6+u
U0pNkwIQDiXMmRbOsWCnPC5nnd/1VZ8yFVAO8Xv5ov0hxn86h9cmQgb2P4i3DY4R
B/xSQqjHgzcSEkkiNaKu6qNYhy9aKUol5iDS2z2+F171aOdbMocWx/i1eBwpsYrS
AyfBnWtJULWecwRL7RWQmLV3zcELxQu3dk/1tSIdCVUuOTF4WgiFHZpjvKSG5qL6
8oWTPceipzJUhEOPREn+YECafEE4ah4zep1b6e9antdnnFbZSRcMJDiFlTzUCGFH
F9giuwJvux6XmW/nJHx9WKDXGKBxRhIvnHqg31LVSdCNmKJHfFHZd0Op4a00iu5Q
z9ZlDR1XGUVF62BccN4fnPclWrMO273Fssi9vJFy5Ek6XQ1Q99sEAfCQEPOXC+P3
lEWebE3aeskuqGZEEnUXMTIEKx1manJnaf8jO/C2Dl3OtNTkxXuKotXy+Yzqgst/
OqwQuP+Jne+9DYP2LgP4UB1L1lnFKt/P33OxvPyaZs6TF8dcZQoBuYvoORzVqSqd
UwNasKYQZyAI5gl3+Skr0fGukN8boGq7sy1ZVX3PVpRUUr1sj4tcZHxEzkr9ybUc
Y5NQIuE1vQgehQBcyEiW2S9zTQ/cs1KzisLVjuE7T6fFHIITXxiy2XADyUK7qua8
4t3bhOuBUVu4/z5ACQmOHwhTB8+mgYh6KjgdavkG3ofkh3oHu2dcvwIYD6g2RIit
hZ3OxNmGyPjXj2YHhL1FCrVoZgA2zQCT+hAFoJOVSVc5KMkr2ZT9e2p6MPKBd38N
W4LHBZtrS3OT7If3uOEJFrSmM52Xfq5tpSAhI2tajt+ibSmJKUYV2t/08fYExsSD
SRiVxWvTfaToe5fs6CdX0uicKgM+7ou3bRh2rAt3aD4dccwnZ4vY4DSRjjz1D2VU
5NHXcvJk8pQXqdcPHaDzfG6Pn6JdsoSo9RFDuxGcVSqelz78FaF8sqJ6X/rERLpK
vwg0i0GN8die3RBsgouXgMsen1vLXA3mC0VtoMsdMi+HWBcPiTrxcwN4KkzLabwE
zAGqQVcbg9cwMj2WztV/bka1kSZBsEf4vY6Lmvvyi7cwtNsvPqqZODWYrWmMtWWI
ISvo4JkbyK72EdDLIHOKAxeDiO3mb43o0DyQ9wi6tVxy6kbq842CnTHWR5Ic6xiF
GHMkAbRJrJGro+eVMi2G4QexEXHxC2YWXSTtU06yd8vqLpD11LMOHqlahOcb9VhV
Kd7lJEXJr7bv+mf//4kE6TlW4NhGFYWguDZ1FGimTb7/e6JYFfrBSMbTKzgsw2p8
vTS3Tv+Jo2V3IQlT9hRWheLs/nPOo1/RLQ9POpKicflahYrcjnwhb04w2W8ga0J8
C6aTORrGsmpYRrpMmX2SWhufcegAc2QUPMADfkKq1cyjr6DqFbIasmqhICIuuIT0
QczTRYPBBcBxHzbctAV2wq5yU5AXNPrzZjlMVf2FpERraeeNHSLGmuZh/Njv3Pxa
VAmv6GdKmlKiEdXR7OdMkkVlsY6e3tiPbZc0/RIvWJLl5gIuLsRsMQpWLvRluxTL
7x68KSfqUzK6xXVDWqunu2vtCtzBWqrNkFPgQVHnNJEvBhbHno1Gs8ROerEyRF3L
UlP9yeTmNtu+PHrFcBTQhxVCVjVufxeEiFOmuHSAfeupYaOfgjw/YVxg0TY4BrcQ
dLNuYSA/bdxlXT/HM85L/FzD3c2vpexamyrgYgozp394DV+z0oiGoII3UYZy38NL
ec1eiTTAx0e3rLB9+8L0Z3iqz062DTxcfcPc8q6lPpnBqd4XLBOjDciY76d0Gl79
U3miMiqq+ugKLfW51klcE25zC/twrPmWiMuluV9tvHqC9FI58DHtH8HZWSBhxNze
4wlGXvsfi1FHGT4r8MOtU6ebop4ty9BXc17DcCeGFOe4eS8bo6aq07CBwSOZYAN8
tFrOZnjkYCt0tyUFK2W+fb4wlBIeFczVBaUCIEVbJpxqeegF8IQs+VqpNnxr307P
8fWB5iI7KCYyfpbr3TeBJws/VSTOdy4U8VOpE3A67IeDy37QTh2aMK9jIBYkJrCC
o3msj+1rPvlILsMaR/7OD6hSlHLaOVoKhiehfktkb5iwiGQaVrx4HrnoUZWLA9KB
LrWDlocxoO9gCN1j2caCgsho0ladmaQbjDqwZiyby8XI0mp/2kXE4Gqnv1rIGPNB
k4umcZibCOMBDVPfR5OnKDUL1kMca2Ir/F25qat06JynWoy8dWaxdqHkJOsQKM7Y
3qEuAG4MK81ac1LRdRW4TRexyVJS/pBt58TDfJCeYybjg00wlQVKi0jt5MTdKF7z
+IQcEerM7yxQlM2zB5DIkH5kzm7BIP9E6qIY5uOkPxWasaN1IMijk/u0bsWhXWlb
num3Rd548rtMCxCSQsz21RGxzVpaz913mpcBGPh2XxDX6TO2reyjTSYcejCIry3t
K0+936uplPLXzEbYYDn8tY7KISwCQxIRqbUc9bIdDkyaGoKQTXzM2ud9vFDOgwqc
c5JEEbix0jG0Ru0EuLmcaUFBE/NTLpFcs7LZ7IOKePk9pAaYvSwtFkekj3ggj4uO
xweYBUTOEh4fsUuNA6it6CNhdl31PBrWElVgQ6aIgAh6kCqMexwHqchEKKh/ckxA
4w6rZ+E0ErXFFSt57pj5ZHiVtF5277IaR40VoV1tWv5pVCGBYBUaCbqY02BErQC1
KrTEo3yTgh+mKTsnNaWIYnV6K0zA+b0EfJ9lPmocGr5A96A9nfyOKij280X7g7XA
XJK1AcM2NAKfDko7Sc1x/ACaYThL+YUmC9aIUobCkaNR9GNUDObV/5TWptItwoFn
KVhX13FJpJUnKglxlKBikFw0Ik9J9LUWXnGXQOpLUFD2OeyG6LoJmZBjdU15Co/S
XuHdGQyNvIO24Mxe313R2FaLnwYB/u8O0gSZVwAHlVTFHzNo6YxguugFm08X/Mtx
mrMmmbnjonZNpa+auLj3Vk1aFaIna4Q2TfX4qBnIiEsriHpZupKKSgp/bfUM9fGi
yny6xNqitwGsqcgV28OLUXkwDjGtUXk3Ecy0fhr8tKioodrXVRHbaZ7BsZIsonmL
Ho6ZWDQh82Vov+SV2DlcK+ZinwfO6o64czJzUsKi1Cn6EbtJlAHbOIOHlRWOQP0+
5HBtvdRhD7tXfLm1dT0iR377VjIzwl9bmGKU+K6Bwd4O3J6uHteczIlCpTj2ewYv
Rd/3VY02YxoZWajJzl+sLJ5DBvkHwZo4BGkMcwA0Y2Nd4WbucREBCs3srbUeIutO
lIbuitqMpA128bpeUhvXopPh0sI0Iurbqnk6cAPCpqhyu5e6kxBzkF1M5J1DyZ3k
OZ/u0Dt+xRoSgAHAdBwgFBA0+UvvzWxyZQeDsipRNrGOJCzGjDj48/yk/NH409yJ
4Bic5hYenCVNZhoS69knz2sSScvrNkTxSUNqe1EGH/O/ZEbCc0WZOUl+SknLzkNZ
exY1zykrrnnXl/caQWu9jY7LnGajljGWXy4+Qwhh4NHECWW4QQHLuZbILU+7M7Gl
9IlMxp+4cBQ8AN/nfK18jwwPLZyedA4uqPPUDgaPN9F0ADUq+4/kUulINhsbJbg6
OIp4k9om5CY11ZlZFn5oC59DIxY+8sSTqSdDSxfQ1Ct261l+wpoLtJaPz+K0WAh+
a9+7z7dJAAVXn26KFoaO6FIYQiCKhpgpIe2uTvVcQAzclorc57tqJJ+QFSIOTHlB
CHK0nqW27VxVFotIYKOv2nitJpIPH1kWk9iHmLkxWQvPb3n+EY6e6NckX8GwEQoY
Sxz9kqfxfdO887oHH4wsLakKqcyiVcIU8lrg2x34Sf3b42uwTKQ8LpPMCtw9Pa0g
aihKMb5A6WqalyhV8Zs8fJo8eE0WVBdt6R2YrvN1RsmsjE56NPPgdjOahmHJB/Ki
9+Azy+RKehpH1qp5f3gKewjAAPFa+TEdwB3zn6E4A+i/kj5MNsvdzVd5moq5yVVl
nbcIpLA1ldAVHG55CballgYgeSPvIpFO6qV6HHNrVSVoRvr5tS+LgkHYUBTp2DOp
G4W026rC3MEWo1JIgj/i9xnbGZvPZx1GZCVF8bhAorHT+VIFkLjy+NY5qhJeENPg
DqbdHAioYIcXlOhLBD5BQ8dX5FkW625W4FuPgwSJ16uxLu42YAlSUybjNuSeNk3G
pA42IFbrp7Dakuwhc3OeIG8+5RC+AZNUzOA9sdjroWlLyb743INkMH6h0Q3KGl11
IDUnsI4DNg3rZNZr7Xp+/4JHKyla7BUAfVmpvcJtZUoswQiulYjB1LGrJYj0Qwgh
96mWKV8UobQj5ebwYVjfGuE4aec6xQIbwbU8qxuFNXZ8iRJiVCaOHbsRy9JxpS6v
QQl832KUhSC4deICZXfBCijXfLgnEDvTGIYYMdlAArw4R6I/LQnnKZT0S41QrxRr
BeGCkS2d6Bbm9GoNOgDIAaC/9iBbY5+SZ0ZEXjuSAkjQ6/+q+SDh7rMMaDWL2b5R
A46ib1YZwEF21OxAKf0roGwjCev6/R09+TdKd0gANoNriKy4KJgXyc5qj0oCBrXe
8BRW266o9Li/a5W9BHS9x1zlo31tdBwVG2Q/n4t5eNvOIUZQmaLPqSp9Rq6avIi+
3SN1wKXoANusW5/8LaV8n+otLcXBVioMUS0cRrlhuj6Ii4nhNnLQTTYWtMJOXPV9
Ic2au47I7jMuiY7Cp3OQsrfWcx01oKmEI12rM054j1FiYvAymIs39f3+zdELW1mh
DpeFEybBMP0HP3kDj5M+8LOeDz/EkjvRayRVsRKLfOxDYPRaM6WshsG2CHZWyd0R
UFC8kIn7hoZs3AAlpZm162msO6oT+bjowO+CIA7jk1qX27Yqbxqb5oCZfXjC+vm6
TsnVQ4TLd8aEkp+YGgvMWAz+/tMO2S3EKlYTHctk6bp0GOI8oOgeE8t8QF0EnBn7
4M+p6PcW4ylSa0OAnMr722v8zOf2MUbMkzAPMIpPI/LsLza3YbUn9DgE9MrJdlMk
IXvB8rz/6LAJgj2RS4pt7rX4vOHciDskn2ggNhzNMFE7ND7EOeWOoDrOB7gkKIbH
67NVUNfLvMDFuYkegGkOPXTIER+ByoRAVjErdIgNp+NJtmFFvclFh5VBXsaf0Scz
j3+mn/eMHd5v88eFoOjd9gSY6DTodYR1XquAu9QVKa4DFvw9MFUmNdKzr3qGfgUa
anDOkWNCOqSsqWU9W6b1odds2wiN9tyV2iIjaBhQxyTn+SXgzSSZlGmC8YfsOUzd
tWu0Rzu6wfmAV7yjX9xJP6kN+rdJxdBfeBHm8dqXRhLz1x9h3n7uThaqd/5Anega
mJTlSVU9Ph8sCMegtTt7u0mzM54oXbDAHnO5bVy3h9rAjUYKu/dZThW0WCKmvMR7
IaFaXWaz9AmHfcpZTVCupiE2hWjAi+gmwb7TQgpxQFP5xni5Yqva1B1tX46GB8mf
z8dbg6wdxpySUA6nqpmroeWXzfcXbXXoHh+WDzAjHxIBPMdM268XEGt5Ff8aXajY
cWq1fS/9Ii5DGN4Ic9laf0K9MDsHo97jIRisuYFnlReIi9TfCyh55kccbG+BobAs
iAvdUZK/fDbkaTVktF4bB/zA3/1YssLoRYSws58LqxA6+l0inejuD0fnVg3guL5x
IBARQyLXPrKjbxBz1qNU6QgZ7VzmYVfMInAxIGCzTlT+cIr+jID5cSoIHJvXl/6c
NEch8cCfEiaebRYwMjjhDhYZ0Ndh5/iVRHsgCW4lC9Th9CJ2AxLK2BRevOysv5lk
VK1fUpzFNOorpbjc0hzt9cxQ3aztWWhBYbYvxbW9eCL2ayDhhLaj5VWviuJE+ie1
wxBYmptdFaeRUvLTl4H4UXDfGgAr7oMPdyFP1DeCYgncIBgDdeztSQVuY1Mdu44T
Z9cqRulc0b362mqr57hgQgwIm6IbAmVVMEeaW8TwaWTdCbCRcsUHMAnPHKjeXdNc
CYGN4mWwkNWmVqBqkdx8shGHB9WE4P2yNyFCzY91RZ3fU0GzS703jpLhD+heq+wl
Mo+XM3zdA93BXkYNz1pKZ4ajY6heVnp/GXSnxuB5y0lgy5ti2RGeKux+HEiMmhA9
2vKI7FXJOZOfbKBNlNgCUtipRkLh4JExAjUOSV05/BVFMQ8yMToii3ZLBeCif4zt
E+hyBmK0SdCr9lV69bq4Gg5+AxATA26jr/5LRA2B8kzEw3OC7theO0Orv0GNKc5w
e7N14NsYlV0QRRyZC9SX8NC7P/fahrFG0NEtyXHU3uNgekGCMsbZZZ6mEcUhLEHp
JFTDEEk7v8S+pwOq9Pl7HU1HLEDRjt9vtZaGZQ9ynaqBjaMxD1M8z+A+p1zDuVu3
KzZ7daDZkX2tWjVXCbIrVfALq67+1ibqbtxz2F6hiAKMGrZPDSJGjc+R32D/sh7q
KSPxUKLzDy+7om2xzb3ws4RLMkY0x6Qo1Si+Yt/sK0yqKisRryGgTpOXRB5Ptjoz
oWcfA0YM7yAkpC7779WxjKsGjoMJ1MELkSxlYtpbHCRvXHIgiPMIS7jDfkp9xD47
e5gYeHV5c2bTf/tDAgc71DBG2VlCk8ReuEj4s2s8WamLe2OrvFAGNxsdqZF9OwpU
wlgi7+V0mk+mHf0+M0cCZ/6+Gtx/12juWQNTQg8ChsDj3uRS62ln5tNWbmIQCSTa
fOnWt3fWg32BwQWGs80gm1kj/KfSzJ9l6FoK4By/3HbG6tRuccCHlL2x9w58pg90
v0zCl51tNU4x0g5FkP1MlHCsxpYDmEJNKWR8SCXN+9jJPPHrk3ojh9wEpv4NxkKG
V1yhLL4O1GjPVAdoXfmoJPvnGXRn0QIYI7YdwMaukTfnHx/7JbNxyhpQSbZxZQr3
BFqIccbZn9YLG60bBIioBkxOu+jM2ymfgnhBzV08ln3hXY4I47Kxu2NP6BYLrBZ6
nmqGUpEKFjzhq9Q1JBiJ2qUCybB/i7w8plLaA3P5q7XK0d8Rcp5aztgQQQAgm9nD
4HQ5i/SwHFqKFRx4D2m2qwjgBL+RsspcjlKDxXcwo/kZ3r2SZpSEOiDeRVoMfuO2
kAC0zZCS3HnZBZI2c5l6Dr/gFqw+vP7tedvnx7DrgNv3HDQ84gehRlM7Le2oEZyP
qH31TCZrh5WqxlGlHQiD0YeQSlrrGOMOfKmxuBjkPh/ImoSJIkoShbB5mjn8ewbO
QHW9hmsBy2OJ9b7e5d/9NSxpSrGav8V2Z4EK6BY2KjuNO3JDLJRqHk53YhPYtmfY
MNeSmOunN3BJi7saOb9Sut4n3Oa2Y2bfRokCwT17UHWJI96WsNQw+UwANRnI0Fu6
4vajh7qlAA3fdLlp3A0soUWdjVflAuijksH/2qcibqakCW8/q15MgSWCnLFzIFnL
ogRaVqg+qAINHHZtp5GGscUo0B/KospYud1RZ4WhvleEahaVKJ6iAzvnnJYOGgQD
5XM28Jcm2blG4KVwG/qTwpTjhq2BSFVHi0pDGQjM+rm/j7FHxUD5hYVcEGC2bpnY
hGONNDW79PMuVDeWInT51tmHjSCiL+Zhq0mfPZwuf1H9G49fZttSaut+7Wm+Z9j9
jgEUOHPjnCooNy3Yh2f7kSHlWjfYgKuM1eYBI/vyfufGfcFapiwAR/vI8GmouATx
5Mx35mR+2hY6Oo7a2a6am/URlr0sHootExIZofidnaLXS3P9YQ2fkYttE6xrIKfQ
awnNFFpqqp5wQUKfIewaEro629uxSnWyOKC69l8tCB6OXfGIchh4VvgbxC4Mv/vz
sGk/kL/3VKcenOTAFfbCtXdLFbMpQH53kaJcDHJJtcu5XIz74JNq2bSef3onefzN
c93qqwnTMlHffrWOVubrlYu3OImQ8FOxG4HVBIYOXg8GEQpXtnf+0mkpBpH3D64l
7HekgiHgds5wZ8SvRJ4rABBa0v8FK8p7Xmu8B1XdxOOu9tMFliVx6ChRfZvm90wX
3KW5uqS/t2hsWbl2N5l9Mk995qiaKlCIePrG8MNUNvvI+BMmJgRpl4oc5yQTUSwk
X/6DkeTxH2lop50Eli7u16rzMBNXSmGZ/ayi2XlFIk8XLp4JqY6tVmixG9SFnzzF
dMI5IS1ltGvb2GYcCIm/+p2aeDm+K1ePngyWPl3Pd7ZiWGCj8XNnsLzCV1lW9DA1
NI6UJvhO2WRI0J6JrqQoWxmhyenoLhsSkEAAwdPs2ssmZzCtOyuT0bGKMhxSDlGk
Wd8+K+YU2VUKba760A0Lx0YzvU3i4YtOkBfOenTeLV2bYYiNrv+QK5Pg+ArQtNRY
hzWjedTEGdCwgVUMYlWM64tEG+ipU9cIDfAo1Liox2yyl9ugdMMRiPTnpe5tFj50
9z+6NUB6oB0fU1DdaqL/5/1Q9uTXRYYXEEeOBlASeJXM7LQZI+It1JzHGd3MkoWI
OliBvrvYeWuXlk6p94676ABd5nPbZyrIKfENodHBiJ2lJlOA6sMQXws4pu6OqmlD
QpLFMN12zAgBgbHKcSA00MFmboJt/sIWL5LmMhOGSwM9nEhU/cagC9LgrBTMf4Ah
DVW/J8GdoQtgZ37rTKVhdRyNs1koBK9Lo0135FT36ZolZGrduAvLFsRT6BqMPYEW
C0osQHdS27bL22mc2vtRUUuzHJ9kAoJG0d+EB80zqWgQKpwzc9yrETEQCJLpcr+3
LCXLFDm/CRXGkSuy+U7UCutrLQ5oFNj4owHtk2Ehxar7WzW4pabVgXUylCFZ1WOw
Vu+guwzaichsHIPQwPyuiYFDcDXx2Xh+rfPj0diGZraVAgLr1OgGM9OAsa60qWP3
aosrsXWwE0NfD3CyqzwsbGTsE9aoAzRtDYq7+H3tDVZicMpqKKkU+Kgl9OF25lgR
zb7JnlT8KxXG4aRq1ucug4GOD3jWyFbr4fyks3ONekD5SCXlvbpE+rCnxLCcFjAM
6QnJ+k0x7Cmm098HEc34FbAHawMVvbFiqwsprnWfzBlfKcw5PxHs4a7u/B3eCluA
IJHxwmkN031v1u2b55EnxnCsf0rBMBn9mkt8A+tBMdeiYHnyPFhC6wZcPMIP7u1e
pNSUZ1gDBEUKc2h+kKUfPM4nnuceYgoBwF5VdxMMu9vDgGHJo0J+IH5vs2nKs587
KltrJkKclQJLzQb8dy+jO8sRgLSMQoTNmxvBcNtYiEm4qRutNOt02sQJJbgvFov3
bD8SqWg4DDHo/bjZAKSar1c7b+eg0mbWIZChBHTAT5asL+c7qnK6kZo0T3m7JJdJ
EUYjtgcRWKFMRDvCFKem67pIvXauhv4bMmOSYjWRedg58OTryNebVOUjNGdeulcM
NU3PJwM7EKdRH6cpPhs9+S8pXdJ3Bxr/bGb9Ud3/ACIbgbjhN8ERK+KT5tnNz6tm
IU2tGNR/sxgTX2pn2wEGMHdAGnjLChK5MMPrhXxfBXHWQlABNriH8nQ29+kykcWk
/XQYWKMKSahfHXtmqzX7VtKpggefnGQ+REUQEufts3u9M5BpFtzN++H4L34bG7Kl
9ZRcHZPJ7wQQ2fmXHzuzK60z9yE3AEIDfr9KxN9YnHKdAlAJ7P9+JJ/ojinalqi2
S6udOup50RZcm348yVRv1W0EZ2vM2hroW2tlwTE5kGlJUVl2DpGqbSC6tzp+xKSe
nfz/lmFBiL01MZz/YzXkDjO2EJXw7mWeCl7hJW2NYoiF8IeHEnwwvyldJrTDE7Dh
CDMFlWAbHJipZvYid1r4ry781AZukVM4A44rVDrNZKxA5vM94aPqGj6PotQdAPt+
AedYIjBPFmXqDHntQmCxnZhLHtJSLr+V5lsAfoG3zLZPzCs0JSH1zQshoBhwxC68
E2H9EyOFPqgaW2bii3MvunwAMmkTzUBU666P6GDMdXyO8lBwufmBf2Ms1McsRcvh
bgvcVo9B1Dy+Yx2zpaIt0H9NBuixuW5qoYVTn/L3roa95pT4MD5+Tls5PzFtt/tq
2N9WuGF6dq5p6OO0wNf/67aW3T7SYXBgr8RlZ8SUvHiXbtouKMLSeKZVFtBtuGh2
Mzqrq3Opm0TfVUQCEERPTHFLhAXB4fiQo6/Y/hE2PD4GL9NjU01xWtTBBLYfh2ip
9kfj4hfLYTozFqx2N0wrRuOVCneaOlgu4H9MNgH+ey1/HNflTr4iS0h3gffVGe+k
MVLvOMJ8XPqCjmdAsj8FkI0t5vB6JXFPlXXC16p6BNNoXPJ9/j3gGB9MZMzmPJ1Y
VhI7r1NwdezeSF1QPptCuqbp7fLl5kiEoEHglv8RfzeU4HEjUZLtQdwQpnbowhVv
VQJA3aN4sKhVqJaxl3l2QyLtiJ5CMGQ0yF2P0ZG6CNAE3h7dZgMZ2lsmtO6OKHGn
s7uDE3tBJNKJNxK3LntvoMRxlvlMvX+0twZ+n3ecKt4MHn4g8UA5mlk6u8tRwRqa
Ur3pxPexkDmWYa9w173+F/fNqsTALFODyK1XMNJkfV+ojkLcwHeHu34IQqsjfR44
CHyrvyfMjfLqvfebydHncuWIIqQR/jVCPhCHo+NQghekV/E7zQ708hot+E4CqsA9
2jcnPDMTdMZ/wDv55Wh5L39eQPYXkkFJUluZN969soxhl5sF5/t6H6+6gBlCKLpX
pqqLC6PUAeSV5vJaHc3QOxIRhm79yGytrQ3EuYMTcG/eSO0OexRKUmu6Ue5fRkRc
Wlpr1zHZuVl26EWQhdbVVvzsiXXjjXhyeTUd/3HHYwi8LRFHRROfWd+007Pvyu6/
9GKiv9lELB7lVbd6BQIkujFxOKM9gUSQsuvJW3fZ8M0n4dNgnTtpmfdO98z19DRp
VjfO8cfY7D1tIXYxcRvUl5ToWAS+hUDntxgFXHh3dyWrq3aPTpP2B3jeSjo3DCp/
KUZ8aZdiK9GY4TxPakdzGM5pdEr6V2xeuuBnS8m6eTXnLDR3aBxThuVXprOiyT4/
cUmYh9/HtEg4Efpt7h+MfopobdzPZCx98Y2jYmMnrKg8dznsMv9ogSw0m6qFuOEK
kRrCw5a1/GO4EX+F96ep+Y0ybsrS+aN+5qpo3KMFWWvHu90iu9hfJkEhAFDQQ90G
kI8DD9U3GWZ++x+Mx1sGgb5zzWAZTeKvnwZZr6P/3cwTevmH44U3RuuNl7n7Fq03
8ezWOAvu2WlnDU3O9Z0UFgf3pv/bqL59qg3MKy2onPfUQl3BirwenFBuq75f9GKd
I0SvxQEbZ5Ul6hzlDSndyOCktEq6wKaTFFcMCaLBERhBB91PTOS/8wIYnvWVp5T3
LUB0eIl+QZRQtPmaft6LQQmpKErNEn34qLvLN7uCynZt/JcIiIxbBKhj6ky5N6G/
ZV3gLIo4DuAHfnpse/WwxEMZwnL4DJ5IoXUwbjDFfdAkIs+mvJNEsjP2NUEQ0vdX
/LSG4KQqImx9ZrhrC5QKvr4fHDgXnVXtsdG2fy5iArhSk9cD/NmiUhRtL2MqrSNc
+jfnx/2hnZdYPNVkFAf60g+sse4L5fYdh455w60XSe/sPfNDrn5l8VV36hYb/g3+
U1gWT8rNtziMS5dLmOxKxZl+gSwR1WdHpGmNJhROUXmxhyTwvSvYL9JtvME49qqg
xS+JJ5VQCu5fHWWv9972yB4bsSyQhP4ZwR+KbcJXDskG41cWKGQw62ACd8X4Q6Oq
tPlXgHk6AmV7vsy7SqqhnNlmE9w789jaE409tJ9Zy8FdWYSP6cY3MrhdaDJZuuGi
jtLItEj0obb/T+eRMUUTRE7OibzdwJoHe2OMBXeUq+WGWwuPQfSUHerAX1AZ0DUP
yAtq6qjPa/Ytpdj6xQ/QxTPsrRMLj0RmDQF1r/EZsZULowufR1NMHkAZpmen7jeG
XRhT3nTDmohd8iRRcxMef4QkPiH/N5Bpsaxs+2J8A+gimBW2hyyF78DZpik/ioei
ai2j0QnvbDLZYJ7cUqVHvugJcO6998HLkLlXpnuRZP1K5FHmTnem16yASHUlvkgj
TOS8o8Oh1+hvfZdcvyeMmxnFPpW+k4rECmE2I1LQjwjdlnZ3vzz63WG/dP0FWlJt
m/sH5kbXrSeBbaNNNzuA2IC/JFhZqEtknhW1ygWa4BQJudD5AB6ZBVegXbMAId3E
JqYQd3dNrOQmL43z8SPTVnzg84SObG9HsZiaLtMqDmpv2k+xvgWZ60gSvL5EShPk
HsqMsGJEAn4dueZZgHMRB7apV0mLL/OUMc4T31CFD/qnRtmiLfRq7m92me+PalWf
y7ybx0AT4rHI8HBPNbSORGVJr6ZwduLF7D6MVD28uf+jrBvxqKru3W3SQiHFhkDC
1JRcm/uMEKyImmnR8kFQoyuaS8WYMCBNNvHdJNwlLX0WS11p0oBq5mFyYw2u08ad
Ic5dVwLL6JIBqmeS9G1TV2SKR6v4kc7wEDnD9Qh2PyeicKtW9ypReQXpnlqH32ha
lJYx4dAWpsnKNltRt+2aCWIrgtJy9oMSxze4IreAcMeFgRjIxZmcd5twmgooMjbf
6ldkL57WuW/Nnver1SexNE0st0TfRX/nH37aVNLQyfjc/lyBgaKnMlTpnKZixPn8
iu4HHWO6fppRqsudEoJsUulivrEBaC+8jP9/a4+hRfCoa/E2AGGPMtgAK8fAwwKg
NQ2jpvdiD6FH/zNAMV+cCR8oyyTKuq0MEuxSaEYgTAEDDK5kJtQgbFGXYucxSG53
2vRSFs4TSydaNBpEqnAERkxse+C/sEvish8T5ugbW824w888dktxNBfcyP8wRGVI
C+jB5PLABoXLagbc8OWTmaXTHwkUSBtioBZhuDyCfPldgkCiVh/fn7qh8b3Q7hYx
maFxYZHGdO9ArScZj+QflPRMWSzGV9E3fsf3EeuROGCaoTyNRSNE+/Mej9Nb2Bxb
gY5mxW77UFy7tvaxD3VMZaAfmaxyES2gG5r0MkkRUO/5eiy7kE7w/jaSSlmiwBDH
EGl0F1BS8GzLMTAXpp0mnJ4eXwefqFwP4uwv6UU5uijyzdOEKg/z6oRqkkcAffLz
6xzL1CnJUo0EqjKbN7bgMML9dGBD5MDFgxjyQIAGHRm1zfxn5gSUDjwAdCF4QKav
rKGEWkz0HAwlmupPxnsvNfBWvNcLbpZSDznmssbDiB6kdG+AlmTgx4f6Np6/1KhR
ZXrunndu0OObxzBOQQ6yYST9/dbb3H8P9zLQ3uigzHTKXm0VHJcidqO8s5vytPzA
QTPhbKenm9uvibyZWkTtTN/z5vZvNqO0D8WBimUTShl4zD/XmrnQeSA9TZZ1/3OJ
vBnUybtTKqvuiowZ7mPsATfgyICyerYClqOCBefwXdwB7MJ1kcYf4USkJgmF2YGS
7OBdA0MJySctBdyIGwB2R22oDfOp1iWIX6ZJ2+Iwv5IzV77nEl3sypRIi6ENSvPQ
bjp50t0p7etIk2kgSKVSx5feZh2kFdAf+gBnA5rTN/lboSEp1XBTewJ7Sy9SbFZi
1e9l0/tbcfI2gTHPuTvAUPnpDuUq3Vzxq4oIeI/o7ZwGUmMJrr4KVPKE8TKP8hy3
7BTlYp8/mrIsrQXWsFX4gtkFT9e9lsdcVA5Kyi/hXEv4qA+6woupoz6jlR0FlOPI
DmE4pd3GiR6mHZSMy5xJVQjgqmlFFqW5i/aPk4fZQ9DsRLEXDDePMDTSqUS+ZmBw
obmsZzKaLBP1n4WZTr8nYe6mhekVMj5lT7AYvdNu1oXA2w9u8dMSBh8dQWzQNBWn
frJjlpY7lYAuGvgkYklJO3UdLj5qs5EmpzK5GHoyfHY38ji/eghQ2EAN0+88FQJg
hjUtHMcws/LSzu0TA0sMgI9RQtJUga41cBXJWLXGbCJyDeuVeMD4qF+w/2FJGX4U
KRXZa8aaPx0OKarVyo2Zrkg59te+90UxpZvoZ0BrR0aiRqdXDkVnvbHUzsxvwGsM
h1V1mxKszGqRKTLSs+a8N/Ct4ab82FT+gPxfTmrSC5qNhZff0wAsKULHnZ3m4SW1
v3qmzqLlGu8ECZpnBxyqmYM2HRWETcWIGHuzHqBP350L5EMRYqI0p+bbD7AbXvQV
PSsfADaannmL9t63BeipWdJD4r1AkO6U3Wtlm8Ya3EQKtv2e7lnTVbGW+3gmqq6P
6t5J4mwFyfRfGlS2y8SKzBQfXr1bMNO4n899rROZRBvwCyxT/2YCquKoesZs7Qs7
JgykInB2cJ+r2rKhhZr583JpRNS7zYmp55+9jJ5z1x+hyoxLGkUXVgvdvbPA1Qzt
3lfpgXPEOqeb0albCjjdAYXUhAuL2gijxzXfPsG5JG0rYwHE6iLauf1D6/FuMbcL
xEHv0wndnil8LrISRdk5kY0Bb6WRryN/DWVy7EaXM/le7sNADrFfwqIcnulMhOXt
pFoN8wLv3Zy+QMhL3d+YImPChiQcPMK/1gPHmAHRmpVhz9sc01oHlSkXvT6QOCzS
tLxK5pfl1c24NP3vigRbj9r9YYSnmdrWwMMywCCmUj5UyLUdwkvAz2sLcjW+7bnU
uN2k5n8sbRk/MS/Dypv56dTfxKJDDXrbvU95ZjQD14W82ErbZ0W2PQMsR97kITxg
mtx1kHan4CcCD4nK/b4w/30a6znq0zTvcxhh92+Cf+LD/CnEiKJvgA5xY41eRoUd
tORyGAYvw91+ZiGTRWZrhsNv5UQB/wmXFu8VL0eL8S1yGXh13F/D84WfZh3P9XQD
t34H6YhVq6aOJB0cHt84dW5vbGjz2Cu2P14m951dH+PPd8hm+oUHjm8lVpqRCCiN
d8X3Jv9hq1piGbLhKTkQ1bK54sjOQlSoy4TaSV/mrZO0bCkX2Pn8NovF5vFGArhh
bSaolaxXeLUo56idywAzroZLke3Fa2eco/onas805LbItP3XDF2Lc6UZEzBYw1EZ
ZcHgBEsCvlw2ufPTAqBlQvVj/HQj5HGDpZXdvuiC56jdCT95nu0OV9VwElhRh3v6
NEzhoS7jwQR1wdfEEZg2OX02352AulBX/3udOSHFhHs+NWOVPizaYOZjXoIv3+OI
Bdbi3Q13dKtZvmrtSeZWAhKULNG2zQJTk/ahRxJQVbI354cOrmEXNl8fSodj9SD3
m14sG+WbiWxSa/7GymnzoPrZ5PskoGjz/gNdJ9vdB4k38lXFMjKBOrnKR9BS/lDE
uUZc0NdeTnfgbJlP7mqYRkjH0zKsQ5W8YQOzkh4z852ug8m5Bb4USXyZMGZptKn/
Smze26Djo/BUIuumI+t8DExEvXKzf3vZjLIi6pQJF5qNOpL7Q7/kDeq/CcbqXYqx
Zg2TkW0L/EWvzjrS+R9v+0hjBFMF7654CaY2utz3AnmnRGMimXjLVxwsFaYKkoyD
OxsLeFDc2ybzXk9BQO5pThyiYoJ7NYoSZKswKRl0ALeFqyh/L9kgj2aLDKpdjOcU
waHyetmSaJDIysU7pi1JH5NYTpm3rLDqF5iTrH4cW7QKEN95oNZmGiWisBc+RNRv
5Dr8peBCDCiAzGsrjifWv9KqnbK+n9M4LG78rpHBwowqhwHJmWsIIfMhhoI84if1
SFos8116NtHjCm48OyAKDBokHfV4n80AK71sMtyGPIfM7rjpkMJ+A2C9wuznvdMu
x9pvz3X9dvlDzWzJkrTu7xmaU289STNabBFds9rqqeH5Q2nbhWKkcv2++3mZYHK2
47rjFsYYbCRFpVjmqcRM7LdHcJ+JSX1NbXpwurlXYp3E7ChczNuma7GuMFIEqswi
VBrWeWzIFsQSo8zjZ/z2B6FVkpGXaAAHlm8FcJDT+MmJJ97IltJnLFCd3QUX2Qn3
VIVA+dbZQR8oKg0Lfy7Mmdvup+lno5xShFMEXoZWrPq6cTWTU/sG88cyWuToX8A4
V7y+uRBimjRoUGHrAKARCcSOQf76Q7waX26F/5GSxNBJg02t2RnQvuyJf2x7l9FC
I1UYtBkKRq2cYPbPUJ/4pQka8N2AcXKpM41yc/JYkbGFoqcsR65Yeuf0hL8Aiudu
DSHyhYfx2jTAlrmrJhonK4WYaZUsq9XyGUCMgkEBA7e0snibzeiZePxbGKSpErdN
qiPdFXYrrr7WQn7gdFE3s5nU9hrbxZZvzDZJ7+AkmS+4L4f/NltW9EEp2MvfB7OT
XoU8p1t0V7aq87A9kDPc4twq5J4jJI19SHZL88Gh6gXqZQQRPEloEQaJntFBnoF/
Y4UP2ltA9M3UvANAt2idB6W3WxYUjNqV6HoD6lOZJsfj1kQqT4n5RtpqKUutXJdl
vNHGrCC4gphLKh7qp0k5a3mQV8Bm0LrZdPCbYJ/BxTfoqT0Cd8GUq4Oo6TrJUfMU
FGf4POGFvv34U2/3xgVQ6X1g8uedCrWKW1FlxqotSBHfm7nHVyYJHaBY9O5pGoPw
XfLiyo6ON/+cgbl0WEoIqoAmQgvuCvJudbXb2lDIxvEkAA0UjloZ8d5qDOo2Z8UL
SW3a6dQK8EEsCFeBqv7i14SJMjCidYr2k/IsX7sVckct/vOXhhoQSxwsfCINh9Qa
Ajd5i4dcH3LHdRS0zFDpWAxXgGiXJQumJnsCO0tF7olzoWbcJijAo0aENRfCoYHC
2aEFx46NsLrDr7S/BaJYxQ2vtOtRd+y9up4QQUYHlARYfssie5DBAk3oMauu8yvd
25WSdzzwRB2ZrYKvtwRxzHdzMtzRfI/K5XMd4VXUR8SURqvDRvABvh8XF5WVNizY
1Y/swCLz+8sBkv480IEL9KLJE3VPPQV59o2UjD6ne8yU4Pn8C/PAVnBPU0jA3Xyx
ZPWA4XVFyrMxiQSf9LURTZfBimFKKkw2NydD8eCsfu98KtQe4CIOim1eEHXBA23H
AtNmykefph91PCFzviiYYk5CqpABioOF+PXetX50E8sAyKW66WYcG3t4wm+IeAwl
40++iu5MAssFFSOYqpIeeIaEOPmRJWbeFWY/8L04vRzZ9/chbAQ0BWiWnYgqeslc
u3FlF1Fm17WjkBXK25km5+/e0Q/dCbCe7C6knnKzqrLuUKRGHFOYEMMOIkphYx2y
z7vTGB2989YIiDCiY+QN7cvd5Yry1oj9Vb5uxrCJ58lW/PQhnb/fZJzmcxL8qr6u
nxLXqWts2xqs0gSPD3dQXmlzVRJST0+tovfStncqj0SxX8/pmVTztaciXSTcMFnC
JLxl2ZTxoxqppDOBRxfMYZWUP1pxgVlXWjK8an3p+KEuMY9cKMkqD78vbCpC2Y3s
T7/Gqe6dT0NaZHJgX6HohIbFhTWnlapjLk9gnzCcq/Iv8rPnQ2G3D1tzdG4x+7tt
89smJzy0p30kUNN90kQJZPnyZ3BSYm0eR7ffiW5o8XBix14z1ZbvHrv8XWLnTAlu
PALaFe2B84iRSE859dWjCvFQ0X9yOY6gbE3+3N32b9A436GX/DWQ97dSQzd+YIWL
cK+nB72QFQnFXk1PCNZ77yp3Hp9qDC4HitTGZ1tVmmCFiX/mLSLC7vtcBd1ipT6i
kNEZ+BIJT+eQJl9tROZD64/BXNzLjL6rqvqkEe4JmlKoboYG8i4EGu+2R0wVnHu+
OdVmG39yoJmOSJBEjuu19iezH9Ss5umV9y1Rx6gqVjzz/Gxlr5W7iXroaeVJf+M1
mOH/WZcTCcoLbOiVwmoWXPpF+3OwS236KdTIwZ5h4tlEF0uwMoUn4qkpH93qr4gJ
DGTtcVZ5KbtACpBPh8XtSQ9yB7wHw7TcqZ8EVDm/p+R7Y7QK2BNSq6qEIjMkt3S9
K3Vifa2YjkaZeteLq0Tb4ihiD4r4jZGBymnSTtH2p9Oy3Uy3iAbIe0WcpRFbxwIm
QIooRKJ91HGkVnek/oHisyhobtQ8tliUDCAkCWDfCjIuix4TQSl0z4NCQqEL8mPu
aie0VZyPyCjpxatycmGCydMWybWkB7fsTfoetS8S1mptTAHSVrTED0cCoDnJz1nN
xuXjBibB48vSddBOKEsZIJMvNgEWmPRfgIuBoB50yhriFXVfxOjnPNlKIAjYaVIO
FmNH9EuGETb3KYpbtN9meFVjWi7Jwn1u3b7wKAITlfmPzVmMOuAvIwPvO5vVngP+
b/bCsSaxcJAvOOasaXPUKZWUO9NdgrVhYttdb4aUzJsCPA9RfrXofGF2rjPV/vWj
y3s/NIKVWVA7Na/2N2PT2HY600k0Oer6YNF/WK4n+e7Y+UQ/gKqOCdLlEZO/Gcee
j6rUZTCNiGHJGbSMgxOydmZZJoLQ0420CbeVUs1dClf9LXqjGONW8danWMy3oKV0
tRGNLIM/JkD5mWsVy64U+T1rSrRuxSDQHJIsXx6kukOOrEofwgHqZeWbcBsPF4w1
D0/yRzsLYWZ/8Ct67cWnyokw68PDhxldVwnHzDioimj4Dy4ZJcVIYgIlRKFcR5Aq
zBXy8WZCZPOKZppSakK4JcQVvgdwt0qOnDCMXw6xmIoF3fFMxMozBfpmPfTtc0pz
K6NdMq9ZE5KpPMtaFhV7Fw8TUrvp5kQxKUV6kAIvNTHlhfaw2oQUBNg+c6MKjZ0L
fvosGLJfDPf63TKU/RzM/a9iyX/D8XufEViEoTdwxyWEC+N5UD36uvCQ1jVn+9FD
3/fSyfv9rDNM7JRuT5jYuhdgu/5WA5ceiqykJlnKw30P0JWHJrltBOUAOk83KDYL
JXI3JTaD+sCChsejG/NIJQYKb2HwhLkn8aVzJHYFEjWQvksk0a8hlru1cnslaThN
flhELt81osEwvQXoPUb/lxVY2lVMPkxhVykCaxqqC8l606B0l8sOJ27L7+BX1uba
XnVOITrbZHWHSSkvnYKZz/LFzqY5hO58s1bcGqx/rnZhOZjaMSmX1FAOqSE4WB42
ydLEVb6CdZB/6RXdtoULn3YDPYaabuE4LzZ/6pWOm0ntz/2EvlwO/w5iMsJoaP4l
juCZt4kGdhx1sC8xuy40+nQzAVYURSacManQ2HcCocG7ys8RMu6F2kJl2U8QKTU3
qDM+NPKcWfzDlLgYjqk8zk/nfmKnNLERNjOK3ahf2VheRCZh/6rxXm157oR5fO//
aBTUIRG5O0VfD4PGzCtAD2EfhG+d0bd1zEGolpYHABxj4uxjhbGWQfHQJcopUdGE
7+/j+tankewLlLWbYOV+Zh41NKPdlTkNnD1GT999VFoFLgg3SGPNoQmDX4zsCQN3
SZakZjUvqBJjabq+i4taqlQeMIw7sDdnXM0sa4e5AjeErZd24E6NdW5CTgdD2el5
ddE58PIKt90+CnzSggLuMGFc5ZZZYqQdVP/IxbUzc5tpj/pwICD15qL/khMVV33U
GKa3N23EJqjsVaf2XIblt8kQcZJpAf74PCscnI3un2DCKDiaho33hiZOfbm+7PiW
xR8Ui8yu8oC58lsLPivasY6ARlXGW2TZCP61V/TTaX4IIGQvVKmq/kC/WOYKZNfC
gDl5FEhU3Q2zlLSYQf/F0iCDn4SzMdV7zstVfpFnPeJGOuAezfj7lp3V7zqTyW6b
ZUwGX1RHM5H5ewv3iNQnww5pUS1JhWoIx+Xi/jA0kMKuey6+TmnRi+pLffEwE7k+
GdXM9JRNpNG+tdH/p6yYszVf1rUsivSbikDqZI9el0O/KISN/RRzfbfNxUuIH//d
5o765jmHYHsCZWjg+F9OjOuNnh0AZjndR/dNRW+jlpM8wwmXjWzYBVAIu/An8Aa3
0BsxgzxCZDnk48oZISl5jNLeiKR44F6aUz8jaCzPyDtPA+PGR4DOZZeh6TrrBL4U
EAVbTB/Wmw0RW+dcsFMVT9CTMkOv3XRWWk65H/CwpdeZt9CYOlKXqBBH66C5Cvte
OzPU/nM/gMMu/27BhgnznroonPqnBuvKDKz7htgoIrqF07wTBG95kmMjFfdwJ9LP
OQh/vKLc/HTuK+MXL9Q9vvxCUjsuqz4AGwMHWWvqTaueRXJah86z7DmdiDWgE4IO
h1Z56IuUkPGbXYLf9+X4Kuvmp8zVA/y73vxpkDm3hf3p3Pvw3rksMBqYHxdDb++g
iA0Unwzw7ppHk2nlhJSr2CEyrltg4YKCe5cc/AA/2JSaT9RtClO1xvsPwrb+z5j4
5PG5uCKT06dMMBCMLThtcZSHTcVTdQ6m8voIIgAxGElMMJf5C8rzCwd9+0Vd1WVK
lQCBm8LCpzylvDtxwlXZg4FM4GMaU8+ZZ4pHa6chishW1bHUeY9vZZQJkT5IOFRx
QN4+rChRrGnnHLKbEfsFn45c6UGH3jq5Hrfi12elUJ2ZFe5OUQB3IMdGywbC2ypS
pHQ6sTC4L/T61yCATCTh8jBi0YCTyEybEjKZJ7n37QuAzJl8Ms3H9F4yVGSnuJ0v
Mg7xmI5NNkgNGMp4NosFsXFNBYDivoHrypFJ6hH+MkFZoYZ5jsFd+PHy1YeiQlAg
iOPNXImp02xQ2mpv45ShjrkLRgw1qMZlA/c1z8dwNZjFGFUp4zzDi0Hy7dRgK4fe
TCSh0x7dAPd9tDWbVSCX2sFmwiHYIqISThvF3xCqeeX8hDhVFdEnIWqwHZg2a/VP
hSJWSCI95jixPd8K6RaNEBt22//f9GzJKJaUy5RB6JDDiJCG8L9ZsHaXrMd4OV69
Vt/pwozsCb/tUiP7VaPaYabXmsARQ2QZg2+4RPFQOhtSDRwQOungHvRTzXgKldQ1
MjcS1h7QeAHPQRSzLpJPZGg5YO5zgFnML5SQBS7ixfe0eDhbf0GKM5YKJaNYmgdd
NHZny3BvL1tzaBH27kW0EVhQQfid3XQkEmm3DkNNKcN172SjjK+cUAyzNIzNmSid
rDdyqgNXMLziKzDMKPc4fnIYsHeQ+woh50M2cdcTVbRpRy1qklkw03LPt5rtmEXK
VPii4+Z2BerTaXW/liUs5k2iKoZfFslUk96QfaPqbm3ijOfXx5tfEdpudEt9QiYq
T2yQYsqM/K2TSt2L+hbqd1WSqSg76TqhYuDN/U1BG0k2lvTsIrNNgCbaik+iCoeN
PkGXE+Mxp2Z9TupPS/QE0qrc4GnjBz0JM2JqFi5q2d0DiNBu6CMMhQtPCTjhWqPH
nYjohbPKMxF8UJcaHOEzijlfrOM4BkSi3P4gWAauXL8RFuY9fxckv8c/zlTb400R
XL020UX/Eh7jMcHpEJu957LC4SuhUGGdyEi/ZAuPCzTks94BrGx8xfoxHnwjtdr1
ggUw6yDKQqdeyVCQrqyN1FzbkN/i3kDhXOgBMVv8E7T64hz4TJqndEybAyJfKho/
bmhAS8SFAsiU3Nm7iLcBCpEhkAXxwanAHZrGJReHLzXdTmdW0BvaUYWnGLBSUMCJ
B0wE+hQUrTgDHFqNg/ay9/8YFW6g5RYTXk1nUn6axXZDzDN0frLyDHJLmINhKL5r
07ysMCuERFFIvQTOSbPzqJDnrDq5FoKmHFbnrbYjW2q3j+5QtTzsBtpypWo8kQky
ExaslktDA2vjAp3SLYTNseTSoXn40E65hUITn1uF007E0pN81f03WklYvYuZLK8W
eVaVMLGLixWuw1IumP2HREmRyDiG35Xa/DCyfeB/7wwDSiGH+x7aHYU3ERMRbVkg
ZWtzj7CGuzOQ+G9xdmhsTdr7NBvI0rYoM4KYmZdfinXar6IzIOjgaUwVeaOkp+cm
eVQnB+WDyyWfGGXVvIP/EfaubGt/voAAGLAuyk31c7h8GcBnHGwa00oxtBVnalKj
Nlzb2fSBGKlflgR1DIdpedQaxnNTBB5UVzc2t2LHgKNYu7+HH3pN+ViMtuENWh3j
Ix//Ej3rRkCaVkrvxQFKT5bq7ASnD3j4r3fvO17mKUC64/2lh6UVuAEcfryBTvc5
nJG7XxSfPeGQVXlRjOy9T+Urm2RpcDBKBwzg4w8bD7PnS8IsoNtOM7yZ2tMDbd4t
ihit0iw0frS7KjycyNsQTTgQGOgNu08GrmkWNMCOsjVO4IMHRQ6SVbk9h7oOKqLS
KRpj5MCgHuxfXYjIMFLnNvS1VIfrGX7brOS4Suf1icxTNY9gLYIlhnyo/z5ZflIb
1P/HweMDC7UDEvYt1qYYu2eGNjBkOyYrCpr+i/5eKlNcme3agKHFg/OyD1FtJoax
lKQf+A3km+RT89nZuxZsJg7gbIwLjeFHx3CngPXn4jtqz5ljUPJpWko17ufmFyst
tLR03Mk/7tGnQUtAo0Siu5d1RdHifFwafM3y0hK9uPqIfkDyPZe+Rp3wVS1+96aE
Xuy/47Gb2w2i/o7ICF2r5BFinlbXWU6X6fMuQLu4DQcuPOTidr0ziZJwssRA547e
tgjFiW5hS9mDLxcdsiLfQiKQlYWDq2RluHIt6/eTMW7/vsGppFtQCTYxvg5vOdbg
vZQ1FZOKbyj2k4TBauMQC0O3KZAEOwQEnzxDb6pTG7a4FgR3BRoxVliRuMGwUFod
80MNZvgivWVv+RWJt6DPP+6OWg7rvQ80ZxasGFcdQs2y/UbROXahPIucAvjng9ba
y5KWYdHd70wgoysME1X8jNvjSCuPTEV2V5ICp+Yhg0XhTB5AYUKsNByq4snfBXaL
POK6GY0dydL/AnvYbWw4Vbru30vNLBNnndWCvRLQRvSTS44O2ZYyjC0YkUGyXcbc
PaUo40odD+viyIF8dWddRyu8ZpnIL3V0HEYB0r5wYnPlxJLzzcCb7srsKtY7Bam4
hh/k7ZCFxZjC09/9o1jV+FH2KPwcgj/wDRAUTq3AlPKGg9DpqJAbJbtxU1sOp+mb
lOxIoP2wJXTgwbT+cNAs03hX73xKv48fq+GgCr/wEl65WKMN+aNh1+SD4x2ZEWWa
aANnDfGZXh2GdjbUhMdLSm/2bOyM5HI+kbMgfq59TRiyhRO8BAJVrIO6kodWvULf
g39lrCF8AlURnerEt4BD2pbSGHy8FuqMnO2+8kRYoNKUedJH5Bkz3GKJwW6b5Vnf
Xpk81Wmz9ms42v/VwaWDEaniHTEUS5sxt9hzmVt6D0w509kHqpndTLB3S29h6uEU
Z2wkLHVr0rz5Gq3518Z9dEMyil2gZfSJXQr4I0XyskIezTLSZOzPqEtkzzfhWpIx
ty/TosA5w6AwnvcFAN/XgYCkpxnMz5dshiHnoU53mFeywNgcH/EihcXRDfKbwjVd
C/vvZh3HWAQLS/ef1m7S8WEZ7iqEdfv/oIilMOv2TZRSM8AsF65RmhgyepgrfbE1
j9s1wQVfrFmOFTiPCfMdDix/0JxaT01SQhi6SqGnUxi9nt2Ps0iq1CJ33VHW7rjE
/KA4MRxo60AqIuN/VrbBITSz13SgaL1skN4FiFB0zNMZ/vtMrpBjT5xbQ5LmyaLp
89pBO1ytKvy00Gz3WDH8WsyYhO7eLtZ1Q2emDH/TMB7UC54t5CWmDly/vhoekMMJ
kdWIAvlRmVO7BRrLU9JmQ17dzIUFFsKdKRoCw11J8rfflS0HzNDa4ouLALjsBP9y
bAb2lktYm8K/BRvf6BWPU1lQDjue+U5C3kiqwK2xBQ1u30DTQ6c6GIaP3now34+8
2AaDOmu6jUwSG70z4xcnuiPlrjh/xpE5vvXjGzNh/AyhPTh9OWMvcYj+8KMJo29o
P+D/U9wOPuPup/VAGIQPlkKhErdxzvg57vrQ7PcxbYQV2lBKiBJ6CHvyg8pbDrgE
OvFHsoRsSHviuUys641xnk7sEfB1E/QI01M/75FD0Y5jDDjotiy+AVbQG3Grjkd9
/btIhOyTTcaV3ZBIMN9XEVHV4euQl6ZKzT+kmVW1CL9ZcBkmoqeljIM/LoTFZDGp
2LkFzLADuoPuPWEa+blXSl4tzDCir3P/j6OF4U9KlR5gBM3GB635pwcB3RzzBg9d
ZvUwTxl87JkhVxQstQLtkAC1CjndbFeKnKb6MqEEJVCiaZWRdFzGXbXY/tknGHg4
VI300YaGqDiLLfrAoPrmKQ6X7oiPEnpOVwqjFGcXeg4HHbmgvypWHqNnUoOzvGeN
1D6CT1N1+V1pCR+zYrPvTQZ+wrdNgN4kuiJIUoyPb0A696gjR6ImrbtKPiOsIZK0
Jhi+42EjCgPOCethadE8lEJR4+mrhQy4yMg/+oGpczX8uEc9XHq2XWQaJw0ysFwr
QF4fcYlMsFlz9BOAkv6KMeW+0sCHCFELe7iGN0DRZdMR5t4tUVjK6QfeV+jRK2d3
YmUxqvArE5K6rp/NadCr++y+cgk412Xw7mAHJ9Zwz2hi3Ex2PR8WfntOn+Qljq16
lj8edGqhtCpbMQEY0P81TjKwaQy9HheE75MTXyjfgxfq9INuwm95gYH3i/JaQKAE
E6oqGAEnE/j8/jJ8zVH/1ySYFusZuB0I25+Bqj6TrbIBUthg5Bxky96VDNCGujH4
xXEj7M+GVtAry67Zn7AeS6mM39pnlvwLlNenq6DiVk0AtA16McAByeXoyVdUk58j
NGb2ENYiIDG9tecnDvbGsGsGvFbDJq0ZKq2L+9hcb763xkt5xbrPIUVYQ8/i77Wk
dTUHIvwHxZio5pR08QYJyxHyftXbnYs/OT2ZLPFwZ+t+7M4ZeYj+JspKC7aazpPz
RuyIzbmb+Fu5/44dzEBCTDCqZuOpz+3A1PkDXuQMVXE0g1w7faZa6ObTpj7IOTGC
hvequv3wYgZpdpYXEei97wsdnfrf/lShoC7mP3lZ6BI1/u8KKTlFaftWJji+x9E4
dt9kxoNKgG9uW1CLDCE9NkE+RDpVK4G3S2Vz7RQRPTEVQ49SLc66pbHoldeE/1tQ
v3dletQOs3MyKY857iUXcqiKp328wKzh0mVFA60lMkmTodmnAz8aKvK23WPUAhA6
CU/CrdrLXHTRoxcUEeg4gKeH5CdCmVR28r9QWkiE5hrIMWgoOQUpHKhZVGCI4pVa
wTLTgQqlNMNP3TyiVAQgNw3QTsqgRQq8mMRzxssrJvMc6rEtJGIOijvUjWC1TOjl
jGx8B2U5Puof1Ewx47e1nkoRGzxJdRToP2vI6yrFHzNZnLN/lcbsulQCX5L1VfkM
uffwL64LICHAHR4OD74EX3X7OFww5UjBl0ogOr5nZ24Lau6ALIBiv6VnV45G4sLU
7a3ZakH8pY/gvUWyM3rbGPbb/hqwMQLn4SEGIAYToeaK/agA/YjVQRIh6BH6pluL
Xz7KoR0xk4FeqSomSrrfOq1kOXA7Muv5a+ZE7y3XV86zRvnccvl5ml0OcRVDhp/z
bEGPnmLUA+7YShB7ZaTGTdjSeM4cy7tMugmz0ew2KWKPCy5qFqHy+Yd+M2hZAqPv
JDKStjGP0GPtapXj2Dcgopwmxp1VMSyaMqVoWx6gM774sI/68TzH9Gf+Nd5dnd4v
L7VsHcpeKrZoxY+AxznArA95qIKSaNb0SE0FfGB7kpp/Tm5cYuz6XTXAyebINfSE
v/S9XlKRzJTlysv7rsylOHZe5nLoBh4UUardT3fJUXo3ErXwo+8t1z2ahUZasMHo
T588PL4r03V8GbYRd09fPytXCOVIYylt+XQgX5UsMxCTBmSG8QhO0n3HjWfU4P7X
6fp4GpTxl66dP+g95qadK6zXeoqYZ6Jjx2uBNcZJ8MGnMOxxI4sD5I6W0EOINxvU
5UkMVb1VtpmDEq6lbe7Jr+QciWM0BLPcUXnkZ9rZDRWcMQdnEUwJSdQOewbEBZQi
NbbSchuMpbbwyMz1wUzVYaCw+cYohwwBJGJNOqMkbHBTKO39PY8jLmfIiWqAo+pP
WKC4997ghhDriDlR9bhFILfikMmN2LH9ce/yRl29sRjesRv3y686/gNDtvWtdBw7
rboCEUt+BJAwDW64CY4NpDrnSb8wFQbiHCToiZt7zWtP9p8GJjDsUdG23MKxw+Ys
UxZz982HA4XF2Y8llTnpN3lEFjB37/leCNF5M/FlAS1r/LFxwHBz/ym/EMWCgXss
Py4l8z+9nXF1Q4md+eZOouMcIXqUG4/GKiC5PtnTQtfZ+Sb//BvrpXD+bCTntj4V
hjugDf6sDZinS5cYEp4jUgUXrO/favtCnxxXTUvzMkbZ68tDkiXaB5aLiAz1HOGn
RdLlLcxWyfbjBKWPxtdTogZ3XTKT/BNeRE9eXjx2OKGFO8PkrJzw7YqvcE6eUsZW
/H+Tj8shAeBH7/QogTsFjXckEdggAj6nrY/magMHyQZ57l3mIfE7GDLqf5ZVqq0k
v8IWtbKeNtOrbJeWM/WRKa382bBlM7wZgZHaeMSTUJl0+Izmul1dGDyXXVeKZJsQ
OScCnhW64ZtGpbZoPB+Zou9HH+sYI/UUa2FL5b8W6ZxkYrD/yxLPJCTAMBAUjdqX
8fJI+OqAa16fun6HEWkJM536WQ8aVYdKuco3Rhjsz/4E7+DfTpYxdaCrSl6bD8Wv
j2ohfXtuubMEF4ZQfagfEeEzxJvgAFZg788YFIk18KBJ5JW4dr/10uvfIpT2v/YE
hb1XEsP3VoEOyucgtBzeQQMfbF9n+xg7hfL6LTfy0MnddAfnqv6DneBYavB+R0XO
nMv3B+yrmirHW0dP4lL/A3rgxSFXcO7257nw4ssFkMjnhcy+1OOt0zmORES250rV
GUSmhCcqkIw0calrQrrnBmLtfmE/B/USrDki6CKBu6K9B3wWFemswPHk1XD4BNFS
Q4P5SjY/s/L/tH1llaK7kRVZWJoLru5l1Z7XiJo+ORbkNB9G/ULomjbh4zPwQi0t
i+z8+p2EcV9btjWUqQe3FvHQ2edj4EzqA/McChnCLdllAFAfrcygrhRETzVJF1/K
OnsIRt5T4dsKQtiqNk4wkpfPHl/HgpNq0kewNLMU7PoDN6XxCVWWGp0pym9lOj6j
dVicJROJCgkMzTnJGarsweTFtVtUAxUWAzru+TicyJ8Mh6qgAgSsrvb/BnHfsI7x
dD3B4Rfu8y56pfInoZcPB8n4t7fiAwqMY3FS3dn0TBllRKPR2TGVWqIusRs2h8NL
XOQuu+yl7hPnHPJbRgdjx3226gyEWFodLJCHU6RIxACRc+CzEHB5ONs1zHCXCA4+
wI52/In3zXTJtTFqy/+Urord+etEoZ0EtttzO7vak/DZ0PZ5kCFT1aJaeTjwfEHC
Ro/93EpQZ8d04t6ZuDBF4xH1mqPOSvGn495zqC2kOIP/DK6dDu5hTB+sCifbhAL5
R2TpnYZKEd0ZJ0WSLqU/UVx/IfdU/q+y+TYXR3lWpzxRSzVzTe3NbWfUuzWNhqVJ
7Ecj5LGNY43fkOvMQlLv1rcfUYDVMU/sk61HFsCH9YXNciumUGWuOkd2vX+cBUsd
ehAwYQeBmXzLvgxfYtiA/haP3oM3DQdUsj9i/2FPgUOb+h9TenAYyzxXaErUHjCW
Ui+tHk9XRuvMyGfXlymP+TbxAqMVhLOERdzH0ogu8ppg5aVxNyQqvK0tfGgxFiip
37762JqaFVv/VqoLZjU0j6gGrX9le3Pdane3Y/I9coKsVb61uJai6Oj9qq5O/wDn
2C/x02eQhQME+oOMX7lO0o/aeD4orzxGsRxkvmIfTjZny1f5HHuSKfkCbPya8ids
carbMJTWjVNKMAQhk5dJSaNymdWLIoqxJKKgyJ86IHtmmaRjigmmqSgb5n3AMe9O
sMbqKmQCbrySWnbUP9Uw2FtCynR0vLu7cFfNLPBKUrT4DKwqfzvXWvAZQ+J7tviR
uAxP4uKNRWFOZvSI6T8wVC9vYrf9AmwV3t/m02uhhh96Qhu9H/rd7ZzXofhD6P4k
CfInBiEKRAlFfuXgytbfMl5DYodR/4ClR7o2KpexnMMDm65ItYlNjJeoKYJLUytZ
STUX1s3ZRcM4N48qrC2/4zZyaM5KcFLr0qeuydgHYPmuXCMM4gJrQE4IgfQfSycJ
nTFmrBsNICOzrF/QOrPHZctDQhJSkuiirIAjUlZ+OSx+mac9GtFhO3kdPabM1CXw
lngX5aUjWmBv4LkwoYfk7kT0WPZFNh1x9bZPvrtKTPDuhSVj1hnXMoW9aIEVqrvD
6U3p6CJrZetWiILVVjOhu/RK2bByQ1zgjQuFZgo3B44L5VsnF3wJqRdwg/d6njB7
D2OclajTJyfwxLrDRQeDddpq7Ec1yh0O4Eudphh/mdHVHTP3zmwsemyKjT30jwiZ
MgQY9lnUvvKm8ICbQPA2gbbZDw8D8xr6uSVHML5uBltKbLPbFddnCQ044/mKvX8x
xRg/THxMkCWdUj4eY5PUP0IKKVX7gGYLvFc9t/Qyrbu+Yf5gS2BkvmyTWzzkgC5W
PXa9sEIgFeLsSt2ORxS6GmjFueckJn2E/T1swB76lXI0k+1v6vU7eQauP/ohY/l4
IDY5OnGXX23PqcYFah8xFslPXC5h4IFRTl3F0kix6IVENNPoMG9LjZeaAZpTPINo
krm4vcpZxsYZ+QXb6AVph67JsSpP9NaScnqkbhfM3tPhWvRfDVmIDXkxVx+Vv6kT
cl1ucd7QioU95yRaNNc7fTiNELi6eiivYe7jqPoamx1AJsWI4gRsiDYsBlDmSJCr
AKfRbBFTquid5vTqDrykNOmOR1LjC0E2wcBH/Gl39upcBbki9f1yyq9X/4VkRmri
dVeXuliKXvsliB/4fKwxm1Cc3uBF2sejVxtqT93EmdMYIBQvM7SMfphCFj97lMgH
tsOzttiapqbieJKcwbk2UaA7IBXTLuzGrcsvxJj+oeqoL92ZG8rch1qo4D4hRSPv
ERYKuJebeve5KOvRkCt7xDZ0t7X6ug0C5gTcwZcX7Rbnxw0on0tuCYluu0+YnoNY
YNAtI5Si2fesh2jVPjA5XHWpn5iHFGWlmxOdgbnPUnxOqpkkVzLcd347z1Cf/z5T
2JZmqGWi9oA5NBYj8B2DvzQ+fDG5JEJd+BwuBsrvs0rJqxORW7mVPUwTXTm7AuNB
hkuMjRr+jNjLmQVHiqUfsoTa8aQgHYAnGlPcWuMKERSzqsj6n7BrEycosSELOwNu
gwf3uvmHVO3yb9+WmFAmVmbRAZe5ZEfg/sZboDtxz80FcQfxHHym2ef0dOf/7EsF
cZZl3zxi1HEDXvxyfSKDiPMUZ6lsPPCT6PCWZI0BR4AwdChB0xLd93F/fC18F/RD
TyRCxxuzAwRMj+4kfCpMDWtlB1lWno57RY71uK7w+uhF6/U5TpXI1ig4z7oQJueX
Fk6ClPchrrSDIPpUQUgAoWlczaaVZWRWpIJPfAGEKnauO8mkKDJW990w6ppeVgxd
CRnmcU8maz0ER03idO8idWZrTMS9FJEVIXlP2EU8LMvcIDKMEh+A589o9B2V6nyU
CJI3IiGLunHFWtUUTG9nGXPG11MBuhOHHlbjGcm7HhevSx3AqGtGcZ5u5ZYF1duV
U090zx88l7eV+ayEj+WeUNORJX3cnSgczq5JouQ7hLkgK7BWegKn6WiOczFTQ7Zu
PrYUMFV7ZhXm+tRUnAllB7HFKImrt7UD+baVlnKofqBcZ1Tsx952JlaQPX+xroRx
DU7Z+UYrVGxpAZr2aVK78+r/ujW2VqI/Otg31M2MCJfqcoq04BhlUqRBbCoikET1
o61kCghn6lC/JW5eMaJ6cCj+B1cMQeb0HNsLlOR9+/dQnJaJxm8JMZfd/Nlev85d
iJV3d6SY3HlzGl8s02DIbSoEj2Da+Ih5Ahmw25hHFwL/GVl6FXF1kPbWtYDTECf2
A9xWqg6KM2q5kP9pVbCFWxAxHaeqNK3260vGaWKizv4qC6/j8/O6Ys470GOH+jH2
cUqNipMnOdxCnY2k9bq8yUhhWAU1f2ZStC7CMOWzIbqX2vQyySS14B0hNpK8DW/5
FS2uskZBM2vYuVjU5i9FqI39yx5KQgLHY+3/eEnSJAKAUv04Dx8ctf9oV5ZZ3mKs
lAmoXGYgfycAymS3wK8gOf5HR80FO/v+PfajUTzKq2sEWhnDneTPJ4UqctngmlmA
NtHxjsF3kJPmW+06dCT8YE+4IYF/pvhwOnOKM69zC6102nGy3DdbNLo2+4yiSy12
QhaI9HUIf7EuJqJMu5sSb/tq2RYu4BIQAWThTV7/sVrudLI69j/OyMU8TprVVvwQ
k5LQKiP243nF1KBCrLN8SnFfl5Ts4GySWnkr+16TVUETduT7mdFnzcM+GC9Uozkt
0AFlL8oUIAj2xq4khbXBVO4B8nUg6hOCIFkZ2KWcMZ1NbnpXbfiYbAj9poA9ttrD
i0TXqWI2pwWARo5zSAmHjnMdPp3UN+dW5l8Moxkot6/JzteoBAmcBjU60dl9TDv+
tJaybbDkk6ynQxRsGw1XeF9Hxyz/pecKs3Ozmok946lFXQTxOETY+WAK72XDlGhI
9z2+pKF8SMsE39afr9sRFMiNcB2Yee0rwtQeFFXWROHB3uLMsujVYoRDGfk37LTZ
VAySkGCWOxjfUBwxBNY72wxiUPEv8AHCij38ZypZ0CRTMSIeTY2fpv8tROWw7gUO
DzsOxgPThDoxGYFvcAD6M+TsuixZprjDWpkzjPweJr4yNLbxSSjTno1QFsrV9eK8
ohK6JAKyf7JAf+4au2CvQDpNt/RXcg2UdMP5i631R810qR7nxzOnIK5HJwPszxsK
1wYTa2fUd9QK9FZiYVaxX8Qq0uSrqiuz4hpqKL0s58EaegIra+acbjbNujZ3+lsE
2EWBLtnAHCx6GhDSYGbv4kuBXi43Qz104W4jRn9tj0Q6X/pyVt43nKdrdA4cYdL7
DAwsTZDm5C9L92vo9o7dQ3NH7+u2Iaa1MqHyfqsfSfPX2CLNkz5+HnQZt5N1KGI6
htASWKAA8OxPn25itHNF7xrn8JG/wv4c2RGq3dgSIPQhl6w/gDcWrfcNXvCBTcT1
RXw0d5PowJY6YmnSSqafEBXbUm4RRoKgT9TdrIOMub8bs/LeTUWBR2r/C+gvJIJY
tuS8YHoc+5RDMwlT6Gt67q1/Cb/81BzsS8zy5mH1OpY1iI8++VW7iPTZYIiZOL+H
IgNilFed6tYQNLZSXtq35C4ehyeIadjxfsGRAK33XdZR+Q8HthIaGm3rjFhzZ0mU
9LlHayqw87cFlaeN/Y7krKByfoXGR+av063eIcM6IaamP5c+Hgo2lF1Ygv2wQ1Q8
bt/0ZMlWPAEy5tZFU/1IYngoQtwHjS89/MGaM0V6O7JNdMVPD0oU9RTfqfj7OaCo
L8SdW+0THFm59LLuxx+jPPdgv3ZcYGrfmfLiOeeJgq1pfLwvGUeSBVp4oc27CnYH
mn8bX2+5T8lWgt7/dAXz3PboC/Dgi3AeSSyEi8lAbpmkiyikOhXZJq9EMPnDsmek
fCcF2v+VdbG5Rbl+0ev4L0seS1k5HFGkP8/kfodXCKpn1O1xZQ/3mmq6PaBvtn4m
IhCTJWCn3OBYFi61KdfCVpQ3fPanUof/6vwxDa+CsfSKgQKEFUduhQw5LfIYO6fg
VoeLP4F5kMBGKYW8p+5mE/kiOIyii7W8bUrvQA5qQTvay5rMTD2YaAnQe1pmSB4X
pVHF+ZdC293r5tAjCZbo9pAIYUEWqspFQZ+8AIBuueiMnzi/kkl0pzaCwlf/GJeL
I3PR3Wr/w4GxAujbNYh6HHBbBdx3cDlvIMLC/01AcgGq2hA40s8Ym3kS4CTZ6i1Q
nwzzbn2ncuTN/EDk0tvAnajKAaJRvECzQSOqcD/9HNhMJDpllruFtatIY1x6qnjc
2jbiKf8CneRwICPBf41IzJTN/wTBo1nGQadAo6HloDoVhUzmUNhjZUtv0t9k3P4X
mnFa48hkutEtyvLcXiH33FvYUiBZxj7KXbl1eVAVmqkRFGaC6+0dmGwJJLjYZ2Bs
ENkZppk6EvPskJWFALfESyPc0VYE8xSDaUKzzPnxqMLrwYeYhR5ivO2+dMoDJzDe
vhj9l2dyPM/52MCSIx8RMR8wlh/4UKfJoOHhNUCmF9OFvihgc2fNYejbf+LEuXPo
BbYWi+C34nk2fZYHkSC9Md2RP9LGnKmU1TzAQY+B6y6/t1fzUAkmqezoWjre09jt
FYy4iVXeNYsl5OIBvRkdBtX89HgN/WX2hFZOdxgfjqz8lI688YAQVcqxX26b4r4w
h7SwWvw6zsA589axaMJtkI/h5nkdtdO69sbcXJVsp95HI0DcwQgTyP4E8YADiU4Y
5sRW4jpIMB4lb6UGij8D1emDpvCqgQu0m0pgcTj7SYM1A4r24+pWBFLvbZEJddj1
hPlhLcMU4KUQtfjC+Pe5NgA5XrVR9nV3paYNdhAS4FMBq4vFhIxy84LSt8sqaijP
FNOksttvJC5uPvi3rGwEEy7sVgXIo6JB9SfRKLB3UKp8m32abqvcOmsutqpbHiph
BZo+bRSR7/woUK2F0GRIRdDJRj8ghRa6RvR+ciuB6850VK7PQDV6TbyzWNDnAAyI
GLZrlOCe7QJlN6zm8PIvtrzEHCYl3MrHgDkFcz55ninBhhMr6QWm7ol9YvAlso3l
VZQ2OJLFUV3Z3Wws++1iTxWIIjR3X+Jw6iTLPzvmrMtqdoyYknsyAlVIRIGgEztY
OTFdL65JQ4P8AfIfa0kmQsu1rNMgm8gaQ9lXuJpQhlIdXXcWgf3DYRe++oBWp4WV
d3IsaYJw64OmsDMXHsUjGMbgfvsGB7GzaYpNNHRorDJqs+UD1p7eOczsYuDxOj7P
KEQaIWVvriE2+ubG7+6MHIaPaKRgiOqL6v3bNiGIJEVDb2A7VHvdRJbDEX6jeZxJ
u97neiR/uBlyraSTdK0IEn5gtyu2giRICbcjK4NoXf+VWJmgt7jz/ihGW6ky5cGT
SgmgLEkwipA/tTGrSUSgdqOypM08l4iHRs7dypmpfWuZoCAm/U07qRPrAQCevKCO
QfKaPjwILlTkYEs1mz4/1doifRclu2bhBaapSV2NQSKkNIi8gzBNmZp04RGbNnwr
uPU5bzJkHaIYa6jPvP16fJoRfdtRtcspfqyeAp9j8un4uasqm/oQwrxe7O2u1Epv
zsKrZ9TYrhV9xqQ0H8Duk0+sVnMQOY7cXoJxvlEca/wWVMGubr4yvI7+wXSWKV9O
rx/2ihWSSf0oG3T8DP4XrJb7O+IVpnpphZmX4QcbxZ+A9jjO6qdh5JbkeyE3qCOy
jzuPr3e0E1QV34mAa63B3sAf0YerpMpHR69t1Y0tvAOSnXw2Z52jUCcm0j4H2Bwx
Cblqxc9TI/DGCwzgIlp0+wBC4RU4YTfl3Y9e5NflU4jbS0eAbE10G/SejNvUyjgb
bHxvsqmPSpqv615Z1Whfmbhqu08hy/cbASRTZhDvveSBe8VYAwqgbx6pKePBimQp
h6z78rsUcw6nwfYXjoj1f28DU2hpFNmoKtiYg6yKi7xoCrpAeWM7vjA+5OkuHSZI
qXO+Fby0HrjUJWNkS0TkaHUAS+fFIgbMCaWU4V2nLlxNMDdQD/5Qepxfzkhge1Ir
HGTP1lDnYzQNFdlP4/uX3pYh5FVmhM3ha/OFhh8ZwTxVtoAtp6VWrCYbcTtJTnyl
Z666DyLSjvJeML2kMKhMUY/UcK3K98vJsj4C7pOzIDRjcasIPMbUNWq+wtvMIiuq
t3OVc3lxzpzBjN7qP6MMpnJfjaYzYU0Ck1iUyhMHb86SS/+F56WE4UZQo64uS56E
3yQmX6gKDprTLFRjgJJgd9fGo1ocIZc/85Bs9sUqMoXYPqNYBhhLtNrrHMg3CF1x
19xmr5asVBea0lwwljIp71eDb2AwUqc4YWEBWDSUZyYTh5jEEEIq+9pFCEUnZ0kg
raAsVTTaUzMXAty+QX7wr01AjwH2GNfvbnG1dO8PZtd8RTxF3p0w4mg9Fs1Bgogg
hEGgLpnu5l5CV2b7m1DDvCzaxelFSb/o/aQXr8p7jE7cfle3lT2qmOR9butp56cM
OGinOB587osj1hup42+FawWptZPmLWQt7CZDiBOzVwcrY9AXG8a/6ll0cpAOijvK
NpuDhoHIK0/ZFB5ZA+sFN2mB6YOpwDGs0HJ7jrO2N8NDAWuOtetZgdlMTwna7Pyb
vIgUPIm68SWTNaQAmMpCaqWYprB633PoHaM2YGRkHVoARzI88Mcl8AQrKMqY3HoB
aHUugRVHHxAdVydSgbPQsK34ZbxC8tUIMRQNDaOQTyXbs0RjVswfLcfwa82D6z/O
YT8Fb6nxh89HK0gy7SvtQU4ELh3boNlywQzNLLxN3z1f4COSmVAA+qSu/9NHJCCk
YvokwSKBB6PG/jwAD/p9AKGyk/nlx42ij640S2aXJUrySYCxMb0Pub/bzKr2H6rM
ULTOmkngU7hKv+HU/t50L9WpYkGK5mujQPrrwO9ht4ORRR+q/tcOi89omXqYiQ5f
vSFQ9xhKTiX0WAJYN0+VFRa9alF2bDAy6Y1d9XWmrEggCaXHdpvaxVf0TobTz+hN
o0LKvKl8St/YlqXmZpHaCLhw2nCQE3PZOB1HuIlra16Qyhgs9f9fXbJyEeCsgX+O
1wF/VltSvyF+KpJ/5xTXrpkQ8GNCLXMsY3rgHTJsyk8gIiIvMPFn8KYaYeS5tg0z
KE4y5QOjeUPSLgDxTxYMyQjlq+g/kScP9jrME9c7manE4zIuVaM04CB10uFam2Ck
brg/BMe+Tr+sYC0+t8lwOO9S4kCxA5MGD9Hq9OGQNlfnJMbd2/jzWNGmj/Bbpqsl
Grx50mnos96Wsui56PjoGOk3ztcbjaOn5DWAqjvBxQzIrqRD4NbqjjyRAERJThN6
u1q5AswnoRjlo/LkfWsliKjxy30s+qz+CM+c04XN49CYyvfZwBYXtScNhMtlVAHR
Ds4YOEnMA2JNoU2QCKLtE9+82qSICyeVmqpEbL6dhsmaiwwjYg4BrIfys+HVM9iQ
lav7QhnIkzEFM6+Uzu+2HW7/7W6KdeUYcN/KOF8RUlre9R+tL069owgBinmrDyaC
4CpRuxbL5aiewbWvX2EzA/rw2GQouxBNBWGGiHEbEtgNJRE7V82GgYCvByH9zEge
okCKI5RiHRs4xaV2AcyGvlkO+kP+ojHjqAY7cXN9EE1A0cnPpNdolLMo5oPPWT9L
IX5QEEAkGMKzYA1xF0wXFepkpTrCNmNm/8zKPK1QDkdYu0ZP+G9PJKYAAD0ZNA6k
CmSiEb1xXQbN2DtJz43hMhMq2HPkXvU+FkAtVppjCUeEj/2+rZIFmlB2bC/sRQsp
rdk4cFKPlDff/XUaAvlP/FbG8O7Q2lRgglUKusDLSV840tfDN8JL2X0Zgd17wyTt
wzqtHRffoRQn8ZEtnl8cROiXu4arIvprYNkOzdnAEyvff2JpnW9+q3U0jQsda1Oi
ml/+bXMeyAwZH/+NQcb3pSM0Nu4Ht5bMrAUncsMKovXLrXgQbpulekpCRxL+K6k3
M/3yaDCyQh5CznYfbwQRTjtnCemR49MfdQK+fIUadfGNuOg13ae4F+1nXfu7EDe5
M3LWJByYB2CKzbl6jIuaXH8bELm/PiYv5aUM1tPJ3iHQyerz6SgK2ng0CuJLPPLQ
QooVSVDXQCQjIlwOMpO+Jpwb1Tu3elPg8OTxMP88gkt4mEuGS0N3ccm+YrLK+1pJ
YZ0KNJ6e0jlMvFVKc9LZxJs6YpZtU1FaGfZ/2E7mUEvZEJ7pwbRCkvEAb0GSAu1i
iA5o9YfxPIRo6wCjxHuhU7mpiqfBU7ULocR0p9WPZQbu4FQlrP7ei2EnKcpu8SMG
uxf/cf8FEpjI3u9rnqF7rpw6iyZglG8x+rWOzkBDUCxbBxYOSYebfcMfBD2+T9+Q
3xcQ0IsALuDRrO/a+m0J4iiknTpyfOYmWvPixduThgyhLE/X0gfAltrgbJL//aVW
C9rQ8SuRoDbxuqjA5qKj7KDX02EOgUWK0JKGyNIGooPcpZ1TtEZ+BtJZyi+KPwPm
ZrNar3y8i3LMTnGaL4/oSXuoKNOR2XP61LN1pZoG+lHG6428JgZwBPAt+9mwtxIO
Rh8o3wKQJJjqJ7QD50YsHc0OP57UfMg0OPKNBERTugiL2BCeL7Dj5gi0zr5P0FKU
/xNGqjJMDRA25fgaaS3GIIoFLmNGmLymL8EyjtcCID+MEQhX/OW5Asx7gPtpu97k
Z5pxISxsc/ozUsmTYbEPeI3FEOdcqilhISTMKEIi4BaKVg4RHbRBbkYUgQxyr52y
6i7feWCklbV7WiiZ5Pdedq8tye8wUS6UXAg3DDHSl/Rfvuew4EBS3/S/wDojAjFs
nxnYd/PnZdvcuyXUCxin18xTMj0PXagmtsFPUVHhQEv0cMDH8VYK5JBIl7wXNWwg
hSs24stKHV9UWuL2021tHCxkPaKyuMBUHHzLY+6ohAuNIadlUSL+9qvW+ptReAqM
tusLISne9mPB+ovyEKxfa/qFCCeGoudTx3LyWYj5gGGMK3c9nDmZwZj62xpH1nA8
RtQ1xDzeEDyDmdPc8Y2BR0sKYRm6vwqr4rQcAccF83H3WUrdqsH1H7pQJHbt5GOb
LyoNngJcyJRUYKZd+uGCaicI1gmlCdV+L6VMqnRdxd6GRtKJY1rZnS01E9Zhp5wB
iltz3PdmkiP/imc0qoVpsDXrXl06UJ9adBirSNXH2huS3poulK07oxulmA5YtqvZ
UUdtOShl+nfohOi78wuHEjmtawYU3V+puO3M5X42eDTKYcuH+b0FZ313madg/EPS
TcimYHduvcwaRfKDMXJ0cPR/IrrAWV5kLRCAtNDWkesdctHp/4oRQPXB5j1nRAZb
nhXNo71KGzUQEdcPTN2dSb9GjCwTys33MrOCXvMT5zus/KxKFpvHiUiPdNd8jXGv
I5TFH9N5oD5uaUUc6I4M8dX0mOsaeqs57GvhTpbXSPUJiGq2220boksg1BYLuqaM
E4kVz81vxQoaPTRrp74DQcaaoORYGOq/K8L7rzFllrqPZ4zoMXK9H62OWAccCB0j
LuVERaUsuUt6tOUmuBZIzeydrqxb3wFogyBn4dx1UXkyYAjOvdDm5at7m9KyUDXL
OGECVs0+ian02UO8nxxSCyQ6vKFlsJ2cAT5YEidyCi8oKIpP0ychetpKpiAE26+W
atxta3TIYLJJjqxLdttFUpJF3B8W7waRXdqitE77m+VVKJuaygZiNMl3cmiPkegS
AuIrU5AGpSIZMgNac2A8JcXHDWkEctiry5gevnoPxjXmL7xCjcllK/9mZpNtT6ct
lEhdX9dvfVTEG6/BaKbcgx72E/2iD94+5rcee/nNxUwX+iQEyvG7kX9Rv1P6oVBr
P/8iZ2ZNOn6rBrVWgRYu+Bng+JUo64p70t4K1LmA6bKIJ158Ic5eAiJoo7ZPSpMw
XPLSzR6Nqf/UebH3z49accdGSLs4FUfZtsdWvfVBFxQIhdHuf+itqLrKI7GUmve+
1oqVihQQkMlYY1Dt+/Xl3jf9160EF3TZsUNpNRlyE5JDzspVP9nVo7GADJnNSmbg
sMVKWHgkONmTELC8f2lQIRAOz+LY5d+vgFTA85hqkYHoa4i5Ti7N7mEukR8c12iL
XJq1fkp0xZfZ4TK9xR2+9hr8SFLNdIw8XKzaeIBv8uh3pFCQa+u5SJrHuedQtXNG
N3JTolenhf/Qt6dRbDt+xiUNQo6MQuaM92I2b3H5M7dZYu2MsB1sxV02foQb+XBF
uGJBnwlmFPQpeu06vdJ+cZjXP7gXzWncYji0Ho7f87jDQAvLpiptUTryU3JilsTO
XWmD+pEN1q3clzY/4YuKMPRS7k7NTToZEumA+jtG1cEOjZlSswieHsCad9zNltM4
9435ZvM3s3SZyQ874oArgl+LvNpRUphggb0Ef0nVOkXFszdpFI3rN9NsU4Ry+s+3
6eP9WiO5wYWZvYbC2eEcQEBqD4oZT7+dRT5NmX0JGX6VqIt7lnIY9A9+lpmGJSHb
SNuB6EKCpeU2CbNRukA/oHeomr+UsccCzAkb8++li/UMpREWnX1A35M06Fiu5yF3
ASxxrB7800Grc/eIoqngMJP59Z2a891SJpcgaLc6mjradV/W402pFfSwBd1ZlhvE
Uc/zok4tJAfFPTI0hzadLdljoTaWNmLqPbuiCfnw3yE259PsSzMU3o+//pyJsnoN
Z2lYBzNZPYT3CoFqKUUSCFJa2iODrfJEe2viTuhm8NQ3lvhKRJYUkkEaddu7Q+5Y
ohwYT0f1sFsGyDCT9FhK/RdzvkS+W86vpm+gpEopUA3UVL5LZV+ogdxjoInSbcjX
b2NqBEruyohPcE+tm6bjXCh87OqNAsplpjhtBFplf4fz1keHolf/+LA9qONbqIq+
3goBlT7X/OmJkzF6Tv9qq/MxgBn/x+YWpjV5HKD6MYGPt3q6qXzP4t9Z3sGAl8m9
r2OCbLNtd7dVB6AfGCGtObiHJoQ7X20rXLJdqEVICo04yTEbLZfVkXI0NBxKQBn4
sCrSZhVJhZ/dSFwXNPvuwS4TjzLyOkBdzESXZURayXBnlxPNutq7OijfA3FhLgkm
VldpaIlsFX0XKi1IgMdPC/tuLWluI33A1M6nYwTgVo6vG3roAt0RvCUaRVRrcQbw
eJl/GslTcFf1eAWXg32XPe2JbkFmxunULEhSBBwc96MI8u6bWlf3gmXw/QgS5iwR
jzTQHEfASuMKrwrOXEjnZG4j8zISq4SZScPh5YSSJO7kyPNb+/Cv/yVYfg8xpr1J
rGx9ul/j6XC2NnQTtAdHR0Bq2uZjgaf5qNgcN2majUyxJQGbUwXLQCWZDtHgfdFZ
Z0mrAMep07LDn48kdwfKqmsdms9nwBEGdvYinySHtfdK3caVX0dslYIt+elrGPnd
Wk49B5LT9CPXipNiz7Gm+ZPOti8vjU4/1py0llasDs7wuU71FscTodltQhwcMJa7
oCxBbvNN4GOMHAIfTybgq+OB7OU8Xe1FHX5O4awNGq0svuVxAHQ0ZqD03Isp68/5
s5keKj1TfW/0avkykECLnKKJFE64DuuKGwmPj+ILmDtqZcfjzmpyhG2LaPNR07SO
omgHd27h7sNdiCcE6ignL2G8P+ZmKii76X8CfwZr6w+DkP5+bC/U38Wr3vh8MMoO
swtdZgb7fnBOwdaz/JDw58qyn7YLou3cysmUJefOGF8AfCCjWhQLaLrjlG84qM/+
kXgSjOOp07htfX+qp4uC4KYF0KdMwkjJxNZKSN2LqTxscwkagmhXIcqULVKKshLr
R1qPcYPZ3fRsojYsfk0dL+NrZ3e1ZSvQQhaWFd7ASsdAnTnw6VKT5cOIUf1jYrNG
a4WIzt5n6V8SvAp0KTczODofGtSVQ6R+BbP2QAeiTPeIiPO8+a3VNgXDDb9NgfHa
3zdQQ9k5UErJY6YnfR0ak3bzuzdv8Fb3hLxGdl2RfunbG3p++ORpdKlOJUOweVgK
0LvWD5+jjo/d9U68TjBS4oh4tLrdsRFjaVRMT6qTvec8aWDwqZSnH4PKkKB1vuKW
RJB6F3qSRh01ukjCd8wYgd/qp5XEE2VEMj0iu9QSpeF6O+la+J0NzUTmh3tV/mR2
fZavMKhWLA2482IRgy3+iaeOIAa7/Rxoyx6oI1EENKW/VFp0mkUbQq2g6Fyc3uTp
hoipDtx8oFom1DluXEg1VGhfEATsEVcL3GpztljBwsfVvlPLryii85CQyQK/1BZ3
UYz5/X/2UMy7hH9Al+jb5N/bJA5uZHeeoSOviBqfb9peq+H0CrDA7u5nKZ46Y74W
i75grut4ZYTrizc2Hs9n5zEm4AboVZo64NN36gOgR0f/g2jw1FFUFZTT+CX/Fg/3
oDf/5xJz/DveU81DNLivYIkN3Un01Q9ABd4DTyhPmGJqn+V6leTdpYu2El3/Qw34
Q3ukiJshkJ3og0CTzusEtX6plo+xky36iWmtVNsswzW+HWgt+DRDlVtLvgtd/1mZ
cC1IWLNDsg8aAGSjo+sJYSN+xQodIlyu01Cukqo5mZbQwhBoEAR9m0VkMGDoqqZS
Lm5AFLHu688p6UGYdP795Re4Ier3GqsjJTXm5AiiOAW30arLmdJA1VKM9u3xKBPz
InmPqulagUQIYTEb4uJbkAeGxH2k0MZmWYBY9yn4lhKlmaon9oxZDvB6yRvCBU5Y
h3eB0gQ/etul7aXU6lOGF8btcOb090s5fRGpXhXCbmpxDAvbuVkNo3PMIdv23M0F
2g/SSHWhnG886cv7Mgtn3f4420ISdh1II7FcffHH3teNQm5bfKLTw89fnAAywnA2
EV3lYnj6DgVj+7zQG/OTMFThoYGTcwXnTG4djCIxtZDAKRHC7xWzWUfcwVIF+/AG
/O9mAeWsGefSJRc6HEmCkgrlLSfPM38Y3E0A/u3vYiBF6zjxtz2XfuJJHHUAdlnX
fk4YzeP9zmcbAPq/IpNIKfZEBkDYY/fHNgCOR5c9O6fiRqHmhFSE+cmj5KHWmA1y
yI0LCOua1rbXbCC2bHoQHvTL/0T8bVstN3fQ7Dp5R+mMi3HFWmfMh/yJ1Ab0RZh6
2H4hgf0lsaZ4uSZLPummFng8fFdVHyu7tEL6kM6j9d4JoUHAUX8DHMejKm74diAc
KbQm4oUSaEELEaRJQYtSTcdjui5VLckIQD2GcRvpUMFDmYjm3t/cHwgtLuOlo7GD
+NsOpJs90e7eMDDcJjc9oQDWiDedHh7O0V1ufel5RWI1mXJUXXNnRSDuCewCo9Qt
8BhqONH/4LicrkLLjK76l3I9HKu8Y+6G6L7OyBxyNoG6P31/k/aNIKZ2ACnDum7U
EJKQKRpU91SCxnGUQSHPQBburJ3kPNxM7EICt+XjT6DNZRI5QZ3G1xwf//UtnQ7n
wHqqudE/uAd9kc4M06jTkQnjB5cvUmWk7wI5UPzK8XFVnq7SoVURCHbfrV68Gad8
hq9MsuqvUBca50rGhxjfbiqEOSlcyPusK//u92UmlYmkS9U70XDK4UUHjNNGtuvu
fl2Kqx0h3Cvyj/IZYGolhWleuxahyMMH9b//n74X+C3mOFIBMGNB0uUDutsWxP6O
L+YTWZJYwREagKQbEdCTixa93zJQaRIlTPZZkcJcjigMOu7sFYvF6gSgpJ6oF/S0
Iu88TLL7O1xmrgbQjgTI+KIbOgHSrLeRpe18O6XwjPKwjimo+ROA+epglQrDzWOK
j9zEnWzm1PLvgy3IK4cTyH2UQc94/bpswjGm4TlwrANgeP7mh0Jk2GpU8+OFYvAj
qSI8TmnTldHFSjWi/F1ODr8WbR9XmUFVtWiI2ScvzbE4F2lpx1ywONGzYH0jGhDc
/3dH3ebkPE4JF6Z84YLzfppcdYaa5gRkcKDAwVmkmMN306t1GWZOg26E0NelZyHH
Mbb/NYZcFtRW9XgeXCLere/U+/hRY4jIXZzxz59BLLKbEB7qe8D4oOlPX6AQfxfe
SSAlyMnaJSYF4AXlRybhykCv41zs0AY6tdKcGz6r4uCh5WiB1QUuta4ItDSGniji
YiXZeemhjcUl5QwwHM8g9A5qtyCbzJG9p9hoFYwzkCbFjayDojGlrMYDlwFOy8VC
aOYl2qbohtpeKqyjCAp8IMwOdgJpr/RngjuyR6M1umlRJ03gF9le4nxqm+LZBuX3
Cwn2Zei+/V8sLiHrcUQsQQ0IjdZpw7DF2UTMxRNx6+rR/20Xx+KVd5VcEq0DsR6K
5PIMk7hQbJPEmBKKz+lZve1+wroT0I2GSJPMIrTFIGy1BfqpDdwMA7IrWA/JRAi+
7Mc9MasVkCZo4E7Oeey8072061wIbrvml0Vv6gsgfH0p5698M4w9CAastlsWkt41
3SH31UVjhkJ3Fh56hEjdLiA7C+p3OGz3ySDPiPiXNbTS3/BGlPfxVjuDUANaqVxh
LtOQ0ER8N9MTt0DU813rplRmdyg0UJUsdioufK6gD+hMNWPqwvr3UBkuekTT28Pg
kOSWUXDC9fFz8SkTpCot74dwNnofueVtwcVwMsu6pU2s9znwOAUl9EWDQYojA63U
E3VxKB0SvNhvad3ieae4dbfw4z2ykK27Jr1js5eepybjT9P8t8QB9GMYTGClJG8q
S2rJS04C8N7KLOV5/0ff4BF/sUL0UQrOu+iLTVZYtoVyq68Czz3t4IXfw4lokKLL
O0T/WQrF1uQ6upWpXEobmg3t/FA7Wt6+F96ShtQ8eix5lYCJImpdRB5QsnO037HA
m68wcPAXAxlF2y1cCq/VPEZnJmMNLrQizzs19qKQ52WcNXl6yFMIIXGJkLlG5vLp
g61KYbR8+svil302crsMJoTCePZf5NY1AsZfoBdHSzCcTdeyfQlz8f2xlnb16MWE
7KkvTqQL5tAql6KAyQxMj0KjaVnDuP8D6UEzEq/8lytjUq5opgu97ShusucVRD3n
iDtH2g9TsCaPYEoS/mkbgtpfnD5vmhkYb9ZYKutI9e5fLVq5ixpbYDRNP1fq7Ebp
qLxq3F4r7x2boAvi3sAB8YdDkSjRNHiAV86sxcUSXTy1CzKlnXceIQveRJezrpsf
KCGlKRrwKokgbHZhcC5MCnwkxLZQkHOJjDNiBcN15a4V8vpci+WRlM7piTLCA6W0
m3PM7o/GljoAD8tKcYI18Yri9OkBBUVfSC2NDW31bRJVZe820BhVY9D3a+3dxMYw
vpvkGe9L36gKcVWtXgqRThB6tZ+JlU5iMrCKX30HafLDEORXwVs/OpIOPJLHJkow
zZrNa+jgUuTrC3yRrUPWd5+NzHccu7CFIf3a04D5LL47Xb5LbodQIV1844oIVQrO
fyKqCDGvobll4XPsD1z+cJpHhMoMVqLa5ZwcDIhIugytwXpv3frSsHbVdHJlzc/z
46lvRfGfAU7Q6pwo4d9vqm5NtHbBCyg0dZBADFl1DSpErw0BieMmL+6XVdwbv5Pc
V6daXtB8hJ52akqAC+g4PCVyIhKO+eWilb536TDlyWpy1ZiqtLT7h2sHenWrzHTS
0OLgh/0dSEkf8Nh2xnUMH4FAVBLbEMXy5i/8/Y9ZZpYbEKnhTu2jWJVsQX/m6YbN
9CrsqpesXnQZW2ylukuosOSDN33DjDcb+loz9q6JLzkUGXfNFS9nbFr1YjMY6n0M
5pcvmOEpV0R3OTUzkZ5knWIRJKEd9w+whUxEJhABmYnkWQLkhiWKqCcK7BFTMOfG
2NEMwAGIUgy6tbbWTHuYSdow8wgv3HV4IUP18kSyK8wHnpI/cZC34v3RePES4Z+y
mBGeeXgaOb81ODURpxbHXCSffbD4LAGNEkze4uYwGVdDd51/xKWSgNnjjoJ2yzrs
tmFjq6iKlfaS2auFfRmWJdg/GU4YmAuo4ksiLz/sLRaz2k1k6ZwSB+mrzE6UxvRW
wy/uhkTd2mT8NxC4Nshud7hgojjF1Z1fBWn2H1e7GxL01Li0/+boaCybf/RZ4XmL
cXyd1Et+6dyL7mTamYRVUxkVYnCIpvR+NwDkMtSqxEh3KOu3EPRbKUWSPNfTReOm
9mJkhfknBiufQmc5h7IqZW1rDoVKSSj7uvx009zFp8bkekXUDe+WNCMH7a9K6lvA
LKoJwQgxiXGLwd8RwtblAJQ+/gNEsw2WP8zpNBRnQ0JsCwLwsF1dyETOvDW9JqAX
f69DC8FqsV/IrRcbv5kpJ7OBjqr8kemyWo5U0pLlGW9BZI796fj5JRov9sTFNc00
O/vmlrb5zFyB4xldzFK+eyAtUWdgp+WDtji/IvPU6jeu41OF8boHAF7CzWthg/Oy
jO5Mp/lI2iNZFFtKSLcWoLmmQJQUwYL9u1ElrewBtOhYUNdPg4H1ZTzp79mR733o
Wq6dpSiyg2tXAQ2R5EEWAw3XdL5+erZPKdjus8Rw9N7Bymc3uzxYpqnnPlhVZVyT
rThM2icHYCPKK6KbsRf9tR4KmyNwh7TMFxTJKP3DC4OedCGXeG67qfw3bm9SwJuw
XJG0T0zL+niFSmhYXpgK4KD4GOxkglljbL9gsgsyh3ec4xePXE3cUqjxYr8jErZG
pMlRUvmWM9Hek9Ayda+bcn3QrhCPx5Zd5AXyyivJH/MdYxnovPeNnJ3v4A3VM5M6
S6usnTBADMfaohGWHINHfgH5ov+wottz/hve7PHaT2iCSap+nKB3sSBZkmQywMFo
sn2wUo6q3odYuVbCPTsDr5J4XRUBVA2BS1CNoJXsJza3E0fZ5+Hayj3GJW5ogAlt
VyFQ9aEf5+qQjWTPyEImAOiq1o9B7OSR2mRGzWUumZhGc4HJ1dkJjIy1Lj7oyPuS
FGw4Knb45YG4rmNXtMaKunNMBOuuG7dcQxI7yUVdWeaDZxJ1708a7muxnp9i0ZOz
0yM4/Jgt4od7WyUzTdKM5m1iSGrAfDxEiONrNFOeWjKkLeDBAwpt916GeOCvkg2W
HLQbYN05N9cyL1OHUHgLsC0qBlTyJJ11j6e16F2AIoX0mlzUSnOOu6MMUF3guD3V
PaY9TzUbw0yw0pRa9uDMnW5AZY4n7XUj4vzxf4C8MMCQ68Z62c3+7Y8bYCn7hbhT
OSrpNv9+fdexstoFWxhlnhJZtPTVZK97bbihQgY2bJ1+zwjcbf4d//CBDeP0wvm0
glJwD9eif3gQRriSLb9n8/YTucSs2B/mEnTmkEbrTjTL453u4dYv0uEJyhRGlFiF
qt1WJG2AfQAGwMGcfojhlyntLHx94xieDV0qWD+aLgfFaIBj6TY/wiH5lCr8wvvB
y5fEy/Y8idPApUADs3xoVCUYZpvEwOVRDq1IvFET6rpuehZOOFVeuS0bdDl5Cwbz
1gQvtCRSFd5g06JTqwHoecjWF35N6kv4K1t3SxahYh9uJbbp2wZZTxSkezbnFYoO
EKXNEFfdS5/c0Dw3ziFpI/VFd6b4go0J+v0dyHUFR+MazrtfhUtGP12VjhDuLgDa
uJ8qR0a4k6d++Y0eqK/cdoH4r9rSlhOPAhLndkCqYIMe0zjCZzu4obzzG1t1um0l
iXNEErFoD71fzJwEKk6LcmROwpNqmkqZVjGz30JPzTpzPHE25nnoqj6QJDunvpbd
9pAtH8yvrNwoX+LfMWg8bKsIXTKZJZYcXX6Sg5Bg+wkCBjBr64nIvwN8sElzUuRX
JZPKjqDtITHBWYSNW1uWKcjetsAHHom41CZtrIeo6JIgB5VQ5V6L3GSZFwgR5oWP
7dvYNkTD8BdzChCxJvLMu+ciZi4a4Ez4hEwpUHdbTUZ2YOH8ch0hTsGA8ksTntnU
dLX/oX5ud/7csgz3oi0HJbD4BJ0KfrUqkbgTyXSnEGSMlJuLhj8RsEigv+hY13LD
8krBQIuRzQxyMO63Kz504CoIz7czTbQW3iBCSM2lzFHqc3wmyD9udSSfd+ClaQK1
1EYzPOYEEQ8lVuAVwl5RROOvYlmzxhV4EjEdBG5BFEsMSjZTQCUEr3opZNjbXGy5
gEZaDqqT5bkJZvyrUUowNV7XDSUkjCeYbavYIvV4aAcU1wxsAPGoQ6umBak9RB+R
jOYX425ZdGfby8gWi8/w2vh00FtdIJS0bjdREx9EnyuIjz4+ddUtgQ7TjDeNjR5d
rV0bdDcq5PBJQ8I0jX4Nof190R5xiOfoSm1uIfxF4ozxLHm5gUioju5/pJKkjynI
PI+BUP5e82bc78a9wpbqyUKEIp38KNtdylNQOUHgCPx3y/es71ag/B0oZBNIJsl9
TI419lOTmNNBVDTA4WkfPFVc0WSch3I7prZr224uev86GsDTzKq82a6YGUOvjmnx
opgAb2q1u8qNmpEm7jl0IjYM3dyI+9K4qs3Y3nwcmbGZwqrqejcXN4a+1cBR689Y
3HgzyABnaXCdnNvFen71RfkzsOltLG7hDGNMuAFqYcQCk/hRmNqG6X2J76gIfsmN
MnTheN0CboNSaOgMdUmtglQsAvY9n+Ik2pfq6mqLu0ZE/nVZieQkVrhIeDJW6WBS
RXWJgT9DBvqgaesEfBzFpSEOLi1L8EAkt9XeSLhY6uJKm5UOUZBlWJwp/g0Ktp3e
W39EKzg3OE1ymyhXnRcO2kiKUwjhPHAWUnqxOivbF4UCSKEHIIua004Rje0JqGkr
CyhIZVfcLVH16MJZDdp9NwaKBWx+VkSH0REOnQW+BrEPH8j7ou/i0v4HtfYlca3G
P4MunAS5z2cGjQ0SfGrGwy1cVIx5CjjUMrTGoDcSAtRhFUFa6W8jWYUuLY53QqhD
LYxZM0R0RLZxTq5g1fFiyytDeGgWQNQvfSiyQwgjMjsJGVOIO3vHKgB/JNp8MiKo
AyHRKBiLntfy7wf5CysdeyN/UbBOedXWpgerbP4SPH0GjBN7r8q/03sGvKALpsWl
Q8/FQuVVtKzwwgHtdiLFi/WoCKTb+BrRBQ5DDvV4pP+9KA8plQ1t58NptX9ABTWw
yOiqNqyrS9g1gMA8dlB2FVlgwOC+gVzhAeL2Fjp9Wqw5AXKwgXqrnTX1sap1Icps
MCK7aN8cpbnJJxC3x/aHW58itF0v1Ct/5h6ovMt/dj1oIfgdhIZkB9vQGm1P5/JY
LPB6DGta7ESkrFGcK4a1wzxPjBwIuVSEM6Z4k947Ymezz30EbLh5AhlzKwuLMNKB
PW9UK1SXnlnYMKVvlRqre2cpsTkcu4U8QYvj/xQbdGPM6BPuY7P+rV69jVRqckg+
+uDGBKfXRdsP8odtuh04FYoaeroRPLZO1TbLLmRP/u64q0pSHZuUXlhck9N/Jkre
Igan0hGsg6bQvh5ATdUYfG//uDg3GyELItL0h7x5Lhtk1Gsljd/jt+xOkngkCoh/
OfKbXg8EocdW88hT1eoG3tMFSP2ShiUOT88a1fbBwBBsvdY8HKfBIJBI3p2rVSy0
7JKnDYxg2WQAqluzTbFxgzNuOtc5ecwXzHVr2XLg33zRM9kga9UZ1Qpz4JKvzk4U
VFcbGpizNJ0PpiU7yRWwMgP2VPC3wQjQJ9XO0MvEckIfKD1ZCSy28b1gi4ZVD2hF
j+UwutBDUSPBYIHnN6ffGHZvm6NdbwbW2kR+DAc+ZuAugFDVCxguqnExfdVsmrTY
NWChuWm9DFp8IrZcRKzzI/UYO64c4Rr06gbAMats7OEs3/VXb8GtQPjrwm53pVZh
guCt11TlZE5BXZeAqtYO5rVkThFj6wj2fjZKID3q32/0Ey2Dz2u+c4lNDmhGdWS0
8anQnx+ZGk0bhFngwOx5HqOA7t3XrO4yu0I8/HWL0Z92yEsfUtOg9N7dIqGJKTs0
OZlb0GGIIr0K828SIv3EmzmCbBdVZyvfVE0pvk9OYfWNeVZ43kxLN1Ih5gA3OF2k
aT1Er6r1y4s4EZteOekm7ia+lBFm4D+Rz5tF4c4whPz5bq6jhrLdDOEps5/Beqtv
4m1t/6QWvbPdtyH8qmFVLW1e47e2UdMPbCnQHc6TzdweNzuXmxSevwm8a2qrJ4Nq
S6qHdfGczK5ZTl9FtN2wGx+TkeoY8afiox5TUS8H1qcFSvcg2nfuuCK78+U8UAsP
g0Et2B4rktTaj9F/OJUYjqxulOPve8SjxYEL/m3VvbANnZjmfnFvM6mImDv8dGG3
QJFWkeU5JBTrb0nZUQGuXmwXU/X+GLyfVGfsk7XRA6rkvwcPyl4vZ+zCXcnqyE2N
3IaFKuSKbspKJrOv3vGcPNPLaB0/FKSlAn0loAa5KtYZOu/aIPSokFQWhDKj2sKZ
uydafdXSL8QjOHigQ/TKBTEYmSaxF8j1WTaCDDbdTjVeUbNSVyncm8iVXn9NuVl9
zHMpUM7rFDo+TlemqwrMVyYhK9wjN4U8m45OuwxQha0xt0EKg8miWA9UZ50ySN68
ZA6HNGGzNWVX+JLS5sQ+xpgSBmYGMXPRZFcGNjD9hOm6XrEyoB0zncmv4wfO6/OV
90vLCiWPJGB1Ns90Fmkb+IbEJ1RpSlJWYcBQZ6WGG/qS2gTdB+4X/C4EerMw3u7B
2Mmeir977CXT3QlZ1E5ipwP5KAFR7UHfS0Yc629zfVas/zV6VYRlkAdoTwxDD9Li
lnSg+ehwehC1Ca1NaJKgghMsBrZvMfckAxg9OVgwym6ROCbPZvyaCgQnOZK1HTit
V8JUfI98iDy6WvSYFKqrhASM0d4/OAe1Ks2X0lPBsOwS2zMrkS8T5NsxEFQOsIxu
KFFCyWhlHooo25hU/KTVvqCrakTTCdx2nAhxWGvEUorlBOadfqEUgCb5vm4YrZT0
LWhBUkD3CdsLGZxoYyn2iRu/GOhzELADbwxdVaon5UUe+1vT+OMXDuI/wXxY/IjI
H2mNCtmRqqXI/tQrs+AL782SXyyBP8YNBM8SpwpsBPgpjp6XHMmo7kWc5oR8y8GW
mo0zX27S47Bn6tRPIQ1lN+ieBmqrxCWVWvaf8pj1Cf9UAO5GybMFsa/81/fN4rPH
UGuDzC8sPl8eX0ArLaOWVLauXkgG+/oNQgbt8oGz9TRe8Hob8DAlDCM4LV3AbsUW
oJWnKUgpQKCRDWOMOuYUfNvmpP3JYXOhtQjXD+xXhQtkhSNenYB0s+wv5KiB45y+
p1gJM2vnbSbvMcG/17tR/CVqddcy5plAn904eCvRLTq47W9z9xbM10YQah7+ltWn
FvKw4M4X2EXnNOkQttQnKNOnKzjrGRwl4c8fUJXdWY++z4j3EiYJY27bMVDKVTTA
chfwNuTUD0OobxlB6WtP0V0af5l+JZbEONA4eoxCpjxECjrFHoCcYQMEw1s5Sh0d
nL8cYjhmwjW/BpYykBWN5mWIyj8n44a8RuCK1OnhmYzZzmdbe9e3K8ZOe33yJrmV
a6Rs7QFtv3la+lCKrktvp3sRJwebDywbWWPiRR3Eq5+O9iRd7wQnMNdgCOV4v8T9
pLETysC/K9JnLvDLlRbz7G+yuE2ZM1PxJvJvU/v4kFTp96m+Ig4zTFCA8cftugjX
lqxVOeINdbNP3jQLBqrJ8LYOjrgzuDn3G/2zlL5aRcqXTYIx9BypZrL2UjqGBjxd
eiMyykjX6Y7xjBvAQhS3K4jZ09NPFoSOBHysssmiBGWUtlz3GzjkXpqROZaixlc4
OnZfsyJXmxD/FBhgxaXNy4v36waopJOgvgTVrx+LVdu1CZLxuSlimag9yZG5dr5U
g043rlVs/u48vOvSJrKbau/ikgnLzXC7JtvZXncFigJdUz7dA0y2TxC5xxPQtxso
4U8zYa77A8NYALgoCCbXMNjj2nSnow/7TXjSQr+CQm/mim36qmtSSR28CY3k+Q9C
5M+aYr1wDm6UQcu2SUT/v9RFLnWEdc5BsVJ2Kss9/eR+5/qSJWjIltG+eP9p69Hv
eZAM166daY3RVSctPcfEldTMAYSF/DDNqEOaZ2Cg4neJS5ySBNsNU5ZrvVYvS7P9
FL4EEZGIQLcy2fZcrBWeczsle7VpyiVZg/RUd4siIk0uoF1hZPsO60VPFcNBzSct
Ncx3gOv0OfbfPwzg41KA3A5yymesNx7LQGlKSOeySIw3ZuGuXM+bedXJtgg+zvLt
zimVuf87443CNBSYamURNpxoDPtLVV2vogdIg1ILCwKmBtsYS1wADFAJVhXevXIM
/Qjk5uWxinR4VSEFi+Nj0p/b4QmmB6fukEMyYk1sVuwpxRzqyjN54ZOLZSAbW+gR
8XKvwmax7gKvMTvoPLu20JONgwtETslFbgxOEWE25JQ2dAEdneKZH9rz6ZV4MSub
wpW1BeK4kEaUyjemKu1aF4iij4Zxp8KZKICWHrl0LIjxNbyp7TDkQl/pD0cROsly
rWIBna9S68HYambmmVaBdWZcuBJ0DxfsNBjSN0arpR1vtnbfzdsJXuB+8eiB9Ozk
+dnabu6hLrvBpOVZTUg2DmIztofq5gOQCZQGZQt6OtDtUHLQLL9KzbelwhD7Dzcd
qAIfhaNzCGyvjoc58sLaTVAyNZM3tHoh1OH8hR2D5LD8H6NKvOY4/VFtw3PaOjN1
lq2IImYd3z/H+VeNoxQvTxKp0ZoTYhmzsxas1G1SVbysEk9ZROa8VKBbXKSjOOWg
o9otfRIVDCrL57RbakgbzFIeoe2JRkdnURUHEROOiaQ6AcvRV3wIEFWS2L3/vvKg
j4mKqBp9MZVHus4jfF9lsody97H4aXqnyLFHqRn4Wt5gqW1HVgO4ByrcUO1vShZR
U7boQqi7dMncoonhbvuqsfyU6Tqym1VmOjaQC08fYsB6d8EhUYlv9ozrKtX8WsRz
BSIxQ3x/nb7ahESY0tuaCtArHHSwMKfNMoM2vqZPC2/fBGpxAFWsFeiT/NrqLLBF
tDk0/tgwIhtTB+tgMqJryRFlJmD0S6Ig4AU0tiEwFOk2y0L4O5Uj1+3eJVCve5f0
eVZ9Ju9RiEXDhBB4yXFp6TNwPo1/fZKRO1gCUEYMvjMvxDc4lIsJc9bN1z9N8XRC
EKSRYFMlOgQF1x51UnPt9HY5NmSfFdCNkSYUDlvaoijrjSmgcGzuTAKqtifDN88e
If1nQWiSMj6TrFB/TUHq18sL90tWuYpmvRDc186p943y6Sa79afwWoiCu+7i9MCs
whVkL8ozn4zWCFO24gVp9oHKUBi0bFNQGYSvC5NJk/JOPF8vXIVQJm8ixkucMz7H
ZGSwtTXOHw0jGgmmohcmQqp+TEcbkHda5EW+BUXjzhJWoskZMrZs5tu6zZFOtZbL
TtnZJKoGintateoim39BdhYPVE+JXXgk45N6CxmkSbam3cLdYfg4CIglcF67Pw86
06Wi2Ff1cCFJuVfY6bOrPfImBhqbJJF0FKU1+9jtbGZCOuCEhCZFuSZXRY5TZurL
rLUwcT6OO/jizgEeWT3bI0jZVKXdhoToSKOK6TuJ9WE7EBQ6mygWVdHOe1GiLejq
qllY/QKA8Id0haucP5vaJcGXUbays+RkxYEDDsFY8W5iBercaRc6PzpOXzYeLXgD
gfSpJJWeOQ0MV7T17J+BVunLHfeUp2h7rwdMudGeIF5iFWngy9CJXFSlWWC5inEj
WvDj5076pmtoh8P8yTQ4eBgxsFlhQ8B+1n9i23DaUjeun1XDFBwJpsI0qMDyDPGc
2Bafp+6D+b9kKOgnkL40gly0yJKDEp/CKgrXUo4G905W3g2/72vfHcJEHIr1f000
104hln3QJJat7N9CpgPeeHkQu9VfTBxqYVI+gxMrxW0jcfeg9QhswF/TxhXxhVpz
hjIfEf/LvORnLDonhZDa9Zq1TCmbZQcsY+6jYeudstmRCfFjEAL1Oj+UXDLM4aX4
0eMPrn6mzw/XhpI3hUbcQH8ADrsGcNA75/ICC8Ad+qoJN8xTruLznG4aXOF70QUT
1sfd9SDTMwPA9SeZEX0dmNwnwnn1EQEr5yCdWfPHuDvhOC/8Xs3WFK4wJNkb7U4n
pDasCvaobQMm/1X8QawEwcmx4vq66TU5ry8ZaU38qJzFOzJOS5y4oJpdmKvmU73B
rJuTYS2s3gphyG2UihkgdGT3MSjpF2DJWLEcHkGyfpQ9jObGAMkQNjdNrJputVJb
DNhGsjNydw8le9zBlysVNGNqEgErppJaR05xazTuz+VkZdKwKcHQS+5MKwQtXoM2
PUVJdRhWMRrpPq9BDNSm4UovU9GqDiWpWxiyH2VDt0ZyI8w4a8k/UjieZxWzYIHL
JUmxiyVGbmerepbElpzQyE40nWRNy2h2GpahVHAdlBlWjHvLuek4dq19DxeSyLRm
hRRdlKu/39/Me9g1z6wJKTH+4E8cCoQNWtpr1bvYVSm+gfrMo3OTlOKSvQg5FFGm
n8r69aGuMmwZ5/8BWZyOa0t3JsDLYiu3PThfZ4OIsvGPqHjuzl12T4cU9fv5AkwT
dDZGR+nuR9SZseGo7m84D+sxG4xESM6UxVUPJzbQuCvTjQGhNvWunKQ4f9XzltFl
0JdM6bsZcPdNIdHGJCoPZeb4E1x98xYuqVHJ99k1pNARw8PCDN0Ih1/z1r7uGP1Z
PYHKBCmNqqjhlC0Xu9BxlFlMtxI7P6c3LbGo3d6SEJvRFEkt/n/xIgJoLSoSz902
WGfVnmYS9h+w9WN4DF9l9w1erqS/9GQfQzh5RLDQ+Nxb9wBYV9oOzhoEHw0/BvpW
Wj6F5Z33LNL7r4WVFlrOFi3yXzSJI6nuEWFjnX6UpwATlN2mA/paqyD2OiGcQ89E
XcaUNBTn5xqVNxw2o3E4R1bdkd02hun/QumEuzOEH4/aWI2WUtuHm180lBGSc0f1
TwY77s6UgCnXLdlvqN8ecu3hD89YPe0HDLzW9iKUOyNY4lIpNulNHUPYQV5PMcfN
6UeT5pyLop3AU4dY1/1PwM3wXnd73tMFzM8JLt9TIyp9y8qkjXIJTdWXRS4pzclA
zg75obJ7viVtQ3PJ2fh5xKPyUjODWoUs3tjKk8+W/8vSqNiyHj7Gngb9iVWYDlvl
2MkUTP+HXA7aiMBVvBZXRVkbF2J41lwEWl+8M5ZtZoixPa3tybdn0L6gK/ZPOh/G
nHHDUQi3rul3QPtdxB8LoviRg2hnN9Xcs0wnpD7NJ5ZzuPJUqhesrUbqQHdUYxXN
63TLR75PWzQBbxsQLcMvLJWetlqxl4E6HopxC+9OSli9vx07Fiw93VOFo/EvdXn4
idTrYCatVPRSsDKPhuYOZeGj0uKyQrfcHsAnm7yVIl1c9QeSqxMai2zRlOmQr8ob
+nEhQHZ5DoGiRNRNYNXx+POkeNg4NAkjSXYMpNqWISb6yYcYUvE5Lc2lwZg6BKWY
XgN+XVem09CdF63h8XLUROzqCLIBVbm8SqKy0r0Ycr2OgrjSVDugjNG701rW7DkU
8gQmQLOm8r4rBSsbmJA6Xaw7ZFLizTvQFp1EBdHzqUH48Nq4jVtZAEL2CPqvhHRj
qxvByv2VUxqTg3GzXbq0BzD9k2Ea3yGiS4H0PdYrr3M0smcAz49yE6p3bgnXyFl6
WnWapPD8qdV522uw6aq1eivTpl9VXrkfZfAz8DW6LufMy73spha7MGNMWLZ/4RSs
QldH2idZS16yUPtvA80DbuL4ruPeGS+OvqdPlxnNUR6QSS2VnMBA7PhA6jp9qkA/
25LMGUeBQLTuq6h+tSZW9dGtza9Eo8SEecmLJ+SD3fft+Hn2y9Kppk7P/klr4A5D
9TSPbchWa9uESLlDU/OlYjjZH/HxT3eaPo33CjeUH5qnZvog9V+3GS+xfgyAK4Sz
DQrvi7yEx2ay7fhCzXF5J8bTySO33OS+SsnHAr3oRHBbiQgNBSxJJ9H3Fyrq7JnM
52cqBfxJvouFhB0PE0eti2Sg0I41CpwgwL3CeJz+7aEJIq6rLz5k1CXIvabAzYn0
o0LGtjjTNbCpHtNrHOURIkpBXlXsJojJ0BouI7HbtDC0uzR0rrYlO2aeuEMKPX7T
NqCtxq2efYtBwz0KpedhU8S5wn0Jip84/RHATo1burrsL6BgSZkZN2T70A5/ubKX
UvljWly6pR+LstJFWTG5Qu0fx1pkpOVJJoiRmCJHb/o/psgEN/7vlsNmswXw9d+Z
B5MK7AbESvl9JSfvNeAJGaTFQt/mRvWN93y6QIWw8mI0dauxqdSBL+Dll+l9NGmj
FxEbY9/qw4v3w3V0l4qLxCGP6KsUZsxSoUIyN6n+F+Pp7y98rS+21EV+kzpxG1cs
ZTCFWWkC0jSyXjvtWOC5NUaW9vT3jBIlrDQta4IQIcLTR/Nv4tqMnKCsd1jum6SP
LKv14059XkwyQ22cvhD2ZJIrWJUFj4sn1s6XcZCDqfT3HnfWB70WrhJvDH3Ui++t
WKe4avrN5BFw5lL2qLbJA2VnNeoBHrHcom2PcFRElIsnG/AkE4mwywtWh3M51lUx
FuUx/P/y/OW5eFpd3FG/CbzBeQ4DSZYxgcGW6Jxu0X4Iz6aeX6RfG+iNsV8r+tz7
y3+qUl4rAL5/1foGV5agKyzhIuLxbCVlT1QlSxVxCKBh56rNcqX4QISow1oJC/hi
CzoiNbs5BP2C/u/Bug9OfeLOda2X43dhekhUzaw3X/2P9JHnuayf3bOkiKZpuNNZ
VnjiU0IiNyEifja7GMXJFtrNs2Y8zm4h35JU+diFjOMZ4zjaOxoRVt9mkVEFIgJY
Fm7Y4zKZaIO3GpeXP/CHfcglaNofzsiBaVMQ3bINrOVx8KRvhGwnVpcvhggMM90P
QAEsFG20gobls791MZpHtDaKV1IkSR233bbe8JKM4yq3XTbI2V9FSst9aquExg1j
0IOpyqmiUfNpqFZKacljhCFZsoNeIaWTHFnb0WWA9VGp/pw0bbElsyd1Vg6V6b6R
6RzwmdmfXLVIRPPAvlg7pkg6rOOni42E80t2cpyq0fDFlI6ZORYOKvO/rMc0AEGZ
LGfEZlUHoByraaLi8jCVo5PM4w9yM9X98Nwv4TQFixIFG2BpTbDnzxZ4/6mo7Cdl
p8JiiyyUYs0q4eR6Buq95ll3DNBy5KxyNsx1p6XJ0ClNLmxrR8YFzJLOU5MPbjNl
gOzFTaVt5Y1zMb7nhJjNZeNiPTiSW2Vy+oCWK34AWq53kAWprW9jN0aXieiRSN+S
cuQ9mk+kOdvLLU7ssMlkT5mufG6I6xB/6EK4q2tQBEOR2QDZeAI8/zvMX2Ym427+
8Tep2YefxXD8iM9axcGMi0KB/Ib9jUSlp4YuhhgXCX0uCtHiaajVbtGDpY5yOywe
8Zw0BYD3cKvuC7U6HfvF70149cCM0ZJZp1Q3Z3CJ7k5LdU+Ev/m5Lu113SRG4Khh
nqULyO+bv+sIldkMvIJPEgH2tL5ee8EvH9uCowpoeJ9JcMGTDJy3a0KELyilM+4g
ycZ1JaS/CzP9uvG5kpcgHeBShvsPlevndxEKC8TG8/cRdakbzvYMyA5fxRSDiAIx
8HjChStPE9NvRVMRoXwitZA4884aCH71ah2p29Edj8hIuWQ//SG+8yYpZ8qOIDJn
0riiSyYKhc13Z1ck8MIpBVB+vqesxsQgH7PSvUL2jTE7JeVxr/bYnv9ima/T1VMp
8YVHb5rD6vV+BpahiznUAVRCZnYJVO23fXvcn07XwePFMGvpcmc7+oNjA6vdtwfw
nlYoEXRM1RWlSHiZhcpYVAjCdnS0TVRw3E755gH5szQyO/X/HB1aF90hXbWnGJma
I1086BBZFQ+izpqmjSiQm9fhVPXXxon8gMCL9MOZOCeQNNjJKTfp0JPvtzvQ9/Mu
OKWZsSxUStu+YLfHIS1zr2zugSvrDGP/qB3KStBN54qTtULhFQ1qj69KOvyF2y/O
Ixd7kKXk01YjaMGZGbuJa1xSbh9hNQWlYcZPASU5R2/ka9oSWXXWHZkmyT3zk66W
3AqKebTR6IMt3ARN/tRmRqF1jg6nkrGd4/23Xkuo9z+4hR5BggvVsXZaRbAGvlKS
JXDXgrkjqyfc9uXZz0dRIeSu9tBNp2UUrOVG/GzifMnbTnOGWFAl8KZKhFlsLIT4
Ir8y3UwBI1/UMjB05ZB5sX0gM12Uzdwv66vQgfXm4qe1eXiLsoB4GU/7QB1I7v8y
PfujVLu8sgclKBxz6/AsR1o3+Psp/J5f2NSVU+khs6Z8fFZaR+aG6VcHsmVa3wsX
qHEnBGRDFingB06UlzbxOsYqXRDhJoOOZv3GE47fQMwy9cNGnvc06gEN5X7K6Jfx
mZZasZ1oH2mxeoTWBkRY0DPj/IHwWERiUJ/POKws7m+teHpJjlTlwr4mEqUXyPTq
Z3Q0CcZ/uikTnZUAtXxx6MdwpRLUTvAWsQpzOY+ZqbXWhttDGRRVMxJToXtQ5Kv6
wD0e7Ymv7/6zMq7wG1xZqYF/UczrDlUZucRJLz5TJ5Apad3QHTl7+ci0zJP1pJEv
5wwlebLuf6/KyQ7HgYst4Q8EB2YexQXyPPY0953RdEeCH2kHiQ5x5YaYbAgF4H0u
KJgjgS/fNa7Ml9o2Wef2EO2tOjiY32fT5bvU5VnqaMJ6Eidh/61WvdHo+qcAmTuy
X/MUVzSojuz7WJpCj9122ZuMjognkP9GLDIxr3/qMZf8Cd4zFGZhR7ZwCHtCa46t
dlPj1xfEFWbdgluVMvi9/felhufxRElUWEKeIrwQlOOIWUR7qHJM2hwReBsmlp1a
fpa0IxF9HyBhBHGT/SSJxBv1l/idoXnMmOrDP+mu+bq0EW+QNF99TKqAX77tuKH4
CDb9WHT8TJGmw+Gp2g+Skiv3UFcKYSKIUiC48ZmU2z235jR0q0vQTM48FitrCTKH
/Kg55xUtQ/BGi4D8G+GiiukcSDOXSYtom866a4xUW83Y2dtlAgEgCL2RkObykyN0
iH6vbeKCQtohOnmBwsHDBq4P4ch0TVxEmBxHKUJQULj702I4zT4cv0EX8Ip5z7Ea
HL1rv1bqHu/bvsBdJCN6reXeCwm4gK+fW59WlT4LQnHPp4kbCiuiiS/zHK+40ABp
8RKZnpxO8lneNLhxacU3/JZPeoYcBZagus8G/ABmfrW00Rfk65iCCHx5o1JtlmGY
NudEMusxp64QYUu/P39VDLo95IzYNSacnK01e6RLTfaLm4C2exNV/0NFYGNquuNa
D0H61Jx9QLbWYT6GpMqMIGSso3JjMLUMEGIgECCf55dktc3odmNJ4PN7uUQhf2c9
pirkvuGKN3vTjkkGdv4QC5d+reCCELA6HbBE81cXtLdLGm3OoQH5uY7PPbnc+1ae
zX4pG9WZbnVKgJxhR+K+BG8ipthyFuLWlOQ7/RsJJZA87Ga24UBxt5MalNz+vB3g
KiwEyltbSzyPwZRgQ+bailqqZ+j0ncH5aGGh7A7Sh5KZ9+LzVnsFePto5BgbtRg7
ha+tQA7GjNB83B7qfZb6FWXR5XWlgslNuLGJhm/RIux6vUeQaV8gCPZNGYXNMnd+
G9IqMtptx5Gxw8rLSLbO4LouzIuoxdtbBcJrSsUjnt5GFcR8tq1BLxi4b0rucW5N
2Y2wSTzC9GaQ25xzd1SEm//dDui+gIvCTSzjXVxDT4142D+WVr6IrEqf7H2TO+DZ
gEjJAdWl80ornGG1Fg3g9lFCvpVZJEKEcjDnuSFZowuqQSZoR46KjYtRXcgr6ICV
qIcd+oSLlBqOXZEMcNuRN/WB2AgjUBbglOJOGkFAy4HJUkikEzW+n/SFca+8etP3
egp409ZldrqkIXuQbVpxxgNPeTOJ6QIKU6OC4cut2bXnPwysIJlXG6a7NlS66Sso
ziQx0ta2rzbBV+AxPdU7TgyvvjxkdBZSwZk2c2RAREKs157yFeyzKoSbF2kCTQ2v
O8rF6tqVlXEjGlY9a2sVw7MI6MUN4StIMekq6rdXrgzUoR4eVCWVlLcal0XkO9lk
97qSpCPgcmCZ4IFX5gS2NWgu0Ulsl3NUCHLi+V1PBn0gV25JCWiwHaL/uDKrca5x
XlWUUwUOjdWopfuh/ISquJ5l63UaLseoI8mHAEaO5FFJ9aDlHlnbaim3+1iCLVbW
0WRRrrbuuhcpIL5Aq+Q0TV7zFcp3MeX6FHyNMeeMWap0tmgS3injYx8jlPMWLXb5
j9+WFreSpH7klGPUPD+q0bA5JQHfIn11no9+u11m4T2ZMHLC+USaOgcCwT6pDIkQ
ldhm7rYGhG/xFYdWy6v6NNP4YzU9K3eU/1gkB+DfryhjOpzZR2+SE/2LhXXohDnJ
T9O0eX3ppEVAa7wj1ItsElpP69s467mDxvrZHThsDNbxJpnA1gNwLdLdNvjgwVYr
cQ54EFAQrgXh+bkzavVZK4bH9CR0DSmrXmyJ0uTZBW/scE680mp0EvNbPHdQ2tjq
wP2rS4lLI/a4+bNBQ2dsar5cy+lNYLYXm6+3B7xS5ZmTqkHt0hk6d7ggqtUzmz93
z/egbYoEa7pgUqvdcgmr+w2YYdYsTVcjnjtJMwdNX5XApVGhD/cEMX4+rZMAeHx1
34NOim0ENghFfrNHahZv8n4roTXd0BS/9Azhe5wpkCdOeIJd/Dpw1fAoqVNRAsjW
tVRBVvge2z2Lvhm8Qjr7Y/SZso62O7k48hDUoeomahAKQLdGnC5xOFido8WXUsFy
+xEGQV3qQpkWeRqCN43/aWoCFECqQW2STwVGMLALuSk//CpcnUf1FOBfHWxsSUv8
ehC1REqFsZqFD3xKSvvimGN+Kv07FtDLpp4Yf2x98iCYa/Y5wZz7ZlDqM8mDlkH0
VEbcoMism8IsCbeZdmBkSLxZHYQ2ZxIkgvmhopKhgn455Kni8FEwLYNQf9ZEJYK2
yH2o4dvrBFdiD/mWzE9XVycjD6HrP5hiExktCMG9w3ptMLAwAWbo7X5DObPib6Kn
UjhNSizuKhkdDeKUG6tv2+CBPLrXVYiDfQYgtAawYKb/cFJiT9tl8FbWiaWuZu3m
QTyKLKDYxspjzTv7XTM5A3majP6TrAXUJqbMeQkM7xxgfHWjpZFbU9eUbbVf9zA0
VaLqHgxHw9USeXNNh1NXMDWvZTKo8TpxV6hDx2KTorZM+blo0wawR1ePMEJDHwat
mmCRxN7qFuQwK1EHymp4hXuKTHaq/7kkoXZQbUxgniuVB9rFHuxSev4ZpEBPYWjZ
eq1aKC92T0DrmEsg6sawgGsNOXg0LETrmMvMZPrhqBoIM2vFgLXS4cVNJALnV2j7
5dzuQgCGDg7lMmxIhS/IvPX7Gr9yBjVGHdo7vEkYAuRvOhKayY5YagDXZBu0ByDG
Tr7tvQVSzA0xPqbnyh9nDqogHCVWSeffqnMNFH4tHq1lGDS7lVj5YXoMg+3JPch5
6CzPLi+hUe62XK8RasKlM84b7z0CU5lA2UWddW/PfDpQPrp6dU55DQjGmVfULtcS
/Ia5UYhIMLpPp3vPxximtvhGucsRxgvkOAust1y5jwDScihZrj7UpxLZpGo3W0LG
pC+QUdjMlrtL4gZF3QWjlr26WXL27tXMTwAQp6Jgz3yubQghmYlIU7j6YZmLnrX/
BYIoO28BzVNTCx9Xaq4fJYwEMu/QI9w8lkDDfMmhK6Whidx10Q+u1K5S/IvlW/4T
7hb/HZ/fAHUF8EixFtVYWmTGpA/MVGnW+/LHPKuMWJ7HOWjBEINtC87aMTM6Tqix
DqUo8UlC6C5s7fFG1smx7R5/SfX3b5ZBIO6T4r2pbN0uvvdBPyBq1/UImWbu5Gs+
bVEnLOwlbK29tRDNCYrluZ/w0XXCrP77m4l34I/05+M3vUBgUeUlg830w4vAXFRl
80jstk5/jxZLjUt67XR+uU3mfkpC3BegoG0gqC0vv6VWzr4JCQ/IDAtKuSKRNZQD
6/4FlgIgrcvBJRrgq3iYYNhYWQ3Qb8/bTgBt67pbd7C58wIDY0mqkpsiFX3iacLM
gGFvE+Gco7UUBgtJqMWPeKJ44o7UBqUY2mX1QDla10d6T5ScAqUTNm/fOZxUF+An
5bOhX2usdyXoIT6wV1g4KTeSlqk8LwmdMofHJM+ViZ5cGAt8VC+GhDSDQ7WyosQb
sqg2O8gP+d8fSK+A1/2Mv68wC3/vzz9ha1YW7OCQW75I/YkkYFua3Q6QiFJb2KPz
/bW6UCwmYOerC69kpCW6HQJHF5O/i0F09wmQmSV5SAwq8AnQ1XF8NbkWqUsWW3yS
dls7ko7vUfe5liIfiQOAXQV0Z4UCcCyCm1oQKUgZkJgVP+Z6DaQkwNHzvenEzqRr
Oe8qPgy31CMIVzGI5g8QgHPujbN5JPe9cXVYLUAgn/GimlMLFSIH5erYi8Tkjpdm
4eimTMEUfJvD7A466yVI3KYnlZV26yvijXG18jE4WW4tIl6EVeJlj8fNciIZljvW
wqQ9hMfQjuPlv2Tn3f48zwmUIDnzl3sb9RuLN/nlCQZlKJGJIpJ8p0eO+PrI6wpO
qXdw4mZ71PbuI8zIoCv+LtF3Eq1UM9fgIIaZwnj73ShtcnCongW6rbWiL15Zm07Q
4fQ80X60gYKn7GLIbmkHEiQe5L0RSEBu4Vbhj0mWEWFw3Rn9/BSgsezT6OtqM8rL
moGyX2ADcSCYf1O2IFh2xoLsJKBh5DYKsBlSLwCU2tDesFAA3kyhh+l425D/UuCa
zykHeVS5WHw28HOyAnzs8eCfh5WwMnYyARD3g0LZgSsYi6QIp3RZsUlai4SSNi1N
17lD6gCyFrA+ki1hbLLaM3MApm68qdGORa/5+f8rmxCzbbjeSv6qc837RRF4O66/
diwIuJfywbwPwTsz8AiY97puAsIt9zxhAWmR7J3NY2sR+FXcDnyDJBUr4Zyo6Qch
Ws+AA7TPthoQ+pgFT/XRGom7DrjIvPJtebVVoxDLk/pz2k6mRnq73ruDYPO6fg9H
sL9k0Zh6FNDWFVMNYEhtP6VNZ4QVxppplZeaGEc0mWavH2RhLIguwQpdWGrXExHn
Ti2WOt9tuscoJROjoC8jV0EjQqlkM4647d1y0sC5kvDHgq6CeeZP+pWz3/E5rJYL
SZskk4WEgr/1+9Oml/pIV3OthgLC0q0cFeleNGhKvV+dHkR6Q40VtBLQATW8EbiZ
omKUf/6tdLNYoV+8osDqnMYoxnA9IBuI+PwHA9IcQ7Z6PtJI+OHNERhKrQJ5DYya
GUB76HL+7J5Zc6d7bMHLfbg3wXna9C2OQ3+N5c2DAiPplDJCbXqNzuZ9XPFlAkFP
dXkd7gOpV6k3VKA1/Maf9E+PNqdqDTnCvclnVrZ+2TqWrL7JMYfmdC3ttOnpa4hG
bjjJ3Ma7JSaERISdp0AWxrx6wtKIxXIOiDZN7OrkSTDO68gntPwKT4uyKgH/BIDj
2qJVoxUMctf4jh+cFPcqBhyRWovV0FeqkRfWXUgyArxJjvrhXB8F3PWFezODoPG1
pCStZPc2fjNB6UJlk/y5Ye6JBapsm8WoDvaFKF1lGnAvBNGqcVrOQgfeHbDQFuUq
AV1iFEAHI0YolORuqtGvdVgUTQBHI+v09q26sRGWjMMMBBmeFJUc8pUU3wYCmEmI
GaIZ3mZ3xtemG/mHQ40e7Ab/lxznLTzK5wFMXkect8ChZT8xTuyrD5idj+qQmSDq
GeoaNh01/0wCRHCB3fEa1pMZlPPhm3x8YGwT1zMqcdWOS7QMo4GX6XNUpZGFc3n5
7Rx2N1L7ezZv70CyiVud9KPxD7Ugm++gNj9MOqA7ARCQZAFnNwOVkAQ8ID1hwLfc
hO3ujF+TsgdiuVRCeypbwX7La77s3KZaZP0dmGU0AmoJxcxwUV3iqd32to5VFR8O
n6c7unkbIw5MfQodMK7jlIgyeHsV8LwtfjLFCS7VTChJHceibG780YiVMIA5Y9Wu
QCxGA6b4z9h94ANeZEti/CSKK6FTcYPw9DJfGyfglfw0jdH3XSuV/5Y3Hw/2zwfP
vqFEPs5Y9Y3Y4wG7+weq/JIhSsYDX6z9LBlvzFZF3rlqygm7u73LMMrRd1d3HwAI
xgkPsvLpEcMh0w0+MIZr9zSCU9E/8xvHTpjjcb5qHV5Htg3VOROczn3qf2GDF0xX
epxpLuMC+3ldZ35cwfySzMU2S63969yELXQmYhNKyRUj3gOWbACKtZ4FWe9v+Y9p
Gs1Isa9R7TmXTpBa7qngAZj6Sr1J0ejCaOaSESZ94rppoQJgjmwohfvae26D6JIa
vQu6JuX+kfK5dO+CMWeBMtGTj+ynFVYHr2dZwDd+Ud5sNzaRgycf5vWfIFP8VNT6
maGv+N5JNjGkfTlz22G2kw0lcvpndlRoJXK2CvA8ELLWE7VSY1e2EkZH7NPjSo7w
VwltHAX/H6HyG8Cawn990jDr27rgeuVfyOSBUXuQ9dFhT+ugP5sFBgkumTgTUuL9
n1WbG76dC/Raeck7SWdS+LsyRjSTdZ9l/xD7E1vNBw1uy2n13N37qtbgK07zQ+pT
YhCSxBVtaI41l8H6q71xzsr6oVcBfEb6iHPrv+3OvQx24zyCjDPUtmfw7W2jHCHz
K5gSfzsF/lyyVmcQa6I4h1F5vrAosRGZPghGeI/Ya7lg6YldJtiUlxp5mTIbAHFf
W4qZUAIbH1EKp5VN8Aojlcwk5ZsBjJPVPnGw6/XVIbCneLlNpdCowid5g+0Rka5/
SbILeIJnuYjTTnClZyMEG+kh3va7/3zQUEa6FaCnO7r7brKCZy3tw+/NU8FA5TEK
QrnSaFNnSU/GaiVFHjCXjP3u3syd79YYOM9ft9YqPnkhaukoFVDXl2Qb31LU2hdh
yJIozbfcOu/h5hoFEoq/EVLvslwZqs7rWjzdLJUncHntOflXgHpY50r7LBNTBXc/
xGihTF+B3p9km+s7nTWoNJsSQ6clWcOdp/swqI5DdJcchzGHVTruY/UEGwpVMEA2
wbdNLGGMmhFMGJf8/9wzy5x0/SsqaMPVkb3R9QghZANzWyEXg62MwJ5PbRz+M6jg
gYu6Z6sbiIAZeyTsN9tugakTKHn33COazZidz2V4zV2mryKdRABT36Jne7VkIxu0
j49P7nVoUYPhaNeQZu0BZYlUDptje1mc1WZW4LIEYXuxbDcR0hyFS5eqspgZR1Nm
VGApxRk+itke470Kx9axkI6bZJvKUtvasJgbiUR4hD7vbzAJ2ATVsC97ww3wHPMV
n817+/+w0pV/U4I5rNl9NBuh6y2JCWBO/nlHY7XQO92r2o97iZu1JiQxzyWsDAew
5XmehMXKoOrXuS0Te1Uef33Y5lTTa2v80uci5BlcNoNQwxCjNoZKgpmC0HL4I84m
DTKVn3xhIoki0qOn3bDCkg0g7c4IGNRYvaUUsd7UDuAavuWWANqtNtJtk1G5mAi9
1oWs1CWJg7OxZPNwNCCpkGzlO7Iey2mhc0uqR7RzhCJP6ErkBiXcMQlg9mabZMl7
g3+MQFrF/Qa6ZBEM79LunZPr6ivO7rzXCl+AmeZTCyOHPvzAZ9CoCLn2f4RAc5Fw
Gz5fzycAR5wX1G4WqR63hVvux7CLVn1ZHmAYCYVvctl7iF16HOa8Yy2wpbeYxMr8
bZ/V6SemRbpkdO9ghF98J1pHAaBceo1IWiVMvd8+YDMT/tt+owPXv+GPLupTV4HH
ptPP0fMf0/G3ozGyDh72Cx/5ixYXpD1IIzsx0bkC8MWPcyWNzV0Cxo0PQNPL8l4o
emublx+gsmTucR5k9mDxVM9moSAow/I3/6tuHAmLzEgsLrEfGrP0DRdgny4ejXgW
8ZQi1bqdCb6Fi5JL1W6MoBI3TOGkFhuIiaNYmKS7VxsBB80iieRFDkvG3hFQ2bVU
8j2EI630HTdghIADSpcxDj3QKrP1umglfF+egi+CoVnqponpigxQXHgw2cakzDd3
0077P1XMn7xGLEziozlMyxO/g5g4uFQMxu42EC3VYAbXQZ8OzxRYFEsRMrfD5bCg
dm87I217586RXUehDHaSFS4LdfwZgLxVuIrNEldHS/LHHw+RW9hCVoZUu1rj/Llc
zUn++/yBUXz0O2X433SA/tIaubde/25KJnX3dK7/ONL1aWj6S7Mfgf2UV18IenLy
xZvqK5XSbFWAA6vlrp3KhTxOZZLqVDCKnj15VvD/pGOvPJcfe3qTEJSxSa1dA5FI
eo05fdNaZN3Bve6tRjvdSjSolLTtc55M4GYrDxbF+jR9oT3OaFt7+rqIeXbRZgRd
lxSbidMbkqNLI5pZ1qnm25QhoiW2x7hLbAHZDbBSoMpSi8phNp0QqKTmqcf2eMQw
t3tPzLyg671yZuPiFbLr7TW2r8LK8zzAoI/c1QiEqlyVTR5sMYBZY1F7lyQ49l35
nm21ddXiVyp2bBqVpVxGFDpLstnEIM4LqbrtMwltO88KsZBluMxrVSQ16KPmgW7o
+S3n86RwjZJpjNSKfwXeDSX/NuwqMwUA8RyroskAeapBZ3e87Jf0whLGTakNHVSd
JmlbXfdXVCTdhZUZulypAHCqW2GCPSwa4Z8Kjz8t7u4hK54jr4c04Bv2crW8bO4N
JFmtjyrcKLVp9tjS+J1x5Zb87F1xJ+ZrQv+BnUgr9Xe1EDB/Se4Jq/k613TsDF1A
Ly6ukTsB508FIdJCsErDsR2kymtuLh501FNyfNhnFaW2/zmvZnAA3w9nbuKnTiER
EH/ESX3GsHMQEydtkvP+2iki0KZwk3/M2mkqxRi5br/9OU4fKnXlC4SoDFHECISm
YT+ON8QKFQiSKhFM1ixy3fwn8ZvQg/SyzAhAORLYbK1+/xHhPm4DoOwXN1mZzh3u
Nx8IdVJCrTdPbZPN4azVLgFnEJWzZlzpcPjjKVT2MTzxeh5yl3qcvANIlsotXuja
XU8UFBmsxYZM2lrgY/yk5ukcgud9CbneYByTmOHN/eIgWgtw03gO4RUX6aHLudQ/
NkfdNkF88KIIRrBiZk+P8OpjhXM7/MhVESfucgeUh4FD7JSnPMi6Q3lwOxVtyYzV
TrI1YBXJUKMelzfax3VcKrG7FZvjrHEASpFfAiuRNC+6xpquUTVdfG0mosKhwOfi
Klb5vHCW9vpi4gPPJqzkiz3MAj/FgLYw2QoHJDkemRlnT589w9nb6C/uDFOn3T6x
O6q14/+wZdnFjH2YyZ87pKXDHOW46wkckUKHnPzMppZLECXQH1XAdu+0mt0l8/SX
yYEM+Y0tUHYbEUOuutTJpLq/wAI1i8KHUG7CvcDrt9pV7H6zPbVq5Pw2FSye4T5J
qdohACrs9GNn5VH01lYpKcPBZAFVreAYQx/Xzorp2F8nvQIUUCidGqW9aj/SeTap
iylCD77pWdjDBxVg/3XbSIE9bdWZid1G78nq1xW7PbgxKqvK6Rqk6VIkOILaoC5h
WXr8kriKF5nMzVWVnuV8Dc/Z/TV4A/Oj5pxBv2xLupc4f1AKnrsjwb3SpMpVeQs+
t/IYv0SWFfgjVYja30PLIHH01HVP1BQmuQuIk258s/BI0/0UyLRXVIXRTx0RXE+X
Ep/01U58NQE0K4TIk3nk1OKTqoTmPkRDPEecZIyfoWgQMYdpgPbt6upHRp7VrLkA
7tw/zhuAyIGL35KdoMYWkXV+xRaMBtgkQ82k7wv7Dz7j1JYfCLdFGtu2Qfa/zq4X
7QsVJrVQu0jTLjSWEnWjUe98su8I9l5ncc9B19dHUH9YD4q34uGnUN5a2BtbESFZ
RHJH6JgkuAnGOOspO/yc625SMYefkYLX1OT5Gv21TmOFw2DIrIgTYh0uZ6CquqFT
3DTYisnJ+0ZXrlqBLgQoTwK4fThQHYG0bgmoRG6gMvONY1BRbw3oSQbfKfAUlC8m
GLQnx0vhHLbGtPvF0pXZS2uPicPVxmwLdyU7cIzQ1GpAPhyKxjKsaTGwVkpPIQqU
Nhu6INb+jeLMUUP84Kes8KzglERyNndFoa/eh98zbh2vFkSkQ8NG6tJfYGjSk+8p
fwgjozgVSJg8v4/TlBAddjEWDhFlGrUdfwOkmkWKc0zRKGQAAOmVP5l1uJ+fsAwT
tuQHKUtkBdZDhS/iJyDndWj30T99y6MVAoJSvvBsPTunuUEj5wohaRD2D6hpCj4p
v9BOj3lBBdNWtfAZMGtdL5bJhkpVPn7gTnuwqM5f8oMMCAB/OZctU/L/v09B8cSS
pUhoriURjYxoHMS1ew151kCVr8guKtS4J0Ht8mNsIz4lhpgtWJvunMlEHeoByc8d
B+JYcfx1GvkO86MvbW1EPuIaBp1tJciA9vlomShtHTM34iIYqIIl0ZYHF2xrCu6F
p96V0xQQiAJ/XlQiEPz4XpwrLn8ZndhfVLxptHhWPsW45MNOAr/EUjWSQSEKjmN2
WFkHq6ohXB3taVSyh0VdAZqmKARZUfBdyyC20KpTsCx2S7KmwX+cdof9hsevtV8X
JjW1RIqinF9ZzKSRVb1ayJh5Z6wyFW/6viXPSnt0evpOedR/7wDQo598egeYpQGW
5v525LzvFwhwXp+rcHp2D+2pJD0ULuXUCMq3sCdNjpU7H5YCxynzfZZ8BS3ZSqd6
Hy3lpRAc9+/bkvpV7iCxH2ED7D9um0LF/vmP5OVCaLyxiAry9a3BsEIQQwEZ/qse
DEsUbB7tE+uh7fwd9rbocC4EYP4osGzecDlUpI5ttRjdZN/DxutwfVMb7G8fyq2g
VsXZOZO/BhR9XVqbXSoOWQtEjIM2hzta5dbHxf8dWFHr2dvitR/ZBxC4zmxyaI3q
KFc4uE8LGdQAfEp/QHi570WUciEXM6UU6Ji0ptzyHWKpchDJgfp8EERWUMzChOJN
3SXhv31jcaCL56DaWQuPAFBigp5inDHm/QiVMEKsRWkd8lmS25grHVG+8DLz36CP
25su/kjfTB9fiAfvnfynFDZ599PR2dnmpJj/ebw1W4ZEZvvP/MsFt7SliGmmYn3e
EUcs5pkTuWpbaXRz3hSfWQoqP9Lqr8AaBSZ/IYF2Gwoemelp4OqFBPls7eVlgJZr
HISGQLBLLw5POBAZE4GYgkpp3KfgEY0Dj7G4DUkLG4sfbKd8m3OcYcLOix09k+Wm
XQES1X1Gvjo/ncd7bHTJMbddTCGZ4ZyX/h1aPz0EBhS6kIoUM1zVXO+3bfjmfgni
mruSzxjk/E1zLGytzEvUSjI0oC3S7U+FZ5GjrogalR8oGHEYRL0jFfuBXvLOdPqO
mYY/VJIFr77zN8hpMO3T7mVp3fuCo4N6QHjeTZNz5K32Avfg36SIN5GBnDj8uFOp
ZzH4HHceYJkCrc719mz44IQjLvxSikrP5EYT7CQhWf0tKFOnG1q5tUXX9pLGYFIr
GROOGtibiPKWc9gZ2lryRgNvkE2a60L8eBIV73OFQ7sSQ9Nk3xrejoIuuUF52+0G
d5aMqd8pwYqSnOUuWCnJ1Rp5Z7najzhOiDMkVzMrTd0mbSkZi8h/thDzlXjfMqV7
nTyZL6hAaKAHAl4sGVh56Y3Va97JpeTsOpAYVOJcDuEq/jA/FhOKbJvZHptWd3PH
/JJNuRPDxxbqP9Bm4VQKkWPF1C4Cp8toDFG+u8p28/NTfuqHEMCiTGCOZFc9L+5t
OxPnK4LKpq7Tfijoak0zt23i5C4S++XnqxdiiUuzRnfbxstIASmMYCWXlKN7x7cq
XGX0V9sUVOxT8K9l6hi1O58Q9qPn/bfReIF1rlG/AILGk/b0kHt/8Pfygud2PEnM
5Bd/zb0z/AGkCg+1ufG/ZSsf45Zkv+pPNVPHmlmQn69KHIhZ1TcKew7Ju9DzXGFW
6wSLutgpxnlqOFaWPLldWCee9dkmgOScAz84CxHqePHdUhmSYx0hUXIZwcsKql8y
3GO347+mWrNZSKgdFnx1V8tXK2c6wWxmHvZ5unBj4UhcFD9PDNdl3quEA1cJI90z
m+pxjoJs8VRingp/mFTsskS8ZLCAHaOojYQdfwWPpEIgVl+VDB216Y73F/Abomtj
z72ETravvi1ezsiQmaOQOHK5MYYkNtWX2RQXmT9C/j5SUrL0/kkPf0DaGt3Inrzk
6OUsDBq1doRQhLzEQzVQCBdlb8bgFfpmn9Uh0n19HlXncGOAGdWLN6nRfzCt7zUQ
dYwXffyoZr+f0aHnmA9+g46tdN70P5Qc+VV3Q6P22Z7u/ppzzBjgooZazk4hceyf
LGbD5piGtWZRmzpGnCozHn86CMhmeG1H6IZX3Ql68YTXubEAQQyjivjpTU9NJGmt
HUtF/hw1r6mO/Z8Mob4ES5hA0EI0elB2c5DtJvqKCNTbchA0OfnVMYD+cqVGsGG4
fTpc6D0jOe7HyC2nY5ALeskxmFCxV+bnSZvjEZTITYljd83K7kj+MFLRqjJJC+kV
U42DPCLRjqgNPN7kPhAXyAWcCOQj2p4GEqn2Esn/LuCtqKKvL7V4HF5DYNEcpRcj
YZa/4EtrkWTtC8aeowQXsp+Be3dGmkXI1xyRvYv4bCAtp67xrecWYAo/j/7gkaE6
3WNDTCrbWTUiXVYkFjYjG9u7Xk2i5MTuczCJSVFE64iJJqYAW6LR4xqkV4PtXdff
jXN3QomUJwQVbvKcqC4maqZq+iGOJL8F+2iWb2oe+XMYzb0tuhmhcxOeteKD1IvU
yv2mbQsmOfIyLRAUuL4zi5NDNmXdjIJX2J43vMQAI+/5YefitPB9D7SI8QkMkdG6
FLWzrHE1QicDH0mNCC4zrT3gd0YAVnjOpN+dYEqWQMWb887F2B+icQVPPDej9y2H
NCoHLp9h6LGkJH14BRc8o2d4Iy4LNuxL6p70tjNmyA2YukcIQ0up+QeLod1EvZwe
+fP0ionfGGlb4Rt/PZFXuHg6Q759Q1iKNAy10bxuBAgVIB61ne6brFL4pgBm+CG5
XlF2BjPVJx3e+Cpcsoj9dzZzdiAcuQBL6rKzlqZshyuJWgaV+Z0vl4eoN4V3Qyv6
nWRIp2MOwMO/HAWCqdyN1okfKitC43+pa1zcTubG2pi4kYtxbpBljePKQVn6lV7b
C8n2peI0xV4Da3Pn3s5A5B7/RJKINnAA/PY7gkeZsioZj6JZPx9BY1hb2+mJ0OOH
PQfb5nmycOhDA0jlSSa765SxtU5IhSjvfCHIIODqVUmqnQgzMU8CwZFxkJ6xB752
rpTIiYqIFKd/Fdno+UQbLIgguOdXy4ibB5WVLlUWYHM/Yda15xt7+kTRaIjDs+Ep
WePW927jqSLZssOPd4WWTu0MJbGc5cWQmM+/+LsTrTRgmoWP6YXjJT60+83NtTJw
rUjqARukXfDo9CZ9KoB0knltULt/F59r93Qu0gsCALGybnN3CJMq8yMwdDdpnkdT
5zChD6kJKldu4Toq4iDeFD1eyPLjkUHzzU8ZH0Q2Nvbh3G/pGxCNec+1HMzzU26i
fg3hwmqawpjM+rSBmNzV2l4H0ZYSb4DdY0F3/wFTdJPOXr4XuO4CJ6QGE2sYl7qb
teKIo7vGDr8nMgzaQiG+/Rlnilaj6lyJmO/Abn7CJbTtlV+9mQIeCNstNMlLI8KC
Be0LUV+fTqwG8mLZZrGtcFlSkTOWpi0Yocp9TikuPUilEvAtJxf/vx/T2W9HQxmx
snmFbm3e+qypcF84EcD47Ra4ysvmnBGHa9EPYRe9MYr7iUufc8mBShKZgnrjPkaL
CXBJrX5/zqDXuxChT8vi6gGt8JUb0wX3k0AU6R8J06KOZQmLSxnDjjsiVIGpIlvR
FmyLNvniWW9uZ1fde/2wjuev7GU+K81NapEwF2tP+Tf5tg4aFEbXMeCyYfyFszrh
USrghrf8O0NuDQms9vCMnzBvYAh9W0vZfz4YM1+XDHQKSMKoLBQUuITBrGoNJdlM
jrA+UZjvgTwDysJDnSN1a0BZ9gZPvv6fne2F50Mt/tmvKTVzcE3P/zz/T2Qjjabw
joD2C5pIePosUFxovkjCg+whTM/pfMZ7L7uc4oHbu3d50irUX7DpiQs9kS0Wlauy
tjc2sovbe1yqOI1kXqucPgBY18/UJqc56k9xXc2zEw40/f5TA/DqhO+XaGTwotTX
14evMSEc2gI8wLPcKHTtEJ+WMkxdQDaiQyEV+fJELjN3ev6/xkgdMQXN72gNedKA
dEhG8LuqmJfw8VRbJ68BoGxm4DvRza5uA/c34YtxsZbqJRHxodqsoKJdxO7I5akR
W3YD3+5rssjjc/uxrG9BHEy0DtJkimYzvDgMeHkVg1CDBdokh4S+NNhbboWe6KZl
hlmdtUnyB2l2/g3rBQDKTJteAjUrQVV4KWDBBdaK5H8BYFElbh7LqvdO13bUp7Co
KsgOC+MoOQXVdIE+ATe9/dXz/8jHyHvY6mvrzGcKwR2h7IKqqmfEo/rqtRmP6XNS
iKESG2XX2dPR0c/w3AfHVw/ezFsgR7ElDVgSYD65oAPfuCaxVAlBXcg03X2rfUkw
s0kfg1W9rxM1yZ+R30FsQAbzT2Cv1aBTwbeEfxmJhWEBOxZgKEsKniH+/5MLr0UY
ObeNSgO7UoAeDOW7jASG5OYWKLqJEbjaih55s4FFKd7cdfc2iOQGRiIEa5k0yBAR
nDpFvLqd0+otiXnbZ8uG8oatWL2+5eIH3UBnlt8UClPU75xKyzwbMqde3+ajDyde
kzQJkh5Dp09i0HLsKOh314+BlCDG7iCPq8SKDEfZjIMUp2uBM4XkvgNN61g7eq7z
SYB0zMFNlAd/qM3rH7x9dT/lcggkULGKKpyAXe2GBeZmQX+W9JqycrtTv8rHiI8b
RSeG7HHOZ7ZMcqixoe2ZAzVaZ0DkzyxQZii6GuhU8R4T8fvePACFXUeIiI14sx7u
/ZKmgPXNM8vDlZkkQmFC4217hiUGfhbhSeOO/ixgB2BsF6DPD6I9AO5WioJ3EifK
l8UIVLkpmjWpsiNwLN0FAMTeARJ9E5m05jAheQ8gtWSFkQwx0TnQxpJwcc1qflzJ
J/Ok4GJA5hJJ+ldb+09Dl/k/DdORunEROfDgbB7pj6arH8bUztcyn6+AfqF/2AQz
ZsrfEozipQO5LwHiWsBJpiMB784PA6sy8MARq2XAOr1kDbdhONmGvLOI6713hcWO
ccy2os+I7DirCy/xVMn/OhXUErejcyiPHgQmynUVajYx65DuqVc4ToZoIRUGjW7K
jc3HVjOU/oTUSNHHiifKh3rGujq8IPrhol3e54hU4TNSfHWpsnyB/G4KEzZdom8r
isrpxFNuA2JRKZ5IphR9xFZjzbVdSc5cwdIGajeSpUPgYtEAvxYkLE8+kFTIHqeg
T6O47mfhKuq/XGHdWpKT9XqwbPnEHCTQFOvr21VACmbJ63IE7sOXFT3tmiVMGNPE
QbcPDlcZjczcOAgjSVA5HVOmJsNNlU0Lb61oj9X1O9wk6l0sg6F4nIMm2bHqKyMV
Kc/KMoxYPbyODkMpvEvDtlE2rMC8Qp+F7zsNaBnJLL1nAATqNoIf8w0am/mOTPnO
oLrXYMvVFA4eDHBEfzqy3yEK/HRk+K9xp8pcAGQjYTg7a+ALh1TBOIbT2ToROojo
wq8X6MI79yQ2oyWNFMuRmyLpsvXtXQZxGYCHzz3FA8Ilbqcw08dE3ELW/LKEapSp
+3bVHiDatWoXDI3zmlMSHhc0QzZzjD3gxLDX2TVpbYhf12eQJ26M27g5yUc6wv1P
iJ/dIuXuChJTJHNKbAe/2wAregjPpJai2UZeRZgXE0Rpght075rTPmK310BF421e
am8DqFw7shxz3dipjyMsE9dx71Ai3b7ihbD0Qg5Ul+Us31gtXAC0EtGzAK4nlzth
phFKYovaqPxa/ItLSzIr+Mbdqz4L73RMTInZ340g3Z1MlUAQ84PVrETZH8gKkRXx
5coesf4H/Pq43bSSdHAKxSWKorknqwC04lX/+AfqnjrJVILc8iJNEXIvyqOO+4Ai
CxToLrHUEbLopEz0QSg9gFDvBEjzn89GYTdOjxAJCU4lIXhSCK1bvXba7MrBTfFx
bx2LYiH36tGmNazu9iDn1necJvw5MbYrXfaq8ZX7LiwVcAApgH+NeM91E7IW2lCM
g/4DkGeCDMvaOriqDx/VHHJk/hGibdDBMy9GODdnGvMaon+luAXOuq6SU7+8RdNA
IG4ICYW9hiuvs52YTVHBCm+/mzGNNX+WA8SjltrV8ZdJzs+NA6rgvrrvdp+Y3URP
T1v5nOqL7Eq+3AHJ6MSK27kfq41Jfz4AxgcnV/hEjBaFd5W+4pD/zIJ5NvCrhcFx
mONwdbFiINFd78OFyuDQ7mISlRo3tkO8Js5GQ9re8JM0vw/gNtYaqlJS8vQdt6VM
OtamPB9BHOs2pkp+EQWElgwS/4fzQk69QEPBU3dPL6R8t4GND94iL2qNgmCBrAfU
HQVQUQemfzQXL2e3ihsNDZLXXBF2JvJ+FsnFQ1UX6OGXVGsrrBhrpJye3GvUHvXo
o41Uw+7MlDCKXILZJbclWr1QgtQtl9+3NcdbWJixcE922WtUNrxOtx3X0Ik0b47w
U8XVPKlG7KLP2p/7y9OkHxICued4vuyv+CDANuMl8RS7mXVnfiI+JjU5u2s6UEC1
OVbu2I0se+hNTJ5MMJKKNJchsjUChTkx+zLj8usg2ydGftcw9EGDVNo0YzSgWBzJ
6HXXpF6x6N1iPLl04XoNK8+FPvlzYCiU7Q6EOAr07mvs+GSY4IrMiP1R3ngz/ql+
D7WU9P5lWb7i69ZNCxJZmEU6YU9VyN96m/QK+06x9AIGahd8ENhqlYgk1p8xo1bl
9IFpngAjtvtzxhHz53hJ6pTM41lkliVP/h5lqBRS2cFEEJ3U9A9MWhzPxiU2NX57
i+1PiKkpE05+pV7FxM7WfMPH0AfmflvHZc0WwoSIAjezk2wc0aEQ9i0EeEbrs4zx
nESEwW3WF/w7D6YVwJXQNtyGNWvD/nKZl4MLEyXleyJriEYma5TOZw3MzFPjH3v/
q0IjkAMgxMrWqMEXgTZ0jL4vwKEbnb2bYmlujxgeYmHVJY9OVYHKzYf7JIap9rl9
8ubrIbzrNv5iU9E1R0A6kolOJgU8zpiRksm6EV29jVyHXwsZ6GsU8ZIIAy+5lUrm
12OTHSq/eoPJ4ReQZ+uGWftFOV4kQLB8Lp2Jg+443KOyxldvF51D37oH0lqRhwlk
v+VZD3KwehKV+fUmZLNbyIGzc6feTshxwG018oKbc+vKvc4mS4OYZfOwqEjRmp8C
alUdPrda9u0hPQ3s3RlmwBo2+to+t+i18PfIqjDUKoF6rO133lBF/qu9BrZAgdxq
EOeRLNvzB7ErA4CpGh66VKun4p9j5ip6HO53fQ7x5BkODZGBCzWnyADuvyW/4T9n
zhBLwd7UDucQaZYbV2rM4U3kXw5C1y5VAHyDAPzaIIsL51YJJrYSulQ9YfyLnWIl
3Nj3+1+fjXPvK2eIZfhYz+bjJXeDy56j6inoX1zhmZHTCCsGkGwRP7WNTaDZFcpM
pJZGGKE0n4yyunh9eENfvtZZzK5xhauqsL4WarlIfC7q/rxpVlhB4gdvJEmLP9WE
Qr8QpbKNhi4BbwuRLnxwqJTF1gSwCJPb97nIsI1SAq7Bmh9NQmxlyUI3oWtFqQTL
+pGQ9hDSmLz5+7ORXU5qsSnGLPF4GkRLUgrrC0DYYEpZQBjqPXQ6lqoUqyIqcdBz
q3wS6QOmfuwa9NBD+gC2c17MSHLaRp1waQCBvjIBV+hQPoHvOAaRQXlBB823DgYU
ZMVqt07mp+URvtG11AN+KcNRgus9FcqbWeS7N/wj1JjVMy3MBdCrCi1H2bzwiXVS
J9s/RRCoWZIbMpGJIxWqw5EDneGoaXfBJtGkZXJEcNaaypHmnVNJOluZdCtq27pf
+lLFdf6z69f0LjVXgAhxYgnPaWKIlKdTtP/x4wa25Yn9bnXkdKjzos24xze0s6RO
lbPVbslpRExkZqqptwBM6spId33c6NBDKvisfUQ+jcmiOrbrDQSbrCtOCFvz0fpS
yiCSC+o9RUSDpyPvWy8YyTY8SQZ85JmWB33QAYIII1/ZRSPm+qWCyPhXXdbxWlxg
BXTB067qa0DHFVjbem9hT10xzv19tCOjvNxmA7sFrtNWxVbyNLIKOq33YGXlh4k5
BzNwjXX4fgyyHz9jzfdq/pUugHD9BBdxKTNX64lhoUxnbSZgMXSkBjrtqFU+bCxf
y7R/gMwP7hMdKXTBgPSczYUEcs35j76yVnE6Ul4KRU6PmD/wGe10/Fzqz3z5JeAQ
nndHVY+59afqOYMy9g966Cg1xfi62A3NYUT8weV7MrrRytmyxbiSpVoPP5NAi6iJ
i0riR60+2T0AvfDLPc42daZSYZ2JWMSL/aI5h+C9ljr8K7oBpYy8QOzhh8KksyN6
NJkXnGi1MxiLniSfU2goCKdQsj6Z+KhEX6O7/E1QodYsYZQIX9I5Zn/iw/qoIGDQ
Zjw08gH0q1FszRARQHIAuvckkIyxWiR+zrZUCAs/pOJNU0pmOrNtiyQdAiHpiVV7
HXIOjqn6Y4GRL8VIRvJodtZMHP4n61BD650agyWo5a9aHZ1CRIhrqBeSPyB6T5zY
MGAHLIiAcMe30mw9Py3MHWJxhcvK+ISIxAUk1EetW1CLlh6RzRpOFh8fI6ztGnoT
wnTre8QNYsaey/chtWs4Hk97hYIPJOogQiV88po/0DD0Ny/I7IYZQwyBEBoFbZBi
ziflYZZB9rPYiwX1bWa43Ei1YqeAJqBIP+0BfEEDHdYs9pdsA2Xr+4UN69s1iadL
OCa9CLDMduGhXHmg60XJzl2Ken9kAhZRI+p+2xzlz2fy2V0YAgx7/G7/b9auJfRC
QtgEWPBKeWKJHZGPVR0pORZ3QoHFg6jqrVt5GV01AaB+3CUHw4l9PFdjRqUQvMye
jE5uKiMmrcG1aRKkkYvJH2Hcc7jl8WfozupAx46bzeCyHhdsD4MisFZgePepak7E
qyfarKTOrjdHFcwpL/3yKZ91Efz+xpjTTpHlXe49p0pmDsgWI8K4auZ0xNexdc91
T1YhKCw60PVid2xo/pGBjzkeVmTGiunAoyAvPFD1atW61p/6HbIm/NjsYePXJyQy
iqeFUpKHdVRmrsQAPgrIklXveFYjrKNFws0SJrUZR6BrjWQnXsmIXIyflDAJZHr2
OV9invd5nwemO5Qx8ihDkztLOSn+cD6S60UTscHqcc2G7bBpRC5nfhJwTiSNK86o
1+rJBr8s36O8fhQC5frIdetrqhttMbn5ADcqf4SXlql5KNwcJD6DdRPcl3NTbkbO
cV+irBd/KN6MCMZqpWqMkTGx+8CbK270tpPiMNnqIXaPnPnUIzzk23IsimfKFj5p
fR/w0JMkLDzGOl1JUdBzcHBL47JB/oHLXvhC1NS0h/bo7xUpI4gevjCCpgdXDJlW
y8wikAmWnmHBIoCX6QyvFK+68mFOD/8h8pATs/eCv2ICaLU2PUV5K8Xyo/TRffRK
MGlQ2H/HpjHWXjVUdXRJ49OyMiVkmFgNPx26vJGdURBMDwJCtcPLkIzLXvg3dObc
4s51XybmWkGNcEta8lkfg9A/O8kXzlZCriSz8D+FP3V9hhQW9Aud1DiGH4wpk+ry
bad43tcoBt42gIpICzNdDKD/LYTf9tkB9I0ykUGUIp7/5Uk97nOneHjF8MKIU6op
bJGBiGdbOsNfidbUFS+ph0wc9CzYyhOz/X55DNgpUCNA2nBJy27U1BgBRG6qGf0W
grGi4A5WB/kOxQmYydagYgwiWPnJ/4E6Ku/0pV9AJC8zLQ7hluXQ+Qa97jab/F0z
7JC7IPEqgmQTXSUtwQzPv6+e1+VYYZgLinaM3cfwmUAe8ADUQelQ/rrL6GUXNt6i
Gz4SDDzGkOKYs/G4n+9XiDxb02BEaCf1YsZXWhZqJhCt4vK1iV4N6rwletnxXdxv
VSB/BwZ4qkmxjT8m8947ZgxlOBgEsPRkap4UftKJ5mb0FMZ/sJTatVTri+QpRVng
IeZikgQoGHvIxS16NyR03wxa27t+2U9AqUv7ryw9ngR9n6bqTVGMrW9Z7/bDwrdd
h/EBxa0pgooJZQ96zh8EBmqK/yf+646TbQwc65Ba7mk/ORwtOzat2hq5ESVqSbow
EacH2lO7jhU3pnADn432KacAQgeYl6asmir78I40q8ugaVkUwooHSpNnUlNn2pkJ
zHMT0zYUBvdKFRzri73k/eElj1deIQsghTaZFJqrhEBFYW/SzTTBfPSwmQOfx9my
r4ujTSubXZ/KiP1d8iSHyoJPzYu1Nenp34KzwoTrErMDH0OSNhlRVj4bc0N1eu43
h9yDxlTfY8M0VtCMMvgo+6LLcy3JWiJUeUHDIyRQqEintakhfY2viirThoHAe6+L
b/3KZQwjNBiyurVj05D50dk6Cm3LLAj3p/YzzGk5XHRP2A0pjQ+hC2YPpXffAgga
TNvtlxO5q033v2cF/3p9hXuysk+2Lfuq7C2CQ+sE7oZZwKGtPTY2brYXOzqXaUwL
9hKhQKiZUQMFnHcXAGszWnCtMwcMp3VnXSBDAL+nhTPKuC5W6e7p965szdZ7SMhp
ZLgq6fi9jjpBGCeOxDDlio2Hi2u+1VgJef9ML7u6QqJwvGxJIC1TPNxUeLk/DH0q
Gj8oDnXqYW/zOnSI642tkPFtS1HLB+vdwsBNv9BYDIRvPC0jBI0IIPWzXGO1CKC6
ZjX7kJiNzpZ8sZwD96UtYEE9dwNks1ts9n1Gjti5JNPv0BfPXpdrn7PByoan1Avt
bq7MaiHL0dS7x5qMZjBttdWwpGsh9sQgnhOREj20aRsT6QdM02WbLjWOX+uJvb+G
UXU17uY9j+kePoFxQFFMDJiVmW+Ih2TAdD/STXPagZub1k0TJAer7pSYF604mF/0
tuxGHEPOpdZ6kr6fm3twQulwRSlBfep7OLVM8qNpHQyYz/1G4tFF5lXgT1kFEtjf
iVu5LqSvxxk7cAl6FGQON2hf1O77BKSatwlQ3+EUHNthqrReDDYjXWW8GvrRnyoi
G8ZImWmo1Jexaumjb501Pblwh37ydTAW6g2DCnvI0fwBE5EiAZxhZAf/aRgsjWb2
eO4GdqTzDpzxJseGQjUoHTDeW+BqSctwMFmLDh2Z+a3WWqm3DYe29AhGGiMI9hcZ
ivHn8/JzzZ3ihaardw3iW9YEsmezJb0zexqlZqxtJBPAjaCHmc6PS2xe94BBfMx2
gJtgqMOGJc5LEDSyGgSv6kxW7IAPmZFhMBkQHLs46H12zoBfIuEWKsGpRGVrMfr5
WHLUTsxLWPqHa/+BZLhzH7nZzxsQ+rf1VBuXAUnXV+Rij3RKxxR0zseImZ1XzON6
oS0ZBLnCX5JlZ1NbatZmM/lXr+qatvmhI5+DkD8RzLh74iE2LE2RvyQi8TmAHAre
It5W+W0Gc3Ez7iKycApZt2AMuDzPL8j5gWpMJ5kYWsqB0KlWg2a++jJAnO2OMsCi
yFzW59DgRjH8oIHCRytuaOdpvV1PRR156rQvsa/k9vHgu5tTkjGepeF4jgtVI02G
RWfyqLn0qDTI3vDxfcda38aoe3+IB6lbXFCnHjNSsZ9c6M+NdwoWoChBz3i5raku
7LcHuQJFG+85VWtQq0a17ExkVfXGiv+Q/OVG6RCwBoeMMt+QtD5wS1WoE6Ckhzc9
OPI3TSfYVJi3zwAt8t6wN60SCqtXDTbYYugtVv48/c+eqGszF3a4XBWHLtEGo5XC
y0uHjENtZNu9LqflR0aEwxg1DoBMORgDpqES/G+SyvsIN5h8OUb6oh4n7ULKnSnc
0hyxKE55hatzLF2RrOYStnbvJ/SupzjXtZ3c9CONy/Hg5dbGeuqbpZe9mYxkB6s0
3+V+UcRkWbCw2HcACfHAxqtBD7LwwFXFFE8aVF0ZiffFeOI93tYRcR/Q243srG1G
f2YdNHR2rfLAih5LPwQoBb+eNGAow99e8DzE5WBk9lP4CSVV1cd82vXr9NmBmrqt
3mdExhmd2ZQ0j/1fVtbzYbtg7orwtlAJro2qdfopKAK+34ihpuTkS+HQEBGUI/08
GzUvha6H651hsEplhpHJGqpjjAPMY4SnrDBWY0Pdn7tApxiCVtkH8ANWJUFbY0Eb
dhgOTzEFQ8fLlIIcX7e3N8Tjt3wV+8og/MTi9qhkn8FPUCvLCRnRhMlkSN0U7Qkq
d1tq1T2tOcUnFnOi7OTbqzRHADSt4ZUSC2dJwb4VxGpV5PA0iQdGEbTtkQ0d1qJU
DHFMljvMxfpMXQLs45HAx1FZSzXTPnxv57DKGiSMf1Ee90cpjKCZdpdRVg7fDKXr
RRaYzG1lPSc+sKMpLZuXyxiBLnepBVxmYCey5uUi4x2wrxBymaeMAnE87JX7q7bw
ar7CHiAQNymOd8nGeFeamQX5NYidC3rYWo2IvU+M4qErEBDBMRs1OULDpmBG7sK/
/ZId114Z2oTUnqA5bahQFyDYI9I3xAZCH1MZ/YJNQf6NYl/Us3gL6I7QIuyotCeQ
1PExSWsowgZlJv/gh9zV2HDRYF9eEcHKEh/JcZfKxvRCMhSqrRx0gZRXUAagGwzV
t9Aq8WwtHu9nXafoQEY4ahn5lATiQGJW+rcjiEbxnzZb7p/r9+3Hg6tITFXwgFkw
Nakp2ZMFOFKOhO0jxrQcf0O7OTcr/YzQwi9rhaW50ws0MNZ4ksvwAJYfb+UD5OBZ
7Jk8tse6Uw/j0lQIRlsKt7t6oNEnopZCOqTZbFlaNfKS6DSkspXcSJoVg+xWngz7
QxXyu8ONaCCE08jetm9tHOqbS46BuvX/XtU2wk1ylyLRg4iLgYSb/ekyWw167fuQ
4sFo8Bed60q3iapP+YwpfSdvikrNQJq2PYJ3vtuVOqyA0et/1Jp445/wbUjsUyfh
sVCT8fRbwtzpBl17SJV7er7BfWMPyEhEbiuv4+cHssGoTqoLrPopWreQQ+CFYDEY
8kUzyp8MR4TcE8Ra2KoArVhk+I7E0iY4D78Quz08sL0GIGa6MpEa1dJ10qSwTQeW
Di/R6Z9L8omUnHL/RbctWheHeYXjcuF1JAqQoGQtEEUwdFSLFo5ZGoAGIiL3eMEF
hjo+3STO0nsky2MZTBByEaVcKmRKmTmT2JiezBSHzfS9cwDLzsMAip2OI4241x3A
mxp9suBzVNZ5KfhAvXa1qvnIo4FBAbWKsoKJTbp2J5TOjZsuIE9cIKOFu0poboMF
jCiX7x0FOBRUMyYUMu9CbKPkoWzrIJUM71R1TMgAD+ExlhV9F883WR4ZrwmB2XVj
nrHJHwd1WCKvrwYS3cRELaZCRHQ5S43QLG0sLwiFBW7Kb/ZhLzlhnomqaUSSMXcx
OVOtDl/PW4Zr/jhbCEvKJguzrVftBGRoJIeHy2vaXMk8bQelAe2LWAaYZaNAWSiI
r9he3JdQSHJosGye7j6UH6zs6v8rfHZk6iVmpJKWZ4Ab0itSa1sqpvhGtt4hMgiQ
6Ss+x9GretjPw+LDVI1Fk3guF19bJkc/L1sQIMYMXXUEs2oOdteqpp2RD8e7LDOe
8H5xw167DWO3zxa/zj6tWCHQXjTsHZqH6zgT1HCDvMA2mc5zKwX3ivDCYJwjf7xH
2jEVs6pAUX4Q1IhFGow9LEOZMXtSP40PyJyJWXdShkLZc+7s+nPaqaqQys8+cZPg
Jz1dIfp8t/i9gMMfzyGV4ZrFDaQTy4+n8w3YBjStBL3KU6MV0dgvyfi1X6FPg5wX
/jEeT9qyovz3OWDb2YrKcSU7q/roOEbqxUzchkRql6ImevDXboERwIkkjpofvbOe
kC4KcxfDIoe4QOjFPcqLbGBSzhaW8y5cWN4MHDmRVhorXy+nZ1ZbgIuL7Ngmiy3x
E1DlMV3ExcWNzHnc9hKWkZsk9ZBJ5ZJxcOEroS9gYfsvUMC4WeCQnYwBgI3Ge4kF
QULXk6B7HOgCkn/gZyPr3N3vBkw4swIn3+kOFdInkIbzDqYdL9rDNFcsnsxtOk0y
eo5lxb76BIj4yzNilEq/d8bUPv387duwm5H/0phPrvdwqeRm1QWGCwzvN3tef8oy
UvOj3++2A86gBY83AZRfj3kqt0KTa8G98QRoTGW9GH/zb2bY/XzFSXJNCJn/Ov7O
kh4HKAkGARkRLoE5AQZHPGEBw+qmEtrcVdJCZrJ9bjtHOdew+R01ZGuBzJjhUuWa
BolE59HHIWnm2++bDtzPmYAeqlZdZkWeZMGzirC4zOP9EYI/BgVt03g7w6HUEXat
Pw6IQ+KitNZsHtWb1GjbcitsioxXYrlPrLuB9LA0pe0hyxUzd42MCQU/PT1vGAQP
88uYiV9twmo9ONxDmqATZPhX2gRjnkhiput+/u0ZzuTYU0+0iFAAZ4YC/QA2342V
jIIYGYE9Z3ZWqAHEy/q8g95RSsWmhOSL2IsngmWmJKNSQ54aL5ItFZZn05aBlZ70
pjb0crFMl5F9E/06Lyo9p5VEfr+Zc3BC2olLuh9QIgSFPscIKZ3LxfPDAWdUL4ST
EbXOD6x2LvhLNyAHnY4jke0zlSd+LkeYc4LmLq2XFRb97x54hWgoWK+4YAR9GjAi
k+31gFqbvpS0lWDi8w850W/dxayMc3YnzBOss/RID8RXSBmSh+MfTOk+Qw3lX7G/
mFbIn7u5inDA3K5xMa88+q2JLmGEhMPhszCYS/YpSheP8sWlcxJ3ytq/lBjjWo+K
79J7ZMAl9/Xy492/XS7zE9Q7vdp9D2YVJqSwCzKdOVo0V70UlT8h4eRItbR2kvaU
1hgYbxPTl5akaYTN+zMMhLKlYtVL1QMC6FlE491lLtIMf4QY93Tyyi7+vNmZ1kaa
r3Ljrgbw8KNpfZUUqlSsVWeGxCXkQSGCppGtykBO0hR8dE+J4Cvo56et5agXWyFt
w3XQ3jAiGIztuBIWb+dhsqmct2UWQJKjSyzPK5eV8Rylg0fK38n9T7MWv4rwf0ru
sfu+k5hbaA+7Q2nKSwTpXv4ZU3JqYm7LflCUEpPRCwak1I9uJ55fvEYrjqSobZXY
jPhUYFZPVxl71QpXVSE+Lr+Xo5bd6SFbSWG87MJiIV11xZ6AyimnWERYx8VU7CU7
PCkUtHaxHgAFqVyL1B5nyYGcxZekSsknyRpt3PMWBWe1zQp+WAXC6/uCnNrhpLoJ
EBkO1h3DSxv/m/4yvCKqRJVwRhbDwibjisaVvRL17XHPgIb9J0i3JI4ClLJk18WM
2YVNvqvpBpCEHsrdPcmbPRNV9SHrjPJa52TZtCniu+fRROoN0g89B0MUMrBn3NI6
1+YRSalXl/gKALSVjWWjhFTNRcLv8Pf1KrroU8v+EyFeOZ8/gOdYvBQ8wDHDmpdI
AUffX7MlC9Yn9xbqqTi1V6f9mtsWKeof9o51I/GUUFUCPvB0BMzh1ywxJehqXSH/
KLBHQ0jkgnOqFmhM6zKxFHlo4tJues8KA6kUs7L4Gng2zRJcdu6aDMtoABSvi0Ag
wAr8jiW49LZ1hIJ3OTHCQA5X9Hu1YV2IHJss9MHBuqtXqgv1NDw/QRmVgvK2gAVA
wilRzpDO3zOAwGHqHmiST9ItwyTjktmi13WA5HHU4M/jFfpZHLCpuylD3cYo87pX
x/dFVpCYfScZNZMk07OInPOZGmSEa7rXU0Opg/Lp4tf1uYzyFh5iiCcpgT2Q25qG
snUinrSbFCKMtLbBonZgD69w3F5Ct6A7gZCJ5jRPh+dxLVAxyRPzBGY0FvtFRv86
SxhQzDVQuxwibNWahy5DOEJ+rYwSLgzBnoCjPiPane6DLvRCuRGrbxR/06II034X
h77WVE3l6NDvh15UHUuwvpFw7gIuhIHH74JVnfZl7tn+duYVDbWyiaSnzR1eVvni
PbyqNOH9e6UxVhfexxkGE/vdrZAs0TZf8lnECbpzqbDyDyRuVzRSQkb0lzIqKic3
jtyKbBzCf/ELRq7qjZ3aAjoan1MABHETldbJZf1dOZWS7sY66sq7oFpjpf7a8+V7
PwwMTs6smPZ+OMVzT0fZ96L5Q77ZEUXLLQaDflIjjMVWKTIwdiTwt0fQmmLWUWsq
099Pcx7MtClPtbDfgKBXqIH6VAyswaZcB/gzsF7wHt4Oh1TYIFG9STr+/9QdWaRb
dXts+eY70s30N627HbuK6N/sPR6hkqtu2+908zrN7pY8KT8WYMxsQGXmd11RfN6V
bGn+tbUZLbkmjww/aBVLWTsQlKaCjlioDpBNeYmFjGkSybC2xdYXj/UC0ReOzBaB
D8kSeH33uUmg9jbdfcdpUekZNNRXT3t6dMCxEGfmE9vuN7Fdk6n3heHfe4dw/Dw7
fx7nbYImh1VT0L17pnQJ2cYtZkxzCqPMcum5ky/Vj3eA18W9/7jfBPJy89VPaYvo
/AY1uc5meja09WHN85iPjxNvQ6PlAPjxJMuNRmoIAnKfsxVn6QtEt/ZQXmD7+CIJ
45txIUBltkVmS+ARpxtTE40xMYrBfaGLmzvs5kFCRJHF+KwGHGggGLTXR0nzXVRD
tS6OJq8H6lAVdG/C6M4uO2WFUnn67Gsi0ILcRXavQaS/DOPjdZa2Gm4bbhrmwjx2
8K5jwyRdovk8fFNL4dHwsfXMcPoKQg+x9yl3ZquT5U349+RTTdYshBByZ03uNOGc
8/zkrTUuSJhyR8oCJeu/HWMVkCZrOzdFVm2yiDyPXp9VjDwut9h/llcTN01YeHpw
JtBs0VrmV/Kob1/GlmARGP5Z8eZgyhpvRNyyTswczy2r1hy6WCe3lYmndgmaSz4B
topasWpRA8ug5QN9BOuffbrbofi9FF9wMx+lelVKvyRABclcmHjM4mriLmtwVOwn
NTCNqltBfxwskJvT5zrgS7lLykHn20Rdu0QyPtix+cgN0EnosudH5JVH9md09FCP
5wX0tNGiyjPkUkF7VpwqvhPLMLD+qkmTvnrl1zLDICl4F6VJ0QVt7/tz6JYYqUGF
a9bfBqnnB9w2HRw7u7nvvcd9YQPTB7UyzIQfBPsSUlz/RL5kVghNTYhKafqr4W2U
Xiz/ACLEMt5klGb8trkMvQ1Xm1r82ViV+QHeSWEX5Yis6Q5xTQYAUEIqz8U7clGV
Jx4GUwl5/WZa1TelRrmOkP81MevgZkzFk9kdtbFfqbJ/uJ7H0sDbW8ZqNr4cavlm
xZouuW6Gvagx06RvXpVH18Yo4tikVBEBM7InyB7KhTI8U3MmhobpXj8SF04D50xf
9RVLH1WUT+w37VzL3+nYvkxRXCBTAcD7HLMXHs3vQNMBKwtG4/JFFECJ+nL9uEuq
T8YulwhA6Gwr43cTq8tTGq43HOwvw19mMYtgd12hjGZMeprgXxN/lQ1UNikNKLN/
Movozu7B5sFQQdyg0V65op4Rr8xkBhppymjeMtWPlyUlxBPAYtKPP8M7YokFwIcK
jRy8pV+yXqjYWGx3tuaiKtRMCOLC/27xAjDS6/J43Ism8yA1M3NxQadzTkEDsYra
uTFPGDvj/+B43mpykoiH7V3wokmnnhsRB+3CRPLmg734A+5N+PCWefLNXtRy7QpJ
9915knNA9hFYsGFx74gyEe7/abFTB4Zt42NVDzZ43tGZb67H2CunPf09S9vwNr+J
dTVdu52+6QuH8b5NEL2Frgvz9VYhM4JlFG1MVw9nWL6rZlZgBiga9n0hT8dgPeg2
oPWt4Yf3vPXR1jrykZXYNUDjHXwKQVyITv6t4qJTXyWkkQXYhLgCPrZA9yFT8DnT
sUxgD3pfYoBcx5zM3zvDewt1Ch4w70EL/KMVWAsyjfTf/7u1vGfj/CBHmPHEj/Kd
qrPTuoPCxiF8S3/Iz+0kfh/Ap9n1cAd1YCqZ8oi6wpwUaGc6Jfl8pFGCVAEu9eZq
+rS7FnabevIAqaFYLI4s6D+2PK5ODRyN7m5nXuXaZ0nyVDn1TSAGjSFkfausHnQx
WN0GXsj53OAITJjrN0YAyOwq3giO/pKjFTQQH2F9yKcfN5p8X3xqLvmpdzconq/E
SPiLh//wvWv107R5/06FTmEW/7L7ghfCkanSxGewQHJfoIbsSPLTD2500Pz6SarS
oFc8wYMlNXYpcXjSZrpHjIm6jBL6VC2MmBeRNWKZ6auUsVrUkbjWWepc0wSW6pdH
yXmz7fvodO7rsb8C8oSrYkPVUK+7lnyO2XqPhz/VCusFyoDgsut+DcwJrejv5Uwv
xQOQBW05wGfAKZQWcvngK/ktyrHDCwGwA6gdnSaoIM6KWXkOF47Tp9kEuICJr1aP
ZvnQSEpvEN/SjRrMvBkKXH3FT0K00PHpdPFA4St+og2JalXuy7nHXBEAAm/zyBXU
cZczVVW8/dilWj8WjMe0oa66dKVv1QNFjlLgkp+0atWPfLqDL8ho/DYYM1KlHKBQ
JbIRy9+z6L+AKKiCQbZusZU6So0BcZnMmiSLrYY9EoJb6vM6Egr6X8jvCnfAeZgY
26vM/Zp2B3qKHlIqAGWOvl94c2KRxZ3wJ5Gczd+CQ/fVM6JX2cBMRQLidv9cf3NO
mQDcosFrtc5/O1ES0QL7igSslQdzBT+NsIzMTxuuY67q25LS6u73JIzpUGsXTXvF
7A7xSw13yjhbJG5eWCCTM5SwLPxdLOt98oqg0CDXCwlxfSwFSlN4Hg7rb+05/UE9
M4Eor5LLQdhGMGFV1EulaOgOErf75CTv4ePEPpdRqgyV6Zgn8JG0rl6X+GMPxEqD
EPIODarkCwqCs0osND0l1g+0/tKTiuIES9RKCSjTIxNA87+fjwDwglNzBuC9A9g/
OAdJSWxOWp/97zs4zkfazNUxZcqWonaTyD9AGCX1pKBXxhGUFq/qoxr9bfCT80K5
P1auRQUC9P2fi1zs/pYQdOQ0Qnqvk5Vf4F6S9sHt81VYhx8TwTw/TcRbabdHb0Gb
y9WpDN9XdbEEgZe8FHBp/FQRjVOh75NNqyBNXuYpms9VqWaBFGUi7Yx365lsuCJL
9vySf7CTaxOtQxK2msa9SsbnUDQU8yn5qvrG78UsGJ/mRgyc02h58hS3ugZWT70C
JPL8y/ID1W4XIWlzBb0+dO6A8vkap+3lfIpXgrTfPr2OuPvYh4vXenlvanyKP94E
9IDj+6mgT1yAv77If6Ad2qFvyOCI5OwN1iCV1NBV0DU/K+mYDidN1pjMoTK0ShRQ
ztLMU0+kog1cvjBtky/OS6/COsKZyVfCATfHpNGUnoWH2PC4Vge0xYLCpa4bSqth
sZocvN7TqlHSW/qgXIyK+tU1Q3xTL4m4G4K50Sv/s51X0ZJ6hd+zeVNHz6H0M8+V
e0ggRJfb7j1fgv/cg7Fjqje62apq4GuGjIIngUe62/XGghuEjKPSTlCZRJsprOQh
lS0Cyw+9gyhtbkhQ5WjP1RU+dqprxNnjdSRolZNR0oREaNmZc+kQdz+JpkQFbpCM
J/C+Esm39H+DqobahAS90HBvFg1s8RPlqG064pxTBFD3ihWb32hWNqhKPOCUf6Bv
UkXbLS0IuVvdT3S9RLJqFpJeUPfOc7hx3gFPYak6GzA84aKYE5W47ylkFZCB9eq7
0r8DYHHICz1zEGSUEivA9o5ZAojcovWgZRWSsvVXhlNwG7uaN90BIKlEo5pM95VR
/80hpiiLHnBS6S1jzcw8vXJrfKtuBfr4nC96inCQJEjU2HX1oolDp2+IXBnFSf7Q
BC6Q89DYKt30wKMEoKWYTdnBkqeOnyTyl3Ygy3Qg/o+LNQSJDV+Innza3PfdfXv2
HmevbMkc9NRwf03k59mhITPsSyjA1br71/rEK9dM0f9dby6p665f2MP5TuVu/ksQ
rLTmYJHq7rfU9l+0fxEn6ThFGAr0DkxS+uttPb/Lg/54lWI0Cfxg3migSvAFuXgi
rvepsIVfMJYzuxszeTKg0X0zJhJucnUnlvxcwYU2evGENUd+2xl5WDIkNrLTSepN
lGhnCMPK3ykxe0SU3WEIbVomBUa7DZhT1yIMMl4YiBR3T1XfpiW7r4jcGDHYMjzd
rqftAmE+PSSTRJwkbAdQbGwDX9jDw50HOWmc6a6DaSEJgKbgK99+pzBuvmg1/n+I
i1h7pmxrCg0enHfbkjkjgTncLNqOTO50yONRDET/EV0rROtORoW4cUYr7aNsQYzj
d+cCut9BTO+AL8y7jJz9sTEE+8LS9woUFjrjJ6eAvNUK7WkelVw4WcqqJuL3rjA8
tqyEjqd+uTF4t4JMonZnw3FDMe7sTuPUMxQDUhDEX0cyglEsMRGG+IDtXJNHdB4o
+ABOxum8UYkeDzkdkyfXGCZKqe6zxzNC3UomzYXaAvUboqDWoibcWH2cLLwFBhKE
efHLvo8jUfpuFyVEFCe6WnY5pUbjXKX3hFHIXRkmrxhFAhprbVFHwvEHDjx0UTD3
h5y+J0VN1g+TPw8mGI2QBx0EjAsoMhAC48f28ZDC3ylBxA57dha5VhDjBqaRWaLE
dZj7RZzCPH/m7DY69p0Q8DkcO4H/pUOl2Iwx0oCEG33Ozh6BfMajg/Rgf7a2EJYb
EpbrW+quRq2EtbnoAAMEZl8tNXZZKHEyIN+wM49onVQP+a0iGSmA/rVOW4M3hXLF
9lS36Yvsl1rp8mrEPbLRmMdYEMq0UUTsnqT+SW8LSeS3+H0NVYbaxlWlIZqBa4VX
/ba1CapDNdOQEOLlbbclcmohOuqGmcSiumSYYwAastRXEWN6big2MnofAvxDR6x8
VkoCJO/I3UvKyGxrWqlMrSrnPlT5Gql1WPGVDtBI/PSikYDOZASp1OhYBjitEI3f
Pf6ghV8/nL4uXbvNjcPLXoDkbzxyg+mbtsa9g8+0JLkoagDuFG09DAu4Bf2CBN5i
o/e+CvLfQbBhgIgYsit3ThFqz2bhIkugkwRx7dAAQ/i6vyhHSxV9TGkYP0+Gc6li
SetHBuZnxb8iE8nd5rnk2iqsaGUcn7MoZDFFqoqp9Trbwxs5orPIOSvUCWBufS+D
dEyjiJo+7pNzrlTNJPt+gZefKBOOXyHHyKezbHX7wVeosQWJR0jXDOO/3ZgITfXk
Dd9T+KPJdJvkGhMiwgI0NS/mS+PSGAu+37FDbs+/py/4BSA7uGz5kklj6AhVSYq1
iGQzgj2WeDL3CKb+cXRLpb9x7A3bKDTiEPRIUQk+HPm1MzGVtbwMlCw8VSBjj7sx
6e2hxVl5NQ+t5igI5qPbhy891y4vKeAx1TfzEo0Kkh/uEzvbjQoV7u0P5nMsEdtW
HIto0yvtPaV8Ctn03USFa3Td9DXxidReK6SL1VQyJhdIJ/cNmwkP99A3jE88mu8F
F9WXneOPT/DYgfIfo6EE18Bg4dpg+hTi9WUybzwdEUBESNGoyHRpfA8ckeCNAMl4
1qVukDGzW+uqJQvQpEx9xzEcQ4xB0yjq+TTM9NbWX3+5gygTRgEDjUl9DlPvP7p3
qJ3JaSL4N4KUprxrIwv44X0mQH/IxXOE/ucfhrVuskNeuNqBsfO/KfTiEI3w55Eg
LyN5k603TpmQZdSvkPpdQgF3sv5vQCpcTLRqggAuopLPZa18mJmnxfo5CXRByosI
dis0Ue4FGlBey0DXSv14Aum0lpm1SEQeb5mGZw4ARnMINU3FT2WiByU64qEThkGA
7InbmAna9leWnBhOf40jb0J8FXQDi64f4FZ1EuJ0kjyZBhDxaj5a9xc9yPm9N5I4
ZbP9LaoyyRL3YAJEGBHHMYeeIlCCP+7pTFmPRW8tlDwDP5XutWBWuRUg2g4oWvvD
DTdHVCawVTq44d3oxaSvrvMpm6xkJeXxL+OZlFo4hKzr1fWjdqYlkxEYw0jGPv6p
YiiGyOyPTmZhYKO8yaxosEwuEAu7Y5mqvcTO8HR/6jBJtDBFuXEgUbPf9nH9OvYy
ob1OoC6RieebTaHx7nu5feEJdQI/DOeiVO9m+Wu92o1r7QhQr9CazwS8PRQrvgUJ
3EOUOICZRS9XiC0C5NaiPkQ+l4OYhi5SR0pArefnFVbV6NZ3e1wZM4iBrRaHBGzH
bzGdZYzsuPeuxdBbSipYlqvzJfxz3nKwYrTXw6x4Yp49w67LLivf4FzOqmhQCwkL
NFBAijiVW6tuihpi3StwPsPIgpdd9F210DyErCZ+z7BE8L+yoQ1gjX00owx1FlVK
/9huGLB2tZPEvNRz9BALOQuGAwhWY1SFS/K56CzoVU0GhvzyL1giO8sB/W/HpFqw
gHdtp1hRM81Up9LAqVRCykJDlwHNq6EjPsbyKE3xrSuDF9roe8BjKD7kNMHO//BJ
ZH19xT64JyvCIiurlsumgBPUz8IPebfFUZoJb8oi50AdgHivxLfzyOkKsgq/fX3q
3t/Io12lpP89oyI9vsKOYeEF2N7CZL58X+kqlcxrIPwAkqUGHok9rqaSxW7Kykbm
dimFZehEOcHN2j3irL7+iSy3HGmrl1bswANv/p6zJIuhEXdhLu4HVeECo+TKDIn8
pwncgwVav4YL8WFIww7b2XuSIMU15GAkV6bu+7Hakpp5hOFGi2FRXW1yRQrz2+Xw
zX7Dg425F97qr+Su/iiUDF9mtCov8qjR0077KRdT3BQWznFZKStybCAGxCVMzidj
4J5Wjsm78lZdPzbzxnZRiRiXKG5js3jEY8mJhuyJoQX0Uii6hw+rXgX0NpEFOPbm
7PpNKOPwB3a6I6rf4Xk/T6anIREDfk5V1wVXQ8FDxYvAdM+3QV6EHe/s7g/MH72v
C9HZUEVkji5AQ+SPr/SK5z9a3yejKHzKmEmKCQzclkPql8bGD1bsdf1Y4ALnDeVp
6lDv3NZVWORUvD6sRhARNhjtfK/DCY8GL6A+rlVKQKFXnkKnfFEoyCGjA0N1xOe/
mpkX5TcMf51tsbQf6gDQoWhqG/7qAMfdlxEcnn+BBUM/IAT0zsMoZ/teRBD6uzUR
InLi2pPZKBNm20UMdqEcIE/qgLLPQGmg3CK9ke6vyYEO/eygYmUiOU35E5dX0nGI
m+pz3z0Navq6gNt/p9unJOkezyaTSPTfu9OcpdDz9gRehYy7+V3/cPbjhnVvQto4
Xn76dg8Zqf/1w4rTmqyh40m3sMCkPetZTfnRUxaJ3+VJDw1IYHVZ4SJj6pPwQwzC
mx0HB+8HE++pxfCxAJT2p4kEFNdY8mS8jhkg5SKxezsvC5Wzk/7Pe1bKpuJNBGjt
sR9gukQ1LnbwSYYEvLyMJeYZ+kkA+qjs+UwAg37ZWGm2cJH4p9UZC5eqLpxNlSUo
ISFY6UE4WKg0e8r9t2sm6P/OnOr5TGw++10NyY+mYu9Gcok6L9XLeeLL2rnLNyvz
Ce8YQH2gXdSqpja7790mgvvzMWzV/wJQmcTIx1tUEYgNf2i/UhLzxLgAFfNdjFWM
SVin/QFwdCH7RVJLw1TDEQDoO0VtIXuquBLYlF+fkp0AhwdJFkdcHndJ0sXwhQvn
JSXzAWYtpR5TzZt3nSMOZ3/isEeYme0nMNEEAUCSiiVYGC7SzGBpHK8n9HHoXieU
LFR1iBPZcreVOIyydwYcg2KHTlUjyHd+xmy0cNKfzo/LeDg4at8LyzUllyInl96k
mXakDxp+AyiPIvP1r8BOVs4AD17YFl/YDE/ht5GSWh3ozs6AdCyPwYdX/dGa4tCH
urBAbUjkL4bY056VfFniBynMYRsNE7NqcrvO+vyjU2ZmhUyRWRG901KkH1eREu9t
MDjN3GNGpzdYq0zGs7RmftLf+cL3udKN7jMPqoTaCNmsoE7YDAY+Id3iLOPQ6qNU
ne66KvVLacRb4B2tDu2Sl7BVF3IotPiXfskfgG0lyMsXZhhuPE7jHN/2pTexwxj5
rsZQDiF0bjsE1Uks/rZ0YvtqYC9EmscpAnot+mI7r4Evl0ugQSVUgXdhTOvfkyqI
3OI3L76BEmjcWeJmy407Fyjs6/BSfTMC6KBzSssMKTqNJxEdKvxW/HUsjc8g6AdB
U2Bm3UuIR3EzA6t3vJ4yin7GeOTWvVXJQ5WFrG2mqYf10tPQUJ/KQHN2GvtuCwqR
vVzsQp6Jul7DGJMnrvF7oGnkbuBPAq++h6rN17AiSb2LO01gLmhPypL4zOUDYiGa
FpewDcTlsX/lesgVzHTAGf71CRQkiRDxvWlL/d88S6GXF6DP3MaTDVXm7Lara4Wo
rI9c2ulaJpwW3m5nei+VYWkiwL6Eo1+Y69a4N0l7C94mrovnfUKBwOM4crLGrAcH
Nf2tdnQJcOni0RxmXfsI2NTUUNSufBw9Zc4++pvAIxcK7JUAATXmfu07shcIFaLi
upfUZHEkMspGJqcExF9hAb84Gv13vrZAnnyZ5byNpifCAQOGFb70E5x5Y11EB1n2
IfgsNI7Tmh8rfmiGIY7IKRTsul8VS8vNkXHHowoy3beUJULEz6qDY50JU5akXNdD
sKtyt05NjIeHPAF4eSE1TN4EFX+59fijCH1gDSjjo+2XATBN6iXXnKC6nUxmqtFb
Tgb5SLINN0TPzBtSKQE+ATHqvAL6VW6eM6n1F5lxfyxJnRcqziFntwVZj7gIlLmz
pw9lwPhg28djpM/5r7xcIPq20ymsw9vigrWefuQc3Acy8B12YP9TjXS0Ms1SrP0u
fbqenLbdV/XUBLc779m/Lh2yy3Ac6cjiXUQrYFcgwCclievQdgRjTjtJEFyNcudS
OeSJlQM4HGnAkjuA43KnQgAV22mdIWEzxjpVfSfCt3uCsV87wxrRJm/WdA9kjh8B
nv+TjGrsGyw2wi7F3ANoRpcgAzXOYPgjk1ZKRPczE9cYanG2VhTRH6HsZ3E4M7hq
95g2l4tGqSUMQ4DwQybZoYW2MTtZT2yyMqZrWIgEPklJciWHU95pBpERFxu0nwTd
BwYhXY/z6T8lF9qJoVFx3ruREdoS3uUyBfaEOrIoS/4TTOqOeM/QelYhXCyc5K1E
0HRK8nnkjmMY4YqWJSkPJs7GgjpXXfUx2DCwxNEn/Lk6d6NyO3KuEO01vH8haLLG
McqZ/bSTgidcj4u5FT2EGn/F62pQS5FybcvQ29eihCJNv3aNRIEmZy/ITgibTGTf
0h77Lh8PAqU5xI0eUa/gXvKxTpLHYUxRgBlFS5usGPl7FPrsnqlr2thiQL6MgY0G
SMhkbCgWgSZmUyC1DGptTZoMPEN39Xrrd1X/PZZSC1Mv8llecngM9VqxB4oeV5Wb
ZxMd2S3pGu/3S3e6tLcg9GvhYH+hR26eTZriydGqO3+3MAR9UFGQDHJaGbjFRSOh
cFCoiLESzGKDt2dlmX3qn/6U6MKYJ15c2KFLPzaDg4LhL6ljMqdOG/uLLEv8IQEe
BTfbI6DA4nNvMAPXD8zM376RPXquEDCyz39KZMm0YIf4QvgT5WRMJHOcv9O23oRc
fDomZw/cgSrwdVs0i3WAp9x/IP9lXNJ8VjGMzD4zaDC0CDsEeJtN70T2e+0DvukO
xZWbEQzN+cSTEZCEmwRgvENwPDN6tH5I3wHznDZBFLVFqOAG6d+hqDcUgjBsq1eP
mHIjfcM+Nbgi8YfhIwhGSuJ8lFlDwXcEWCZACjVxwgSAzMPshRkAyRZh9JyMPdtK
POeMhbQBTc3IMBHUrmCx3pg+UrPJBwYip31RrE4qdYUHQSsn/3rfHep9sF8ymd/s
cSopPnmWOu2EJbsfGw5XQ26vxy/ZQCgzXCrI7FOKQ9Tu07P9GFaVnrOgFwlAXKSh
HagK9xYac7wUu8jxfN5yMppaQbOTOjT3p9siWA1EXPVRNKc7CnK6gi2LH3x550A1
xwjxn92YXqkuU04VlNUBcL+n/0T9JRlHoaiIQKx4I1A75T4PPLUV51kYQiGMDXx+
YyjbnIr4KnH9gosU/TCEq8xKdv8ywYwhKIUX+0t1aNV0SAZ50CaW7ECCgVd1xbpM
3RGWFeLOcSzBx5BVJvLj8UywssSEEHElytystCJTMZ+Pb/2Yy2gWUNhiZ38Cv4Dq
W3b8oLvPCeNthocg2V/gU1GHhvBo0AIiULiNGlRhibaU72zZlSOfwx8a2nKvuVGG
VcX6LPizWfZhgX+Z7t+Hs51H6strallJyLLjvqxVP0Sc+8a14zU6tT9q4EfUSSGz
ZkQM8BaGOfDzinF1yyhoOC22natPxc3E5Dx1EXIKYjO7v9FU+RYnCdueqCzuJaa7
qdvm92++PZn8ThpgTItOwlPVzaUZrizOH8bRJfAAxMdOVP0BKiAC8LF8s/Z/34po
fhJKnwi0S3e6nT2CukU6gVu0Yqg2rnrcFfUrvrT5a3IRbOAPAIr30KeWUtu9kqmD
VJ2pUjs5wa9W7GK9a93+6RwORjfEviQJYUbDD4/SfeE4fYOE1ORGKHgdy2tL2ASd
1Ipb/Qr7TaASMpCQ8jcahrF6U28YwCQyJ5PouvrbgQuG1nTmqK0jIUfiVtJs+kly
I3ie5R8O5U+NJYyEdnoDOmOhV4por8ebGLHFomXZ86RTBNzsprigOoudnxsq1ry0
7AivrJvggtiEaZvj8YQTS+xhLdtMuJ+GrpFzV9HUWNppHpeROCaAcq4NaPupgPuh
G7bX2tmTu1MNF89MAbZTwaqWDmYMLJVpnB/wGAPCOGpYQpHPsiYB0cdtFCkyRCvl
WXgz43H9xYa2nG4nOsAtKlArHEWlVCESRxR0THzB1fdTCUrFvkqKDbrIfCTsD4zb
TWYnzK1t/VZi1yuOQ1hSr5JAXtGT9TtO6Q/cK1KB8l4kdIsG/VrD2r6+y0eX6nJX
FZn+QaRiOPhoH0AIv9a8roYE6MoJx6nekvmZnbXklDvZHq5j73cbAl+Huw5kfiMo
nZIAyeionNWp1BV7fqY3djTQGGJg2TN9y7gu2QsQ//2nk4wlNEyzljb/PSceOVcO
rKiw8jI5OLVFr84uQdPrmGFpwMPKXHLjN1rqogaVhldbIgya4x8JuYWs6b54bKFD
idy06E0rnZHWSI95yQ5eS87bxW7Gu/hPt6bFsNGJX99vHw0bLZw90274A5g9FlEE
ZqHi4JFiEDHtGOh3msRFgcL40TEdoOpuHm+OQqkLht8HGjddfpsmxjhzjYBgkq44
Wfz/I4WuaihF+abQ8NJWes0dH5LSXR7Qe/pwcLFKwTFAHRuwdPyRuCutGYRlbUAP
4PkzoRRJRZMIUneJWQCDf+rLH64/iq8AQ1K+1VKLiJIkXi59zRnHSbc/dMS4VHNw
qIO7wOQB811s0xdK9xcN7pRLz+xn19rhGCZTVfs5Maq870q1oOuQNQhkGGc/psBr
V6AQ/aeYQ/rli7djGPseRuftWAAcYlWBjpfTz4LiIdHmJThL3E/yQxS3WuZ0ccR0
6ggboqbmGs9CGyd6kvQTek1eaRlGOhPIN3p/dsaPGUXI7Rvf5kPODG/JXUEs03fL
kpq2RxR5YWqdtUSC3ZHEI88215/QXXODjqOdPgGPQ29O5IvTFTAcSP9VhZu6UIxV
ncQnH2bwZ10FvWQxR5f2XUkMQvfvB4RWsVWVGavnk1upldiwkd4JdZ7F6QKxO0xN
VPnWJTrCJgkvF1QzXC/2dBH3J4CEvgXpG/5KFDL7TJnZKf7Uz9zBZRJURopjZEou
CNMUPTANP3spEtnj5/KmvT6SgsnG/harBC094Xa3QMdv2gYWGNU7sFroLy2xUhKA
nkHFQkIefm32pSbioBzBFpoj6O6H5Gfyw53u4YkqYu0WTKI7bzLxWu5TNOY//NX/
ECG68BLio0M0+YMWRdBIv1MRQOkNXB6VXJRZiA0G1jWhmAkSWeAn3x/u+SCFmsVz
npQLTQDHdUHjc0SW05MgHACOvRH4+kVRoJC+60vk0icZhwl8AlpoNumR4fWsgWGU
GSNlCXn26UsAr/DjZe7Bcs/oHWlveghEslBuD8o3dMW6bv5ZbU8l2Uq6R3LjYE42
qGz3UlY2Gny9KbTi3VoJ0qvNFDasVwnhmpNnnNTdjOkwoPaGlF7wWDBDXeTU7Qc9
ei4Fv2W4Pjv5bPZ4ug60PjPzntK1eiGaLnLVJMUwomV0l1cpdL9l0xEmLOWonQbB
LwfkIRnzp+TyQq3E61qJF6toTqYGwtC5suPLBo6Nr0FWbjMDuwUe0hCunsSeRF5e
Ns/pa6YSPJH2u8vnr2PYB1Zul8v2AwYB0P8pd4sfl+gFG0kwQpxMCSZyySf9QQ6F
x4nbt0ff+t0Nt5qSmy2BJ8Hz+WO5BIgc4vlwkRC6r1pw7+FhuWZVBXZAXgwZ39X4
VvIYJ1UwstRB83k9UDQd5Gp9gfPpyEkuP31V/qvrkfp15szZwrMHDyjESgvYDMrJ
6O46TnjJGNTYPW9jCSumkj9w3RXSD/QAs47mfalAzWQGKNhk3e3n9VbwgE7R8+aM
y0664XLLozrj/dHn/ceFEmCnO2XChkR/aWlQii9tCxeEa5Q2QAiCVpaED9SKfRQt
lo7o0r4fJauGCZ+b8c6cBK/Z+IoIi6lAM5pR4z2NFYockhaqg/WBcGB/qnz5B1P0
oO3W2VRt/F3epbk6w0EekyHvsJKqaepkN/Lv6xaD3Xd3r8odocwZU51QpccWLdbh
/km3zlF7uGKChOZo7rT5Ndl1Gcu6l5gjN7w6R48qTZU9OYKAANz/BIdy2Rz9kFdd
7wjh/3ltmWYfxiatG5PVxioZFpWTZeABTOGHffKaTKeqSGbNto7piqKzmQ8xEapu
5gE/pKtlsa9zeLEeN8t+ox+a2d8RXHQLzYaR2vATZBLUUsSi9YbFVFDxG1SUgTEu
Uo+6xzaxC2eUZEaaS+DAwz9CUKxNPMM+m8hK6R9L3kCkwmSC6rLvIbhvT8NKw9UR
1S92r+BuKoMBZYroylJpT0lUWWl6RNlLsr0VFp1HAdwV2nIeWgbqdlGyQEYjoDGl
oJTZzOdB+jZjSd46H9sJ5lODJWjVGUz/PN0EpVkig8r6mf6PUfllzjrhf1ZPeR6Q
8/TKCflSIgfIfl7GZwSBUyR4ZfCsoD/ZCZ1AjRDcOkGDlx2oXu05o6TSUj+nR2IJ
CxAfygWk6+3OY0I1ITn9jO1GNJu054a1Okj+cUcK/sKJ+QWaG3yxaU0daq4J3fm2
Ymbi0VkC/lGY4KytZ/Xeb8zcUgeGh4KCCnLEW5wCuGbE+Mp0gTqRbWMeGpTwSUP4
GmFG1MLDX5eziORW9VSadHPqbPGARl4oTBJFv+GeI8RJVoknQae8rT1VzcG5lp2E
UJ1ETNJb/Ww4zVMTteehO3nyfoUj6uk8etUzRkkLuz3MoF5V0PsjH8rjHiKx6GIF
EoUtqHQQwro+/pNb3jHtuTj+RmCrWKx81aBYmIsKwrDr49td5x02JpqbdF7LN3F3
EM0gvvCM71V2p1vzrWz84lnA9ZnUBZ5rY+TqUrgqWdq93lLwgsw/ij11Lq3cN9tB
C5qU20TdHtDC55dfe70JrxJfR3zqSx5WOt74wTrCMe9+Nr52sCoorEicM6LmOtT/
iimfmJtf+jtHiRf0lxZyEsv0BRU0VYTS/T53apTVvuuzRkh5wyY2blzj8j1mr59B
tOMmHnKenWhmZTuOy2/ovTHTNDIaZdzVs7rHkir5xHWVlY7VhlabrIPqnMaE0LEl
cnmNovAA312DEiS3P2cxgqgy91fGJIZi0iuAf2xIlD2GjQ7haZaiLx67ZdjBZhOZ
LFLEeHz4+sJ28Js9cv60d7xDROlx+hJwCgx5EaYr73aCDB8weT0++e/Bjzb4mTaD
/X2G19ZssnPZEgZQaBzbV6QTlTKEF7v5ihMZl76Wl2kIti51sltQ/dgwPGwgrGSV
Cj9W3txE8gS/vc9J9/XWq63fwddj9+aJpi6zTSblvtx0xgaoCWlyVQf7keVijDAT
RwSJ+zG0iAmyckHrLDk4ous2HM/k8md+MYBgJKl0drPJHkbhBteZqDeVzayqXQ93
/5jImzPZI2l5yE6TAiqBrRGHSr/jcUoX2hSQAJetp7RRHF4j4kcoYTw5ZMXcsROf
kncylSCHsaIYSbPj04OKKyZJuzUf5PPkkfYs/mW15xcRlXlv9w3ZH4EKdimwfJDS
DewUDnLGmdYMq4K+HWqRaX++FkaB0FA32EARenbMzBdmzLbDLIXUA0WGmo5+mDpF
iOz8BK9Sm1v8UcPqrDxirvh79uOlbXPC7lV6S0t24ugA6lQ3ZB7O9BafAh+oxLOw
v/FFNv96/bSMl3wfWE8rqVKBSX7kx9CjyYcxi7FCODpzzqm/i9GHK8J1bRhgGNW9
CmQnMJ0yIk1ayRG7wTqd5ysWpZk5aKtYthpcCio4zLTMToemb9ffK5hKPCVVEFv6
B44A/Rs2aMtrZMD8VNI83O/GWtOYYsShSgTXQ7jPYh9ausEedFjR9KbQmLlIab+W
aDL5Q3KLotTNvfLj5fwEvmyFhZ2oygS7KpSk5JKsgnhvF9pVlzKVZU+s/uWEFaPh
4HcYT9YkTuzTNtzTvJHC1DLH6oq/yhWutwnM+aEpvk+57HEg9Zsaqd/i/1YDVYTf
QwKauzukv41Ob4hVHeD5zWtx9/ngMBEUE93PzGTT9vufEtw/cyHJRPqfPlXRZCF7
kGSw2bOR1YmwyiYvCXPfNd5HAo+Pqk1baQ/iJLCEIchfhsoi+M3vVxpgqNqTdfQO
GB23HZqwH8+RS6hwrsLlGMgY73FPQd9QyGsfcjfvCTnuQ1c+4WSZvd3n+iSl1qGO
02oWq1Zl351mgWZuaMxJUQXSMPpOGIYlaoNqvkLgu1MJVgo377X8rg/7CO+ICgRt
XdrT3H0Z6pJhTKlq6rbTzuUpsPgzHay4NUUgjUpdrgx2dYLnRCktrwA6DLIg0SQm
O4tcFajT2Bs1lTJ1N0Fr4EI79ddXbDbs2h2UHZhkbjoG+ukn+1XhJsTThq5ItvNG
RHWbWOOeEmZXJSiwb6prDinJ/KhvchljMdZgeUWad2pEd19psnr0CaiF2ZZ64ruU
8YcSH4JeLDbnMaNfy2beFFX+KjkKOqcOfcHc+zVrkhkTRNAES1a7nmnD2YSf4BD7
w6nPXUFdmB3Zr6mT4xBZYXv+GfHPRTT3NqD58+Y2wvT9aYIj0HWPiSlccxOINwHE
J4ILIbKLRbHqGCJDk46wwfk4VkuaL86jpA5ztPFV387HOxzCczKAvEjhLhhBFb3n
oPnzZXBfgxVBtdqlxc/ih7nmeHG6v/rqYJxk7jn/b0WPsfAg7eTJ3w2/gpz1JhhF
rjas5XXrtTB7taMg6G+F1u9SGmYcSXPCkS93DA9vlYSR6CpHJHoUG+j3W5Tc9U2E
Z9YnChNhukRio+5a8gWHHmjFkYa6nT+wE17MBV5hpride5AFZ9UopN4arXypqQw2
6uCRUdJTJwYeuvSLv8eXJF/89v8iw9sozupALfWJFvMBuS8ep7RVZTWW2QK49rbW
2i8Lu1a/RomxMd8OZzft04wlzkBVcwT/Gifa4FxzrU2S+xtgZ4b9Lk3jxda5LtMt
FbFQQS8Hs4sa/gmOAjBH1tc1vlQEuqEkzECQCh7m8gxHGQBc/gl5TPNTk7WjGcPu
Vji1bdbJUdFtjuSvmMMUVmY223ogPGYaOV9ZeFpLxHNHAsjXXmEvKDz+WT4cFivy
ObD1EZi+nsDPqqQ3XkTVfpMIO8OOp8gS9UI6cpoZQf/AA/PwgCZCGmFtI3PuenPl
YkmOiSUT7TrHlc1X+3ea64xLJCzg3G9/sNLNa94l1bgqLy0ytXmxP69uSK8Emg5O
3uYsS3hb/mzH0wWxIUYNlbBMaVm4VASDO04eQpuQEfkkAd3QCD8so59Jkl+o0HEQ
HMTBnnEuP4EQHY4Ja+QEwQos6q4NoAsg22k7wHyFcRwvOt55MxYSQGcrpxcet9aA
CfqaDfn2itJyWA8ZlJoc+N2yjz25rHMUnFDq2cFupH9CDStAxqOsle0IzqkB7+eu
HRsPdywVr+2Lld9poTHY8AngRT+Vm8h5R1h76eJkSkbIz5dmnyJFnNv1cjVrHYVO
Q0pIwiQUALOiDEkvkcBqjcTmUTPrlk1eQ0iDnuFuhIG+60OtyhqvjrSAvDC276ml
iD+ql75cSBLNXYD+oREr4aXHKJsTlMsaC9L92MHey2Q8tLhEhpcKZuzQXO5oAx2e
aEzUtpUhw/f/lUJft5UwxJoesVtlKuCjVEU3Du0IiffcCppqU1WDmigyrc6cbNPc
Cpxm0uYcgoGk3y149yIRTgB0VVMNO8KcRaO8gPU+t37Da1ofE6Wi7mWe02eazA+P
2BJj70Cv+2iI4thwVNPn8pTN5Q/uZwo+jjQboBodliUsdT4ys1Hq6/DBJ+YjZu8i
VHuGUX75Y6XRGrCHQOFWNhSabhuiM7ygPYLNTYVLJfmPaUDu/3rvdOUaqYbE8zaW
BxXhOEsx6ncgVVtPrrPgP4R8Hm+lq+KvmqYNLjSaxnUWonHa81iOWVP96VPLBFk4
mINVHJcNBJ6OXUEKLRgru5r191edsU5ZGffsuww12V6bXP5XfVDqMwZezlzxSt0S
J80MnpQS8yGtdwIDkI3zomIwrrG3sNpO62AavWoGBSNpN7v8+YKFXix9gra+sLwa
+XoA7AvwvJEbnBWrbfA01UgeJsEYEVEIsRB1qTZVpVmUko+vBReGmc1jk3aXi4cL
7qfMtCSqGWy75fl7PLKHVtun5nRNyNEJd1BTv2MmpecJQG+5siPyXOZ7eHUa46W2
nHKn4SHOHTWkYDdEVgJiDarA2p8VomgRXW4d2qLtqm7a9PmQHtQAo200YMZfgMRW
fhUQW2bmfhKzH/BAg1K26zy0t1aLAmeVcG9M1heWuvC4z3rcB+IcB7CoUKYBxJid
fx6QJHL3IaiAAYuVuIv+GCeTjYsVOcVevkqRJHPxbPGK+aOPZq8JrBqzpcfRlgbt
8VNGqodZ2OhdUYIV1V9SyqcbcHK0QsYw53HB8G2gbDWcieL8j/3//FAMvBmZ47vw
soXcM9sd9QTGMj5CbfLk5CiWrHX2GYzwUcUNgf53F+LEXJN2+RvY1/alDnbWxsww
L5y07uR6Ncj9DAW3eYmpYkzfLur4FzVOeJ1GBrCOypYls1spZiz9W/5jeum6IkhQ
YC+qeLmZTTjmS+alTp4iZ5AJI5m1hmWQEflNgIPHsXbXv7RPCd9mOjIc677+I2Ay
EEArQAb19/91xnuLOJcIYxLvw+n3q5SPSMumG+v6YMDXTAg4BmRbt+VruRpPDUOt
KuArjvNGGH1yuTE7lUh76TpjNcaSx/5rb2C6oKGpW0tTOuAiyRrefDT9K1tmDaWJ
ZVFVYyyteCbqehqavyDgTTtL0kSAzv1Oy4L6OJMhcET11+SSbFhOoes0D6TZ9ORz
UVCIL4hbL5oXIEj4jP4j6S4iB4GlvWy5Mq4w5NvWBIynG5qWm0qPJyF7Gr9G1tXe
EaFGUKTc+5FepfsWebPou/6HTrkeVRys/1oci5KwnTvD359gGdtcGGFPYJolMDtX
dOjGn7Plfqiiie+BEYV54qO2tioDqCopa+3CZGAWDtrZ6VKB4Tc0WtV/nU9HH3WP
MgPZ7+9hzpdh3iJ0pPOj8GfS4VokiKIHbk/rhEpXAN4KP7Lkp3k+oS8wfh1OJpqt
nNZXGP9thpSyGIaTvyjVRKnvDXqwHjWbdqd4YwkZVRiS+5uk7S194af0Vn+WTv4s
AnbwAiyu/cZ3wKC3Ozru4hV/bf2O3mVs8LLdMqwQkYzcxnGXaRaJMtWC361lunwb
Pqkh5EYXZGSG8m2ZYyv0zpTSaS/MgkdBJDwvAh1AI6azJmjH+x55TBsnov7Z2AUl
M3H976HKYQHEPb2Fsj55in0C+p3VoyiCdBs0cLSHBs0qm7Q8Wk3ITiRhuvt+0Quz
t6WILY170BdP9NpEjl6KyWoJ307TPGMBpjpVxUjorxqireM7Js/+gd+OChFFPcOJ
SOG1itkZ/EIQl4llit0ZhqiGN/mW6hzIUF0kxGwbzjDWZyeBxLzVevU7a01Un3Rt
9UbszOA+qtGNE1262qEW/6bC4Igq+TeZlkA0EMadGnSfz0H1hvOvFEXRSE3vHOh0
ZdVhYvxa+MFVxHNMntTyF5NHzQGdt/VYH4n+mISmVeE386QiM4Us+jUNo01FZerG
ZrKwnwoEupbyjRCh+JuIexGuAdx1PcfIAKpe07rOtYBg9bw0IJV/LRp8Ur9ylyA8
1Y286ZNWucUXVWqt1z++uKYueG46ZbvuzVpy2HhLWaNBbB1RYYEe06ycr63jkqAA
BRiAHW5j3KlnR4t5rekG9oYJCuD6cvNNR2abim8Hmo1iwZZp74Fdncx9BKCYCDKo
MewPFZyP0hwqqU8v9EmOWVcWd6trjJ1eeZUtj2Gyx76Q5zko9Y72pqonmkm46/yR
RAgAqZBKKeKF27i5+EKv02ZslmY6NSbVmJ/F01MeSQUeUI4wktcH9gKeD45vPFky
V1hCcnOE895NqEtJVBABozaz34y6GP0zLYnBUuv20P/BfsKALcGfKcUAkhrGfHde
3ZW738k9QjXx50XWiOsEMEC4smDEikSWPoravx/mbUXcHtriQ8HJLP03xvBsHGgz
1RcTlUhMLiDeHWwVzIltGXSn8tGFH4WDaIkkSaUMTUIEDRHsePYRC5L7sbg1JLGZ
AL94tesSiC8Yr4Yj8IZ+DdRUzehvI8G0e4A3/yk4MiYvtCkGSY8z8nukRLE/DGB7
6SO9f54Bhj23G4x+yzwoRjzqzQPBuMTKw/pAFAlE3VU0nRcUnNUDd9UcxWCf+hx+
sdTO5PoM3e3DjAqiaM7r+gNDeLw9L1VtgC+P3dNUxRxdgtTMg12MYLlDTcVF6Uxy
LISCsavMd+PtRLaKIy6FTa8QuHAckxFeFyGgSdFJ2SSG8GgofIXzBmmCopoj3lhk
WfzqKcdZpp1xnUo2Es4ZvcZyuRBx0St4BjXyZhvk7DFdg5sAghTKeeAjpkAy1T3b
X+V87smBTxIz0yy6/eRtN7n8NEOT89nAQrNrbp/GhJdsC7ZiY0J6cpwKUK9JKdPd
/F4Qk0NNwAt/b8Dc2i5sVvLrR7XZ8vQhnvPit+KGNlJJzoswv1PTHlBEDVLYBTDd
pK2RbzQFTSPMyMZwuaZgSO/8ykbd28wJfBFIKaHXpd8xoKnFa7Uc8USwt0jhNMvF
ABPm8uLAugM0XqToSYGIcMWrK6AOmvE3ZZFKfednjjPa6x2cfSsi98SDET3V1qGT
fkR1pqzpJwzi005qjNGXL0gzfSZm4DuvgQBDozGNNQ2Yizuy19aVAwCnlq9Tj86t
nbNKHXnXB8AIcIVBSP74mMKljaeMhrK+kypV0Lb4S6yHQUiC7BX2HcAlDGtLSpK8
4KcdMgCZwT1TJEPB3NLDiIQkgVodRjGrECw+tFWxLj1Z5J8J/xbCZWmcUpTxiH4j
B1p+lLCyxEJbqNon+4ICyrGPV0mtS68m8vfOEC4HA2ylqyL8+Zliolmx6EalV+KR
b+GCQ36WX9Z8J2PTtLPfnYANi/28GuPxnd82UQDd7xGNAFn4qWZH7FjxVib4dQ+Q
amXlSgMS+phfuqrM21qM3/sEMacVrryxHoyYKrXVr/F7Z35dtzFkeZRi7GSooy4Q
1euJu1dHRcCT43Wcd7rnVN7/Ok2BpEWgd7K1Taz+wpq/iyS+Im53B5sJ1hf6YI9D
eInCDEv+Cd6sTHELn0Oxivj7I/JyIchvWy4u+aIzBgW2RaFVZl1MUGwFcnZocJfC
Q/lYV9aiGEyTaj0an49DQKnNMgtRFO1uMQojgewmHQ/yr90HojNjZe+iH6x60OPr
ahyNQt9Rvah6sn/g++tDq+xB724GbYyBohgKviQmZ0o2f2bGQNPfXByI0l0ESVTs
va9j7nm5R08Fcf0gcmM9N5iY1SGMyKVSNP4atEUTu6gbgBjD6SSoGDhSWckjpMij
bLsnlvcc3kPG2qyYjX4YH/2BvsFDzwswKGB2xlcsk0J+bsq7Rm6fiGeh34RDdWLr
RJtpZdR0IhZ4ZQxKJhbEzghwGdlOiTrQJyFafoKvCYS+f7Z+CSWgNasX8NOY62oA
4jw1savd39XvCeHewWfWcSA8AS3d4iQ8bvic8kGT9NMmBK4212VcbpYeImsqnBL1
/N4xnA0HhKsEzp5hIzM8PEXySbbL6ltKiRVOxqZWRjjW7oJn3kzaOH/u369+knPf
/JVei7mKq3i7s66RNZAO2JR1yVyr+Q1QwUzPNdNqST7tiUDLU5sG01DD/sirmIUA
NmIhe9/qBLPONLmOA34gewU1tA//nxJkMLIv5Wb6FUwR9pCzlg/zavMq66kaY9bb
jW99NNQSypIqhPINPHZunZVlMGmZV1BU7RMAvYWPn+4sf8rl4SMehuUVfXgc+tnV
0ijXdj5m+g+U93zFm3laNJLsXxaSF0NcRJmWDe4rLqEYUvARlcIdhSSn3jHYhkgy
ZcewH6h4fjSBOnUB1N9AIp4yc+7lfv/CR3Yd/T4l9kSoNUAy6Yil6Q47fnbsC2wI
vilWzvowkS9xtAdoEoMJWYrdHg4kdC3/3l7aKq11u1/n5IqFnLOLRlwDbvOV2epN
yp7KaS5pVjPIxH6N9gl74Iaa3N1ZSTi8tyfeb2tfX3pLx+Wgquju8oR3blSklHKO
M2Kbijtj/F5F3KHDRAjTZIYhlEB+pJcDN93y2abalvdqiBoYpr5r6o00Ll6N9vqC
ntts665etVVmS6MR1z3PyRL21AgQM0nKZuYRrM8NUJ6OVXtNa1WoNlV4TmIxK53P
pPiH6WsClz+ChVoZNeGDPBGzCURyK577AoEnhSdtc/F56jD2AsUWZSVnSFvtnin1
mMaC0mUf90Agubu3jzvHL8vCF/hQyazK5n4He9Bx2xhPRl8a4CNayftPxIYi72Ht
sQmHBuj4sgq6lIUs2UQ9hzyENvq/HcPLjwj9rsbY84gYLBxCoK120aZQJumFfqsQ
VJJvOD/9hN38yQ9ucJtIlUkVDp3lq9psPuP2hQJsVheejXPpiRngCYJtOVbckVvX
mPFUzvOAA3+nvmkM2R4vkNieQXjQBMU2ZN0z4oxDuUnGVX1Z7K/WJbYTIDX2zl57
+sNuzOowzIhUEPv20tdquledh5fBpNHOryfqw6i4hO67w713MYljXdTb4KKTqyUD
ctUcJj4/U6VbtsNS6UO6by9n5nczUwasPldfau5mZ451Q84n2T0XKvHvsPBYxFVt
v+3Obcvh0eGwDx90jDjbCEGnHuKneHlqG2UlOJR/0feud66b2esP90vflL7sGrik
5oAXJTn9a8TnLEdYJteqit9zIYAPL2NH/RaZ9/C9kHZv6ewzCPzRlotiYtnaX7e5
ufR1kbbOB+OqNOq8AqwhYWJbVmB9UOyM/psBBxUlQxx2I6TyJf6bSy4yjC+OD0Fr
+77QIVVeWqlpQmnZiNq+hRLnvlbiPlwDwpbmD1A8K3wMhNJX6Qm3IW9PjKHZbmun
ch0DotF66HS87WJm1GMuK3SEBwwcqLXQHOSVBprtUYdCvfzAKCyCqQ96vdLzdPR0
moC4C5a0+qUBvkTBN+YP7hWefFk+zJDddQWy6/fAGxxPEy5Z5hkToHo9Mahn/MCT
/b5ZWNuUgCuYdQOZQn8XyK1wfB9quDZYXtlGLfOwiJuPBn9JSeMub9hpTGRAa5OP
1yR6dPk7pr/rTiIktzmhoDZjKoQwgRcIoqg+mBDnUm37ynnGYYY7ELNzcDudNul/
CCHZOcPH1Qdi/+lu6fgbqpPklBAznKPsUC2It9LkEkQCZk+4zOlHsshjgmHqe0Y5
vtANM+UpBXW6EHRSXS9IbPXYelQC1+NbBfjDvYuVcfZBTFX8eo6eP5SgszTVt314
HVATw/fPYpQRgywsJV4HeJKAR3xynSjYqq0j3Imf1M2KXjnG27WfT74Y/xHDDALt
AqHx6pHatrXGiqpYxR0UJFkpuhcphPLf6+s+9dMWq2nMfMCm1I5xF772DI+dfcaP
CjFPxUFGJOnb7WqdM/F2dFga2l3bh/EVxVliyxw3tT7pzIx0qn2YRxe5XXWbxY/S
BZxlHxGaz0Grqd8sgK++RFR2ZmodesXNINc32Q3bYumyIvFn4q0XHqywohxWzYe5
wrxLLMcx32Jywg637gcC0TLacgGyk/S9HGeURUaRLAzYl3oeRu4M5D4BIMmzOWL8
S4ZJi5dNWE++Got2RJTqDB8AOlaGdf7UOQSGmP5eDu/ubtLB1WGHptrPepLh+Z0I
8UW+vVAWX2Qw5Xh6Jcl9mowMVN4P2mI2GpoyAb9nlP2uydkDXPeJ8XfRN1Of4ePf
DCTXu+Q6KmpulOO4P/LIZ1E/m8EGs4gYams+o9r9kviSTdxnRTz8yUzAVqhMjkn5
LWvaJJ9HLdX9XHPbKR4egRqb8IUD506o+Hy/5Bw3S+YvNWrMSCHK3lN4Ic2/JeB/
NlkkW1TNSn2Ppu5YtyXAlaDE9u4uX8QfNBN8GxGTr0bj+bpQtUdwoBvAossBBQDa
xtv98dZaKn9Pb2/zdKL4YWx3Zi802LrOhjpTnSdDrhls4L6LPpsbaFHHQM+dpqVr
oLvb3pEUHhmEUu3dXlWK8VyXWU7W/IwXrgt+0Zv4sKWdQsXOdwYUWIHCxC4lQkwf
TyNNLM75IkApKux8dtDvo4BkksR/Dp32qtabE5rABvWCDC+UGNwZPDfcro/v+vyd
+0zsaKzCrsd0R0wIQ9RBj0wq8noROoHpVm9m//R3cZdYJ3TzgIBNpxtaPRfSFK2L
ev/Qr4UmPTmVtcJHWcB+SZqxzjLakqPVI65rciCRFqeeyayrZFgM3rx/hcZyS0/S
h8FuFTKN6TPL3cMSJSszhyJ/nzHhnVOHp8imxNdklHJZkpBIhb2xHEzzRPBE/khQ
x0vlJnMlzaxoxzvEbUhAsGQEKJOt4EH1d3UNTfDipSEca5NhQzPIsFlGrgzLWBIb
7iigZcLP+fBDGxoKUv9JnlP8rMMvEB6seeyGVgnx+hl5CEqLdQ5Iu8Q6Ozvt2TrZ
ngBQAGbaignRLFH0+k4Nom7wV4SY3DxV6tIPuLKlu+vS7IMFil86/MLA1U9rsPao
cmVITs1Jea/qgCHXLL3pMlyk6ETzU1fH3j+KpfRWKVKXEeD/crtuvhCmZt3+qNIZ
vpgxi49H7a9ettVz26buSw0j/YoL/JUfjB0yLCnaf2UOwet+z7WTV+Qb8/Ju/Kqj
40mVbW6xxXJwygAoYrDSl7WxRtAGsi4OuEsMeEKWrvd3g1Je1ILeZQ56fr80lDrO
WOMYI1AskGkKPM0YOqRemKISH9SsR4K/fonP3BYgu+ELrWUTlcJ3qsOiFDI2heZt
Wej80KXY50Rw11m4/dw3dk6JCClJSMNHfKGPUcjKqjcLTH+7jRxGi8mMiQVN22m5
JgEA4f7+DS60/9RxyVZxCV3O9J6SnmL5yG0hJJKOrEfFcXVSJsyrzcu27adoUyxk
REVBxoZ0hdOYL8PX69wZkyU+/Zf+csFX7aMDK5EGjfPZFIWkAv83ZHDUe7TU+o8i
PkRZqgIf+BHpEIFpCQIDGEWCAEPNY02BVWjCPKT9P7C6VITnAiMeTgMD/pohIA0D
1hN11emPlMwCOo2Vvcxfw/5JHyRYzgH4bYXylm3BXClh9DT92H8rr9tJ7elCqEgb
iidwZ+UWh65uNi8+ECVI6v23NrXZ0mB8ccwTygh1vVG/nPhhOGOx6/XUM2CT4tcw
u/cqP+kjZIvXwhZNhKRIHD33PH6RZ6y9uSL0Iz5Kvu3dNh+eYH3pdApTEctd9Ngh
cvsIsfzbsFYF0tZoO/zipWfDZ6Yf/cSzkQDYUeeFRZDUEqekwt6CGCfVwKWyPe8V
eJmrgtLDaGdgf1AAIY0rFSqTngGXorOt4qKMEViHfKuvZV/W6Guina9XDKKj/8SG
rHa9p8ParHq3IILg55/QI4kN4XTjja+CeWALpKw4+x0Z4Dc/PSC6fz0DZ8vBuin0
GvwRBteiivqr8l1PK7b32BBKcEgadITbr38TL/TaCcQ6/JM3eAFCXJk1RWOay4dL
Nk8PblIGPO/whb1BklNls32SGXOqhiHSWljsYNLGM2+4iOYEPUPvh1ZxbuevSytp
z9EhBBA8CgVQr+wFvb1hYImz0RFxyqka20GatU6PAqUsA0KgmMEMr0r8WKXdbLLm
t5EP+2+ufG0qo4mH4eSwJ/oZoQNxmG81Eytn1PIPOVg/AvZb2sJg0lWX/FEGo5u9
whz4Na3l8NIyBo5p/fATYJrEiY4Fgi1dFRKR3lVXfOyah1ZR68D+ZqlE+MNVVi3o
o6aMSGt3/CnBpi0UAqstc49FXE5a4qKdYtBoRcoWSRKf5s5wq/LdUo8k74qM7FYo
LRNJprS7gM7PnDFdRDFVQiRfAFFlbO9Ehbt+htYgslZsEHPmnHgV6+kuVbx4qF0f
do6XOe1fueMtHHTtOa08zzLWCe5NRoeEaE6oFLuy6xtvRYkYK13dB/8hVKH7yA0Y
s6HprET3UsFhjWtvX4lH3D3hKdi8iSIKq5e6zT/XWvWougZtrB9zTWueEofarCL5
PQJak9xQmKgqlgctcNG4cngpnpdb4r5uvkNjmSi4tizDw8+dnXQYkH0XTYwWSAGI
Y+e2YOK4CQ6dp4yMKZlDw9tOL41qbPcaqBPnJWEhjPvIS3nQZrDTvVodqs82EJRr
3mASLB18/0x1guZiYKDuv5smijo4wcn2AE14Hg5rNqT1rgFaBxTJAyz1BUiBPqJD
wRRAwlftSk2H6xPS0ABw0gFxjYFgk0eTyc4Rdmj6itblPRAhsGNaCBC+NLtQN9u9
DHGmZFyrlGwcTb+aMH6X7hVEjOpIs5LrxVUd1cknyt7JXp2OWbpZaOJ+GTV7TH2o
1QUzTcGIOn5wTYy92AFDCYsdAjGzVN56sh5qON6tydfUDHjG9x6MeFe7EVaLwr3o
pJNIxdWKJe0D9DJInpibTKUBiZi9XLsd6WrYm4LQx1Mgf42HRE9HcgMOYzIFUklC
qD1UsHYbiIx7KkhG4aeSNWgfNmWgRe5ckUWod0yJY7SEYYDANEd+6iZb/j7hqgl+
kQ3J2UbxSjugodtU7dO39FBrdDosrZOc/xt3TZ4jdJP1RTe4CdfVJKb/bXPKGjJC
GZWRHMPSf+HjUzHT/X5t2j4AgZF9BWUWC1EcPY7Ej0rI4nNBp21hzgVKQpkSiSQe
W5WCA+t6fEQoI8RaSlgIw+He5sftXuBxblWd/mRiRzxepPI7lHpmyxWqgiAzb6qb
2Ix5+3CigU+/0uppJpt6UUDP2TyW7y1Hpjs9PfiCWD99BTA/RXVul8ZEQXrqyEUm
gebG7GekghdE7GJ4/WVmk7IaDBZd52RCdzehDaZ+KOt6LeVRHmfMboU9OyJABlfb
3vCB1Vs2xUSkSaNiUe5fudsz6WN3AjiYV4/ClE3BzgEp/t7KSlusS+ft/vVyH8z7
1rpm3ZAkuw+NBlKaTDrl3Cib6NzKRafDhwfbeqcCrzeKZZl8pInAXuIKKJEi4l2L
/ls6PMCEIacMCsFEvVynoeHrXGwTWsrnQFwBcpDS7MWGX6vPtIVcK1IRM2T29yZJ
HU9ZFrBG3qpvsOM5IwnJcUrG5aerSHMfzslHChx3g+wqQoRK/dYTsLNf+Ol6IPOz
gvADLnZJFi5fs9TUbIIk147VkHwCv31e2ufAADS8ng57SP9gex5ym5inbuF2q0di
aoqLUTEmPeZgGSrEp1WLzIE/795Et4XyuUATwFSr2OqNc/1AXTInmzz5176xLrsC
66J/n7wsjfbJjslwOc2Lx1QB6xtSQ+i9fU93OoX727nxsT/bBwPCK1toeCXU/xmy
4RHrqr9qKbeCeP8O5LcDYnuay3aGaSFfdH84WcPQe/B4RUokyoR2ldgRuUiTWvTt
8WoAmZUJbi8pp/1OL7aOF9ClGnv2QCOL9PnduJ+rbkWNEdkXeRLzuvD3buxZWHyn
4MdOA8/vhM+Uct65mfzpEv5cAwxcTih8XTfidt6K33mcZzgoHj650y/HvFM2H1ls
K9TWEUcgcyxJok0GEpHEa4gUwXV6Efk4tfP0a0NfvK0E3TE0jizrPWZYS2MOOFeM
63UrpKwGoZGKW1uPTvERi8wwVNM0DyIPG/HBNGOViJnpIjbfi1ae6oaHdPwRFm+z
0JZrT6k2mJbTXP6XhSc0lMnPkZ7iu8SCK+EczTB/W3Oa0FdHHMOH735RiNXPIdkP
oidKh5WXImecqdkncwsDP9KCHU/3C7sXge6kTlqQUz0XnrwIg0q91XjcsGuGsYKB
Jv6BoZnyF2fXye0GcPLyfhnCacG4dVCscX72Tru5ndy+pu2FeTdydFQJzMc1qndR
v4IPgGa2jIHF4cbCltW+T0cNLNi7gM5w0z8QrD/q4H/o/mjCraomhqNzxBjzgZfy
qq3JY+WneFlxojEWfgsHS+xAPVScU+Zhzwz+9kmeKnhcwR589Ow1UtiCSnAMF33d
JkGMseZ/zA9s7Q87J4M33Xg1EfzfPGkcvVJXjIqPzVl3OM9FgdqRzwTje5mUMblY
WS6XJdvenis9Iw0MXZcco8a9509yEPWrecfW0/4WlHBkhAuEmMqmFfODoS90I97m
0vBDNbCIQYz0zQHN9HNccR6q762NA/spInys78T2ZWJ37s5Gc32qtlujqpgq1dtX
iEla0hAgoIxPUjIzEfFCx3Za+sSS0ubUQbssJDpY7P+Av+A7DboNVZ+5AXoRVUYk
CzXpDpnb1FPcemTLh6w9djRYWdDbD7/sxd7u/TlfZLE0O8u5TYRnIDG1k2t+0HVs
v/0HfM7u22zrXbLU6Hqk22ReEBy31Fw1BnDIBNnDAxj/6KRnC1jrcKKgez8hbJm2
OlDJTnFmoWvGFEYSXEVkUfL0BiXvIG+lqkWpRTDbyO01BYihOTvIvH+UdUekGYvX
PW+RY9/vh7b656D5jyerKrFOD3y9q3+7uDbKXjDDjbbfKDCS0BgUcRQogxFvIdl4
rcZHrOvsPbtu0H8wXcj7jjwh1ESKA6h9jjP+zkeZZqB6w3E7pi+l9/o7VB4Bdi2C
zqN7JW3FRN/VDiYlYqIwKau2vMJcxQ7MkeCWeC/8Hf04wvS93CGw1wnHTIVE5UrC
p9fuEMe5YQNeJkjMAIQi1DOMGQQyuFZc9yB1oBcUE6jiBuCUiK6x5ZwVMuB+HswG
1VhKT4FAx0XtyGnUgoGXmjWdGlGsX07QckzsbIj9LFbaIabogwCKHXx/NyFJ+y7E
lRv97DKQwrNjUveSvhNPUillsO1n+nI8Yg2pbQO2j264k4+iG0o1q1+kY57Hvz4V
He7/eVJqYFNVlo6jJ2XUxmGtLWmk5v8itnoMQ/3svAiLFLStXAHiScRHA+g4dE7Y
/ctD+ETk2ox3AbswisDpvD33bTBwUgVeCYwXr6aIk7JpDJIsHxv2uj0752jYLoLf
LoTsfsHfHfiBifMNyDSTF9MZyNuh8VFr08fE+OuruOX+ZP6Fm0xXvd466tfYCj7g
5xVgPNg9bcMNEHFARkICoRzA6mOc7LovCxtr+BONJUmXa5M9BJGDtNz9EBt+5zH0
PYnxXP8ir3swYsKPyL7Qg8gZ0yt7jF8Q9Qo0wbavtUO40OvRuhvORR2gDcl00N6t
wVVoUIx9OZfXV/2cGkBOnCoZdD3c138Aeg6qBbnB2Yh6835CrUUC7VDOVtd9/wCj
c4A32jXNjr6p46Wqzu3sSUK/rSxmxDzneDO8ZtHxhnosmTrXvqKSvZUGIAKV6t8p
UgJqgY0hUOlS+N0ZaWurO6Q8JkNJMeddytQbJQCMJmv3FJSMtSycq8SazydSp+8V
xcDp0Z9HPJv5KwtisTQYipQ/3o+Vyj6WoQGrzNqfvEoNtZ10UF75z1UyrJH9HW8B
Dni87uQeMovUAGdi45pvQWV2CSrnEaLZFVo5vpd/ZVK5e+L6bDvTa9NjsoI4Wryk
hTLQAgI/PcqR6IKfpxYRJR6CmA598y/boIYNLrPvXCJohu2gbmg+TlAJmjE5hJPM
SAAArB5PPDZ6x99L7W+6q9aOT3PYDXE95DzfaMuxfqGg6jhsPh4MN1YRyG3xAjYX
2ra9yu4/8pcLThf9FnI193V/qCOWtlT//gbIA3yvdbCF+y4RaHzSxgC+1p0LJid9
28ehBZgDlprcq5Qsx/1i5dGSPsbRl3SMOwsvNV2pk9Bo/ExBUcrO4bCcP8HQmfsw
78hTTCqGC3zsO/orjbKzQDs2+L2JhbE99AvSNRysXpIM46OE9z06IFTpgoKK4TVT
Zly1A1KvFUZs2E32cbGzr2BEBEkaKKjPTi+MXFf0TDWUK0IFuEEMwwS/eBMr/5Bu
L3ELag9HKipDgYx4VzElk5gmb0htlnHX/hrDHqOoCGDKzgzcgvGuPlBRqR3fBDsc
BJyWkCXlPEik59DPdtbR8CEsy5dL7AxrXneStEowbZ/oVtuoX7Xf6jvOJE/sPhPE
Ble7ANSbOXnCicExcyMkftPUxNs7+G5O5jJpgtdV/RtQtM8CshPcmwh/GAnmk8Ga
ZUVnnqsFv8JXMnpUaPMBPxYuEBFtYnplAxBgBi/NVloQsoFZvv3S1OoQRjZTFbtu
1acrl/VPMi6jxJMOZgVXWNx19JIpFYxDDt00e9YrbIK7x7qe8YZQJwFVqQUzAqjZ
d47NYKx23PO7SH+Gmx/e8qB50vRezBMUJHHCnyB60XYlhZ0InX2scgfF2PpugFJ+
1Sw5i66EeHQQsLg1+4AduK2ehVCw2bjCdujT4tcPd2V+kkmBkyRr0wlkI8I6whQH
IRs6p5T7FUJksekp8qw2dbk7I7beI0yo2KHolK1h8WcazGGAd+ZuK8sC5aRAHVbC
L59Eb3ETranioRZghBMmJcBfcrYlDyqsYwifTDAG4WDjQIvCTzGiS3O9EBFMMO31
OtSX04BX+qkyBy5yToBoXOXoZqhYiiek2xIqTx2LbrDCrQQmp2UC7HwBQZykpc9j
5j6N8TquK04z4qC7NHCgHRU1hT/s2042wxr5UK3F3C9X9NUBny0vur0kBdRajNpT
52m2KyusA6YEXDshggvN4xfldTWF2ZdYetYy46Lk7Ep+ePrg6sBJ29+SuTZST7xv
iM8KGRz0lEje0NeQO7RVy4TmJ5NoFIX2OawPZEhJeBRIIkyy9dmiU1A57EQmHI5B
JfU92FUUeLyBZndEMz9s3QF7T3f79aR80Z4boOLiiSbSaZZcSi+SsDDnwNlCWnPZ
Cee+Ffnuoi8HpFkCheeK12tRXGYnLxbi1VhZBYarhotOaDPzovMGn9s0J8SofUdP
erI7WW3yeSpI8rkvTFY3iaWzcgPNS6wvrCnDGB8RNei3B9JvmGrjkFkxuoX3JXVg
AhAfMA18XomVH220g3hrDHz/2N7FUnGUj56tomgwsF9Coi8arzqPQZWWIbwfmo8C
LO2yqfYTMeW+kcFkfaJPOJXRulXle8P2uRJnM3iMH3dfGdn2byx/vDm83h4tBoqZ
gun2CKPkc7Nxbca44gDhWtTCGAgN1rHcs3M8TkFWTd0mOWi1zk+4975m1sABMuYZ
QZom+mjWuIYgViVdOJZyCNGr7cok70g8e5M0xzHK1+z8KPxJQ3Y3Jr9rtmbxXUJA
/swWkPBKW4fFe9Up1TMrdp3i8aa41grXjccVxxJ/RnVk20HCtf4v8QmbsD8wdQ5O
J6lP7N7ZyaI+7OYPUltxgtaH0bS+KB2JMXReB1y/AjBjKxH7LQ1uJX+PPIOh0unj
hDYWJJ96zJC9brxfO8r0AmJqtck/sHuo9VoBvUfmhzY7a1Gu3rcAvAKyfyle7nkg
gBsYtMgtJ+nzcb0A6Ah59+Yt1mnfeWR6KbtWSn/8chBfWlcs/yM6pl0vRCJG/Pgc
vjKmTeDk2Dh6rLfC4lifgg+/pVXl/Ks21Qe4p8INkq1zs1AisX3nlgvbtlsOT7NG
IyT2vp0Z24EQJbods8ptXlHUNL/5B0A+FIG+woE2jvdmEJHdKQtHMk3mbSyjD/jT
2AdpDTSxM5M5twDt8zbnwKCQsjbzmgPNCTuJFP1u8Xd2IxfPeQQ6JYFXO7bWWeWj
01NNtHl3r9jV9YvHQf6oTokJT0o+rEYoQ7AcCrZM134gjjUzdOAPOR0eo7wbtKpq
K7R/guydHSqTY/r9H3iZpCDuHhJf29Gw/oOpaS30qhp2fgwx2IEph58lZaRxY4zW
YPAK2PZiV8UMq87gdKzED7SDHYtPaxBPWweAT2aDwR0HmBf5m8lNpl4JJ98mhLXQ
YP303c206J7ne5WIXQe5vFt2GG6rU9AXz/eIkOL2t6zg7zkLwmmvxPCB2q1kH42O
Vs51AX+B7TZzrEoRoepGccfks1KZbSDvJuSu1S6Te80bb2FYlmIrNsP/Zi3xDzBP
y8K2lh1rz4rNT+3w/2t1TtbXOhOdL70k8nTlVB0fZksTw+TiADVL5jZ8UsO51601
xRin/RpamQ/9UuKl4YMhl6ii8hA7ILwowHYzeYgxNTW+SSVxiy9bvGncbiN5P18r
aI1wXA/DEQPet0CzaY6pQ+mL2V3vSvMvFaD1sIYxqVYXEi/08BmF51+QjU4a6GSA
uB7zMdRUBUOSxno2/koX24em3ysSPYQ7AyTmoKOLzfAxfVcm5vNhGdq95FvS8eEk
adFcIQ04TReVQ9YFmHlxhMc0bnZl/JQVwF86L7E36C+OvEhDSs55IL4aR4/eLdSA
xg895FLxPTpSH8hTvnAn8EwiuNZL3sohVN5e455oJp0auVBu12Kr0e+to8IC4XuJ
EQ80oMF7cbrRl9Xtc/Am3PjByqsK+wDGeLLEdwWlWhO8PldNy3Fqns61DjwNERct
Z1er78oJE9+ijktDXSFpnDCSiTn5E5ImRgyRXAjsBULTNaua4y3604fY7+XAAH2r
6+r7+/N23dDo9GqorKpmop0059kkmRfK4u2/RJAjoewqxSVniIJbWnPnUXvmJjVf
sE49WPqM/t/7TsZYl8FEAMLoe44hXwC1L0QhqPsj8Xc4nawKUzfK2yTAP1eW6lAW
6MBQPBooayxk7qgU5LcqJEfB4y4CIxHQT1jL+PL0PrEkiNnd1t55pXam7PR031kh
c+KF/07i+gLyNlFWEqTQ7JSRdo6HNBmkGeDrNGnrI7vvNZhCHownL7q/JiCKmgWX
bSLZZhRGAgc8omU7LKFnRczizT8rqZPv8zcd7bNxHCNhgozWDeMEueLLQ6clMtrJ
ext82RBzC/TTDJIt0f7RcaEn7pCAnOAnZ0zXQ8SMRkAPUELa4l4qNMEmKUy+0TcA
aXENu9mQHJQtgPxtFwtVpmSMZTbgdj493HvN3NDUZDnMV7nS6EElw7JdSt8C+o86
E28BcLhzFvVvpyI7CxrN8nhEmpgWheu6/nJBmW4BfwJbctbOXRF6WkECcWS4DjRO
dAXtz5IKPhZIrNgSMgDtWlaLOlpEb7oah1U2C2hpoFTqiIpVMF14aKvC//AuvgUD
IkifNuBoXQE+r7ZH0L1CRmdOJdamJQUAoY5mC5mvmCkcviKO+9JlsmIYQRkluGsc
7d/wykfQRBSrtTh7gcEQe8oVjSP0cKAdXZc8DAUZ0kiPfprrzuKV2ZX006EfXbWH
12H9kD4m/VnLCi7YfFQ06jCwQyTvqdhiYyVLn0RXli+hTHvDrI7Sn3bDswZvG9V9
9CkCMHbeY6TRSAfjigAmaQuHadbEPgpVxvUCkSnJ8yPwnBJ7XJdNhVSgDUp8zkIp
arDWlm1R2d/Yw0+XIwDJ6q6MGCJ/mpaqoZY5HZPPPBTgOAuedTKkhSJansjzKZDn
4yEQGx4sQMvBnZhQ+RVOD+snTudcnmszwPf2HslllomkH2dlFwv2DVkUPnZQyoTr
zjWogUh2bG6rKVC5oXE8GKx54vpAeZeS8MFHYXI7PeOM1qw6SvLJPAK8LLRelP8t
4JtGOwPzp4PyaDv/WWh2hH0rznYya0lHNaYJtg7eFdSpoFJTjSL++myjkHL84h/3
8IvwS8viysd4nnZrm0tDhDBIB7vNX05iRJUn4qhjP396r1xhENhJDT9/jJskeAbe
LNcmWusYAORIMbm8/fHCkXbulAujKqRxCtOq52FpxNvbOKAkiT/LS5Y1XiAtJFhw
VIqD/zdc5t62IJkVCa3QdIfJzRezXyyRdv8BfBU0/NdBI0AljD2puoOdRyOTYFcs
kE5ZRwG/Fkvr3B7XdjTLxph3uA0KzO+QnLvXTz/jaLgsdyWqQ4LaIUpMefAy5ZSJ
FmShTiFdavmrvICvPHaM3SfqpNkyT2FeZYjebo00SuqM+JJS7J0RQcs7wARLyZtd
C9e6JVPCpwFtR6Oy9IQ/pwRgyda+bstegwrjyxHsAylt+tfYahe5D5CnK7/3XVZv
GxkVfWkXfOL5Mz3wXNBBi0aWKJhMfiojO1sT1wOlTy4dXcxjqHccFzlTZdR34pla
gXSTDvxuXaoMZ05f8SlSRrVW3waHOAouvNZep838o4ez7r28bHbtT0x9YicieIf2
MGZawffKcmvgNeEaMQlT0vb8Z4XiU9E34Rl6CAy4Izg9U+ndT26nvCo6LquqSRbz
vCGx678YrByo7d+6UQi6v5nptu6GzcskbpqTe/3nviOID86PYf22ieJtpKz1bKgK
vCmTowf1husrIQq36RfRm2pyGB7RKvhYWo/ATq58Y6F0B3FazlnDmdf/xgjscBvR
nwvsy3T/S4JqltmFgXQMjCsXbwT8PbqdJZtaayilBXu3xDDSwKXp6LoLXwPKurrj
M93x9w8QgmXDijdGjvVFJGSwu1zqXjmZal9DjvU2AziY+ZHN28daXV7PjXpLHwoJ
t5YfmseO2cTJ59PBPjl8sEFAX1HfID51bzYG/8AikIoq2P0+U5Ilb5ifLJXn7Hpc
DXDIGbtn6+UukNnAFcKHFjt7TsqekSTYdDPtMYgXFEqu9VDZoMyhs7J3FedH7zDT
9/7uncAsxQUz95tCx+oEF6OSBIGZCaPXUz52SIB0CesHrLGF4l4Y+hDz+CTfhd4v
uAhE0YdF0g9NsBNHH1hGEx+y6b3swniEDUSLx6NC8fEBa0MNDxXZln81EX2Lb9oX
tUsWnivviUYu2tJiDRCVRAF821UhkDsW0yPlLdyHyg61lz9xsbz16mAbYM7XTURm
TipIbULHhY/IiqzTcJPWZUi+747GQhzoT2RwW56btSXeFoalR5Y9bA+1IbBOztN7
3BNBK3nG23a+RFTd18S5vvuKEnogJaKSY/924L+BODYOSbfS0BuHXfp7u1jggXVa
ptyBUTC8gvgV3la9563vH+DnWEV6JmxwThusWg2RK5axJdnEoKChPpuVUGRv4mL/
lhsinIqnzeMDdKMd7voaxWVSai640DwS2sYUWQ+tK/Nn3GIIR+MiUk5Xsuff5nzP
D07xsaQnPM3Dw03Vh4jFJKzYprQj/WhfgG+Ksq59wUNmrH1ketSZ2Tq0/tXrd+Mj
snX2q6HgOD0/uCTE3q3KN9etcfhYJAd3/2k4fTbf7n7zGe0hvIR19ftlvlkSF6Jo
jZJjrSOBOKisRI9VbcjXEyNT764VG4ykDSATmGRO9xlKKSBRP/z7U17cjgP5KeBz
bNUjLmixW8zgY3LZfANg3wv4ESgFGNAfYxjUp2RGdzasCUipU1VBdcYc6zPF/gWk
KTJRwYsjrFKOLNyD9hPQsDLi7XUBA7/TEzXxvahVvWy8H1U2aHAW6QqG4E7bt6K+
6BdZb2S5dm2LV3lkR7Jyrt7hAOmhVf7PL4/J2jt2meBrsOTCJrrGwx4Fu3+ixOYe
bjE6T2x/A3Ku+sIXyeSO/3jBXhUDiRtVMViij/4axHWBdBSjc4m6kHcL9of9z5eA
/p4U7H1oI+MdXQ5fEBWonimCnpUvJcm5hj/E0qdznLqBLbR33M2bLESLKYlSgZ9r
AQU4f21vSOYWFSqVwrX6TGGapMMLb4e5J3372IzKS8h13ZQKkzE8WZcKMVpYrTa2
jOBl6SZuipXw3qkZe+caKwJTr/ja+SuVzOs9LP+v06tcUtBJFBYtD3evHolMX63r
a8wnxC/c8p0CTqvtLlEqyXx73jpMmjK2E8K/puYPAOSllyJzhFhEU146/sWcN4+K
S0vwnvjs7Lr0en+tOMyJXJspgkMw/9Fr3GJdac/vJth3BGUmb3R/3Q0LfRH5SOg3
6NYjhl9PHipQDW/Eap7RzTnDEkoVKCdAzGEHra3fr3ZZQuQGd9VZF/teyqjlVoXO
05DslF6gYJ0VVVLxHlQPp8NG5gdDFOx+EVNCwCjciA9KqN44bm4lpQ/xwS+DLtoO
pbfXNaD2wcsep0XONlpyyKzVj1LrFXYHq22dvjQvHUCoaI5AcnoL0/v9TULqzjtI
RIQbpK0iUKAsn3S/cLvpbsLcksUgxs/zwcIsJy9ui+9t1m2qhXr9W5cIjm0YL5KD
+C6WYRpkeU6xqWoH2Slox56X4LcCX5NEXvUFw5CjabssDfYyRkQrV2IvhZNRdkvP
Irm4u/qoCI0MTxmRO9cnbHJgdFRDSbLDarKiBLYvZsX3tNd7N+SdV4MnG7ZA+1Py
kY8MR/yIpwc+tBwH2fYIUlDTyEul2etYDpc0WnyvO8o2romVgUwtHcuF3Fx7OM7y
nNjyjm+kUh6frrJbjr7ewdl2jd/gajjmlejyZ8TFYqKXRtY2Ozzmhh+zv8UtHPOB
KksupOOlBR3QoV+9w6qoMTZIOhOZuhuG3NjFpJecNcUSpLQ2ZRjW0xQ96mT41ipI
pAtVLCx8nXwaTLSP8nWYzCcA8BorhyW83Y25n6JY409gnm8duBpmvaiqkDRVZr2Q
dhvh+49UZ1oUZbqCvVrc8IpDd+AG7mg2zMVjEGeoe41S/raiYVnoMh1C8ZO9RYtA
kKhXwWipq1N2MKVlBfF9pQM57fmHVS+B9rWDJF0BcgIyKQKFBIfcjE0ZPIVylU6u
itb1JlDwfkrjc3Rwuo/oXLMsxZNddjLG/CjZXw1h7OCzkQfF7100mcG1lMgOgdnb
xMyNhdCBUxKCuZdZBocRzzRNSZr3UdON8nD5Rr3q97DnARYhXtwRfnlvSPt3xiH7
Ei9mlC+qKbkTN0I/xJRFAiYYrysV9BGha8TBHEaGAIxLYffcP2XxgIf8d3JeAIqw
5uM0S0Muep4MmuKC2buifE4WSgSMLkyikEdoq4uY6HCCoRuOQcFq9IrmGjMwlIbr
3nQkrQF7syqRH5bYw6D6tv9bwKmJpG5GNwipUqtCxJ6XsF+IWDEXMgiayNv9zo46
q7zg5DGRGUlFZnStWR5Y2YN+tVriD3jJuJz8VYdx3OMYIagKtrsEsZL5SgkFlFVA
ysEbvjOj52DUAVVbSBRm/MbERh8asScCVfOi9PCwzjXsILp/TcxzUly+xbEVsv+/
f2bqUaZH43qVSF5o50+FrWjeQuIm0v0KmtcymHMoJpuFBFdTL+4rYsuuj0Igsz2l
8L05dzRLRthfIhr5g0MwmWAI8G+wOrMqudZHeq6vqxcKS0y56LUdyLff8JX5+OxK
R/m4TET7p3S5ENT2IkvaEapo0IFWz5GJ2HIdXMjRwXzKxHh1OD84TJF9IaPEMBTj
no7mjTMhXL95iLFfzI5RmgIAcwwuzBVG3oMmifhHDRLyLVOROgkvDzI/ti8Sz2t5
LTDGrAx2vwBIg2TMNIY7SPPNjXaGL1TmehkixOMsukwoNqs4sOiXdbCrSq2pz8r8
nQzYunuhgwUwuYVwHJBTTDOhNaAjOIiqBdlHSYdco2UZUkftL+HShwy98+3Eo83K
SsHF3vcfEG3tzd02uu7R8ohrC97KSEcteHJnHZ0gjR5Hi53Uh7GtdbVy9Ijz+ZK5
GvzfVT3h4oiZx3KM6NUA8k+lVtxDDdZw774FDU6TbkWz5tdsXa0D2vR9yvj7mgA4
3plrFyvHdgRQbUm+nrxfZoW0srIRIFsNGmN+kzW3AwxHFFnb9Q23K3n0K9+SIZN8
IwOCN3w190OZw8vP4nB0gX+ppRWEoUeneediawkvGbXDSR8jjN3U14eMheUCHkVY
DjkzzitzMSCf+aX7kiw27rk7/bIpfOoAZfgbRla+63zPSlA9gIxzGbT4s2t61AQO
0UVDFo4OZpM9OAUEdOfIlOwgQYBqbIdWJB/7ypGlLuO1GWKIX9xQA00AitQQjBLU
zb+spFJ0DS0tkK6POW9aPFKVoHAKB3gM0byovunofnP37aV7yMrE4qp5QQFxeIAA
Rv1+z/9ReY+Dq7VV1ThZmSIVv7I89SdLryxj5F1iHeySE5fkkychgaldL7bJD3Tm
FNaMe3tKQhIUXwPLeN4+uqzTI4w/GAJBAZa8jr2qZB6LklNpWs2ft6idO/9Yai9f
LoMV3m8/AQZGFCCfoLfYAbWQ1ma7ElxRdm4+ltVy/5Qq3pdbO11fKRuiX8ssSrY7
6EACDw5bavWwIApsWX5nmKh/D7wofdh1loD0mZ33xl3UXnZ1n70VHekravRbkk12
tdKWwzdza6L6imGscgBgAR15m60yNPaLaobkd6Lvz9XioylMh/4WxGcwuhrJvRr1
Scs2IuB3QdW02jNtfb6xlIX5DfI6l+Y/oAbPlMQqFyAwCAktSg7pJWG20J+vuvn5
Vjg9xhuKuXD1GfyroYO3Cpx4giIA/Ray1wEhxwTVSIg4Opp5fE0XNkQrwqcEAakN
8KUuWVvziJo2+TdS8B4sWY9X5GeHPUwY51iMMoaYfkGGQxhhO3FzfRtNN79BK2yC
Twy2rDCpBzuPX7kPkR2xbAPDlmbdSpp+A86do0jC9erlzAcRRmjDg7MnBBJ7xJmB
/gGm1G/E9NHAHVRcDI5EOrtEFygJToDc/mr5x1aKeW0CLPUx92OSGWpGMgwqcN3P
aF6GwN7fwY4YWhLsHKg2EtXXL63XHl87Fyohd1YsKink2qDmkLs8siR0YiA0Z/A8
4Uv6jjw0mYQlNLmw8j17Hd3N44W1GvPTR3lLHgWkok5cSIp4fY/I4fVY11uG0d/0
o7srdy/5U6y1K+8XjaEDucDwV278tzcXcAvvx5Zs5FbgS3xdAvRrNelY0Ly5EfLs
OK3olbxD0tdokWEVSGsK/rsymHzYxtfKHXtNiPHnaXeKRDQpWQuiAyLeEacfweWo
eh0TGkDeiWoQb8bM8363UXQQLiYPrxcmSFdMOokZKNBxTK8RV9Y10KZY22UEkTBu
28HF30xh3xJVlE8xVMKC0ZGQ93WnTe6IJ3r8DDxEjr++SZq6oj4mMgQLNee0Xp6t
rmxQ4+be/Ni1fC3I7tLEQ7DuwGKXiKlO7NJ9fZwpM5C2LZf+E2o8sGMBWJeGrSxI
Ik4kyfOcvhgBc2Ml01x7+9fQd5H/TkWl/4c4u+Q0qfPyrsqPppm4VjgQJNfNDmZY
GLDSMmWpZ1McurYpkB9q90jYwHs/N9TjNRrmZbmKU7YpwG/Squy2fP5NybjIQX2p
4oqznrFAIp4aykcIyUhSfMtgLxlU94ECkfEDWIztu7vvXdeT/H/jlO1aj/XrWT0F
ZHffPSmy/FgGotaaOOcgexSb5KwhNRAHrxonM6EreNb7325HILEn63XBRCBO5pVm
XYtfH7QsDi+9BypZiE35gSukJt0icamx3KrUrTkHPCZEQODHCceDXnwZWRKSu6Mw
WTYcg/aFqt6Obs0evNzrRKnDis2GQQSrGP1726WRHIibrcW4NQ1hVCFiHUugqFwe
1UCG91f5zXHTK0h2xq4MRXQ0CmgWJ/wNvZF2rm+0n3YBO1c8Fz2YmyY4B1QV2RZW
lEJzKblAE0UN6FxslcWglaZWtZ7fAADJ5H1xtpLvKtdVpDO+xcCF8Cy1xf53cuif
V4RlYrlEJSYfi/EotK27TQX0+UNTYp8wLCq9Ieyu+MuBiRf+F4UPEHv3XgmV7C30
t5Q7EGHXKVhgPsqkFYBR9iQOvb8AcbPbenQdH6wP7D6ZKcXNmyE03tiHAy3yoAtD
iQ/3xILnHMm4hGGbGD+lMU0vqyb7tq5+CxyXVqh7sdNVqBat+LqoKBOAFR31EPeY
jKuuq4Wau707Ef1zlK3SdOACQRcrjYKSn2pnAfiPODJwlOWKQWn0HMUzuz+A43Mk
FSBkshAlw5Jkypv3Gh8P5VRuPzz2kfOWQnViiDsFlJ8ohHLMFiKDA94n8IRUf0Jh
nocKF9rpXpXaHl9L7bbx8EwgcHnlyXr8qmHvML2gLhgw6/c492lV0WUQ+yQ2B6MR
42DAQ6qnOTd9U6wTYFif+GCl5fufdVKzKBsaqeKTklFz+9xSTsZSpAGuNXdls+68
PGlJ8UP5Gh3tfVbxXtasOu3J29hOMR6k9lIu8N+IKg6MWzakEQNlk3uGckG5LQLd
mgmIzeSfJ+2x931hVOMymKZhLem0npVOZwWD1k/XVIWAKIeaSsbUCgRty6KtdXSG
Yawx1k3XCwtKh8XHNgkPqWKFZwG9BgzT1tcdYRUoyK+f1kdirbGgJ7o4UPUNLrbC
PCIc20NGa3H117EWi+6IKrh+S15splt1pLwliQ/JMIYRklDBGO5ed/uv/pJ4qxFO
PMnTA7AVpJdUX0WgFrpHBxT1x04RiUVeckKkKYLLqmxT5leX0RODQnz53HQfRr0J
NHATLVXZnQ85KIuihmsF1uXw5VeGDT6QnRoyiHSQvndeni8ik9/tLF9aQVt4dnhe
vXB2DD2ISnZ0+vKsISYm1zmmrcvu4yaX5cBoHbMZLG6GMhBhLhuoOF7HAoRFmG5m
YIVBJM8FBgbjpeXWVwRtY1NbtOcoTSYNnisFUh4noF0MDboHQKKMtq8BjeQqqddB
1FFDFiBwJm5zbnvmUKMu1nrpuS5z5rFvZkFJOV9QBnTDsrX5JCI9nQHJbWURWsaV
1lImFFXkqHW13DQWokfKvuSq2tHzavTF5TTodCanMF9X4cijVsF4/H34d+RWJILs
ob6UxeBsrAZco8Czhd/WdxTO6Q/NPOv22R/n0idQqfSkUceoscFPgdbIhpGLCjVz
qov9M3kwsASPbynx3yVzUJPRFxQ6Rl6pq7perP9YkcrOC6+ZzLzYOmXxzcX6eeLc
1oQoburu4LtIwURwO0Bp+VkzvM3BhE0DF1ZOiE1209+MMjo6w2F1vrCa63E91sw6
gJn8eZn109veW/IALYTFXwUFbUSWI3UclBBx6zgauldgguRgwEyYtqM0m/ljGsxE
sqhZfnriuTwteYtelWan3p8bcdcHDRjysxINW/dh9OedyH+Cn6greAtfZ8fkl6VB
LgomYrH742Ga+pSZhH9ho7bpZbDSYHFQj071PA0k8/xgjNBe6U93qMjsWb6j0gFf
VaryyrKVCfASNQoaDxd6pcE/PmD+IsgjFmitawXGVy9b/aOZlQ8Xs/Jlqz6n0yhi
loh+klXzcERcoUzORVrXSN/UpOpwxXx/7YDYDXYRU4wouaRNZMEVyOFT364AxzMg
JYkW+5L4ggD48NFdYuVZLYZl5ft8TjQLvcbOtLAWs0JbFFcPTt7GcUIcIXtD//Kp
stDnq8X9TeFuxFsMcZXry0nFIAm1egKQ1EsOjf49cJwcdVrG7A7yTs3B8509FkOa
Oa5dVlHYCUjziNICAa+lfBrsOOU4pSYBm/GU3YmSDv6XkcWxF3uahcBRRsDjhi/V
TSIXkX/5VEFjFPDyyk+5D8cTvvPQ6NAUGAShY8B0xTgzadYI8l/1zqT1f7Zy74Wf
vhVFGHNrC7RnKH3rsWFKF8lO7C6XKyGNEBuXY51MexMKLUhtFMsYGbHD+UZ/6J5u
2qrilwCkMw/O3DZH7Anl1VQNFvNhzDJdV60CupzWxUpQPooB6jJGTSMOQJBCTeCM
TMkchEnPtorU+t7QxRBjUoiybxo2pbAUJIRry063HTAmI84dMqaK9f/KYMLTba62
vac1/xkQtdVZcn+hIs7vGIla83sJ3ps2SGJbTVJbTmt55hngovV26d5+I8Op/dpn
ScZeWtW8V25DcWfIxw8Le0kpG8vKNxXFNuxpPwrhnan2MGCM7W0lQlDhognwc5QP
7LNKDEoaHPrSU9JO/bAYJl4pwN5EQBt7J7FGlux7YZe3qygQ6KoYDhR4iJVvXyoZ
mhQ50ymeTgh88NSRpkQ9vLu8zgAuRzhxW/LmzCnNcuUGCZtzwXNvWgPirz5WGiZS
o+3R360XPrz6o8dd9jwV+s1bmZ+vl2uLftJNyUFULG+G/MtXa3kJywBYclXZGTY+
VjXji3ti0IZFqC7rPiJlOFbltwUy4vMQd7kaf3im1m8A22dM0LVusjZRe8a6sGp+
eSjd05X3ORbZkOXiRI/eAqNs4eQleV2F8pt6AWLj3Iy4L7tQlJ6SvJStEk5Ja0g6
z6ub24mvkxH4Fcu2vvs/usRmW2z5qoRN6Lms85qnZL8EfMvJPKAfNecjBKV2LGx6
wUzwClB27CcWb2OWTuKJHUUjz2AuDqISmvKBAIKMDRiFGtfJm2GD67NrpAfMad9r
mVFpI2RsecM72sgnaRQkBnoNMMhUzQQq3/CsUdmQIEEv87RHQ4wDbX/jqose3U7g
aBJxy6VVFIqvS7nut1xt1KuMtJqoKfZ5jsCMTW9ncSe/JsONm9E2uNp9e5LJErz0
TMtD5Aw3oEKe/K6nSqMopnPDpFN9dmZSYsq6FCTUnZrdqdff+o/4lNYOGbqq8YV8
vbU/fg2heSQ0rorMgEApuueo+M2suQW7EyaS03R4VOAHyE3lt99K5LVVMl/m9R4c
KH1mmvf2xxjjiAY/PvooL2Cqt48DkK05cr3fAaVNmY81fd8cmEJe4sZH9BxnysNe
1ZnOHgAm2u23wUWqSb6d+0w/nMteQXpOpFXDaM5pXJ6dvpZvP5Qu9t3snlhHQrjw
G7AC1G2yMCNus9HSj4qeLSCMnTdhMpfxGq2ZqOMPYGwJivapfCNcUhCAnjN/XjRN
+jacg2htzERuPKenxf02YlXxOPlIEqrnWizZtS166za6Pkkzngm+Vylz+Ty3Ii+n
hPJM38uMijmmPTCc1NVDxRTWEDoMr+7uM8NBPuo7SW1uTA/OGyFpxChHw9ZbwLeK
T/GKeUx678QNeZWFEnjICiKwKYaxg1rvpAK9PXhyzASr30hrieE1Fs546h6ItnM1
nn0Ar8YvoTN8HVMudCInC528hWgupMkCrn0WFK5fCeREGiQT58T67DQB2zVdn/Lh
VPGx1LklJ4oqBvIAnXD37AJuS0E/ubUEyUMtvwNPyD/EiZ8lITq+MBL12xNeFOtg
WVxSN+ESEq5ng1celjrvUwQMC+j6eUP7ZVYO1QpgnirU4Hxi4Cv75EZtm3lPAXWx
76QvjjTveRIfMgzSkrZ2PdcdhEfUnc9QT7P+3zsk9iu7WTJtaSOhcW9YlrfDcsL6
XjNNad6lPLzxvcCB6nwXGMhRmsLgNgStDuJQlJt/yZWdOYRXQyGD47YV5D7ZZajT
uA5ApMQbS2K1qgQH0kNQtaRorr5dgSJSdoy50c+9DaWgXzcY1JKUe38fs0r0t19u
/BlCUA4bhxiAVy6C6s7juZo6HU0VPgHUPPJGnJvieZixiZ8LkRs8SvBkWjPbN65M
ImkBtumqP7VTKjxArKvr8T4f4jWtFr8I9snU2JpGK9Su48xvPc7OMWXHQi3cxQdY
Jp9wJ6gALCBEr9QYPG2FxyoZY1JNVcJiSmSyPWkGukjP2dgptJfhQ8Hj8oT7akw1
pm7xrFMqGRC/fW4Gj6+ppAnumt+C4d8BgM1nDVXff4xWxG66FScpZLeQ81Ec6IOp
iUVdpbDMDVEbTs6axQVdbifAnVlIS6Xz6QqxOOJNijLEy3aJCULEsW4WgCKAlh23
kxZ9PiVI96PkqaWvH3sCYpKPuhVd4HN8YMh99hsJTAtrT8ExYvnWCn3Fa+pTgZuS
1pclfez4ViQ9l5GZtHVjBnfrjmKkaVY3evw0qqKnGWW892POQnOIAhEkdPJ6MXxb
bKq85s2ZR1FmOhELxNMOVWmIGVB+4Z9yvahzsBtOKprVftm8zKkfJJgcCwXxVBt9
JFXg8UU907b6NKRNAXTzSQvmswr1Sajzj+es2zvG8IQTbxJNcuqlcPhRnQoZnDy9
HFgW7s8/SinPagrD0SIb7rgnvPffiVtP7oKEwz8qoepkaDSTzkc2topr+sjiNN5f
pV2shgFwlwp2SlMHEog0qEZDl68th7kXPhKP76Spp/OWK8SGDemF0kKb2QYLhvoM
sP3PaLlqhLUmbQa3ulfGUthpjKM6A9rwr+R/eRkSm7Io4y+GZVpVPCHvL1mKz41Y
M2WApjWAbp8gqORpHs/zTCjnUJFxb5zqcaygUr4V6tpUqNvkFzY0STMWA830fIfz
qG0ALEA0GxmDWumeW/hUvMlWWyJ1e+R8aoRUjQLBt2DXMITdbIl558XQ9dMi8p4C
OYpW9hwMOOVvbUygszUo4CYHIgPyVR1amSgDLvAfT8fH1NqaXvlEVDy0sfoOoxZT
AXHOh/4u3jaJZiJrRYRQkm9h63O9fAFqR5+NmuQLpnxTUgBMwApaojC2CDu801e6
9QU2GqAzMHzmD3cHmP/piZAOq1CoizpYSUaaijG2H4LTIdV+w7ACY50SQ/7KKWCU
dS9t8+OngxAOEoMDZjWeDHO0/oVMbpFv1wQVXhDRXk4EYGyR6h4hDamglA+QSJSM
tn4y/qbBuHShxs1reU7bNbkO4dZhCRzBIZsrRO0y5LqW87CFilpwl/ptOsW+46Hs
AETEi85Mi/NKmL392Sol0SWG4w0KCRqGJCtPtJryGQKN1htt9nbMy4ThhDk2GOYx
IUb3b6+8RTy6YQ64a1zQI6VEbYe1G26rVGiSj96ubY+LZYj2EcOkYFMVxbN1NzxP
s4SgO5dqkDTSBg+XkiJdmER9HYqCRIw1X69iAte6o33O5dYRQM/dn4Z1qDOKhj3G
ELS585/z414aPrvSWjUIHfNZ6oqOIrgnbPmQghDCxqS8Nd21jwhLauLXda9EXEhr
EjNLL7rP3XoIFklZ+adbRiJYnrV67Cpsp2lay3b2ZQR/VXk4w/iI9AB48OpIHV+v
kXkI2Xtcz/k1lUwDVwyFAOYAxzSp3oXKqNAjJMYysrPTwaDc4glRGx7sdciEqJ0A
hf7Rkhh1r+EvjLisQkQzk6nzzw1POjSfe8swFjCg+dcEniCJPMCq3cAsJQ8irUX2
mqo3WOcLECTZvsiGnLt45XW3MZKLeHLyyfemoqO1GbI4oVVQcx7GEHP68rpNbhkI
PwFDnZfuByb95mjBLvReT9iYaSy5AHWU15tlLvjXRBBeesyLRm+7YfI+JcelkItj
fD3d8dJjEUdeRG42LDN2PQoqLFG9lo930xGedGYMe8XZu6CWOjJldQY9jcONfowe
bEYceIb6PPoUZy1IpvPh10jYBJGgTVy0/sTvrXYR9geo6z1HRS9/yBlquhJJZhe6
k9rtz8mKHHdXzWDHcYeb7SIyTvp99w/1FoCSTwc7F9eN8jWKvG0ZiT3zKDwWKU1l
bGweJwyag7Sc1oQTXGzRTgqvYnYTcVqGlJQMgfoIA2ht3y1YFShZccwK3XfkXvjX
H4eXyj41+sseCXWk50i+XRXhV0/jk03lZIOJU32SNQJIPUBHnP0VMRPEXPXtWRCU
5NrCZ1BBPXJP8Cos6BxZYO5U/2XeLevDNnPvblFhs8z76pbSXDfo7gQcx/HB9FHN
ivA+ql/oosrcB54CCilTfxNQMldObNfY2NEm4iho7O5sR5pLjAPBhFZpZYRVLtSK
VDrVf35/kBgGsmM5AHT/Ed3/v8kYLH/IVJORtol+8ReW1eHgpX/tnSwlZJFRbO7A
qxonJ9qKA2/eKUQTXx9qzVFoeTSYdjg0Ua6JgRecY1lLAjsNVVAou3SLb71e7Lqc
c29RmoGHyF4UIF7gH8lU3UG0mWtJrrlm+tM1F3sot/v1RRM9rHRGv5p+xL5X8Lde
SUuZmqPJbEifNpHJ81iWQ0Gv2cK+GgtNcin0pk2wedjTAzC+lfjiMIve6QLtjs+I
T6eP41wA09HjE8OtxfGJtcnAxtyDVg0SICCPQ8A4swO6xWZS6Mk9Z0pjg3l5x04S
UwKzacNNCz4wLXnjIIomEsERBeVyurqqZw4MUQqNRv5ctItGkHbYiMm+arCd/EZR
I41ZoznnFqI1H6NN4tSKfx4waa9hGZvuh7tvgbnOhcI6f/aqhwTFTp3cTK2CUp0C
y4PRqEjFtWPmWqC4WLlj63Fn2BcqCQAOJYlFcigWdpnZBf33EG5U1omvsjuaFeX5
/WcdI0YYaSu4vMWHnHOaHUW8K4RpE5ufFisBptwWUOYIORckditz0QrFra3cIz5s
qZoGV+U1pusnKYkMVp/ftIkEqFx/mFryQPveuwkCcCKtw/g0RJZ+KAmaf2rWJlMZ
wkqtCnuXUbEr2z+n/q/DKtDAj9vOEg8pLQGG8/O2A3eN81+bMDhy4VqWKDv4WYGj
itM59yjNzXs7lwVf3zdzEglcFG0FfO+c93JseDy69XzcmJsGE7laaus8Fd21+Mq6
DRipYmXeWAMnmX54Nn4mkQmqotAHHeRUxKBKCQ4CAQnU1R2oZF8vBwho+6teRSyO
Cyo7SYVVbHMa90AeuP/Ue3MxAF+wdOZ2c2/O3wsjXBYGA3ea3oheEutjeJAjGuRl
5xdT64McKN6FX8GLBUkZ2Ap/e5ZGMm3eiHQR624Y2HkVZW6JcGE1lYDXJZT4058n
xYHBxA8L/iPuu2FtA2/qZJ5UBoL2mOtZ67nCanbzgr7F73SigJls8pmARvBstyua
CO4ScepUGzsJRGcx47uBTMsPMoAZBdrBqABQMH94q99H6vJeJ+CLw3AoeMONzSWk
BAu6iLfhdJRFS35QjVhwA2LMJJ+3Wkg/qBbQUHfRxYPnrLPda5UgmqsKG48pIK8F
uBAeE4OmwHZ7u5YS5ijVWHLUghj8NDe32RP2Eb6gRp+dvFypTeSaearyCjLRvqx1
90bQjmUzMO1R9BPqSbOKyKSvxJHBuAenuJ0gEh9rgvQ+P5zPQDsazIG2Bc4NPyrK
iiLCfPBScxSSkRdhssDC7jD/Ld+pkWG0EI46h4wZMFNYEnRmwgHGoqFQMPOazQ0s
SWq+dKQAbYnT8kcylUYU9jGBEQAvEwfo7i6o2ymO/pnNwtdjcSpxV785s9CUeyIi
ViYAUsV28GffZEBLIn0y5ajf3PJroOVFApJc94X/uTYT9LK0kp3pGlisZTbkWdz9
L4U/XMYmn7PB991Herj1II313vMupy7Vee/7kA2BOPQmKypqXmIbHpdfmrgQVhAD
IHVwPLs7JwygXlCxc78iEmHrdJg42WbPJ/Nyj0l1xgBsTTvjdOYea50ntnXbXPly
89r7Dr+xsk5cxWif7KsmcfWJ5FooD0Ru+uJfEEkZrjQ4xTJfx1KGptT86p7bzoaD
uviZBI/yUyv4nlvDblT9NTYD7W7erlaTGYdvvgWjwYs2ESLd06/d7tuCU4Yn3RGN
Bju0Vf81DCNL7lZcjAyIdn8lvy7Sjw4887CJPtWfPF76ECPvYW41PtfdmVOQBvhZ
GiEKVWOc4SPHCRuAE3gTlXOAIMpEH03phvu+4s5751WWm4mUEf1LlbkVmQecu67o
O16ST+oTNd1JUvTjwH8ZjriZCPF+3oEvKrgOcc9iHgy5Wp801DWZlaA3DZwGNO62
CHsO06BBpcG99oqwbeGFatUW/bKau1sZXxO8gzxD/b8TZhpMi2ZiUxg6lAAkXSua
mDs3RwNssgIrWrFdXraUzQZAXjtp8chlC6T8b3HRPX3uCDCyUp95MXuSu/ZSLoWe
eZGPgV51aTOtDM5eYfTqU1MnRyGRNqCc1ph+Pib4v8+6jBQTIwDZ+QEBwuS113Kj
obCbV873JFQxX4R5AHvwv5IG2DXKvQtbA6FjPkypxLGLWU1J1VHF3PW53M8cCmgk
sUsbr3QrEnxXkPU71QaoBZy+UbjUV30+YHUBRczBxlvEPCa4DB7glJIbGmKhUQub
gbG/H3k2D7dN0wvnIRovX2QEXT1oiIp9yvyHxKhQTJCWOwylOfZSn1gRsqXytYgp
+hobi6E2HLCmHY+HXidZtbHAhS2iO62y9NqvdQBBkoRM37K0KbSJ9LXR19p0d+Bw
sHwH2It5Js+E3ZxpHU+bVwUdNaUrEyRMCeQaPZjYofiAeGjcHsH1Gkzd9PxxEz0V
HwMb0o0UqN7ZASOJdw+PSwQjsBUclvAQL7hbFnIyc1+CFE7OM9ZO7LBrENxZt5IF
vnpUjRq0WsMy+WH0VaJAgXTBcTEFXScGES+zMnXxJvN76JjRv7Xrp/OjJdE/KMBT
oCUChKcpfN6U9dlGnTY2Ffd2qQp+IMiLC01vbo9f+Kr8HjwSRIGE5TwBDhIBXZuk
gwCNaZgpQu6C3w52Nlq7+dllwo61c/qvmT36ZtRpslSZP3U7UA/gQT9OBkzEaqS4
RDlk+6Su6FroQb/vE8+mCbKgDKMTA6hpKAS5hcjbQv4JDpS6P0jYQiNOsiQUtDHZ
U3eKs8EJb2mvXI6CfvadQELT5PHHP8mptplkxhSiIfjfgqkABJf6FDEE04f9TZcW
jAJUYx+Y+qHAgQU3K6hT05Dzn8sveu9r6dTvseY5sf+Phii6p4stmRQq5vx9bn/2
xmiVTJo/6/m7b/dkzUw5rG1VWWv1cZczcyY+x+/2Y2rSza/ppL97DKH5l0DHYTdd
VVjlcKIBLVjhA/paPiIBo8oYIUvAyt59ghlhNYD6UzUO0VKYI5+ebym9qohc+qJW
BC4vEWpc/c0+dzEGSJRhUUAx5CZ9M6Z6gBVeM1n9qee+sDX2VXb3jw6exbP0HVx6
m+lDq0YioLeNwoo6nOIyih/dh90CHfs/6VSbojOSZEwVfC3D1Lp1LvI1l4Y07VFI
w9k+NuzqKteg12+YC3r8VwdmodUP1e+6fjXjNweRpXczwxaYtMwre8+rkfgkqkkf
X2Gm8l5Sm/Yl5cRqJED01Y1SSmC6ZMCSZbzbZQ+1GxHqwkgPon/SKYqpQVyGOAZ1
LFIt18kMJWh8PKuw9Uvsy/NAeboRfRMtrHc+t1BPXgRkoQdTla6beVfaijskMlpH
rnbf+xeMKnv0TuLWm7OvUqD1tI5qHLFJFp1lrj3vOlzX3KkWsbf2yk2DJFBMMlri
M2TvjIw1tBXGkGjZuQIWTtEsg64cFP+A6S2+xHYaGY0gFLLEK58r81/5BigmDxdV
qLfBtp8Q+NVDtkkQtRwPAJwBJV8f0hzU9JdCzD8c76qPLHGpSCfgJinQ1vMUzP4q
S0aqf6rIdmvq8lFaPZr4fBis2YmbxAWm5ES/NpXepNo8WBTOMZRLEu3MYAhQ3CRV
XcJzB650MUz9PpZ2TGAH5b2p9XCtSOe5t2Q8dISkw80s8Sfcy55Uk7buM4Iyve1n
r/ML7aFUWcno0xqgTAehsCgtjQmqKWAyLkelFneyYKYqIA9rNt6zQi2Kuw7g5Gvn
qNRBB4XwICboxfoK5cWi6nb0oR+p5CxB6mNC/YSQIb65uOyldVuhvGquK8E43Nm2
AITMOK+BzHXVKj3+zn6r2ihC6OV2rXl+YongIEw4tZM6425fqeamTu0wvZ3YFogL
wCGeqIymUloL1JyQfEHVvZcGCmn81UFVyuUhTvICwjsp/9KPmbEqeKFLeAuCtVUA
i9jBMe3SkxSA+k2j5aj/Rl2m2KoTpN6Ewy8bEgZAEQq+I6bjbgM1p/r+o8FBX6i5
3wDxgdO24def/ZREoudrZS1M10eiEN05c/hzs+ninEBfqkUOei/R7oZrtMpzY+qH
pVxbhf0fsStI+7Wc+aHypQCAQG3WIoAt7Z0dK8ut+HKy2mbazbI5c6FEexE29i1b
dMSGhxwLGNk7jNKKXUtvY9HDMi8GZeX+jznvFUqoN/9Sf1enW7mJvqiGPvYXqc8q
aaPB/SweA0wGZQQthAG3mHXSwF7RF3uTh0KKbPgrkbTzbFSJM4g6kd/TcAXeU3g5
7BqxDZZVRyjoOZwMAWPzs5lqciQ2+cq8hxwKlvrRYB015qTD0mYAqzlsnfPhcL3U
/6uEd+UnHLOmHuaykzBGUAY8mjLnjqp71yqiKjY1YyVyrjRJyin9yAufGVHb4tU0
QF7ZNFurzmtcDQyrxrONvsJdxYl2FyGJbTUDoUHBlOXMX6wXrI+75dLHLc5EaOwn
3ypazZweTskw9I2nkJnWwn0GT4jOf1kmkmiqeOgwqj0NXHGFUu6us7Ill6SEA7Gq
LatDHvSckyW6TLlCmGkjkI0Q6R05Ph3HUOOOKtwY9ETmjrPfo/0tdqYmRCDzRJHp
2TtOYuCsErz+S14HfMh8Gx8OytP/lPeQitVmoPnGzXGMgBog9BstQGo7KKSoQgMf
p7RNPUr3mjdcStyh4wGRhAjFTUZ4Ro+zMraGXpl0XYjf8AKvILGg+tJJtutV+KoQ
ijspAWzEjxWw83jOq27qeqp0y2D64z6VKpFChjOdYvAp/WsxLLFcQVD2kTxztUKx
eqhSJTz+WGhnBxBGYIjU7cgU1nEXGCAsctq4cu6HX/bTu4/RL/Zmp5kferOBKRHg
xA72wrYhrmUD4mPgWcCX2cutRyYXi7NtM78pVDj5YMQdfZlOUqHKD2JRSmJCiG//
CNYoLyU5JVLaAA39wNdHynealob8VMySmR6OZ8I0ip7eLulOC/CDIIVfJXGHiNMP
KhPXVg/64yVwXEnoNs8MnSrQGoGVw4d+yRXYTS+YtrxU0qLBESohzRRAgclwPPxl
DdgnqGfIVnLHI/8E3HFhtquzeVivFvk7EKAWK7yLYByT0i10dgxja7wmEHlKdVQG
bH5wEVfLbIAM7NlIm6tjzdiMJItZCAEfsEA2ZEKWSNf1ZYxdXQqlWfsAtA90kxu+
QKCAlZTyYWB0rE5X0N5hmzWcLhP7o9EiECdYnMDGhTrpBII6HyUhVk3x7ORVHTt9
Y9Ml0FkWSNWwxEx2Nk+3imeEj9Mjxv9mGcmtPp8GEh13V7+B5dOceAkfn63X+oLE
/Fgzkd0LCbcnWxRjRkgnfO3IT0nGi1s7y3YlrSUB+XCZ+Yl/dsDu4gXB5lJrhkaI
RwYgXEcn/XOoKzEn70m9V9aBd4bGyX+j1+pWWilH8DlQqQKpPsJ5qb6cKTBTGr+d
NsC3huPLGq57lpivCRAEghFYWO0yzrHeMvL6biQXlItVAjEz42sAjwMCsC2dzFJA
kyRV0oWVYkAfZGFZZXgVilBVAl+4r3OCBVtCubpoeAeyAiRnz9Jkc8AKhflb6CNY
CWolvsbcciJdEfUYFs/fHlDLSV+twkcGqp7vwUhUzuKAWomMAj5RutFYy+S2Kt3L
dC4f882gB+bwe83OXg53Iz42jDH/2c9LASrVxZ5RXK/Xpj+DBEJL1nbCzFMK/7QB
jp/zdej/6mizokLiGDxBIcoHtjFuir0jFP2gzJN7Fk6wwJtPXQAbrcyc9t0h1nKg
/laOZK1vytJk4eXJPZjQkDj7u3IpuuS1ZE9yFE3u6OxBu7M+BcvqvWWXm/uIyMnV
kXSeKMQx7Fut4ht7ri4XM2bAfplDtjN26g8j3dfMrty3TyqtWFTCmjtRyWgqKGeH
XugxntXHyhiuV7bGi5jM+WfMzBEiXHJV6/StIQ3alSzUZV6qvpbjFFit+r9zA9Pt
qlxLoCJualc6jhBjTZv+3zkQDFdmtwiZZWx+vpWT7NeJ8YM0YZCcBYb9/6lPZQqo
pltmQs9Zj9TyIbUyu/su/sEM1HAnGNLDYrEIVfUaCSA0AnsOWauRhY9TiHu+LFZw
A/ClYEZV65N4b5mR63dXKT7vpZTeKYFtKooge2/IEZNnqJ1688COcs3gNfQw5Tiy
Mq8Jw3XMjZhRdFrjkQrYddhf7GNMsgjHN8eMpxUovOlI+xwJDygXslDxGW5ibK7K
bKtAMSwlMCg+uymm1S5lMVMvAq1/os0R//vynkT97I5IOGJY3AamsfeQp3JuGq10
kZLNos1/mKPbeyxLjynjrkyCYq/14uQdasTjjs1Hm+IgJ0QYJT/S+hdrNj0ARAvD
/Y/wEmm/eolT8kcKs1ag1N26FogIyAB1RED4RQ6UKXoL3jwfVzZOFV5dV7I0QJrf
3PQcQPVjsFn+KbxNr8KBmkitPpU/fTYlx4YJdkpGUxwBXsbD8/xWH7U0u9NBZktD
H2JlDutTKXpz6o6Yo4DteM0QcsQdJkEXtIEMRNf4AW5ZrQxy7yVs5vzVdK1ClAzO
/JUBNqDPGbm5D9Kh4HLDOXL7k9Jsdr2jBXAsj5RiAi9qAOnWqNbjihQFDwGyLB+P
3dJQAQdBxZ5CFimvqOG+vUIadci83MGk78nULxNLpoVJtyaPPsmGWMpNiT/A9pn3
Su2Zi0nO74MBbdsBE+FM2jJ7JRbXHYddRQwjlievmygXJ/3IKP0lSmKymIeS4G4H
gZLRlzl3m/BMDJ/S4eBE+OfLk37/EjIh4q0dXxOxUkvLmb9y+6rEnDZ9INd0RELX
A08mf2vK3q3BfQidcDZUypnGcIT2La2G29Wd5CbzmgBiJ+6C3yNGCyxeVvPwXNlW
mAQLXm6iHisuIulD8JUBTPnbXoShZfko60PHvHNsw6jIIZPx4g6tVkEgtEk95Udz
adiJYiHdLzgL4Ng/AhsaRUcMjhLpHB6mKs11UWaHJml/zEQEHYXTPQChXM+b+o2i
15AwxLIqhHz9RNPzkYibYWhwCmWGfbpKSM8DaavVWULAkgwnL/TpecVKh6mx0+Wz
IzIBfs1aUY03QRdn7xNX4+B1t4kLAw17itA+2mJIWiliIBnpMcO6LXn8gQYQYWDI
PtnZeUgQRoidFHVwN/5zrcNMbItC6elt9urQG63SSHhrQePzjqr26+KxUii8LSOp
Dn3pZstJcWM6G7sGBxZA5OWC5nMbb0a/rzO8Uts9J7unnK3x1enpWqRPJyHpM5uR
bgg7eSkZbFSTHxy3qRt0gOeUNGJM4+c1aNzm1QOqWh0JXWG3/XNBq1jFnoETcgNU
TFw5LzCpPtoiHZeR2TjvV2GHb9Mw8Kasa/akkQgVO/p59vltuGuOCHw66JwPBNb9
7fzJGC+nlxXbVNNvb9A82zfXl7LB4gGPaxqgukQLg9iQuYWzq3z8THIaXqQ1cuyE
apEz+a5gXm/wdw4pCqr5PBHvoQC4LEMxFmN2qcJlV4DAXaMvlFkot/P3Pq4ZblRJ
wI0xXIHWwVlYB9k+RCkV/hQlSTfcOjQAyxmV/ErwCg8WijT2Gh8qLRHGv58vuH7m
riXAYcr0ZaT6f/Jgw/HyNNK2eCmA3Zw3l0zP8vJGMBXCDQ2FGfT8IwTCnI70erFE
KxE1Mq50/YU8wBCUBWzs99kp6F/o3poCaU/Z3rJTnbjECdYtPfE/9Vjii96VI9ew
RGnaGSj1v1qPPw/FA4LPS/60kf3vY9QPhdIySrdQdLBqMHQ+sJfETOWihCJRRkiJ
FVC471XU8dEsZIYoC/0N9jPagOwh4+iRwz26YV8hJFJqKLM0DLrAaGG4rsYAVpls
wgkEc4k7uOCPFKxgWg59u+O5Ij1VObvrDtrKNdkwectqloPYz/V1HMyXVtol727w
+bcrJ0WQqxVPM9Sc6Lgt+UWN/4MDwU0MzbcuyOJARewjjhedeyav70GoUsrOSwME
qDyIfayfpntFFwcQmqDpGKwLB0b1SKut01/fFNgk96RSybJOMEvKH7L8670WmgVC
5PFeIm6SPuNygV7o4iiu6PS7aIGeoD0TxgHMybI0+OPvrwOdklxpj17ZFX6ysD2/
dOmmLlwMTX839Cz61NTqOvF2lyms1XZ4Jj+d03v4qqFQjmpA2dqsJle4QKCK89lB
AMQQmU9ggLeBOnclN1TNmYQV6UfhVI2IailAmepYEHdN5Jpj4EdYGaHAXzS9WKD4
OHjxpbilAiy3u5lK0VqLm0/ew9OUDr5Drqgo/7bFgE4hRU4Swfhylb0rExiXzScw
2ro4yGJ3Y5SkY+4O5goOycxCf7cfhy139qQgIXBzUzNd6O5Z5rsuyi/JxEnT60mZ
K3iAgNDFxKvkjCL7FQdGQN6C7YuIvu2Ih3D841sDRIJSzkStD4tSSb58fH0s22rk
ypYI8TzOm+hmELh2JcN4B7lYBS92Y/fXWLPqtKEyY782pQ647lVeQEZ0mhXjuf7P
Cskvnq7T9yqzPvEQwyEOVzRhcFZ5NYlCh9H837+6+XupdTfOEKoV1iaIRV1z6w5v
oUTASld7H3u+bUKdgkEpf/fbOjcuEJ7e69zflGrzY/CVLqsm8IMCZPpMOZAmvFz/
TgsIGodNoRWPCLDF0qpjwKiQoxl3lYMGou9tqgU9qoR9GrMg0QpGkG67WtNiUuYH
Etq5hkQybCJZB3LmEmO2VhcQ294rlYoAeb60Ykk2z8PPRUfa4mt08FxVdLFbqwfK
umyp62UCW+0hTR6L8RRvUUUjXuc8j5JDahVCNcZanNDKYg9gYDyaYJQD5m2jRrpn
9SYfQN7Kzap15bkD2b6RjKElfvgKNvQLNYN1Rmma5j2AoV8UXdu681t+d/7FzcQc
BEnUZ4cmUgU4GxPzp+HSDLrzHF6V4FqzYlA7eMnECj4I/xJT5g6GJg4Sk4tmOynW
nH+REE6aErI5e/kfiuP8Dm6fq7C/9406qi/SoE7W090M2QEZvBfH1SX5E7h/q5gR
9c9EAwnbAPWgJo78ISSNxiJAAiBEDJ3l1j4Io+I0YMhkV6Xyhnpw1/BZeqPnJUhQ
hUj8IsfJlctJFin6iYDURvR2Bhau/0/+MIgZqGxCeXV80aWlmlMIk3yBmHsIrabV
ILI178dlDlyEImwqjZQT2zrlnaNk3IQM7NwxyGgGoDFTM1Nf43Tm/mh8TnQEAtwv
kJ6bZhwMzVrqds4i5uWPdNJwL6UIcAnlzTibL+tIsHnHoWv8cGXAvmJT8yYJ8mU2
+H0rEmYnF6AW3+wf9v8Q2w5Vtgx6jY1UQND8/QAgktEVdU1mobixKPvJkGHVfirW
WXWMwvcmZOQCIbEVPY6fHKrxdid6/bfHMA5xAzonjqWpTjMvK3nU9vTSPbMqtyha
CQZ/NU9RuT6MR0SUJD7ITmc3T4unMSi2LYguRVv6+B2NaVk1rLk0sjTXXRMOm0Kq
/MxRGP7zSHSHyuG5c4CVFJLHBCSuqk3ub2u01oWGL9erjl6CUOWFKQ5OGi19l+iB
zwiJ7oD9AiAXtgO45oEFLg3858JuRVSz3IQCmRINA7U+PXlYfAEGCLNTEJX+Szz4
kFEewnAZvjEIUoX6p+wZ6IkN/8Ey/nSwYTC6xOqG81J1fqR/z41d/86Z3+Mejudh
Dz1zsqgQur35yVbEkhIwxFqOlP/bMM2KkKY/hJ/9HdRCP7k+9DXAJVVtxCiUfGu0
wznx809XScQ7i7L/d509GBQNReGYxP7cwpB/KHa2s5i/nCyitO4XZTe0BfXUoJih
QGLXVrXeyvrzdNV3pSFnQRtlEA8kF3bk9Mm9pE9rJPjE1Ns1Bk7YAwOGJsIFYNCg
hQdfQyJvZ/obmZl3zMoqap7jsuo8o616s4mLPwtAYcy+QllunSiehAewUKOnu1jl
YvBN19ErLcJXpwDJwu2oEcxcshaMI+LW4h6T8mjZgwuwry6EMXg08H/ocTzy1EQW
Rd19xAmRqTaloyUayN0Zr5v3Yyl5Y9LOWjDE7qWiRF6xiq7ncbyRpqSMz2YoGtNc
KPYn5gTzJe3SVPzsQCR6yAB+9jAe0Dzdf8aEaQKxGRttjaI6b1DuqEPJzNxfI7mX
o8IXqxFw21MqkhpIlSBH3W5pJpjCKd5kp300daYtCDr8zDLbrdWOR62QpA2yl0si
OXn7GxwmOXrn2XBqulo2MR8wQQJxV+QlWi3p4SkgVm1qthuhIL3bMeS6teAcqPUD
0+ji9wlSDobKrwrGcnTTJdp0YrP6yWl6LHznxap3ZLhUAMa/FmWdOM3eT/4+PTIC
QEbM1w1FV++0drwwAD3kk3mZeG3fQyh2ViZQN57+hjdpEzjr57GVXjSdlpm0Pk37
oquyp/5HiMd1dqsGk6ojT1NAs7CVQDCkb6QNBuAH4eboHycvZ76AzjJeS++u+q4W
V12lLrPG3gwyCHtTssqJ7Zf61M5FJHk5oIRi7MFnvvPthsrcBrdOIhivrGu5reCC
u4nRB7wZ+qlo+22g+KdWZAaZie5kIUpd5s3XXWWkdJmm8coYJAWDNsaJk/N7jG/Y
XhpofCyxBgsu8UzH014nW6Lb2I2I48HyrYMX0lJGt9+yVOfT83vtqYtdJeE8GfM/
O0si73LTLSeTtkhvV+CPrtUsBPeEqXXo0J75vEQMv/OuZ8cgaaVDAEUlt7Rfqz30
gRq++rLERZ1YktZq4/xn7JLfM06B/vYhQJTFnJLMByLMPt4m40tmGgkA+GESvPqS
IT5FNR088pfx5Q+mOYHNiVf9yvl9t//K5zCP3HI+4IU26pd1NbG2wBSbNxeTmQmX
hGXcF2NyLfok69f7mxhi0Mbjyzpk/00GjrQse0HFLb2yceLaQ6fTCsCgFkgiGy9S
Q5CqRlnZ6AqC7HzkMIKkul+ycIzpzzT+G6uU0sf4KjGXgJ/bwKB5TSe5rRDEeOzY
aqgt63LP2SUkzlFDa1VItLsUJqxtM1PJjqqotTggEh9NeV4posOikf58A6ZP5f+b
LuSLGuzaM7Og69yUVNfoEM1YVh5wd/wU9hbt+cNDTc2GqnV//EPVcAmN8e6ug7Wa
XsCJDKcCMgC19Djx97nqZnvewQOwM9FQV8Na1M5cEVSOIdLG+lEqEIsCefahUze2
Bw2h/0ZE8McgyoJZle9pRs3L76zvI/aTQ4Rksv3GlKbBR719kCqSNWhs4kui6R2m
srr9tMjA3epsAO4PrWFrO4G6AX8TesEAdCBCaM+XK4g0tIVFpIbM6pm40yz+FRI3
VJMFDgryqDpX03mh+EtNVuRwivRryhd0SjF2CBoRp9Fcqu5eBgJvUsZP9iyRn22n
mV6w/VqM7Ifbm5RlasmQKySO7bp0hJd6jotLTS4KKooPdMlzXt3emu6zeeXUsz3O
JKfONAQdMaNrbKN7/ROlhuCpgsFJZeYA8yxA/5K0QgxXa43feU1URFEq4/1G5i1s
reAxjiPiBfyNRu/c0tQgvfPiJKOaEUEdpsNmX+w5pLGPzgWJGaWREfShvCqfzYCN
msLmslHy1OYEzULO4hbkLv4wLCurhVIFnu6nb6+t0vAg4rKh+wmBo3OcdsZ/yL+2
wL7GmIvWLSy92FsHE3LHkhhF1ScKqWn2EtzXJybLj2okjeoe5ssf2fxeczLMmYVf
OHOBurt+BAf8sTnEG5bkwsj+KNmu3dQEC4xPnKeDUV9mimy5Q3NthjEfbaWjPOyw
IvYnSJA6aki+wLOI7qhz4AaSsGpG5tMl46oAF+S/S5Vt8rMfAQQhjOj8mqfbHHLf
w6c+U2cEAN4Ci57Wgr3FLIsemGUIz8XzzCIg7BQgvg4dcpwLJ3A2eSxdvjUtcD3j
XJmku1xphO8bL76s69lhJlKhfZHehMoSblMwHYc2gLwKqxmbJ+cTE00jUjOkl/rX
vdLCS+tzxIJ54etZYcBmgeR5vwFamRi8ECwCPFC1roECOuG/cqgt7Z6XPKigQ1e5
ptMw6KUXKCbJpGP3H4zvJP6WRUB+hR8Hpor95TQA7g2Eh6Nwsm9W/XVpqUv9X92S
Z4cAXy3LiSD3LM9SAbApSAUcygIvnqYwtVVVzAaxbG1Y1e1Sw1eP7fHe4FWJDVXj
Y0WPlX0QTN17h+J/mN1FidVhN/PjbkuHpXpfMDiqXVmzm8/0MbDYBqeF8Iejd9+d
v1y5AC71y3wyOxxi/pq6GxSkPx8nzbCkzq3Su8Lgy61QXXKR1urOGK34cy5iXUEE
+v7Z+LQxy9OB4QK3BByKEjvFarMkUx8SSY+vriDFPKuUQU4lBDCH1PMaw17c47q0
HvXZ3Q9z57MUk0oat3GjSzM6NNrOJ1dZpPovdWVrVBSnZBVQ8Oqt8DFsNtH4IZOZ
ka175ZjV5PYEiiWgCv+0wNy6SB1ujpZq0di3ndgeNvl/Hg8wjfwKJigoaZuPOpRm
7fZ8i0bUfyFGzJuk/bQNHAzfV3cl2ZkM4lNpokyEu490qhARl95QiyHdZA/xYRDY
dnC4TLJT1JNun295DSbNgiplPjR/Ig9qU+xLQ5Ulm2u6eJx6js39Xa8QZXN00pg0
mN2Q/qZCUijFC2przaItBtWCs6FU+CrbWTasa5kS+01F/FCb3CNJJyy3vAW6FMxm
Y3oz8UrZVQtdC/pmr7rAZyPol7Hv4cnEtDqzAtoOtpC9fzc5GCkZ99WtCPGAN0D1
207FmwgboSjlxbRDCL/SUXyr2xjUKZseJzFtF/0JBM4o1wZTxCOzj+fsht+X0L0E
LxR9P864GuU6PFoztDtDhYC/bxkM05GUmxmeAcoEr786UHv7csmcgf6xlR7H3iSx
pHmQT6k001V77bUzkFvMFUxU8eFwT640ff5AJp5f6SnpRjnWLZ6E//VL/xPktOf6
qLi9btZq06MH7GkyEtDTLYDzeu/NLSPsAJB0gt39/nnWWcby3zLkrqNmLtpYt6vo
9KeMEMGPx1ndu7O8l6q24ARf8vw2W2o2L4ylJF/CRepe7ZublTYf8yE9Eark7V1o
qkDhXIL8b5mVbGTtZKYvegSOHOpueSfc9bfgK4ILlvheL473pvWkgnRJRJWBuUoF
5OjGh7SK0QUdE4Z7c1RYVXe9yvrUL2cX8fhFjE+FKu3hQPD6c5TxMbJdv4zLvlBy
OXst0MO5t14B3kdoUtjWqbwNtVyGCi+SgGOBLjqORPOgDhxtxZFwoTU/pCdSiQ5q
iJEi0Qq1XW4nSEXUjruTcKcskEfbGc4ibkzUM3Jl/FxNfJcWoDZTHtYaYlqsRyYz
3SULTRC6TnqASj7kQaJfvR8yBG90l0MIrCpcZ+vPKowOc6yNrl4Z4JaOh7xQPtTG
5yzHh502Om8jTauktNh5BB9/G47T4uLCyBhMAUKofHaimMUk3UuAmolU5NUZuotC
gQbRGVhAGU53eVIZp1NAdBICdBKJ388GLKiJpQc98c1wcqXG9OV/ntvtJdyBxNl/
3zCJ4ZC12c+SUhlIlBBlPZqrFXa3E/qWRi0nWLk1DCJ+eJz2RbXEQ0PUf2zLim17
xOIc73IPEbKyOIWlyHVXcZIYEH3h6kah9/LusKS16Lc7k8RG1FSf/1ztvtXQP4Wm
pcLHwHOtpRo6sgIKN4cn37xw0Lwq6nGePF/yScz35R8gBE0MKGbc2gQ/an5PlP8A
ALiVUSnJ6rPTdBzJ3Ls82dEcT9zsdQZjnQcG9lEligTq3C1MyY6cfmimQRYeMzxN
qY0J9kvKOdTAca0SLiK4hZhYN169F50+TbnLTB2trKBtOoEqEcYFS77F77uCdGgl
hJ8PtUo19gc39ssgC6ukslCcZ740L8DUafUnwPu+4ijaYws2lMn8xTnQSxM9fViQ
xWx4UX0alhPJoy2PAwLdvP9L6QJD2CN4u6Sc5fBK6/9e2m2NjFpd+KeVxrVFEF93
o7zn3StDmeqqOr4YbqzgoYePk5ZA9dZa09mVIIclVyd343CZC4ehX0R2mVXh68OD
AVJ0lQj2X4oe6lczPh73gLXIXENAgkmxC2i53yDMXtizmS0tE4ob43VmxT6cf50c
0zxdPtqsNzBk0PCUBqkPXcB3NFuKu5r91uoiHD4AgLYzyh9lp8PxzqmBQFPcA8bM
DSjt4cdY4AYeYI75jTUIMmBJek2GaztZu5v6901o2K+Ch5JPM5FnUye+ejY93WCi
gkmzCY7KQz9GKtbSMv8E41G2iR6r/bhbcTnBDxL6bDLW4LbIejwZ+XbxuKdn+IL7
olX6Y99qQtrXMLVqQbRQ2AK4rTIOXs0CVZ737sOVFvcpMetF3YNiM5C6ZXVPMRvj
U5SS793dMGvjyO/BmQGg9+ldrxlXAPgL3xDIPzy0u6yRwn/UT86WhM8IB0ERKTW1
iKwhsFi+Bq9J4A4W+/ZZo8BHJiTGvoWAjAsSrja+cAW9Wphy18EjrS7MEe6fHFDG
0+XWpkI69SqurRR62rJbMemz0TGWIu05vv3aTwaDHkqAkrCfmqBVnMRlxEtWI9gU
rIWiS76ND0tGMNmZ8f55cHIH7LPLoXkM2P42y6H0w6N/OQa/3qoqy7vWbeZEsbbE
oQHsSq508wgQSGtJBBAuzotwYCiqdSmEwdEk4baaGmBd0KzBtE+CrxXaygqCIV0U
VjDhRmQb0tsDx6XGs/WZx/+PvZfkaG0jO8g6wulzm5qtWyTTu0u6T9B5flF4GzZZ
E/F9nBfsx33NPpIrt1hlmCTYydj5IeD47I24W5cNKqjy1NDw0cySwq1AcsoTMfm1
Olkq7ihIvAMBDCmPFHRy5DCLc/sS7nI+fMY5NKkki5qeql9m328dQnb/rxmFzxwy
XC5uxNexIgRwce6Ws31h5Xz1/AJSUALVptzqbzhDzTkWTFPc28DP82MNK5h4BWgJ
jHntGtzsIlqHTtfzs+tTeMmoEuIDsFa2trL/89SgIyfE5ZvgZUn999YwFdli2jKR
gNgJ3F2+UKPX2CUhht6tVOVvaeHgK+ZroUsDKr2isH1nAuDaa4plMXXqefIQauCN
AygHaiZCkGpM5i0UrQvhQKAzk/3EJ5ZZd8T+wXAmnWZZWk7tn8H0pIshX1Vm+d4y
j3StcNR0QLjY3G3jJoDbdrRX0VbuLEtuzhi3pemgK0sPHx2N2vvDZ4gh6/sWuO5x
5FS3eWVSpTflWe8n7hzLqHQBfXY67At3BKmQRqjV+84NQIGvdUmWmlM0KVL5fkk4
758sieg8X0bSD6WI3pm9H82WuRyebyEpoqu10JYn/Cfp7rQQv2QU+v+CWtvi8Rc5
swZ3kaGedhVKtWS2Xz/9rEYiYh0vtdM+R1ZoW8SFGUF5REWzm6Xqup6BBoNuTjzl
xWyRWxSdhX+f7r3oqqt5+JpCmdYY4BYWWej6N/yBUPaOn6bUQfhzkm522KbHkXWg
/+UArIC4tI5Gby3ttyYuggV7DWUJ/S9dZIC8I9L/z+q2Yf5Ony+obVDnVGRZNtSH
15qWqFjrKNx2N4qVev2lPaGcED9pKC+KlBB49URR/dJDHMAsneuncNYwjJOYpTGO
fP589eeBDXctCvZmkzmN8yMdpPBBUeJvKAZlkKRHNAxLxht81mxkFr3+meEAcD0D
ycWO5juUf1uxwY+UF9zpsyB06iojB+WXsGSLYQmHsdI4QDystlgx17C9CmZLHhgy
o2JGN6ckPQvFFnwhl9abcrsXbD9dGAbTQKXBoQZUdWZGpJ36Wx2bkQHE+EQqUi2a
WtijRrpqdBP20bmIbp3ytx/BlSTDWTkr2/xEcSP0lTo7EU2+I4RsqMOKTiTPRWPZ
yZ0mCqh2kTQJax/xeixX5aVkdKrl1r9z6zcD+CXTE9xUC22xL+oPbdeDkkfjIGNn
FkpDJRcI32e8nTSBFbHL6c6WkCOLflo2Fgi009za/D9bAfKY6zAVXFood60l+e3C
BfFDZJ8Iyo2dCXUcWExdAaVrTjoZRUrA2StDi7KqZhiYFbqFrXHVQ3nZeAMPTK6S
MpVai+4XhP5HoiWDIqIeaKBylzEmRIaCYkDa3IZqpvUajYoYHdycGWeiEx32WAQ8
7JWi+Ie7FfiCanH/fIjTYfv/kqeRBKN21hsebT10Tbb90pYGT17KGN5lzfZOjjAV
sW+l/eJaHIrZxbiXMfOROjgliaMxOWtOcJH4LQrzZ8I5nPG0ruAAbIWkteBiYhwG
QgAGAtTxycTlqnmzGS9aWWSVLG2Z1Im4mtzZEm+hXJmrdbae0hGzu/7eoeXDl1w7
kXI2o6zurAzqmGZj0iTP8T0hY9fckyB57JF9sfLazXyeyO+9FWJFN1PKDBrcq09G
D7Qg8dudyLYfYYF+DuBOnojT2RHXE3RUqDQVJ9n15/cx3xCE3NAUzuHtpHFUQU5g
LFQwQ37Sj7ppLYy2nhZI5NMP94Y7h2ekAK4/c7inPdCVSSAYKlQbU9Tq8M+DQyyH
9GOcQcvj3+YMehlciXON2UEZ4fL8zHEuh3JoNyzzEzQAT59taHokHrELwKQLduPU
kA2BeYygZ51ySLouH7GHsKVoTkQWqtn1Nr/WlTLod+3F6wB9+yp4B5gxoQcTfitG
YJPoWxWLrd6qfVmEbNNuyIC06o1pfvudnNb3FwzXL89q1YL5Rv2GWYmszdg4wk5G
4/ryV1vZ5tWyh+y1YWycFUrU/UqV16pMhNtl9Xem9OY09vrPWbT8ftj6pZG5rjW0
pQgptXJv7fEbiQBIFXs4MERu6sD/pjEK1dEL637NYYHGCHW3nWG3CRiO6Dco9m38
k896Tc8zzY/yyapeyTDK5HuJ2byhSNMYlDH8UAqJsMQA/9e1KP+3QmzIpgOJiYJF
VnhrLa0HoejOVQlXDq4v3/UwkmB3eQkrESrGpeButJxedV+Pf85qVM7anBFPiYnj
fHVZ9SsOHVzpHsM+W4dpmGsjVrb3K4A2WMo/BGzRp8UhvXTJkoN1MK3XVX+Gb1FB
4juYFZfZqwfKBkFTM/BLHVwrJfWR4WDVPO7JzHFGupmBljg0pktz0bmlsaAIukQb
F7fnZtPsXNwgcztHJj+aBxf8OrM4aiFORpStjGUM4FQUKYZgvM2WMY6FvbhePQGz
Toe7xwBHKAWm1IigYtPFeqlunptopaEGA0SHjhhtpsua1BW++eALxqMx1dqEaH1d
3HvLeayIEBRv188DWOas0rS1CdjOICQBWrRl7ixNIfS3UJomRks3nliJV5qpsQPy
M5XlmKIrpkYGvxOCuN+e39S+j8MF7etobdDUVCVqGziahAdRUwONeodXxumL+51s
fN8J+VXUuOQLJJX6FQRFkPLmdnIjk/yxxdTySSC56tnW/QSJ+IWG6lfa8ZSqDFBl
K5fr4LLymoWHJuDfBP0+vzqxOYku1Je+6tXrDSldeuWQvJ+xrMXkM41up1VkMgmO
m0f6JU4iqOtkeNe8wy0mLuBdLTv/oqOlwaLfJ0HXEbVPxFR4F1RoSdvQ0w2g7VU0
Mi5kE8lLbN6UogzsPsOG/963CaZgGv5cLWfpHtWeGWz1Buv/Seim4BUc43aywGhm
dpKuQleRLfTxAWLrcRQE5bJXalc3bu0gJljF5vfxz3MTloiHR3H1sIE5P+ay0qXM
owKxwGYadbkwA2hNzvsp3+2HgOfaDY2ffXhL1qKE7VjEv+CKPqfBzoMMHeZdoVxO
r4lBBZpRTNdNFSyftlrRS1vqLnh4NIRqjLY5AAHPCCfoLvbW1to9bmo+bglNvprh
5J6rSmKfnkPvNjVgNDkQKWu04GRQCqiMsa8loGG8bHO+2ufOJF2rN7lVdwGDDIxE
6iKUxp9BhiJynXEbw2jEAu32NXMyc4gyke5nM2kz1f50x1n57XNzr39r6TaFBx2v
DsoLykLUse4HGyIfkHH2d7epPYkdTTOOjciU+jYrSmC0bQK7G+r/6dGmY7Nkqu37
flRhMbL7RNEks/KHtKH5fFGvxuuQAlcOEs9EFfUrqeU/HNz9phqe6UNQ227te9Fe
ZDWpQLTTFWPKLYSZqfgNYM6ttZl+/Agi+qi457tCAWXoK7IT//eN8P60WNrjdtzR
XyNnia8biuqqtY82/elpvr9lMzF5CrpepX7rETbHLNJOxtGgVxlMJLVXC2PF16DU
VTrryNIam9kdVDecMfOw5B/bs1KPlLyxcAOVqy2MqnNVz9YbGmWZbXyxPSoMOZuQ
LvUiaIeJGPv1nMX/+91lDIy5tPGg6Mud6i6pt14ZFpmdGkWYK8/xdEHWoVpjJ/k3
dng/ePt3xX4vhten5178FPrnWZAp4e3YjJiNj3UlwbJHwN7EYDiFzpNSfP67Mc0N
RWSbGhIAb+IUXeN71EwLbLDcfLEHwZELDm8Wy46YF+djwjPzu99nFQ+i4M245QVv
nS+/c6unF7WjLOvniQLjPzEnGrhpk6gtvtj5G6ad6E7OBmcpKs3JNwvvkZ00RPg8
OwArMqFxfLTVQ5Q9dfNtuoeq9lrtJjtu4QVrO1oGVj1DdrSVK5xngbURZyulItB2
nsjr9CcXre3cFoG66REy1qdnf1CTCTaDdAIaqLgIkH+Qck8C/22yLi2tZ7zK+Z80
tz1wD+6Q4FW+uOuvIQBgZCgvLBD4TLM80e6I2jkjAJDFT/pL6GpZ/whVIHichy4O
Ev0s2mcRwhnryOYk2vmBuaBMtu2dudI/46HrlTsNcTAWLs0EgYhP1/xqaoabLHuu
A2QNR8v3ErcgYPyVg7WpDvmld+/17z8pOEM9YRd4JZx5NS8G6RBQfEIh+nLmqeGX
RppGNEHT/mLdnNiwnOHWkQIYYw53QyixE/eUxtQ3j8dhwIaKCzBoRVuoQ/Q5XRi9
8gGUERWqHUteAH0/Go0uL1UxBrX7y73KDr8XcIuQ8IrvT2WMNZYWJXfX1clHwFB+
wF2eW4+FHYVrx7C1wV3tZfsC+L364kO7GC28LZPduMLGZEcG4aTlw9I6YrmApKzI
NjXbeb/l0+fUapCRjtBxLlUiahIV4OWLxrbn312G+MGsTnk0U5yaEh9JmZkndkkg
6K4xFturDVnUQdgwhWXE7uuxm1rj51KqdYfg+H1jAUPvuS4Agg3ab3Kx8hNWSeo0
szRKSxjsNvXanz2Q7tKpEIkj7Qh41D5EQIL9rX+wbv/2eJPQgf+YrEUbS40c0aMm
3C6atJyzNSjJBqinSLVLcUsT2ejGRy3JiIQ5RBamOk9kpRqsSJwfzNWEVQkMI6YI
W0fgxDsuasb4d8HyHlAsP9sXUWQu8MjA+ovDf9lQ3p2anOTYVSVADv7gPn8Y9vpH
V498no/NMmw8VhY0NjKCPcfmBXZE70Ox+no2n5YbtNsjAxBJ2Bb0iAyybMYXuG4l
dcBYVX4krRQ7pvQfxrSL1jga3odccD8ai97T6Des3gYeSXlg/BgYzNMMiDormWwy
4o8Kun+IstlGxnzwRlfHsRO0xQ7nvZYw+AlWf3gnV6BATCStF55aRgsnKtIpOybr
eqDo+uZd8AilLZfxGVirmUz7T+t+91taryCvyN/PrWevivEFDgooEeBpA6Dfh+Sc
2p828N3Z1bTFeVKkO02NC8WTfABmJFwl2shx93NeifJgOYZGwFKKoW9dfHUX3BMs
DwE8U7VInJ9/ZzlSH4W2Mdi++ts1AXrzK7By8rTrRCmZGCt08cOLF+OfJHmy6IiM
yEF5khgMCV92o5r0gfkFa6lJNc6tJ9LtPodXKBU/w2Oq7mRnV4/tiBtxO37+iHYV
xWiMu/glBCRMOkoKwF9pVWDZ59pT6PTLRbIJtYxCBAMrCaxwZKp9Ju7ENpCl2McI
ffb+UvL1pLmqgU+S+xJ4KCjiJrS+B4ijD/E/Q/1He2nAT/vjZyEb6BMZnn3rE/oY
N78ZfafX/cfFmt5xvJQEigg/HKof9V5hwLqHrBGhZBskrNig10ADEu62TYIU3Hec
hsuDL9ZfTFxrvtFBbIr6Nk8jynOAHNIvWh8WY+Skr1Mjuaxqr2lLPUPMyLAi9yZh
0sBPbxONUlwojF0FdjDMuszN8lrtHoaTtUYFZ2yo1WUCaCFtTdb7rjJliX6OVEj8
J0Wx6JcgPdhRn5YxFjdR7EYXXCzU1LG/6qREvWW5xHhA2fAwTzHnfaU/CS9kzPsr
e9JdeYMXuYhC5FEUJYNq+dq3BgTeSD5wmEGyJy8zWkUBnvKLS54QmLvCdcr6533R
K/bi9AC1OSMRFjdlFjay9qJZ55CWxQD5dYwJ+878b+0NmrX5j2FzBEHZxipI4TCn
gGq4wudV+3w6jIlrehyciNRAF2MLG7hkeY7knRLxFkZRZfXWeIg0YTkjcVA2zX0Q
zyCWD2CMz+XRLQ7gqLGEjD+jtNDkJgkPRnovWBM019R1y7vXaxulov9gHAlMsp4c
yNxfBdh4/k1QZJYCs02AZk9g+RWkLxeqvhKENtF/0iUAyFFt1b94AQypoyKclpLf
N95a5eYf7pst16SFwFSWCfm2470fxE1ssmykVyPTVJzntxBloY7MR8EG9m62xcF5
k3/YZPnEPqJnOXTprFzKTQzkxwFPdt1vcA8DztjOQkzSN4pWmzQkpI1L56fbRYLe
3gHpgFQEgM3WbkOoo7/ZilZisgONZEDSYIjjlNrPeHXCx287hQOAnFXJdp4wl0wm
+nlw50XrD8GqowWMkUzmYG+IQijcgHwwv5vsYoe9vN/vSSPhQCEj4OVUEHCAajv8
cpxjdCs3swhR1pRi7T9UczPUDOjhu9Q+cG04Wl1H+x2f/8+/GVcjN8ObSzgK5kyf
FzfnQs3yIaIEyH64aaXCxVZPAX2hJYaZKA/Q9WYLRX9atMO23SsjAY+LU0UrZakL
NnDicpKCJBq/pdEL6XljoFMHiSb159rsjs4RI1uGk6NCviecOMmiEkurbnPm17Ww
M5IOYkybpq6D8nLAXjkkE7icdaVWYykGLIV5EqSx5QhoX/GyiKaKq7TcB94WSoUv
uduoGDvD1hX3z4saGZPjNZTUp+FMTSvJNMdDoV+LkeLeliLF08CQtSH/sS+eKq+B
UPvfguk2IE/meO1eiHboLDJpX7DGG9YLMtqvpkoDrOd6Uxykvb54XOxoDzIDC6Vy
5awfaWvWtaaHqf5jswJYKOujYDLsV472Zp3e9ZWAXdXcjbR3hZtyXiCImY88mH7J
bt3V4onXqSF/sBZVkGuedmU+X+iaRFK8MdADzm17EdLKxX7t9JqBrexipH/idtgl
MtmZF8jngPLUhaRVaKMP+fSDbNs/6wDg8fCITLvRRwOTLZEGhULV6xzeBE8/iB4D
xZn87E99bsR5ZyuLgxjARVG2VOMQ6OFkpDzmvRikFGHdvjpmBW4SID2uKX7zfdhz
JtCINZG71m3d0RUUQnHAaoH/tIopkoyQHAwochsJ7dbFUuK7na10FtbyLQ2DCsf5
oVbRootFQ3QCjMzcH7KB2+hINcAcmWhEfzgsqmKcvpFjOq/xnH1ID/ETLA7C4dbF
i2kqy0p3BfAj3dLeh0cwWrokcA8WNhR0g6sZFbOYXEHdvdNGgpNGOk7tamtWycxF
QLowakQ5KBbdUo406W25In3u7U5CxvAvxFoSaJhFKOHpP8d08ULRqL+MZuZag8mo
p3iIwx6Z6MQuR5fDbtQgkmMwm0Xsr3IvEuoWTNbyMOKHsxRJU7BsXHoREgAkxlmI
gHnJIf1Z1nKGExFR8NYuOl5xxjJiZ6k9x+ynS4bV9NI3+HyPTYPEaOZCcL2uIEjU
KcrQEexiqu8hKrLMojhHUL+yNCUB7EHDCmRTWNkiYt5uAraSBrar2PCoT/5LFRBD
nfEXlzTdeqYBjeoyjHW+6iolGZfMJBFpW9ieA6noSN0qOtBsHTTLNaiDiLfM/u9f
InSUl1uyxFuvSR0UKaayVhYA8kVU+Siew/vnob0ShuJajnfJHIUl357KbM8ZSXEo
ft7BC9Fbnsey81IPtn4ZRAmLdSA6VePZBsd4urtzSqmitnwo8VF4JgoSbtX6zB+y
mk1ia68FZHHyklMvXO51rpw7pJ76YUjUG5Slfu5xsb2zFuWJ0hnM+8fUhy5dNjkk
UDHmCFwSLGvxfx+390lMqQKwk5y2F3D5xM0sXL+jigDi8PHNIOEgPAoceaJ4BYMG
v1itzrSH8sAIF4vTnLJTAKx3FniNhM3PzPEI/COu4tqvySP6NbByqgiz3eBdY4Xr
FPEIEZTJU6VL7Fgro1NrTArmwNp7KrSFsewZ/B9kvzQaiYuuqVhy++hebJxtvFal
cv1rvIUol1WAdfYQ8LawWHyYQ31sXqAGW82NHQ1XhdXLAojizakW0MHgH/Dwm+7B
c6zDN3BgkNv76vZuH0heAjPUyd+JzYktPlbz84xUyWiJkGmQ3+/xIQUvDEvYQHEc
G/79QR3ygD8UI8gJYlJ06C4CpJxDMzSmgRxvW6T6Ih40soYWa6XnpAwAE3OLwVOo
EfwKTEjo0eWnjXmJKJ6CRmS+T34lKzi9yN7mtxAlBo2Ts3pKdwGaiyADRcCGDXwW
syr6folDDtmtESq3WQBDvIxHrQKam2QcHLJCD4QpcwZR04xYUyykrgkjcIBiHcrg
7F3SGLWi3rvrmwMVuDUuiZOB6DpgYgJEYyXK7nkK3LdAstIuShU2nvxnSoKoB7w9
S9XhjPCuWVd0M3AnUPMlBZ4XQxZvSfRUUBxVfXXAiueqsCxmGeBLlF3fdj8MRzo/
Ba6QvlEBa4BRNjdHZG3GpeIoQ4z4M3kg4YL4M0nWvhrjNlcANUevYJMiNKQrqOFT
+PuVnsrcHXbbBr2AIdn5krypFqz/50YIxU0e97M35Uvn3eJeUJ1OGAXII3m/Cze4
Gp6bvdx/cFovnc6aFOsox/XB4ygFBme0IxtfBqXuZWN3z1CDG/NxbdLSIgMEmK27
OkXON4jwt9qf23mxNt62rIaOzLGoebcJKY8YBTw2bhsGgoRkJrYxueh2mktO6JHi
wkxwsYG2gOziuHcwxIQqgR4vKcVJ7G9pbR0Yk5A76+ckG39jxxFAssNBL5aP/mDb
Tp6Bxkg6KjRUXf/z5GYuYNuCqBh4/V5pWM/4kLgF2JW4k83HqFfIPo9RjRLsUxBp
BcqJ6mBgTozmh6pZ21eHYf6YMvlCfPsWrQF+c5SGbjUPvsRQZFWdpK/k/hs6jzcE
PljRajwoX2DnANDIoQLnQ1Rp801sz/yXyaKSyJw8V0YabRI3eBsXmPO+9+lvyzsS
mSUXOAeeRSFFilOhpo0KWmkCimZ6+E9PVo37pX3GcnhwEcu8AP8V/KCvZsCQuLN7
KDERvIeFqOHuRe72FOd0Qmz419IcLeN7xcBiUEkRAjHe16nPxvgI3b+1B2IUazOr
SXeNxkpXKfQa0a5tCN2cLNIyFwC62sk03XrrSBWDBNG08ezOnEofeTJoQJDZLGzX
lJJmwa/ydC0veuWOfWab+bNbRbXNb6p4RKd6lo5kCtg3X2FMcTdXnYNOHl/YQpR1
ygLbbcFY1QK2Bft36f+aU5ovZdVb7FIWcXQfzZrSLQFZ/6u6x9tpk3UZeCF1ufRD
jTeW0rpiq6ksCHD7nhdm2MSq5neoOq79vex2CdzskVqNOn46xrsafm4lR6L8V6Ne
hudoFmSsG62rMN1qzE8ZSjiKgcN6BM6eCoMdqvddbGBtQOxlLH0bvm5DKF3AqHwa
aqDK9cDCMPB4YuT6PwNs1kFDa5bXhhnVT1QIkV12UZJ10fKfu+KMfcX5djqAwDU/
Ycf0uRrmGRmrdMdA+ha5KPT6C9kv5lzqsCW92BjV0Ce0Znk8yi52Z/dtLj564X0q
+G04wGypdXAdo+twRXiVDnBlIcWOr2Q4PVk/o5VB1+3yIYELBw/QflJuvLld03Ts
8Co/J1C7CvhYgm5pc/ZFopAJ/lVtoMr7driwh/+k6TLs5i6xUsyfAKmT6TekviGM
fRaerS6YfMN2rMcbUndDcOPZizV1oo2s+MEPw+lG/dfNjTCttQD4vqgHba7g3OQc
Hp+5wsIrmLygRttSTVcu1UuIK0DZidqtum+zRHwR4MRA6+dyo4Jar48QxP4iOLqM
3FA6qaiRfrc9MOEhAweg6jjWtmmynlfCGHttgqwqdO/VhUjPjvm1Qz5OUetWzpjn
dWXBNoCi5YgAZwwAsh6qKrCPhMK2dt+kb/w+1B6jEHL8m4yJmtS9Hm4weW7E5Dj9
Q1UYJ0ncX5hJYz/YABDxNI5qQ2mtWZXNjNAqAbO1Sv4grB/6vbVGLJJs6vQxayj2
RxKi0fIZrh6LJN8+B/ougLbCtBFZ/ISL7ds/i9v/7ZKSkv0LWLMaPwHNLxMQ/fIH
vYSsDBSBMv82OtUXSqGXUSz5zvPyqp71sZDP4WUHlMYpb4mOyvtrdsCztSEQ7uud
YyJHOcsgzVjnGTE5y9ly3i9bxlRYYoQ4HIkgE846AW0Ntz5tKWHoWmZ5UaO1xyrc
F4P/3aHqpmv51Y2P8bzgvDyU/LTzpBlkGGi4qJTpW8XAIcflEILkoedlYMSGRf4b
oIMYJBMb5O3Mqlec6K82TQWSq9gHXihvmNDAcQg8Wy1Zc3nzKwWAL5lMGiY1OxB9
b14Ve6hC2zrz9+oHlRojAwR5Z0ZFONjbFrLCCQIKh2qjXlJ3IFFMjvpWWF6zzEuN
PPFBeskefSAuogpLXAj2jz02jbLeEWoJ88eBG5Y/02Asxy9zVgX+P5HN1SGQ46Lm
nZaS7wkccAOFSANRDCSNatlTIMRmYbxN08dV2biHLEvOMacNrUwvJDrzYn7a9WjW
dhYU3Mh/awc8Owek4krdZgTNtL2eOfXXpxbr20cxJSr1kZ0WmqehdqcUlgZUCiC7
c8huq4brGb35raKIoDPD//5jFd9U2IKeno+28xZeRU0WQvc1p9FB8143x3Vt1OgU
Titd4D/gVLmsSNCeVeUldDN1GOQU7JVnLiznDafBG/Cpmc1PkQjvU2xG4kSTNlFP
pjxN+fzOXff/Pzk9gOw+eVXdG9rMChHP7VuJHKR8l3mFkp9P2ONiz6nH33mGS/+/
beug37b/SF92sPudlXgvrQbtSGgpK7O17AkM3tFS4sJd2n8D72cft6EAnV1Z7xUT
s8fF15Hv0BTxloEKzeLrqGhn8dOCwc5V2u2FgXrcbD3D4VEkdazZIPEzr9WHkFXn
SLjmEtvHAsBDJNeSn5ysI8zDT3pLdlxomwdcUp6qSRSlWP4jAKxv+QAZplKeMyrr
7JcNwhSX8v7Eq5hsXopEa38Hg6oYt+qb5PeeETwASBM6XA1B2g0WKJRDTf1xwzk+
yRGySfxbP9t759QSuA3wDhiCkbyn6sGhf79vacoSzfofyXp5CLAz94CMVS1AjWNo
iCBrbiXgoII67AfaMGTU8BqbeGJ2KnCq7EC28lzhNLz+9ACDhDf+qwYMO/sp5c7Z
//R/9SHGIf8blTyZI1HfVGQQo4YxuGLVfPjNp0J1xQxAvrO9gM7QUe3O1reJF+Cd
d4IvtSMiFNiEacRd18lD5bHMFLRercWL3cKrxKP4qxxPtsjLGhCMcIo5tgo3qdt7
HkQEfPfI1Vfawx3DV6KrpCij7AMJluVKfPgFBw+V/RtSG45fQr8FZwGHPptJtyLB
818BAhmW36mvkBtohpUEjruV9/1eM4J3WGhyp+rwHjOuG3+jwoPUwmMRx7oKZ/sJ
ChBzjT8wTKLDsoo5q0pzAjGbvTiIhPnZ9rQMRHpbg52EPUdMXoWx/bkjjMyVZieV
64Yl8S11p37Xf5nkbBHY3WfxrUnNPLOkAA9EbJcA2YkyzYDZzU+xEldEviBYc8TJ
nWfxSJDd6F9KPKA/jJjXZ+1Y4syMKPpHl55UZQt2T31JN+eS9POJR4Q/OF/JgDTk
Fk8kwF2EsEyJ2GdB2Pn1O48u3O+XV+6SyOUIUsDfVueqryBHMCM8CzzfaIIWXitZ
ZzHVueqb3BGOFOrqqwzsrr9Z7i+Q4aoVmOE4XFqqJBp7szXdFCRbKmvTrw0manll
GBwylpC23iIkJkCeBpNcXrR84UDLGnCtNc3HXTzIFyDVJJri268EtLYoC71p+jRH
oZmDZgr6NbuTo3zKwxkiBWcynixmJIMC/gPirVhvAwvH+5CcN0DRkKxuL5AcpgGH
DSNjbfnxHT08kGpSt1+2sdY11Xmril6pEPYD1y7qUhJ1mK2cFvOxdwgefoWpBTu8
QWTICP7rUKzGjdLngGqsSgJsNaTa2MxzvBI4FpT0cOzCvhQzEqDDMGF9RNaZfctn
mqcpZoSEsKiZ2Znl5sbuaf1Y6n37LU8SdvXvkjvbpEQ70+4jmhgaqNxD5BDdAsdp
Ve75gXnNFQztScr9QZ6oporMjFbV3xFvqa83QToD3SW/md5B5rCuvqX9lzhTLT5I
eaFYQgWpjyNXKdVVZICw8lHkEek6cMULVnuCKVglXWk9q5fnlTfouXIxOKq6u/LP
yr3U4N00qcvGvq7pTuvdHtNv8suTlhKWZjf9IQBKI/vhMXSkHqAgGrRZS9V386XQ
gfVGSWAcVp2x30rgMVHvf4HkO6iY89HsvNPZK1s0nNXZX0z9wUWlBlM6P5lGfnpI
8OrC0mdh4XeMbD0bSNc3yYC51zB4eqvN5uc/JhvKsco/w49afzUHB3Kk/5fDfk05
LBQ6masqjqzrilZeRa8cRLDwMome2jxPPI3rLghgthDhIHNoIoXEq2Bt62KMWrfL
p+gAQpNeTYq9BZE7lNbN1te17UQx0jtoHtZkTG8ouiKYH8p3y8AazIFptQbFme3r
R0EgN6xIEwBd33V0sJ94IKen1dAioB8T8dlfkfPvJ5rdr2zwLw0NZGeanXE1cGvX
eafSE4yjrrQJmr9UIlMP+ZU29A7sOzKZmaXB4txnNsRq/+Af142AhRyrcntmlyU+
ZG0e7ppZprQb9Az1nJV6VZrF/YpIxi56XTRynrPimKtDQoKymSirail7OAOFT365
CMt34L3SDvP6JzdsEQknLqFNc0E3kM2v6vJaOpOZUlXJJGlWbgkJ0GvbkU6okGaw
bThuA/siB9wUVA45Jbowyg8v617JYo/HKVLYBjWABKBPFnUPrUkNmucUxzvdZMjL
youJRjcU9t3usSgIDU4e1Iu7gt94SJqXuEj56EijKAufI+IeS+xaySN8uFWy4Zi3
48Z6p2Vo3UPAnUrwZMSrog61ck0dbgKvT1e3/BoiJXpoBUxRm+z/nxldGUO1OrOr
RTsule+00bJUSj2u/sRXgJkk2OK0GBGncPY/nGHc8ukooisuqY71+66Phy6Wep/w
Ac+/rMJDNX27V3PkwQGAG0dwiXo0A6ElpqT6PX5PhGEtshOSTW7LVCaI7cBTwxfM
d9rCseXhe8Pi1aUJfRuUm+a2rEXaklQDmCNBQmC2CA1KRGrFwN0uBQliWlOsQf6/
LA6ABJSouwDrDToriUj1aaUKBl1NtlnmOTk8PQWflVBpxLkgRqIeypSRxyjvyRyJ
GgWDYhudyHRNrwX0rfgIVwSIQrsLIIryg8QoLR3Ar/4bTY0W6NudHTRYjQv1hJfA
t2Q5Z/l0pRhWxlX8j5dkiEw7CGQAAde0FrJo2Q/RABFZV8M+fDteeEPIYvL7dDRJ
XM/x+n7JiJ1qfSrM93AUzZekIeUFXwMSSEhxE1rYRQvWG2iWOKSfThe9v4iMfcQw
tIVo4d8/REsrBsZLcszJhJMiW7NhItlclT1ShtoOZkaMUGtOONnjYVH0oB1PSCpG
Kj+CehHhr2V8oW/Vw7uq8LkCjQzyEnDUF1phOJfclhVYaa/TZ1gK9TsGdxxW0dDj
J1ISlwomZAmcZ905tvka4uc3WpMc9N6x661KCHgoftb8yjlodpSqFpv0NOoCKuVf
1BJ0XTH2LZUgqyYTX1TZu2u36vPBlTP9cfsQPUJXDtiYPrNBsoq7OwC7oCLwzcxk
UK9hX1HJKOIJeQFCJiqAZBPcEX7sPs0drnqmpacX6bZ3opzRyf6YgW//cwVtOUT8
FskH33VkAL+HiHdRfyRP+r4VC6uSXL0bQJSH4l/FHXi0NLg/pZ1T3MOeuYuXyqua
PC3xmMl435HukZ+wrGyvarozrocpxV5SmmCKlti0mae7g9jAKJbMbxOI/XVK8CRc
FoY7lZrNwpKB0Xy6Ke6o2sW2ZvU1jE+eM3UmfWmxJbzu5+Q+Ea8Ht7Vjm3NDiAyn
eG8SqxfMemOfvI9PeA5r6bK0SFD7nK8LGcNJs3ZdiTa1R8JRzV7pdpG5ndxT3auO
WeRIG6DDbOv8cN881DrJtBBmaKY5Qw5+3sAAVMC8yXmbrLtr/azm6EaFXArZ1a1r
fCicbaFF17U2Y6DpiTdP3GQISVpDbgBF2JC+ngXk3tAn3bFu7Xkjm0J1hruXn/97
DM5zg+S6QYfwI0u/4TLkqJWcjaM3rDGsrf/6xMpX3deQxBSG3SiR+Y6ftaWG8fvZ
eBj6T6ZyqB5qSxSAOxExBU9iwJj7bpb/6mxsy5gX7dixsrFxRx2ZbIhXyvQFJPdh
9HOsP8YZ0ed/QuTGTnwqJjyDQ7Nq5FLMcpv7nRJMGhPbV78uaEzy4Z3Ahr618UGl
8ZNs0udvnltLRKpAARiIpHwPoyKDvDeFF4XjCBswfE4e/UxneCR5KBvD6EdcJ3Xp
AaxO/PwehSCY5KWrwKiMVDb1HHnvT60T7ZC4IwQx+D1PuAvDFYKO8fsfvj15LayH
WYGuWyf5BhDeEFulLnTACxKaofJu3q8soN9Il7Ebkdg+w0eFK89DYfQkCFAJT+u4
5lBZDdEYL5z7XQdMuSW/lMOi1PaHXi4M3qy0infwlXAd90HwJW3Sg9tVnUL4+nUS
18CUXFHci1jSVWaY2IP43cnZXhi93Km/2eEo7afdaAQv5DrGgrkQUHfC39gSzD5m
ZeFr9xiqTQMkJo35BZRFr4CsJ2pw8DfJ7P5t8Sb3fQanzZrlMB+kOtnlC1Kqw7jT
fQf+CJYhN9frsK1jGhJQun+08R9UZLM/dY9ydw02yBwAMrY5Fl6h6dqgewdQQ2ST
isGOQHB9sTYpZjVZzgvHAD0wWIkGiE6hhJ4Wz+5e964A3V/BBlkZhTvzlpYbFMB5
/tUuXnuyF92RzbA8Y6zJ9jVCNVpUDk5q6ach8lNPa/rXo+gL4wzyZJTqbi47pXtA
TkehVV5CzEk3V6InA8C1rzi2HNEu/qYCKYi3lihoDHRkpp6OGfHVuxT+Hu1FHP/Q
oE/u9TZy9KIXfSVMS167azW/EeIXu2ut7ms7LwupsKvSc0mHGoW8NEWpPW5mWSe0
7Z9rxa06KNbugNNPGU9Qh2BGPIJ4GZxIGKFFCUbc6g9TtN5sKVMDbu/g7/cXyzfj
/XDTE46+DWz4hBcXn6oe8LMbtJ2Oz351MhKiVnU0LU611ARZWQ3BHvTJPn0eqYNZ
ah+tOh37ttJmknH+TOHIW4dazaOeb9PX59QxlE9cOKBZjOwjnRfCa0O9s/lKhgqy
GljlJ5sqcM76L3bT0kzQpom1INNVpv5SRbt9yUXvWtjylJk9Nn0uggkGjV3166Ac
4LXy/tLN/1aif2yjstAYsWSSCtfo41d0bwIakuHmumQv30+Gk9o4JvDD/Ea+lpqb
2BSf8d58/Q7sEVpgCTrn8aHf9dpxU0WLWf7t3izD9m1pXOvILTiTNnDNCUhhGAUk
gxP/GxMtWES6I++70UTmrYqyM1C6FxizdS/YJjv9yMh6I8rh538eea3+2niT/mR4
AfvsQvMYEgTgiR3qzt2LDZ5pdxZ12Tb7HWr0eI4/dkerewBCXbTa7spOGLdkc0wC
1EfHiMNoVlvV6oUZS/GSnhw85WP2a8XTozRVS6mCjG/aH6fy/IHjFAM4tvDEz0C7
0J0zmJ8MgK4hzsSBcjxlWNrllYsINuuvIsqPQQt/nPH1iyG8M6DESOdwuZxOu1SJ
KWUr/sjN6mlNeL23FJ6RC8GKWEsFY5rjkNqJOuM3ScOq8g3Dfuvrdw5FRgRb7KHO
DxIXPwuXcX0ZRamTZc9vmKy8JxOUT3U/nFJfF77okq7odiPpBUd0YwZK4QJi5hvi
46H1T/oMSj6rJsm6R49YH/cAWc9NmGwdr7qjxmPrTGGGdKDsfRjnffMX4Ilz/bNy
bzkWcCmQ2XmplR6d/om9VqYZ15hyetFct0iQlO0oMGCtl0dBZBFOGaeRFbhe+bsK
bOWKFhiUA1GsBxB2jnyV+AL8rh79uEaLONac+LURftczuI5mnczB78dRppnxUXWH
4Bs0CcAESTcwVn2DV4/hBdOjrzT2NY2WITJoLBk3MJIjCMTfTqL3ORHooC4nlgI5
7+y1gJzw7lH5p/vE2S1DvF1/vT5RbS04JjuImw3a5C/je2g8oNtJse7K7bbKs9Le
1kan5suMFK8pYlHUtO7usrDaoIC34oMqdwaLWrKjF8Q/O1Q5PorfdEvzmLj/snkY
4+rSnXRSTldO1KiDCRnb0iUHiQ9tv5SAaztu9gPXO8o5GDC2rsS7WUYJ4e7+ScIS
KAqiwUedTI5IArjZwfF+TnzaQG5RbPuOYvmJx0Q3kNwK0EQFMsLgZV8nSUyjisC7
ts9/bIONhdCv8BvbeN34BdjuL8oSXeKfHAOTuqOazwBB/jLgBQ4uR5nxh0Gc8vne
RR/UC6H96bNnLPCNaURceFFkscgJ8jQyxoYwqAjJ2JX7VwoiptmrPyEBImDdI5og
I3BdF544/L4ZGu3CtKwfSaGIH1h2+ZDZBuRTAxn3fyMkpgP/O+mKYzd7M/t7bcaW
CMdEblIUcW02Y6x0O1HFFzHGMGF8Ls3LITmfPNu3LjwQnlJhhDC/1BbupvEIAqdO
U8yWt0/2tcvkOjpUnbsX01CDdK9lW0QA6gEHeid3cNYdsBMwxihaBxOzfQpU1kkx
jBJBjlwHE6CLtntqT4HWtOpzvBw/EB610f11ccqHeldj+VpEbrum38Py39EraSRZ
4d+uAbzaBH/Gvw7qxShJ377b22l58AoIhHPdHkh0wkK8QL+/f8nOLL9rAc5ckgJa
lr89W5xzA27Yk9/yFWtESKzRG9pphcBw/mhJmvnyIWRrJDCNkRbIYkf8YVcDn90M
YCF0FQ6yOBT5ddyptNDD3pVrXLCgxAUmsE2DxjNIqUm2FZv6E6JMq9WcJ2+zAyuQ
5R832Y1gP86cD38r0P4WQTnef4pPXE0v+8psAjZlWEP0RxRRBuFSDxb9t1MzDnS3
yEp4tTcZP0qGJ6tHaDyGS1uZfi27wOEu/eW8nWyM6X/5zOtWBrG9uk5DmDsRzEJ0
wCl86S+djYfYHii8c3Cc2AZPGcA46GTB8VG0oH5Ql6mo6xz+3FrK9suuNIgtEXOn
3c3U8f2eo6Qy0tE9yY0B7UVl0Pcy+YcEEk9GwOf+6shRu16vy207GhUbyfvHy5cg
IYZwhaFmCWVoCagdeCYykISY2OyzLzHpB2snX/7Tj69yqSUZhDq4RrEXqLwU+ol6
MNupsg0BS5x/0eqim62nL6SGGynFUx9R12hzqHedqo5wQGafwr/v+bSJ1FTZdAyG
r0JwPhqcOnp4UAADd140y5Kj+DvMVLpV4QnvyBhTcftBLhnHmaTQ6cPJcMMhnwXJ
JxfNvQPYY9bkbRoszyCT8PXEfQ09dfdJiWWVpRFxTeYwG2rfrKQRsCAJmxNAomEG
cuvlDSrVHyrUBaE7M+y6sRO3gbltMxXB7XV6cc9c0JAuoG8JYtP1abkzpZnZoiah
H5cgcvNqqMvVpw5s8TDLgWB7BFVfLAXlBFioHLrg63gluf4+zJGbVUhPMV5XTqXI
rq78xJFkwhRndl6kI2Q++7zsOq3EDZujThTqYsbAPTyEESrpgARNRQzrD7vBaKQH
osmR36VYyA2VsnTXyv+LNki7uKCBV1stLcW/dZPcq07WRqFA9pw4MFo9+gCLfkuL
xxJyA1biSzvA0suWK1f/ojWDeetqq0UgWqOLFQyz1oP7dRLrbcLsUybJVIxWNNud
+9BIFzG2If1NyBY38WL/eOn4jmSi3yX2B4gSn/ZH7Uxe4XFjd7tBSaEFBbK+JGMz
s/wpBJgDAvdtEr/T5+jZmvBxLoIyo6RUS6NCUIMjCheLuXj0Kffb7pJ9++54Fg9/
/tz2uo3zUQgfHdLme0l5IZRgpOc40pkgMEm1KerHFv5YE9z3uDU/rBYyaQA+H9P0
pJav8x4PUxG7QjFKrVLTiVhSmpd+CND+7RwK9ByUE+LE2oeLfAgpG6i8hMXL7Kt2
A7Bz3OGaRWm+Zl9XFYlCaDfuCjuyiQJBpK+2g/ETFaWXkDkkmTBW95uhPIc6FCtq
nx2kwix/05x089ZJHhnXdSso0Cq4bel8RXTR1vIT3MdwsLeU09ksAQkwvfVfmGrl
6u0UaVZg23DC1YD8qdXdCfWlMybWnNMF/0jMAyL2pFad6YOCflkd57bJDNUbDq63
peg22TuR5Gy2r394snaNhEqV7GFvC/9CAF8TTVoiBroN6IuuIH0n3uGtmvDMCFSR
bPFXvhbymXUCLD4Kv3jmkUCDaEfL4Nv4G9qj5MEujMTkqFfXl4us+DV1HDHWxKkS
YUHLD/GKcyYxSYQH0EAVx5w5aJ0GCjngMRncPv32gDIj3EkDRkk+quFJittPbotv
jZrYBiCA1DhkpQKGAaDgr/lO5v43qDr6NH7nD9ynyyhUVbMPvmCpD4GwxoZ3e5bp
HVdnmPlI3ECZ8avOBSRnfTLs/+TbdM8Jw01D3MEDH5MVK0tQEZ99Idli9YdeOuIF
k/QdJjcdIsALXpMfpZKUMN5metmh7rAf7pYmqcCiE10HRiG2xHvCFVT4yh8oLHIU
acnOg5115/WiCT8OPfwFVy+u6RNXO0f2SZfNZAo4KOkC1RbW/MzksJl6+5DeX4b3
jkr6vjV4qEKeYbJK3EuS6Ksgq8afaS4ZoxVVFrl8bQ/3duPKc886DdCx//zVISxy
ZdhnTsCSKivDDIqn/p8+scq3gfmqsNXpXM5tsMRDQFo4DgzBUu6MPoWxmdoLi8z3
JwxbeNDzDGsN8c9JbMvvaUw9YbKmliMjhL1BspfLR0sfHlxPMb77/WShRh3uIPnX
FmVcpn33hg5TD2T8mWoGg4rcvUeATfqdOw40/OM1vHxhfgzVgQmVr5Sc6F6YdT1i
58uOqpbWkfptgqn6LoyRkOil0uRGFAXV5wFdisce6esSCazgT2KexjEK7bHY7UII
mkdymxvm2mATAPSV70dbx/FwYMERdLOGXzUghup93BuSc+QX/cA4an5liZ5stVLu
apwGebzwao3b/VniwJwOko9+RKsyOJQ1HwVM91ZzVzM3UWd6ueIYDVTt8d8xpx76
+szFIBahcFNb2DCQa5JP+V68bLi0dlgt/OhbRzzmZMW9FGiWDDi3h7qfa2Dh12Qx
5ekS50gyNwvFENwlJ+2nuj5sKhIderv24UJWkvlvf1EgwgQlG750Slm4odQDLWnX
6KrPQbF5Qncy1s7Fys9HXgZ2MZUxADooQ27I25YynIFFn5UDPVcc44xpPyvcbDs1
kwYUToY3j2FaDlyygD7S776foUS8YyVNzyg5GmNYZckRTetRQc6E4RN5DtAt84+u
gykF5KGzK5EL9Fn6kqwXWF2v9uS+zEec3xEFvakzrh5byfMfBF6BTZl7gPKUKGEO
uTsvnunaPkaZ2daaevAUitv/+pROaMln5SvitbeGatlolwoWksugw3N+2C8cF+/O
255JI6qkyO3KX5E6MPe7XdFM133dm45rujeJsmi4S3ZYVZAf7kVdfCao0EVTvksJ
t4jAfz9zW1MQapeW+sFay3oLGhd1DzMdLMT894tkCDWDFNHLMxa4KGSs+ud9O9Pr
McWaB2teo8VXpsMZdb5NKsyoTeQZBG7d//dFh5NCX2jmb+lht3sRlAiiTXYOaWs0
a5iD4LLyX7B75qcnGsD+65m9IyTmQADYfHkhI1myuMTBDBkvJa/etfspk8BpT5V9
rnjXo5KkW/eQiyzQmMMcnYpZXZif3HWq5p+O4zy5ggPOCYSF+vDr1gO1yVw3/m1c
7aEkbroeOMGc/WCLGLB/gPxhqTIMhPOKyLQ03UOsuidoDmL8BBTBzjglbD8Kqrsv
Ge7Ciu6PJ4K5cKKt+hTJRqI4s3Sv/4AuL9hiNi43D01pMFFroX3iU1LQyAH+798t
d8fmotGHqle9xDQTYDFa323F6fzXfqEs5Y6MQuPoxZGovP8Rjz2fevKJm/m1+dAE
+GH1v2CSHzJgdownsTeWahaSAYev4uOi6EdzV7pP5mhhFV8/+79WtK3qaTk02DDh
Ow1u76zyOprgX/GB3rY/XOhtR5oiMV8B1pbu2tHcZ6/lGqXSKV5vKPdwBzBYRKoU
gOeW7xf3Wbi9uuytZcIXOT7Ct+/AxM4dUBOLwhFZYYofp5YH2AOpNvH4wMRsjWBf
itiTx2vkC9xDPiJsUw9f278vo5tde4pA/0TSiC3uiEiLR8Bg3cKBBcjhLaPEIORk
joDLCpE+lpKHluVvSNkBECHBmymq4vsu4vZ798uQGhKvIofKOCslcXWGwSlL0vcc
buzop692bXz7ElQ19CtiM8S0+oWgDcoHb9b+qXc5fkBw/sIuMPTLIBYdev2hjpjf
00pqQpnvQhz/JrrbugRRbMSZ3hpNqBRVocgh2H4+Uy9SLMFpG3C79kbYdnXPqR8B
3GKj9hDOzMfxmzoN5rVEN8ssC+/LdjfcjGb643R3bReWFXMad9/CSA3vsKy0iB0c
ToDi/n5S8fhlwdSdrm5ytUf8hiN9RIi1VvFCa1ivik2xGOUIghg5nIpaPJLR5NK8
k+mW3FtCobuQJ/SMwvuZ3R1TBR80bIvNy6kEWPu9udOoSsHEQA7SS9unSrDRPyrX
DPdMnYyfCdmqS1g01y2u1B6uCfyorbUVq5a1p4J9SIhrqmKDP99ZyhEENjjQIBG8
v2L35dLoC/B62c/CI3bK22F8dPZeH/DsZz3N2zF9YLC/jMxIJ3k6YBneEY4zbb70
ojhtsyfFedZhxrG1fkU+mk/9g2wKhhg+ObFcttbMHr3jCKyGDcBFAmqg0mAPfBcR
N5q/KCgs3F9SKK79kA2RcYSbIGF9kGVlSbRYdsSgSYVEGpOkKaNGpliayZmc0CYP
oYAxBSnkApU2eN4Q0IPY1YpCSrmD9TXtZX5SQvr9+Xdzh1tQkwaIvcEw0OxvFyB4
kgr+Pyh83L7/GjlxG6LjxXN99dgD3kcedFdfmyJsJKglqzDYpJcB2eR9JyKrYDqE
B35o8pfzA8Alwd0zLvNRkONpc483bLjFV4L5WrLQ6CtmVsGz7Vxvs84XpuPvIRNM
F1Hda4udgCV4v1qceyYGKxtUFP0HP0rtFg0Pzh8QKxE8Z/fpXZDvbhI3WhLSXJMC
mlm+FLFk2k0yreVgH16kHC6i6hT8G5zcYDsc3G4q8fPB2PsfYWFG6pEw9Mptk4Yz
fTKUo99d/kN8pLYegJQ5k+PjoEWQwHax2E04mD3o6tnhHALDcRpvhzqhlboFBmxx
2mqtxlVzYnU2yYsBG4a0cgWQrxGrqcWQvd2vLeJCY+Wet9PFf4jUupUrgUD15X5f
77dC1j9+Axt7K6TXZLn2D4LBpWrZk9w5NDidlfduD3d3YiVthvJ5q688gyVSkFyB
Jx2lVW3uaFbwlJP6uHiuyc3ZK3mbXvu6hKU1SzKXYW9m7CZDco6t+lekPwhK6MA+
f2X05RnIbF77uQ92PnvYGTyna24ETTfeOLsqwGqhTQYaIvfp/ohyDJIH3k6HSaaH
aXlDHin35kAhBSYN4CTOeVaqVZTM1QERvq/eat75CCWiMjs6szVPv+ypcDhHAMME
5wVHVVDkB0t99mom7UynJu2TqxzQoi49zx5oraV43azKVBUh9zp/kAT2Vbv5yTig
a977e+DazPeIg1zfcbr7v6Wf7/cfD+w/HxdrVokDMr+N7iUkOB9fkbfRJJefImLg
Rxu0cwrjH6k1/S+scjM/c1eTADX4DgQ31em3J6ABqpvfXCqcDizrPY2DnAvQcprb
tVjARWPorGrfEclZfmz/eNKx6UDDwcJdJpAfaZ0qe5FWNIw6l2kYsjZhneu7xZ5n
1P5a/GSB39Gvdjf98pFRssAVxBrsvED3PDvVJG5zjcrHYpIlQZH2N6FGcJiFi/PJ
5yzykXfNPZZ3eC313ouyOrXWgrWC+WRcBGG4soCywEKSAvV58UO2xOZCFexN2RFl
+OXKhDvdaF2Z1YXGguMXIhc58rOSHNj8I4nlvErnuyrQiXUF2nXNV/uD7Ww4U3jz
5XadBk4RJOCQMLECD8o0m3aDTY8nL7c9d+x7L9Z2PmwVhiBlMaYHQkgULBcqy4EB
PKht9oyuBNTJDAOlb2Y7CTpiCD6ussP0VlYSIC3q/DE9hefFeUIxuK8zojRMf6Ei
Qocwzx6DHHjUGoHo64CWt73wk/iv3C5KtHOGVqP1DbJ/TRVaqWOdZV3nxvfmbtYe
jzFiqMPJzDbWY9pC1tHr4kMh4njs9P7rspQXV1sLXPsV71N/b8mivmG+FsTg7sMZ
X4BT7AmTOM8DReJChzVlzShnf2awDDWa7WMuFOLmVUrw0SwkQb/7i3pWMcD0sQys
jws7xofQEcmgoN5QOhGgc10oJkmwRMlsdKOxlEPUqm6oaSThABi3zuYCBZVzKK4q
SU+e1QHgMZkXHed7jm5eGX8deecAQA5zFU9FjQAWzr8jrji8uw6KCYtAfJN2qMAt
j+k3XERl6wOEuWYr/E2pQe2vfC/G7vaGwM64nK+1vZxK/SMqvXFPalVlRiO62Hb4
gbnmYtIcuP2cxsBmbiu00jOu9k1A2tjhb7a+B8DINfpJlPVOFl999AirJRALkx+5
BhmCcxB2yA3gK8B975siV1kMIc6f0UNH6SubvOHBFbng9ik2SrnBJDu6+k1Sbh8l
bAVN81GQgi/ConEy7JkPImlMBJG+sFwtZ4SIpZ/rl7ZL5uRnpmkxrANOTCVAdnV3
fvWsU62xKwwdDVdngsu5IL37umiS3luejc8XE5cXyNoqJJqK7LIasCulWl5D9Bqe
f34r89Ybz4+fnxq34J5MU0CotaIrmPA+WprT3gnp91SR+0Sqc0rJXTdx8Bznnbz3
fyGNIqEhCIUdDYjN0/Ms3BXaj2d+iDaMBKhiJCqq1BxLGjJ8LnGGdFvdc8d0iAwc
CO5QEPpnHsTfa3Ho0DxWXa6XmC8AJHE842gst5UD7yP5JVlnj+1tNRrxggzffpcd
/eaN/8qPq7nDHlLegnR7uGyIZao2SI+RuLw4cpp6hz2/0zreyMVpa58Rfe3sxJMi
7xdXxAVaT8MENJFGcBNNKzaVLHeT0za2c5xM0lFWiRjgNMSe9Nbw86bToMaQRjOl
hxdy4r4tONbpifcCI0RijXml4gOeJWyE1vr8MubD0fDN2KcqLabF8ghU+1+6Q5lb
tT8uocUQ/UGJBOupM5M7aFVZX0QvmgpgdQc5TkD3XrPW+t6Jl5KXLNcFlX7PnOgw
tImnyiLInuN/REKm52yJA7l6qfZBFTGIsTIdlTql5q7J7llLmLkvwVIac+wmilLd
uhzG0SaXbMs2N40Z3H4qZb8dW8maHWBH49yqERgs9FB6NmMbHmb8b+xjy5Bf/pc7
okQBYouD8MG1RdZ5P5SDnAcmNrBRRHzfzZOtPSYUGNi0iujU8dhSwehYPhvfleco
PSw16T9lUOgnQXR3+sJpOvXXpEkgPjoxE1NFjY88PaY+QUgLhH+wbvEkZwdf4VOl
aMeffm4/lHCm8YWkd4CHhHlFGd8wP4WXNQ1M1XVVFggLhk4iBTyijsIZeysgqvnT
X+CZqhSGEbTEeURRNz4YphYD9WzcFH/ECASlX0MR7tCpjLAAZV9Dg0kr3lADdkIR
W1loERM3t4tCq+oy4+I3J7pIz38jUBHh+XclDjbJSVungf6MdoMf9DI/6UkD46fn
Y++x2fJAVtbOmPJ29rjL81c2mihKUWOnziJXspkisEN5fzxPjAbMEHVS5kN9opFT
H6DBxwJpPmSwXX4zK7S66B8XQna8jhCUZeoB5JqQbgWiJ+q58gXb43SneCNVngKs
QG8XXlN61QaMLkHc4oww7FMxGIJxlxtUCqqIi7tCzbyXDFMzy+ea1Hy1klxNdjsb
x66rONzaH6j812vppuQdeYEBzPFw5kwtEZNICbxxVCOjVPpQWdSW6TSaPii8GKVe
FCejXhy+10oMZPfc4bKD3tgZ/81godLsL5cdK4DqAsU/q0s3XTZpCiqXK+/ktRuX
UJEIRQGbLiN7LbyNvEyQOPm2fIF3K/VwzRe/SXde8hgNJBStsP9HzhvjNxQwClVF
qdP2jU65lUmlIdQpuTi9yLpUCsmBAv8cr9ZFd3brABazBZttOV9z0VqQX9ioE6R/
C95GAKveu6R0p5NWdsC5pPGRxPsFlcPcXZKL/bPXWLBEKRKzkIHXYTIXYoUmnVMa
ICxnJzoluDTZ0xEQ4Fw3MxPhN10bYjH6V7i5xyoY2GsBWCRBJ6v9k5EMnob5hZmU
DU//P8g6ekBUkqmIugxD2PweRqSUQJby4tIqpMn4tktabIVswkFfruNcnLHld0lx
QtqWvq7nswz6HFpUhGNny7p4OqPPRMnDxynxHAtwymxVKSxV221w/IBwv5U2hiKD
yQIQtw8o817MawnLgUu8Q8/G3KoC3+0jCvbBxA9H27zj3Rq3KyZnk1+UrIF4SuMq
KnWenV41iBlMojnlcnezQ9V5iWgbp0QdH89qvPFh4EtsTHB95PNpvCcsMDw38huL
jx7f9giF9NoE2zENuTRfOtUdWrfETuDOrFiSrPBJQ8StnH2HuFINAsqdTDrhXcY6
2yQOSDz0OtPXSwQOdd1HZOZSuvN3qzZ6QH4NriTS2fmCwNXvw4j7Wkun4D6irZun
U95wZJlKUjuWPSsQtQxFb5ckOVobZnyBL7mccJ82jSX2VNMYi51pNbT4Weulu5z9
mSz8oSsielnWWB3br5NZLvuNZNRuuws2p5U2iQ1fnZ3MBJd4M8iAJoqNDve/pUng
9oS5LC8ywDBvvS0WAP28MdX7C6PJ/gYk6mcimOfXkfAk0rcOt+5LBTHJivCj/LJ9
W1fXZZpvlKmy/UEPC6gscPjzrTMP7LiF6wvMvgcABybOolcVaI5jEySeojn7KYlW
aHcaIUEYUrHx+UxKkD/evXL8c6T6YQxodTNX6M3QucOcoYFzns34XqeRlQsMxtdf
bmyEEqDD62XcfQlVTN7wEF3kh5vP2D1ySbusGDvXGBUCOz+wQCSgvG6Hc44FYn7V
r2v/2xZT7O+XReM0a6xijCUAaccyGqdpRq7hFxVse1II9sqIi7WDjFNVUxfoyQ4m
oxNAuSngBqR7HKtTqJ21j6B9Il7MsXPoL2/v6a/5GcbKm05WOBEALZaII8fgp7gB
VAy129O7AsM19DMVpTeG3ONBcoqQmsv2n3m12tT2xI9uPPmNjnEUk451DVY6t2Oz
I4Oe9QeYrq2dAK3bxYbye9DHrZWRuXL4jIjJiAkzvKg0CQxAD8Pl3g7qiEV2KLBA
LmK/ypbnpU9Grtw6Qz8Tdx30k4ZJHF15Qry8f5kdlxOGAkyogxPVs8PKZt9prscP
7lt8RM2JxqZx5ohJDR9FJDsCH1IBJO4YYaYckSOZ98m0w4/62DzeI34ORa/DcYCw
XqE42h2hhNkwVem1IX3KcApbhhjpmG12/dCNGjnHVZo/kPWq78Wk09xgHh0BiSSg
0g+7qY3LN3fj8YHgfMcEFstdayEfLbBGoFZF18xi4VChsC/fweBOYqkEcYkvkqoS
tfe38/k5Am7cib5i/LrecOny4lLoTyVIO5JyNqCEeCfHqrTT0IzpKG6b28/bJlul
7DXmUcLMRnV6k6P8X6RA9lBCHT1TKj/6w9ov68gamNWdohyEqtkamosuMs/Lw30O
nV5nQJM9EloenQjF1io615bjDD5xfzEUzvpVf4nplgcKVs3i01ZXg/ELuv7FujPq
B+32ZJCKSAnlx7yDvhsLTg8/1fO4ULJUMtLlyNhYJJGGm2IUgNzfFSPq9T9dbRaH
y1Otc1Q0vDDK6n/nFYVkW6FUlBCrj3EsTO+ScgHH9a9TIv1a37LKHmWlCYCnfqUi
HzFoX+CyVISsxctjoE67RyFXAL9Uwm+V5P9AW2qef9kKygLdLwK9EMdmFxksICVK
F/Hl9Voa8E/aX7CMiKh9V/N/bxE0WDNhpsQzzF/KPTuSH2InAoRzKFZJQMrE6bGo
pcrK4Mr1WL3IqHOHIUBk7IDevdWmgJaMZDBeUZMvPPJz5dyv63yw0GJMVnD15j75
XJoFhctHYv6aYAFuBRVJn+uVC0z3jH7n26UQc3iwIoVWt+z1AtlC99Sx6UTFQ4tt
1M07gXAXafAWdHXImP2euZ17o0aBz/U5zsqLNGIfM/p1n9gjVl5c0cIgEs63QEpJ
AjPKsvfaWlejYBGMSWc/9gnJeFwUJRqar6FtP29mMdG//czfSDlXOjTB9JFIbU4s
KwTmFmIWFipIP8UtrlvucUwAcSI6w1cWvE8VnoTrFZt+In8SmL/iM+Jy6uZd5b/v
kDEGvmB53GJlmpCbfaNtHQXmsaqafub4/iF6jLmCYadZNSJv/PnVvpEX2VOFoGfU
baG8bQh8S4F9qqsoYhpzVWdQxLKYkic11t4r+8yAxTqOQmt/U+79tK19+uCjCpXm
0CRMr1ugzQKj2Ihbv4coDSeuBi25tWK/yHA6QSNxOLI2h42W3EE7Nys9tEX3JHP3
43xN8psvDjXQhNZdTLN4k2RJ15jZHZsfvsACkCRzryFTOBt/5HT1Kjll/HVewUNa
ho4huqoHyH7UYC2tC3vwoR4xwpC5KVRCW/CqfiXFD2Ykfvqw9Hx0xCsHKC/3KDgJ
vSZXseV/f7tAlrs2lXiqpVTgzVVKxdSm2I2bcU+q54Yn7YOCAT0TxOphgRFb6tF7
NMedZIUqCA6Xz1NbfU8BkDmFtck5pKxYPtYut9bLkbW5/vUNhQgU5bXX+3FVb/sP
4NiQ9eFg5IZ4ea2ZT8C4sfEQQr8Onn/MfJAkdt7ovgvmu3VX6MY4DAfhezC4YCGZ
1xkpusqXhFGzBOTZWzGmkNB6UUDCMzVlYx82Wme4Eofzd3U0VilEThB/1sbltqI7
TRAylC1jT2FCNLzZAvuyWR4tbj59Y7j+QwzpzrFDeXoiApt//80NMSBlmcoY4i0c
xEXQ14rlK/uVPDAoVZpg/anz70mCGiY8oPr6ClXWJaOoyz2PTNmSMB3TmICaMLy2
RjCOVG5og0DaCQ1JBCt6ck2KflIeiO+m4cEksoOJZbKQLlfRPiGL6/VkjcO4gj9u
13pIOzWZzci11JKgQQmgVMLrXi2JLEKWEQ25LZDR9xq0UZ2EW/kMC6bU3N9B6E+S
6WzqsmmvW/rE2yjPvxnXiwLuyyBtxEjWvJChEkWIUSOEU0sArPbOxgkM5D9nW8/u
wUdTojZmzoTQwT0KnqKR+65d2KyQMUsD+KBh5fJzLEAAG4rOoNBHkQ8kmVLCeJTb
KYQ7NPB1qCQ1/AMXNRTvI/GNpyuz6tltfnyBuAk//O9KNWjz8PRwcw1ngSjRljfY
f8ati+zFUUOb+23fFZfDgesgcUDjy8bZOkOBI3nhiVmkTBgiwLki+y/ftzuYNSbc
CsOQZAFDwIsncQQE8QW5vV0fCzUsfQZxzRwCPterDBzOO42OAf3XIll0GO8ETCUR
bql4iI9QLV5NHEGKQsxARgvuHhSsFOydLa1G+8zBLun+ntPtoSbk3B9Bdvrww+aq
y41tQH5LjC1OWiQm6Fnb6Gvlhpx8v6YyZWRoX5WeIB6ptxUuClDn2HJabwNRQcdU
mv5bEdpD+fmiFxx/9ta+VMCyxlhPwmqN83ndPsYgp7pOi8spO/8zXNr9s8audqA/
3yUaCFzAZh3Zvq1FjTLSSkRx1vfiQB7eA/7p4pAxrJY8c8O1y71wTeh3NmrxoggZ
Av7V4Mr5wMZ0MfHYcw1mgwB0kvJVntq4qy9BaN5k3uZqWxONRImJGws9I/tmX19S
5SEnbImMvxI0HvrknYUTZP5TPDmulRMFD4gqxE0lHlXV3ERT74/LKEkuSe5EFqrS
nfqCfsrLr2T3aCsk+YSBu+Fc6zFk8T4KXZg4Gwnd1lwsxymZQ/1TqTIUFMFbI5nU
t9ufsj0C0XN024bsynfAjUCDxEL1JUGe6ZPevkJcauFm1dSL939pIxku/uftALfP
wALbGvgINQ3yWh3q4ZWM5SmmoWrU0Y7MabV3OrxPRwUhIcajN9k6XokquqDnpWX/
pH6Z61X5dDrYQh2mg7/NUdjaqSgQWIlMrrc5nRNOtdguxx2UjZHjuDVY9C4ZFcG6
hmn6GCdtHlH8TESrTT1FwUqKo1xleXUn+wN+jd1GrpnNPFnf8P5ZlYPRzOV0Z6jV
7GbAKNHoXOfXzFacR1SCZnWxHB1gTiH2pWMOMM454HG2o5uI9j183RD057wDq87X
3WmXkZZBRnm0zOZCW9hxT+0rnf7JiL8o4z7vZzlWRailg6ZhcVXlzmWPxLjksvfG
pW3EieqbiQrW5VnmyabUz3rZjzBo5VzFlmQLl3KMR65zjwX8FmKBkX2c3P+5FYra
kvFlao+xbWSjoJmSErPX2EIxONjHV9TgCQ1u9EXDpbF8Zs/hVev0iaAobyMlumIc
vnrCPWrFzjg4oW/iR0+ZTXPo6DFm1ZZ4uZyk0DSCGoOopp/hrpyeSBh7MqG93OPy
r2r8748gTIz7p0wu6Vr5n+UhnfOAjUnMmYIzHdYn89tOPVkHAv7E+S93sGH98akl
pqXs5q/z1iWJ7EkZtEVt6xtlcL6W2JgfW3vH9OfqMlR0lMxkQh0jssT/u5TQaNSd
jgSQOd3KSMdVyJ36F6B+SYlIIs9XBOSZ49/SAQUGBWA+FAPJs1W36dn/Ff3gejTq
zG47m+S6haf0eEJthxMGKMAWnIXm8BZDpMdEJQk8kcViqHwL8nn/E+Oz5Xn+Y9gn
Z6I07IzU0YS64ZgnHtlLakUyfeonvnTR7qjPLORD8okIICXvrvDxIUdsHU3cqVYA
zW7O0I9QZ0pJ+Qv6lpeAhT/pA6C1Q2SLdRH4rKZp/64XX2tpzdhP2eO4wtjaVIIH
osP9t3zfRw+FcF6qB7EBRuk6LIQTJJp5je7TC3YxXQgGnBBjyWtj52dGggGZTCsD
6/tLy78gB2Ndo1Xlskt7yS4vwx9J2AECj1xYp4y5l7udfbcO6wk2Wlk5spbR7R8q
CIm6xn1yFx8iMWuvFhmpq5rfTEyG1WeI2QFlg+5WEO3RRjYOxptjM8XDWrWZ07ys
dJBQviuX6+8D3Qd+zA1e7qD6wocstac22+IPBmLKgxpKwvwp3+yd+qHlD5UVzO1A
zICXgmaIWHefO5BgboberV8/MwhQn2z8vAofkSWdIFBc90K+ayI0kZLwEsMBCiLD
cq0Xb4puhFqHiaAQMq6OnLn7iRqixSGTx/LjED02+ed5n8Azi5oxV8qVbt3p40fe
jYI9LW3UUPMRTb/NHzAVWux2mi07HX2sF3wOsSsvWDAKUkoXjliio/TWYBQaIT6H
FAvJNZ2YBJgZRE7oWuLQhWXNNXTBvd6UZ9Jk+Y+HR5UQ2k/+jd2B2xK2r51H66wv
ljLjdOGvcUU+lASbatqVdIrKyixIAj02A9xWbQZ4LHvlN0kqwgJ4MQJz3fgLDN1x
GSb3JAPFp2sICUxVjAf5AQjOJ1xj67auGvMmXE6ghSLqy0YSZ6Qi1b8Mzs31E0wm
XClqVdShW0ns0eRNuStw515z+uOpQ51xK1MzbXfTuUbX1r7BUYLUlHhw+2RgP9cM
LUHvcgzAaUcnNlxy7fQjPkAh6ZSxXCxQxyZ5wf+Q98MNvNfryuZED04CRlJEP2fU
cqo30C/qiIigocK75jtZ2ze/FqocjxtKrFryV8YAJuuYXxSTARXm4gzgln5Sehq7
805VRH9RYVU/DhK3YpVuUcJFXtSPd3Aosf6H2aV09j3Kzue4C87zBAabktQpZSpZ
PRn5dohMdlyK4vb4UBpVMLyxoW/2klA/We8GeJhyHAWnuooaZH7OSwX2A4qJJ3q3
Szoi1D9QzoJ+jZMfAFk1L4BFYguETEIOoABgW+DAoddooRG4uqiCD9a9tGPoBxvJ
L2zjTJ2ZDgfSC5p1izDPRLTdQRKVAk2D34yEjdcF5wdWUTTG3dZwhtlp5ISZphsL
zJG3XEFiJEdNc3opjfSoM8U7zqljt+XL67Yw+uQn6fIjP0eGEnKucQs5N+RA/mDK
8NaGxoKaO2cpx7EtRzHhcrg60nOW10RbMyOTHM23S5COWAbM2vMzEr3yAeR9uUw1
97F+9WIfjE5xwFsXST7uCz1VUeIU2wIpd2js7exxoGLecUsfs0TtfceYRFuIyLG7
t7py2C8J4sbVilVUACm9vxCPkGHGbMUhuPZReOE6KKsSQv+Pag8Tb1mxF915u1fS
Y4sCyyoQy2T0fjje9DrtOtXHQvwWOVWfcTuW2MrzYfPk1qOmrjBhkTfAgFt77+Yt
6lUcP4nw3mS6TvNDp7yedBKyczhD8LZ3Mqy5YuhS7c4KpZqVCdlENNlyoWHJZVWZ
JRkPphkwpyxB4PZ3X9ro5SYR4bTkI20Cx1ZPp6N4+x1VbhLjRZsLNNNnC+o74oQm
7MEL0aGdILuJkFzZiEjahl3yr+LslQsy6+sNzoRiiogJSyVpWRxuOkRkDC3ntGRa
wVC/vP9HLMOD5+4YbEFUUwDEdxak/hAD8qKmUbI0hmCQpggFBPINjzMLVMRJBtAZ
CLHnUZCkVlSsK9UnRqKKcW1De36fol0HYalUIYUKql7cDyeo5IfKV/3jsR5562Se
Wojc5MAjnlCefaCE9tUsfELGHT0KWdaEpyS1LShoH9s1t7mZwitCpQMIpxBd1GCr
Rji1K2LZE2diVHxEkJCq3rQwx/vmiNKkhuf3xuF12AGihwFJEWtjhiG3D1n0KXWZ
lvQALV4Dtk6l87OzWIRxNPZwqhFN4G00PC/qCL8RoBEpBcV4zRZuCIV8wAfjWmTf
oXe02fySG6Jycje1edOJmOkNF6Fba6tHZTuOqImKhM/goRUNl9Zw4yhO4frh5x5e
MAG+gKrIHuAjXv3kDZXnVaYl2qNDfZ1PvX7Omt2gY9t1w+nXOC2QUmNiTgMt3KQk
4xi6kuL4wQZGyPEFAEl8NOR4nvbQimYurjbjIquUKguQfOe1jk9zQf8okO9IjSaw
R/6BVTboSwKajcHXzQaYcqgXcjn7GW4aXvjZmhB0wsT5V5hpl6+u1kiX2xESKXFb
4HLFZf/el0tRgQADxx8sz3RjJG3Fmpl9QKVy2C3zFTXejzEzJ0Ub6WPJOkewJIHQ
iz1vpIghUNKVIZ2GfdmBESfozxPQLppOUz2+b2yvjCrF/9DurvOJ68vuSIlj+bvO
qddeIwLrdrlXQmJ09tehhGcRHkR3tV7MJhEl5C0xIg1AUIFYXZEAKJ797i567vc7
b1zWYAdYt3KmuJiGZwdTqRU2tfgQo7bsvtOsOOGHp9Lu/MbomAdKw2ggR7YPRCu3
dtuyAG0tJS5sC5rHHPl7sZGhsjqRK2j4ufc8qIMxVcQ5xBBhlRXwRJz1rOu/5aY8
O6uUHGkqd415V+kPi9XHK2ixDp6M0lIuaTuCIR8LLNM/0ntJI4On2Y76FlQXAlsN
BxPebWGVQ772HdXoW+A1VDnwnlBiBZo1zZuO/V8g2ohlIC444/orueESInZeCXvr
Jslsz2UhcyY+FPGr/JyUnYv6d5T6ry8WAJQeqEWK78XKueGdv99POxIKc2SVD3NS
0Yw3jcwqee6SHAg/lxxb0r4GlBpktGRR/M/R8mhnM2Sp+4g6DYnZvuX74W8A/Vfp
4C0Ws5/8FSdvLuYdwtKDeUGIvXOLjUYaPX3055F9i34Cm+/u62x6gzbYLjoSpYcn
N0AjA1sSFPGREpWKgt44lqQBOtQ3V/JAW3M9L4hIeg+/dDg4Oruxczrelw5JSCyx
pMS+Go9gSA8yomoLADvJBzAdxGja4eFZ0sOlsajRmuyyS9MS5TjU/G6+jtP2ltCC
N3blqTd12Lv2Rqwk19kcnnD73hADyOLC7vWG1wQS0tXHTygAlU3Fs9oxjBFfz1qh
XQugKlk8fFxeeRpXI+aVa1QPc5Vz+x/+/eSQw90zUfjfhRqhu0tovUh5e7pVMMe3
VMJvUYut/ozgM94Bw9nLeXcRNThIIsDltkbP7wIyDUsoWB0IPtclq41IDAa/Spkd
yFjEFr8pm9aQtfpLoj+LvzWxxAVVR4KWtWAK5xZirxUTrtItC3ENG5F9kKRS1IN1
QkEoMLmKmFYt+1yHUyHesveRHaHdeugEAunbK8ugde9cGhVN2q8mQcv1DRkdQtiG
F6+I/+9SwtJnXGPsygzyG0QmqgfDh/ynRwj/2c6uNRbwh1b0/cFtRcHoDUpCYHPA
hvt3ZQkzevc6sQOVM01GOLKNd1I5AZN19NXFxP3Ckxn9Y6O7ufnN31kFvejjmUVZ
ZVJvUomtSW+0vG+er5RNtkQbZrcNHp5R55NAYh2YwGGeyrCXRIgNbtUdErUe6tcW
vXlSiXKXNVVw7N6ZYzFl+1QZDwN3rHyGezmyBNWRjipcQiimV0sLP9Yq0JCS/EIR
SnNoE441sycohTSH62JAfmgw7QeJuVTu/9QR4QlJoWMz/NPf4RKdSWr4D8kRzprN
FcAx2aP/E4H3lq9QLVDS0wBa8O95fdW5ADyze2dj1tR36xMxkkqLhGHFZrBH0jW+
IOLGEQsPZYYmKnvPGEs52dPVW/eFD13KlS8Mk6mOr86cKIBBh10rAiSKDRKJtBJW
SCpwlfzrmP+/MVIBqwJmgs+FIhNd6e74a2aRbl77nuL9w1U9CyUAnIABftMyPD9w
XMlH9/kz00gELRD3Uoi//2YCi+nN68MP0o3b8aKpZ4yorW9lS2s986FrybjtEJ4n
RTZiyVlFNYveO9EIVWzcN2SdIhGPzpwUKit1zP45On67ACTWQ63kY6iQtetwfsJP
KcYDEituXZBvfP/NT0AIlXQH+QWxhhqrLjn9zbSJQ1t2MhgeXkW0MTEpBnPA2Pt3
KhjE9gIJxwUVvt3V0l1Pptniv2MMJyN7pPMMtIZ8fnN1K9HMGIjSlUaeE+SBOt25
4AmJGEhbePkFYgWlgEru682uCEo8TOH85XbszgzAwEO22tsiwU6yMmXbRj1056pi
yfo59u4gv/UUR3JDxC6OuinaYgmiPkDbQ8NIQqfn6mZsa1Uh8OM81O+4qt0HkWkF
B3qhJ7fcuTCS/6bxMd9myPDoaU+cbOyaqiVQHM3fbsX5vx007Vpz7IdFMqMANcTT
dPxCBmc4IIn6NbcLc6oCovevkMol0xyomtwGsIfUye4si1kbdIuB7HGYt1e3WDRp
/WERJZFTho8lE9VVYp2J5o1pIgUbpI0NIlkh/y37ZBYp2a6mwIx9xbFuRjKP4usH
xjBvWtgnthKw1f8JFNmvae9TeIHGDowqks7q0yYdMe/V3QO3eFahAiE5wyH3p4zL
t7lWgx0xBwbezzhpJF0+tjwdOXHvRm5WmypKLXpuDZ37TFJNztDliQqQAGpEMrHa
C04V8GgnSTxNGyM99YfrITX7bEJqvB8nGSRPPXwm7VUlVWRYBw9mmfnf/gDsUQkC
7H6pxSzSsxhm/rMe1LBZVqmYVafXOCFkE/Qm42OAIDCmNdIEAB/NkZGhqK1iXpNk
FRlEr+SQjWXg93xKTaQDJ/JqNqpQFycxpvrBZ6l+dP6bfAcox+1paFfueuCq/u2y
cmi7f5Htu/7BxhFPuc/UAdQVY/CQdDKqrxSCFOLlszEMnkV9QV84a2jLbPOCy3bJ
mhSy4TgunIrjXD9yY1Z8w52ypj6aLsPVIZvxK/7f4S8wHN04+3SR636cLqrUdqFp
MKA7JXC4WfUtSb59Z7v9bsz6GPl/9APbJP+17fbrJrRC48eix2WyC+oLcAC6zgBK
giAfWB3CPT/962+hoiXxXrlNUcInx3zsCfWLuuG9qlRZdsAdBW/cnnZtilhoZK1p
NC5yvjgWmXCuX/6Kg+aYViz3hhYwyUrikll5iUlyjDVHZD3qACxi84Pthq52+OkH
Sdk8nl4IhbMoqPyPVjFqJKUuVYSk46yLO4j0+L0qhcP5QSutQ7/7J+geLJTqpEpA
Q7IJAm+AVAVsBjh6asFBvz+u5X/csmkTDqFf2wWcMsqSuYB7NwMHPLEl7Hj5OT/T
T8vk+a1h9J+sAw3qsuRngrsosUwBP/mXU8oMi0bAgwnqTxdoBFHSWnF45+QMt6tS
7c+ptPmB5Te8p8gYVwQH8ZAIhTXz/ydkE1tkH1OVap9CEi1FiNjZAmYj2mWT3mJH
7GrUp+3K1wPM9cFcol+0036RawO9Wxi0NhfBExqXAFGZZpTV2q1Xp1c9lFoc7C0W
dyJda0WnjL5OmI7j2ictNkLoHaVayNPXTBhH/+hcvTs2mRMeWwbe8Lld3xlGg/di
scBhWXl5nNbnYtn1Am0k9kxJ6r5NhbpDgEtZeVjsCa9PhiN4OKp5G02vwg2BX3RB
2SGalq1t9pDEJTNiFSBPQ7ziKCFt0lAK3u7Ei6t1bqY70Swr36WmAs6Se0ZAd9XC
k4aQuV/e7XqMHoLuxjvJ3VJDoX1O6fjKiTlBF+TTO0SVaIWrPIsd8SeIv1oPdJDx
h8DyL+YG9CZkpYfkWY8k18JL0eCkQvkGq4pNNv4ZGbhI6TTyjsTw+zYIcVeIYmB4
/tLPOgVO3QaRRKdmxn3I1KgRCbn0AgFW5rF31YaJukWySHRd+ij4BxPMFOsaAnUa
WHko9zgMfuA7tIW6WHn6sMlhQ97oEgcNRYZ7NmYEfbecLaq6/Dtypi2DtsuISOj+
+gwTpvk9N2MiN6zodEtq7SKMH1OrBDNHCQPWemfZV8ob5yXTAlU3a3Uz9BPzWqzJ
6mF6xyxZ5ERwVWoIqctZKJNEXArNUsInEJbZ5G3HX9sRrlXlbVElL+oVmEKq4auu
gb2PHhlULXJo6Y1OfemSiRQf3kLggvL7NkmKbnwpEr26hZN+2AwUMvcZwFhMhWX/
MY7VkK42qifVbYlNkoWPoaYbRKBRVuZq62c1QwPHmdnlh1tJlaNOEe3cFQHwakTJ
qEbhpA4/XpoS997AZLG6cQnvne4jG17cF5CjRLakpK47o6Q+rnNj18hE5SG8sRa7
1sbJyjhaRa07gWVpWJJSvkOKTl9elMcHbCgwFVoeSVow+89CLF27DHPywH1A4+TG
ub30IDM1jQjmAG28HEUGzAyNHbXX8YJhjx0j9puTL4xIHeLesUwgPkCvvW3tIXBR
qGA1uYZX3uwRqbBlYj4dSQTJdEmubSuz0/lsyeqQdZwYsmmYPbsEDowqtByjSZzN
PQOak57lSQmQkx6GPmCkxEXLH5nuEDzQgvo4Lz/Q+9iZyKFzEUEyhZKXX0BjX6sa
rjhdeUMo+JDqRnD//W3yMm965wWMGlTQkfh57kx8slanZ4eCptrIFmNjiayZwFGW
pkuu8ZfwoInujF/HeIAo8CJ2Oq5Y4uZLY32aquqeOdAGEVdppDMxjG0Kv1KUzYlC
Y1Y1NPNNpuXkMcgrM0qS9R9+Cc+qi2ub50dqe7dWFUWonwIdFCKU8vSYF836Mmeo
daYyRe9vkibSLCVu6dsddC4bXCXitiDS+bQxh5dwkwPWi0xmV4CdbnJubds93YVQ
xNaeMFDfeWMxouMN8Z2gzaL/5tbZ5S71Kv+tOTiLjv9TxuoSlChT+hlelDzy+NFm
aZduOTWC5IGwx0P0FkB1fRnICeRunhroc9JR/4mbSwzFgTBij+7elJjRtuJxw/m+
slNuRhF/YqDmyc5nshiHKcEoGHXWgwnh7rBpO2r6WOzGM25zIMm7vaNUf7uDkpWn
718TggTZB1FM2ctBoeKiEBxO3O6v1GslFZC1MWxDsmmd5KrC+jCXKXBlLY45vbgU
/nd7oF9kpfAJR0OkOPEKhj4XJP//otlr9N4nAy2cmZQkX68JtA6rE/Zzb0cqz/lf
753HaeW4B6Y0SNUc0fsho/nx5G7vgepmp4sABjEUez/dZT/s0j/IZUZQpMsAE/q3
K9R74hUv7uOs88lhDxIN9Ckv+hMi9695iKapnN6Ght061mdu7QSXi+EZegLMe1Pt
yTC6hP/yHPwQ7NCei/ZP1bbi0T28xyTJn9ThlWttJBamya9nINn+l1z/cm++vKg8
shOpooKp0s3/p0S3/y/sy/uP9QuSlBAmbeWdwweJrlg5Ppjsg53YUIEPgbK/7CQe
InG1uv93y27cHmp74xNqlJetLxB1tLKQy0+ZpGox2r2Qjc/ucG5Dbsmy5fvAvmJN
3Y/OGfJ/zdBL9SgbxN7xY8AXIyHD4JdvFWUmJeXedvyO21gvCR+i3y06dKhbdPYB
KsioMoC40zwD7aCTBHtF8bP0gwbSvFJ6RGC3eRvEHu1pNXrgKixmEdAAoAif0jMn
9AYRKvRD56/tvgWM1RBDTmM6GG8vzdvNOfZQ7CHhdTRZHAok0JCT5680NEgHrtgz
W6jrz1BEU1ADexCB5pcK/DKkDnC6wQ92tMFpNLXYX4pI0hHPSEj4kO2rGqc/FlHJ
0iP6pipJiBSzS7poT9AfyZpbffQtEz6UIrpPEl82YDWAt9Y29pyyGWElHwvFdtpt
tg73H0R0qN1qW7IOtOz1vw0heNjNdm9syvQCIf8LWaK2bY79CmWHpyVXX4Ien8Dg
XzppXb+uFBDWVMy1BshgI2ZwMd5WWCOGnzaqiVvB2aDMXTsIdyH6L2ClikEKIxA1
QphFMfyOPvoMYHUcPppfuByzFHctzlctynnjcE3l4TMCLqUNu6JMi7uaC9FCJIcB
nS1/e+eD5hVXpVXScLJBLIYlCiLkqDwmFw3HpJHUgVbiT01vJfhItcU3SgnIANmX
cbCALzRG+cju40SkckGj7Hr+V46uH0Arl5S3DSPcd4BYsQY8ftQq2106Y77Lt9Y0
31tsPgDa+svtalnibXi1JXgms8JaeNWvsLMy+kYFAM7VFECQJhQx0c1VQECthcPw
MAaB+gSt2oGvjdAuXwQpltu8cs+NodvoPw3gvv0Geyz7oU348MS5nxFk1FTVMgjX
KNFVZZG3BEh85vB72TrBdr1LfGtn5jTS6NHZB/UqwApmN68bKY6bRqhKtN/5GRaN
VlWlrCah5iQzrltgMFWc22UuUDFK5Ff1Fvm1zw3n9C/ng5e4jAXvjn/OfO3+68kR
5eMvwF4LtvSDXnAZwuY48rR+9vZwScEzCuc9BeNt8d9DN2srs/BtTaisoArhn99Y
60WY6NwNpLOvZvoGCTo3ih1v3RuahsfnuiI8xkBVtMwcMzCxBU9B0jYnHpkrlaxs
VBiZUXBFC3NpPqBi2f5BrxPHjzj9J/cppHtCb1KqHaG1Ib1LvuuIbrVH+EE76opl
u75fg4M6PKaBspHp2v9T3dNZXo+Mv7sizkHMgSpckN2H8IXKOji3nsos16ou4rIi
EhNbnqV2o7+fHAj5c+MBDz7MyLks5C0Kfo4mD7tm0SaCStKPz5lEqGRz/Aqv6wDb
2IPTSETyU4888/GUj+EhojluD7J2DpJqXwu+RTwgGmdklVsRtYxRIqeq8qk9JPGW
ftgUOlCWNFOj1vzKVJ+Xw78w3wi9YgV04eFrIl5yU4UlWEak6NErWt8tdeBXBLRZ
sy6wNyj8QliSd9acvZ3g5teF2yB4mE1gIi4x0W0MJH1l440Z5l0PxLpT/E7xF16O
1n+q66Iw7KuBHPtIAt7eSUK7RS6xKN1us6OjyY/DtzLYlQVZGcHkZkAYIdqpHuU0
vTF5f0vT6JnZrf9QVTvNhJlKYvSZtuYjhOtSZ6RhJHJtyGoIuDHdmqTzt04id2aW
pUTxeNDVWDyMeAZk0J+RLty4Exkq7PSW4RhK67/q4oGckAAzLDJeyINvKOMCbLP5
ASe2RzhNTJGQ7oaw+duymVuD7cvParJdFdCCGDtZTh+wl5vHDJu2bIpONNBlvTqi
SQgg/BiFzMQWp/ApoLdXxahuOtPCYZO40GqofM97HIjcXjkr+RuwVvdRe8rf63LX
W6iwTbxUtPfRnapx54iQygSN4Xnp0n9hdfeNNALTLeBi08RaiAuKGBqZfkh1E2QM
CBhn9exPQq1c4SfgUQJ+NaJA6L0j0inLL8Ylm0Ot/gmdIWXZw5rELWv9QdGKYPO4
MttqNqRIsZbZHS5XWY7hWFgP6LiciigOFm2PQsensUy3lZuj9UoJvRUhi/iC7w+/
/pX0VTjxJ1/cciatcsmWyjbU1U8YhYcySLznLRi4v27PIuMLC1JwFDU9RmKNWBHf
zi22eEus7FFwrwyKDc6sXDE+V22QQSdtfne09FwFPJv49nk72j51RZ3UBlZhBZPP
LmF9HsQibqBI92vuUyqYb4Q+BZ08PInfUgfHWzd2rVSqo+NjHf3vLsZE5iditAJm
Eje2EHCeAqmak2mr5Zbl0I8J1fWroNHBkCSGShcRDsMPp1wblz+3NfsC84cLLrJE
L49tCgWv13BVjBH5QM7+Fknx5L5LCqUZrULHDiIAjSo4t2PepsZwXiudxpnY5sQ9
TmLA9vM4FBKwkQpH6/WvOoWLntuDZytpsugzt9JYn6ZuSD8cF5J9ijOdkHbUzCZx
4VIudCCPuEMxmcdMZJzHt/oZo8glEiCNXxNnq3NQ2IRPC6eftmomZ7OEBO0bnsgX
jf+ZDmHoMBB2R3m8ClvMK8Uil9MOfkgEMsoWY6MeycObUv9Iy8usBIERyKPEQXsM
Q9VsLLUIa7J1+PIYk/GypINzL1fSQnrKOJT/oBYPG6QVOsVYF5vx6l8KhMeAfloz
OxRWkh7pI40gZtAW5vO/jRqAzyMUFhtyHF0MIV/xUElmhb8gBWVRcbeNbGyeAfNh
uahW3D3KOpj3SuVJO55Uk9nEvVRtd6d8ybYuBpE17BtShN4KAPm1+FDl7Nmvuz30
qIUhVDsoSYBMPGwpmU4QXy+6VyP29xwZVOZ7f1cEAPui3tufZKQbF7yZwxUFBk5C
hpRmcB7K44tRv4kXvvgvwpPsBs8F1jNjX2FS1LoCMwBlfpjUpSv3MGxpd+oanR/L
ur/jhgVtMkhh3DQUO2BrrsgoEpBw590r+1iVjg+lyJG21cifr4iNr+IXsPycYRNc
LEtb7HDDeb4zV+WdiTy7MyuzRIiboGU+07qHzXbony4KSS1tqNWCfj4aS8nn2RWG
3UkayibCfdyCsyQcLIZuktRHsDiCtXRol2r+OWF3Lj1RJEAC6U1BX/mtmBWvefrx
iJ6CBVyIFU/QyX7ORVlM9sJxeCwe4mrwJPIXWBg5RHqZaIz8YBd5gl17z1+re7/c
io/dWr56AXjVUgM3POovJ3S1N6e8Tto/x/gQpPmdna1VAmDVauE0bdJ/J1Dijt6Z
7S4zF6u1AkuMHAUzm4IfB4FrpzShx+2XpzbYuLgfWSSfbCCEfq9fDVjuItAsP4Cg
7GvxkP+XPyw6Gv/HoPuinVrxmGl9Ka50bmS6f2XooLHi/q34iowoIV0gWGyzyu85
O1Si1B+vyr+bCKK1R+mpJqCYS55On/Qz0Nxl/rbP03izLKN9wum7lEN5SGqo9Rd1
YvRb4AJDO2gv+aYVxRA2qCYeALE7uPesWzSPSs/RvdwGXrJpEJUlHQmivu5FTgPx
9n0gSfnvhfyVmA83fzdRAnu/MLj++0nV2x/cd/SW902oMFhRWE/j+oACl487tKF5
Jt98+NzGH33lBOQubyBhQIQU5UyDhrgf79CpkalTIEAykcfDjS7p+q6sDD+jt1H7
8voGojwOD1vKD5OViBwUIkyei2o7OT5Kd+7axoYgycA7Aq878z4bpKMSvS9CFnSI
D5eOQGx7DFt63rKISb9zOtq9dANBxZufuGwZGHKn9STcreG4IElmsTzIlZgoNww/
9qLXzFn4ERySxTzbMPI/k18OvlNC5Bg8ORd+Hsq2kHvI9FLvBRpMsJ4gb4mZwm2k
56E7YZgmklL+G8hLG4eqxzxodsJrs+AV3d+bzZui7caU1bC4o+h3hTXaRwMe6Xh8
Fmb1wtQYI4sXSRtBkPBL3TvHVNZgflKHiAFSvooFBrYFkzM2Xsn62Y8e3ynngKWk
9u6wRjiW+FNVsEZxVKi0cTKwSXKgDMtPtprklWlvyLcp5aIUOKFZiNBVenTBDCKg
eSPOcSer1cKTexizqbvuZThwkvy9yctQuSPt710HokCAQVDVQGk+Ue4ZfBkIQcND
QGs5H5a33m4zZSwWDI5RHZqFCkcDukm1s+OUUeTv7mwkbCJwwyjJoVV2tbThI+6S
nfPQV4CQkHlJAtACuVnscj3NMgiO3n1cZncEnigsB3HDUSBSznSVsMyJ+8bZxNkU
/va7z6ht79yKN0VbmAKZOi0xucQhv0XfphovhbzQlr/tE+oE6a7DQ/IG4QPqO0bn
A7BGv/Z89Giz2Eqze5S8Ytwj3xjRxYvk7WKeLRBHScaZfuLqszIKt4GSuJqfetxL
7OVZjb9rWhVqa9X+uOaHE06JsaMlOZZQGGlb2eYt8oOXKm2R0Y3jBQUc4oJE3TRX
qLGY+66HwtO7+R6hf1PReajSvMi2Br5LK4UiJkpGFuv4n1YF79KMaR2Q0nYggrtQ
TGHy2nfAV1H98SCgPy6mC3nTb0aBCzc/kPvxDXdjoqzY/8QRHe2HYkx8HRNIDZ/8
NIsAJVYy5m/fBjQJ8SfoszuCe3cjnHvIEeCDciIZjs/h7S/0uKCVnOY6PslD/k0V
6bLo8j/SIV5CJDp13suOkgI2i2cL1FfpY+t+fWIMkqVnWyrSsQ4DdQ/g3XNu+jB5
OZFUFD7C/nftqBwxkdx8dIkPukDFTO5avRUHgACdjHKnC8+c8F/9MBRohPkNfmw7
0+KLk7dzl0z+gIl9rogIGGb++7QmODVQ154JK+hqUSSWXQxJgiE4UVFKzZXoiH8c
TvcSGwAHTTLedkJJpqRkW0zLAlAAJyt0ScK3MkpdUYRZtC1TvOdsOAjPW94cCGbJ
/LJfiI8Pfc19xoN3crJ66uQoiVA61W6N4gFFSTGKrc8wF/Prw+llae2StNCY5/Ne
Crfx1cNuEfXVl7NRhOrbwt/6hjAwUluG59w9Ewgh40ej0WjEz/xz0A9dPfRM7nsH
onuTB3mi/Sg2v2IN1RCJ/Zu0kTsffboF9JDTG6BkquLt1YvLXxht+RgrZTNazouT
Wt7cp7XtMsqXaCAIlkHreYBIYiDMsycgfBv9T8MrPi3B3ssqwN49mRskOT6DzOOe
AyUlNH96RHQGrpAaQz6H5aaz9qoEAx8g/cXbujq9e1/0/4ROpdvD0WDDQrk4YPhd
NYPpg/WEC8jdNHlJhhmbRtbUOZX3rCti35e8bdYO6kd5jEcSOk/mA1OO10loGC4h
8drN7yLp+wEJxIRHcnAulRTk/o96UXU4WTq5PW7UGDPXIIFAc0b6V8GiEP7jIGE0
psOOvBYPJLfZIFxD2gaL1f80Ue+H72L9jfKn9uYdjB5qjFQ5uNV8vow5nX8Wxnm1
IeAP+Q8mXCg8Ja4Q0tE/GhjToh3GjJ1NoURvYdkB2L814Jt5ZfRcU9vrL+B6o/nb
RTyeOGvt+Of2STCNn2/u6G/VD3aE4xVhfFRD2ZCYhe3B4t7Iw0DpCcv2VlOfZePX
wEtDAoun+EYsrovdKUErOjw5pS2MQ+6jTIqoYIYOwFEu6hSL3cV7ayBn8zDvKXTL
OZupBU9sP+R6ElWv3qXC1wpXcOHq7z1JvFz7zvZtrobVW5NAj9f+GEPqiKdchmB3
U1G6V0ZxUZlOedTxNR124r8rn4DuQk950Z67owCq7N+PS15yh/+ZpFa/dIICtbjl
42NIgiHlDD6yovp8Be3OTWa+VV0RMawX8ZamOo2qJNKfqPD2a+nii/Li+0Q5DYRT
SKRbHPwOtWInPJpI1MTfeHiKAihJrimFfuUp30DJcgonqcjlvvyEYZNY2QcwD8Ke
emD8ycvV/preQ6JmoZxgTMPxFGYUItpZlILbBPvap9fZ4efZDqbbgS5QD61i1Ka3
+yblOqBDTdOaefWE7solplxCy1SWsTzyDKt0vhBQPuNiaf+NjzMFlCq8iX1+mpbG
zQcHyqhSY4JXknrUlnCp6pcOBTfkZD5OkuOCglX9W/RknrXAjZhfgcRcL45oev6Y
qp4uLx0T8p8ktV1HpLZ2PG+GOXZC4fmbAEtk9sqd6awF1aTMCwJb4chsu685I90Z
Wa5W2VHw/ehMMLYT6B0CuVlmVaL6NRGI+3JyVhvAa0T3w9IEqm7UhDcJHYydsC/j
QMc5HmEpUI3FK0vUM2P0GPVhC5gCAxzk9BP8vIU9cED74wK6HBXKMYiSFU2qjAm4
V1+TGS6Cdj9qpD7oRtQyJToZC/fAKofL9PSawJz2ZypjdmH71kJtxbSsf70Ltzck
lc2Fsd74337BcldcvKXeb0mJDHxh3ycMLiXwR1NbFnHBK8bwpLJgR7cq88VX1Cfw
D26+x1jWmfbSNlWJwcEyer82mAgDcG1nXqNYQOL6I7MstGtRcWzrhTAT4zKzrAHi
xFfKoMNV112xkzumEZNIbtXtEKN8OJl4QdWs9EFODLkKtTfD8VggmjD8O6PevQEj
ayggwJV2famIPXeiJyCIS4BXLQK6QjwMSW0rF4p8FwArFQumVVDprEN7HaEhqODI
OL09iQoy6C3jlNv6OK3PJPzCuz2CKmSNUHmnK4E1TPzqZOOrF7ZKEUwg0FLyN4l/
FLn4A04dyoLRy6nHtTibMQCQ/Vqs4Uk4EhUN6EwH6F8rkKTJlVwrypLxi1FFtfFe
Jo4+Tlg425zo0nUKDOsu3oRvg3ZVTBad1gHfuTSKYfcG+m/067qZ4BstGd71Tw6v
J9s7ZpsHhJ3GY++bPyGKrCx6Ln/PV+xQ2f3WUP2NxKj2pX7AdgNOAW0TJwtuJuUD
Xbuzi/yfSWmceaMrnBV5EBEr9nubPfWZ0S+wgpra9venO4lv4MRpBviN8OYAqzVK
8O1mraG+CTyfvKvLaJxkd96P0lMcxw4NFiatWFMCOgc/MoZGmJI5TW5/eXzQ/Taq
FRfTS7IYMWwIeJg9iGXFXGEvJIKlYy4V3tG/CMmUL4Sv5ga8PRFhJzo7uFyZkM/0
W0l0MnuT8kb9J8qIFkG295j8cGxNOPoX69x78hl38Q4x7mESrGpG2V4WUxsxaFfk
HG3T8MNaUtsfELg3uijhSPDzXKZtzHSSaGZ9HTPMggHlaKYZJ4V3/j1yVYkMhLDd
/350EGxPlDT+gNOHAp84R8JQMW/dVOPaxgHyQKXILGDAYqOf4GEAvKyXbncAkl/j
bSIVHKGOWBMrk8vRfuAO93xRhlsN2wxPnyDLUAcYormcX/MDb+ebmi7vtEu1GTxL
jk+SJnI8kQP+YcsppxCgTnN8gOfA6hVBWrNf4rbGWmdzeg1SaMCwiJG8XtjXXb7V
gF6PLL9Ts/iIxXnU7iEQH9w1LPI6OA4zFmoDUB8rl0Rt+mndkz3QKm7pW9nErwyL
MEm1Ep6x0TbNRhXXs3xutz26hw54IOwlhMVirnvlaNOLU8Ll6qOs65zUeR2doraB
YW96ihC/tsTelWTZPn7U58SwzT77FwT3ODpf5gY8FuZSKuXavXP54rvIdiasBVoY
MBNSIy8/XquN4NY29J+cIwaACf4QmBd5hiPxfIw7tshOvnSB673C+MXz0Ojtp1UI
+q5J5jIVHeGePTcXrY3cIwwjfGQ5n8Y33zzrvtTALej0oc5N1YV0YurV0PfrWLp/
vGMips1xq2DxVOaGaWjjCxJdLmEysqh1xQBWHhAxtLi6cJxizwFMdMjagAx2YOy6
GrUUVtmFt21fZZoeXFGZN8gVTF5QdZH8/cuzXPorRgAOM4CwUbMECJVj9BxQOuOG
bCarMsz14Tf3lkp4z8ndUD+X/VmKampcaTal38WJ5SV9ckhOtk2HPdFAyVkV3JoZ
8aPy4QzHH4HAkOGRKCQGJBJX5z6zlFLa4kZn2SsQMH7N2DmngRJ9sZe4XjSIcUbP
s7w+3MZgCg9ryxyenDxDU3BTxA0/fxt7MsnD1ByPSemv0VkP+eIQp1DT/ZsHb3R8
EcHHptGrBQ6DT29qOV/wQxix8OACVm9tJeQN3+BgiXgKtFxDyHek+JLOxekUE1sd
53p9wvDuYhQlCNY7qPC9Z1uVN/6jZIfz0WB520LT/G60WhwLrxofk51MCfYoZWmQ
Q362heAqrHNSyNY4ccF3WJz987nDaidnziycIzRajBLDxgjeUERMVRf1XyniNju5
R56kLdIFfuWn2ngVSTPC3zy5o4XbJMJsu4Dlhu8iuWkRGb0FSIAtqS3vBNElN7le
gh9pEQ/Q8OvO3gVYEEj4rIopftaC+d5XCSYuG5aU8SJLTILtST60cbn/5WkbDuh3
nUBo6E3gQak5HA0sfjtAlCeHc6aXf2jccq4NeL6ETfDEWlDyJqd2pjtZ7HiTskx+
Ym9PWvdDb2XzLa9Rw6Wfv267WvwI35P2Pb7dHPYCFl9WU7acly9tirnpnB5N52lt
87TdgD2MkLOJy7+4baBvx9DPlGsaOsH8XGuN5Pr5apXUMUXU/Ia257V/nTyyep10
W2OINkV5hgdpFciKj1G9UPWvXfSEqzOKkN+Eyks72fIY6zAFqfAp5Xm7tVmXTKtZ
lL0jNOx9zUdBzxVOtG7tlzLejAcftBqdBB9yp8jJjzr/LBrNMvHzqdMg2fWp0DDu
62ppuPl4tGLMCwQQMBnCU1edz1cpb8fKP6Pxbku/A7JgJpkm1SDN2+OOesc0LbH5
xMpHdUOxv/ze4Ufv6g6HI66G/sGooqmUv+RdzfMdi+oXLgrGykgmy5WgJbSiGAVx
guNByFAsiZ9UAgIHoi7pHyP3S/suDoFw9BQFeVVeNgia7WLvWeoyXLGGIa4hqwTz
736lg1ZwrFlL3Y0RSYJd7yU2BRnc11cyYuvB4FG+ydSvt42axtOidY+RpgiWGsJR
hkxKNOi1ENyAXFtoYPCPVazsW/Z9VihXQZmT8lvC/dAAaZgC4IWc22lIuOLZTeHt
0iUHhcXzAqBiq7FQw5AsexjuPAzszoL+WdhcF6ViNa7lFmPHXW2wvfhnOEGy5CvV
UU1JLco8JIHfKvDy9muQSQggQf5jq0KWmzHoohw/xq3Kz7KI5SQ2rVHbPiQdSsJ4
GWbx4xTYKEQ3KUnWWokDttKkkBiGmGW1Ll2TqKFIT3PYRex1fJLRgU12hojEnFsu
4lq1wE3gljlaI7SoaVuGp17V5LMDbvaxj41CyDuG/u6LnZylycikmglgJ12gx3yT
+qU8OfmJ8AOV2eGqEY3ZXpU11Ls7cXEY1+dcoGeayMlFYRDZRgm47+P5T5ZQ5RQH
1aY7Hc+osmAKLy2nCXqjpqP2JM7RE1LywZx4ELHcL7aKQo7r4bvMQfb9eesCLlXC
+X2RT3dX+zWcLD/J5j+BhAXKPMiMjivtXQiC6NJgv1TByVlYUHW0pTqvG373cpOV
XahUWMzW+1HugS/EWYGIe7CVwEPZQClgw7rCK6mfi4RnSAiyaHoZntNWZ6ijQB4r
/O3Y0+m39xvqrgF5mwPjvv7RmE+iWc2SBcVFVjPtuGdpunmEO+WfcrRdxUhGpfgb
gk6KHih0o2oUw9PiTrdGEjNK9fpgoyDAJ3DAGuUcIVx0OYavJw10Jp4yAPzPK1Hh
VcbBRcqosPnS33GzDpMuuINCrqd2BIiN/UNry0b/tsvxaZbXJRlvOaU6SABzbk/O
Vd7dI1yhVRCSppw4yWMrdRHLcSpkrbmldq/zrHw4h067shP0JQHQhYpM7sY2kOJO
J4iGbVjTUJ+gUAQH2o5f5ed6eBwcvCdLphOyPIsq+sREnrB0qju2TomXqyADG4fX
lzf3BKDiCGw9ZfRxYe8DyJG2RlFVIOZ7GqUniUu38ns5lGA/LnYN/AY9Hy64g4pL
gFCvXJxlMh7vN/Hd0cftMYVUqQGJWm4iJAOi5ATF2EhSnVMqB1fUt7Ct1SfptH4y
Go+Tb5gG4NzhiD9td6zQVKK/xGd9e1/wZl3YOIJTU/91o3H+gZKqd6x0czAcY49z
iOuusbOQHSygi9qBQTGUSWItYZPoc6K+g5tXE4+DrjmRROHWowmKJaK8/gl1jCt6
+4skA4FzjxKQXhnTR4zqd58FKIvGHQD71AkVjPCB0yeCC5AAJwSHA4n9ljN/hY6o
GQKabJWsjQLKdHFU8sHdy+FL7PcOn11sn21vn7BQl4D8bVYPIWZ1xuYSyruOI2dv
YiclfsY2xQG2ns1sOf00QgYpVH+vn8jGBmtHpCPA/HJ8B6u7gZX49dNCqjq1BGbX
A3hTpvYG21WPJRiOWB3ANl/vI7dfJyNoiUURFwDMcCpdsIZ7Ea3JD2o8kbAbOPPv
eC1i1eal7upE3DZvtM7e06B8jpAcKNaQFXqx+2IsnxHHqQhAbxZ1x8Nw9d+gGhFm
Qbf3Jp1dYRXM4EOTked/bwSa6WRgroAIbGxhYxK2Bt6QjDPI2PfdI8LmgvX/crUb
uTtzSnZuv96zr7IKucCgVjce95ms4V28KO4rJjU3vgqyO1QOoHxEAu4rOjd+UBZ5
QaK2lsYreKoUsXRV0Pri/eeh2SMyIscbD/z0To1LNwlDhCCopbdWn+bpaQox1BG7
6Em0fvPSecX2X+VQKnZ5HSBK2xqDtswiVXqHRtrRaVJilorbm6WN6KN900ih3y58
9fV889K1A+Kz8R4r2cFAaXWTMfz8Cti97aP4Jk8oXR3aFqtIJ7R6SdTDHso8bblO
/FBvSgDPFnjAQjJmry0XBwWH0KMySZr/kfrinqSU316re7O5HN6eulQboeg/7pZn
IOdV7gnlvIsgdcs+xDnVkzaXKr/CRHsmWNfrK+rtVBuS3ARSLdGx3sNPLWKOImxF
SZSHqlEkMI3v//zqEMsu7wVxSds26NFzhlN7PVWy3VVWDyG7Y4fctwrQSOmIjH1z
vjRRuohZ8NTRTfUwaW2NJxcAjVXg8MeZgzQDQStslucUAnRFOzezSQjyxvq6P5Ru
4w/YcXq76XtLaktnsTB9m6YwBVWUri7+meQdYO71tg+aNhlILIl1OXWABZU36dUB
4ZsliAUeiTcRP5IYUQ7nHHuIhWYgrk4LKsvnXQmt0zzH1whegs3UJ/187VJ/kItV
Uop3hIlcK9rNu00hbRLUUR4ifGIcttwtyjZpiusYr0X+sxbw6om9/ecemKKWIrU3
DQganYgvrukEUMGQnolAK5H5NvQ5rqKyhUP7bvk2AFTSOaeqP2zKFI69ps3PtwLV
G4/jSQNuswp49tPBHM2zVnNaWgJk/2Ci7mmMkNYwUkg0sxgWOeTV6GnNEHTBXFYm
UwYQUvprhjEDnX+dj43h2i5NgeFv597PpB4lW2hJfgsZ2NfYufcOYeG0IaMRT18W
FRj3jaH98lYgzqUAiqr/3nWaL5J1l4XK8CKLMDVgE2IsdqhW6KHL4yBqFlqVRN22
sow7NQjPv8sVJ4X+ujfw+sDa/qhDTU8BxfpHsUNbw34OXjhg/bkzbsnlVoF7aJyY
z95VUK/g2waCRNIkOGM+B+N+GI8nzozazDB37M7mly+AykJrOd5egz/daLQPvoHQ
8IAiAd3fV0wuLDC+o3MJTminces2LRb9biu1iACQAymkiX4Lx4am8BweCsolanzX
v/3RFVH+8KOg+ahJWIeYNwx/antbLln3qUUI6HdQmVv5gKzegoXSsuGlMw4rFNnl
lZxtS5jqhSg636h5LVmtojdho60DZvHmoTnQrHZk4jDW/N2tE/7Cf/vZnWRKhxw2
mL9egUVXvtFnhc274oQn37pzLfqXqizJwSqq6eYb4CkGZknxJ3BAq6tPVvgi75lD
XjRsK8g2EwF2+OnekklmwH+/9H0MXE3vW6ffrlRrN7VjS2jlZoWoYRZAkf3ADBB9
s71WqcGfstEVxU4m4KoIpFAYBB8fbAUowTkijOwv7Yoor3rupooWqgjvqC/VKl0R
xBLJhGr0vhfWSHuQd3J+mdPcNpBej0Sdix23+GNX5mrpdggJLBmheybJt2kNx1pB
Mzky/+CXDv/3eFzALkQYmcLPJbCt8HqNNuJ3HkRlZAywkbKQq//uqey8W5dzt4y1
orSsPnOvlMigHJHh2UQD5SITsoE7Xs0Cbrwey1gHb2ruXISi+5/jq1McAcgnL8jC
XI5G4YptYrh+DLUE6l+KcBoT0e9hlR1JAcMj0ori5jjqgdhbEEli3M0YYScHc+Zq
w3LdhAGdwiMgspNzKjOGFk9k/31s/2fdrWwH8WSzyLNj2ByeT44GWFOyIzzBR36P
dby14De7MfGv0Z2TBw3k/dwHQuhh3KHudFNiJDz8CxmbUrcaDGTAJCzuB/6xsFqa
nZsOzq2mGnSwfLvjmgVheUJHK5HOzKuLTpebnMyuoNYg6Yj/cNdus9w6WSBBguN7
3qK1L93aCVw72nN2ON1roqwYYpLUyxu38Xj0dB7NKqTpTGTcJUEOguCghnUTspiV
cjTYRlzKWTTJWK9UT3SvGGQQWivY/CD52xmdhsyzQwwyMdrlIENduoP1ZpgW/WUW
n51t9W1hJo+4O8eKdiylCQF1LCq9kI6d6FTPqqSTDt+filiSe2d7u/2JTBc3WspH
cU++YNj+eCG0Nsq/09bYOKfvTmBStVLYXSuxp2MjTpm8Ed+8Vo7R7MVOVlCyDmbm
fsbChX4kZ7sdFc5vA+y0HhK884N9hkTeNYMZag0P93r2b1xweRDpr+XBx57YqeER
iVG1H5RphzkGoX4kWUBDIrU/eOhk44OFD2eR66EX2bVmTuPNdqgNLn8Li/j/3D+U
+jG/s6Q4TYr2wJre/k0AVLE0F0/nMqIOuTWIhQga0j4n4s4oBZ/HV498lWZHmrad
Ih2YVo5HxdxrtPb4VEAZlquVNEkHYhEvbu6N6S446WRpwBhmslB7ORdM+eagrRZH
PhH6pyVSvhQ5f4XQ+0tKsUrSSic8Ha3graCPKyf4kyTbOI7Ykcq9u5jy45CU1SYb
gFCo+YOeMGCyHzwdI/dV8qn27aNOVa2b/kC31wHFutsbzklI0kI6OKLWOjft9mlN
XtYcfoEVPdTXLJhi2rn/qtImBHpWscvbDh/g8Ckr3geaPIYq7deyVv7zRxKvG1F2
5uXPWcmpNWpjqdNd57w2nxpqGVQfejTr5SuyVOaH9mlRdWJd2uItD58337/CcXiC
TMtmfSLNNV5mtTV9VahG+xxVeqrrRsjFjsEMo64M36kx/cYI+UGgEnQIrkmPfRAB
maz47JB367RlymdvvFV3GgfdDj/HwQ9ms3q7s871L4maEiQZ4MIlBC7pZ6HUxb6x
fibeprUL/g8W+hf+lXFs6R0aV0hU9LBRkS+Xezuzyo8O5iHdGT+qAEGYq0EUWwOG
p/RgS2PoP5hlfsY5G1h27LYv5MVOWAqNUD3h96Lmj/VtFL8IQcS95s8B3cHdZts5
iVti7md+UzbbXqVykNYLKcumVZmYXl1Uagpgoz3h+P5mdSiup8mgwP05ZgiL/UFw
5PNasnui5D0vVfml9IXmQll/J0d92UaIOonTcpOKWcEyeMP25Yxx7D6kucmaavJ1
HSDCL93VHm1cfzOjW0cwcD58YNKY20oE1dYEcyLDIuQS392H84DM/xBNDUqGS9fK
NJGvdJgP6kUZJ6RRJPcZcsUdZ3Jo1sLlLFxpV5ouoBzFKcX9bYbPHbEJYa8o+ecB
Q/PRaU6Vj1Tr6peQNsC31O2YIl1FDHyXp8EF20OFvhPmsKL56Dg4qYdtD7vLvZII
NmENQlQxs6FmQtSjP9Y2AodvmGE9b2Q1Nqcz3YFYch7rEBa6UVdsHZeWy81tXhHo
XLjYbWiGOj1zvGK8hsCsaio2jQLnuTrx28/qCje6V2IM3hsihk/vIZKPpMABYFfN
fUp/IaVk+hIja2yy8WGsVA1MckCN6mStQo6Yrff6ALZyX/dtkZYBbCktEsfPJlPx
HdrLNtHIPLPjxwLP8kfC70KxG4D2MeZGErXUkrf5hqNybgKQ1rRUkneiKnVmx6Ma
tMFwXyiHMG0GgmGTbC6YI+d8+p2if93wyJ10wxCTBEWKSGajhyEGR0BNE7346rdy
a5N3/poXM+TInl6ZKjwIkF4w89ikNC4u99REhHjIwghXNR6cJtzgxceGun3+AQ+R
PmHXcxdS9ToV6+pqwtmbzbtgEJOt3MIx50MiOWSBnuMHENdIuSViJsbqTF8G9F/G
Ljd/Ogpubz5saHjEnNAFtlutmjhAfJqg1As+e5Hs8TYjQSwqbB6XOrmABRhTJ6oI
+s21k3Yq9NAd/Vn8DayXKgZfERta/lxh8CTRMYiI54UCBLUMXozTi+dJrTFrCJkQ
f9HwLBD7ebmTa50dF5XcM6NTjhvn2jqcWbSd9JPi3X+pU9W36yABxYAz6IGNLvHk
R+aw4UEq1jSvQxHj9aj+PJdDkbEIwQ+GNhHVc6zH8LNby9WbOrKmi2iv01b5K+J5
sigTi5JRSqgbr/HXRtO60QTCSNGcExnBev0ZJaoJgzs+AzRtDEy3s31aJ6kiP7Og
wMB7qqr8hx48BXXV9dpYBqQYI8SSfM9E91GPE6kHYzc35Zgv4EylRtBKlHMlPY/0
mxG6gYHGEBxwxSDsLg7XZlYau+AAiPkaTTq3GdtW833K7j3aX20L5XRv1ll/a8Cg
lbNQd5rNIs/sn7Ef0TRibvMrbLQtYNfJlf0tXrln7qKyDmTsYnnPfJSBQQLvh91i
k/yU9UMzfMJ6iypASz5e1nBdYsNtK2lb9JPmoKUi1KHJIxJ5GyU4SuQyhoUAkd7c
tnWgj/tL8t12q9Cr3bUiQ1zDR82QWPTfnlxxgAU0KWWT+YR3Hqj8j5dZ1WEA+4yf
GVh9yT/17RVW4OcPxI4JEHzNxpeuojQc7Uh+RVu3rMmGXYDIAdcfAfY36myf5IGt
MuA69BhA3ZliW1ECr3CnBCd5MEzPqnLkxhXEWc6+i1E8LchjrIMM9ZCz1BNj/T8X
SND8IerrRRbU5DIgZlj/7s659R3IvW3s6R0dzPLYnjyLaoRmxaog3TZjOiQ3Kvcn
hx+kpn86LWHy9i1fad12ySHCywvi+rdtlV4iwg7zk/3f9BQ1a8K+k3HmiRAil017
w8GcFK+iius05NHYCvuvMDi4vYSlgBQdnmNnEF9Pnnx4NrTBFNpHyh6yUvJUOUic
Pj78ew6jRwmrB5odk+prvN5+atE5s+etyhe3bgqbGRFtSrEKaMJwcOaIjdjYzUt4
5MhLCkl+DvPFkbUnndQzZDrh2hW5DunWpvzc//5vST07zFKvU1d3L5bM16GZpHUE
LCmS9RDfU94weZpew4PSmWp/pImYRpd94Oj2Z97MndJfxvs1AV7tqpYiG4tVp5Bv
auK2kyUlkStQuXf7/ZvxTeKeiXi6kr4NknQJMVsJZ19lY8OMBX0nbBkKw07/owo1
0utmMHeFrz0J97FxhrARbLLIc1f4fWU/8rgrPHz0/QxIMhKF5kTnk/uN0zp3Xvej
AaFp9dun2Y4YDUtOtIRD9t5ualTxHzL88mOPNPfWZgnomQg3guiccma3IXfsQX0B
Hx1690VXgmcql5B7NEgCzV3EJWRMQRDAXouq3d43yeqpMIsNVHCYUwZJdfsPFFup
uR9ZWuorm6LbBAEhL/7wIjWlqdZIDt0paU0fOEi/EYcjta/1iNpfiX04QCEr11oW
t1f2/FtNPQ9Hw3b91b/1DF7PCYIskYjUM4mxMfJWPrdgrgdghXQM9l3pNc2PPLnb
LsM5COhtAE9NfZN+UokJjiqTUuDG1ONonYgfv6VQM0sZ0wfA5U90K+ccFeXuSRFs
U2SmsT9QREo5yAnbvrJUj5ZFYI1rFDYwwjjacRXHeD10YL210kcuM9ta/Yln6q0I
Vq/NCBBcmmz3KxKaezeelwMLq69kSW0djhTjoV6tvaoCZ+GNOmr5iV01pnQpYHJO
oIC5Pz4m8DucBhMSWawNPo5qbTNg8ABV6HKJH/WuKyKW30Zs82ODkMWhYsJqUdAL
tqWHk0TihgJMaFfhZyENh0GAPxQJyOoGBncbHUtywqWchTB4r59K7KkVpg3AUIDX
EHiSm5A/pRwWnpfbkyuL31EBm9txwmFEzDmextIOZM1vo2f32RuSBsLdcfJr3Iv7
LveTpcBgfmw0Fiv04IL5ECS2ZWW5N5W7WjM2GGT6Rv0Win/q3M9OjGSDFsNEt6+9
G9c8Z2b5klmWmLAccLHxDcfG2XHGfrW7sSsuA5QZjImF85HpWilg5eu1jWb1Iuai
SgLKiHNQkmQmJbOVzubMJTGeP/TXZwAmB81yI/l1VPYqxALYyL7MWp0V2sB80BoB
chGKtlhwAQ5ICjq5Z4vNbv6YIYIBN/kwYQnINS4qEYdtna8V/UO/Phgg50CJDN4u
yxWFKDe1wOegXIjwsEtOfIK3bsgAnz/OkvzVRx6mBcPDPBD76HQ6U17wjHhY22Km
kJVJjP3Opumx7zMSm10oGtsJ1gl6JJvevBSojPOAu8lPmGGZudSHmOUnBldf70Ku
XzuDU+BgGDtqpcxiz/tqZWbJnYVS+/M0RI6FqbQaZVDsf8G3LqAwsD6n0LplBpJv
BAVlwF9jaeduVaTGus9VIjvv0BfvqeU/YP0Fx2Y/RTd5M6KdeYghGGpYt1+f4uhi
/qdw2cBMHYW0m0Cz6qSjl6yn2984MWk0p+bbWBoXwaLma5CLsRK539VzZnZCSX/G
W6DxcLumbH8ISvO4fvjUOVe6zKMkguIynZWiBjERo3RCjyCMW+5IxZV8WGRBJILt
9V7Nh38h7rJOlpEyDhCtKGiO/2nguAYmgY6oefAs4tZrKHWjgj4mpUggAzLxtH0/
Xl9sgYRlQKS6qd3NlX9frqsRjgh+m1sraXT0/q5/v+Y1KpT25Intr20d2m9zYt93
Xjm217XF/moLSg5CoiVinpJ36b3FsZD4yAJQ4nQQSEG9HpVd/Q+zG5oKc14QjT1X
wl2Dm9qj1ssLLRiw12AqA5PSyxLqRIfiOVvLciL5bR7Efbf6YB0lmi9/my5NWWwJ
nGiDfZMVigmndlQX/QSK8h9ZJJ5rHUadnIneuC2s8lVtUHQ2nf8d5bWYp8rME4+6
IVeIVK19xUqD90HFnSJh4dqOP2jYGc53lGujbo8zeV3HGSp1HCC2c8nleYEpTFMq
m+c2dMpVSrtRvlVP4LwBk8paP16yUH496wjr6n405PQgKNJybl1yE4fDBrgswiop
+C9vjnVtIE/MTi7eiei3L8YfIbYL5X2KiG+TUGvakRfppVbQZcO1okouttqHNYWE
6/hswsl8O/3YSf01csHodoik24QnV+R1Zk48Van/AS9HYjUXIiTMFPt5VQTICS5y
JT+0/jSBvkUFWT707svTRBXIAxSD1hj71tC+ArBwi5RmHMAELMFougzy+VjAj8U2
yuUI3h3akj2DQXrk0gNPHhHBg6U13MAQiYyQ42DwC+hewroPcgW9MUAee27TGB3Q
AyZml0BySJ+beQkHT9z9s9eaHZj1t1+QpPQ+lcsU0UsnlYYvmbd1ZefzP+MTbhCX
w90zrqGb1HervxTZ4OgnEpV+Aru1mvgfN/if+pJkFe54khFkVBvBwXdt5LcXvSHy
9OFgRu9Dq4vy9l9Q4/cYlKJIcQ1R+GTkAd9qzj793VCnsGqTzi01r3AERbMwBFq3
tNa3grxZDPL/5/389+h0dxNj9BGWdhAob/GtZg/E+GlMMWrImq/oL2lctxbGq2mr
5dxl/FAYgUxrK8Ndue56YMnNXMnJbfXuZfeSwqHRmiEHPjAP5tJsxCd+NKdmW9qA
zMSJK5ZMreMsHh7ekE3bU1mieVCq6lBmAxrVr6VjUwhrDD/jet1BlFdij8Ko8kAl
ZbMQWsKPKK6kPliu9DwlYs58HJy9u+LK+UCD2sDHydappuc6qhBAQvTw5UfmuCuZ
AKAce6HDhUu/wGBw/LsfQKewp9i3giXtilSqHknT36W5zTH0fUPuXaaH7BvFRcLf
eANcF6y5yr3xLZQLXQc+tkGhRxboX0uw1qgAsr8B+uMkX3qLpiZv8ivSzBxXoqbp
2BGhyJGUpOuzj8o4mxWOIpgiu/7tlVDfeSGo76DT2C+8uLICrsodv86cJjp+9ReB
WXblXw94FOy2sfZoPRLQF3EFA3ZYGBKyDtPo3Oni9DGB5hbEx+3Kmzbj3L7+8FTA
1DoJOtWfH2SWQ3jg1P5vW/AFxvOjOHw+l4Nupd4WEuEVzOxpoIIzbF0GXB9S5pOl
ozCRP+t5imIXCExEgb6mzop3qZBABFT62ZBoTi1GMVJuYML2etDTY8quuvWtitvp
Nv78Y6wzWtPrc5fofktn2H89K1yogi53PTOKAeFOo7Xs/s1C5gu4CriBXVaNNFby
UMK0y4MJ7Po6Q6lWnSm0fxIFN6LMhlZwlWGWHtaoM74jZfnrPdYVSUTP8cU5Fb8n
rHdWdhY0qkOi4Ak3lfLfb2RsKrvDjplQ50vp4Kd1D+DvDkvPsl44Me9Zh0BSjsd4
h70jNLoA6BD71EXYR6ZZsMj4BiJFHGo35d18IzPhnoIE1yNNt/XmIal3t17O8rd2
/1NLFR0INk5bswvrIMPDes3lKDEePC1N4fJdwLLpxpk0FLvzCHcYPxHs/1nOpI2M
U3Urt4MEsx10FELJ/AFmy0mbX4+7vaAbRQY8JRzuvMpUY5UR32cgN/Fkeh5EHGTT
zc3SOGQarxySdgsyX3B5auX6W+fMjlsd7WJDGT0Gs4DVwCBZYmVDCwbIYndT/CA3
y+k7bLi+kr6leQ0U7uh49FUkW5iKDqtht8eyKRyLANnW1DEjfjM84aDfZE7jvXVL
PCwLcpYc95OL4JLw5HdRfCKxg0pI6UC8fpL8/KCDsNtivt4utWUmnX5prNQWRw7i
oHmpBZJBONXt6tHZbQFXfm3lU8YXrW07iZlVL6/IuCRQMNjz/Hu7p0evd9tSdrNb
0AbaOnGfyyMTvcasbEV5v9+ibWRdSm56+hb/4YOClCI5sbpuOqbvvNUVs4Dca7wJ
iAPbnYfHzmM2Tcoo/0zwGbbpAMRRq4rsD4SIDgg0RPNjt5RTjKo6yOQpTziMqBs8
RzxctSRoG81u4/yGgKS1fMO65V3TxTI0W6u7x+lUxzSsuV6BXmUSHBPD2uQjtAER
NME1bL9LMHaBNj7c3SAKqG4ew6kVAQlbGSiXJHVUzC1+I6tkOtE5fj8TvlK0/FE4
EJdN2fnSqSlxtdiRdUGgQvbGG2vlMF7ajuztGrk64pYwbaswDrP0qu7L87IUyM6m
R5jYAvKjYquHIo3U7cuigNHRx3DV8fxhgXsWs8cVjnxBSgYbTl1mTwAA7bWAFkz1
hGcpujYPDsrBKzSRQDuf7Y/T3BXdSRq5FDVW10VpP7lnf0HAeVyI8MqgjaW3+DKL
4BQlakyeK4OAjD4hoOBuYtPlG36U9HUXkTrtSLYW+XwZhCP7rVpeoactwvCiotIl
k0cYBLyJ8P/2TMiHm9tFZsQJkmZtvTJYdDA8yF9SH/CsLfmxFS2rAtaAFSXK5S50
bn+e9lGlTBDvpbHfpAAlxmvqWZ2F7iJndn68l8EVRWBPRozXj1LajomCCRJYmy3H
QBX6M3yL+jgU98T9UuyJSeV47F+RpYRcGMm/kn2BCs90GDAWwfDI7T0GPHB6BmwL
TuEmgbel5NYRR5BeI8qNpBdkZU+2hNPC0zPH/ggnSIybaf88s0DM87Rdn7s22P0b
bA5nQw9IzgAVQKIXFUj1qm5BN+MQ1DjypTKFbfh+HoNHaCCTrw3DJeeGbvbAiLkv
t7XbxOIDAikbkaHmqoUfNlmc2y6cMMKAW+nbdwH/dgREsQJVjB7a2l4pJhfB7Al+
+fTiBRclgLlFelZHO98+2ryRV5apeRjyEmXBGzz6cT2xwcVIuTMO4vJUPW6CjUn4
rKmOuVFNero3kZPINX74Wdc6grPFxz9nnD2+vejlQ5QC+GPZ5mgDYWY2P1e2Ft5f
9OMG3KxSzC9g8hZY35ao/scaOfegR8nOLaXLpQr7e06bpkPWNa1QywEF1uU5R76B
S8Vt850ZovL34xUh0WGy66PSkiycMtttoojIGNBEUTfcwVbS/RzqMFWFBOcZlU/X
LC92JulYepUO9FphI9R0v7toJQAht5yr1VR6hFHTYkb6RREvKD3fX+rZMaT5icFR
vQwKEeZyokGmUV0prkQh/oW6CeXknpB9Yag+WowzN5CO9yIj3JoAN8rXIhRIia+5
GmM9pIFb2kuVjj6dHGppHegg8q2hxcMM+V4dlZMB06vwy6+p89wyTf0ZQoNEUzTY
iF5xF1XU0kztzhxM/0XabrJvrExp9OZcL2XArQPaw+dw79pR3xlUyxbi6KYA6ubZ
JJ7sIdn/5PPWB+ZFLZpQOphxg4GNd5ksWlFYa6U4IuIUQdeaQukuIlqnkFEdPzjh
bpL1hSMApwOxw/jxxn8YFgqiWxm7R0Cn+ou7RLIP+rQhAfBTNwwHoU+fy1xxswIs
xzXlnhdZW7DL7CbV/leFDCD/zmcyD16N6JP8YpJb5W3DI47y4FJbZLhd+68BkoQP
NT2cA/0bYD8WiSK7gAPLIiEAqejxu476RalMwqsy5sMn7FOn2BS6CVzjYCNuDmAy
wnsIhrWDssTccRJsXKLSUkpO5384WAGYDTw8hRsLWLltOyYFOJQMF6ZthbNPPUdH
NYUzx1W7s/g8ygvj9YZUa8WBl6LF/hsofNKrsSUIPtxz5fXc9/mleaVpkBwSWDZP
82F76TvTqGlKpDO6yKYKGOQZXbdOYd45M6o8tCGJepN+DmiXHXmPumuVGLZkbYgz
Mll3wtm5IolkzP2zWiDGpzS5RI0AsH2hkc9T4bNoZGv+rEXWIVAICKRn2rHu2EpY
HTkh5z2Qiy8XzDTPW9+2TK1gmce1jLldowZEfY5BfEMQcg/hx2pfKJK34Utdofkp
GzwDAwCSzr28lruBCbIikC7OernQuWUzNp99gnOSh+9o2i58uzwwcUnAXOp16x1r
s7sR1sWX6UO8PlBvS56CzoQOFNO1jdK+H4OyrUXUIu0B0WWgb9xS/12JKeekpDCQ
ZhiFJmGi13n5SeLzc+zIGprOcnNUiKrop5kJnfcCSjVkpgn1bKlymiTR2oXSmB+h
upWp/O+IGEpXuLRBxRxS3GEBKn2wYALqNq1hhE5q6ZnvkDjDnDEhIygkUDyd5Sfl
S+/bIThu9hFL5ZG/drlw1e6l9AHM2c0quqerDSo0IViETn61XOZdLmVScHH/OW9C
DiPxMjaN7JXIAA/gusOqselevrMG6f8E9XvzTSUqoUrFgudSsRKmXnhwGyB/7nfK
kcvL1pqxeM7rfWy9e4WbvnqV2J6ev+TrcWhE4RkzvG+fuxM0ruZdwGbn/6dDbwnG
y3xUt5dLwRJMwTJYkEt16RWVHb0Cs4lLEbIOvVu7/2ER4ZLEG0jFXQR/ZBb/Ji1K
qoW29QEqMdVkSWR4ZcruE+6EbMP87MGrUnX9xEHZ4JuhABX53zcFtsSROk6lh3/K
Nka9W0et9ybit2Rp4/6n53OKMXtK7ov69PLoeUQDNWpHDD/T/jhRWmFDg+1Odovu
IVJwXUeDdkW8FYMchFmT0G557qw+iABHO8QLXrXdDEWghZvFfKmP8IgAqdw6rZqW
NJJDF9UVqfWykxAG/wAEMlkDc8Y9wF8nlTwgCNvdiSzy02+XDoJu15UtSByT1EQR
uQgw58N4DU6XIMF41gG/6Py7M22s5aDdLT69NNobp6ckt0Qr48RTYH8F0wW3FMxm
ASp/2Nkcltcw2b5NYtjm/8dY++aWlvKWg3P5uMAO8AdgcYRGNpecnXkgAQJTDbdo
zPoN6d3YLEsOdtwt8uu/Zqp6+ntdv1VvHL2RkjmVVhOZEhNfkOHosvXGAbT3S1mh
7QvCbhZ6N+RLebDYyAg/ZbkmkNGjLUJ9RHZCnexMRsy3RGKqzI6CGyVhFoURXjGj
8KgLV7zsKpOiHPQTE3LHfIV9lIr/dhYNq/OBD3P/1sZFdXFs/cWPNPPcoH78Qgx0
pMOuVfGg0VaPrZZyBnB6Vy+ANNeaGvsUdo6/w1qN96YDd8IeisQ/TGrcgTmivG0Z
18wrbRuD5FdMi/6E82BUK4rrK5/oVzKudHtE6pdP5ueD//S1docHEwsn7IX8rhps
VtRv6TpLOaWWmmPrikaWlsGSGEy9r91MFe8S4ZWsuqGqmiGSv33YFClKkcFrU3e6
7CYa7/NZc1iyqWrNvQL90kLmLZq2JemOJo7w2mcL/5ARxWenuQhMZN0j8806x9he
LW2Y+yUBnj1NYoa948xqFA6h4NNSKe/F2e8wd0j+PW5v2ewaIyIHKwnnl56AzUl+
BV2Mto6XiWaLDRsOWFDO3XT89wxavuSAhDY6W3H8LdxoZYlbWVuKaRv69G5r0B3O
tFZ4NWWZy2riJZrDKmPNGpxNoNDYrdCB2zTVob4OfOULS5aFhxPZQiRFnK4tZkOi
isCK5H7JtoI3L8jrkngqSpKcfXArF/EYMjm9kRnRwxqlq5Fd9clxPszaSnWf5SKa
7to4601pBlFjq3CuIKu2HX1edlROQspj9F6p4+kn6VcrMi3aP4HATaHboweeyLEj
udW4kjGtb/RhYLx+mua/U2KEJN5vf3jveYSIzkM9o5M/h0Ozb9g4iEXgoST3mrOj
KzMbyUjb+2aNXSnAfZDieqiMFjYn0VGCDd6przCgiWzFQEWB9rGz8Db63fSEY2Ek
uNa5+zV5pOrVkE9BVw8FWbkcsFcArzIo3ZbEwHWGkWsgWCPR/DuwgYT3QuzqTEgy
wHfE5bf2k9R0VFanGYLRZxcWcIbSP016RyV48MgArYGT6FAoY6fRXfSXOZdgzDqv
WSLaucWJvytYh0fSsGx9CRHmpeLaDQlbkK6PmuhZWVwSjV9VC39SDPOvGg+jRFjt
h3msF6qDiBREYLhC1CXwYww7IreDGv3EkkzMKLpOvnCbFwTR/yxb54YPedy0vYbz
MRlnH6Egat+DPqVDOESDBfgQZCe/vKHXuYHJ74Je6MNrasvHr4d1DB3WL8imeNb0
arpDzhiFhCyg9BLTVA0lcFBQSKgHjTVhox/7QU5IRvNwbAM3KyI4+uo5M8TzHvFA
6P4WbY6ezXQX+fTdiIR9sQmzuCKxEkwbeyI8b0F4tGa2PMeOYKWzGOamYgDdCmhG
rUEBgduyzwHXJTyQgodUyz8kHMQKcyIEOcFXP8QUSnlXBuwMJn/ZGXBNso4jvCXf
0O8rHNQy48r0NgoGIApYhmmFXo8JNbfbhIU3BuF+/HVszLC2OKzYQEDfLxTtZM7h
4fytQxWqIerCHAFWBsHaByu429x7CNKRvGzba361VVvJggn/W09Uc1X3QXU90ty8
fNslc+1H2PxqEDkaRoKdXLUW1+zKDGJ5miBLbH/eh5YY/d8OIFuvckEvfG2rk8vK
ninnfCokqGP4XsRDlO88POH9LL84wLWayEEMRsImg8DyTKDlYmyCq995uEpPokky
YnVYIN8bw+ckwXEWbL6gmc34BAn7mgBap9oo736y/js2vmL/W8IzInDqxS5qc/o6
iW7Ol+pxftD5ROVpCDlxWACAoHinpqZzQ4TuBRvgQpLm0B7T6qthVXXEZjePH5uw
xJ+4cDTnkAnruSpWR+HN0/4DC9whKYlB85irll7s2ZKUiKjV06isTvyOwgQe6NLm
HiIFeTsRGVs9/umEd1Ag2xE4D/+qVOVc60G0I7uAAk9Q8rVa9jUJX/iMXyN7fP7o
cMVJ3wPfEqpPBpUG4EQWj3tfUPMXBULlPyxM7IW9Tjn15YZB0vs+0BJElV2/EHwj
CpX6+RTGDKVIWFK0xGksQNgX+MlDUSo0ekS2/HNgnQS9SKfGCh2ZaxjPHNHfoFGC
rfv4E/HeGZS9VPHoEhdUTeUi8NLVmYq7V2hLQtK8TklOq7hNblSsvq//quSXyNkD
UyKHh3StOZDvYcFF7tixe3YbKXoi24lkYvs00rly47puV3QyxKSCT8pJ8c4lat4I
NlFiTLha8VNnIn7n8Y4xqnTqMhqmEw2oUbe6PF3jZt/R5w/+BSJB0tasp73mRi/7
JZS9TKWuaCL2II1rjEzWIISsDMMkgzdgNENaPh9d8DgKe/ZYfOt8wxPZElhx5BxQ
AoJn50KWcdEqAS7k3gR7tYMjngtqqKF9PrIAghLGt8zQtzkqQJQMhpd+0wLpXTqi
qFaz83RrQenK3ImArmq5mk9m7OyR4HfMQ8Fdav1rcFE8fsfBY1RK9rJrQoaYsq63
ZlJ6uPEWFBWUA+T3D9nGwOHoTv4SCFwzD8DdcmwC+cYP07aqcBCE5bEmu9SYk3Nc
TYGBTr17SGrTg4jBe/wqkgsc3kwKgRCwUR6m0+qYfqMCLF00Td0lVT6KULV7PDQm
WpcvR+oYMeP50lEyRkyLp8Ui85bG12S4Htpvmk1XmDcdiGBe4B4Gg8JDu0gTfab4
l7pawr7rCHl9o91HWW47FTBrZwHhyLIZfZLqmjpgZzLzMPFrgbFIVCWsF4Wzu1Xu
Intyn6qh/veutb3EStCu2+oWRuG4/AXtQ1AnRARvWa0KLkhs+YQOpUlEl+NrU/qB
2r9fWL8/UC0MYXxYwL6/IyjpXOBRBTf8op2b3APFxdNjzmVcDsZzdx1lPDm952cd
2mcXp/fLxvRm2GjQBRHTGLMxOWrxxOnYBVRLEvmK8U3etZNr4QhPCdAdNSY05utr
aH66jIfqgYthe1Mc58XSx83X0EddoGRzdGP/wcMjmCfISqSPINMJtMoV/1IRdQBb
Z+7KDj50iSFV2ryYQe9uboPvlfmlOPumWA/Pp2/jTBnFRxhtnClvy7E6cUJtmU36
06zKF+cMyt8VuOat6gRGxnyYo0DJysSG+ElEyHql4XRFiXEd6rJje1ej/KKpHfTR
878EQAmcvmNV0fK1mx0spXNBNaukRrHogziGzEL4N5bpo+wuq+He/LIwY96/jGaM
5mt6TZueyIrtfSKFchZ1nmcw95ROxT07tAst4l1Q5qLMc1LZHie1kxk7tnBN0qB7
TvnPVOgIiSOwG3nnymolX4FwUSsB97MTxFKvGxExdzduqjmmsfWlKlzSC0KVeXAv
A3Tiqruu5Ebm9z3W1UKF5dr7fvf4MjQ3Ot8tWj5i7CkfliA7L4gM/jYCt2h0aVcS
TIBFWRuI/cxEIRS7zxHkEy3j8RdokFQAAZBgOt/z1QEWUqpTEuIR3YnL8QN5/4Qy
wJb8HkAiJ9P6GSEo3MDpH+yknNGlLAcIbnVKN1XtJ/4B0mWvSIi0OS16DXn70LMf
+mnP2jRhGsGWzHNCud8IwWnkCMvQDM53/URnXN2GukZRZlWm3i15zKpO3l4y9huz
M1SIXU5LoJCD73LDQ8EN8gF1OhnXkNV9wapSTrw1wQq2hYlcjjssnJEFEYMkBczV
pNTdDXAkg+DkD5lZ7De0F+Ntyo7lZpheKwjqS8DVcWT5h4rCvbNJpjWHI62lubPi
evBnyqWmjj3peH1novQwEYDMqqiJ2YNF6i0st0ZBtIfvlQ/kPP26hkm6nFBdxtqZ
azvCSbaHzuFeivjHxit/Dx2s68hEYKpHanBysQzQiwGkH2E/+Z4MsQ7Bo+kRKl+T
QWOt1t7qZAzEu5Y4g0mCWU50TAKPH+mdBjpgHEqiH7JLavWRohHwjlvi6hibxCip
jItNzTYzIU3Wta2VXLcMq5c2HVnkL8bRL6uLtWRnhdze40D31LHPYSfrE/dS7xHe
CL4qXOuw2zDc7jjtteBEU4L2Sm52qkM06YEDyAXCmiVJkRhxRMe097Us8pMlCD6y
SGOi2ngl0l0SsagFISn53iwlSE8KifR6OT0/jhuKTZded1mIPP5lUsK1cAez8qgN
bbyCt0g5CC0aW+KtdtMfpiFZqFiOD/nvplCVkgiSan71mL238fSf1vArf5drj4rA
PydX1vVowLbmkrlTdLJq8Xih3DJdCMFNJ3B4ExNcZbpH6hWZbuPFR7t5yOGWwgXM
9+dsQ6vTDUCD3n3+5cIOdJsuvjk8D0NDLVwc9nzqNzCk/2sqyShYQAfW6xmBUZqU
fnY2Zstsog05cTgBL0mYWl409ss1Lo7aW8+6itdiko1rzhet2pjfAP3y5ifeQJoP
FQRKQvaAGX/2iqXcWiW/1BgYDPN1uOfBQFbnv0mm8uJnVHf4mt5MBTtpEfqK0w07
eYMpK23ddvKz8T6D7Ns0GbJ2mxxyT//XFn8Om1WTcwlx+JHJiWlC8SB+JvjdmNlV
BITiWjEETCFElVa2uZJszZZBt9A2W4KSR241VRP0q4pLyea/3XRQtVmDajnnkcZi
BX0CcZCdAkT6bsrvx+h2B3DpvCxhF26RIg0o6VhYzLvB0e/GPO0RFP6TNNxGKywS
ImIYCdl5wh1Fs7rStuBzA0NgZeqwKsqTgefN1/HAILf6kZkFDsCrGJ2AmmuEFuH9
D07R3rn5xcoq2tPLCdpypbWVxEgpkIFwFaGuVDlnFMYLJJ55kOxrwg5JriYcFD3K
d+TUQzJHWKeO6zZogk98XpwwkcU66iVUcRaHPsuLz0XDT5EqzZMuZwByazy1Kg9t
S7VXjSRUYZ8R2Sei0z1ka9DfwN6lBbIsXir/tvC4XZzphkSK8JqUfpOIrnykzI1p
dbaUazeAZnchj5jpoddMNAQaf0M6VSXMgXpFam5O9nettB3Gbcco8XKJgDObX1On
kx1uWh2r9XIuYCPtxo6wW3ytdqVE++lqXR8rXGWbtRrXnpG6H41tiJdHJ8MIwUDa
oeT5tDyKO+kTidPsYFJl7hC//th41Lrpi1cMHM+Mb6SOIFtexEyOfIjYrCkg7yJD
haFz9U4dHgOKce27G2laPPRY2Jqq11HNWXMNaJ6H7Q29rfOvmrJU0grGhVTvUk9P
vytLxtMg2XxS1ooxbscDOCHYIY6zpbMKjqAHP2BVyxehaoBotaoqqcXe8Y1vf6LI
adMJbMw6ewWZv+w4mh3Yq+6KDTTyME0l8HtXZ0iUlTUYRrZH/YDf6klMY0iextSd
H2KWvdvlsup2VP3AhSWiDku4b1lVxpspJBGkVfp0VdVA0l797GmSFo9PAYHrEGCm
dos0vCcv+scRP8x5WHkggTarZeAFAZs3EZcrnVPq6hXeWgIKtRoenw45l7xz2sOO
Ln8c/mIJWRttg6YtRlwUXxaJlPTszlxx8mWZGZveM3qNim6iD3JRkgBgOAqDpnqc
lMbWEvdOx6pNsOLC76mFFwBHfW8fXcIcbnExJbqgkZZcoZnYfSySCSErNJNymtV/
cnRLqpXwIfJohye1bdKOXqYQnOvOTmKe9OvELeqHqqPWi94M7+k79uP6H1G+c8Of
WKBps/KaVj83Kwd5obYsq2fLRsfUOHrc4UBaRT+cOT43jv+AWuxaHsrFVWPfZPOE
ZG6Fwc9CpmgwsnyT259rhy3Ku9cku/MYT2kA+FTU2oCIOmSbnmWefKliEsn0C3IB
IH7hjqAMJJJimeO6hV1KQSQvLXSBUGJeohp2KgB/AZ3ZkIh7mKiXwahR2TfdQHPL
nk/i3+VOfuf6V3Ls3fynD5wpzUXyo0O9Lli7rTAPleYJLUVNfuwvdqECUXBCtQqi
XEwI8vWOrwEVJnMD8BsCMmc9o2TVXFFt9c+z7/cOzbHbgZpuYH3ZbD4OYz3ehXHS
v/I96uUl15hAXRCkj2deW9czIqDvnDAY5nvspkz4+q02dD/JHnIDFidyPDeizDiy
yRfARrSAI7XhcRKOZiiowqo8cT4CJkjZDEBg8ugdvu7vMIMZi0Hc8FM/tg7ULOGI
iiLJWHAd8C4jfHNthGK4GiAw4Koc2dzoWsU171O419EYamibbbzetBYJnT7MWxVE
WLS84VcwS0V/HHN3EXYEeg648J/eb45ShOqRVCFYykRhs/K3PqeojrgHZwj1NB4v
RZPxINIFJoAnp6JIDomwjJnW1NDaIV68Jsd8ImD2GWjugxO4t9D6oPLbIIqAGUKv
8tYUPVyI7Cz/AoJAgQMpTkY7+Gn7zGZ7UKyyeK2xgI9KiX5LJcpGovw7GCqhOExc
xRyEwkjXFuqfZ2800s8tTcQJvVJo8A8n6EQ4OMOgP3MLM2nYybYacjeI+HIe9n9w
x0X8UP4kBVfYZIIkjcfBqN9f+HiqIp4kBkdHj5Uq0krfmDe2F21cq7+cx81SBmO8
k+6OSG3MeFjJM0j1wNXRVC+jt0OctXk03WW0S8NdJ/a8JtB+1VHhtkhL6gNrIfcD
MnZbSDPjCEKPF7rA93F3l6LAv3Ll2mkJKJdXxsiYtRX0As96hTAi/KY4+IXDJ1Gi
6zAs2e5LNbe+TvLo1agA0gAxZI1JhXOt+WrDwUl01QRSfKSu2maYcqhBXKhK/fty
VkjVO4VmMyk1TX6DeUhNHmNmvQzGC9bQRbS9QYp8ZUqSZWmMuHicUErfzBVNbp+n
wmRn7XcrpgUcrgKKaBVVPI3gc6J/drMzpRzyKMld37t/pKYzc88CL8QwDA95a8v6
NRWFh4xEPLexTrX3pX47vOJyG3eSIEyE+cPtlWY4/FF/z7S8dVu2RprGx7Mfb+P5
Yt+12WjWjA34hfxAZX5QSmTE6TSuUNKI4BMOjzTNT280ZFyTLHD4vMYb6B4sXAnq
VWUCnRiILsE73I/TAErBB1k0HmpWgFt70jK/cWsNabjytmL/Dqgd8fCfc6LVfQQX
8ZWIdbzNXjeIGBAMI0Q11kdMOl46QO48NaVYeYkT4ec/UNrTXuJLl4gFupah9nlH
iUphSUGeFOKEsB8Q6YzHPxfHIp2Q0utCcvl18eu+zxtMBikqVdHVVx0jRIsIXvD6
YFvHVRqbTDEXZf4E/tZeAAyD03yhE9Drn1G/OfMGe/ISJ6D7itUBu+Ixe/oH9yWB
9h4/CCinVmsEFZmFs+r4JmMzCrTo6dcos+pWOXjTu/Y1Hw+cR6nkMwz0AHogE8Dj
aZWVNvL2Jlh+CPicMXSh9O3GTDS0VwalYaQVE5j7b1H0BNHJr6ltQzOu+VTAobbE
dbN961ZDJj7aA5Y6BuZsKTKP4pc8m4Wv8HoXrfz1rW2il+DCYQauqozAnAKxFdlT
QGfqpe5rnSso74ZxRlQpyfiU2dECMUGxG3OlyxR5z3czeA9yxMKsVEYEWVf74t3J
k07lkOkbbGDOS+4YQJLflwTOMVwHIwML69/zsPSd6eNRY3gUNjx7jI2UPvHngI2V
15siUwbFDmEQ/q5UDdu8utnOUHn73Tq2v5nkkCj7SIprLxz3C0Z0FdQ3Fk5lkIsD
RbfdLqazdvifT8kxA4hb7C5meVnizxl2D5husOmK7cTihXXSes3Had4Sxg5EKs47
TemmiVOsVjUnH8kEIKM/LKYgaodKY8BjaCTVXs3P/L6Tzdc7EwpOK4p8+le5GVOA
y0tKLyk9uXVfEQuX1oji3AKYVp1v14c8BK1DVqaX/vl5g+agPyJz8HpVC60QyJzJ
BNBRtEVzAPlnNMvwCu5Bn9gMhlVzELHM1RTpbunOLk2g3NODrFlIFGgrGwbw31Yu
fg8G6hCXnFa8q5YdD+sFh4tTlWUkw9HtMPIi6uBwkgdC0rwOzHmnIwvrd90loPVA
DyUlEOUXSklTYMOKHmteJFb0LFmAAXF+T6a0TtTqSB7M8WHF1iqgGo7mck6UtdqQ
j80MMTuAFQRrmtktaTG/Aavfh09CXbJlMV7RqHXNGOt+gCxpKuJ77TCyfYgAEYSz
5hOavMVaGhg09uEIOm7I0VooEN189gNs+TJ5owa9N/O+PWW0XXEl32eGIjx99xXV
jAaD8Q8HRH8QnT8rq4MDZPptCoPVwKnzEkvh8i9ZaKSc0Uti6ISGq1s5SDSwgctw
KzT88ZYuyHbCvV9grV+j9BQHG3T5BiqkBdB0/mNmxfB3fzk4c+hbyNK6HwTNApU0
fd2SwzeekEq/aQMuZHi762w0hAxTAYKeQYxUUjzvmN8bRx7x1o6tv7Di5/KJE/H7
JSDKY5oo4UvaMA/O9ggNj0SJQvjDP9l4paET4m+yAb7f2dQUFCPuketmQ+f9d7Ed
aHiCx8TvZPHetDuYIf0XcOMln0l8ugCDzjU6Q2hq9F0PgPlPqIsbFzdHE/HjdOMZ
/6mcI4gZ1Vs29SOfRoHVr/04H+NwLqFzua1jd6T53ViV/iTylkSijquZPdnxwDSE
YkblL40hKNnz5aw3rxyeQ1LOXVQ+koIIAWdDftLIl1E9N2NVFmZXjtCDKPpclRwR
sxOmQC4rGECytUFeNyLoAljaTiD6JOdYoeL8nKk9N2C4cpGsbXscCwJTs2Njlm6H
zpE6cd9orRtSnOPsP1uQ5lUyZAxQw0QiHSHRjNJHaLCq4kg8WJnQtZAGEZM8C59f
XlwVrOJnVJJ6wbpnDk8vCiz8H2whHq5mks83yp+7+qjHM9vU3yiPOSIQ3QIbAJ4Z
J66LQECywwn7vB9cISjuvhmjVSn34WnKy2sK7h+LNvkvvX9PHXMG8IaKEW+7DhmB
7jfwT2H330BpszhHHZfXKxe1oXs4YgaaG3jYGbgVZlR9Tc6vpUDYPp9UwVftPuBI
mdLxvMF5OqEAXvmQ6AwayLCO50QkSDRn24ydvEh14Yi0Wrwawo22NmK+8pnXHt2o
0JtCAKvZZkqzwpbPyVqaRhoR6l5xgdSrm8q4T0B/yEERlU0dYjtzf/wvah+qxKZv
qXlPGCb4v9Y/JlSwp/yB8YL9lc96EdFrI43o0YrfNKLiZg5iN4ACSrgVzo3s8v17
p0qy/O5wvn612MKEC8TdzuyobCR2PFOEew5iDE4q6RgcRwZdGsvFPWKCFmlO1UY5
X729p7VCeIGbLKKmSiLK2qIjzrtA0PeTFAdt2X5OLdz2BhOXEHRnRsiOzxxuTFIS
ydQDyBaoMDW9WeWEPznWHHjpuM5UGGOvc8VimDUM4Rb9NwTze1qsePthChOYWttc
Y6lQ0WhG84JshJT0c7vLM72N9yr8d25JRsRSUKDCZFT5MMT6ggnXHTywDwrHoHWr
D6DTRi66tRfX2MQAkTyVD5RyBtVjGDb98kevZkJb6FFyOIjr1j13JxVzIujYH8NG
mnA+XZRksC/FyJ9hzCWUGQLS65hOhLi6u0TiTRW3JjtsTOZg8GRV9ZuwrISnkgFY
fZRUA7Oi0kO0pzq+dyxNKYLFactD2V7Q6JmYVMr04qMTtPM6aBUPrCeRad/NXP2M
Vq2LMdAtmqGrKCTyc+zqkb2wmbWMhRpHcu/VSOZB8gU5oaXSgSy8kw6M5y/tboxJ
K+VLNxcJgJb1O9yYCE38Id3I9XKiIGXx2k7ifwlWfcw8/NWoUxfmpU7HTiPgB+eY
6w5Hvok2RoqBGfLol5tm0TJ8rhyelikEjMEhBmkPE6TasDeGMPsgX4YrLGR1Xy2t
IaswB925mIMTPHo8Vl/fBDOufkHhP0x8tvZYuE6t4qVSbqRwpByBiqfbCx3LodWo
jbPDDzkj8yGPr6UEcW/W2Rw0tLHcnK0zrphg7FPxBAC/nkqb4zHFTCFgt266l2K/
8dtFqKm1Ezt/+tw5PUjFRDudbVlPHQgKDLLASy3P3yR5oaay6/UUnsmtpsRTmN0g
9HEUIa2vNbxtACvBcO17pAMFzhsCCUBfi7RljoDSSXBOZfhRqR9LLV25tmHedGAO
35rNhbsqQjzMojepg+Iy8auZhmCGmlRwYBtxfPz5YW7ebBXW9wGw6N1trqNS+Or3
iwhDUlDG2/px3Qu81YC0p/rsUIRV0/hlT7zZuPq8lGAXFv+Bj7h3vyZP9fwp5I5H
/hiVs57teiv2+xfCjVSFxPrj/HG6soxC4/HOZNI6g8Le/HMvd9rePf2UAZkO+C4l
xsHl8Fx0Me+0bxDePaqHatNmBYMvDPsvxaRiYCfdrHV7WB5fzy1iLWwU+RfmGU7q
zT6E7pt3c9dEQDk/+DlTheB8M89qGuNq8UXwJ+xNKr7g8aIeDysDZZarcu2eht/y
zUACjwGE5RDMy0tc7dM++GVhQ/PQwxnEMh1CeKhF2MoSKAQfH1gaZAAOpvYbZBKE
72CyOPQlvlNhoN7GsaHdauqrfAK+tPaUzFNt7djgsx8qlQObRr/zVmAeM4pUd+Oc
RLtYjE+GXxep0wFL+vPbdU/B4/pRQv4fQNJFKjsE80p72gnUOK4fB6HdeOpaYkZz
/3ZnbEnvv+71KaEfRbkqtYjK9kEbhZRRjYqaup4w3jHOot3TyjC7LWas6yDhwcpC
FkLv5yFZoHqqRaRb7kKUd02TmtLcYK1neGAEIldf+BkV7I1sRCKGSiQDErOvU3dl
h+OnNjRo28EDTiuZ607U7U3Mt1tFkP2VOd1FBXq6lr6o76Q/D0nS4yUamvNJR2T+
PHwB3424xWOnlNgy07yYMe46D+oi7OqjfJFuSFM4kjOVxb9TIpKBIOxpohDzZld0
BRKSBWaxhmSks3s4Ln8pthP+YjXdJ/w5TH1siSE8HaqZO1FfycyQkBD4WAAjoPVs
41OIuy/8QyXqWXeNCUCk8cwgSLzUPyOTbw5zroBVJ7t8Y+nHLb9icJPiE7U62B9m
J2K+tvDJyCEbL3zna0WcJGl0gUYsW4f4vTnLlateLsGUYXpALmwiagphYqUSYvJY
AtCFlQIeuuO5GD7/lLCC3zd16iqJoRsuUeQJqo3jonna52yPeLVpD/jKIFvaFWhw
CYGdpnOcWvepWDj2sV6JKMF92+sbxpTLl/Jb8xdtjoWGqBegQU3BMhqiVQIQ9M/S
yZJbEjMIY70jY0cRnE8zVJg/hIJe+0RXmyBa9zI12kcxkGHkx8PGwx0hlY/AtOpQ
7OMypmEkBNzoqkXE2uB+YBODIuPtM6o7ZvQ8RMvpypCsKU8ZV0bAYKmjE1/P8iVM
FmFffU1vxcxxT3JqtFTEcPe3W5QRy1EMnyEAVtO2JgOJYnkEXVi0MKLgIrF9gCJ5
GIRfvh5eucpmpWLxUOUWj4shF1POjfMO3WE8CQa+QLQ4rLyodSQDe2dlEKEvbG5l
1FYFf3LuaNQQcX+aScDAoWoX47dnp8adjZg9VrQMDb6MEQ4oSpKOM6wKX26hLBAE
wNkFfaxf5snPdVqgvQ0a9cdJy523lpCo5oUi/iVG5cl9fWW/QswSBFV3ePmgP5G/
UXsBylLn2GwEmsHb4FaL/2EYxZVDZVZGM0WtEiNQQ7ZtJOoOeG6H25SmDN6cehls
wb1oYwOMuyBI04m0c1ruJrhh0xRt46IcyyXY+6LUkDTrX4SvbSyZ2Qy41Bv/XYz6
5gKgXSIQpkYmEzjpmQ/Yeofbr6z41U7HQHAUmjo6iHMnU00EdtCM6XNos9UXWT8+
Iq3Ol7AT2cSD6O8VKKMgmigG3azm/7rnm4w3TQA1/GELCDgG5EM0OUWl6PLHC2Op
FRFaGzoZ3QvUIggsXPq76JU2R9s3VgQjaddwYSRsZGcMq/zBs2PDzcdUyt67huER
7Mp+fh+4lKZIDEoXKFn1SQ5l1oZo2OEf/9XnA9oDvuWa3LGTi0wiZYkH0lR9E6lN
5UNNaDjZwxU+kJVViqMm2xxkiL8cZqeOjO64oGRhTDQHxwb5pcMNxayRRCr/1FWb
mmiDixnzjafLJRBH9OSdsRFLjsoTmptHwLNRA/bY/2aCzZnORO6m+aAfkk4DeS9F
pFgq6hqB7CE1hr8QVWCXxpo2+r6ja1+UMo5niltFM0ryOyNC/SsKwF5SB5po/CGv
R+GUqBEGGf1BnhekZnLkdbr3FBL7el9REKr0jCHyz6qaRwEoTTZV9GJPN96jsJHU
WUHj+v4upNiXqUQuQXOHYdj/8gk5ug+Br60iSY6cHVIbrNzJYxrMonLl2DLqaTjX
YDjiSG8okkgrmeBF68iBpnRZVr17zUZKkaARWAu7RFKOCR4ZdxknV6VgVlgZe41f
IqpnpQO9v9t0v+Fb8Bf6yPgRG3EpATJsdIhe2QL90dJoy4QJkRWVSYb2IaL9AjfO
+3uqExN0k4p4PnzY+IyUyTXFup3w17VS4Pr7KCEB47/zro6rXE4VCksONZtlXzHm
qQUKnLbEr4/vxHukTN1/k6YgVOPrJ0Vy3ZElaBUJaEZ+V0Kutm3UBUN7phwtULUd
MsQAAqO7b5J3XMA6kfegB+ldEAcXirsXO7eEESGp3Ja62It4E/kEkTdRQ65qJ3T6
i/F6riPILn9FqIj02P4ilQD/7wsbEubr2MKSHFZqtFEN9URPvoQf1wb0sZPPTlXw
v2oOPlMC/jb4Ymr22qfnRh02fjfL7be4l4Rff0XwlaRAkSJxDsMZvzWc/T112lpt
bLPb8SAz+yJhrf4IxYJWpGyI2Aj8pjvEp9fSYUR0LMszMrSowLIFsfNesHnKpy3F
16GtQy3xoQyINLs5ec2fHPq6vbK7VjthocOlDEfwYqK0uPLCx6EMXaxPFW4zp93b
HHzjk8IwqRaz5TliT9IpVjOA4bc764nR5O/sE90oJgCBpEcH/DOUmy3Yg/hgSmav
HWbun9ipYFK8iMKMt/c63lXdzFi3mY1eXtalMJQ06NbcQQwTaab0EfEIDYnV4h8H
3xP4dNoU+M6QFVJZMsr8/2OUR0as2USCxcDhUoWZzho6RilkorKIy1rnIbbm+QqV
Ds37q13ASXUw9zODJrvzuAuBZYvtL9NNrurfi1l3yu95ApEXRaQXaGCAl+nziuSA
NyaEQK0jS5H+IhIsJt1EX7DpLduHqa2iKJwYUxDuFxbCh/9Zi3T69FoPcgS5OrUJ
OpfE5e2gPNOw6jni+uL0z28eQ80M3qwZVEfn3G5P63R2T5uJAh995dGNNVWZDh5V
U4AFPYZdmiTT0AeRYvvL+zeJWPBrICq43xxx8IyoKx7casvd0uiUk0IQDAHA79+L
+rVH1HiALJszCMS/mLf+iyROb27GhtmWrmtlVFw92v8wM4Z3i55Py1WJFRfM31mO
0f5j3c3VjFY8kM16cn6jzLAuN8fyGDX5hIrgRtSeMRghSTzFqIC+jqchHmcYVv/9
z5hlP5kjf95qV8OGK9whqo7qeK07D69+aOeiDMlJ9W/szeYpjIDnQjoP8DB4NM7i
do9q9bAuxs/N8ME9r3CXyD8qh3SOw5kT+4siw85MGFgH3YIhuZTPhxuy/ALmY00I
ylfMdIDOUQCiIYbjnojf0YpVb9u3GwSsTy7LosDWds9RCqPQRHr3tEr/tbLtDCzj
l+nPbjCzZj3l4bSDoF7+cWlzJso+3uJKBFIl9TdDk102aBX1d+JRC3YjFalvdVdz
im+4O174fX0J8CqE9mX/WULaWIiARIrC8iqkAr5QGTbzOq3w3hRgyt6qCkB3zggE
1zLRTXLVEqRQJjhtGzBflZzD6TTYeNWOeKevcmLSsRfqT6sERR+TgB3W3P2h6JCs
0e7Kc9HrAvYGTNnw6zI1I10cZfneX7LEEuxMDm3AULMb/GN/olVe63udSUyg36zA
bX2q7pvb8Q2yOBJ+tgWshJJUHnlLAI+uGyOzXAAM+CIY1m7TWgxK/vd4nN3/f1Ay
/ZIdzp6s3I25M21TamhOvSDq/o8IM0DqiZb1UbKohFBMocCP21qPI9SIuHAVoNym
GRM1utyiuo/t7oLPloh9StCGONwMkK7laYF8SQtV4n4BsHmdmz4b3gJVQoAbPyWI
XxEFFXRD9pV2xJEsuUeKcFsXt9eMLDTU9au6z6LllYSKiafprShptY8HIUdPTJ2R
CYZxJkdP9tMTOLShrYHp4zKt9zyWoovoCIYUUM5DB/FjREQp+dp4T0NmGX088wYq
H0QaVaIfkUJ94Ue6vw/RGMgyCkMkx+TH3K5TQcQ6oGY9IMbkw7JDTA4CCvD7npef
mLtsdEsRZDsI091Vddy9p42fzsxDsRBzACQ6/WAyPSyWEk3nJSHwqXqQokO9wV2o
bpvSeu9C/vfDPIzBgAvRyGogO88atpk/dhytalcv8E3WqyDX3yfB0Ly88Xh+E5zH
WJHy413tfd1hBaLserhtwOhuAq7bbIwTs8TpYgOK9U7Q7hnlF6aRegPDuMm1zfkI
jcUouS7I6NTgYmcgkdZlo1eu4kMiFQ94aMyDo7nGbzSKHEaIzkh2NSzjoqjxkNDi
wM/fI3d2I6LY3P4EG43S1WTjvtrR5JO/RzMt47e7FynX9eu6FA8G9S82MoBDW1FC
/zNYE7RpG1UU8SFgThJu1fJn9QOkRrsJNZvsdRrREHvSfFrHLn6oTbFa9ioUipkA
iXu2o6KgZpuVYOCzZPcMyOJNcOZP0qc8Xo3H4cmIL//rBQisfmEVfU+mdn1vjei3
UOFDtqlXg0yFmCsOs8NkvKJSKo6eZ8otkTVSofK8+8Il5sje1Zg98VmmoxeLF8e1
aR8gY2IaufDz2XhlLYW48TxhFlDczvzLI3MvlPQnH9gR2h4Cxz4Y/MPLKypJrnj2
SMeCKCzqlbIbZ1BZMADJT9rrTF0DaENh0vCxvVPdEOFkyzjgL4P3p5TZ+zDvn09O
AluA6rgIFVxS6I2TsocDvRnJaBo2BISQ+ULCCHDeXQ7lTAGDTPS/1l7OFTE3ZwjW
9h5IhLEpYiE1XXf3aQzb5rmk1vceNEoUG2FRcmsbjD2LKoajozWUaSy1+RjM5b4/
4TT6S2T/yCKPNuuhS+w9qMscru7w0BLnPO5C9QmHAiPhuccJpxNWJgJbeqE9KvHS
bI6eZOXaDkXvpdETcctSywXC+JmkrpOx7YPFmxiNR7/mPew6YhP369zdOi4wWGFy
0dnHQDq1CUaDm/lWat9IHZEZ1iD6Xmp5xGyooRapRfVYlfYh7g2y06e61bcnyYa/
TCYoQmBvBSeQxS3gymrpPVXEIr81dQZr7vtxOiH11VvUgqa5YegnbBK3d1ejT1x1
CGbkt58CgCpAIvAym55acWP+aHqh441OoD6syGbBYwUMEYAwLZtTtr9FI1hG+DbT
gqPOdMXdGW8P3K6oDvrU/WGGfF4AcpL9TAwcKF/0HJa0RoiML3S2aq21sck84LgV
vM7O2SYQylRwQnh/HpOLvREazxPz+u2SBFulD2VQXcTIgpsQaVRCNJy+YNZYXkLl
qZfDjk7h1Lgw6K5P2+GRvqBlHxAZQPzfrvuYDBtJ8W4OnkP23YqJPGuEcIapF+oz
Np0wobOZOrR3a6dG8926BXYK+ea+lwyz3C3vy9VWy6jmvQXri7MPShgBHECf5GTN
n5SNJ5vTyVHCpP6ZmB7qGMbnlE4KydfRsa/spI8VXQJnX42GU6DdnPNbfYyGocNg
J+0aMWscHHAMkWb7qboEUC9fy1iKhbou1AYJS4OBkdDOBLV3ELOfWqN0V4mJxRXk
LncL+CsAAEs60aV0RkIGq29EqZ60HYsIaWMV4+61JBc/w3nbs5zXfcft8LX/afn+
AAp1bn2kuglGwq+uFwT60jG1laBMvesoC9QX7F0Paj9bwzSwAZsqDBLEGnYegzzy
pXXGSax/+GGwlXBeDfrTJQVSXbmLOwBYaHsZj8iKEGaA1kiqkIBheX68hrpedJqk
LBDfokY8I2kKS0fMzp9Pi0sCzmkX8KJBmCBKOd+i7QjIKpjuog3ViFtqVmJcISkC
TMQQ7UDJux6NQImfz1acTuxbAB5i4HhrLShRO+1Y0O7DZ0Dc4y6upenwpF+/l513
0utOnEydVROs+PU7NDKCISoscEuRvnBtLFpaCJSKWBSMJV5X2SDMclhF00dJZayT
jpTezhGmHjKuCp+gaUy++Ng+pfF0gAY95kxHTiE6ucLk15ktJATqNaHE33iY4FEf
ota/lGTF31isjK7oIOhRRvBRagVcMshSweK2IBvIocr7J9OQ0tyPSi4JwJdLn5ax
kQQe0puCcHFHPIVPwf1PnsS/AC8+E+ZYnYn5jn8WfMOEphpLjtM2NZ2tX/koPy4/
dT/jhaIBUJVSdez98O5kloEZ77A3KNY0w3UjdoTqk+7deI7L/ixUmAE7w9m8p2cv
Ui6s/i2CpD32iLuE81xTreYNrR+eUlnVtqn2dRj+K/S2IAyJa4d+NAH9KgdibTuo
lxfVylDhmpNh0j1a7Ecnfz9ygwPFog3+SggDJds0jh88hAAOLRaBnf6lg+m6gTip
LiQytZQ7VKraVbTi/pJRn5MdxbqwDU+OEqI/VIpIZ/LAK8+nm1aLH6CIZsJgejzj
j9t3ElhJMUZuyHCj4wf+ESXWakgznM/w7Zw66bkAJnDnfkncffpg4t+Xk6iHUUqx
LRznOqNw0b0h/6hKg28mt1Af1fRnHyqnMdN/CWq5Ywv3GChGp/+bhNblOvjmY1o9
51f9k6hE1PHjRigDxSaO10HwTv6coKrViT2pI/2MnLPnpkYBJj4sCA2jToMUdWUU
/vClo7G/S3rohXU9iWQ25sm5jRG/13jKIopaonRTokJx2cQ3bogMKNYU+P572Hxq
nb2t1larKPv86kNa3pHjN3Ed2W77MzOTvCipT7pp3aDKbb7sqczdKYJ8HLXj8sL6
vfoQZU/w3WEQX8mcgDtFCzw1D0/1MS08Cnhylb5r6xHKngeOGCZ+XSh58W4A2rUD
/i8trJmHxgUmsB4GjamEAqPaJ5viJqxLvDyQbJYVc/8kDqAGGpPPGz0TPISkLxId
APHPcTjqx3IeP67Y7rzLFLBcYEANUdjwoZawO29laUEAlPX/s2cHRk9MBSXJDgeE
Gw1fzWzcLp2JDM6/vDtxoWQrYqRZBiZQ736BfSSRMJqUwDJXXS8c6ciLhBE6qKlu
0dn9euzaXmfq7hQ9CppfNtVUPYCfAvAG4pVyQlkcfsw1E8+ShmJWBflNZx1FFACv
kVsKJDFq2m8Iloq9oA/jg4+RrD9S2Lh1xWRrPOQODqVe8sf/OJKU6BcJxSs4I7Bz
5WbPWeizWYC7ARpF7JsLnmGVvG87WEZ1gkHA6R1kB2ke69x6gtBJjl+1SQ4rO9ap
h9bMR1qcd8a3dReweuYv+mk0lx3qe6Cf5Kxcs9+4UoHBHME9WjkeTDDQPOq2Nikd
lxaus7JKkkXIsIjIU6bgkVMR1ACeSgB9mBYl03znwbZHG/CSH2QgV/bublWmwMyN
Zli6MZ0L2joqwfYXMMRgNZ+CYvSwED6rapr0ugQU3a3cg09I6bTiuO4Ys4LvKJYz
b/pg0Sq3ul+gT1kpKZfm+ZoAe3gckXW/V4Y0hwMLYuH3Xod6Ar0+QR3uNTsaygxz
S7xgeW1+E6EqFClgXC6CM4HXz2dm7u4tunmvAQ/4J3+2K8CHErnQt9qTHdYq6y5T
Ce/2D1SGRdQN5BoTUpNlRsE/SmbLtaDz6IFaAdfIfOOvjA+PY3creWH1i/LYFUvf
ylvdZO0yeUuL1V5qRi33PWuIbWmhRKROHnNwbT+pot4Bm27FZAxlxU/+QBZhSdZV
MKmsNeVqsl6dP0X6MsAWAZRRgfnzEUolM6PucsWsulVtrvilRImjP+ABUxeGrw+R
vSKqnSoG60q7GZ5PXJEYpfuqwNpHUPFB8CQfgCCCZVb873uz52TsXFEovFfOsEn1
lUClIHf7kmYOfsW2egCY1h3USLPsomG2nV56jx+bw2h3c8+ds6iVvabQALBy14xz
ME75OlpAnT89lOJje4aYrzFPQDy2285mocLva5/ifsGu/+nwGXq048RK+HmgwuW9
1dPtDDKitkuJTqn8oXSIqETc1ot7OHHJm3aN9LXPKEKjU6WqT26EP31yT5t5aDT+
01Ih7zd5t1wOQYB9HalNfcsgR9AAdeLEu6nO5Xnuga6IQK4EcY/StiLDawftxoth
0IskloFYgS3XqWQKNQMBLKaqlTYgZh8zsBcVI99PoZ6/IJEr9KhaZ/DQTyUqttuV
Ofb6pdhVqvXdoLTuGSAyLMSL88KJqrqPSVr89phjxa9YWdELgdGMhL8bny1LsQYK
tC9RAvzyyUEOv9YKWBLfGLdUbM7xq/t43YsQUKJee89MFrUWFHRkxxGxAJMrQojs
GDFy54Xi+YpzYiBu2TVzYAj63GUAF8SK1KZonw9jSiRQlngq4mtZKA6tYpmfD8Oh
xTwQU01OeS6B1zo3g7mLV+KXJmNo3FW0nZlsdc9A2lDTvNqrIlLSV73BmseMUDJB
UKYdSVrrqN/pyfXRGcstaQF3Qlsp5O3A8ETfaL2OA1rkFCmVGTP3cobBT2Xk7qtO
PLR5rjq1PD2rOVfUiuPkyTCzOCl1K/4OHHA6bQr2IYZQD+k4DUgVav5czg9Joi89
pbvRRT2sa5xE8QpzbxiZUMBrYsXqJH84LnLgrFIqrgB22NEmXO9agz3Kvv3J3sXj
s5vzOIp3VpUEKbKShLNb/O+auUsCqjhLBOUKQtNt6tijOPap+wdYm70AmosVNTW3
kBl1tTR3XutFViRsYzE86vFBiA2y9QYpsRKM+5029cUcpTb1Eos0cNdNLchDW+ND
bJT7L8IQcxVnZ/8aBMDZt7+75p7In55i2YY8m5qBVyyd9qxi3TQN5v0ctcllT/Yv
2oX6suQ6WOXzwLaHfkkPiT6xwLqWwF6wgHpQtBXx6SAwFdKv915vWL/YuQQgYhog
husi8cIhys0QCYX4Kbz/VgBcsOoHlP4tj2bIpkbtOvLLcwgQ/xr5RahAgzmrXbf1
qk809YQDDGbKjn60WgzJcNCGn5ShRGx/tFoFks2rzYUjMaY6o/ZwYlDkf5w71Tph
s3v9yfGK06DhEyFwv479La/Th2lDOmKG1LChJkSebpl06qqpV81XIEC0d0ofCCps
OKW6lJYCcl9y5QF3YcAjc4R+irHw1Qz4+jrGrBptdA0q7t3P0OWlo9syGNBgWEkK
KQe8BaqcPHEIXjZ61brLlih7I3k6M/jIJcmasK4sl9uruFZjWOAbK+n+rOkroUPG
Xve4ArrjoMGTce4fkkpxXXdZy1P4z5eZB9HHmLL3nyvLyjWcmigXPnm5LTKaMfUm
7ZM1iG2L/e0YOpe5tyzycCttmbq5MmJwAiTE0LB7+o2D1WJASQbq5NjJHlXKDg3d
p0eovSM+Dv1JbbxSOPOYh5CYsFzv+tdD1DncjzNCzeOxqEgqCyZmXi/sLjao/hCl
Elie11zZnm6fMCzOxGZq6DNMcRtbk5yPoKq+rX+FnBUCPjW6hKmHNnQjOdMDo4zH
av7oMya28UUac8Dn0qRvuBCRe4nX0XYYUDhwstC7XKHU7kuZ1mWxjlKSSOtM9LxY
fBRPtsno97xgiMALJ+gOQKLm2+dbFmMaVdbmQ3aH99eY0WFfKKA/ZFHiedfv1HcL
dlDPpMKnshntbG6BvS2/tU2OV/Ng6c5MOjcVfbNmzCbloFfZT3GJdUVQ6WoNejvB
9zyzfjgICvuq1Fe+9RAkQA2/ytcYHf+ZNCw5FFxLmCUBQwWEN0Ipxm02UO4ixiKS
lPOyMNRjpE0zaK50Rn9F3AsFYGZ3wn0JGh7KtCdPMk+W66VpZGpVfBK68K1iy8Pl
vNxp8u07zzh/aejwlaAfTlWvDF63QDEN+FKBA/1zQmnttdj/V+ZNRxMe3uHYbM/t
T/hkDdO5h1EfnGZsxVhf3rPcfOPF6stYPzEn+gMslPFM42FVEEVf/UhCi+PaxTTH
LkprmQB7VTUJM102S7XBH0wkRNhi6x6ijZ1G6hqe+frwYA8HT3QmCpU/pR8hTHH1
0T/6T1VGLIdpBajPRWU357jK0cbJQI1TAUYjqEfkBObp81c9Wgfp4eUr1UKz/BbF
aEHwnS5KTpr3oWTyognUcTpzpBUtGaQJCB9vlVfnT3GqwogTRukDllofl2xDhDSC
SVTCYo58WRCpLzkqZCO+W+X2Hh1QJoCMObwcZHjKyBcHhJf0LewwnRIybsuXXu2E
eqY6r8KHlpiHw5JHuK5Cj9xoZE7XoBMu6WRVwuYhvAg+2YJvaz9M1d/9+oLqMBb0
Xdlisrvj6neJIDhlpZS5P0g4qx/5Uzj21jzhZo53et8uBkWEvxfc39S8YreVvpdY
N6zINO40AdKKkh8DHtkzFY7PAhU1h74Rge8tBBwKtnpgQ9FC6wORbSim/SrBxFX0
DFyhJACuyLHpD/+QY0JQGVpkGvn65U5DhcgT8VegpGuN462Xn6Gkgb+ddYJmDyRM
u2PJGA+xAt3qP19w47Si92QxCgQZcPx1Cr+jkFCbyPbJmD5FT3+S+RWmQ6lsDowu
NyzAbNmexMO8g5IMIWB4QLY+7hCVLQH2DVlAa1r5gRcIYUL11mtMd0JrVAzKWdSZ
KS/otLe8VExh3UlW8MLEDqu5gqVp08h48eoZwTXTztfvj1oLVF8etlKlIhyxILR3
aJhwNdBVR2RPk/dfG88Isle40p9YlA+5/tkxdEdUd948k4jWUgw0Iq79VqALbvmE
7wXKa1xD67ytyFyIGWam3WOFFHrMdb6v1Mi9G2Laeh9p/9SrcU8h/k5fkltIJb8D
avPfuaOIS7+7TRWBsQjph35L1XpEodjwmLbR33/l8G74Bn02RYrpXSB26iirYv+H
kWwTVhiHowj5CcorRRggYKRg7fQxi+mjVCKvEBfFVAM7ZMQV0MxrU+nVela+vbfy
85sa/8VNHL/0AKmXRTnsi0FJhKRskSPLSXA4D0F+qzQ6xaqRPzN7o2sWbHnoiFPo
PQ+MO8pnDxtlVISmAE1ndEa1viRJu5dBukMc0+FFOA+GgUrHkVcxP3ZQQfuJ9IMb
UNVHm55Vp+3tLg3qg8IVui+pdtg45e6zYz7bv4/rGcOXzp6n3c2+EE9GqR6XbSsM
HLEM4lVdec5X3n8XcGxWOcx4NNEQlcpVBxXS/4w1SHWjuzqzhzgcD6wyi8cv6pUV
cMD3gkVfh8CmJ6pOkW9YpPKPjdgXTaCrecX3jlhKo54urYRkYsmWVYQLEG3qgm7M
DPxvk6oe6vzK/FKEezJNztqLhewg9IrJhoqKzigU362jsBSEIfc5Upnb0baLlgT6
PkeBwi3cnWkRuFN6s/ItEzeKX548lP5gd1QG46b9hik2KIaqZPtRAow8ER55daeN
TtkDNLLqWsBkZuY86RmABOOv/hMGdH6MRWMFSXZORdgQMU3fKdxQFmS+Xpwo9KzS
gvoASaApmsu83is0LihIpqoZ0pnP7ZFrS6747tS7vNLRLHrrZ6YqNp+F2g9frt6D
QUviX/uFVssnAHMaSTpzg3lhuebxC6WyaOd7DXJYFU4lA2M7IDibG/4Rtd++sY3J
wq4k91lOiQVVVxZoDxuCcRVCGsGK+o5HsSZ5OkxKsAs7525tyD+3ijpGDk4pUiEO
SCoAU+fTtjNN4Z6DALAzjvth2nkx4Gj6rIL7CfrEi21VXNAWGKFpeUjUUICsACR6
uEefYP2W/TzfOOdheg1+nOM5ufU5zh16UUD882ck0V83w6vZnhvAmywadV5cwNVX
QKNfirqLSQijhqi5jWW7999IGs5NZVR0uM5C03+dcaxqHukuznIn7x+T0lJmw/+m
99gEhVj11kj/3AX0a/KwZiNdD8YO1qruF5iBrUFNXiRPQsaNhvx6neAYdWqKCCQz
uVaA80XexVqD2nkCXD8Bunv/9kDm5OR5Ty38monjklInVoWOeSbLu9mVUa4LAA2p
LlZbqiEpOwoLUwZa4iaute0MnPnrlaFF4erQZMLagXt7hWiVbahqqeBY5Dr2UH6C
YA1qaHM1ATkkLechnFJHT0S2NiQOR+UXP3U8xb3hSqj0VUxxsaxxIuS5z/5/fiiz
ttxHLEn23H9gaoQnQQSD4QzqBtnQssbl6+/paB8wVi9w/S7UZjhy+apDaekcYY/j
GO6FPwenArqCUs8prhO7un+3s6jFGwB29EcmbHVhir5wNGkhJbgrfhFBSo3EGIc4
0BJkM49iwZyc4yZW8CLrVQru+YziJpRo2mt4jMuqHpQEcRcCkt/u2Lx9bLnl6pp0
mRqly8NKtozS4K1uMWkzxXvCqZonV0p9kJ6vdPtU7Vn+bRWqxf8oMkkKNj9nYi66
W3EDmZgmuqbW+1taqqJI5MRAP4UyK+9aLt7SAwE5184Sl5xSSdlCFaqyLkJcIqFu
FTzMHybgpPzoOkdDdJ56/5TX8a7ifAPocX3br8MjkKy/04NVLLY91GPADOoKnrol
aV2zrMIdVzCGC3j+DZa5+3i3jG+ocLDwcjW5EfmWgpMfGJFfW2Jf0P60XQrKUkLK
viylwwJCai3CiVu50m1FnMtuAw1kR/G8tnBwGiEMGQR8kiVCq4ArlU6YrLZ5IbrU
FtPws/5VxE9U9JKFTddR5wNku4MguNgJg2jQag2/W/iTlFLlseb0W+n5jE72/2dQ
5oDILzD2HA36uaqpViTbUykZkvBNLEKtLeWjWmSRVivAfPsvclO87dqjU5SBAst2
2+YXHnqIk/d850RFJcu17ItYvf947WPU2kK04zEINKxornjDLWrF4hqrGv4RW6uB
/Hyke6RD3Yn5AMmaVy18wr8whaphLD7VSH8ibhxCQvVAfIUtfQEF7kje3XyQtVD7
mA0yjrM28mqFUBp0UvgCZDQX5jpGpcN50HfFUEfQKa7lclzoBNdLxHX0RGLH1KY7
aFEeRWjMIfSoduckeVe3l+ePRaqZJhBoyVprTrcmMkTA1tgHMx0gW5W3ZxkgFsOd
hv6dhqZW3mC2lRWnClPBN3J2e9lp36tXI5r4EeClBdHql3ZkqypNxIpCgZkvDS8M
N0Iw8Cohhdwb4bFPzw2tj/FIN3y6LdNX5y4R7Kw0ZXP1U2wG6JeAwr5s3sxGsg0s
vAlkuwXrviezYCKbDYssDoKoD+LmNaw7/SIfCoiY85hkBaa1vvlFWF8fFZ7x0dwo
yARKmvyH28xvUCgdz537kO6oauap5vPoDctmOOreVff3ux63Oh83VpcPzWKm7w6B
ZFVfkcMzt4dOtUI+sPSqJB4f+RU+PLo5YubuxLvTfGSQk2mAEitnPpwxDlcj5Jsr
GoTWRqV/H3x3IDTa3YJ6u9E3xpsxYjRRi8eFvhfX+50cKT1+W/e59oC9GKn7vrfx
QbrxRBDVp/iyImNEI1SlwRn75bAqlMclrFMfayD9cLbLXyccwtS9LdrW7QaXi6qz
dc3Eksmgbe9kEdFpYpBbaEQDaa4fFr71yKUnzxMbAaDTM2D9+C1ingFaC0g9m8fi
+YNGmLseSvCVBJPcXGWB9/vC4IjszxM8tbigt/7fJjSPdyfqkWsHZ9OxZQgLvVux
digow0lC3kl12NZlTQjVaeAA4hr2CLXWhtcCHemgAnjsZHIkkQ9gBLVdX2bFQ/i/
ab15xBl+aEhZrjOHnEOedUULyHBruPeonJVOcuCGSxkG5TK1F9wZ0BvEKOY1RIVy
JhIj5TNb4xxSDO6Q4xFjN93WCy3y++mxcLh/xqQ40MWQCrJzkeJlIvr+nSeSxIMo
vgXFE3N+CxqXubu6nRsST2RXdSRLDiac5xSdfiIew0f1n+t/WCPJuuCTdRETUW2i
3W9X2xlukuFgOrM7YGNXIq1Aki3HQrg4/9P/PMWX/+ZFHn/eS2O4bv1rnMMxbG/7
lXjgDEGBG1B8m4eBE4qulXTo6jv5WFQVzvFDfdd6rLMTYF+0C8oMsZatRbWYaB7m
dL6/zPfA/8BSO2WsgM9gJa0zk+NedbsZf+oHQgOBSaZiHEODyoilJEUChur81wC3
MwDgE+mShwkTPAkxtgx0Z5ITRK0yMvNLgIW6WAKHLfj1yOCSD4fxL5KI4vTiSFv7
Y6xexSs7F4Ak9F+dgIp8AACB1NljRzvI6e+1H+GtJgcO2kVdbKaxlxTIXIqVqE7x
b36qQaifSi+mlEkfej3PL80O+kf8B/6vXx2iYpM9C7YQJFAaCXeu9nIVM5dkBl9M
4FFDl0dwuRmjjNltNx0gNRrqXWqDp8/RTSi0cjrBtFQ3ncLnlVFKSXxvTETuOJ4p
KlNuZ1aUxD6eRYapVSUM/U+cITZPxIjari/CfJWxVWXvw3ccvxxiYvE3m33cTXCp
6Ad1QUGsfFxAWPSpQhXN4PVvHtxPY1GwJs1cNv80554NW9vKUO/0by2NPhe/7p2h
OZMAsLNl4BD39Rmw3Mec1DThdSifXUMDRkSt6RvybwkTYcp4NQBcWBSJy90/hFbA
cmUuH7H3k0l+yxNgYVhanFHtQrK9+8P0Z5AtFxnp4mNAxgL+hmgQ401sbacGMOjD
FkTj0gxDezeuEZOJYX4gxP97iDYBz7MO4biulyFerQIRfFuWsF+j16mlk8d43RD/
0xSl5tcSyJbF7h2+QRCNCIlG/ECg2NTrD40bq/Rr4QHZr94nSzbHG4XQcuB+G0H4
U3uZpJ7x2xLw4UDRlFoFGmzclFUdazyM4VburgPk6+UPU4224SrTfUm+n/2DxxZG
Bha6HQxCW1h6ewdfj/KH/xzy98Tjp+OpJLb2kPd2Nx6jw2CGq++YOk2VT6Dv9jLz
M88l8dAEDRFIGOLDDkFN8Rtuu52SdWcK4cpq7kAO8McXBcglK+muVOE33umKXt5/
qhc/nC8KN4N0uegW9DbdX2wwVCAjh5WFOJbc8Nt9itPIed2jyHy31GZrYjw3rMCG
GWAdolQYozkC30i5/PMj7YdoXgvx++QDgDNpZ9uRNkFV0GSihvXi0PNKfRVOVoCa
1PmGhytb3CiGdKpVp+ks5x2mGq2F4J4Wv2Yp6DVL2JnBQsBEiJsp1qiyrqO5kbkq
pvN5g3EoOYsm3Djmt6zWy6vcWyzQL8z4w/lwoM0majDV4XyDIOFJPaCKDWUmBCoQ
7lG6vRaTMXjfNNmSRV2Bl74T+ZawEyOJwqRxWnyZBMt7YZG9bgMdFbnVbc0Tsskf
hxadMArd4BucBMMBDC2LBJClI+AjS1FNb0k8ztLEyfaNZku3gVBHP+7wAC1yKjp0
3ToeC6cyjGTehDcgJr99brD3xREeEDyofBmoLoLtHtgfoNZhI1Wyyohr0uOUgSaJ
oSndBp4fL2qY1vU59ceUb4B3hy4uxfydpGekH4X1ydAYFsxjb5fLy1MUHGSkWHna
R+wUh9lg+9Swj4KjjQMyAs6gm6xHE48BdRS5AFgOSqGN9G+6pj7SxpOsXWW8eDMU
PhBmoprdEB+VClWDv49hUB0iL5U48vqTcGEb1rdnGylz4RzGTvUf8N8iIrNA/8Nk
WQlPbLLJmfxAEg7rcl9enHMTw02BRQL8cYwdtBAkrgDeAxFnCKXHMG1CJ0W+XBfi
n/6oCycWiNxHPgqYazTUv5RG2tQAWUDSFvT1144IeNIWOJfmvvYiyLWTfOOmV9Re
Un/FoNfvef60M/Shj7Km1X69H8c7JuKmeIbMYhAtdxEHpY+R8cB+vZjruFKhU4g8
HTWwuhZXG7WUkzU5uDsd6HENrYVTKhSngE+G2lVGMBKvmLMM0O2Wmib1VbFLKCnX
OPPR6O7iCDz98XsH/DMtSoFLXXJRrn/XX7BLs2ZBNqaCaEJY2nYRMr1o0zEHbeRz
66ZUn+sRPCneytXEBO3EV8eMTgCC8/pfo5FqOw7tF49in8FRzrGa+0mpHvwkJEWC
0asSLm2qqT9td25ic7gJ2RAEcInDk7eeniCp8YTf06JTcwrmT7Aw8VLZYX/UsKj7
Oy2CyVhoTda/s/T5Gy+Pa3unkz4xYmBlHai3gSRRcn5mJ5CSoIuLuv0f7DcCq5t/
/JY4ribsCDRK98on+Y8nJVC6npqn1iEwhEKMVSVWmfbqiq4FO6PnlsijCbZ2q45X
ELKkSGcIN7ZBDEPyQw0LsaAyD1kITKN3m1o0yPd4WG+ARyA5U3/4yab9Wlul8iyA
MGc+7JFcYufDtGxHUvM7lYTkzYiU+gvSgioqJOPlv4EjZpqKUff/QciYSTLKYDDk
UHu+aOrAWCYK+xGSOiCqvDxx9NOG1ldm+uShayqpixAjWL7ggla4J6YNf4eA+9Hl
rF3xuvVNpDhg4KTyN3cFFjupL3OJGTt2IN+kWWd6K1OYIxK3YxSi6AOupo9EPWxs
R9JQX+gmVq9hPazijPz2Sya/qZ85YJl5OCqSTiaCw+waj862Byp8kRym2cFS0BW0
mC69bnYtg58ZJiKPlLOCn6JYEgjeN2OqNorSPiq4G3Py9fNqfHG4ic4H8p6q/wVJ
85RP2/a5INCIzKAPkvl0ApLr6rUHw8l7PiyZyNtgd7b8NBaVHJFbOGy5PLufB5m0
VQrjcTD9kmD3bQkJkf+GyuFyZr4vy+T+rGafW3AcNJCVQijWaQCbJtP0KQTRCnGT
7ZztkKToAVnUF62bZmsEKyt4UHV3CCtHZLpnTialMNiaf9Wz/a0n0DyBmUTKfjxf
YYdQBV/l9Afue4c1Zy+rfIFX6wIvHPP2CMX4LVVquAZot6cxNQLF2fMdriyqv/Ml
K+v342+PU0kANeMfatpF5IXyYvafQUBwF11osmnLQpdac/19MmtL69/bDKOW+gAb
6MO1CZxkTRA9/EPYOpjnCngmmicTmD7B068zx0Y3xbJlAeB4zSuqRjdyQc6vZ7Hd
ONEzwD7HwnRKVUjVcvIlwDie3kfwK2keCDtI/5OlOFWfFbRqXpmOK28e+w+Cj7wX
dXhz63CWFLDvt+G/nE2/r3aKopPYaKp3daTnpicYgsFj/ajNbJV9wEximdSAtOoM
X2ANYJVq9aeVM14LouaZTuNVDaAgUlejgjDH5C5SKLYNkdXS/zNfl/fmsdlaU/Fg
qkfNljoxYaq+Mxxw6r+O3JC8Ozn8Uk2iJm1/c4KNxJ01NiPIoLCA6J9lk71mbmEh
9xI/appwg4HGaqNjwMmItDN5t7BQ9vAy8PNB3VGHPNdjhddm4ZKPpywB7/npaHHp
dP5LnZz4DxJuH6xnCv2BdwYDHn65tF9YlBI42gCxjrDLf4q1ddUAnMhQsF1WKpLi
+fATBh1VBMw0g/fiLQn1+622UnH8HRhIrMxedKQlz5CCsHRK65OTrvsHqyhRKr9s
j63zTCJjrQ8J+lnQAGE89sUzo8QZnw0siDO7GvQt5PslzrzavvMBFDdmAIiKOKln
h9eWKNcAt+ouYtXPKsJXAkYMA5X5UliBmk3okZF7zASBmFrhi+d6M8FG2wlj3fUn
+/yoymHk+4jQrVANLHusw1vZZ5KG9r+S8hWlPY19GuSTItZJc1wUi9sAUJZA693Z
rF7RLql090pAsCAYpwIb/M6e3lq3j2Xa/3VOb9ZmAyOs/gEutorImImSzMaDAJti
nlbxmITkv1beOlePGx3+b6FQrINjkvr5yb3okaUYcV2CrkbPpCpFT7+U7XKGkfsc
4A/M6I0FTOkXi+Mxm0qtIMrlQZzNH/1OVGzdcoYo0qTQjxzQp5PF3MTa1SjB5apt
sqPWQI6/A0UPPiJ5j2fK3Xe7RbTEb8joo4IQSnJAP3ufSOoEVH2Z75tmBXY3Fz6q
5iHjWGx4QN3GT4OGFnWjMwlI1NAOi9JJmV1VGMVxdSJ3o8nYiQc+9E+dd/rIZFry
3y925DG497Hs0svC1MtaHzi3FCzj/0vaBW9DHCXbmnFZUc2gaHIB2y8a5UtbY3G7
12/KTAJ1uz5xGtzgTTymnPxRfvEfpf3xd09Vypm5+dbiFK0ClcuGr39xWop9zg+g
uv7n31Dm0m4q5b7tdIuG0qBTgdCc+A4XZKTyVAE6kXtnC6cAxsd1UsapUEcg1a3q
QUf2PD+f9iUNDwY2Mf6+Id9/OAwkj/8vk/gQ5uFTUftERg6e9ToAE1CaPCgp06xJ
gigCPXGN4b1zMDr2ZvL7JvS7qffrUg/uaXQWXzErcubZwN2zCNCSKwqgY32sWIjj
xwjPon70nn6BlE/qIdpZaSBxBy/7MCQUlcCk2k80xbuHdPYcmILpxXzo6fUVLPzS
W2cVs8dfIDcV5lGwMzLh/LwA4milhAllVNvY/Hr8tCTmP2GdvrCx4hepp0jJst5v
C3MangTCUezMX+kUs4aTzPJEstBf1Aqlo3EAUCjwTev+fBFCIEeec1RX6AJ6Rfc7
qE6yxPpQLBT5kWtC5jz0NdbCSGZKqFoNjA6FeD5D7+yIxXiEVpxHGr3/GSXsPjUM
8w/QFWKwVvcSAUskQ2DoBdbp2BAKFdJncMOg9O3qFoK8yFJ7V/BRHCt7TSl3AlzR
RdFqH9EKIYUoPrFYUbwS8suWPymdjT+9JV0UCWSrsYGx1tnyFPotg2WgzuUNu7qv
+cWB9YCFAo7n3niLi3mtnsCa2Kl2PRWw6YUUKLhflB4QgbsEKdJKc2WjnVLCfSy6
APBRqsuvnBlAG7ApDJrsBzek+z+WEmpbmVNO/qMmUNqXCE+Siu7tvxRCDCVrPDCS
m6fgeiYdyULUn9FNrZYQ+x7JoBR7E5bUCHNx7N8Rw8aggKZV/nPV4s8+4jvex4E3
j6vtq3c4qobok3u6xH1hlD428UFhvGRPLs8djWrGf+Eocut6UH2StFvl9VioyFH4
JtZDGogVQBsTV4nCic41+SaTzArm+GfC6Ojx2MGpl/OKypvgTl/CQxpBb1HExJwH
X8XH222mMRDFYilXASqrSssq6JvxIEKzPInjSC4sHbbuhsEPvBSLE94DgwnBaf/N
vmWS0De9BEF4f2f6UHYQ+5sdGHbwekIWbwr6y2+NJKr7TbnhkSg8gHvAxzI9TErY
ah5t4wxz6qlG4bA3kxilm6RtgswYImSaW+G6MoXX0lPPTKAkuU+K+6LlQJKDXrAl
BHzKsucs7/kp972EYpB0Cx5E4Jc4CMMTtDFhqj1K7vrGwV6JhnSCgRRe2m0LXYC7
UNBw1MuaXYrwEYzbSH5ISojnAEUTc1LLJWTztmiBNR65gn38wXsbvlu9pP3G8Pz2
idvKP3gS6DGibLbnacftl8Ak69OgmgNn8HVh9fUxdoP4Vq/aWKYijzTgFXZbCC7n
EtM15HQdiwQrXoTgqU1HheOggiGvNWb7nTWCYJlgmMcSKmxvpzldw0E3Ydlwft2L
6rArx7EvOt7AANDih/lDHfXlmHPClYQtw6wIKRXaVI3SrbIl83jZOhR6oaIJpI1w
m+H6cvriJnUMmyGPrFTJf6f0mEUW6pVN4lIWEVgHFpOUu9D/3GI+mvYoQhjpSTWb
X1DiTMZK+mpHvljZHLUrwDfL37E4vHDi++OSI5ssH6HKuQSgIz7SYcTEeXhmB2eU
M6vy1NIuNS0Iy5iEIgoG46MNBbFqmcphvMoPVvUDtzEWD04kTafx+Pp51M66d4Nn
DUUb2pUoSNCQk3+SdZCbtcTRcFF3PkRmd2aT330RBdwx4X/UfnFLHUFy60K0kVfh
QaypwcKJ8qbwXgdrr37UNrtIz9u0c/Pcaji7plAW2qrVDWkdybFWhn5p3o+wHYSG
9vZOCdZibSTkYlgTdcN38/uGQ8cRyRHljmw2gfRJq3IvIFHoKNAmvjxDXg9+PqXv
yTCe7Xwhvl5Ll2H/YgFAib+t/mLcxVx3bcsutWkdyWg+enK7YcH+jlz/Texo3JWh
IjoFd7rRmp5EVxw7nL5VhhBaKL6fVvBPhITein//847Hmy1aYA6JIUkvpikQdaqB
zbThzDQVMUNx8diH4b11s77CqKKjSkmbxPBTcuBC5O3ejcftYVhn9hD4uJBvP77l
/q/7gmLCs28XPYnU+zKaivqJHHuVVaQKey5SBTyf9WXn3sDq/8WUr9TAP+tktK8H
+Psx7WA/uqlLFqXiqPIxgMz5No2LOt4FjWLnyWpfW+Yf8t5wpq4W1X7WImWebeQJ
UPpc+cRZCGwprUqJphB2ANuwVkJffhgM9SQy4SfCjnUDq3CXULGOXFbY4NrjJOFa
Ka5lmcpNCCPpRSU2tD6QJA6iDa3tLHgDnd0Db9kUd10vFIuPMblT6xKteUD8CezC
DxzETCFSr7PIHEYH2BHTnT4KsbfFn56JRFHNWwOlBm/gDnouPYzV14/yGlv+eFGr
Gx2cXC+CbgFtHUAGu5GhXdg3vh4QLBvlEkU+DZVp+aJLKwCd4BcGvXyotm/su16H
MWxbBH18k+x0IyGwYxM2CqGbNatsNRZW8t8/5S5T1h4ufH66GlXTdX8g10WoGAcx
gkXOQSyhi6wBtbHmyvqd+tqwEGCpNdbNatLF9bp6CIjmui89u+VzIbs6Cg1v9FGX
IvD0LuXxpxJkK9cIro2LW4KPrhBwZ1PF0YJ0xJGSLKdWEJ4SFsFa3fZT12i/jf7q
zmv7lYD1j94kYS2LddWcvOkfnJY4cRgoizQqRTSvVXLzV3VK6qO4wdoMjqx50LCE
8mvXIJWePjAA7DerTs04BP+Z19rLGwOfqlTNk6fuZhqD5GQ+feviPkTos5VUEE0i
DRY39sMxB3SAvnpslQZk/5FGOhADfZzQS4Vjn6HqL4w5MGwnGdWvNmKP3UaKoJog
ysL5WkatN/x4RILlKNh0jC2CaU8vuhQt3J/tk1sfcIH9Gh5vC4x2hXafFt+JFFcj
YveigvbgaHBoKYdZMihn33BDa8+ttm6eEYGk+Zj+MlzCNWcJ9Pp4JF7f35C9UdA4
0c2QkFSz3Tub2Ka4fL10fjX7sXBMgn15KXS3yc/JCLyvNdP9mb5yEqPuZ5Y64kFq
HiXTeW7iNVjhvs60sRFZPimGzqB6XKrAZK8FbGN+a1ZWOkPwpBMVbK/IO6H9QIGZ
yxKvNWSbNzxaTCR4ZvRAh+XxTmfnqzgb4rYv6kgTc73JKax/wwBLdhziMdeY+O6W
ccQUavyccEU1o+8+ic13SQamwHONj581UhfceHoHCRp4rx82ENS9sc4tN5xto1QH
Z36rRFpURM/j2B48iPhZkDL5lOQ8wf0aBxuTZHsdjZFiLfLdMSX/j27ASlzGWZXr
Nuu0lJFixQSBqzP7mKfoS2Gg5GXu5VvILYzwvpJ7TCPQD0FCYbwKhbipvtp9jSGR
OZj+m0Ct02vxCp184SnIgYz1/rv/ySbMh/BUhf61nG29mzdcY8/BA/mUW0GtI6Lb
bDC+rcdam1rYOZ3Rvz7wZ9Iozr8xVQ9TCxRtTXCktuHUca/sc5R1Ksc7ndqDs177
PDxwwKg+zQgfdnQpTrW0jQUN8j9mun+ipcTVwHxTHdJg6FwsXhEGixhdF2OFq8N4
iBq55EvYck3XDTgAQOvQji2gEFBKp2/6WpL5jb9Xj9N6TbWEHD+58JKIZs5eMqF4
4RiT631tDiXQHcjYdMuaR6162wE31ohDfk92xctGjRRllr4Hu409vSBJ/AVRDMRq
LeNow8esmQIRvDKhI3m+Xv2vQebazJqwVn792Hf+vZ1MR3bDo12wJmYJlXce4pOh
c50l6jATvjsJMQn4p/PFt+Zw5X7KXHWUYiqd+CIKMcTCMpFnpeYKr1IYjxXhW1i/
D56cCvgaR32jAdXqM+Kh3Q445zNDe2B+ocP0pjfy0DVa/Jst9YmFoHPQO6RaRDdX
4obuntsF7sXHZblpDCLoIy8WJMP/PGnGSj6Ow2N7bqdFUnmhAJHj5c98nxe2MLme
4s3RY/dHP9R75skljUFvT79j9OgBQFyU70xShGjT/ldlw3w0RxPpklH/j1sidZCg
jd/cNdpGNC5bTYU+VznWD0odajlj1Ar+ZjPE1ve2nJmDyFQvVsNiAxYHzfgcKAXh
a32lQUZ6kdiPqHEffcvUW2ckORF5hmGU8wAc766pMCJH/tgOAl+Um3F6E1fezt8S
r3BVQQuFnTCMptoCyl9pQNiAuF1T9Hu29Ogn6oFCRtiOv9+/9kOzW+3motv2SP4A
J6Xztq5UD1Me2lM35LVdcUhI3wu1JjeojnZbBJYuIVpt8RmMSJL9eOm3aP2q7hhd
wZG7cpgz2mJzne/mM44pNRj94NDs0DU9yHMx+/lowZyMPHvNfxqUTGjiACzN0zKe
QVEy6JOf7VLTngqj6/RNonhrLhs+FMR8mwV+A37isS50pLBpElvLBw2Pbl+BOZGJ
H24QpcBHmvdFWBuCdjN+aMUszvsOFeCOVjMU5Y72S/cMW99o7NauPKUeEdUa1hqQ
9Xv9FW8eziS7Tl09m06GJjJqEvW1sOy2pS7rFBopR/aEEe1yk+bWFXVJKCHWWUAv
SidphVqyIplvLocQLkju252pzAySbEpdIdRKAIcrJZJWok1Pe0ZunnImshCkEyCP
yHmusSLzcEp43ybZrCDWTVWWyBESqEyyc7796zcw/TEecL2RoJVY3FN9CK6Jp/MB
V/+dp2c0jr2/0C+gR7471XE1x1SRapCKlICsAAYy1LGwdt6DYebSoxycze9/gOBJ
/AvsJVdDHPFVlpcFCdHSLKoaPQRj0Vlh67PvmecL+bwfgPuzwIyAmjVpKMrL12HD
WU0qk8GLITk7YA5esd6Z/rsYHpNWwy1jVkCUVIkW7NMyQ7Gt01eUtAHg0/nfxwqJ
2v217cv3QHO5WBedDu6GeGnXI3ZV1WC/TeD6sstoolyLigigCEgPa9AGwdxrwhp5
P8IAvfhU34Ha+5dTYEK5/g98Mnfp3RQCL8jPWh1/Kj2RQfAKGuVSZeYKQ+WcKPb0
MUZSJa5sPhD7MzisK+u3DfCMcwMmfvK6yxyHfOPZmOJtQhVGGoeYjFYKiMVh0pSX
Ni4ZW2/XBBJSjoYTRI8LVMVo4K3uaaDVXhsn2SV95s+M+VtEIGGRdM2mSnliF6TX
jnmuq2p+Os1Rtp81XGjtn7h5Y9WF7McGyJtSSzRFbNoFtJXloLx18b6C6qqvG9Jg
bDqjU1drgk2Z9baHu2td/g3DxsXP04E04pqgI71a8BLVqTNOZClfn/yHLaF0k/D7
uqub/Hbci+wpsicZI//6kv53T2T5iQkT5NQ8QL6h+92cokAifKIQt0biMEieoIje
V4xiACpOC5Z/f7dPqlx9K+L0O5nMJfutAuzzG/njAsVEWsSH/g8x1JYVJlNn3L2s
qjFnocem4WEptLCZGlI68fFkS1SF2+AZD9Epee9+aadqZvxECQu/+d9+k6r3cMIe
qZXJyPM8IHnwehoweDjX2gN1Z0Qb3OTxmHY9iOuuH5u1r/MJsAsV6PLbCy1jnje8
uk3T9q0QIEMHtrf3xGp4uTgFKbem5i+0YegM59nCuAhC5AUkpDUz2RZZchdnlE+9
1evzW+BZQoH+KQTGLg+WTRr2abCgNgVqhBzoEKnrafuddFg1IptZdSopxSRHR3Ri
Htq1dN+TzxdhSGmbmtau+RicHzYoA94FR1U/+35EY+5OvCksEEMr7H5iRNTvOUPB
1VS5VyWz3017ywueBd5sIAKMf0CwcCgDsl0rr1YvJeebI5r8Sq2hDt8GdINy1ZOt
W9dPFIWP4ZgPqzaljBAeeVxsoz9l1MmLwMDov0Ghqhve+zOYCd2wUk2IwcVn7yFJ
tnn9DUQhypNjmIDTp5gm3RiszgmczjXh9YjCLbnaWoHNNiUbCF9QJfECQAcSwqmJ
aXoBiZiqO37Nf+IwhInx4I+nmauwlqdfsKo3ePj82LrO+rZwL/VVN092stqdta0O
sa0LAT2GFjz2kucJhoiHOM+2Y99xZR/t215R6gPE+l6QIyK6IMRX6iHs0Zz30Btn
JPPjBXNXuXaq8ad7ZxYxVvIe8skfKwd/yw72m/IDGQJL+M1qqgLst0ltVgmpXBhp
99G+K03i8GAGvFLbVx4uJRg/J2eI8RQVkqS4wYeGaHhJi+avzhwF5X2ZCTjmE3VA
k+5EYuELFJIb1Wjc+Tv1jdoKg40mkC8RrlDifddsyl4lL5P/dMW5AA4OYKXhjtKh
HecdkKSRZcDUBxj4MN4OSQ7G+GhTvL436VpsZ77DPYgpFxTke8skajWR2NZ4PlUx
EC9Lk/GbiTkb/ldbrmGszTfLSR481a72kwXm3tfduaWTjVXL5WNMso6hJOKa1Hfx
ZAjVcu0kK15UoV1FoCbTWE1jAsMaTc6Qh7p7z2iHKe4eVXmSf41Za2GeIlXl2Hq0
XtIaLPjnnabF+kiza+wOmPSd6hcTsSF1G3ctPqIXkF4KpMfgENcuPS50hEyQ1uRe
zxrJYnYrDIYwzDoDaH9p8JJFt93AQxh21E1OEQjNb0dxIQ551c2CblfdwPbSB9jJ
JZwhimsxULDMrT6mvHU37Eui3FBUzlXMBxo7rjBIPva31U59GwJFGp2um3mH37bn
VQUEKs1bZRtwSl4pcFMUFsqEMeJgOuy4G3aPCa+ElNuQEkDnFOIVqVjj+o3YSpnO
7IBTiHKgMDGz0koni5aMhdk1UrRwmmvnJRGinFUtZ3M+kRbYOI9OGJTDaUA2qY9S
w3Qeaq2JIyPtdXSzSMPEGmaUluc7ZLGGAm+uINKGYWFFm9NeZP6LqpM12qLOBsQC
OkHmr2RprATluk7Temb9xosM3exZT/tCUd3X086gUjFic/wQLoVk0e9CuMls2W8z
jWZfDX9H/8l+AgdAB5QtGkxUr8crafF+NaIQBsiBRTBvJwfb7tlxP6lIV338C2B5
J80ZCtKI5PHNMz27Nb+bYwLEpow51zV3FQ9WNNWSa7+Au/+QNh/hhIg1N6MBi6er
7+yK7MSUtGf+S/baR9IcvgCaNfFSI8ODSMiAGpxq2otLAcJP3A0M+5qKSO58HxVx
x2V+s0L3uZ/6OYg9wdWkW9CUHRo0n5hxYuj7ux5Ade4o7Jm1erxZIPmnPWen3+1V
f7QpBAkU22rVzKBQs/vn854uewZx1anzonO4+auuyteugjEufThs06TER3HpF3pl
eWLqg6kCeGcBPRoKKwP6JpiasjWW9csuCUDuT7FNmQKxdYrR0xbfCWMTTT8w/B2h
QjPG4UniXximnjHp32MZtiubPoW+V6VaTYp+M3P6U/TtlHeKcy26YZK28scgJNUl
d21L0u/rLEioYtMVg400UXAGz1nK+ZR0a8AV7WebQZrmuoEJzfvuHtPPqgIphs+f
tcrdZxt1HKyYN77x2lOAkHJorWp78rgiZQSyOS6HbaaO7ClE31A/sK0MoizxQkAJ
EKWtAFkJnnuZBynoMA2PZUeFfeAZVDbPtpUQOdiqTgrkkT5xOeq0jYhnEF+dLSng
j5PkMVD8KQ42uOMxkKSamPaoelqCWSN1RSRBAvml/4FoTv0igfsygFew2igU1kJa
ckYXX2W9650Vrpw6ADHBoLbA8bnzU1AkqSt2AC8YsqCpqRuupWL5vMiq8zboq1FN
kDGry9p9WJm4RLxZlIifPLSCuO0XABZlkRM4zhD4x7wpkhmxxiSuZaLX0nljxHNL
3KNxn7ITpZhJwC92mIFQZxIR7JKDd2wFGm801QRuz0FFE6RxEV0t+ATo3o4mf846
VB5CWovL2tffdS/RGFVjoW659epjYYCPRgYfzJS26jqxQwk0MEWCwFoJLCcO5SVq
ip2VXTVx0rmQzDw9zU24OOaamDQWs9lPsdGIAmWdT6w009s4obloUmP+iGjlVyWT
fSMnT85SYqZmQwDVb354tCk1O7haMnDmktq3Mn76fp8hyek/HLPN/qUH2gs+lx3c
nDC5o4sFx7+Oh+UudbS+EkyV/mzWkgFjb6Wvblv6O0kukqzSD+58ZC/JrLYC+9YF
VWLhKZjw001eo6EitOOqRHR6qBH2CeNLYTQtS9STRmwV51VO9CATuwsItVmDoNjR
uXsKu7L3ydv/+zF4QNvRHEoWYzgqkJRMq3f5WePMrAv1LFZ16DvQ36isuByyglsg
q1ojvYeDqI1kCj30t6tOIcsT3i9TpMlb2FcT92hWXYK57/YOpzyu8csQCYZmb4dJ
VkMFl2kYl7HYqNnDKUxPjOypo3nG17nncKJDTBaMLXHPBfQzb47/z3/xYBAPEZdt
mGM9+tb5JYRtKYm2J/8Sz6bysV8h8+naQPz9XaQFwEpXHfD653x9fffRH2a2XUad
mzyaGEzjb7v5XYovWy8WQ+lggvzAiF+5F3K8FPyxCLlfM/bDHGTgcvVU7q2WfPC3
nYcuYkLR0nv/o2l3VmiK3h3RmONElRlqP5yRONaaERaayK49bm1++EeI3twsuDkI
kN1PgYJl41zkyu4fEdwPkBFtsRCfKA+SPQBUhnt5p76hSPx7uA2NIHmfQyIPRghl
NNto0Jo8CQN6bH7MHFvO4rQDm2xXnq/yHqGTqXGTTwPcictSB7nnZfRcglkmTVFQ
8d2yZWcsBju+iOh2ewetMXcIQPGuidXtxDv6eMNpS6fiiUT1P5iuNEOF+VbmAbu1
V421QZkH37FgpRtRaqYZsGLM/GbDeqs/9EmbpRo+kvAcOjJhAh2TKTB4Vy9gGiKF
uMPnxnfvUboLWMQs3Rl8u/YHJdi8bSAj+H0fpIAHATHAP3D91Sm/XYGE2D+3R9Zl
UEbuPNAkSi9c7u3zswo7WIfrBTLeRc0ElXLM4P6A0pPItA9LcMNcZVIHi9Dc/3fm
sNaRH6gAxN5Uv6VQFMU90tpMuKy9vZ5NyZdWKBaDgcwT1/BeVCQvWLGNfxFoWy0t
4RgLff57tRxgN3YyDZuspkccz41CFOIxvDMEndHyiR2cPluoErYx0IppxoL4KG6+
3ijSwp2/Pc1Ii++aq5IAbPaXEZxa6gzhP0gsb7ExQXU9dw3vZlYF6DRGBeshrXzN
g6N2vXytC4jR92fdHLTUTYo1HhH8EWWZVKp8FgVkesWSsv5czhp1+noDQcDaj0aQ
rbCBQ4PROo5iseUZ48leETj0jIxE8TmNEXMHaTb08lKVox0w8G7VgtBKTJZK1SYP
NYPG5ljx6NgpjKg3R/3JrjL2KvdNjuNO2bsSSEY8S9vtACdWAY57GkC6tbNondif
h4OM9N451uvZmWKEA3EsDL81BrrTE9SjoQA17ylaK31yAeKObOfnJWBNZHY7JKkI
NoRnjebzSeEP/BWg8gdGIxcDQ0OeZWiVF0ylUBQ1NvEDt5Mv6McS7M/yl28f6EMF
Zo+v6xUebdV+jyRDYm/HasYRUiG94ivO2Bj1upELWyT9V+Ou4vsCKJoxC1snglp6
GueWfSVpFOXVt/gCFobqOfShkTMnTjURjfbw6Su+4veBo+W+Unj/WenBewsL67Ha
lVhg6PPOc+Uu3M3GynG1sMdFQLTMwDuMApoVphs/bK2zcIx9TjQZ8DmkS9rFblxA
vJmI8/NGViq2+ydlSOfNUepQS6kfOcxCxBj8y4QyjDyOQLZeUUU0DtxkP2Lstw7w
C+AbiZIN4wenKR7Z/mlY8j2xWG++bVL/TxRZqaAOF1hIpTRQkSkUESmooDnZpEXX
34ErfX3xMt+pNeNnuNKdn56sTr+Cnl96z9jn1LyqIqyxjVhpp2M6TKMJyc1Xw54o
gjIebAXdZ/5xcNX5GwHa/dhM80EdkOkaBHfSJwuOFKI0yM1gGLl5GIe9Mc1oxHoa
PSGgB/zNWEaYVnh6qcH8aFA5pdkcXLbcjcI4p3QxmEWLvSEiyvUwabprl5agsF5S
8LS8xyN6rz0lFVS/Vb3U6HhumRgV7bAE0Zbm63nll/d0MHayVSVqM2JNITnE4PlE
wqVeu6uSTCNlwzhvoNFmP3/qUDYXZhe+OHwR0GEMo4NtWJtqq3NM73ULfrQSZaG5
Br+EltgFsJcOAnFodbp4pr6l1AOusMhxs05DNph7rAySaQVzw8DtzlhpbM66WJRJ
mIG4JIAGBpCfH+c+fzal86uwygIWFD+PyndmKJofwkDplr4D6PheZfFwlCUmgOpe
F9QA8nA60k/jQoSBZHl3CQeCYf+1wEzjO2lqv+RNFzUag84Ymc0R0y4oqSWVnmYg
aASIQs4IMx6i0v4tQx3CQiZE7QqZgVQiQFzo1pEy2a6cYL0zaSrgIabEkxC3/6BT
z3Ca2ckppG1TFCOeJIPS3F5UiD7otqHqKHtInjFYExXV1ORWnvja5BMd2rKVNYCf
qrb25siUqc2yScvTpSq5W+qJqVUyFxIyiwlvfNoAkzq8XhAevgY7A9IsyDu1NrY+
A1lAygapqdGsNhmweLN4p3Gh+5KBE0d/eZ5OVZjjnhuAfeytKmruaK+wYBju4H/3
rB+aEWeO18FTp5gM+NFPKp4qGwXJ/EM5P8TwYHqb/tHDY8xGl52DSXUU3n1DWc2F
TYsjDRayexoU6wgepwg4DqqVQsdGuau2zqB5uM0S3JEkHuj4JKiWFg2SeLg4SFVE
ve1lSmM579KxOucSpi8cOrQ+waAV5XDuzwS7PjqDLioQ2TYsO1D8OcNja0XrfXz6
LiH4UiR5ESYTutVf8VbFeSgZafbADlX9BgDmx1xpaJOTq8bQgpit6FOZ0dC4uMVe
k4EJ76RludK3O/vYSzytsKJUpJ/+x4/peBWiVbZGG126tH2H84H4K9vzrafWGN41
8HG3IYOb+aN2N3h0gJfsCeJeL95R1WRz56pVH4n3BubBRGrAt8bSbiqCImKaO+IK
uAKbrmaMiL7iUg9H+PuOOX87rdjJziKGafKHlCCjWJ1x3sDwiAe9c7fSNQaa9MIj
dz1PlLbBeunzjFPGroqVueKt6/4t9n4PsaojnDnubuqKlCTIyq7dw7fGiux4X66F
CgcNPK7ncxcvBuTphoKM84gy81QNCG2jprvw5ybBV0IoLxQK6gRZ+UhifEk6Zj31
wvyQDmwJ4zUSz0v8JEdisSAWCSKqIDSV0czvXZHEkauAoXpOZzqEXFtA7OxEVgsE
fBufNQS+bAxNnR4zyn0txQ4nzi05g1YpqM16oEZpz2BGts1QcFYumZH69kJXQWlD
soFBMUB9U0UzaeOYbmLN/GA+Sq+yuytUzouqX3g4q/Leb+ChL37oQtyzhaG9ZynX
q6sEs/KWyf9xi3howiYD4kQ3GVDzrqlTyzVwkhI5HhM68oA9eV6ugz/OqcAvR8wr
JsOL7+FS/zx4DgEnqgZ0zLi0cqJ+w9kp7d0Kj7CdyNcDL7QJJH2XKcyLyqCx/3LZ
nVpb2s5tWK8qgpGxW3EYq7ZDt/miQS5HeZRqcp7DGCx7JZmHCdqAfC0YhiE1a8n7
IDGwWNTf0gu0MHvTOWrAU21wuwFjqC3eSSM405cExgvaQRm4c6dfU1DdAMI1o96w
gKmywhepJkTpemX7i2p6marevWlFPh+naRAn/WZM88juxCD494R7XuJM19p7SsSN
S+wglpoa768TvSGaluG7XR+XuaI5X8lS/gLatYfZp/ISj7D3+Lz81QLhYWQ1g4V7
iVBxDQZWhJ86gux1c27065ScsD80oPCU0doPdPDsbXOW/y46sPrxyrXDhgmiIKax
kcoGFUKrLLanldddpLExmmqICjrFGkSKbecPuyNtDdBMxh/G6S1E5tCU9ihYbCEJ
L0QNq9vcOTYhIHNxPDdT0xJc/5lYESipW76KO7J95k1wis0fzzJdwAjETr5QZRUa
K0AZtgV0D2aEOJLkOLTUD04kzsNFg7pHMT8NEzR84KL7xnKNMTjMEMFjnpiYpQzr
aXQoGOQJdYQ0g/UkrgKzHuy6H9Uo53hCBkaQZ0jdb92GuJNkieFlxuBpvaog7Pnf
KWCLChUxC9GXMbvwwFDGGZlwFuOtr1VDCLso+jXlIPlDq/2TZEr5yIsm4WCioFKW
cpXxYUIf6QlCPOwIM5UGBxGHMDDSI8m/J2f3loZ0j0Wm6Fivor9d2oCnP1q4xtQG
mR6TvZ0nfXUa8y9iWX+GknA5KM7LSaIyAbC9mCdQ8QVTCovQebp+LcN2XqrofmPS
jzWx4tzQqqe1MLrpDiCssmCalSGoOTu9WI2ILn52JhAKEmpYMhWpcTQCDEZVo0db
jMultiGBYkFhdzIL+L0dVeWazAwbrKgLrQMC0c0i9pGqX1XGdKqESVtVZ5yC/ClI
J2/Ik7Nw5Wp1nBUqTQv91qXadGPJrST96flrgEYBkNIKGVZvLMWvZo3TS5c1iEoY
SZwpmX88zJJ30VMnXqzTSdbvSdX1jXdhEd8iAgREqmnmH4o3kYYRyXCmU5iBArgn
AfkUR5Bi5RQzsyAB9cTmpuGg4ZuQK5b6MW9KmdttAuU2YC0ZwGHPy9CDwuROWaZ5
tI6PebnOLmi4D9/KggaPYrkdngEtyBbqYAtQXWESgQ66zauQhZ3LTA8POfpjXXjv
8OBH5BCQ+8zJo6HicpoQMIHrSrBQPYdVGKC6R5MqEwC7ISCMR4PvyyzvdXalAKIW
Ccfp9wFAO/7+nbWFS/Uly2BbwEN4cvnx3chGMfHdGRAulM+Eb5ZwKvPhVqjnsDcK
TR15NxSgsrlVZdOTodDHi+J3wMyPiVmYiRYExIEsquKLOlKzZgtoKE/icRxW7Mpv
l/U0sh9+Zedvvx7V53Ag+xlax5DHb/i1iCgy/n9PAWPXBDDGcZlE4cJzkatCiqa5
w0kejOmTnPw6aQQ7BFbV+8ezRaHZEKX1b3/+m1elyWmVGiNMikWuoLCTg/ICiBuJ
+JFHLGig+6tUw9kTCEr8PeDqq1oK0o2Tpl9dD/6V1Je5ZeNZKEzfKATjSN0Bl5PB
GfmCZeD8vKlcmmNgolD42DbnS120Cf79R4k4H84AN5Y0x4BBbIqCXn4bOyjf19nw
aPne8iMufY4Eb0kWrV9rUYkbZ4qCy5oHwX/7c8XmikcA4nkoxMKdWmWj3+ZS9aQR
LwQbgZu3jQ4rxML674/hZAqMDWmL0MynrcNP1gTc2YJr9oCCOAHbbwFmpt2DZFuL
2jxWggttx5uYIAO5mwt8/r3YygxwkpxNgtDSSo4W8nQapCMcK7p4cnD0kA61geP5
n80ipdJQHloo4tAYmyS342W3liaols5fCVV7YFISg+0C7Pm+1kulq+4ARilnJlUi
myQCbpOFo3hPybBCadfIZJcBdaeGjvX8keA18JLcv9d2FsuXr5dVdZw8r4NrvM+8
4Qkat8kl+TE+zpp3skT2A3WGedXaBrmIqKwdCYge6tREky5ozfoNMDlkk0REQN9A
I16ho8ln/xqYHzeAnb61+Wq4P9D8w1bQPcgcsQjXQ4vknG6Mtx4Q0GgXK+MEEhZZ
ea9yt1yqWlloK3vrFvdIXtrKu3c20tRzYfUI4g74EBp5I65rjTuzqK1mBnef3c+X
XoV4l9da/LX48oz7+lzh0thRmVKcGyuyqJ2kff+SRhAKdZp3ZGiXDxeWRnTM0Afr
N8Mjbzp5B8pu13ONRmxkQubWk4BZUK/6ZSEKiZB9M0mSx1bKjV5xEiLecltPmyOw
f/QqtxpBBqL492g1kmtPQbcKiRypjZk6rVNWz7vVuME7D0OvCxGAr8tXQF9/8VPG
d+WEGS2MGYgNe8MOJv83fIBWog+89vPNgZ6sRr82lcjcRGV+ihFZYnEwSa4b0Ia5
NTVuu97wSGlVLjJw3HQbTQ6KkTchpJErjTscioySUIVPTy4q/H7mUat7AnQCCrb7
Bx/aS2hn2ytnkCrOebwMD3HRkaxPcHneiNXzTOqIrZYrJPVKeuZjJhT0R/wIiFOm
N4Yx0222Q9QtdkIFfBKyVzIWieZijft8d+/qRkyJ3lsX/9JRZoqzUkOVOUzCxNRb
k1j0J3aW/oCEahywVy1foGDpGdUN29Z4NruuIo/GdIO4rGVYNMAkpHN077PQe3U4
lURY2uZM8x7v0JMayp39ZSmMzm9RTtNqDYjL17c6HtFGemEPxiJuSC80mquv4ZUT
Kela48/WvfHTmCY+StXs8Dts07pXI1ABKz9Hcb7zoXsmVy3oQxfD9BtH72qRVinl
V3Wu3Xq8xvwV8CK4AnUTadMiHGSiX2e9Yif/9vVNunV+4dglv8I5lFURWmIfFD0u
2+c5GEWBaLp3EKS0X1fKlj5UV/bv/mGDhY6X7hZxCxpHGqdEKQfewSuUeLF7dbjP
jnSdAMR/czPWZaPl7xf0v2koUraIjB6ZJa0VINv++XtRnOfs/VnnfZqM4KugNvgV
8GbP0PH0JtZ07GeY/X38Uf0gaMSzNdOuGW+M78M57taEsKbtv5ATnn5MrZmCbuho
zFITGrJunNh9A3FWEcWpifBbZB6nP4DSM7zObLFnB+qehh1tsD/0Q5A9/jQynaMM
25lN+aIrf2uCC/7NNPSfWkNGiOiMheBcYxfrK47OaBFEjxed1YgZF87+IMJhm9bG
8QnGzojlTIvhXA4fhZd3RarydMAo4UuMXMmYGU15XZCHK332xjJ0kOOidUfbmH8j
nGfNsF3HsiOe4m9rN9gLcgaZAgC3gd2eVLQolQQeEBd79VFgvj+yxEcNaGwHrO+5
gO5Rzrye5AL1youmzvQygURT5Bwz5GpVpcwFT/xk9zUac1uMiyoQfqUJyhx+fFGB
Zg2VTpwufRyV6nyt513GxXNWOb2qhCMCcPs0JYjDqLD2wLQZryOSzn1fScpyOilS
Y2mBreGCTIA2yqg+ez9RZtYmZloxmt50+nRpWqIQmnHtdpt8kUGfSq83G5Rb9bmq
rxRfrndDL6YoK/y1B3k0p6bBDyxD+I28LJRtPZGT3nRV8dk4mKdQOpdFv6vXuKLI
mv+iYTJfE+hSmFBZI5WqsOzIEAHsObsWEntgmOLobFAyqrbhvsMrqVW4WJ9L2a7s
yg6NBM7oSc8UVQ3rMKEMEeYnG3M2DaL4Jt89AJbbtJPpvhcSyOqCGh3RxiqizBgf
CnAn9tREUSoh5uC49U+rmrNpNmWyIVGS9c5BoskUo3QRiqSJ44WZnI+NtaipBOhP
HTg9ReZfhMyjhYXBzhukqq+tEXKD2JpkdUbEB1b+IYZhavo/orvEFbww5ewad68f
/sXUdsYlellTcAzIKuODMsodb30NtsFay09MleCUtYvtFkW8321nBuY7uVUY1Tyk
/72mOgT1MDKW/nKMFO0lwaRFJKcFranZF90hbda82lS0bhITeuqa9oRi3pZyZDsa
wTMm78cfjDH9j3WNAKnVgHP5GvEb6p76CkvPcAHkH/QcqQIqkYpzdl2lw90Bp9IT
oerLwhWyqJyr3Ajzjm6BzI8q9idwn++hrYNTof1asceuZRrnZCwQCr4isU28T+WJ
5bwx5SG7eKixktiokuDgrvjAvTDLAlfxYrMmc/3NBhVPVQtGMtub9IETwASyl8/y
I5wFUtVBY6k4k6cLxLNn7UeeqPwPLDAHmMRQzgCJlInDAj7uHP40dAUwnh7ly7xq
HpDAK3Xgm/ocIMSBCDOHQ9Kth7pV+G3M9X1ktQGoIX+f+m0FccCLZ2jGF1OZfFNq
mXCSw9AkQA9Lm/k0c00d4EKcjdO16wDQDeJduuJsOGwwVN7flwrGkLlqIqYwDup0
uDG9zI53YCYillpPMakYXQPNvFjH0uSHanvXjTDZq6Xj3yZ9QXQr+RYnAn5MQbTM
EyzPpuXZlfsoUq6+NGKKMtnx09SsMggssUh0kf5nF+PAoEiypkOtakDmOdHywJ58
NsnrVy2jHTrzVTTC4K+Yet4jD4NEP1INw48gtCwkqKMA1oy6e3pK43Do9YHwezmC
Z9u6bJvoCLZM1wPnACgiqQCUDQqYJ2egsK+RmW8PxdZQ3cHddmXrQjKuqMAfu+Ed
jnUrzGQspdhMH/SpUnVIARUqseQI5FtACJZqB6qQU4/Mm92RZHZBblHbbSXCtWrl
lmYESnUdtcjRm8iL1Nq64jVWDgy9a+yhTIQTFD0aWwpP2YkGVajvQmDEVtnny15R
dnUOws73+8iYqMN5Wjrh2uZ1r8rw3nqKnYFkMbyzH0IReE6JGLLgfIi3eH5Kp37n
JopYQLTGaf8a2ZuHNum8gl9gT+4lLmxEPXaP7Uz4psXGQmumuBzn8CDrQYVOYoq8
HttftouzJB9s+bdNVAjHooLXqsyknI0AMbAgTUD5BEUdiyWmed8cOsSAlYWBd5hl
MpoSd9YrpytNdXWHwM7JoOXdHSuwWq357zK4bhjX2JQdbIrO562unxwrUBHxfIj2
oU4yIopbRwG9yVNTaATnarkiHXkX2ZffwTWcOnH3cHdCo2UXmeKvy77ddNTM/cF5
2bo0FHwvGjTS4T3CFbZN33Q+TIcD7QeasDvnBKxikG02aLe1cczLjDHk9/D9h2iw
XsWUXNbfpGa0Nhl894hqczEwu7YL7bR1RrEwhWL1Gno5NVnckUiuyACfFE9q/FGw
cFvbwrNz4cbz9NcqnBeTbm+bEcV3x2bmlY1qsxva7PZ4Tu/u/jjLjWRAM2lLBfj2
oLwMNkP7fYBZfBQNmbVEO7MVORdQaKTYPO9ShQ+asWS/bLKSfzrofm9JhtETq4cP
YTH10WsIIxZ11JYouXZhnJIkPQTLpt5yvekLBawltZhP5jbzfatuH+7nqzHqnlQO
pdhL3Ys06PSbVLNQOOHEedq/ydi2P4zmrJctSGHvkdqu7ttsfU+9YO+AAAJpRky1
IxzW99xsAe4gMzT6RpkNz9XHqhMs5w6uga5e0xkc9uPmqZUNm6wXHbjRIXHNt6zv
XrdAcdyf/N8XoMWBJprJjY5h8PN0x3yhxwE2d4pXqLv9JgxCl5LZoo5vCqbvI7V9
sp04QQKxE0HkCnU7tD9yqkPMwjGKWkntrKtCjJnQ62UW43KSpNZkYC2murITBlV+
Hhg02vPss2aZiqAsma1mH/+BxIA7RpgFR5bXF3DneKvR7tyNOoQqqnnEGVDgKBXT
v0i/UbuKoo1YlatNyVVKY6d/GIQMTm8dnvfo361sMov3oVfAy5cM56xT4J0MzTDz
hCUyj4S2nD4K2A/T9P1Y9+o9OwzqLre7Chhao2bjVF1GVKmvJlPEKAcVpkOVHYzl
diwUpyFEoDdxvUjB6zkjIL5SBMqS8CJoiHnD9Lgn1pTo0imGeKZUpEIO1lz92O76
6+twEG9RQPUywdq/E1Fodp+3k5ZI5RWQeVBiRjsX4H2bEZcSFhj8Yu9YF2PtLJ3W
NFjeeiA6bRYuErUpOfJ4YEaL+1dRQqKt1YeBoxwvHL4mWvrcgp6JxGl50ixfFFRn
U7ECfjmYM3rEaMuDEzShRtlVK1rZdfAZnu5lrHivOxMy+wUafm44H/3aUguLt9JA
0lFs93X6yqie4eUNmNcdr6haubSiU/UvyNS+FPXDvpfelapvBdm1eUSB27hX23ke
Vzp0IFZi+OO2cTZX85GyNLfcg2XxT0wLmM9xNBpO4MQTbQwFA3439o44/DAa2nD8
XQGSUjq/0inF87JtiRkLPCpCoci5G91T7w4uNqIomW60fqlyko06M4xgRgJNPCst
ToyfwIMmsbQJa2MF7iKzqgPabwKltH0rIt2SdueVGUDvjfEEhAichCdFEQDNRJUB
LeQUwN7uRTiJnw7kCs4TLx9dklK5EIi1I14ihQZ3+pm6joD1o4BgdjDE5tgDuZp3
tQyqaqAONOd3qgY9QL+Na6MCssRWFV9ydhaqFjmP50lJHrJ0NJhDkqiT17FVrLWN
5s/vMpeQ2tSOamzmfnDz8thN6HUisLWo8scXwdz5jl+0Mgit1OLZoaFkxPHG3Zgo
O9C26AjcRvYV8a3nFUc/OPPB5p/bj5rLaSmdKjBpbf3ElSjhgrPDxRgrQhKr+JT7
RWIggWTLh4qmrKMm77mJOX3tDLcK+Bv82iBOsJWlRyZzYWqouxxmNLyhdmTMMssH
4c1tGfTEdLQG0QZ0StIOQ6VK/Ka81mEDjae77MopZyjs63FWyfawiGVMFADpc6kG
aLe3WNswlIDAOLOAAS/4qO8KhTT5Tf+AuJAipdIVbSMQFWMFDcNaIlhGqCsC3hiy
G1eJLKTNpskA/AJPu4OP3ljRQP1D5tIyofthdEr4/zPzySXXwuQyYRh7uVxp5Lha
Lzo34r1zE/xWcNpzt4tkldU9eeqrQFNdiCLq1kCWPufB/17iEuXRuUOFdHcUa0TN
5AQP+FAtVvyvEn5T/aOzxkhePwXnbL3O+d3Fp5vbCbH0/x5jD8Bv4+qKRNciJ4aa
9SEmak4FXPNOpG4fdMpEWfE6SUvdo4liph6DnGnnJ82mKU8t7ACUX+hvWj9wv+CE
hM2DO23O3HsJI0x0idMoWqYLn7Jn3M0pLFAWYMQku50Amg8YGc/nuLGHpSELdUcL
uIDPDY9ZOh/iCdI/aA/iGgkJssLyVpqSYMBlWQDafrS4iO5pTyrKaWCSHBo5dq3N
ZcN4ORCFTa3LFfRvdHLpLsgpjBRNqu/ZnQUWf+GNjgP9maau1uLVCRhZYCCJTlaN
/WkfnGE65teJNvcj1xYWH+64EsBGIA4XWQWyvm93cwVFjc+xxbfJbEFOeXMwkY8+
EWfjGn+BNT06jtqAD1A7FLV05bJOrgaqZhJ6O29dEBjlwzofhPq1akCzT/2mQ2vM
8QM3V68FL4ZtIgWhZKSSgHNbjnZtq5G1k1fqUMu9XrbpuorbUjifnYdq+EIdS/b6
cmZvtV2nbmmcs76N7eMw2R6Mk4u1KVCBH84DuW4oNsjKRWbyU4/Eh/OfKXHS4zUd
ikht7gZq1JLot+Jd5xkTCFsr3iL0Pf7kknMLwsqPDTL3M85S6j13rMQAnzPa/72z
NpGEFZ2EGtK6MtTB+egqXCuIfepE6Z/N0UxbXayLcR1wIej6m5+QNd8TzgqFpVN5
NRbwN5s3/ma1mttz+FdcAu9kNYKhq6W5Mh9TdvDigdpBcSMhZi3MpbhDfqEidP4G
lLLbxE/HXh/rt04hmarvsSzQd/vMYZlIN8deZZ/Xlby0+5XQo7Erz3ska9sglq6q
x6vHQfGBKR/3cdIxV7S+xB1u/dSeY11dpHhBREGGpLg7JIQbhGBzAvbEpcX6SweS
7keHia6+TzkxFcMWqg0/fHAImlePLJy8fuBANmbAJo4hCqNhUgk0Vba7HNATx3IV
ftZ6xdE3MgBgqNYAXEtQBopg74av8IeBGGhv+9wuW4SDogPT3nSODTBCUlDaltv4
/7qJHSIILm26NdibneTaHcdC7YNZtgzUOLMvrDVx/Rtsb9Ekn1T9LzaB+acN1qje
9Xj1eIAdXcDh2S4ns0iEDbzVhcC2KuOvPMmfAD7Y1zN3YScgxW2DjiciAh+18Jpm
QSc2PGx4Zc2hovu9nHduDKfjYq5FrexV/IDSNU8l0wyqcS2xowWZK/FeSBQcdW4b
ZS/0rlwerEgeca2UgoA5Tt33z5PFDQCevAEggq/7NTTGUJoMNRbLTIQqFo4iJubf
mSuw/spLqSOvyRdcB8bLXmAmZH8RE7NbCg9N3bMUtE8IHdDULOjLsENoyAzhBQ5b
vwCu4ZrYX5RrsoL68kG+S1kWoyx7otYLnmncyTeX3kj9cTt03YU1DlEkTkA3eTvP
LcDuEIJt+R9R0UNb0dCUrT18aXhesRYIre9boFoaqjuIANkdm6GcLoU5HXDihW+K
yRerNOqBWOxbsnxd4HPi5e4xx47CMYMR8IU119ufqJHXEueU5ONmXLtvymKVGvKa
NrRrd0/rwK8x/zWGTBgVrMhlBXxmAhGmlgxfQ5Weti7bFCS3KKOxRrG7zeBkNKGF
0czG9WHNdPoNmjZIDhJ1VUXYbcseDK2u+B77MnKBO2ezCJRmrrybZdtIFwAkmrq3
jKsxNzoVBpidqNLEWnpNdDkfAyij5tCYPq11jIirgQYqHpqMH6ExCguYDEnIYr4a
NbGVUDoFU/C6lSQMUQGU0oH9UEIRkUbnl+XMAfJksMNkbW7Jnrfvx5j/NetQmuum
BwunmVw5xy0d2iLgvoGyYdxjnfcbYD8l5Obeg38cEX+SRX2t7UtBYtkcSjh82g/E
I/SLI8RJhuiXSeIWVtogiG+p9TcFfR4PHyE10yIIJ4YDiDD+vfSh//v5MBVwjHnY
dqNI4te76Yu76zwKIlyHmXqS/R0P4/O3b4EH/k3i1Lshx1EttGdVBZS/iZo6mdlZ
4UDS2EiWmF6dK3UlQ6KDmiVnVO3qHuB6NT6QdRFbilkz4YD33BKn26vM6nBeP0hQ
52+aLg+nx27pWu5diTd4fa3DdCFscFSGv1hf0krfkhOifH4kxqeqwItJhtLzps5z
A6ZO+PJ5PKH2ycJ+M0K5GmGlSi6sbLcJNEXdqdTvrDbIGcc82DkRgIZB5DtT/CjN
U+n+Sm9BxTwssSdqdj1LsEa7QzF1cYYqmsGN2tpHc0Z+FHAK5Ycw48MXeMjFzARR
TKyYd6zh3VwsBki9GLu/SSpBuPpf8UIOggnHt3waEDs1DZAOA1NC6r5LgJFtzPYF
Nv/y8XRxNceaFzaEFKELUewX3OjQEwYBSvYpuXJUiUM/mCwXArJV65kpugCVjPKg
LuoISAoARHWawEzo7dm7sYCqRTc9izJpB2707fOTOQsCSnSJ/vgcUW6inFzIG5H2
frt50bJ1LPfG1CNl6U+HzMZC/N4YrX2VP4wWAkCS63ruhhgC/79hOdyVXVF8T9D6
xLkF9XV4/9C/XhilAbDWSmikGAj90UeTZUYQYuCz6+2rssRA+yqZvYn+NRc5YTKh
0WOrWbf+nzDhG7/1EJMHSYqIzgcXBsrrA45AkFauXjcUaKQ8GahxH0REPRoEynq5
zyGRHwjefWauSaCcVpzEWOgtgaKl7dxjJsowwYoEkqnc6zSwQoGLNyXgTXd3uceF
NfLDNGeQ+Em8bJV5cTpvOyY8RPFqCUuCEzPxj3zioaZzFFq6ICf/SLTdDcHXQita
SxiHNxSYdk76VLnigg/jLavppgif3qttqTIn87poamEhDJ9Y84Fy82KBXEbfADGq
Xfsn9DZt3n67Q6ApWhbfl50lE63WkHiIu4ZWJW69LVfmTGna9MicUy+/PVOTfY8P
JxDWOZ4qNcnw1b33YNfXauXLfQTSFaFWoNvXDMx/Qikbq5BnUnp+A+DxDkMpk+RC
y01w7eb0PeY9goq2Nj0jV3FqDL7slqFhHxsIoYcrmXn3mw6/XD7m0P3En7IbPPkN
DpaBQJ8l18QajDfUCupdXZiMFJXnMpMGSxC+WUh1gehzDPsRWSIsUlFtzf02Z0Z7
mXsfMHcHzOCu0VS7ORcop1ZOB6K3x9V21LmhUzrfHGSJGYPHCPSIPDwyPVkTFyUc
C1z9isRL/2fI2+4Ss6lv/ZFpJQsThxgdL41kWeLjqNZElnm66n2x/j1o797ZUJZP
2iPlVhK2jNJJ0AH6wuPhnvsx0PuuvW0rA9lspEsaSMfVcRFbzFK2xQLb7iyKG//0
xZ+J2i6u9y1XNsfHGbisd19j8PCG9KUMod2PUox9u0rLSTLcgZliASQdRXWpnJQB
5QriXVl+HuRkQoHEcb/sDWzGkVntkW6dtEExvGvqt8hu8LogTJqy9Hn+RZhimpWj
Q5ECmmE6otMhfOE6gVh+zSRqk+BtmkAFipBp3DeMXiQhRvcei0fzPUx4q0A69DTu
7AhiITW637XVC9LoP8D2RIqIkcrKwOb/kVO8rtZgDSWEsjsWHfS4IYY7oWlht4mG
mB06P4aKsLYGtBbBvQU9QU42bKdHyK0sJKsfIOeYTtpfD0N8HRlCym3vhheVmfs7
yazF0ERBbkQLjpInSfNy9G499ltqUtAkxDuQKVaO7g/xnmnwM5gacOEHdVa4FrZP
yC3rji0I9XCxXhnw4d8gGGkDS4mcShiw+Mp+mUNCPr8mzcmAqm+lXOAL5ebgpK3W
+T2uGxzV7xLSwpPnNGlZ5Na4Pdas1qSIu/Tj0DOO4gMCH8APAJy8Xdb/FLN1/gyI
EM1MvRlddsGf5xNYl/D+fsdyK5U4prRPw9aYbofRlfHDTNwSpbA2oKHDFtHi4uhx
+n+VwK5jC+H8EOyYdlQKQx2IOuxUIoc1LXYeKQcQ6hv8b+TVJLImAiRASxI6Ek3Z
c9gcpFrmM60WNYrr+TnIYe2Kq0unWBc1dflXB2D3DoakvZxk/ae9NPKnrJGkpjxA
rJORDTHkLRLyzhTR0GOScpozvGV0MVgcFoay0N6/q79xcW+EQGo2Rzb1Ijh8bAts
2b9RfLVgYwtyyBp+liahLRYjTXvtZMeq+hmY3dOlYzWm+sIveTyyb4ZmklY6rhQe
EuicaGklUIE2i5cP8/CrcOdmdLAf8zf3Ba1DoLLXkFbCc2hCaVE4ZbIwpzlT2T3B
Cj156YwtMItr/bngQV2FFKwb9DlT2EsJQUUifBdIICJSSGlKy/9SF7I2kG+0d418
t3G7meSUWJqkcRVqUCW8DiRQ6PXqWBmv8VbyONb2EWsdX/D32jhX0R/zUt+EqFUL
KcelQ06oezl+tDG7iIDK91be8RLqNnpB9pMKyl4yx/fdm5ipw7kUYQ3VjlN1TquP
ZeGSOpS2dJW62nbwXbl0yWGtnJ6pSOgXy9XaMBYeKstqRUOCqThrI1Bq1EROpLRe
/DRCDj+HzKYdsi6gI1KwdkVP+NIPOWh6Epxlke5RUkfoaoMtzE9SroblzyrpX5WW
aE+LAS7GtHTGf7J0thKuO/TZuV98Z9pPPwz+b5wt4QLHMys6uHC2s+Flg9v+aoZj
v9uc/3icIlVJcj+AVTxZwcSP4R/+tYIZHrZkqti8FqLYmttGy2P1f0zHrMUnt9KE
eIRtxsOiWGPBY7yMjw7puDMPE7CtybYSS4FB/f4aMWvuPQ9CcvnZR8kYvix+9hZo
98h/GEqn6IrmC4x4VPBNYFCyaVIILBxwhgAuJNDHx8+T56SCVi9V2M+8WTl1Qrjn
ntFAm3SLEn766kHNFw51QwU3ZCjzKgPvJip94LjGx0L8TyMY9ZrhpP4yLCURJNS7
t6mMwTfho984oWNQebY2pGCTTjtTtZniKvqDkvef2yWkK6xcxTb5SGtGJKsDSeSO
jA/vPZnQI3O5WO8wDILz7teaD882SF4Ojyu6Gzr7XB2ZnK0efGoiMre9deugBcwF
JtTSW81g4U/6n4WC41Q+qY+pV+Tum3RiFwhIFWeAcKmo23TvgNNoRkG9Qiyrpyrc
ppwEqj8dyYR4R7A2UbP3LJl8sJNFy19uSfLE37XxSkfdd1Vme69uiSBuqSPSH5Km
Gz0jz52J4PC0fsicXF3BtO+7iODrAwAt2pD0RlYXcw3jmN5qQBM62Kwbg/diwDtk
1HvH+NXGdQ9/z4ucn5BUWlDy8bR+mxDDZuehSE/3n3dQDSGGqNPy4e1y2rRBcqiz
CAuBpGVRBWjA0Nd7KcOpXGPGMdBAnxgMvMEYYfv5d7XNW0wy+4rGeCRngkzx2ULt
WZbvpWaTIZBiA7iumQJD952S3wsPVClO4lqqTuE7Q7vrexQp9Vl6Bbpf2Bo7bQD5
RV2hPqvc88ewIrfqEqNj8c/tVveZie2eOQwgV3iTkRbK6SAZ2R9AxVqkRErKWO9h
DkRbqFnU1s/hT0X5R2cvArG5HNhLLy6G05Fo8OaWFKOWj91cWqSqGzqBa689pnf2
RqTCvhiTjzpESv4iGQqlP6l341IxOo93j6K8jBEvUiI5YS6qV3r0ya0/EiyfV7Z6
+GcULqnxQOzC1YJz88SJRNodkgDZpJBSZu7vx2abCGTHDLKt9+RlBJi0XwGkaLNc
P9xSlnUrkb3NRPVTyIaPGokak2ot6PC5r+cqC2qp+i/WIFOd/zeCjHcQbumcX9X4
0Z0ofLEI011EXbwDDsZNQTiWaXtTYmjSLouxb1KDBSDvoJfB5rn0lO08ZzOrUgE3
EnLp+4v/r03gEMAEPkp59NmCdUaTyxOTX9BXJ9nvxe/M+7tfDwNnOY+A93h2vifS
lvmwHibgopgerdFANzDU63gkINituyKLAANRaJQ0gQ3dDDFz33vlHkoOcaaSKCil
DtmHbr3cIx1Dg0xjbJcz05kEzrquuErprwI5IA94cGY6X7bTQB2vUFi6itRhQfaf
i2vQ/m+F2TvNHZVwSgmLIupghtspo86HHHLWBKS/zsUaND3YKuYGYVmVUsV1QC3g
03FGUYAEqapkjvZN0nsE6i+0QJ90h4ztvO7rSrb2UGKE5zR2zxW8d04+LJX7lbuL
ZTO6Dsc+sY9Tc22+EqOpAKaJ+bS/96m+lLbgo5IT89KjNK1Fgcb0XmhAJRspElvX
Qf6L/eOAA+m+jORJ7Op9h+P7jg5rWiBz9V+UFXK9RjHu9dJC7/I2tRnC4jU3a+j4
qXWfGTtUNf0B09cNMMl/DZqieMmB6X7dDR3wvrg9uKjG/GzQM8yzER6HCAo09qKM
xc9xle5eukZ5YfvN+CJP25aqULph+oLaaeNXfMMjUlF0EAzJUK5WFtcJEkoCJfs+
Kmm09TzpktbJOFijO7iPSM3cx/uwBBskbeCj5Fypwl3ma2R2MW/VRIHUTZZoBq1S
RykW2LwrWja8cHut0E/eUNXhtfqfOibS4UPwYEnI+pgjCNCTxP1tKxqQqVVn0rrZ
7PD06lWfAJf1SB05dteUTAjT3mOhKD8znC3rL1Kah4lNo4rcNna6H33ZaTVBEXl7
ACcnoE70o2RWtvqNX0qO3NdOMbU0CihB6JexDlZeM2A+ZUCu4CpR/EqbmNCJSHn2
Xcy869uvyY+mnikhxd6mjmgL5GFf7AWySM5fmqTPBA2JDom6hJWX8rzGnxWaWYA6
ZpEWI3S5NH/kSYDEY2ZaNWFPq8oa1xZdM8JqJ5w7jOz1ZztSISZIdPd2Iv1EslZL
xCEo/iPkA/hWkXHqPnOgaob/uibLdjGrAYvYeAscKgF0eGfhxRrGp3+b9pwOznTL
xbsqyqpG2gb9uNjkNAdf3V0/b+531Qbxzer7CTDLoVtV64zXSanwzatgYiyZdMoa
FjPXRv3Vf83k6SB8BbN5KKpkHH2eH/KH+nMqKbq5tKM8zPzKWL6/hl1DaB8YoM2K
TGxCT6jKrn3T1TGA2UMJ9n+4Sb3wCm7FEMpq4viQrcxmNJ3D6dv2+atJOl/wq05k
4+QW0flPk494aZJ8gJOTm0Z2I0y6lljGL/wBBEnCEbwsHlkfvo82fW9Cz91EP+Fj
yrwdYrmTFF7vpanvxZm6Zj+d2SbBn5+PFGMToKyWkVyQXI9jfG4mjWoKX2geoADR
lUW/z865LGYiRrJavrskvJ+oFx8WE/b5sUjQp5G26aO22xcisZmsQ4tT205YGS2N
3dWKnBjW7Ld/nckCeiFH55tGBOoCRCZM+50SN96WokYCEUgDafSOrA2+zDIeRttd
Ov5FMgvqYsRSbTH2z+39ht2duVz1WVk6J7jtvbuu9TnX6KM0kN844nPXUmjHOrfQ
cdUk7xk9Q8OX8Vg4Go3lSzLBUgaULak8lKRySQFZ/qLiIxcTym0xCnT1hvxFjjE0
NLgfheIig4BRwMtpCBB5py3E0RZdcdHZcFdQlhsldSgRVB7qndKimcJdw1WM0oL3
nOI2elsEByCywTp9kA2NSadW2sOaYBXQHRd1r8ji/1bktndLEb2Wa5LsT0Z6Gzd6
rF2AD33U4sI68L20YWYZf52h+C0lr65GwnWU5s7UnvsAo87M0qDxh4yemyVJGsrk
pNZsqHJ4wLczjHS1yQowr1MetAhUGUO9GE5+3PD08xz9rHUe+rLay7e9D6kb0O1I
ketC717ZyfKLivh5EzFGQ4ea+S+K00E/9SxAaoH6U2T13G93RAHx1FxPHSRAIekL
wsPSyGBXrpPRgQRIXMA9CuJ78PCnWPgcYkYqExkCQ8aNLvOwt37zJOLFktmmWpXG
aFfPbp75S+8h0083ZmgRGyFnTNHrJhxVlMp1A9TGZHhf1A9LP5HXRLg9gdPi05da
YOAhxM7eig5fBa4rtHmIWFZvQLWxeg10TFCAVm5hTWWgWqkeAsuN62crldEOunXx
xMGBkBMU1VK0Ul1CECC7gNBc0cxefV+vA4vJEmDqq36A5GOwmb3HD5hcbMgcw9n4
7NMyMB2DifEv6yfjISE4yLVjzVroHAkW17Zoic0hoewwfrBir7+TrJpSixxnqIaN
3mIbR7H5OCyYPJeJFuwbmqmXcwGTmpllqtCTpMCWY5XYNyh7PwzcJaRO+Gt/ubjD
y7EZCtdp4beDtciC4qSevXR+tN5eZhNW8XNJp0Gm64eGwdYAzRBaLXdnGYfLLvLt
Rx5AUY769Lspg2Y/aWVhLIHjXr0dxK8JP6j0yLBQud6KBenhUtP3XNW0M6sg8mEY
TizVWKdJhkcAG044XWj0GJG1FMbiYqYI/xYJ8xwiGVlzn+5MquOk2iGqUWlmwZwW
W1aPUYGYrZzpVLJCkcIscPWHkTPAn+AStJHPPcAcWGtGLy8r18v94b65JVFlJUbQ
DuqvaYcSrqiFPS5jfO20S0WxPTz1sgXPFDyaZokFHXHbW3yLuPEJPLnJHIxxEZe+
xGSKvYRWhu2nhQaLEEbtoKtmuLotUUHIPu3ChpiUINF3rrr1DLNm/raPIPhkLVJG
aEJ+in4FejqOtXI0Udjkuy5sJfN66C3qYzpKk2k4R/ff7MXBSkBme7fj2vnhNEXV
W5WehrjbN2/pfi74KC0ByERg5VtGwF0rLDNy4Wj3OBaEkcCDSrcvK6BJ0lcRS+ua
JbGL/5u/V4N/x0X1LB8UsBojIPGBa7qpVSlKP1Q6NulmGsD6v646aGUFKWdQkirW
kkNaxHpT4/lKW4CvxqvY3fJkld6QhDWRMUeD1fVy2FoiAxGG+4vL2+/A/0A9Lr8l
MAAH/dmIulEMKh8tdsxVoycTh4aKlXf5HaucmpgBZleOf3E79wKxP3NN26JNe8aH
ptV9SAM3PBA5ysLhcp2o7OJc+/juWo5/WNze1Wz+yRcCidHrF0Ks2d6j+AVWkpOH
NaGtwNqQFSZDvIjcq8teMkqPB3g8aF59+wN1SKOcTBRKnbqgdlww9C0QcyhGSNhY
62AXzrego7Q0TmAZ0zUYZ7jlCteh7YOq7SCOFX3Gt8mRW/7Zj8+Tg6GHCcXU8koh
xLaCqMNLR9M3q23NX/Pe/TzQ/8ns+X62rWMe1zWzvoCu84W84rWBk1l6MmSpUJPw
8ulKBDq0EJxcbmDM9rsQJpH2jx66KglaMSgINBZP7AIaTiBzA+V9NifLpbGdecNh
d3FnByrhGALKLnCqhEY+qNDuK4lB76V1IQLQBlQnKhP6J2mO/JOGNgalcdrRv0ze
BmKIfwsSsjFIB2UNSWAXobHq90bHNrpQZ+7oCUDBQ8DCX3DqWG18ZAKG2KMsR3qX
pEJuRRJAot+pBrfhQH09xlZ0VpkHPrWPOmgbSvtNKzl8wE9WM2JLazk8O06WGzRa
KTSZoa55MQw5hGVrQKqn/SLoo16ZElDjutGa9IcqITfEZOjdxZKdK3v1BwzR8OOY
KAw4Eu0u9VkoGmCJ9kAcWPJJ/E/dBe9TKUZI58bJ11l8EoyTMzW14uSvOSCrSE+l
nDdTXp6+QtzV2UK3QL8vqWJDFALkfkw/KzGMsVTq+CDdIoiX6sOIs8hDnBcQk/lu
IPKA0pFodEEdUrJjzWPdUKCZi9b5alvfVDHlD42e8m9S8wNvJrcMwM3ZhJGhZc/A
uOXUftqwst1NTCn/ll75cJIsZp5npjN/l2O7ARf3zlDTZaMajDD7znXQOZT5cs+6
umTu6xsmU28w79G+4xafyZEVF1P3EIS5+9uOU0Dy64Zw3IdZ7QSnoNpnpIxBG8X9
qbFjy0b6hRcNgISi9a2BlNrXZj4to1Kp5fptCH08qNid4uneK8PmlFo4LtavEnX3
WsoJbduaLoOMRbCWNgoN9yaUd3PaXd2LGf82K9hbMF1VndQjfInniQ49xIlekV5y
RI5Phg0bQxtZkMI1lzMLm1D+Tmn+wYY3cc3SUwide4Xp1JwBt9bHanzcQXu4TC5F
qtvTLAmolIKGHrijcIwQTUDzQkEMgg86iBcuyl+hKkszNlfPPfmjHJdSp6kd3fTl
vZ9Ty9oCu1RkrzTFrDciMnKMVvZPfXcuEMOu8FIxr+bHVu3ih33KPIm8AXytOYZP
htDSeSYLkQpPvzPmbw6FcAe+MZZXDFvOZZBlab13AQ0jMd69uYzInAbXW3XWJdK8
bnI4i/l15baFN9h2+fCdVb7t5hDSqXmLtbO32Mh0FcApTIKZsJkolKnh4j5EnBMO
QmWoR72HOSbz08cz3iUdKdxtk9hXeG0pYS+IVkhIrskFWh0Jf2bWQ/Elf8UmYZaC
q/pHlVTOCZLTSIeMg/MPAKdH4rOgVuOGHmi5TAL1gxDBZv3iOaxAspxS8ZoprUZW
OE4Xw5KRwDnYdCrArcDgj6HLcfoZsbE2vp8I2V8vbi2/goVBG4d+z3/pvTY7WmdJ
yXyCSdPwSjgvvoQgVoXVQ0or2t986k2RAXTBCMH7YkWgzSxEtJmPCqlc2fYb/CbI
6qIp3CqFizgBBHw9TcRXd8gaBHTQerOvDWrNtfkGGIWyTs2y8xs7udsfRIRqW+3M
ydvEubB5Gf8/Kqsg9UhUEH2PV4xtO1HnT5v0yfQpx2tsA+0lqVdDNc2pZXLEfV6s
m1ui9XZfdZNQIBOKrqcA8wN/YzRPC2cDDmlpU/zZ746gvLZ/93Hc+NoIzz1NI8XG
+zZMRZLYydwGt3KJtf53cTDBdi399TXW8YkncQdWPCv3eKHA3tYP5LWM8xm1XJFx
YFDH5jdnnCHPz75d/8U29WkycoqAdtVJgLM8LtThRYjR6VsQSn5D1HtLKLs3Fb4r
8BOvEfeDyBPjcOHK7ImnvyBgR1vWW7kVRptJYBJntJPF/0UC3qA1voYe6SxHPB+g
SRwDZEFGBy9rnntiLtIcwVAGAAGk5hrrG6RhPgFXAObta4seir+0IgwyX92W/a5R
Sk2Z7LyDzoZPcP8N7ZT/0HOznNTeooIpaQO7Aa3EUcn0wEMNoE6D/kCZ2zZiV1W2
S1qgM00OE1LlolS4SObXbACspOSdW1ZmwWqmtOisS3o0pOoDFVGvMf/HpX+9zPNe
+VBiokt+AqGdcF/8Y/bymfSIjEEfLDxfGwmRYAwzvYJXtx/75KoSd/Y1YaLrAWfJ
2nCKYEZqVSUNxMhgIaFLAG8iTyyCEISQ4eByJ9ccrMcSbPSDX+urPD0yToHRegyF
ohXim4UPWWa3L4qlYLnEj+KbjneLErx/NVFz59zAZr+eCfKq+GjyidqhMyHAO/sg
ZXcWYetcQM9u10x/IQyxyGE6oZXZpPm7MdgFYvm2DD0F2uWdrpOF1ZhtjTMOn8Td
32wKZJNTt/1HQEVC7tUfvp1l384djcAT4SNw/tlgLjDBx3a60NmCJ9RJ/quFwZpR
K0II5VPe0ubPrI254JeRnz+sS3Sj0CCaa8jHPigRQ0gUFd+9mJOWmQDSgT8o/GVp
sBS7D+HsIrOQ96THDF3XvG27yTG9OA0dwlaA1cxMhVayVvgYWqY132C46T1aJ0ZQ
9CHDn8+7aqa2uO1ejybFim3ZRapP4DkS2sn/kGMemASNK8PKA2z4cYGkHXNvrcyK
TiS9AccCQXWp08Ff+bbq25KwVaOA8hi5Pi69hG+UZhHNtT5lT2T7xKqPec8OyIxc
CE8EOLsG7HOYKnKbdcWdRNQCstdSfynBPBGWvrW9t9HEtKsrqes3Kkjo37p6vEn4
qzwsHTGrr3v+7bQxhOrW/CpFLmiCL3WV4+SBPjxlYxzAaHrcqglzefqDK5UfF+D0
UeFjLCZU4IiZQ90cWrGHFcx1Avrzb1ZH5Upn6w0Fp/9F5SIka2lwEKUa1VObz8Yw
wwmnsYW1lBpuImlYxSMyah7CPvUlWT5GoZXmNKy3mOm6kqJzdlZZ5a411N/9gIVn
bYSg/e286PfNuCeEG1SmKcZSMM9Fxoqkbb/WqKFxFpYIm9rEdkm+aXlr8sDoajAH
5wC2lel4eB6+CetHGfu1MBOoHRM3JlMNnNehzBgrZCFqzhqPZlCsSyIlCbZY0T6l
Queuw6iAxKxlZwktnNM1VYeOJ6PhPMrWCXa9P+KYn0Gu0+2IF8aY1JYRywFHvHst
+OLbw6KJE5AfzJIioh5/IbLdgdb7XfkZQDXtFiF38UpPhOHr2ErhrNdZTvfBoMQQ
YpVyXIb8GAvHcsnxvF8I0fJ6cL/kLPh1ROJR0a9X4Im7KEo/Qu+LJhv/I/GTDe/Y
5pQMpHvFAhxJsonQeIz2K40biMzy9P2HDyX4YqSmRbsIiAaq4ph4QDCb5q/6Xl4y
Tt/FPaL/sVpvwpvtinvJuKxWBxHTTMtOMuRJa10bLHuTJftWqZ0TmgGtCVsmr+ul
1LSInO8iebyE16Esl+Lm5opNwAfkEtG+bWmAgSek8LxfZrQEuHjAPWnJa2KVd2df
Wznc4C7A4baIgppOfItie3/vWWnTGTi/MUMzP422j7WIY68LghTJ1LSpz8+kA1nM
4wbJCZKQ0ydj4N/P3rlZvJ+3Dz7d7exXPzkVG/5zQwKCGTxMFLMMRF0qtJqngnb+
EdNeL8MMhw+Zn0D/bfzmskM1kvbmEb1oMcfcudW5KPzJsDC9saBb46skw02HWORJ
PIE0c5cqmfOZQh07Zyrp+Z8kzRshEx22q7saguano5VKoPHxHjouRpUCXNePbIMa
bQ6Vy2QdiPPOcWR6JsZkeaN8CyrEiMnv2EmmvfiGA+OtIF2UYY7Wgrp+yTSuqapY
OM38kclC4kHxsQXfTnge7Rgbr0h2Gp9n0UutFV1rGOAWTU/MMT3tTrADXNpDRDx9
SioWVViDoQ2yZAIHxEUccXz+JscJJwP3X04H7gblL3D0KUMaPxvmgCZgVhYSE2jR
RSfmV4dBypzFMi94QXWcQWyxewnqFs0Q7ejNOpUuvpin7i1lp/IYJpj5t3nXDBQq
fpxy6wH6ey9biAsEW5Nqas7ej9adBf9N1CxvYQTidQLYoXz7KM14iOoomHxg+PLV
JQycltv/NnTwFotdRfAwkinkRx2Owm2/oL8pMpw7i5wNPrtObq47BpqxvGfT7hBG
X0TliBzI9Um4a176QXySIeE2EA3SPsc2G77dy15J+0fUCMXESIoQwS1tb8kDqEJD
Kvzy2PkjZQLr2baUcpV00U2bkLD2Bma5kdIAZ8N3BiQysXSye/gRXfLJQZE4sGmt
pJkJ8OBBpwj0Ro6dxlzLGETo9K4vsdlIXbJ4xIhdPxkNWveCzccxGR+sOFYmxxxV
KWudC44fgno/JtOgrM5a9dWg3D7msv0XxjdRXaIngcY04R4okfrGr8dy/BkFjgXK
jKq7+yiWaIU6SMa2uSzqp8WhAKpPC/z/tRFqndfwey2kpEJfOBfATWHHiXXBMLCh
kM47h9teFcHrsiVw5fZizdKNn/BOnw0XDD9S0ayrFnD4cMSAeL+tOnZKLNIKrLeD
Da3LrZI8qdE0ko4e2k3LWOWfZoj6q9OyyNyt/3R+xGEmD21jYIm+Ud+RW7mV3Mmm
YQXPIqBt6nnVxmNcNQSNKooAUztpvSg9npwYq5JT567SpwsvktHammTE5muh+Lg4
+OS4Lujm9JT/PIrY3LL0EWUdK8IDjdqX/Cjnkh7rOOmxnRkQ12XtadQ5a9PqLd0m
s7yPQZDUuWK95mGXR5lioOdwcQmZCOrOULGBCPg5EpqfQihKt8lJCco7DxgFcf1C
wVYT3ZHcjbaImbPT8Tsj7SvcZBcIfQ+sxDeG53Uh6nXexu1BA5R7CRnWnEMhSiTs
g26IXlDywSPb5e7JvCVlRrDpPbXksCbU2+udNhisWMVniJhjWlD6mE7GZrLKv9PV
cLgEBoo1oVHV6ZVtTC/FT+HgjR9IwuisXjPTc7i847+hPmc71aOQhI659nb9f84t
K0uK13TB+5INKxNppxGkb2xUi1XGE4n8KpMYBtOFDtn5omPKVOVmYkzymd4HKpqY
9Z5oS0DcsvL9Fobd9JyT7v8XUqCIK6Uv4w1xoDfOBu4fyv+sfPjySszDrOHKg7Uz
4PdqasKzsG/wjAO4GmaY6EM/hGiz7GHw6tOyWOibtT2sKyv7ZWr6lGZ3D6cnL8fl
IfsVYqpEfgwTByOw5mbQbvVM3rbhtUc0Rj+koPoZSchQ9xut71fDDk9+Bw+dILjh
mJhnutiPevuYXc67UKsmhy+bI9rD7joO2p87wr2yzZqs28Dqv2j702CqhkST/o5B
4NsJ6Uohw2nEPy95al4oHV4zqbCB0eai/6EIQi+vSEW5QV5KyaeAtMadscge3K/1
QYpES20OZptW0vvfqjsDuoazKC4BKXnJvktbx/BKrGaRQzyWebNtQs0aWz6MCpli
C9ySwh8OZEzyc5pChrTqBZHiRuTs5FJxOZ556nrvU2V1PNXjp7b/pWQP41PXXOoV
xRZ5oT/bUQKDeHK76ju6EHk7ZxX73PPviXKM1PgE2g4BXaXAQDvS4487Nhmo0voR
fHZxgOCrfCVii8JwskYhN/e6BoCokaW/6VR9J0JzQzQapbd+wLV8whEUXsDDm1ty
tGu13efapcmligrKPHJ4QptVdrg88n5f7Cgh+1DesQYNV2RK9VZa966tmi4Ny4s4
XFbpuWl4i4FwgaQXqwl2EgfV/oxUikBSdagHW2AOCsT6P1/YO5rQ7HknhDXyYWNT
sCHNy/CkVRW9JVJqMMJYf6/kTr8KNszcr+ek6Jy91RA1y95iYf6vEQ2b9uuO05aI
6mVfk3LSljYAPp9HxSSV4fkM9fDTkwz5k8EWgmn3Gy2oNaHNeTMIsvWxbxbHEOuh
XGfWQ/jzMvLIjZdSJl0Mr6NRJ4ARrhIQpMfGjI9yMSBm9y4NoP3dsJ1vOrFUZhcl
RxWfzDH1Oc0n8ukeOsAvXrcRTqrpk03JJgUnkMBEmy7ROsRFAI9YeDgctHSLyFTX
3DK8MukEajN8TGzQwvmCout9VLsd8W+M6SqfAAbPZrLYnybxzThv3ZtZ5J2EJfCw
ImMwvqstbIfxpngDeUgOzg620fo2VFtUSiWu9yJigyheNL+yQf81ugjWYxxi8hHU
ZRKdFtNiFaYrsKAYD87TF12rskUJf3XEB+teVGpU0NYjvx0yAB43HAtOCU+PUJgz
2N0NmoJ84f5bwJKcW2HFbguf0MOMiVXM+FDzogkBNONy2jlVI5w2lvpNlG5KtNpV
uMJF0M6DLUR4LZNz8nc5lJNtxz4psdqRU83fcmeszddp5WuTFPyBQ6aye+zWvTep
nff50MTeAsgX7BTLXzSfegylyL+XoZvGQ7+RJXbwEytllrNmm7ho9qEKvCotbuHK
VAjNmcaU68C/iCOq5MsfmXn2xNhlSV8QDSaFz95L4Qe/pOyVR6WtrSVFaOdjVXSm
dv0AskdS2MybVPzNLFdtr77v1pZIXeB+Ngzx3Sf4sjKpUl+W+e1pYf5XWnBt+yjX
OtcL/KiVXOR7esrHUzj7YLLLWvckpYn7eGRjmi6kRq/elbK/gLxNkKs5laK8rfEL
tVXmKZpRQv6jUhiFspn8aTvW/0+ByHQ3k3P/9fJZ2sJJQlurTyl/l1X15YoUZp62
pelYwteLv7emNuB9t8DCr/zXIJzZqEWhrtKLgqwtmYR4djLz5LKBuA1nqrd6t94l
9cewSh7k5mRXD4mjfay96WxzhYkKXAE7IDd9LVHbcJGHW4MIfZMDGD+3C5p/t/vU
GYeKGMoXUyS0AeEz7o2wKxGnyGUcJoYx9hkejWGkb5csU+YoTF43IIF3VEl6RQmO
rBTdCeakhAnNc3Hb6xhvC1yrDXdqT9BnHA/NvXHzDegHVrF4PsKYkeIQjN3d1V8t
SqQB0Za5dHz2R9fcka/71SM5arY0NuBZ2q3SaSYgFXBth65QQwtXHegdxjkQo1vw
ZtA/B3EsXNgP7sqTh6P6yuX1z3cnxxie3gdnJt1SHOWGAjytgwAOCrF8LLbh6Z3x
SF70tiLqNs4yi5tVZFOPILONl9xAExxG/ZAMjhZbY5eD3hrPj7RPNN5ajKePqZ6k
4QdmWoKu7/Q5x0F1oXu2ShIPU5+pzGJh/Jn8uDZYZzCPydnRAr2femFEPg6J5E25
9m9DiNZv7+7MOy8qLvZmAkt1yClHwuHzDLNeUu1Ffskrz1Ez7F3tOAgJLiiDsNKB
S4F6LiYXWxANMAPdWRxWtaK5mHr6ZD1lFjb3D5byPxRMKaaEaO9VsbWL/RJTkqQs
1UJTrIK8o7gBREFwj0X5NQmZtVw6VpXdT1+Z9eQB0R2qzm+DN5Gs3D+ruHNWiJsz
L5REtZ1F39eQWX7LwJX5s+L4CAMwqZV2IwpTgisU33a2wslBJfY8lWCBjPFkoTJx
BhO66WExWh1xcNbFZCSPOBP8a8b0PLwDJB1pCDvM2Yp2VMuxt8wVk7YqipwOpEIC
GlUyxR+cFWfW20ZA6KOGl869zO2ZvjI6xITdIDuPFVgygeYeNzkwLvoRZj9rrwkz
DOx24DMObGf39c7q1NRB369gSVcTtjDRyEQuhwK5ay2yf+WuAG1Z4wj5pTi88rHH
m/2eMCAYBvu34McD+3KN/vBSOztrDhVXNqRH3UMsZdyowjl+qZ/RBy+w2EsJIUFe
QOO02BsCz9/KlbDfSWAeV6kW1BTf4pXJjvqnoDFxT193qLpjW/gibdTW3S6WTz0x
uN9hhfvqm+ulW15rTEPOy6L+XXAYRE9C3RCtV4H3RKbpxdU4YzhFZxMej6XPosv0
aR1Q7bBN/KmLIosuVEK4fENU7XebEXjiVuNOA2NaVQp2AzoChI2jGEWHgH99YoVp
yLKYJ0nP3g/6aoAVtRoTMYPZlHcUfWs61QPzv6CfTW8p8RIfDnny+v8FT3S7VO8U
eiGQ3hNt/5RUSZEu4dFWTYKhlhIgXWzw0PBwrptuRqbMyeTvQj6+EmrTbasr1G/O
FMmf2fIc6QX1rHDriebNjl7STtoYljBK5PxBOScKiwb6mEfh7xWLoH0fJDEkY8xe
wlIOQYUKIOR3KSJmA7eMCu8KIu36Qgkjh350426ury5lGmv9f5JJUSa8As6frrNR
ZIpUt0SkCJp2nMFOABWpbqx6NQwYabunjwYp3G4e1HaDMpUO4REgtsPRptn40BdJ
WrzGEeLWebfNLdPvD3uQkN4GM/e9VQe8dnJalEoWhweDj8JPCErhKwaIfSrPz1Yi
hMkFiSIokcY8HMSpGfDYGo9TV3M2btWorPQa1uxJwlSgohul7wX98OBqUStNHX+F
zqrRZ9earzvQcFBC8NZZ0M4XX419IEQLUj88fkWt+7lCMMiU7rL+dCOLRyUvrS5W
A7G9kFUNuKFzy+dRRSQWy4dDAs8ThgnA4OVwfjXdXUHAOkNnWr62d2RTM22vkLcz
w63q0MjLc54kB5BQRqBvmU1ay+nlNvuB+IxgFzQ491WlPaPv9EWB8Z+CsdYk93z4
wastJj/oYcnOW9CrW0jTGc1GqOM7ie2JdFxG0vy2B3Y5ioeLRIwhcmovQuXB3Fwn
UMKTmTqguR9h5CDvKFcGD9811cvJdg4Jm3Pe3X8P23XfPunCNX2JbrN/QOrPktXC
NVpgXjnDRS2WOzLTIx1d9VPcwRH4Cgnz/E34dmgYFuzYXtjFnEJBHPm2DWOgxmkH
7ywn/coW/etKRUYUEV00cjaF99Ew6uDwV6VvI4ruH08j14ktvxhn1halBANfwVGD
5RUu+NQ8Zo0IONUVx1SBleTNbQCgoASFP23fNveMjiRYaxA+AKe4zv39GkU3k1XN
5XMIFOFy7a7z0fMsVx/5/Bs+n6a3IexEL3/g1a3FEHW9C29hohuQ2l6k0zhqZqXT
+K2N4b4B+zloT68Se9va5hnE4OF7FMIKoi2L+UeBAhfNfiSxMKZ7BnbHtaaAEAhJ
CMx1ZEe4vUztPUcKAuendh/Zc9+VM+H9fDZBYg6SgcFX6bZbzKoWd6GgAC1lI2sP
ajGskzMIWGEUh84wjhQfw46EYyiEUicTzT3CtC5vr/6Ju5bZVJZTLHgGCFZgfT0g
lGDNOj5Ub7crB6E9a4AvtyUvSj0mlh6RaRUKGI3pBuBRTCsdz/mPLJXxqjDQXt1d
JGsdYkrXS40VPhIDxPGHpaMdITtYyVXQ90Kg8II/bBF8uo5Ja8dYiWUQDS0xKv+m
czwjfNWjtVimarYRC02kK+Zn7uoDs3k0Zmg3EXO2U7xXS2aOyCaw2qj9ZQ5kIbkv
2w2+4GZn9Zse/rbL6iDN4Q2uUzKJKXCmVxwrP3TYryCiBAWNYTKgSacZxve18A+p
Id4NclUqdytjDZ7k7xNkDtn23Tv5m0uaGUwzZm4uKEBmcabE2U+nLmtG1nNme1QF
aVY/JpHhC3eAACeGL8LVniqlVFMt74mb5rYbAUiSGe2ehLU3WNGH5n7qWPK2ZFAt
cYa6ZID2y+QpwTgoWni76h+oXSCDEEW1Z1Wu6kAAVioTRoLi65A5DeAxNA9dNcCp
Tw5WwsYEo+0hdpU4G1tU+4TxZiNqauexdmKxVOVHktYPCC+Yy9RtNX7nb3QJXr3e
NKcgINxH54qEdEppHhHxq5PEG6Nr7t+Drem/wGC3b1Lix0WZL/7749siZTSoJhX/
64sFePRRevFIIvz0ZlBuPlu8SUph20Vp7RM4EW3Z59ucZmROJv88mVF1AZsAEKQ2
NuynSmpCwoymwb1BNhmWVGxc9lBmXnV9dPCOF6puXzLojF+BV0kaey7+s27wIGBo
2UolKyfaICkWocLzOY25PByWRac1T8IYjYDV/n7OkWkYFWitvm6bpvgTI9UZFy2C
4pQkphdzoUjRKfpnGTgpYeh3w6iJKujMKTOHmsHFyyaVcCfQ1RWC6TjNsFQNjY0o
jdWZqHu27HoLEYXuYM/nfxjOQ39oCajpbRVa82I2wh012TAM1VxmT2VqkFKsNDqX
gJ0RIx93IrcJ6Wn4hrZGVM24gA+FAeow81fSWx5TD6s/LYSB0WKn3MLqX0oP/AMR
VkLJIA43f5D5Qssd8HsA3oFvAIcsHB7EuiateG4rRiBwAJLDCfhGNxALLsa73C3H
UI8eyB3AWWFZmJ0/2VLb1wGZv8kCBOHlipfNjUIXc/V152WQZIV0VHK4y2TZjVxE
p1qnfIHeNYgADl5u2Pc4dj+w/CPcdapd73BOTRB6FJfvOdP50S7+HZ/D1nH0euFT
088aE+Jws+mE2/2A1Xm0CGDccFhDAtylJfuGWHEMhnfRCWYJjgGErvGU40Aq5nGM
EENjXbMbkc1A/BCmVGcUwVSt0BB3Zly9W9kSv1ngvPXrmCqjDbFzHtXdp1sp3QHq
eX56ysasvCEAWEb+OSLBdVL89A0JeODZpRED/3eHs4RC8NcPJubs3obuzMbQFBjW
ML42dXXkyUQGCnHO3Z9F0zQZVNcHjzM22j1hQQrHxjSBSrKBzdRuW0lHNeqyCUhc
HaZnZ0OOLcpDs7+MLHrxj1aSQVyXsb/47LS4+ZwrbGqeaZxW+OqxQ8ppSah8vTKY
NxwV0ag/Nsb2nU0uzY6vlS3MUBzbQk/zoR/OHwikDqJruADpGUhxYsujOMcmrrHf
aSapDX+87dLtsmtpObTwBm7lQgsAWMxwnFkoi6vgZo4qX3wbdbuPSu2dyP5Rdqmp
wdUSQFgeL5TFn5W5uTkKovIfeYXP4pzSr9YQgk8oOR0SLsM0AuIpx1E3H4JLLxGz
btzl1X4uyechJrTNxYOTWzz1pna73/IBlQTy9rRFUMlFAjIuoccw587dP/kjvzOk
pGMme65AfSoYV69TljW/PrwGHxrWApvcseW/Ffxq3OSFpjgn0L5s9Q37fTjfqszH
EGEmv+wU3sQ4JABqAV85fwvtdFbJEwsKzUIYMFaaAj124QI1rEKu+4wjX0Vnbn8M
iREPvmcv4IXErynkaCr/AWcZHfopemoQTa7yjDWoGCQRjvxvtNFT+v/EhJEbnArT
VnorlMjQG7Pl/whQhlSdVBJNBSctjASM7pwo0dwxjwzeVXIaQ1HSuPVGp70qDz53
JEFLktIAzuwHV4nxaOJUXW2C/3zOAxyh8nXS80mIDh2hrR6TYmKQnuM8zXeKB5tH
AlddqbPWHyBUcVWZ6t3ceBNy6ZXGJukoLg+EVaXF8dgmzHnKuJVODiTT51/OK0n7
iS+BcnBHcXFhgaYqnKl7zt8M1P87nLeawAlch9xWyMy+SAyLoRD3NJ9xmV7NWxU1
rCN6vrAFJ866DEHf0XoS5ZjxwgQHThgjqH1+Ai4yABG3PGBWkwaSN6rVVeQHG+qC
ehvuHfWdGR6hMQU/BzjEKzbkYbhz0OKlyTZ7s98HB6YKKbzP7VrtRYjO5K37OKPz
NUz0fhRJENCwuhK6m52/nTl5Gqtxg8dRu3w5MNQs03Csj2pE4pQZmhWgltiDMb9I
hpHpo6cr7dJZAHeL2Tx493CD98Wu3mw575HL1r5SEczLF7XqSRbhTi6wmVgriFRN
z2nTRscC2/0F0WZgnns9Vc5Ar4qgABu8J+zAISoSCNRXptgNVu72rKRLEIquacpj
2HMcdIAcQuG2f1f/ANMPxpxu1QMp2Y3L+6ndnKZI65lJkzlYzRjDIaKt+y5Sp+wG
mXFK6wvbJMdoIOm6GsU/LqqJMcGYpRRajiL2O+YPqd7GnDgxYDJl49PiIjI47sad
iJjCUyKaoYueFg5UJcJEMFqaWzq61Bkj2a683Vb+Z0vZsbc9oLGnDTBfVprIoC4v
9bPcdE5kNpU3gAYBREk4bbFv6Z844qtwSRgElJ7hDQWqQDhHPTv9M80GAxGH7I68
KM/ElWeF1IuYN4QlPHYnl3OWFqqly0G4f7Z6ibY59Xl2R7LDTSdQ88+qoE9+Swf8
tntgf91tGfb1YOe37s3WsizfaZaCpa0u/QClAcssjQ7BoXkw96m+EJuuPISVxM2R
Vz5Ia0xAmpnhrjJokM6OkJPNlMCtkDzAjQ1BcTMcegPdd9ZiQmae++NvIQtFqN4i
CZqHxd69sTLKb3PPeC87Rc8oU4N6ccHv62FCe2GRdLnIDWzwZfP2mCb/WzK88d55
xP7I5d4ufAKY2ab8UFReSopuNdIK2DjbkUQwaROvykzex+MeTCKg70j8EsPv7+A9
SMsDS5MCs8totYLIHJdPsrFEY6xYFDtE66cZgSsgqCOxNZz/ZL2IvmfBUh7PFeqR
HQBIqCqQ09zA6sznKDyyT+aJiAPgSRzehY9yA4KrQuAwxt4SW3JHGJFbwqgtvLvc
qk5Z06d18ACn+P7pTXcLY1wjuovAetlNh/w4rq+MdhUbdqYBaamZOFqXXYsQgDP3
2H8ar6WqZ8+ylM/n30HkJ80GWZYNbOo07FMK2dJPSblGFQt6oY3N0iwHF8cgRBHL
/0WK0scmInlHrvkT0mHEnJCZkylZdpEJFBeDi19cHMX3bxIqgBTEsMAQ18rhmjP6
qGpUbxhYTkLPlE5sGU9gXUgsNbsOzSgb4UNjZhJE2bZpHrvEdMXi7+HlM3ItYxNL
kdo+KhL94Xa1HpwbsL7aouzwD7GZD5LuIxm+HArEsadDTsefQNksomfsVdRA6rt1
ETzcUHVi7lQcv+6IshM7KoPzlKr0L1z1gXw+3diZVvunOpsfLnf+yo8+lckU/iPJ
L4NYQcFkLHN6ZP+fNiT2WA0dBxNGKpCBmBzDcQZ8xLfOb44qMsmZfsFMsaW9qv8B
G/jHHzGj7MbICtf1rvrKJQvp7CmZ9W4PN6mc4A+K5n0cyxFsrZhztpdzPws3rFfc
t8UdILda4awWde/eQhZLiOl22N3WXp1WIabZ0Pp6oTRWODClIVzLY1mdzQlRZIrz
scUn4umSdLyS5RGYV+45cTYeHfmv5koPN18A0FmIylkqX6NbipWeHlCTHrW2kq4z
F6XPUwxMayp6BHaq6rNCu3AyYsmWKrzucAcvgAF4MBduF7nwD+l2YboQs9rEGFfb
MxyxshFpmIK7T/O0kMDeL7M7G071lB5O4KXiWPlAX6IYV2PMdJjITcDr12xMREkz
MbR2tU+kh4U6Rb+Ikcw3h1D/mHZ8yL0D+1D0HePCbKHOartTLNeeh6KySl0mZITd
36cOnbFtmPMrF0+GMcjn3yNXkn/FAOmhiBaJ5v1T8m38pXRV6+ILT6D2CPdYdfGV
F3DTH8Kewr6RAbD0AYg8QCj4ro00PrbTsE22LuRgKPg05WToifIWgXi3BXCPlKFy
bsFqCMIaSEzJY5hJ9QimYIqoLnOfwV88RUBiONLjZzIMm5rEARkU5usS3n6d/zua
t6uxQziDL3AovejXCQgfvPVRvGWtVJjpEdrXty8W+ZBhLNHvA2XbeqzvcFa5jvaW
5AqupbRQud1mbfoQLEZqffpoTiFX3H/5HWKDvr5Ek5ezNrETLFUsE54iwPTJq3lx
Q7kqCvIJwT4QgxO4gOA9eNh/q492lo1ojgvPdcZq/uRDBJ008+fa6V8N87sLUMD5
QE9h2iC8IO8MmW7ga0L6UZxRrOowPQ+S029FNDaBdHftjqXDb542p0C0Nc4PPX07
Jdy0yQrERiQdVPeDswbdS3sxB/v8zpKpLJkhq1INPOwT+EclL72tthxxjUDDlzlS
I4yI4+UCVAivuwNZOZ35QI9WFmL8vofko8R3NRwV8TRMhyCZfY9JmPWGxGP7PXEM
UfSCd0Ow9PsoJr9NRYtypSK7pwsGeWkEpO4HtGOCB4QREtSsxnnBU2GHVyfbUt/1
WDgQuoJAVszow0sGN9i6NoSdX/RXV8frUXQeRUdgcCDaAEj86DfTbV1vFA/SWL3P
ytBIaVe/Uyos2i0c3fhK1uykshus0VpKcbqvdZtVf1Gi56wWIcVvCEGuVd1a8DbE
n7fO1vIZR7g+yXHaBYmRVcYCJZfU01u3gt0kpIgN1i2cZIu5aDHP9reFMkkhG9x1
5ehaHyN1jwgo2zP6kAyXsHkVbLxssyWdyuRK1a8/LqHQQ28nt2TpwHZ3O2MwVMOS
/iLe1VJktNHI4281fsijdKz1fK+wVyBAAMero9LTJ7ciPX/oDf3lPny7UHEKyfwH
C+TIB3Dvg/Eh+YqVbk5DTeXapNbQKgGokcxrt9p63CbjNGderOYuPcwbLg63pujH
3laEek5CMN+8yx1jeh6njBl8x1aQ2nBVeXvcnZpQRp1Fs+va99k8UtxHXDnLrwVK
5OqZ3HsNONe+6yhDaWzvTbviQ6Q2ao737lYV6FnnOO5rigYJmh6bPSKDl4Egk9mz
DH3Qq5+WaABGfQgWmdkFDj7sEsvEn/RGeqWeMFX92yqfQXgM3O7YNZanpk2FTyxU
FcrwY81FLCwp/yqBUOjna21qUqRoDjR5a1vSiRQKM/4TEXphPS7nmpWz6Dv/dQyh
hcSlN5b/SwXwiad1cmfvL4y/WyU+urDmzqMUC+5BayStHVjlWfVc6e9LLfvsrPxc
AIxfDLIC1C0utTnVcXBWYinAmFG4DupnWDNSbh69Rq4wG5iy6tnuIJBifM6ifWZ2
lM2pGJX6TwR/MmRVrKSiN6l32HB8iLGXuwID4OCdonwQOdMPEylbUcdOV+Egfcn1
57IUZPRVZ/kv2o0rP31glqkLVA+TJV5x2nvshSjfFPih9P4YRaupl359lcWgtHyS
YHzN1tADfe5XOw1gzf0z+jSmTshC/sjzLudmROgJYc4s2L93/I0G0Q8eX+W/mgt2
o75ZQxsrnkviHOe7FvIE+ytTLwSMWAqw1hqp3S2OACz+KG8WsMAvqKPMFmHx6+wB
soBtpjvJACUsOp0oa2iTSSXvG74eIE2JBAa1/barVx1ib1uTlB1u2Qqi/9U6yf30
HfgOMxNwuKOgipYaNdjeHYQxEQ5Ym5iSYQ5FI+AVkJeb6XAP5tk4b7rWmQO6BJ87
okmJwrF8/6UEoChwxBmZR59Lxvq2ICmwFmfpGRxmYHsXG3Dd5e07P0dWjw6K9LOR
BWaA9cjBCn1JWOqOWW2w24pYbKyFZoyVeyJO11TvjA4kwthdDy4MLS5OSvR65jRt
xrXUVQbzDwL6ZMKYeZaK2TJZTh7/HLrCmBc74x6H3ZP+UWExzzDOLh6qi34R/dv3
IATZ0AXwiva6uC6ZGMeZsTfoidRORdT7YFWnWDfjKoKG+SChdWNy/dAxJ6Do3OK9
xJSzrzpUWRHs+Y5Kfilj8KOI+s/U/rL0mYUmrm4CDS37sCntfJUek+1UZogrBm2m
yaOpuabtqRatAG/nxdJ5mDR7rNoKsXSoqFscLJT/19gELp03IugMxHcD0rAbXTaV
jqSwrgcr0ck/Ps+HabaqoQrMFocTVVteHmINqDuDLkiTI2oJQH6n1EWdq05AZTME
I0qNejOcwg/ellIm5I0qPyxAZ/NS0XqoeUogUZ4eyJt0RuZTJw8qEjmVfWGpV0zh
L+PhiIKdQm5bQ3Baf+bXtEsqudywM+9YuSW4n+wNhBIXlZ8k3LoVKE7wtM/OFXQ3
Od6/CdH2vNg18P0Q2BwlgsHJyJnDZcfwGCFAUca82XdFDKYX6pMRMYtrI9xIuh3I
4Ax914AHItVo6+xD34t6KDb0S9q16LWhPQvS7jRoLXxmPcqwTK4oeREYBtAs3tgD
3wy68SQw1Jt4s5BBScT7DdkHMKV2UdM4gOYLfWVq4jzh8uY1klw7oOtx0g/nWuNZ
CTE9prr9XlodS2mZd18pbwUZP2JbFC9XVCIFT2RfdUPYAaqEuVjgZIH+OEBeSx3K
mOFJyOqg83V7PjDvUcztFqfcBz80cvdunhEMLwkf5Dv2CTp+qWPuMq/n6YdSl0aT
9qCtW3R5NLsYzPnECxvnAyhVFUBc/65zUbZX+DEJ7Fo375tw4PBO5D8wqdIP8P44
i9y/54mqUr+0PpbFved8R0bN2edFB0gOsaOd6hk7vuf0aCRZLt8VTaEtVJ7asbaH
Vo0dH9EtSWWicCQbABFDHZZzfwINgDkapKQJwGw744ELAamMP77HFvuz4Jzzz3OR
Y/73zkjfjFVWCmCgYX42QkJblZw++NzkKIh/A3hchBa8DDFmRR+GU1pdPUBV2YzR
Xy+VsinwceAj2jMYUO9aAw0lHco88l6t6H/+WjhsmFtLaeSDLTb/Vt1D2mYeLfhT
JIMJhkdTTBXw7q+4RdQjKdvofEoxUym3yao77eoMTepJmcqjPEIFbS4V5HFgKocS
kbr+X4BqhvJsfIxlMTsF4Zrhv7k1CRUehVWyb4E/r1teLuD6dVqgGDh21JerIonN
0KCV9NeTwjqs3uiUYDMs4S5Y54E2xpYsr1p/jS0STWuLYpjpEICBVH2de3R2SGFt
lpslZiAjTCPkD1/s5gpp384E5jqkI84/frF9CFQ0XHcd1wYfGz4qB/aKWkdiYPoV
XcLejfuk/0edBoj2EcGrrObfK7rFRcAQ7lhxd/QEuzI9J4XfK/X7jO79uaANFmER
9Ot+rv025Y0gQ9ca8DdXFj8q8jTkH0o+0y5C6iF+MoFuoFJS2i8dkJW0g36KyO3s
g6WYvLzHAkNfkqsRsnA4nc3AieCKi3rmGqz1jpgs+vYjAWw2h1GTzo8/L6EA4CbU
ZatqBhecGVD62KYOjeefiQM7PNtKDLLEqs5S5er7nNuByorjLd4k1TxiHDgZnx8q
fTmAT8Ed6cW4imdO0bley5zurjo/b7kFMZgJiToVXWDB1HB7Mk6l8EXUz7WkVhrF
f5n71Wxol+Kx8b3Be9GmAF6wdbCK/4QXwMhIhVNMLuk6PfjNtBHopecZpHUsrLl+
H/ReMsYW8l6qN7o9vvAelHlXL7vdh6el+KRwf/WaXLPkVIDDf38UoDWYrZG0J2Rx
73oqgWLIZ10hETHbeMbrvGefwfi3/5vCvDrXVP7Oucf5NIGmbWeLH6wlo1qKKRXC
JMg4ypss96mtjPemceIJThfmXG0YjJ1iAIlIZlaSLTQpi90tOp6W0AdfhABT69l3
xAy8I+qQtIUJegIJKeaDE2lusxKU6IF2osKQ2evmyOAsS0Gx8k6iIzWpmNnDcyPf
6rHtmwX9/zb20vhAvGdcpqeEgDAZ93jmhQb6H3UQ6szQgiaGJJGX5BckQXlmuAfl
6hOsaokgNBpqgEvuks4gldBLau8pDi0DQBT9+ISxWhcKwCtqCx67W5wvFn36V5ZE
IX2m3Nv0me24+o+8MnAfbseqCrQfGoNx9iE1WLF7GpyzNsw1BvEXQhEEqyl/PKAZ
YsMEcED+ARKOoaDQQIz9cJ8fZo9O5qnbq3f93sH2J/8l9yQ44V1kHcY65DVCrgpz
YktpvgGL7LmB/9ooDinaaXRZnAcaNjqFqL3KHs1S7xF5X5UWQS8pZJzotZ2m5jiG
dAADCjSdfaEt+Zg+iZwYNKsetMRxze7F1BLkQ8lUx0Y1dguV8tEN0Rbd7L9zFWUU
4jVLYfat0SQJdOy2ihv81X+0Wb+hNuyEQIS3Mk5vb9rTmnpTrShWUWbmkcZ4FKxf
lITltyvHTy4IIub69QSO6iToG9NohJeFtXnMsTLzV0U/ZYLc4V/csTsKutpG4kPW
O//PH+VhRyyuUEgrei9Oq572NWCiLxRY/dNY3QDxSwmPQf/gHINyFa7AoZtMdeTf
SsFbYihktI28uxVO8fqBk+Z/tNyPp4bT9hGQNN7GHaW+ozK88AyGapAEvlVjQgI9
rabwCumo2svla4WmVEzt5YVsPL/VZ2lwaKzeRk3CDSRamU8I2B6nzwcLW13/15ez
4gJmHPCWm0jQuCG3aNWG5i4sqpEiymHSEm9kpS8sYBEtL8Ydqk/jrcXEezCh3pGd
MtTe6UfjBpchORjWJwxaGgpxmtLEmpUhNCUR790oKLj7pWNtjw2yI0rLiSpvwv1U
0ifp0f8LiJOHnDfB7RrQVS/r/3lD/2Y1XnUaTvvhL3njxsPKQydxI05OwODUUdf8
Oei3GDyxlQYgkgwsRya81QnAGIMRJZMG0MDH6N60V/uZzQTlZ9c2+qJdDF6Dj5IL
MPjt0cnswvQbiD2fAw774Mg9jUpWMH8j6Y6xK+jPh1Cts5smOgDBSz4k1FvZ+yXs
FMbXVimVOB5GbNnBuQUbG8i2cdZ+cODSN5nWp5NbFQXU59OF94WDLNkEBrU9jd6j
wvCfpg42kvQVIGVPnwJI5PyOcnpV0Re4gmle7yj36rvZU4zNB46hTZROmx/hn3ki
zTBgDSnG3Erd4aLlcxHcojYT7MlFW85rP2HEYWGcoPv7dQnuIcMIENLFRQWIfXUX
4njsldGlsatqxmLahrNjP8sPvrUuy1hrHiSLu+YA+34qOWbojoNJVU4scsSgS288
xqAoS/dg+CLoDt8x7/Y3WXenqVyB+XQjEx5DkA4QF7bV148NH4ytDF4T6JOqRzbh
jrPAPKdJE1ycmBqmStAjWnAXk8aMv3ZdLgdofDgVdGCTpOtLm/wmvG2gin/Ywsfm
XVxFecsawy4X1mTXA2/eGFUylho/pWuP3H0jvyW6wLYaS6wsh/hLiMMDimQdvabq
8UchQ6Jw4Jf0nsFywfybvKTkLSWU8T++y8ATLEyx3V2Fju+EO5F2bTahmUA+mzcK
9DZiDgXx5PGEBiIVs+Yym8g73rsEltpgbvozTaY/g/9fHMhUzHfKE6Nz2GLBbBzb
d/fDf9anlVafLej91EGznMf/AcalBFNYcBrVN3sdjr+yYDHfyVq4fRVZGY/N4lS8
QEnLEO0891LhAhO8Vx4F3+L2Q3tmHu+GF4kaObPUdJrgaJfAWPIDmLrCXZdxtcf/
xFQwWyuYh+9MqRLb+CHN0J24jr93x2IComHDNqbFpA3VYcoht9b9+267UrrBNmtU
2Y9bBd5gihzyv8nmSXV4s8CckmwlSYaracwEViz+cA6KslkAoe7S2k14DdjBag2j
QsUD/ADp4daOfD70cWk4j+MoX9qaC34u3KaJVTYOdpQT+vnjVevDrpHzZ9zs/xVe
9eK8ntd4P0ugI0/QLXYSs+Q3ab91IsLqfRwfkN7RuzXSncLPvFvk0a4WBB3XOeYo
pvJfe/LhMhm6ElgtpXrPzPZaCw/e9dEKTrQqkPBF+Zf4e3cagy3SppB06pzZYVva
RG9iCJT6NMBDhD7xi2ez4ejh6SAcL39VjVkagCzAfeqCi4MLnx/aIur2SPeywCMh
/Xv1vUZy+RFJJFkLXCa2y8izF/mEGc+uWLxZFoxmR1FibSGP0ebhiuiGK1f7MIWI
/MaeE6yqRShrdOWxYdASPIs8e0UzNZl2l9MCP5EDfAXtEeEmOSxcOlGDg5xvh6Ja
Al1oPeSVPenPjlkRG7HITBZzZc1QfPCviWUIihl+ebJ21u9p8q8hI/ylR1UqFSWp
2tMrYEs+yUFKEw14HzR94Rf7+orynJbXqa2vecZNc2E3YVZM08hfadlluOR5w7bz
n9Q0n2t4JZg/XxLgsSe5gSDJzbIT+UqEKEmvhAZEHK1OUOiVe66h773KPeK+v8xn
1Onjj7pbWjw4HPn0SUAtzZaDyWBuTBs8wKzy9saldTkGaQ7pheiDHm5cp7UHDDkY
JVPOXYJCr78bczQqRDw3hEL6R5eV3JzjnQvwJySDU84YxqWsc61J8sxRNdx9azK/
Vbz9imoOjbTg9yS+Ju40J55lvLnSycFcYDpms73z24xkaoNu6kDLf1TnUxVUuyJA
dAWPwqdFvhvCOUkNfhfM+h7YhIeNWNda8J48nIuY3oN6kEt1NoVd5Guv14XzO8SZ
7DoFyBDaIypRZ0bkBfQzGxbpgaw+vnyryOJULdCF7t10L4w+pEY5DrOEu/FKmpTt
uxsI5u9hpNp+cOgB3/+wDYtThswt8npeRAvZIJemUgVJRczdsq0amyRcW24JN+so
ZSUUsxJuda2AfXR0mOHvbuRaNbiT9t/GvkrNdquwc0wy+sKO9AtowN0UHkBEK6m/
0rMgLR0pmoBK5YFaZ7nuhLq0LmN118pnEhIvaIBU46+wT5AzVj1AaEfagR5A94QE
lq3ySIN3bTWdwd6RybsiAociKDCm19ecMqFSUrgm5efJRkeFEmqoA+LXDtTzpjg6
XfKYIg0xT5u/EI6pBpbOCtJifVYtygd3SAdGkN9TGtGB56OGgxL9ojztxe5ylt5p
jeAQGRk0iyJ7w6jqTlaus8TY46jYhHvvK3N5uyVxCSfyWKpJtBrVnsDAJHq+ethA
tk7uIOZ3+uYFl/eZHgQEVdVpnRG4R+47Uv6UDgGwXy72kp7ci1nx8yLEZzsSO4/6
/xvzqI+tq7gSM0Hr8W386dbg7EnNPUtjLu3vE7McBFRSzrFx9SXpkKKqrl2iXgtS
xApV0s8iG3J8sldagBp2B//PzxkAI9QMseEF9ZG3PLIEQbnugp12Y8nuZ2qDmoxc
dUXTmKrBMVpw+ZTwW1Q8Zdp0Jp03/ZlZnVjZ1XtJWWcDXCSD1JVn+uZ0qmkuGYaG
SU+2+UoBK/CXeYIrhF+6ljtn8BNjE5rYklhtjPSg3cJ2Uj3d1gWot1UXEZz9ILMb
/XEARPIznmPLpQ6YIAzPPYj+8UDlKmYCNep8Ebgnc9d6EFKfTMucMYc8FxgofCaT
e3ZhNtri+P4dAYziyTClIpQkVOcjM+4z0g/Ntta0H89pazaLsFYP0RCw/ZPJHRJa
8qj3zsNfbyO9w/TBPp1p13NPsnTmv5+5QEAGJykYjYqvUsMBASHaQbBTg/0NSnye
vOxj0LzKnlcwUfRvm4gEoRJ8Rs96EzqCL/9vNAXERr8qSy/L86++EIGEoimPqdFI
GDCNyOJNVqs1h5GwFmPszHZMGxgp/6GVjwiBNRjgcdQHpOeveOUWeb0vP28GbBrl
hKG8l5bpJsTrWm7EE1VsH4oxYl90remFGi33lQoDINKiJ16tv9tikrxNR6uvv9v/
7MNBUvSbPXrKJgqDtRVCwM3PThNFKmI10T/2gAQ7HQtzKzxhbV3fiDquf28mY6g2
KBoQYnCQKzwwyixWDfF7cKKHIWcESkC+TrCHo4DNJsE2FqjPRQa4H7mVm/rIVVrF
GyAKIALvnfQRpfxsSCUFRkwmyNWU19T4qQugPXcPB8rn1bzT3vjGxynirTsNjA4Z
tcaV/H0TYYl08kgMjGbQsJ6X1foG3GdjNJE4SiWKlk2eYl/jcgMD1YNquT2IatTY
20oNInhwWy+pXeQhHcj9YZuZpiESf3mSReJNy2RukFRdX/bxo7IJIjabPkBhPIIy
ipueQhvyAYzBfC8SdvavhG7Cm3F5NgK4YCBrOL5lpGEFmJY1L6r697U8aHCsQ23V
LT8tKnRco8gJpjrDZtJdt+xb43c6qI3k5mqs6BXPQeOJiovfZfSMfBdh0j5Rt4Lu
PnWGwv4pHIm1H8xjDdWY6IquA+i3t6Mks+3aUkKrwdSzvexsC3dwuzLEKmsyaSD8
OQkb4R3ND0h4F/9P7mrHsgNh1a9NyMgwVV8zaH5k+Yh+fE0j5+Em5LNa6gf+BNmN
em5oSoCHuQ4/3Bo7DaVKBqsr1fbJ1Tg619mUHJPugU8Jof8O1DOHg7Vb8oZo3pmD
9SDoWcGNblVsB6tXVaiF27t/ZEkeb9jtpkckF8DjCm3iYQbed9qFdtC3q3mi2Kzl
c4BkQWh05SREWuc3YUdk/B3LNVCO1vNJHDv62OZDlMx5b9oFWGKMu6OEpl4E/pmc
fLHnShm4QQxWDcnjfsZgcH3vLw8KCoVbMaMHs9Lp7dSDOmGxh7Joh7H9SryUOSEa
rFYcSlZBpn9AnHyF/w1oObRKGZxB4FV4/dfkWlh5C0j/i/it7OOsRIEGdbjNnpNS
x2mzLo5J5HtrtDzfzlz8XMYDHaz6P/LmbAS0y3U0ECzxhl8En83VGJ5rlgX8mcQa
B8PK5gLS8eyhC+0DPSBYnLg/h68YnUy79bW/ZTJ5dDateBOGitOXlfAy0XquaoEu
dI+0rrJEcKpaQJcQnReuSD6hzMaYhViXvSCypcKTMZG8X/MrOWtVeIsFrNN2Klyv
SJ71iMSt3eVR6Lc0Z0OkWhlWhnScWTT+bfMCBpuPaVtqLFhv7cZe3v+Y+IB+PFR3
VGtTjaSK8y3mLjs/4zXTIT1TnYMXosURAzIrrudWVq73sC6lFa+M25R9G5D7Oj1E
7iJFdCGyzrGkSLJ4ERSACID8HstuXcmIdGNTA57lHvL9G4S3DseNDK5YEJIgyQND
ZQrRI/yavfwEBN7q7GVOtZPJSf60eimGwrruccOM0rel0GfEq/P/XPwKtVBPkcW2
v0Bj6Df0RhAVAl31PO625pwhAnF56MUTLEuuLAz5/Z5oMsqKPTzyRtb9PZ8vN+IC
SSeZ1tykmN+XL8uKVnTUTonLxYJ8fJwCPE6YHV1TSxiDpqNwr35ae6RyQKQvmzs6
3siQkqJ5/Yud3UaOhlvBXCBZAioP4Pl9aDkhY0MbA3rDDFo++CLf58uNtScKOnzw
Qzbnftuaj8n1DfRU2Z9D2FZo/WUA/vyQDYErRRGiLUer5xf0c91SBUVdjQWAtJsF
xJP5o8trR9LK40SzNP4F1fy2jgmAOWF4wC+7FnYICefDrX8zt/efaJFT5Ys+jzkl
l97SgphACnBJdue9P1RVnO25RCER2VD9Q3QL9uMNWs/kKnA91AOijdgYeTLJUQDz
xOZ2HwVWURq8kyMcs9ww+vwaoD06hHj8uWaMgAgbcDHlgsyErat0RU8c6CawefOv
LxitLutPeIKdz4z1gMGaV+8FIFff1ibKMay1THZAo+1+U1fBTwAMmMwYwT7zP/dH
Y1bDmm59giWELRvPFmW7xPhqjPXiHkbtQUrYpC+nMDH3WYtqINJuNcoAhsuOjzsv
JpWmodGz0kPHFmmlAU/H1Ghj5uhCOsgZK7YjAjEamwzzjQblDP5eZjH4bjuQuW1F
A7cR4uZ5Ee5ftTDqZba95WKHGpzP7ljNHER0PRWQ1qqJ7zbLmGD+Yxki5XnSag9T
2u7JgA76KClwtDsmlRNeJuAsyDg622O7wE/OQqVf1Fn+EtkQEt10vSt2MnPMBpyh
wdp9OSi+wF15Glp3ajfEsEhZcVjJo51f1nKQZh56SHfOg3BHGco2mroOtG75i1gz
9nWrggQ4m4SIU4k/S4e9Lp4HItExtGjRkfYPenIIXy4JJLiPD92LdyjhA6Jvur3Q
5wNA3Ntnagh9GuFwLiKxAJq6plmOoJe1xdv0Xo6P4ODUkLOHYH7uTVfPndIS+2Mu
ZjRo0f67j9TCnNcrGeyekW3MlpR/FLdetrNyZSBtrBHKlDgmICecxAWgIhDxzWi3
GpKAvPX6ozfXim+mJoYjg0Si407mXUhNCF0B0AUkQI997X4Ec/0dKiU9IFxOGtBt
jBz5sYVZZTM25AG061YAn7p5XLmFRxxPHCkYEQ90YdkbhW/NVE14xdmNQvRPStPG
oMFSUOXlkOKdAfmrJkDR33EuQri71SrhDHh+Ep/pqjImmM2XvPyWoc2rXRaBZXip
goTvgDcmYzV9bzPEf3E4rtrL0FVWehOmRjp6ohjOXjvF0bFCCwB8eLx1BYNRyQLn
XK3Uu6Pz7rJElHysFFI+HR20DUxJeCpTF51JXomWrE73PU8RlhOH8RBFtFjZ3kgk
/SRQ6NXXVPf0FrETbqv5eH2awOUGySkIBnHys8P7sNCC7EzCTPmOUVXbprLcymeB
o7zUJlqseim8pPEx+OCpw+10yLqzaAOqlZdK596DjWhYRoRslDthznMuRcfjEwu/
hs8BCKoqrW/n/hCdVyUFmrkaxqjG1RmwbQ858D5PphRQx+57+bVyxGCCSvue3arU
YGDFA5a60R1MT4Mo1j7NcY2o5sb2KWHrRXDoICuC/4tyBXk7AdXiYLqvPa4VAngQ
3D9e3b1ASrl4nexymlsV8Ad+xqXYzRKZheaR+lvBO2sJc6HcZwzLe72fxky73wL6
9b6dN1/crTFVY4QP5ztY6AKC0Z+s6esPfYi+A4c342wJNfPEvyZCGlEplXKiZHkp
CJN5XIGNLZTepohau3FrMxRbvihSS/FhCghGzf8fRhR3eyG+3kEW+vIbgV40bxc+
CTxzhoDX/ta+ABSF6cmwllVdiwNaP/bJs71nxBCimrbpBG08akNdbR54DyGkQwZ+
A77Ph1CN0bfhS5POXztBCnzWNgSb7e5FlWARAMubNGJfYW1jTb9iDQhM+UZIboeV
6u4mLMUaQLS+NfUhxbltxqqQMUA5GwA6OniJczj5dWNnvdZRqwKpEyNvcROozQUh
auejK7PTb0Yu+KaWDbm5wkl/gXQhr4N7N0ZVvveSCWI1IIrFO7aPJ7VCQm/MufPH
fM8rKhLeo1ONBHmYBG3/kAbAxB6IZeElu+UWsF+qexKqCdMTtucCAAWe0sYrXr1f
OtezRGVcCGI3JlIrjLeDdGzNbS1kfbOo6qOsa7meht/1Mow4SVfN9c+LDXvYItv8
ljr2nhyUWgMDYeTbRnxsbw4oZOnc7NZ6qHP/JmXFrjcSTCYUZxsKKRL2GzdPTPbx
sieVni1+AXjxcmdREoMll/o/B9IL548LGpn7YirO2kOilNSoj9ZqvgHVaBeT67Ls
rCuWoCgPYQjxn/EgTwfUajfF34jUuaWgQ9Qe5Jc6b/Ca9T7lDhKuwE4CcXhERaKL
5XfeWO0xuAnCZvk9O4FVztjRIPvkV/1v1EXQQPXbJoOb/8n1qdoDJs0F6l4wp3fh
5hHVlqtTMSFrwT3M2CieXWxvbwQYBfgKixXOF/ubiEQzrn4VI9BqcEhiffRFBoon
DvPTqkXM2ftj325E5bZuOZ6gSm0wsRgFmgkbv7WN8RnAdFWxU7pucR8qxbttMOmF
PCBdKmD6FGV4todN+PKO/5juiILooEW7AEP38Ao8aBpAmyf+AYOKGdAl1bUrIjue
GmiEFi4eGP7iOSrW1XbjmZZeODrj5kObBTnNqjqt17WxArCG95lmKInMKO5a4Yax
yJPKsuLLROk99srQ++VEXAHYPN+mx14ZT+na52de7dbOkQjRvJ34AFg+5EreYtR2
P1XjB8umVXplMjf2ix2PPUMvpVB6zDxUwpv6rWBqFECw50vRy4d1GaX/4Bjh4ppo
cKMiCnIHxHqn5eJBv903/d4i520PQjqrYiOykVT2G7EEztQ0FksesPlLaYNzDwX1
oOzLcVUFbA8F4ZEtEDIrhRO9sHvWVuCVCkT1N0Ggwn1CuPRmbtFA+MC/xIRIskk4
EVd8hqdZ7UVAmTXG1/mXpwR/g160IxRCNzuwLmjNKz2CVYTBcsoj9NLvdDL5Sh5Z
1p9B6HTN2ksaf0zD8dCE0Plfoq8NgJzKlu1qzjYvQG7qaD97I70oaWhPhRJz1QYY
V1ltJQyUTRyub0Wj2OHnOYX9BRs/ZRGyZjWlRsPqdmVHzSc3Vnn8UgMYnd7vqffZ
5gxU6yPnumIFBwZIP8IF7zHM3RrcgDF2RreVDtTw3tQl2yHCdgfGiHHe8hDfeqY5
vgT4PylOFesJxUYgYjm3smmyemXtnErEAtHjykW89UY4sFzXwQGb+Vfo1a/EFAag
IQEYZp7n33rM3pqipgQLIe3OalEWz8z0cleAAdISMJoHbCH22rBESYszpYov/qwq
zRI9vhYQFnZ3Lrs0OOaLtQqLJs7epLupZh+UwMSh9VrrDnrboy3C0Vt5vHiK4Xi3
DzUJ4MPHJ2+5LNyI7d0/1pdn7a+ReJW7zbpod//C4OthvkNqJtEfgngUhsQvYak6
Jba+IRnZKD3R/3CTU2yGWRhf93+2LldojeOKdLga2/tNQ98WMap+wxyPTpHN2lmZ
hyLwVOx0UrjmTiJei4l/Tzn/EYlNGUkFTQu9lm4XqqAzQpzNE7csyRxHsXi3OTfm
fbLFpOj8asWwO4okfPuIWsqrxHS9Ul/eIHzUlrQDPZxaTevEzp+/bwd4qD3PcVZD
05XGLKg89wZHxIi6pUP3tEwXkgq7vpkFK1PWrPnPyTq10CZL1/4/UlJso5igfe2J
IXwBJt9mS6F89EDmeWq0RmNn+r2n9FQipcr35/8S3Uzx29VVaSeLIooWJnlXC85z
gmIoYDhDNrLkDzxrrx+h3AsRLgcrtSVPEWlcwpqofFD1crhuLENrdGgUEOM7rUSh
SsVuUT00eJo3G4s+CQO5mZAEWJ8L6B93XFPFj3nmKJqMzqu6dgFMlbi5h2ktsGPA
HbxZ+OO76glcXs1Wt39Drx3zvSoQFYTNxp8xezdJ9TMD9/r9eHxtxpPVpsqsPuBO
iFZ4QTLC14yGPUufGh8l3JO4IZx+fW9k1SazH/3Uy1u/xWCFSGXc2NjOsbBEVB9R
BOUC41bQyAQ8mdlVhZTIJ0MPmbLXV8MT4ezJ8QPmwDOt4SYP0Z6XXLjT8Se81W6R
+oTKbqtwgXMJC8vevP9PjENvUAa+ryRHvWqQbHSXEXqPhTP58+4JBz7I0uupri+i
QE0f1HTY1YNxn5hRX/heg3ncpG5ps/ZdsEjLmmw18w+DGCiZ7Dt95JOWEQm9vjk/
ubibezUxxogjqAlRTAAsmTcxVI7AOCS32CKeH9190+50pELX+vuNG9h4/Z0BerLM
VFuoxR+N2c7I10Uv+yTINlK1ktIuPG4qK/qTFNSxjshUFkWvXP7S8qBBY5Ne4U4y
w5a4/fwMOr2kCCibs+N0fx1dmMmS/MKUxKi2l32MDyCziNr10zqo5ClCnEu92MnL
jcqaiABdyMoBuj5jH4Tf2L4AA/crTmg3jH58T1WjOdTFJiUQkeLvPExjHxhUcILi
Jim2batELQj5avyaAtmqL8j9EezKS96vgPai5G9Lbtn4gJG9E0vZWy5M1awdMzNf
RZOrQ+ANJ4FLnrYt3O5M+OSQBx4K8wH4oRFJzE2Vm6PbRtFLF8AqYyRG1fBcrbsr
mznCrtWsyCvy47vYImBth4gSItcpbNL0z4gghkaW3o7H9oCnrllB58qNAkX1+1o5
rl7Hgo/Lzv90tBpqEW5qMPbhRkVthv52Iwn9ukY+gMfDeLT38Mn78i8Wr0Xj3JcB
GhpA1t5BvsqB7CksDOAMXK4KxOOGBay+CclmeuaqFDKo7xVCF/qLIQ2r58Oi9CJ1
pF+5mVlXvefuwWFTPLSSK25eyHKjpZU+RRi/OThO517MRpib1zHKN/ez7uqITNFl
Y24BdviP8DfaFBT2rkOrDa0ZfjhrvPhRCx6ElFNYlDmW31rkCgKpAqSUby8YK6Y0
lmiCipSCAmoF9wUbcNDp4RAnM0DoLdAQDXH6kcj0kJDlm9+fHxrniT44GSZWk7Ec
ypmDjPO4Nz62Vax4xcY9jVbVB/5ZY22AT1dCYyvRP/V1IE1B85I+eAnPUguc1kJD
dmovNXcOS68oKb4WtYFYww+aUimtzH/u9nLX27l6UUeeZI0hz8HLqV7wFUgpPzET
aNGK6LkuD2vkZvJZM67lsqVt0AtPSRt0xeGNi+7qYvqID1cqhvt1EAv7QfVqf+16
ckVA3ZgNEHsXAbiVfTUlMleijif534eC7V+p1yHn8pUxZzxPTJyX8ClQBTTXRlY5
k5LM0nanJHdMZ/nst71QHWsrRL4OjGbAP7js5tqJ+I+2q+prN+KRaQ5eEHt0drUm
XKs6ABgekesEn9qZyVTSaBFpCkLyDTT6dRWOTm4CHUSVYhUCOtEs8Iek4kAFCF8W
vVVfqxDtJwZVKT0suaqMTs/wEmWcW7BNkv0Bv5ZpICeQaQFSv0lQByag8FF5K3VY
KB0LaI5RQD1FW1qKjTpSzAnfWD3X/XUwf+pEIBEGhuXxwcAeWIP5jwwH1I/j8TzY
mqk4EpQ4FHSqRFQFxRmo+mZ02FT85pQ9FilZig38eI2zrMIBjITLf94TLAKvctgH
/G+BakEd+1IIdtczPbnuneCfVMhC5HcUDp/AuBBWLJOu25eSwvu01yjRXT3o/OGL
epWKZ2CzmlsKJOZ2M4/A0OkQlmQpP64LTRy2P6kN1FmQMZRunqXGFv/6efkX7CS9
4VjGiLbSHuc5XCvHzd6JKiYDW2iBxrWG1R7rW5z6Z5raSMd8SZ32ZqP7fa8tLfSN
DaDxBk5lwnNx0znBOW5Z94oH+Xu6LyI5SxDc1swjbW/TCRiZCyLwSz0BOZRFOFxa
VACneqw02NygMnmJpN8o3Sd79bWo12wrn45+7/RvJgLG6YEKDH5sTZxA8HhQfCTU
vItth7kdoZD9AxQjG7W3h437AJUR4Rp8zNWIU7a6L6ePqHpdqIoihb7CU0NhbUG/
jCuTqvMo0RqWLOzpWObIqn/fUcyPPSRpRb1KPW+UqBcJSHKdpCWivdrQ+ePLGLSR
q/4r4NLvaNI/Zr9yLsfVR2Wt0pYipSrG6YIyCvoSYfNfr2G6SRE+LBnUia9ZTWJe
DqJ/QMqmyltd4KQ50jInykeQIE+QixYSmk55azYV7PhpeW5bFL0tcEimmiJtOrYP
58PVl/h1Ngc8ul39v3Nx3AF/WZ2qZxNV7cc5/lQAa8vo1KyaaLMPvYYXBbYGDc9F
klkK/1hs18BH+xxqluGuw+qeT8go2DMSBeOHbj0KZaxaUs8ri+Qg34TKs3QoidZE
bUZNIZHszJbJ7sEWsC2tmF/ExPnhYWGmebRIRYmm/UiEtE8pTD4tZe581moAa7dB
EZydd6Z7nWZuXcchpdo5jjwQUmzP+a1GlWUuTyeUohvF8ro8B4rt3LwACOZsRxAu
NRUT14ksz+Us2Kfx24zzt+EQplEQalsfg2t4XiahcdU8A94vGXvqjZV8AzrlmYIU
OdaUY4RMRFEBkC37TZXGJpI48byG9Q9TuvioU5Fae1Bom6oxNvmrZaWqa7xjqdV7
ca8ih2GOgu1H+Ag/UVk6gd1vksyQthK72AC4RwEAwAIXm8KQmFFWCqgB/YV1a39P
mEJTxTJsyjGJpoFCtm3kgKG3g0aSwrCjJwkSrP+FjmtEBFi8RUTV3oYjJ/BwFmBh
cOQruDgd2tO+CMxVcv1qSCS/iG6ugjNczBf3oy/joYE99Fy2Jkgs4khrqcIRpZcQ
QCyxJON019Kb9Dl8leVkPafrmeLl+Z6qM7jBEZDMpQ9Egg+BKCUDEPWf7ArqK3Ec
1C3NsF0o80alIPrGBHyb0Kw2vEo7gx8nfnMialmxUSW+6+aKP8Zn/0Zq7btdRGdc
yl5W7l+WDknQDt7uPnr/ds+o+XnfWpB3hjqcyEcXsPpcjh/fB9evkhy0h8nHvWBF
YNcLLlEZo6VpAfCZz3PO51lP+m7Cdprd35uAR0DlJNOELox8sxt85fZsmCcKZom5
pPASCie/XUBt9NZwMmyIvw11yTWYIwif2o5OsG2HG40hxi2xj31QCkUFC4iDG2H2
ETQEts8ZbobXOE7Lvj3vf21SKBRUvI3CYYZl8rymfzuJ4MZPkWsqQik31l3jlz3W
/RH0IN5+PeGCsH7muYstNrIFE+YShvhokIz1A2fywEF0DaYGGA9JGSXXAUERAfvE
mkRFtGz0zVQdkTTAEaxywmJ70d7H+KEIX2CBWd3mxOE1RcVWDI+mcQeEh/bvixWV
hSIeJeVi0LUpyiue0kT/rpV8gPUh0y0uHVIbhJkuSKjGGPgWinX1o3nhymXHquC4
9lPqGuqeNo5EvWDfwWZqMsMbFwreRUL8h7exwbsMNeMx8UUisVpn0mNdp4BhWI3z
oT2lBb7owg6SK2Rbz3GSzrDSxnK77lzKlSxVAzBXmbwHiUgmiV6280SGEGqTlUnw
YDGKv/SUlWrXCLNqJ9qVCPewJ9lvHfYd/0G9oTST/pEq/eRLHVd7U9/aOMKTOzHy
ZrQvNIRMCo5MC02VtFGdP8Beurlf0r4Uvo/4D4eAuiI5wJtCvyOwmhq6KtKO315O
lZfRZlx+rYi43MMR0qrVhJb5oHfq34DuM3SzlGhdxrdFOuNrr3kFB23GmBUM5NTk
jkP5rSPnRJLHk+3RPBYOMcCgvVLD1ruFOBzP7fYrm9CrvI3aLGdXZWiCqPaVtb3j
TYftBhoF2i9r7F8Mgf7PDhctHK1h8YWpa56n6ezMZYO4X943zF+gB5wNLYLi307d
SGKkCzKdQKVpelw5grhxa7n9aSsAv5mjHchP4UaR7f4P5XKhdXSyxQ5iPs/vnsiT
d+/GD4xUEvo5gdzMdOVI1iOBo+FGe22GDwVONCT7WTPyeOB9IytH02Cv0US6lyFr
jESFNprLsCqvH2ya8a9lRVnop+uGWKkNr9dDCpvAjHvNVv8GO/vCXx9UUnJN1ecQ
zitApMtoroIC1Aywvog/le4VvCxhhBEsB1v00Y5NtHImK+u+JQQBNVZ/sW95pK0Y
psB7GUguXkt4bRfKgHijat+gG7UN3kLLhimlqpcTdFNeQ5k4jWnE6BUfnRHMxRRd
wAJmkdrdH1zpqOWM/5BhtuwwokMNtM8pZ9z9W24i2fo0XPB70tT3bgOhOz2J26q1
w7gBQbZ6aSzpzHkNgXzxmnHGVSh6ehiUDz2iNimLoz0pblsYyhvrFJXs7Trq227c
RNS/Y0/tKtM2x59Dzovbis6BW0thMhQeuFTvFbCqcr/eIZK21rQ31EdKigdtX4Bl
RbF0VDHinsleuO2kTH+X22B5zqqIM4TlymD2oV47uHU9qKUk3OBYa7j946KQwqig
b/5ssv7mdPOiPaPm0n+VwmwhvYjzfyM54Fa31/YSCZY+EgE/LieIqNr3tdx1ruxm
6+eAeDYRfj+1ataoYKYxSKSrKd5NW/Sr3E2wj+fsEZIH3kVN5zVPDo3+Dwkj8/tl
F/30XtukXZThtpH9egDUwjuQ3zZIasIt4huxlnquXvMBD3aSnuA3cG0bkrGodbRg
Pyzs668pyFQXKZaUFXA8oyeM0QMcEUq4L+dFYzFpPzUu2kv0JFpyEh7Ma1FEXuUk
H65iv7CNeesq2nTSjP2QLtjKNWv2PnRB8x2aEG1ej3gRkwAFOk+LU2QzuSgBy+ga
J9TCgqOtEb+uqJx6a6lliUuOUoBVdsYaxSPFhpPFh+vAZ+PkmGWUPFtFwmCOz3Oy
XCXPlynxs5FWkCwqL+9nmWeh2Th1blGIwJ9CvfwDolkksTqhambfIqxWNk5Yr9lJ
YPtrMk47KmvGlFyh1tojPs3eWtGizr1PJa+sBPYLWp5khSQ0STvPxW21MuBQMuQB
127CgxbgQI7AS1fG36eHswJ34+Yko+IpPF0sGNWmcT3vKUAE34vTylliaSiKoU4s
SaFl7u1OXVAQ5DWqFfMl3WFTNDFq3x1vYP0zPvzc51S1R6Ddz5LIPvNzNjPl0lcU
dat/gALRcv6slDLI0d3LxR7ZoDA3/gYjvKR5BejQ9g4wXlOAXZllgj0rXn90UR5z
iyRhTgLAH3dpkipvf63Bo58YaEdqm4Bf+iNfw+rzbsLsv8bGpYPjmIhfFr0UZgAz
+8WqCak4Y8GhXMPcc97rm2m/EXV+dgOo/WB3j1izLct28pFvH4DJVtpqbUO9vq9f
AVJ/umN8vLtgGImWn0fk5a6wt6uY9lidBoJJ3AGfk9yUz2RuCczHH1aSl0isnawK
axSuJ5SJ6iIHGYmes6HZ5GYwq2Rw8tsQLb2SpaN32pkxEb3rNKgskHqusFeg0Btc
Q97gT347YD67GC+qbMzuhs3xmIMAIV3NeOq7lFz6g+3JCP5QasoX5yzDuvTbptOs
jcRawwbe47+NKYnBnT3MFIWMM8tYVILVU0v3mjeyhPb14MTbEOGgrDsC8nls2faO
ruWKxUkcVbebLOT6KGe+c8vII9yJ+1L5v8N+sfV794WNzTOo52epOHV4geYPSaLc
h4RXovJdpyhWGzaxUWYqwnSVpf9Sc44xISymlG37xlgEATa471ifylmdqBj1+WYB
3aTkyuooTAhbMzjix7f1bBzhS7vbrQ+126b2RKn4zhptWUd1OqvufXrpHuYAGgys
yBafw3L5n64ArUdTfxNA9DynLHJpZjLZgtkClyuXvK8BETrI8n8a36kRRllpAnNH
tFc6RBHvChPdss0XzcIpbUxyf3fDj70zQhjEqRcVdO7DzujPslpzeYVcfpxLT7cu
jyGqJnh1/EX6IwGo4EI5Sp42LvB61mRTsU1UL5czJ9TW+iZJ67XyX81Zlamc2JV7
obTx8s/z0TcJbrKbjIiWs2ujiubeXXYlj3W1og1FFxesx3xg4lroGgEzlwBgcvNV
ykrsduwU8HZS6PjlACbzMhl6/dk0NC1LwbjFaFEcLraiHjQkWb5zbbf/h+Qj/+CU
FQVyOYUnwc9AhkCJ4sQMaLvXyh/zEe6e5hPKC2tGtrqNYMKI0Newlu6YN88SoB1e
cRnqOWk+j3PVTWW/henq07NolNcVJ8L4u8EQNf5G5UbOrz2/pcKDWFWHfpDQfGYU
9LmguVCiQ1TX+LPivVQtZrmWc+aPfupAWqnp9nppJaOBSPv2/nsNgkod/X9Zhhzp
c2Ie9M3DMAOnL7B0H5edtODnH/A9UjvQtddfHnht+Wwclc4wjIanqUdeQ72Ganqy
+J9p9TBSY5r9mKQ9h3kan5lOGgRsiCpVTzA/X9JamLf0+vTpLIV4kX54LxLQfdyY
s0nhUrGW3ZnEImHIqc5rRap7XvCnziIg9RDlTEh4ASNZT2qvh1B2HIA4RVRyRQlC
mqh7b+qgmr7FrS9HZJrVYy3yChjiD4NcmIKVGRUwacXMt1XgbMpqdpL6sl+yM/v/
kb+LxVznn+9AdMBdO3Cvk097Fz2nSr/t0dmVpryMMjSibvKgQfj7i9V9P7uejNzD
2TssifTCj7rxK6C+fWqxEDHw9rRYRUfJJRWxRQAA17aRaAun8utAjImGFDwYudxw
6OFMXQDlzbW6N5uf98dBEpfiA4Ab5I9sSoi7ZxCqxYFAlFwATFUsXHA/wl/1HFPz
tXwL62+Nlrhpw/wyiFe1Ubg2pS+ZNuxdsgUXiDOXTwC/7TFsEqf14MQXAELzZ9Uz
hQ3kNvN99s1UrDbhwisaJmjxkLbcEHqHX+uLbK7VPvJWyUoEmUTtG+EObKTcYPMj
ClF6b28PXjHm/vgtRQKLF894RHQDmclqaXb6ZR8B5+1nx1uxGzx91G60XJXipVj1
n8v7LeQcxOze/oN9trqhkhVaemfWgnI2PiQz+fMxGHhtUhbONCKXi8wY05ZJXRww
4IMX15GAwVQtJ0+/YB5TH/JfkGI8sByKO45rlDFVuy7Bz8g8lAYNyo4fCiE9H+yg
EIY5kJaQUwsRh9r2ZrIHZiaFg8MSwuOfs+fDCjHNQYANYv0pqWg+Gkw978F6pcuJ
z8X42cqL4ej91MLKpcqmtixog7jlqrE37+WURWF5Vx+6724ZN43CPnYgHN0fLH0q
+XV1oaX/dyp9LBPLzJ4+3diu0QYAVgC+Upaj238KaEiFRzBFXujMJI1gj4ze4MZA
Ud1EYwHgUwf7VIH3ZHGX+BiCkWIG1Z4exCC6Z7cDk6/0vj7TF2arI6Evjmvufuli
KQWc23msbqMD3Ya1kVoI3vr0z6P/y7qmW2Sk2wh/IaBq6jbCmnXPoMVlhFpu0kaV
g/HJH3bSjHUuT5HQFg6YGt2WsjbFCI4PE1hD+kLbEmsIbrFYA3WQ26TcWKjXpYlq
80b4lG0Ug14zEenqGOnZ+OckzQeBsJt7LGLPphM/KjJpN90b9S7WoJaXyAQWapYx
/xMQx8VdB3rWP8hhZLmcamLJIH8V2BZalPF2jeIfry+Maiz3fWjvlSDSk6kbEhMI
lFDuZDe9ZN81WWoQazhYyxCIam6bkVc4xbGtEhPbcqVJ4JO44iDMgkmiNLNAZMd9
/pMix1ub7BGsc1Q3iR7WFlboHKocFCZImgv10Svsz/L5FRhbwBMNAhOiLaKZXY62
0Fcw16z0bUKnco73LZf2uwPSPgEMYAd0AwQnLIuE9XLXPykmC52/suJabTYZ+r8J
1s7cvcAG/R3CzJeSgbYXu5Ot34Tg7AANqTvD6b8BsBZbOtdqPl9Jz2wQoog392jU
U4utAk1oteMn+9ohQQiLJ16m1/Grhyzhwqrpo5Zheov9vGCrCEn3H7W9mfNjc0qn
sioC4iMwsqL25eQ4x9qCpqsWN4+mcGlX8dZsXtfoB5lu1cKbtoDcyB0MNx9aUeC+
w7aLwBlbVqxklKE1ZtMqNhfE9y8vfE8fG/izmSzCYowyslypBRd0+yWf2o41X+gY
ikIho2fxHGZwIQ4pGqFFyfJQIjxNUkkdP5J42+UKLNV8CFO4CHyEtkPCu0koe9xO
PvCSUAFpTZCBNBJ/BtWwdWNznrbwtizj2fxXXdLyFHX/ecxoR8upgow8kvXyKj1h
LL1znzcvA76VoIWUdomO9hoOaTDhNQuCJxQzSPHhsby/9BsjR7IpX1SvzQ1w35n1
kIYpS/6/tLz5YeewWg5uqpJf4Ai4jUjvs0D4jpKN6l+S083ppK4guB0iqG2u2CKy
WeOhK+N9wpP9HCzYmRAqtE8HxNRzE6s8f7eWkFxwBwfjPmpZr+Qy8OaQ6zKy7lkv
hbbF8zcUK4UAXKCPVe12+frji3GIqs8dQaYos+bsc0uXbJTYzZiEGvUzmWrCiuC2
sas3hPL/qtwV2XbaEyde9GQ4u9u9PGBgy2F8koLect2ou+H+RJITpq2lvVo7osd5
iSsLMCValpebl5Bc54tqvWm2ZhGyRz6/tcJl2xMhMBbVf57TqX4M/fPoy9NWp0Ax
7AfHWBVNywQ12yG3tesWPY+qq25WFuFANIQUpdHoa4G+ije/4mLGBMGFRxQnH3IH
p3tGRPZ/WyLX2cjxKWlnQOagZnfsuCiEZzLKEMt1UvTwOj+edWVvq81FiMOxREVd
YFYLZ15NFz6rcNOdyvuo+JtkEtk1LTMOKslxRL0jq5SM8p45RR4Tmj+WqO73oTno
0RYjRyZODz0BIZ78ZNiavSi91Ax3apjX3+s8rJECe/eRjVOOHjheXpFDt88HFYia
urKZ8vohEZhe8SbEACupgzLhC/XaLKJ6ly/hiTteame4oZneqtJwjAw6flTLGiui
omPfqHqtGZj9JRipF1hOjljNhHHG1+IYcxVui1agmf+jlmAR5rX7umQr1urkNdfB
u5tORuo2EfWQmiOavcBjMQ2OBWO1hzKT0r2LR2nWT5b/H4eLbljggTilYlPYVqto
6E0kiHYHoEuUUiaaXgLQfHXTNohZRb38n1itJW9j5hW320Uh3Trl2Ht/ERW15Viz
TK4pYvycoL6Gn80If6tjxPvMdDdyqetZNxAh62ubsExLBagWrTgJPNX+u+wZoTxw
ZTxrxGQ8cYtYRhMgyCwP3QNs1/xagBxUkm23PUsYMKByzLQmKW9vhLUfCp5ebDPi
viFeYQNQGp4Z2td0H+2Hs26/M6RfmMgTfFzvTt53lRkiVzIWVQvuqjBaex1A9JnE
81V923hl8lJ6nKdBXHfwwH7rsTrcc36vYBoQeRiZFVzHTiIR4IFn0hS4zKWLP2Tc
ZFRcg+4kIMjmFg4NC4cWDmNhnIpVT+u7uNbLT0W/Ym0a9LWFyr6dHf7Wbr2L/xNU
qd2YxGURt9kJeSy3rJtVAQYhd0lJYrfD7ic/+ycWm6te0S9k/oIU2ofDyVM2i1yu
af/nwoYRRn6uKyDC1dw3DefmZt16QkFAe9N18YbkFQ72hBn7pyBYXTO6Aiclk8J2
8Ui/3gkCtQAoIGQp3UzBz8ndML5poGARXnMZd8HG4ZwjppNKRkGtLmV1jOG4OHsp
5yWe172Alu+D/lo7saE4/Lokkifo78T8r/APvf4pokCdg5WuKeGtef22rI1813VG
altCBYXhq+mJYnheBrS8+aXDY+xnjbYeQSMaU3e/4xzMVwDZlV/mcn+hNXvsnTqT
Mwdeyn2bPwnNxbmXYVazbhbMQbzp2gFEKqfq0w4kObpfAB2RSCIN8i90f20E1Rwx
Xqymps/E9S7f0+B8QXJ0qVzGJFfprTg+Fe7aBeEKfXP7PDcnMNw8hXO37CFvh5DR
yfLfEhNXctOa/sFl81BfKVHvrnGfbQ1ZVeR7VWby9Cl4g/XJGqtUzsCAePVH48Dn
WfBXXdhpV59zkd/f5jzRhIc0VtiiEaDpMnsWsrPNwvG9oy8/Yu0irajq4n80lTmS
+/7ihbIKDYnARKqGRZO3PT+rTektVt1OCTC+uOH0ZN3Q34h3IHHlfgQ1Ss8cSVoc
YKDAZbqWFIQwno1RF4oWyuhZYU18pO5qo8D82UOYbh0tPYOiedDO03w7qjuIx3c0
Ap7oxYwUVtMCAP+vb6b9KyW1W/rBKYoFvzC5uKuT5MU5QO6bjNIP/2c8rQ1RHYO8
vl94K7Y5W4Gm4fXblzb6rMp9pw7tyAHKiyuqU0JypnqNOkaEaXvov536oODBX+Pz
kP/vBZYLcKezK3GlHibww8fIOMP6iyP2xsdQq1h0q1I6iE+Ki4C/PkeKi0Q3ruyv
ds+gx/prb7gQfp5eHXhycp6ZYztxhe9MUAKO3WyjDXk6HEyPo7finvmcFDZdj2KW
218KIp4h01D0dtgZLSY103aH6MPPhEnvQDyran5OkHVL9jBbYtjuG80tJj9gGU5y
HbAUqRqeNWfesKZGyGX3qj+eInO3EpT0YuvU8m+D6A1XnSBZSS3ArsggfTp6v5Zl
r9t91TO5HpoDwnS9OTfDWBJrmIW6MBu92PhvsnbU23NF4DeSe82x8AZDaS/qiuFF
lrU6S4IZIMDQZMlg1zIFHSAorIvF7vdDPyYiAn5l6HlfVJnyV2dOZW6N1dhW+NCD
s/ijhmzfKqD77a0c53+f5/vrRugAVnzAJz4Vgxj9hNnKwPRxZzdbdMAaL91PbpO3
d7vHQvO0YOZ8/KI4MNurDdqVrS05unGjTgpqkXTEkg65QbJNFLkTshpRyOgl6mT+
EfnysMxcG5BtTaS3AuGzeKj4Z+dFwtTMQ+Kq2KxQtb/XCptBgsBcN/L6ZfMVICyn
iM0d21xAUT29+iUyWUa8dfkFBd55PHPbh6zlR0+2ZZfhTM62BcV/4ybok9BacHtM
eH1nrm1bWfcb4IRlaE8S8r+3yI6BCP9l+hvdkJ6BMKZKyvSVe/jTb1OvXtlEcVim
Yoyjsl+NSoSDMEDVJjKja2x2SMfTvK/TPpd8tn1I1sB52Ovgy4KXY14L7i9zaOB5
Pw961UKwlI4THpoCVq6BRipsKQ8weUUrr5G1EYmppceT3OF38b0NVY0OXQ28pdw3
w/OXqLFBci3avYv3/JduWNjTThGwJ/zlPQshZ4jBmYL/zn+QhH27iPaZJqX4FTZX
Zixp5drMq+IkoL813cD1lZ70t/3FLfOBcLGVortGchMb+ulqloo6A9fTQXNmabhl
FCdIXAsGnF4zoZ2YeMUkyZ6vQAisDp5o31fl7ELe60EYRzzuMJPZ+JUdq0HUcEXv
1YnZH2omu1ZddqjuzMhfr/XimW2cVgHLmOzAQGNT28eKjvaVj5h8mdY4lGZo/Q7a
15vtQwkkjfgkyHuvtdwmgd/6HwB4eVkYszI2Xa7BdAUrDPowb1eY/22Gere6Kpy9
8YdFWps9xXjC6ftWvep7Z6DEl0elMoSvnB4P5fziUc6xnR7l5RVvbYn1IF69neaR
jhWKzHjQoHeBGhCzCCRpTTyf/h2DRRLGBgHJA5By5rILPm/sM5nFlvnlQk/Bu+NO
+8xbev1AQTbdGyfbNYLjFBZSQEwUu2Z4G9JC/pBbu3L+kMUWVH9hrM9Xe4CL2q+2
/51QRJ04QirD5LdLBdrHyhJLeZZ2O1tyAXK7IP+ohtUQpi7NrAMypZkjOjEk66iI
VNL6sG9jpsML+OOILrCGjTb1Y1tsvpG6cznAX8OBRFRkd8XQxWcWLmPl1KjtBcZ2
2ZiVKjy1LCWXbSVr4OxY6TCv8ss/KyY0QZe+UcM31W4XPaAJoA2uSuzne7hKc9X/
UxXem+cceGwRo8ziGxsCe34pjAHch5Q5MC21ok9OZ1u0x9CCUw8yTbstReR0oSqk
/HX1abr+ooO84SL8xVrhLAsfRM5ZIOeWImuMG/iEXf9Qbj3tQd2++tXtoKuQa3al
11B0VuAdu+2HTp00eI34QFNSpVqUa3rsDFXvcXzXdrbkwWRQzzamH/iBdbAc+OBd
Y13MNDQpkjkDkO9L7GsVi7LO/Qcc5+BcSK7b5YyP8tX5jBii/W5iNZ+lSoTUhIHZ
n7TnDUG65sGZs3ChpKZZonW7jOh/2FTqr3xB6+ELXId4DprLDehEg8IfA6kNZY6D
52mRC9gjKNBJ9PO75JgL+0C1X/pEpXQrzqqHEuop2c+FjcTZgIQlb6U1Ge1Wpso8
d6ht2/xJ0f+NXGIzui6mLi2fvotPSDMLDVWXWEGXziC7OzVPI+wex6vxWuzbwn94
iGsQtjHPfxgLgwcEa3hf+5HxJPCZzQ6/2dqxf25a5nyBzXJbB+In+UoiyUi3Hcf7
zDQunKsPJ9LW1EwGV+LZ3T2MH4qA6DBFLr7NZP4dl+krl5BhrG36ysvf2ww+ORA0
/zn4rJm+UdnxLxhNmYR1iLLPMTEHlUqdXncS7w8/OYF/RNXgSW83RiEYtcLUQzUi
KMDDJF5SvuYddbzgU+QrbjXa0RTmQb0NKbe1C9M8QDB586ZX9rsd8Sl6PSoTqUh6
478G9I/jSHalPGxQCp1wxVLrHsb7moMO4kNRuyw06N186BUmM0eWHD0wIAY9F0k9
RFwcDUynceviPjERrdB+vLI45usyhER04lGhGR4HAhpcRFTJEZFSfs+2LlnO2DCm
cjYt8W5tzPYjhdfMMy/jz2R2ZrvaPaFftZzxX1ZyzAbRgj6y/apMYpNcCgB2Gt5B
NcQ0biuEr2fc1QNsO8RVhYoeujgSkCWj+/xR1hLWVVEippBQzKDhzrCsfTr+ZNKf
C0twWXFVJf//63keC1vB1AKcD5ziDI1iEHwrm+NjCai5wYkiHrObeyqCNhVz6+yH
nFfksRmuOu5ytW9Q7iwvEcXvJKpYi57bhMbXOckvLYCzP4T6btIguINqS+IR43d+
a4oXEhfE37a50osKsT2cy/h2ZegnOCb1MrrGl0IMAhkQg42rp0t5xYZ4LlKOVX2F
JATNsRSJTbLI4cRbfPsrx+VYNlpcxfu9xAOd2iDzgN9j5c58jkJi3gpgM34mDomF
nyFor10PWZY1aVm7YgxS6m9XaalvA8Wy9tSxIODYRkwUvlT+lRnKe1nzkSfSbEXc
JDB28KX0AZPdUPExso8CULgMgRaLw6qQtWN4ag95fSz2cIAT2WzRuUmHLVs6BL/j
k/YRSSyNZFgDBerR5PgaH+ICvfmhJK2fvMVytcxw5EjG1dSGCNX7ilywwri6ExYX
jGFiUfwHKdBkCSqcw0hhDdNB9b2OSKxEZJtsnzO8sU1iAJe+W0I/w+C+83Mamhwc
mH//KODCzhJBnV94vzhQt7NoO4UZ/ltGUyuVzDR2QQflTu7icA+55E00vzZL0ZPU
XoeLvWRcI9jSHUt2BLRZ/VjZVndCdotCnCryz7sLEkbampa12/sTKzbgqG07+gsv
fpUOmRVR8Obp+1vU/rqhF2wYCQbr/4HnURWpYQ3UL8U+x2lShZvxbpCSZmeoCdJR
9UMAWWKffYCluOSGaPx+ZtRUfHRF2sUc7aZkg7HCSx0FBgaXTKn2LdIcG7bPDncW
X85mjCFrzRKz/PgOBI7KBiSEPNG6GiVEa/u/blKlrxFK1yFtQVGUpu7q5kFQMBdM
sk+F0DcoT14U1sot+9wrASd8VJL3qmT8Hh2PN2B0rCbP0zVbpzm/OC6ejEiHQHdX
hxxDgo7RU92Av5Kb8cHKPknMnW4PUI531r2zCWqFe3u/5d/pMK2+RmS52jZqJymG
BLhs6fb9vXzQweOZ9eR+AyqwyEcdKJxDhu0kr+H2hWCO+4b9JT+eT2MPavfszk4n
mtEx0eNUE9GXillb45u4OkQZpY4XZYGy63iol3a7SmlFK+fYPL4frylIEonGEAXu
+0bNT9PkerGVoiN7UNv0vXbewFNT5gGf78UL1ix4jOQfQxmWW69suzaPP/Ex7fo2
gidRTBOt/4yZXXHeNafJEMn5+TDPWFB888NcR4yinOxsqmcXkSe9dHgWjL0nMQUh
Ocuhd5CGH8RVDrdGbX6bNt1i1Chzpju8G6rrCU3beW7/xL+1qjh4vf8XxpgnP1La
+cFzhpnQNILFSsVEt91P4KFxgxQSvWXgMTgOdiBdwdcaGoq9AGJfZgKHwoGsOZD/
wu1NlDTv1MwYwEFiE0hDf2582BC0aEsoReSFa+mVd1a8ZRcziFQdjNNgw/QZgPjc
6nJfD8N2/jZoh1oShArsUgEBjQdaqLyeFsBcVmfS9vmj3SI8neVxWrUJUOG1HFD0
FyheOCGqLWIWAfMzE/2z3wbMGvG+qzZ2YGIVUKeW4eJV7J8lOhvN9mR2vEab1aEd
XSBpqGeZq8NV4zdafYiO5Ngs+qbFK1ES8F0ByaiEFshcu3hbvR++xVbbzPvgKkTA
f5gEk5R0R036nfjdIdXk0mw5+2ZM4pwdewOO+WLoMI0X0fxLvJaybZBnTKqA+TgY
B79/9xTYtpI3/h50HHQ7EMuprekXhKYhTfbOKvQ7rKanCO6HVpFG4+u8XGHP4/dP
x2DkojZ4X4BTFJtBcOSEOOxDK27RnXFCwlp9hvHNx9dr1a/yhQPcUbf0mu0NYbfd
shcpnLdPthraqXXzR+T88OHhwFTWejpnHsLQVwYia4sEvl2H3H2CQdzooX8cvbDh
wq3KiSaIfR3ASn8QRqxtmyg8cuhJM4On5ow2LA3LuKky81odyFNMWiTp9aekpTqN
Pszyw1NzPZcmY6McnX9TB820+G5zP+IUrnIdChgCE8zeGcjwVlZOo3Qhr3vO+Oio
Yq90vyzt5O+e+LBHMIR4LGbxzjEqLkW2NiLWiAVBo7HvRwPCYfOzSBRXvTAG06jM
bmkrPL8q+p1HtB88OlKpkWS0KFgKHGS9SB0RpIZIe+Ml2fmSGq7DmDJoSQpZRRsr
AqEPAeJzuWqvTkSinHC0+iWz5Fhx4H9cCkJKCgpE0CuY4c8mgy7iv6CPxNe4ramg
rh3yxDKcrPTyEPKhFFsBZt7P7LALv+LHjsUhXg+biLC6cmc3/i2PeFGvHocBmt91
9y2G3p4afx9MHdfEamVps+vHdvYQYdvmF5aUaGwIAubodd9IYB9NhnWV2Kapqkhv
xtKk567lG+3QHMrUs7vE0Oo6feUtmCUcksO2y8zyALkDnZzfyT3Ea0VxQyoL9EeE
EXGj29MRZPAzFf0n1JUw9XNiTPVvFICIbInpOlk8DGNK6RpfjvOB/g4AOkebkjbO
Ru56cmoiJ4cG6SiKU1HLnv+ygVK52x0wqL1egsSIoKZukvoBml8jarnth02Y42pB
7p7LfkwxTrVJlYH41JFvfx+0NHmdeyZ1f7gcNnrP/3F50qDes1S2FOcMirhOQNHP
YXP6LaXc0tkwin0/oU561Vh32Tbs6iolRunt3Aw6dEqgSicda5e7VDaqCQXoE++H
v/1VKhLUAj8ofuP25Z5plY2pq9c4fkux+xDVD9APM/H1sjOPnUFrKjJbb2JUQIfc
bmh4tm7BoN42SxLfK9SwWjJl5V+9LJxdHJYFx6tFmCfcxNAc8nx9lvgMQumc3r3E
m0LVIRomoJQYiISQv2cFiLomcbwWjVGXNQ/U90qmvO7n9waIpcKhxiEPgvV5FM1g
6vEXNsuiKoOXxMFAAOyT3Ni5qELayBfXfu9VmOj6AhvQMR/A729eCmwmrdRMiT61
NlMzYy+VAHy2qSXXeQaPuyRtqp35t82CsX5+cZpNSWZhgwbSLcVYulscWoHY6JRC
I7w1dB9vyU8EkR3p675iXNNVVGHrKd9Nj9nsGyfDR8TOu1r+sW7Kb+qPIM+eZf4j
ygAqnRG7sS9QTVtwyKofGi7FC9HAUE/v+vyOL/MqXzDnuhhqpGGCQsWV4FLjcPHG
bDW+c1DtTiKRrpPv210TbU6RIVZcFz9VHzbQMs0+TYYu18jDagAATNVwU7VEDrFm
jvJRgZro/6xPoF+FXCgddbkBXQoyuMCMXZpoCXvO7FkiDSxbe+AcsKAG5p10NBzy
v+Fhti5xHFinjfZYv3ILsDxGot7bdwf0I+yzHioG7lhf5BwxjBjJX7xGP4DHpqov
nd/qf6UmDcu+trTBmMlO8GChnRLSptzSUthqi9P/2EpyRXlN6sIO12snPdVi71wa
UsLbJB4fX4+7TywQ7eV0fjdn8cPITVQtJUDR9SHPM0sTAzWH6LFGboQjudmHwGPH
GaGwjIHJDiiodBxJRKPSgnn/RZYpnlzkM/CdJVmmDp6ZeTpNH+fJrMq2t40xGzuF
WDa6lPYgP0EbGZnmLlcUst/EhVHQFo0PfFhmBP0VwgVx7uDFYQSqP6M6mb0vLUiT
U8KV5erjtDVPwr5r7JCmhe+XKZOjrsrfb1K+egMt31oN+vjIu08jclKFO8dpN3Lo
NagVcZmBTPgoNrnO05aEZF84weZJxkqIbJ4FEOFpNKS2vtHERN29KQ3I0Xiqu90W
Kt/0GpxSYZSCcI/aBVjiN/9AxSM+epHP/eS4EPqEvE1o5BMy9OlaFlqPYz0wAfql
rnl+w6OzFdkONpkc+w84HXDPQuknjkDUTv8lxNpBvBCIk6T90DaldFIUQGbGbW2Y
P+lYR3vRMSATSPVMSh9FMYPcTeqlpDV4rNJJF+nRsWvup37uYIk5G6gaRmJhBsHc
2mTy4pZ9WlRVqRmZz/gb4ESyciwPoOkL+EnswVNmEXtiGni2IELN7A/XGKk7kTIt
kzgJXzmHiuCSgviF0fqEvMei6XANmEEUaTDGf1cX+3F55E0nNIF2MD6lhVPCULBG
JBU1zNajLdKnWweHp5Dlx1I5iwNbs95izYrc5i5A7rFETQc25RhvZeKzJUVTRYy2
DaVdDkeVXCxRmjEEa1gV+JpMKuk316Sgt6waLBnRgBYmExToNNsm2ms2nu2jgcA9
kRkjuxGEcSfNpf2spHDJVnpo3Jc4SKyaDnd28s6MeTU7Encd9WE7vhnOJrTo8yPq
2YCO/KcHgVaCksnvCqJd4rGrNp+tHIC7XGHi3nOizMV/ag/+yZmFOOmarv7QaPzI
j28GlNM87zk5GK6kbiZIIzjQ5azfjWd/HbUjTgHTCFqzsfsxkZgFTE13Wg+B9uwe
G2BSJG1aJaBtlx37+e4yYf3de0SidLjUQvrXwEBWhgKtAl5rfKw3utukU78aEDPg
iZ1GyGGADuugcAOG7nsi9gb4wu4qUhC7dreCREFXbNAmijPv1YhzxaJXzS73A8Mz
lTQ0XT8u68H2Q5JDBm9/R9z60TIxx8Z+N+/f908MFzWqGwTjyOKE2eWDjbSzVTc8
Anxh7JEwCQ68gax3Qv1/62KwHXOadhUf8OBNLb0yvRJYr7+tZk7BQH4jKRaXqN/m
1rZLnLILr2rfZxhmAhTwsjlcm1l/0+GN2qL/338L9bHerBGA7iv6g1ywKhXM9T5P
sw5Xfocu80xMV/BV3d2Ww5uazaETRNaJNOk6Gpn2v/Qvm+PaSFWcnDuRvBrT7U2N
Q0QovYvVD3n4XCjizOR1f9Itd612Z2LOfM8Qf13lfikLpS+MFb7wSv1vK1nAOILs
yglgaOO1FC/aN/qrSaFBXKNtFK/zJcOEupTvWvJ35Lefr0k/aKf1spqf4L/lKolY
ijhOmuSSsW2XkOwwv+hGnRiHF0UFPfgnk9CqkNeqLf1JqHG1y0mEFDguNKUjtGk+
YKdZsp6R/haKNkpsQIFfqnFJTtU8Aty744HTwsex7OwYyJlp3YtN7KJZedA+sk+9
kot4FNSvSUwpl9UmXaumM+Njy0yJPMVlPO/vKb3s0WCnDrDj2tHqj4c4pytxr88T
A2rbToPubMPqjRo3uzc4+oU7FXXbFHxRd9RjHBbniu5DO3vV/hcq9Ir2RAY3C4/5
tWesLZPHBsEYPxXEL3IsM29ItXF8mYvMD1G+LMM/pcNSviaUwv9L2yN8ug6S/4oK
Gf5yiJecyIuTZsuJl1jNhUE7zpKBaSPbeEpBTtsrZgHH3ZfQMUn8LJ38hktbdpbE
9SdemziRZGRwmF7y5S9jOB4NVmRFEPUKiTd+pQAReqPRIlZc1y3FFz7y9OrDeI9n
4gYQR+7b8CrZWFYI2u+g7h1C8D81QPwiZz0l/Sq1lWcHQz5py/Fvs/tMId0A+egQ
iS1/ll/eczwvSreYXjgzH/aIuWHePNXfHN20SWkFhb/dk5BtcCKD6hRamufIqhxJ
RdO3fyFzh6AjS5AyHpnFBUhjoRP8pjRTXGI6oB+FUEzRNbgJNRZhWfstdsP1R8Gz
SImvEJ5MP0TkJDAFBNXsDd82wWyCNsvQIKaYPJJTTNIgMKX1yDl6fRXrfbsFOxdw
v+EtaRR47kMMQjwXCMLn7L+yCKpi6igmen7jOfZ3qjlDqNDfzctiV/+MhrfwH6h5
9VzpN1stQk5WC2xbHfymFx5kGkf6nl/N7xnwQmnpGqT80w8tyEmH69JbAoIWIH/Q
5oPLsoriFUlEGjcgZ30PF7ZRY7X0sDJEuGCzPwMsZrzAOhQ+kBUIMys43fYB/ZE/
rpK6hlBjojv/YAeIVX9JbMZG/8RpcI2e7E/WgbC48L+uqkQL8BHgxRkK4dbANcTO
goul+sLhOhFQ35UidhjRGLusY8d7nudVNpNlSd2uQVHyutFPnXysoVb4+Fz+cRdW
SV4vMMEbzKOmnqp9d/0UTluGzcs/N2q5nJv2/8gCrUH++UsIzKfrlT4f1yNnkH64
TvH8uu89svUSzxJvDYB/OsWTV6GTxoEEz9T6AqI9SpyK1q+RX+k1m/vsuhUklsug
bWgDOvSntv4u+Hby2ZaksKMGJa8KopsMe34cfWnPrPiFNbKmwoXUbBGNnHp9Fx+E
1sefAxmRPn6GO9aR8heh7Jp14GqAyXhtsxdS7+xQfp/e2nIHMBxqJtDhdbeXbmPs
LTcaVZmsrS15sYtYybV7CzwegA/a1cybyHQsyNowwbweftstETUBArk0in+WqAxw
0kTf5yLtepeBtQL2dgDqhQeQbytZ/J7K8RG+I6PbBS/VSvPrUCHLxKftgheS7oVE
qtapUknYHd5xmORX8lfHjLnox0szIgQYTEKGCGrnqGAWY2VvbpWf+4FZxhFu+On/
8BoX2zEfHnlKDILofm/Yp7RlTt5/RPK2bWXkvh0VzMKKf1CBZGzLPkFoo6q5D4YH
8KZimIifK2vscEt18smLzZCN0Mrp+/KsUHdULfuOyUtS5UQAjqkB9XubP78R2uCW
GmLXZaDivmJDqzz5bTuBJHO+uEIFF3MBkVxg2pMl3V7U1mwE+vRii2LgbZkmJsh2
Ve2aWyRrpZtP5yUp+25PK58/4LcYi5pDJ0ovKH8Nh3wFGflzi85nrmS+8XdDSjkB
EFbq4inbgEVzdWGzVPcJAB8EXcb5sP7/PKfYkbE9FX7ZSxfO6sw6HA2sbcZYgb/1
gx+8qBkBPqZt0Wzj1N192hdZZ1iaFILL5CgPfB0gvxQDPGX76Cc8P7wtlp+kAPMe
zXrjABErwcPVVdghXbQgKSCUUnknBd/FYP3Hf8oQ/WWyR55tw/V5OLmB2RzAsRBV
8SLBxgZGVx7X3uI2gQcnNnTE5yfKsnuV4tSaO6pX2do1wo+M8hHoL+dQnVe5VdJg
Ckhkh/DAmQARi8CQPw/sun8Lk0Qn/JtvJQ61NdECTMAP2gYvYajA5jz9tto+pTbO
5z0RUIzUTW6JFjPsSVwOOAxPkk26csU7pbGcHDwaRCQcU8X1OEw0vSry7CPRw1fU
q6ceqG04w0fZSy+Gie4ltgIAn+5WeHAvijCXutdgM4iu02a9N58RdtFVp2etAUaI
z3pvgC3D+9fIwU4blY1NI0INArAZZnGlklPnLb80jVm+ZPeaTHyEYgsk8ygQfdEn
LwiF9D2fL+huMpo8d5aN8c2tgxupmz2i8VQY107dBYWq/t70qY2pXU/tggtX0T6u
fy+RS4kXqpyG+QtGEvGlKCov8gOnkRxBCi1bpJuhhVUH4/MOeeycyBv+LL0jQFH4
Zh6lH1f2+2f2mMz7YAA3org7A1w8zIxkMDwDDHHdeYHG+V0kZfv09yjd7L4/xW4+
STG45S6vc6HOPugGxRAW63A2T/Da9Wsd/wg1tjoGZwq88B2jtXiF5rHFDvVSMj/3
tulCe2U4FFD62rXBVXLGZYZcOVQduQd1jZcLN/2OADXP2B5YrY2LElbDEFX+RIxU
jOPRsW2ki8ca0slSoG9n1mE0e1kk5L+CwXI8/YmszFqmOmKO5A8BVFBAPlobIaq6
JbS7Z7Qs91pL0HZy/0eYFjYyOIpBZ6c1AKuO/p4jZCjDMs4jUn9J8TT3j/e/Ptys
6E4Ei847EpMW+5P+7+sca72w9iE8OQqGK4vvdOkHqiWsE7PXcpk2lE0OnXRyd+DA
HOHTxa5t3piSlXuow97gehDbzB3d+9sHTUicbTaJdptzBEyMeiOgIIC0Ho7Z6Z0P
cQlmwQjneZ7iOLI6fx/lTPiXnzLqnQw5aQTWNjfss5E7yOnYOaC4onvIUNZZH7Np
q3Ij7DpXleGBSN9pN4J6rY8mXFFFHdJJwjUd1wFuxDW76S0dpad6iNOAF0jjRr+K
InuArjyFtzIVDc71H7/qSvpUhf+ZqSR6wcPgnSZeJlE9D/TDOMMlwhES7zApqhsl
Q/knpxx/U3vKvw7U3gpy//mjyaw+Y253su/vODg1Grnjhq1+8nrcWqAdRxTfE8Rj
SKbZLikivXoTlHl3/fCEmVNqne8mHAawC2Iu8buMDBjpYqZbYEIKQrRCmCM7MYcw
9Qu6xEs6skvViCFXVi6D9SluBcmpHZvWZuEPK/S5TLntv/NB3P1vJG78VuL12fQl
0QZi/Pk270qVjXDNYsVUrkHvCQjengJbKoRcrsr+3WlTM8QSklm+gASnfIUc+LCM
VUiVmuyA7me1lvJ71dyM2f2qn5pzr7DuoQo9UWXH9WPFB9YZugSbi57zXfbO7zW3
ulvJSJTz+KjeDgW74Xh7Gl8rk7SErsv1hzwQsBTQsGByZeYofTox29kdcu/uP2aA
y5ahQWAmYjiB7FR+uK6invekngp4pl9/agEulzJ7QfeKJUu5m0g8vkvXQTcBB76o
ZG6fIVdoXTtaZ8sx81cz2bIrvSe8m2D/ssD3Su/Xfutwwd930SsfXZQ5fGdFBhza
gylraFxU/ESHnk4uiWGk2ZyCL7AiDQbkUa02PHqixc0OeGC/jdyX4OuDS8RSqMa0
V6FmS/04s2pan+U3oFpatWy+tzfKZ0Q1lshb/Q7w7Skbp0zdw7c4yJUm/DlSsh43
PYDPnB3Sk8YhYgRC4zU1g4nDkXiQWBAFezCkGoXFY+950AssNxzbzGUX2kutLedt
qVMc12hO4nhbK07klkbxeKNZMQXhxQs1vb/tuAJdCD84cdysRJWLgnmYLPVBGDPL
7nwkxAWMJrYUUViagN38TrMDjLVikBbCB8Ueo4cQWWK1ToypYU8myr64Swo+9HcP
+wr7AyeNiYxFda7ILdJPWeo3wdWLNVYTKjBFnlg6ARytjuh+TuPlqCk2WEYmxuU3
b+RVxQHSomKtd6Gq+7jtAPeRHLrd2KXs/1HflQNwkZXY0An8OPteFsBur62pLQWX
5Xg2nr9JMV/FyacruCGOK+wJwWcMvZ9Rmfh0mE4Vp/Hhze/H1n2xVj9eeXesnfzi
vf2xHaSb1j2nm1bq2esT56bYWUjV5r8WQUugGYMOLveFWCoAIrIjmvmBFEJWIkYz
gAmLcOMKr0F5GdL7zUSAOBaVLJcuK+DDMqt5sDfW3gBEdQ0Vvmy0FkTD7X1KOTRq
uHf7totamrSgcd2zvTV/CUFuPnptG2W5cWpjB3pXdRyBdnnSaGzUR8F/YNvWiLQL
7N/soujoAj0uY9w8MnYEVPo63wuUjHylJhzmXcMT5MtZfW3xUoVFaH79I3w4sKs1
Bfb7CbgSP5SJIBgpZd+UfnL/wKXa7AAnuEebdbNf2Njkbz/UYMje7hMVxQJXb8Y+
cfyYz1CQ91iVYmH7vK3CQW1mza3uCiEYTtKTqyKtEjOiLtGhklgsOVr+byeEK8A6
+G5ONNMshYpgAVt+YpjrdTydh2yGZZNIQBo+Znb71S81Wz7ywHdvOC2tC5JbzydU
ODI5+8vk5xV9P3Z5CXiDp0boktWVl+NVqzO2fs1ky/+NkW7SlNe0ZYU2RwL3utD8
HwvAOsiwStFKgduS9NJ4zvCDE9hJ0wgiWgj4hhSihsOd7aGJbV9LLYePnPdho0Xx
Loxu6uFTZl/GxU5xsEtjGAwhXoT8qkJT/RITAhYRFDwAFQo4W61CMpiqzSwnMYVn
TdbUlQzSuSL9U+cYuQmXt2V8KNX9ZOtPe2hRu2nN7XBWPgrG+PK05rNGcvlS1iSo
pzurJa2plpdvWQolHAZLnvqT4r4d0ubJ2czaEOdHyhfCOKpN2H0o0+A6aGqd5Ln6
UZyFtABvS8qhK3et7BNyYY4UqgFgEyiARHHvLfe7oUB4wwO5uQKN6rE7OQ67wu5X
BKrWDdj0pWTRiRihwSbtH1ulWipzB0Hz0ptzlJ29hcse5kJr+XL9YP/jJgLzz1Ey
H3PjsKvkhU51kZ0VbOpiekvSs/uaMa447cvGE6PfIoZW3sMEMLB+LQzoaVAto+RV
mKTsq5YKDL5bRia1aRQ1KM9n1ZXtTmryUMaWOnd+fTijLXlpi1vF6fUk9nVhPFIo
+iQB2J+1gUdkifrycBcsgIyzv3TSeaR859OCgPEThUCl6tQn1FOb2Ck/R0M5hmPG
szk0jTtQCnWDBtcqmJVue3wtwp6oIMLbxgusXTr6c/xQKtN2qaZZeHl0fvnmiigL
Lpkw1rPZTaJ8fJMgfqttRIEwAt9J5x9PCBfdeDrlBWwXMrL9foKUp3mH8hKB9Sjd
QHi6jpFbR+atAtYJlVXqaZkFv9MmCzK/T7od3jVVJtmogzqST4Bck6xNwM8nqhdn
5X7rmcKMAPFNeqoc/6UqbQCRzzaIy0DUlzMj8j7bUDI2mM6UxZs0cFF5zogpe3Fc
ZyvYexnVHcp7zegaLF5e740oslVjve3ttmB9i2qv79bO4JY21vUiFXm5ZUFl6z9B
/tIWe9OiL1Q45uE68Y2rVLuo3U/JqqnXQL95A+HHLICjBRSVUbnAwTrojFwasdhj
QiyANjkRZ2FkNBdfpfycJbF7xKnm8jIKzqXKgVNvP4xiikVR07GFdH/BfsDKlCTN
s0u6Mk8YFtRxEU88jaYq4TsT+6SR0+IMM5qQBxiZnSgsiKfC/5aewwA8zLDQyv24
G9IG3e16hnt0HzvaGp5asJN5EyJkGfESfCvuxc+LEy9UxsGMyy2oIADmhFx2Bn2X
NF/rSLWu1+Df9XltHclt4eH1iMLdviAx6G8l/fjrMnBl4DlOmsP8v3K4ii96JBqw
+WixphZb3Wk++1S1UGyQu+W4WW6cX+vqrTF3l/ldD/4tXKHXSwQY5bpUrIv9YGrr
cTmXiL/0/VMmyd9Sf/ra3V/QAosb4gPe6wRP5NVEisYzebeWiciS6Wq3BghqZoID
VZ6tX2A0MwymM/Py09xSGoVLDs5aq/8f7pjzKVO+s9pvv9sqmFRgRnPUM63zZsI1
/rbKLZIKyp6AU3gk730gjEJ5/+OJa8scNtFc+djI7/IJnqTimtqvLfARngFsT/lW
yRSIUVefLnRc7e4LkUXrZdYonBfSBVXaIIdOAOxyjlYuJZv5nBquSp1yPK95AqXX
7MQsdTLF+7mv0add+Q8sAHFtFJS/vWwVCgiwvcG9yL6ZzriUlECrVU0HhNdiv76k
QUKG+umh3e64Q4pDsBAofCHFcreHi1zyx0eLMM5XnH5UiUwstBBY5m9mCuD2ph5M
IxrAaMGgt3ve6XoEggorRF1VyasRjrLX7WYaSBZmCyaTB+dlKZgG0wZg9Sbb2hvK
JSKPHQuS8o3ZbxhdLkSpGdGsXjwyJIS5St9qi27scN5VQ2b6dLQeITvhDqmLphpw
9LkOeywGc6/RuLDbfnWMRgQ/J4AnHzDZOxsiToEQgf78xUNVDgYKsQfz3VU14aXI
a1e0ZvMVdWlxmJ5Fnp6w3hIyYfDM3HL2y5ryElc+PYIFAlTmv4BWCmJra+Wo1zFm
Hr4s643zRoyE4lKeYKJPOdLVYLmpQ62j2RKLhYAiXrnqwlxCkxiQDPpih/GrHP8S
erL3LirP7lxcqltRaGQJCIZzzmuzhzkSWdi9hFoTlsAI1Z2AZ7EfQjdwvcQG6rPc
oGrRIuZ6Hh+4QFjXfaD83omtg+ew1KCOGVk1D51ffDV1tSqAMY8i6ec74wXLQcd5
3lSUc1VHhYxCAGffXGo+HJhX8+qOm4vkthT7lLFdRFrjPWfDZXFPqyFgdUk4Cx2r
nOherEDVNkVRpmdntuJrMuW0ZXZGOZqx9cbZ6EakPmHjtKcSfqJvtx8+tMm+DZUC
bcDXJ2kb9eClGZvhCf8n3fsDcC+kUcY0Uk/xo57EdR5r2kk8HaCzQVQOqMp20XyM
lsp3uaFRo7uemDMS/BPIKFOQGwBsQRKUqdcXxUnV8QbAYWhz/bQVdRTqGlPibDm8
SqV+UyCpG+Bj4w1Nv4jZhgpsuCswIbmcmYJQ7ZT8norU1D8QV0GZofq/+50mZ7yh
itU3vQScrl5Ec3CieGu6y+NPGMo6wra1I26iBLFrnc+qKHmvliUL7Jmguc8jbonQ
oT+LwhQQSK8An+FnMPMFzxdYnQHjAR4aHcUeDqV+xNv8dwEtdLmaiiYYi0ZnM9FY
rcq8dvdjwRkKtnDmsigI799CE4FGLdUuTmpsg+kjWA1/SKuHqnPggmRjPPASXkoC
4a3OrkAVbkISO+kfjdejZpuel1918/LstVfGRO+42iSgmBuB6t8rt2kIDXwmpfCf
g62HoCMApDFLVJ/tX94psqXo2c9gL0gbmyi0CtaV23PETHQQj6STZBBhc5lhMl01
DPHmq3cHgtDWomW5L/3+0P1N6Hwk8AklJUUUUd8HjMeSeuC1ReIBoy0FTdTRM5nx
jVdMWNLYuSwBVvwDrPLEUvbb3Sm43HkS5GNAGTM3ECDek2ImFHV0CAMSQ1YmSCf7
d7L6sO9BMtOogw2NeEyATs+tv5dV8n8nqDYFsfwNSKUcijpzuyRk8KZE0eP8Mwb8
EVwnPvNgdwjRXWAdJRvaXmpU3KdR1cz5a7GPMwypItRX9nOWomRCWrGvyGuc6hW3
2LL69W34t0UvYdjMSBzXOsAbHguA0f0q73kAk/OMthu5CNbx8ruRQlY7FOSxllOu
XJ+fbimLht/MIZgz6MYJuB6Uz7uHu/li8lHkUFQtyCUCzEtvF+3q32RlwScmueMb
IchZmCwpKoOHavE0zEWV+Rg2e44q6qHubIgpDp6WbPmSsHX1kOps269FgEFcOlES
V/UaTuwPKy8ifWzKJm+m7FGSVDalgkmQYQfxD/VtylADhOWkQO9VEHGvDGz65Lj1
0V1QodGMv1ric0IULpNhFeYFlvEXGN7OuB8rgMzWHsNLSMuIhyGnTFUQ/Cbl+Slm
Qlu5327KODT5nTcmhA6m0FUbNWB8yI7TrsS4+PsvKXIeYexmOSTwiUHdQDj2ztjY
uSxZKy/kxBny/E9eHIwKwtBy1Dg6QueIFnmA3can2c3eJbvRb/qNdcJy3vBA8lxS
sAyKN+6QJLXqku70yA8Fx98XtCC0oQ9GCRflJkXBft/8axx0POWIw4Rf4As1Fgnd
k6cQsp6cMyfCfUdMfM+/JjZZP4Ux6MkmldGpm51RGrZGBR4jSzTkzo7gWlmzRuW5
Fus4tC3OBWzMYr5xH8Oi1PPiPBW6AuNHD6SNrArGfiKjxAHWaBNwLO5890ttCnh+
tX84OxjsvHZBNG1n8Q2UzYokZsGWA/P21ovasESM3tkj/gNjTEjPT791tg12v0wJ
K3vE65sww/Bzx7laAQn06Are1twIUpijakO6hvvdpwm2HJBOw0k5i7JAxz7VWxUr
kw/7hRs3TrbAfdbetMCNffHe3BhUrJgtv3hbF9DYICEeNxFByHZCPJdwi28kbkJx
PwYrMNaOQV6XxYK8Sz3UySXfjOAhdpfg+6Y/0qpWprWdtEk7UfE7SJWkLJne73zl
sRAoQF2fxYVet6rbw4WM8H4okxqYJG8A+vXddgV6XmB1RD4izDmTp9UZW6aSwug+
vQC/pU5vnAxYXyip7rYAaZWvxesGQ867/Ugj52nlGMFNzp/T+HLpKJqvPlwdOviA
vUQBGVwLwubl3sUY4kc1y2hNzaHhxy4T3ADP+nqjhJaiDfmFaqcDM1G4Lz/VddVE
kH+kAdjN/YxjzxCrjdOIIeh84NnAEG5Xh74b7Zddfuko51CY+f3Q+rfqrs/tIUzf
X0pbasI2HO3BtrYyPTwD4ogozPz9AsqOC0p4JocX+7bNHE5ZIKw9b3oVpW93+lz5
IDmVlWkd4J2WC0ekw5/6OaSkapKeorIzbGQ7lGO1icFCbxqwsT1jK9Yw4B3qxU0L
Oe78gvTKxptEvbN/3tj5fClNloi/n5oxnMrOmWwKMmcaq8qkfraW/0wJawkbosgW
TyQHHXSPqyGSDwrKurlf/MxghJY3KFJWGLc1cqqE4xeL9+FkwY0u4iydOcaP67pM
9qNMfQIg+ZhUxcdUFfDir9Dtooia4WBeCM4j/+531Md/GquC5B8K7KDRuBmE5AFG
bAkbW3IzaOH1g/zrm9wGE4PPxbDFRXh3pxz5UFFkgABWZs7lOwfOCr2K+DStzWAp
XECETttneHq+mnma8yyd0cdfEpaSG0BRIvFWNFU0vPPCVSjzIEgyYW7jHjrAE305
SKZNra+d3rIsSs7ePV3ZWtkJk259C77HiOjFQz9ODCf6j+j3/TF7n/USq1ZliEBi
Y4v3fEIVEDQE+0p0UvoRx0/0oB9vRjcttMJi3vIe60FXY8bm715mW+3o15pcL341
ePG8ShJYDuQynVTwA8absKPE72bhMTIbDhimlnitS7ogZEgRInNjNHWUwEcU2DJe
i4C9dTmqBpG8+P3EZjnJTV+e6KygTEdunSlkPeJWWqVNfeOyrD0XihBXGYKUjlY6
1/UDQ+9WznjZixwmtgrmYWrVca4nUouCJ2kDNfpAPq3MSBAlS9ylra1/wF8NAX99
o90J+0KhSa9lkW28S/YMAJ65Hs1SnRf5fBK1KOMMdHUa1Cvojw29HetbrIwyrZi/
gf299Jlg8b3hHx6Q3eGVYRebRmpz9S4JlvapflpbYmdnVPyDnnxoUq4bJ63iRIkv
ktEK8F/X4HhHZ+jGSplRiyMdNS2LdVpZqTZcx7RS61DGd5FcfjZGsbC7mSK/RSNv
OWtphk13MrV+cdwbmCZfO0KMCSVdIvnch9rwbiiI7DrY6Jz4fLB1/d21NzjuhXe0
DMkil+rz0v9ML13taxGTJvI0kfSOw1UXb/lA4RiqtXcMn0HdtRI06FgxeaSJnxDI
Hk3jdcUO9OFLLjwsZMm5cE4QuMDblO49VQIV4B92uGXCVhQdHplUep6LQSt8dNk+
Rn4lCMDL+Gd/8I4rWS3WGlEw0u9UW57RHtbmzXCvqAM6acoBPE/yXGsYSAyZRy83
MVF14u5smQ9DflXKD4dXxCVgEfy60uw6OzlLVsurTTMeXX8Og7wY+VbroR8Vl8gC
5HXchgYkmLgQFLUbEdyha6BApRp+SAhAuH2SGq3aupkrrytb4mHtsFDQMt8wX/gq
E+XpDZvc/E2LlL6XnIyqB0QYewuf7qZFiEPoxQouJm86g0Yz3Lu2gl1P3dG+KziP
bNSv7uLEJTK3naIIDxXmQVxUWP4c/NsF0IGuFDLqVr70FkLfr8PMOAV5myhO1qZS
zdB1CJs5EeAFTEkUBmQrHWfYMroSAlfRCsKZfcHo76RB6aFUVOLDMjxFerlgsS8u
7ERfcXDaZX609fqDxBV/y6Dmh2JgSKyq2iv+T91aJ5/c9GHTidbGyufLLCCtXSu8
Mx2wDABlMGP6IqC63Cki7vJyyoN6eg2WUuDbrLkEl7UDls7wwpABu5gT8U+OuNT6
u9f1aa5UhuDMp78ln2rbQ4aVbp/ksdNdgJO5Fti3OfgpqX+Vg3gzLP2mdCf2KbnX
fumDgiSCg3YBAU1lXqccf+YiWOguQBQ1qMW/LSTSAfP7yGONvQ5mi53/mXZHGMlD
c4PoTNlzi+4LqYfnlWYWm1wEUPYKjdiLrT41kwkQGNDzSsSHzpZqvb5N9Bww49kf
wLLNczYHhbPnwfJDuwpiB15PzYum+ZkvoZE6zmKCM5C1XIfqT4cdA04XTmEQnaIO
5EaFbYgDGrlBYjMfQ59KWuku32jXNnPRRZNJL77ZCVu4kYYM+ECqytjAyV/HgmpI
+R7MmW4R0ZoutwXu0bOaHd98T1L2M6Xbe8ySFP6ZgW1ggDopYZt/NK+mZjFADnXH
82IxQZzOrJz41wAPIYTGNoNfbmKcxAlxY/7jFkuaRKrhHFH/Mf7MpTybe94PNSYX
DWPn4Jl6hsyskpEyXgmpvfoBQVyNcSx6P75XOO/wupguRe17sQIiabYyPoUZjyBR
psdHNfmO9R3nt+fm91GFbIsvoawwvwhEOMGYbDF4ndA0Aoy9oxQdPuqeYppx/wiM
B8t/4nqzDl6lWFdbLrS5tSADJ9Ddr1yfG7SK7oRi7EgeLCtst2RxlmJmyMXEVYX3
as9GDHgak+50TDHBznndPViAudXOssyLmyBSNkOQPlaOQBlmn0fY7bpm4Id3njd4
SMgKwEW1NHW27oETZLb2GGg0mLhnj6ib2tzz8TUQMcQZbmCXxNsoquFnfwCMj+op
Yvk3u/mzXmq0bFm+wHPMSNkbDFsTYgsoKSNnoEOqPbbL+VQHMcJDEhihSSlCTLtv
wrXFeG010UO6sy2W0juaB2loJjCEGCEl/0p6WNVfjxu2qZbxZeGcGrNJUSEVcR/l
hmYLeWsUs/+bDRWp9Qc18cbLVmtLZb5+DxjBbTJBGTh7wNcdb6rsxP7dufyCYeyF
lTkcDfrLcBUqY2iPJRLkNvfLaqlnHKId81OIbFTG8KQDL2UzpUsF1DWtyIGnisv9
JQC1cWI6YGqOZMsNTHNG88wWwHbB2YntoZUeyL7oCNculotICsMJy0TuP+F9VfZ6
ozNs7Jx6Je73ILzSp13sTa7Gg9AMmnOedjW40fNqGoUp+p0zF+Sis4F8xCp1hfFc
T3jnPG1kidlUHMLrAG340tL9JIcWNm3u4Lhv2FPDBTdEmU9P9ReoXyBvX7woAHbn
kAysqouRTr5k6hqEjqAvSkXxZExYHJnbgitRfIXtmpeyuQmBzjT/gN8xG+MQmY+N
8y0o8R2qFnhQjPKG32YOXgh8tlo7qjDI3G27YgdieIDayQuW/wKGoCIMpKjehr+R
/vmMpfmVQBZr+gp47QEowxGembtYl0WohbtyG+L9Yz8bYvKosZ5fK43++Po3C/+9
vf9rJjXvcaMFv5dKaaetcNpzfudeUIr4OeldH6EJB1opGMLV2MDvfV/xKywtU4F4
ZpRZhEI3y4tpngIsGO6245Ss0tpWaRHqzcllwlHbNPK0a7kpsVYorIe6yd/CH0Ja
EjzrU1JHji7QkbBEpajcrPUtCnqw90znZhPybPuyi36vKMxkB3gqjBdt3t86VXQD
SxnUb7NVPoZwghFwweaWAod2xrcUhEig9a8ry/VdiMZih/kFdK993PNytmkk+bc/
LbG1zTaSTc/zKF29XCEeYnbl4zR2rFeJ+5r8++tl7uqlfdCkqtRsx3vuE52Wmyc+
RmKcPru9/akVYbAPaTm39w05Kneu0DrxyGd8fDolyH7qc0yoIeTIqTqLa2oMXyoA
iBpKbgBR7HBbnsI5a7iDxmfThQT5PF9asjs6qWuXGWAo07eQ7km9yxm4LCxDQPk5
xsuf2dKEvBn3Fdf2eTaHMIxidJkTkFA4jHyNMkn/dku20Rsvgm5qmt409XPNFJwh
i0OCbA7iem65dvv9NBDDM+3hlEp6OZGhf4je8mR9xypRFGhw7jp8ISQnNo6/0rhF
iAdVqLH87StLqMr5yGAhCd706jCbAnDYB/l26YXI1jsL7RgpcWDtmS8zSOM879nU
Xat91s3GS21ys+JzI7cllxS31j/95KME3MJlfgChlJpA8ndlLiG9VB5edcNismDz
NSvTpD4sri2QWIrlbnXqy3LJJ6WCNMv6E8L1x//7pkhvWQVcKhlkWR5NdjUk21lo
0bBJ3L7dBKIm/PS5Ljk57LQQLomCZte0kZfmkI0gltPaNC6u1a9HNQzV+KjnF/DA
QaKi8wnXHde3o4t8XoEcwYsxuObNhLoa/98ZI1WQ+uq8g8vx44pqfjrZGCBPPpl8
y7XkrdY1Rsa6EeNOFyEDYRJZG/Xj15EFRhL6SQgoYF1C5ecUXOlPXBjUuEgfLS5P
BVvgMEb/xBCj+KVs7sUlKS5fRYF8GUiKs60Xsm1MKT34+e3xI9tsIrl1tcwAVvVU
EkKxZ6d8tgUa/jG51QAijzf4TWStv9j4JiuZl2IEvQ5pZJDyAWNJ3yR3o6VCdLP6
7zqIOlw5JieVHZXlppjapufTwN2JnCAmMSMs23KHgFHrfLNgHzvIccxzz4VG/Ia0
KMnnziCfkdXsechRIkc/QLxQc2FlO8sVLyoBTGbygq3qVfs4vdnKTTtJheRtrFPd
rFARI+Bw3BOHTEYz3jaHR/ZqLtjO9yX9dc845lNfjPz8R+QcOZskHeBYKxedB2qN
0Wl9HMv/eOVEuceLHX60OODo+8ooRvSyLowt2Hv91zcm4SEaUSW7V2bgMyMuaK1C
VfEKMxKZVEq3xfACcfuca5yFejVzn30VKD5boEav1Ah7y7+7x9xSljfjfnV84rL7
fK/SuNQVV2KmJA4XS7wzK/o6GIU/bnx5X3C/nWpil+1Z9him7qAaj1b1ZQC4/pW1
Jt+6m6oRxYkfhd1M4Or2cqV1+ECNxIkoPp7tFsRX4id+W+pmccemEkpyemo+N2/R
H2PkVkbGJGhQ5hR3OA+VcBd3ZC+yjAdj+bmDiphAdAUukz0XNUoZn23UNfmMKYab
GW5fVb7sOiKnIznfpsdvMfajM36JhJJH10MEfzV+OiRTbo9/VvE0GV9GJiApLaWK
K74Q75lTF2YxcA1JdcaE62uQudcyJpsHUCGxrxChy1CBCA37sXH5GnrvsJ/Wq1Oh
3xMFU7JuU8GXQs6PAQ4UmTzXzfQcqzoRrG2hgsWuVWtvw2WQvwY90C7d8ePOyAMJ
ou81+oFuXYmqQ5GV2oPZDYTASYrpoZjSPwYWYvkbgS2cvDVAxrp8UbfOZAfdKz5d
h7Hpd4+tymCRqSfVSKOpS+dDV+rgZv8h4a06Q/rq1sYQ5TiMS17lmFWPO4wmJrk6
rZxDwqNUzPw8NCBrax20QLI/uNoavtBS09uK3Vo9y1K+g6IF/K06v7hxfpZ09ANR
/9ROj2T73cveh5jQukfPNgAKledchCfoba5a6m3LIqmf5YUXU7Fuw8vYs7XNyny5
ZJR0pKDDm7BdKH04kc+ZMZ2Jh2rFrhlG+ZNFBwpPHYGHR2otKttK6j8Kqg6xYlBb
qV2GiFwiKx6Rq5SYKJoafSfoD8bQjTDz37hxyeyDCzcoatju/C8iHXKS78PJ34pS
89Pu5D+N/zo0Vsi49kpI2Z2LFnYLsB9JpJmF6AuD5bH24NsPzkDQx5ul8j1Ald4a
iofUPWks1ip3U/vGGOkOIi+JZRb1NxFzC80BQJ1xPBBGspKaphEaBAs/zFSvD0wx
u0AIFVhP5vPwNjQ5LnjstABPJ9eYPPuvyZwT+U+oCDfnkgLMtWZoWc0E+Vzvp8fw
GoFOnoenYd8qiJvg0jUEBUwGwaX9WVJH3HxwhNg+lIcBGWglQX7wn7Um5wSkPMGh
xNLMYOdSDo/IxzaH0ZS3qfZYZN4PY+IAxfuST9Evtkr/FxSzPxhBBN+BR8xmQVHG
3OltzNUkl3oWlYgAKQy27Xx4ErexqbGrvSwlyoT25jKQ+oCCEn0jZ87UcD5ZuKnB
4JITWcnS+g/wwN+d8z3NLzPOpY7+aJMwLpwroDSyuSynDHsCqjez/KRLnu4ExFLk
CGZr4X+3a1gDFHU2fmsWZLCivXbtszPP5mWg6z5xrCB7C3m5puXV4/kOH7VVEb7J
fMwqE6cZMKE4Q4BwE7M60di396gGN+ldXtxeFQEL4TvIUuZzztOqkwVqfX/IcdY5
e98FJwEfoNN7whqm6PiHjM6yLg9GugkquUbB96kBK4gzcfKC3st4FCt7BYzCRjiw
7h3IJEJTcqkg+jxOcFAESgQc10oybi3Y5G8AZxH8TThd6kbgg7RZMhxVALsp7afi
gBCTDTTcgQOU/fM1fIWCbPKVuYBY/QeHxfTsRUU8PuXQRv/9DAe7xXbMiIgqffXc
N6mmm3jjViTVaWual0ao6lpKPCZJnTNd7a92kUBDX/ZXms9prc+QFtlT+d9u0cGS
YbDsd/9FT8EaPFXGozhzikN7RfSi/s6YqGUPudRvx+Q8fbqMdARStSXn7Lh+PHvI
yq9ZMe1kBW5CRoFKAoCDwUH2oruZW3W9HqqkxT7zFd4ihyRKoz9x+I5LwFjerdcW
KSwsT41KNp+wuc8zWgjeNz1NyUckbNE799ka+ntPkMDUwV3F1GIvfXfOzCz3Zbo6
TVSqWoObNUka7Q/VrCoh7Emns/S1cBgnFe+RoLOuFjNNXyjBuxPpowRw7rWTPsGh
RlyBDzXeKqLaxsVbHf5OiYSOPaMoGDFgvtgKaZoNMrifp4OyPG8nsMbNWvwor3OM
jghYDRaPsgU8SR3fbBJZico8h/STk2K2xmArD7UqUr2a3knUH5BYZpTDiI/1zs5V
5ynzhLxEsY4hJ9Xy4PJAQvdsJdAUqb2hRqd/sZZeHVVVIDsTurPuhlZAamyDY/20
mg4SaULGh1elkuo8VCiDJyqcipfakD25hy5MG95E3zXqOOIUJyV7i0f8y8S0ZcGV
WJ43PC32NzUyPiAIb7ns4GuLpGCx3TBCU2U/wn9prXi56qvlsBthBVKIeKv45G5o
oProlIT9KnD0DYyUDdFyUb5+Ub+zfDap5bl2i8WAOXddItyYihTrw/PldUy/Ix3N
mp2L0Sxn7AFPw3c5pJwWfKQ2JdtyFjw7uTWIHc6oUVk9tK2W6Be/FQ68E9b2pFok
fIiL5WgoeVK6izBnGxQ4HmUcA2I/aWUt/Vw+Wi5MnpQtom67qswuSVHWcVqpirtF
dVL4GpVmWtpB94auXhLM6sc7JDqtPvPBhbhHrYFM0Z/1Nl5c7CvDAnYPDcrV6z18
uRgSWDAazHx1QYYFLM4KhzeG4Cq8ux4fLgfmI+d9iTh2HuoCUrfgIcNyyNlq+bTU
I2PmWKREc7EeHxuc8F7GyflH4QAW5LPDUogbYZtsKbkV5Ek2nY671dh+o8ANnUzM
GpYZJXxq6Qdsniz5T0XNWSKgqIP0ILCf4NrukCGGTpz2a0Z1dbBcj0t+Z9RrMgda
KQm0CAZCcLP5SdXbCsBdJgBmn+qAhxLF+LZaNK7USw5S2fTbLBIpM6EF5PDwC4yY
IghOla1OFgsN9VzN8XhyXiUZMODwxusQ7rjcc/dojbt9eaPdbi50YaH7Wje9BqTx
9v/Pgi64NP5IB2fit2wI5JTJGAeEPc+VyGcs8QQ2t/cRbeFVhxXGGUL7DZrdKIic
t6UjdtQBmZsLakXQiYZZvLQfYensnTe3aWoBl5ZcE8qZ6T9xAoRs3UUmVbGlOLFI
DczTCEwa68wfSDJir1hEoRHTmWFHLzAZnq7wWc0DklIqAVF20Bj5xknypH0nmkbe
NQ/uxhd8yj3IHd2699YC+Is3ZxzbASPmg1lS8qR2FuyoVyBW3iCrKEjuGOBTrLrZ
qtzCnzK5vu+kyZ1/9txpJoO120VKh4xvFvYcMm9dorG/Z1lLCGMVSe48w16pkwzK
1p88W9wtyqn+5Pe9FYEO1g45M0t+JcXqL4MDg0FkfWxsQqt5oT1hglX4+mcENQKw
HSnDopKfblaMwGFOCUXYSKhyf2xPNKzIIGgHVW3HS0R0PjR/MM0jqPJnWA5lTPKK
JQMBzs/kX66IxB+ynNv1rnXIk+gkI3Qv9aCvkHIkSEpz/Tat58XwFqYII5Yhh2oU
IniSOjKs1w9+HSuA6G4GJvfJN3dAzk/M/x9m7u4b1X+SNEOYt/pnTa0C4ZnjiZ34
a1I7gbP9lB2PHIN2q5zAPaDOFPW43UkFmJtyITHQ0To8Leh+Cd4kFmPPN+nS+qpC
/X6uxquOgoZGZ+ar1Go1zXGmp/NAbZEi6mAmuEJZAbJAEqpG+agj4YOTWcNWu/yN
NurAX1HiH98rkBDNP4rT5rJW8nwRAindTQCjqyOSKJ2cjYsiAwNQaOaSmxudYw+7
BiJHluIp2I+L3yt9dWwRZ4YBB+6P8j1PaP2lQKZQ5TqXKOa1K22yI31mpZQur70w
PhFFbQlhfgEz2SSFhGDSxVAwRKo8+te0PhIVkkhShqMno0nrp6itysG9q0+KcQFp
GpB01sjZOfEMtwqE33CKhTkt5tkAfD+6Wm1KSdqU3bVaRYdzjiNvaL14zlP7xEEI
sN/vPJGBeEkxoRsUxFRI9cpKmNH4P5FYBFbhdxmGEUye6MjHPQlFCsW132ZPUc3Y
PL2M9l4Hf43a52R0plsY8NPiKdzBi6PyDmNO+4GmEHUCAH0zPuIs1FMnRAoEyq3+
Opoph1FztOQCqNiSeOiO9RD3E9SjLSYM5Ku4IlrDd4e73hpSTKJxsrcM0sdfjj4g
3puIekiiXGeZYGl795q1jOKQXiWvJOTxhCfPZJpRocg30x8voQ+8Nfnhoq1p92bt
fINKlyyf3jv3fTkuVkzIh6CBMnav7d0GJxI6xmlKxdqXySeZNhfPaT4POnvlfVOU
r6RpezzZwFzfhLNPdF6PlVqrIfnVB6j1uKURE8Kaf+clbf3+Z5noxIwFXO+TOetM
78sXCpmWcTR+56zgJd+0IvnlCjtiY7fgeHgHYtafn8iFk6twpheqXdcnKdeqVOjz
6VVpKwk3aOHGzgk3hqeIinqk+t/A9TKgFrKCowogqNOd5b15nCKiCpQRjyWpXShO
Q+aT81v+LMGL7qQks1wpXpacb/6+WDHFaC3IOW6pzG+cIb7JBwBp2M2g7RdhH0Gz
EikiOCvFkBoB6zd+0Ard2O9TEOUsq82dKzKeeOkNY6ZcBapEf8Dbwoh31zoPkyMy
2PMvgfCkyUDXsjhouk+4Z/rkdZw0sHl5jY9lydRsTvaA8CN9l3rEpqQS24+juuSH
GqZXFKWDw6cHU8ngeXSEEMoA6Y9iAoV6dUZNpyxSBHJADkYlJmHZ+HSPYYEy9iiL
OMBPPi2cLXOLcw+tws3ndr4qU9Rqext1Etmx1+C7o2jr8pT8a2tGG0S12J46Kshw
Ms554wKzdeo/jhke01X4Ry+cPZ/33SWsor4OepkrOEJ9Za+1bhm+IidnFeA21k+E
QLjmXhPL2ABJ8k8AIv08n+crzLC9d/9YHKc67Jb+Sa3xJh4TgLFs728yJjtUhI3h
aiCGWfUGT8oCBYu0zjX1eHPoVrnDv6RfqIo2FDHMKkZsbyTdXIQ1AhYr75XVLVyv
BNiIcbl55/5KkeWpfdsFlXz/Nso7awYcuFgkGQAf/05uE0o4ePdRPY0U0UpBtJFo
bFhuntvZ3PIkMNj4xm7BvmyoaFPPf+DWf2EHv7d/NwmwYx730oeX5by0uHEFn6KF
Aqh+8G9jjvLXLk0/QAOJanGW2Bjph2p+F+KlkfQlA8JDHeNcLYFCRl5pcktWiQa8
RK57WTxZrzb1LkpjFKj0OJHNrMD93tagoZCiQo6UZvt5VlOoGncicyfsStOCx4GB
S0/rtKmMT/phtMvFzTbuiHN6S7D1WKAkP3VKby8bru6h8/Y0DZifBMRgYstlDDjH
zuc2eLNSlBNuCllYrRhnMes1zkTG07jcya8tiFhITXacjeJTLVUTDyrujLibOe2w
huN6DrB0XhTG+B7t8K/KZhyalXaeoGSGQbwGIlFrZncaG3WoVkcYk8gkMMSVlT71
cz9YA7fhBzt1ezFsmdRbQ29ETuKJ+lf4dg0iE6t7LXqwY1a+QLSlRQ9DVdMf9bQi
f9mCshtKcC/mB+Z0/yq9rdF2dP5PRflgOxVrUeDmjEJhfUSvYLdp35gbXgnVKHbq
rDXoo+h9DxZDW0rF7ljYsBMBnSY+fMe7aiUWy9FLduWQy0pxM9RZpRbCFQMYW4mm
Hke3CuhlP6Fd7nGvPgtPZIglt6VcGTP/nms7s7uPdk57YTRevbBiK3xzmfs9jR1I
6qjUI27bXCBHP/RM5dwHMZ6gxXt30kPQW3o8odXjbblwZ6z6Pjz9SewbvyBGRqI8
Kf9R2tJaFBdh/Q1BXTBLV+aO7GkPgrTSgoPM2BKDDPzlhcNVbFIhP59+6sjopWms
wwHLD1WGBm/mbNM/kN5If5CGipuO6kUZ8rWkBoPSq0EVP3wTXEcc82Uo14mHd9KO
DxjARf7SkLs/PoMeALAYRVhBD8N2zLwOQPGPdEZnhdH+dtxtvuEBY1SeuzPYFClj
0yu25quZ2bB4fjqIjVDFU/TihqGMPSJFVuPqMyvT4n1JJjc7NDSWXCIQgN2Nlf/z
6yPLD9UXlf7hhx452Cf9OLebpSMHiK87Norz+coOrpdOdnr7+ShzTMoV1SCcyAud
u4He+NJs4LAWmybhWCusIen1KGURm2jjEg0BFBqFV/7qWGkU4h+AMaymUazwy/X1
H9xgd0FUvgYf89tU3kLe9v4Mq85A4hBygQB2hq6bRFNr0+762RkICpxUhjsIw2Iv
ajyQSn+nriu2ZEyFd3fbJ6+BFCJVOx4OKpdP3CvLnU5EyXF4RRsFAvcaQysp+de0
B8zXikVdIM7X72Pn2x2KeuSXANXsL1DI5vanzhnjyTh43ikUQpuY/H5ja1vu7rkG
B/vf3c2kvC1SCaq9MvyyHZWjVsaGnIW9Usm4pFwpszrtAxPE7FkNLlz+AkjWUHho
qunZXV0rtbOCxphu5x2iz8fWOelIdyKQGdA7VhnD+w9b/1oYnBrmMO/MlDflXNRi
zZaETcukMtqPcLy6qCNvbxQHiDEMlDOqpe/5UFXS+p9kab502jXH5m4JNP3a90Nn
TXcSWYz0CP1doQGsncg0OISrBdmp/A2L+PLxnk2lz5ujyJaEa9mVmKAbN5elwjDZ
wcoNfe6lYCaJcLx9HQc5vTcn5RutRzgo6g+7RB8ZQLCIQXhddsO7ivfCIRpy9WcX
+eNtAQshaqSJqxOClY5ddwbRwWfo6Tkz14mRSM8hhdp++vtBGCmGvGBASEKNs1Zz
MgdSeMlNFbivnZx68DAoupx1yfSiyEgzY0iCVxlfBiFUpZb0P9C+WCO1QIQI3G6Y
SzQkCblstKDQXPOhVKoxdatCcD0n57NkDx9DOinzdkvmQIABAwP11EarVTxdNCz/
y3lJGG7ufSu9AlbkNswwTYEIWRtM7QzutKFMGWrfDnK8a4uCeufJFp0MD0fi66mQ
Iisry32/hVbl9U9eGbzU2Ls5NAe4v+d4CZC4QBCl2thJg4fcoiqpziOkmCgCUvNF
2FFyATNfMtllH6hMTRDTqTtOzHuWe/SUa/bztDv5pMmVzQIyi/YfvQahc0Ad5ZZF
2ko4jQdwmYTsJCvv18trB+HO4E00eMMQl1pzVZpSfO+/qFhX1E7bSbsSgb48rfOG
hpctrqT+M0uh963IJaWEDBzP5E2ClcjH02U9REzZ25DATWo32WXsPcsTb7JDkzMe
q7Kv3eoaCE7Li21Q/PpmwIxalLRpWLbDR/zIayoIaMCDbvhHqF+UWsRCh2gJ9bGl
x2UQ3RaR8EUQaI7+FF48A8csqHphfqKZzEtuVi/n+QGSHH5RS18EEjSGrRlO8jKm
tNy4oASAqWnpvTHMYhT6WYEwlrFc+y53GFiAxVPt4c+epizXMdJixM9O/eUmtbi/
bS3LWqmMEAxMqpIQjZR7eXwDuaTqdHDA66ItFhvylmzJSPh50sB/Ey72UkaDoMn5
EIiufz4acf1689WQduuDP3mTEDUEok9DEYwmFLSDaOPpunihieDqwa4MYs7HBB3g
kjIgbZL4RKfAhah86OtZCFIXCyyfeMW+PYd4om7Giv+njmOovoetXi1D5EQHd+UW
v3r6Mk5cC8dDD3OWhs2/wejGv7oNgEmDm9rWZs1cmuy/1IDwRXL48o3JM81zOysb
gwvb5gSz8c2ogNu/6Kq5NKXBE+sLiDvrmUQfTvqFvAgeBA/D3/qrqZm+nJmIQ5H9
WehQlP5t/nGGoGWTgGJ07FwIRoYeMgHvqZ/sbMVMqaHnwzkcX/zzaNdZL+NLG2wP
hIAoV9HcOnbug8mOYTr9dMK6Nmk+yCRB8d3+XPghtfxhqDn3DHtxTp9+J/17YH1O
1evhaIDZONG/y/KJqFlI/zjLmqg7d88UlU85jRUg6Ujo3ykneYcSGhxpY5tX0v6K
u6P71mZeuSjCwXP/vnH4ZkS9ng37octpxEi2pZfnZBUmWIBUMGGgBjRB+g4C10x0
qxKUC0ypyC44McrvFNW6FfG37i26fVGwW3XoZODqEJN3YHYl53z5oWpZIemf/5xE
IwcMnfVSOarIE7l/mTkbFycy+BMxoBqcZD9ZJx8dd6qBWr9H9jekkt5SH6j0NfoU
cUHOXVehtQGERGw1mXALZ38EID1MSEqhC6PMVbW2ji+RGL1306sqLyVzWLGD81ku
WvsC5LECE//PhfzIyxoxoutWyMetcui06qZMeitaD5DvniOz4JV5XxTHugpJoPel
0VJ3nvcrYeHX6cJBvtCuq3Y9gXHIlC5qRS4PwubTvDZGdjxNdwvN2XBL/9hrM5gA
rxqRrgQ9DTeLHWuZ2UYU9dKzx5T/LRLShNjE7y58sBWCzYvW7eWVkj/zb50J/5eR
+LLRFvAFwOuJdaCmjIXbFH2o0hWLkPmOkdgVPNldEJ8jcQMLkbGqkP86sb5R26xH
KlNlw9vLJ/PPHLx0qCRkdVulFwn49vLqFEEEB/8sz8f63ASj+Z/aGv067fkaPCVD
5IEnlLgsRIPOVCO2HlC++x6AZnWrVU6SW4/6iwtU72lPMJONTfAw5NpfLLb0zVyi
1Ic+GAZs4vCu9mBXf2SOB6Aw3oVcXw5HwQJCZhNLgWA6DRf6JWqvppx9CyydI3KT
SrkiE5d8fzjWPE9+56AhTx0XcrSBTUYau+hw9/zE6mhxyYbkqZBmtMkqB+I8CmBD
nAlP8q4q/K7oy97f/ngtdDM1Nt6Ax7g/goGGeX7I81W5h4TalNVwn3iew/qb1PAl
V5jfQ4pFZSYaSWlgeBjC1xm5kBsb763sbdCKFYlE8ey1lH5gVQ0raflKko/ioVtF
MoIJDxAhWbPLk2Sy2YHZeWA4TxwWggdiloSQ17ZO6n4Ypq3oVY9gJ8fhnYSEGm+r
8ixiZPvG6IE8dZ9ZlDsVXjtJ5msYcAmcKs7QknU07SU1U46D/YTBV4r8tfMkgQQI
fNxcVORo7NdqS8TI78Z9sv65oyv3UfjBw+/ICGCcWn7llh9agh+pLCMpSx27/3ZY
/osUCqD4Wthz2ztADf344AeeCVukwoUGii971weRBPpwIAruer12sSPhf+7fY+3n
+kba+Ws4fc40Gd7vAm4FNUI1U0XdRfioIIYmxoG8V4mRwxAetLyo7CHSEwu2CPJg
yIpVGFm0njcOGxT3KR8RB68NG0AqGMgWKzv9+eU48VMiXaKxRkcGC3RoIdeJikWN
EgjGhyPqe8NLsgD0Dfc1BT3iY5312gYcDUvzxPFiYcO+iLU2D7PnIHwpe2SpKuiJ
BgjON7UprIHva5uFRSCEkR1eRR76Bad3T4HhTtqsmcd64ILwDcMZkMxQuVed/FBs
JrdRYfw74whoffTWvuOW40L52IrfD5BoEaw1KpYT+GnlhbLul2VcZAnxR7vrkY7w
hDmEtwUwx7EtZcKsyhHwrOql7UAj58jObluXUk+lYHN5bcI3ZwD3R96j6YcXf3Ws
gpFfxmdVrJaC2aiu7TNTLK3+2ZxxsAgEwG3Tbes/sj2i9cXWyEUxn/D+aV66Lofe
8nAZ31mmPxlppt7FCSxvHsI2rdTxjdstnW5JUOSbF+5AwBflGjG014vw9HopLTNc
9zBZtcr27d+EnOJzZXhvO/rYfCR27sre3zWw0ulNxyR3pyo5k0VbzVPnM7mCcFIB
0LE1R3BpOPQznteibkmvo6Jt2oI8jUbHHMZHiwoJGo88v6IObFkEsbI7T1YgWEBg
3yEAmb5ukaU3ZP1hM7seJHK9OJDQcuCiGBLI1lvIs6c1YnjikzyWcUmjSSPNxUxg
ubRc52uHGpD8u4bMa9wiK8DwMjBXdk+gQMPs29mgCEzlpdxjz8zMg791IR23S677
TWmj01yZvBGLAfB0ZCDGlZyrSsd7kX+UmmDodaL4PVaUnzClEqh6zCWyNh37VYSW
oQPQf0bOkA4oxz+PdbbPlVyAO5HH09q8trLNTBgLrJLtJsKwuGt4J8RwgMr0t0gS
q6N1mSDDnrOZm7gTq/XhmwV8y7SsL7DWncXs087zd8tiE2lL3AacaS6D26qSk0Lj
nQl45oVuJmYY8KBrNGaio+c8ys2Npx92cvqxAfoyZpp9zKGtN5ehOvKiA4LA6/iU
YaDj0o2RskYLi0bXHO/OH/0+alrAbLz+yb2t7aX5i9oGujrYaDMVL/CLpXYKn61D
ohCIr7rvhYHiqGT0KUkvCgOBs64qN3Bqqw0ZdNmv1uFcdXqw1OpvXis1mljamhnX
HSlC4s0cflR/qgaKQexwpsu24N7iZFsgQhw2cLmp6uuIF+elmWlrmNTSXTOOG0eU
tLZbEtJvhwBeqOSAX1Q4g7kL2l6K4KHKHep8I9/LxapKq5QC77SfCqywqrhkEwHm
X0RDpFlHovfylTRsTrZyanla8c7Do7TSPJmV3d0JDztcPG7QhytIFrLjTMyLq1kE
khy9KnVfaANC1d/dUqRSmJp5KjecXBZlqJHG5wb5sGW83CAG+25GZ+y2o51S3IHT
giBtCRf97rJ9JSUCNVTgsZIdlguBYN3mG065u2ZCPt3mUMJkJbV/c6V619jGmrko
ke6GtdCIml+67mSpS79ymORusWUlOqbc8paZIrej2if3qcN2GY0a4nf/sVArT1Ir
wUAUL+0aRO4UdA8U0X+MbB/5Gb1GwJRCPYO4P5VoHfI/CZbdZp4LuNspLopjExQ2
6AJdE+/ZTSF251/KWuofFvNUx66d73ZRYJe0IcBf8nlyWLuhqptH3OfEXewhq4ji
+hnSTnfQ6F+HLWwzKx45XxkkjgfMuV7zKmVZAVMeRDCyAcRkttalj2grl2oUGSzL
FAjp5yB7I8n3S97yvSwtmgTGYS4BwEuwGVXXQqOTZ/jyQo4x81UE6CE9STJr2xEz
tkIugsuidvEXsnBf2c2R9PGw4r0+kJ9yHcdyHFflW71GJPvRN64pUM2L9Of6Wx2K
rvlEm06gwf6RuwV9e5b1VYxnakOS0Z4geQoF8FreJUOYzqETA5C7S6QQkYpyloID
4kt47batnQ+Izyly43EC5ad/6KImshB5awCo4n5VKX5Fs9J1er0R6gqgyc6z57qH
Ekhui0PU+vODDn/mcYXxDJ3jxTFhJBaNhFqm+1DFIZgp+nnJgCvsakdcd6deYPWm
OXaSBMQun6PAOksSu56bJnwowFFP3P2FAsaXAnLftJj6Z+hjp/PUZHFauVWSpgOr
fT39fVjW+CHl+S5W4+Q1W/oOkNsA2NIuPhz8UbpwWCuH9mRwq08uNjwk3NRNMSKu
mLp7gOU02qBlGlfdKbbv4Klf8/P7Jrmh28Ksxyp8gjHr728CQRIJW7gi4WyohErk
2Ou/8S4lyhCrEe1ytEvMPQk4sa1PS780GJ8gWcbMyCevMYzuQvDRms4+y2Q3zroy
ep04Gb73/SjxGyDaf8U7DVlpBuRq6TJQS+NR1hFxhP6OU7S0gkYJhNg+pHNtRtI5
axEXoYab12j4uDJUdek3ZZlRvIpjFM+oIZoi9krUACvL+dL3WhaXcz9NXB9F4NZL
7az+ZvXvxNVhaah6qf9ir2S94SK5WJ1hUVkbPJPp6WX0CSfXQj8yhRoKnFL8GAsW
MTY+mlGdYYuEzMEANS48Or6DrFWGKFN8/hw89JDD9kK4R2J9a8j7stFKkzqgoOCB
2w+ad9MO7J6h+I0WIyQ60wpH1p9vYW39MuCM6JjZbZKA6mpkPIOcCDujyJwCaxMM
tRuYi7XZPwzgzzDy5yM/Jca0eMjwbvTgODRrae7AzXt2yRWEtrKPtcbAQA32Dmso
4BWBPAX4LTnmNlh9JisbFBde4OmSZmHHoxAAj96B3oh69twngJKhQ32VH/ujBoEr
Qv3Jb1J6LyEacZN7Z3DSfrcVtMmIm6Sj09NjKAy2Cvtb4X23ZhxC1ztRfdQ3e0y5
x3iNnaCFAaYXinz3K28Patlg2H/citk/K3mEF7nY096CQ/yZPYDlZnMHgykt8opN
hD0/2L1Hmbpgs6IEqMnOQP6lxOYJIfiudi1fH5ZZdJl0RXl0okVewJsmlO0999kA
4fV13xpORby0EDSDuBgjgmQIX36zotp27qgpQCI7ckIJTD6wJhdeAlYgfP6s7+cx
o8bJ41nZrBXLijsf4UqYAC/I/kjd06VpxUw06uU4ycLCBScXzHSffQrk33ERKc8u
QQ+WsQSVR+Q72nZ8FlHaKrOp2UGuzgGgnrcmxwpmoItV8HJzX9TtpjivfcvyJ7dV
kvIPwOSYJiIva89x/fwZc9mEGCquzTsaPo+yIl7Xzsa9THxDpDwiBeyVt4KhNleH
/mi8FN1zCkgQTvm11zqNR7IXkx6cOpoZhckv6yLqbPCTp3y7luyruCZkcF8jL+/c
MRIMLkoAjWRvOH+QVBoIyWrLpwt4aipVeJoiyT/dNuumQz0shu1qFOu2oMlWZyQA
MiZEwc/gUrefZD8XjqPcanVZh69eyeycubDaDJuU5Zd8YGC317YyuchsbTAcsrRv
gHYU1Ow27PblLdG3Wuf3ENIcSwykoDTvdilSV+rE+9GzVMEaIfyfyMjZIU9ruyhC
thTLYaiijGS5CR9T8pjFmETrw3Cv/tIfdNjcp9eY0ax5oiTq9V9BrJZQaM5dhmyD
952frQt0NRMsPazVCSmVvM8XX+UOqtkVLWU108ggjeqpoJdGhocJqoeS66KJms3C
LveZxrzC6rbSLEYHqvIRJjgioBKzM7jZ9xErGVTGgguATykhb12zne8ubqBpoSTE
Y3UNNC9FDR4fCusUWBP+9nzKl0n7wK2tAvvKQ64mBhURZiQ6krN62L5whS9zNqC5
R9jP51463wDKVYVGvxH8eJRnzE0Ij8iJQj8PmU7SkPgzEWZJ7SpMZUNj8nshBAbU
plmt5b7sMC7SHFrs6Y2fs9GH3AnMsSLRFbcee/aKu6POi9mKfI/J4v3HPxUEI0rt
o/mRSIHt32y2T1nsOLVUWIoS9uHZF64ro7z+3EMQP24rNWEQKF78oV47xcQ50QdI
CUBFa68itYNgUyU2g9QWFbUmxUrm8R1VhmRS+5k3HuK6U0dd81boUne5eEN/kqaf
FmR8If89SMGska/uObRa9IlMPFpy/53CSwe2YMxAv/V4qNjIXTaToyJpvEoECIaI
jqHDTCGYNwHuxDLWZleE8ar8xX/7SDOwaAYWOUbmVaoLTvriziNmoO8D4pv4AOhY
k//lkaJXGmkCoBk9FYwVPcOIRV7uc9MokbaYGz/QC0WPBcu5bxsWZx/2UAn4AHrX
g7kiTHdPXvtzIaHedMCs4K+3OrVFeQ9bp/PemmaP0hzYkzm4dwXS9VkLSpqcgt8+
deUxU734S1uukfhYOwVK/UVkub1XWTwjUd8MVd6fGpnvs7GzyN4lyJYBfNatHFRH
HIMd6J+xn93DpWkz7FwgifR4CBjFsldNa7EWgWTrJO2FThdIVowoGohQA2Ral6NL
PNhpSSzTP2LQADQKJoeQe0jxuGezSbpHFDNvEoo7gutWFFDPZIOF7P5UF17BT1Zs
hnx8bZbL/nJOS0ud6Bifw3BIQ31QryHtMZxv0XB+7Oy4dU1oxtPNvyDxuJK14EQF
p4h74YQjSFJEPamjKarOOZkaylvd1gWrToGnAvnAyMgr2QFVBSkbZz8SYYpqGJuP
gODSkRqP71YIr/M/CKbU3qHTkkGHuVtRtcnpFraTEgfZp7Nf8gNHAPzzUvJxnXXk
M6qYm3xDeJEPqTd974GsC7NPeeWUka1B2w5MTY4NILD96r9P6L6YxprGdCfEkXGs
NyTRCnyFLXIQTyP4cafIDZVXzlxpWC44xmnxw/74/QqlU4LP+s8L0r9GBI9dBwim
QtX8UE9oxG4VuP5bkSxJCKH7qYoK4On54sSf018jNjYgR+vOM3FlvXcaYCNVhQbR
Q9JA6RWd0V4J3yaaFwynANadomFzBqOpScuXA+4VX0CBEI0Uvsdf5dWXflJmiGwc
pfHw2PEzI6QibgTgFUefB/jZl6IuY7PhVFYvZUR4maxOZBVofzy/R+ojMiJhm+31
fxlQSvnP9PYe8KZ689MRrUN+mHeqGhp9efNxpHXu4ysZoLlmc3ZahSeqknYo2I2t
ZxKjNDw8epCNksPwl3egan8eMF4g6RNoYd2Zxi5kCx6OzZNLSHS/C4zGRUCwyI83
Zl6SD47d4SgNIsxZ/KC+QbgK1NZk73CDQy1lgqdOtOH0fc7wyHOnXUiSDHkKZgyr
0wKy3HNVdHzElJuihJH1Ycyx1wI8J31n5pHi7eMl3fLOZBq1sIH2weooq44H3p7d
F3IO6dBGSlEJN+YGuWyO/o2fFunQPTZVpNv4+Y/I0uIM8BKa8la5mD02t/6hNHKU
W2whhsm72QNG8fcVoWH8wBPrZUymab9MWvzgHwLgYOr6bUZjZLJyeLDDOOXJb87P
Oo5BC6tDZrc/vSdBPpQBRknOKAS3688n5e0ZpOBTRvCFX4/3mVsd3TNKXZb+HBZ6
HbFIt0b1dPOsU6S1kLuYz3mzWIbU0Ry8skySPSX+ySTIDM2b9p/TqJ0JWS7X44/o
lq5V+vSCUhj6DDW9yCayYlrpHKjLB7K4fkep94CpBySKIkIMCz3sQoTXLnSzxsJt
QlrCBtIedpUsbIthTWUzx9bWC6KCEQ1omRBxEXUh77beKZqsDvsbpqc7EK+pHlKF
crLMEAv4XHO50ySlH2IS3lKqp8Rxx7c6UoixLUexgLKnMg2FjuwSt+J3/4arAO8Q
IXmhCu2GJk/Wb1HeAmKSp5InMMMaIU9lqGkxNc/b2g7O8vja6CcapEow5LWqj4ad
DuDPdyEVDnadRE5g+0Zl4wjC2vGbzeX3x+mW3oxFZEyp4sX7bjD9l4+wfFNqxPTp
1plj/tVSVQIBa5qpP1Bc8CC0hKLRzT4bDoLOVMagLwzirWuMwZ496qSVqqx7SN6x
bPZNnLAbS5DjnbPPusSUda4/LbG8iqcCJH81dkdvoZT7iUr7e4exdP8pl0QMCgHs
1sKFBOvgU+IjEefZljiHz7eS0PW0IspuhuFyKGEQCsGwSAAxuBx6G/aRbNpVSC/s
nLiExoWpGJ73b7E25I+RQdo9HPx0etj1ddWI3r99vj8ejlClyaN37+02W6WV9kGY
3jFWJ3awiSwnYTNz1ngqgVEXxaLrLu4SnvOC0542W5lNdL95SVdDi2hWneS3KcRf
bqnFEwHGPZN0ODN3P8wJBqmM94F0KHyzYkOOrM3CZkui2tzvHZ6MAA5BQeUwvxwr
JeELeWgytDkgVbTWFgiSvUAARaMI1I4M6/VKhMPsgH5NaJigH4GvOBL5caSNvEjs
BG/gNrI+Dvn2WyLuLlJHF3j3uXSO2pfli3BbLiVN6SvOquuIbjkUOXGdrf1OFfBG
iQN/hH8ZELvXW2qBSInLn8dHbVP2Qro9eIhkle0cylmbthUwO+Nuas3AD/W3pyXy
jIGVZyhyUAwgRJxH7GuSPoZL/FShf5TPydM26t1DIeNsvWeemn+/H+BmmlPiiZyn
Fptl53tudiDL52ua3oX13RdUTJexPzx7t7Kp623DwwkPqZUqe6eSOmpcnE/YYTjd
0Xqh0oFiGI8tTr9BR2rqUBqvpyz2ZJaPZieSD5YFB5u9+0CDFVnxjdLuH0AQ1Pup
Vof6hMVpP14y+VzwrWm7a31ImuA94+IL9qrSLllSXoZ8r8Y169xhe8L8HUD9W2Jv
cyft0zs1kA9J0kbJkzAO7LzBS5SAJwMv8RnTCtVAoWSVoAUNCHVfjvbLs0lEfXXi
Owe6+qwhZ22rkuuELvO/gfUnyE0Q0ZvymamISOzG58s0zGXdylJdDD5CjfX/Qhjm
pC4D6MpkOocTuH7I44MUgVioQgw0LRGMywVIM17eRRmp9NaBA9v2cn5IP3n08JsQ
3Iomf6yJLtxDpjFXvPfJPzhDiGuC+v+hjpP/6v1XXuQQdagFO0F55+GkLBstvwc5
5FguNihx/bqhAE+h+K2buYf1l2da6StpwiYsDsvqosAPi7asDaYHeLfzfXZozYSx
PyFVHRc9NDiUxmNcjrTTsnmuAUfC8mUUj21RP/DlufeikhE3TIcPudNG8TzUT8nw
mzUIngLmSESQrPb9Rd+50k3i18xM3l5A/gyB40Af3xBxZ7MJNZxOxfwe4bT1Io3t
22bS8mG8qXvFCdjT82SdPhnWZ1GhFgtLEjseapEqr69xv2jcfQD2qpiearEdk/F4
+tsOcnKiSgrljnjYWxCA7O0cltcki907zTnmAykkUSbAQRTMaGrYUo1nLJU+k87S
gHOf405cSLXNcrbdj8iwwDhQyu+5trbMXdHVdcuNi0sWnO8YNwe+hpn2WrFKPx1p
10ewllgihKhl3SJXOUyuxZkKJy9yjRXZRR6/PQgGId4LRgzAMhp/Wqm57V+HSCUC
/4NBSKc7zW2oMv7wEkoQcsiR63MSd+FxJx4NO69IvHa708nek6IKOtcdTq2O/Itn
WnmUeLuuDR0j4LLXe9fkQ+Xn1pCXe9M1z/TKPUfSGeCG+wUoOsQO6n8YFOigTjym
7JiUvKweby6Vu87FywGZyVSWSvlgcc+ePKUR+2JZamcfwd+wHoaD4KFD5NgyYk9k
Rm5c9QLllGQOiMFTBrn5oJRHeiBBXRbkf62vFAuQgCE0cvk2X2OkQhUOvEciq16m
XDUMvobeRtEmemaZSbPNiFgdqXCkfm6wERWXxIR5uKOjoYjJL8gCZ6qiiYfFZzdP
bXjY0BsPWXZOvvODgSSIS1zKozWgdwoxV9m5AS9m7YjNBCQkV3Rb0uxerfD215vN
rUBhEkeWcucqElw1uGvRA2jQ6PYjjiZgWk9Ug3aAFme1rAjYaftxTV3Ts+qWti2W
XgCPik14pqyUpJMZSzeDnbvQppc48GJrh/0d/VrTpyniIC82JcHDdCz2ZBpA8llQ
6QU02mrJYIB1m6Hbn8AV4EfSX8Gzf274Z/aLOo1GN5c4a1K2a2EYIl3A5FmycWs2
nXKlf+V7HJpAIW68kZyfeSGqFATHbqy1jyd4Ykr2cMwVn9bqFvVlpWQg05j3idDJ
je3FUEiW8ZfLmitUIZzP6ybnxPCDnn8zueDVyKxZ4XFucl1VnJ4ker/47BwEDyLz
tJUsDrG2fF/RELNJUePQQZbqt43kQPkzu6BhP7+ixJ/mo9Ke9h517AHxPM4OFp4o
gIne6s49JIJmbvTS3WLOQoRxTHvUQAjqIrt6KrWpqUp2bMLGrt3T+g2/ujZJ4uLp
HEGi8dy0QTt+hGHIZuMHP/YzWOgRkRUWevI7/c8qfVOGj85VPebtC8mxhLsbue3l
/YKLTwFUWLB4Vpd1tKkLStjociX0R+xVCpEx/Yfw8OG10ruROJCtYUyKVpaw0q0c
hxTtX57bpMDvLm9LzvKB+JRNITp9Mt9mYTB49Z6MeGiouqn6Yqd0QGM9p+r8r1sc
fkIGeEovdApFhm1rczmKT3lXcxoBOLz/Hf2JnxuzVfplSKlQ+NbEBP+wRC0n3cXN
hrVi0fOeEjkWpt5BDUk8hFDUdOW8jGQwzNsthpGffBXgf18Yvog+g1ChQpQ0ClCp
f/XWvvzxJOuDrvu2Q89nq2hQ2dzLMpnj/VAqItdiKg+0yEkHtle5ZfxR0vYryQ9A
+DEH+rq5EKups5jsgNj1CiFA2dO7kIsYMaw4HYiuByxlMKpOChW5jdgkcrGZmIFu
d+NieMywvgYzNgNUftIZm7wKY19pUR1hSS6dIRhyNKX8bZx0oWYjfaviGQzzuQaP
7vpxxWcWv5bI8gZtai+AFUd0LtwRpc07bwKdaiNPeIc5QO4ErHqDAd+OYY3t/qmM
3UzAb+nvGCwfiLycUMVg33KoZaDqIOO4lpdG2s+k9LOL9MKCWk2N62eL8frpE6ex
mh0zX54zzT2myOAUkViti7kvlf68fYwN9W9a1qwFXOKI3WCXdgxt5RbMg2pX6EKI
wz1lYqf1ffO4Js1bIFHGQfIwwIWiWceUEzE2XGIyV1QnXHdTBjVT+jH6DXmm4H75
kk4ozMgFSLVyQR1hunLbnLmwBpHGnhiqWTU8w/VZQ+l28eQvtzUyoOzV6y532K2I
M+hPjt7OzKid4NOeQ60No++6FkKiYE0w5S49cWL52ljhR5bTmJLYchTjWcxot6kK
owQirM6m9wtDjQq3dsq3cVA4MfflicF9z2CDn2xDS2TkmX5/I2+0iRsuf/v3JWFw
uXB/Oxinhz45EQMk7qX0aowBjjIQiktAtFHldI1UDUIlzN5Ak0fEV8/XQxCU9pxO
OyI53P+m485zxXfiYnzZdmEyMhSeciu2tUmTCQZcxnwQ7ox8Ge2eIBMAqIt8gFSz
t9A6G8EGJ8LrMkN8YiKzQ5feMuhIcpVSqHbcKc78K0Vavo1KhcCkLy9E7nA9p3EQ
slX4E9EM5Dvnj8uIl63C2JNas1HP++52jU5wrijiRJFqHh25ZVdw2c61T0tPBUhh
qq6C8cNYs3OOtFExff8zGsyayiLw6x2EcATFNb0xZ4hgiPzVL2kUrwEwCUIiufsQ
VCFCRzMC6oh3S/SNHgYZSTK8dkyneOC9TG7z460nbXCG/ru8/KMfFjKsgmuL+j75
aKYdLk/VaMfIM1C3/WPUg1CavfpfMHDc9w2eVi0OEZHmPtxArsd+f6VvuS603B8k
Oj+Jn0Ytp7D8gnpdZkkVDDwnNXEsCj/aKOks7sQLkEDLYKgXUHD6ohRBeuNkWGVJ
rWYbxi3DObzKnSud2+UtqjwA7A6/ETUN0gZoxBg8zToITFx+s2qj9pCPH2wTwd7Z
wnzBy8OojgrQTy1S16L+/bOpELvaP5jJUAAXsz7N/1AznrPN39YphcaavPHcXIdF
hPHugSMd769Atm8PsGbFgdvRlCHNQLMpe2nC50zYVyEd4C7tu6lJmeV4P9PClGtd
t7Fw9C4UCeaRSvtOblTpvsfAWE3MdCbEPUze1GasQ2HDY+r8r05D8GuQndAULcIu
uaOnPgs0zmSAuIdaBFrirOMNA1tfR8pCR1edK8tzWboJ+J0tdo1tGTfn/CEw2gdh
xMFETCa3BKu8k7a3n26Npm3M3rHYS5qJHBca0sEOBcICqrIOzg0QUMSIs+Z95EnV
/Smj/9kT7yYAb+Kq0aHj9kAD/rROUvtMruijTxCvCYO+HgDotqTGOAZZCJd6E4Fp
Wcb4Mvj17A9q8fM4C6v1TwWsHxhpDz9OaR0XhakYyg4PBT7xK/aBvVDESpI/hqy+
MWoMp2aarDv2tOb13YewuOU57840ATOy3WwtmAoSWGf1A8sSLT30Wfb3WGTZKwKQ
NfkkMvHLFd1gtQRfbrMFLkb+eatx9v+7gvIGyTlYIN/vZiFPfFsjDy9J/IPfJvIR
aiaPKXiais4DmkemH+G2bKvP9zGyQxnFQZCDDpI7uvsiPLMYArPIgXS4VTC3mUxI
kPYfKPpeLAPEM0FdPGyInwlyWxH5gTdxsIj80d5E7xruriPBvlAdZT6CSsFNzIeV
H0Gi5RNMK3+w30U+sB33zODpw5QQEDE5jL9LFx+tGCV/wKBYtSePQyvMKlwmnUQF
eRo5BCw0YKful4oSveK7Ee4eXcpP2/zxBmSyxAqFYaaf0l+36ingyIzgZpCYt+JH
YNRylDgW82E4T71+k1eK9gJqi10J+dEjfESIaNe4nDVxgaJv/sZFahzcsaPM6DBJ
581eJa3socZIU+FCqcMJf72/aXoArGQJ1fQVJd+AH0l6LR0+kLlIRV4Chkh74EaA
9iQ3zxHzqNukrnP9WcUPw7bZKPc2mBbLRHhad/JQ29N9RAEAtTttPozYRw0HZVYI
nNjqQAhmXA+bSi3b08ytouajjdnbSKirIHVUM3aeeHDLhX0lg7DqoZZBJGhIVfa+
6yy1dz9oSQ+J7fjIPqW5wY1ckwLOs/MNbQf65hqVCnOCGWQTKrBSshK4ri5dpNlz
Pq/yi+BquNteeNrVKjS77VrjNxMt7HbPIPMc2xpKYOR57sJaiJNDH6PrqRgb/oGV
5QUq78oS4NeWEFGkg0+b4PcEhIpe2RCpr+iFb5PK5CfBgZuf2NW3omSic18gHgPV
8W5uzfph6vly/54XFY/K77jBLyhCIT7h5dTsaK2UrCaZT6hCxMyxMmrpauTENp9n
xN47P+ePxrSdm7MMdLOUmxQyIFiGFAtL+BNLKK2kbxqIaQwczvnYlKCR9cR0+G5F
La082wjdxMB7q+/qLm8Ij8SVwiUQXdn5Db6+4O8kRvvYRTQ73w4PeQ21SRkDagC3
U6r8AeUy5YVKkDPYdY7Sua3VPh9jsVoyIh0+ygxKcOV0jUddBZsGWLdi+7sb3b8Z
UGSAZyp3g79EFBMgVBKoAXbyPphliHFgn2MTBb1DpI0JlFhnlHhMvpxmfAkZu7NJ
OaRSTCVq444IW5KZ+tomasCDOXLQxlc/hoyKobtEzmS4r8pjvTaYhW/R7WFVATxZ
sz9Ok6W5VSCXlWtUqOUbTM9zWXBKvj2N44W73AxQFVgWDAMJ6k4izgHtFwbBFGmn
WaZYeisPEwjK4oB7xeQvyOw5ovJ18EQk+E2/mPXrqBNZiJTE11TE/iqaa13Tr8Bm
/iM9VEVdKUksLIxo44K9Z4XHY8vlkgEX1wGR3gefs0KIdefCQAfSB/+gDODBucP1
GNGrHaY1k8UXA0MzmVlf3cTauYesGYDbx0xoIr6h1eeLQmk4ZlO2/oNKOBe7mLLn
y3+hDY2rJYzvkfCDK7LSOzx9gr/2Bj1Us9FfFfRqSUYqSaLOxYkVoqoyJ5TFpsER
PY2k/t3yJUtB1w5dQisEIP6tpBuKeoNUoArLakkPjTomqdTQfToSeZIiMdJjup9B
E6x0s3CPJDkru0G8vZZOR0usm+yc0CnSff8yr7SCQlr+UTTJMRwnysKjqKNbyIMH
da6EHCYFzMlJBeSv1gs9TZu3XffU1f6QSSG1yoBas5iEA3BK44M3beIzkF9AtcGL
VikkQ9a8HpfESNdPhiB7SeyJEMtV76NV53CpNVglfUu5Y04AS/vlrZB8tfoKkfNo
wR5kOC1EnruHeZUudbuo367V01tRuBXdusoet9EDDcMQlee40SsdgrLJ95lJQCjj
H/ZJspUx0htXoYjot27e0wYeZUjr+8PE6rOf4kwtWctWaChaDb7uNjdqot98ynsD
HNuQwEye1W9OISMF939qlGNr3Pa4tbyAHsZVwCyYPXXSbXzfBvb+s1JaN6ouAwMC
w6qbdI+GzigDAIIo963ZnOruozmIlDS1ukk/IszyEnL1Ynd13/FFvP8UZFyKbucv
+513MQmthK6vSKYcX8R4bQvsYc/xrQqEItjQNpKNInCaZH2C+rKReudeuTFOxH4O
VuR52Fz2l5cXCf60fWgXgwiyiYkwn44z8td0JTn2KW2sA/Ro4X4lwyzMF2l8CQa1
cQ40iem9gFbn2EKsbms8y2wj+rj2RiFiZPRoDk6jFwEPfeHVpDWEd7IwWnH05eLa
Lj7mW5WpRSFv9w7oneIuSy6c0cTXoCkcWd53GmVTQJCB88W6KTfQzlFnV2CwiYyU
9v5HcFva0kN+p7nV99GZZ5fVf4TTOPxh6PV4gzx4VpelMxpjRH5pmDttatEJj72h
3n0pMJtommpL1HZzjBQVUkCO5Ob2uLXPa6j+TobvTBomGEPRIqGUlNYht4avNS/a
Wze30Rco4qhWhGreRBLF/WFHmyOQ+R7OT/YXzaIgE7nesgoE8CqQpohUaNL6avJe
/HwuViuskLBcpfKMBL9GJ6kuYGEN74O9Ie0Mnd13qXIySyPc1ZEkNEZWEWl6UsVy
R+lzsMvxApv7Iet0bAJGkbpW2uQiq5GVwu3qdQD7Yw4U4hhHgDsM4k+sniI2HDDq
ArJArwJRut99vVZfZ+KtaAJupO+VdbkkVvl31eLFVs4+hF6nYFAqwQ8vXbacV6o/
047LZOeAr1E7AbIdPRc1jskX9V8sG2y/jOwm+ir5BE5jfWPyTbrLsODcw5/atwyG
DlW69oCXtNpmcsQVf9R2pGsVhoA19KuoO9YhDO5C3wYO0RzMDWkRXTy0FXreyrbd
pDfd8Dcq+EM2MBNasvZar5Ck7vYewnOabbMsuGkV8oHxxifs7VgO8fRJNzjyoD6/
YMJ3Hthq7/0dHHJprwPOTidxHd7WINyG80HSjlIF0vyMQsWYx/+LObb74ofy+R04
Pq0ALdfkRt9CC3/dlmkNw7t0zJQVLBvH1G6a04EsmTgk2A8Df1157noZ6Iz/zpsw
rf3jO0GzRqu962GSN6D+GnoNUUNz7Zbcsc042bYqquwbtruomlvjhi9b4rzh0e4K
ojnduKhgE8qDISVK+H9edVlCQmOcHzqJcbdQXcM+9bw6nR9GJjl+X04dcmTqEAD7
FokCjlvpEdWluRMNkDmjf/2z3vBZWj8h05a0LzYiemf+FctGCziHCSOCrIlIVQOK
0EVj/roU3CrKmRCXj09ETfPlch0Clbxv+oiyM8Xj1DPaCKZ534Lrde3IFmMsxmUj
ThlI7SXLvYqsgkEFgLVnVpATtd7uDSlJrnfElhwTUY+l0aPW0+NI3x1JzMuiGnwr
8JckyzhGfmfckQb19AXrR4IDKTS0GLtLRK1WBkcl/1iEP6ImVRKUBVBc6udETrTY
EeRr1iYLr7mtoNcWRyJMh2y3LZGhqq0t8Fts7QWLbv5YGvLsV4qDrmVJT71OoVNR
1lEJMaS4NLxnmGaG8zGhJotoraJZnwdih7uM18eU4Htlx3U2KR0R+Ee/BMy/BisN
S/a893xRPS+bso/gdMDlYw0p0XdS/UO8amC38mvELck3hPCsm/0WNIVQBQSy/COe
jjEjTMVfMIS/oIiEPG9dBNWJbtugA53K5Z25YaCQUp/unooUymA9+KSJbcrHhNvp
YaB0ZB0Gjq8zYJG4raOtuL2wCxcvFaJBuK7mc4y9TNiXcViVQNKdzRqi83ehQ7TM
NY7pC48Hu0LGvuSoOqUhbBCslKRHZQBL4qohtKw+JzpdV9JvLHGQWKYx2uiXDpp/
8xp/rR7wgmJ9KWDYQRcDR/LMgCLPIDxxAMrH9xbxk3CZiAeat41IjFVqjdh8wwMc
z3TmkopCW+chmyMmyc4wQaO+8TpWaYhzn3PNP+WxQnZyAMKM4rii7wphTFeILAgV
PsG9Pg83ePIBsS9aAi32E34PB7KLvu22S6qUw/D1ViOSIx7MFhqzBkHyhR63QcaW
UoxEh5NU8b6PXZOUQGeiQ/+VY1Gz/WGxDKzWu1fmK+5uv7sAl8hOxopIMHubLoap
XJf8Lgs4ZDychMBkHBUi9acBJDXQqotfE8YloooLEMHFrmjzzW0xo9yasL3SmXil
Vh5pPsarWgA2Gv6xYwmWBtKprpxjY9qzmS9G6YRdo6f//IqorPzFrIvz9WDcw7wd
d/M5mxSfDGnaISbNU74AEaKv/nyxpuRWq71BNMDHDiwXHY/vxEuqOn4peKhFrWfw
KhNJdPlew5LVxAhH9o4rG/ZB8wI2qCSuugyPDUhrjjkd0hO14ZqnzHEeI26dTLB6
n9TUvbpg4Gtn4yHUPFcpqkxQSgYuaKyrE1R6xX9xX65X7FkaPqEfOrujdKnM+MEj
ZaBcxs3W3/ptnkcQbDEZnQldsLNR8eeU5oays2any6LfyNNNXvFkmaWx56D5H8dY
TCs6UhWAQvB1sNbk7Gc65uMjjAPut4GGxDBmU56qj1P8VCKYTbiwwunvyC/ADXYM
ofHwSXQFllYhJ4oFtnQB9uBWb0Rx5EY4lkOtyBFTYzG9UBE/ln66SaJiRdlP4yqY
iXVRMJ+X1fNEa6poAFo1BvsoTpSFZWNCl64oY5N5ywESzVR0Tb8DvZVKPWaEuPU/
lQhjMffKzT9Ceuwi+vvMt3cX2+rbBNbu2w7gtckpH/CX1XvRyNTh8+A/AmFBWR6R
DxWRpWHSwCEK1G2Se9PfCdd2J5PIXu+eHkXRkC/EHcmNlES9Fp/SNq6sGs59JjOw
jl6qIqLHxTYXZOw95QXBTpswod9QBfr6Sgd4f9m06vBkDQ1NUxJC9Evf3jyJBtgG
IyTxR5JGBCDapcxPyQPHkIbbSqNF2x4vOCdL1KrN3seIcYQxgCmo0dhliKAHsaYT
KwOtrhM4BTcwMuC1v9H/VE5CoBimw5Ns7HmwPZ9Xx02yhsnhhldHHw6h1XZ+Un22
PLCM2QIy1+4/2hMyz5Eh5bQ9GFfiFJ0tktUjfsxVWhOciaHTR4+csl49ZU+AVXl9
wXA4KAacgTD8hD5u6Jq3PI+6ZXwm925tiqb302VnkBEtAVriiD7ce9sop3Jx4qn6
4gs42lrir0D1NIhXd00766shJQ1Z2qKpuCpBNUpif/HIFk+m7JCSHn80ERb1Fzt5
cCyGxU+xxadljaVMj/I88xf1imLIRLXecAXGNY+ar+/v538PQHpio/fSH1kT4BGL
3GLOyA0G+4t9oX+q8bS24wBgV8+9EdQbo5e25hbWFe8oahON1fkZEocCyyvvFlnF
daIYfRVZ9UkmPFbnyzHeOV0m2bkLZmssfrs5mVIRZT53FoJkSYFoJE7D9mC/rSGq
UOo/mSE4SDWDOQDwo91dOKwyl4ao8GL717v4niK/sR9FwrXFOgc4uN2KgORE7IUW
cmteQhvw4MDf/yDDZOMoEqRhR0XcXETwXUqSriGXZ1vphPiXHSprsAl5KY4SDhmw
sck1oHLKzFR/a+IP+fqc7TjgbSRnQiDniqT3XdCwNJsh4y2fujBJUjEZAs2APLHC
jYTW95/zcPtBEjlnLl/izkfzCS8ss0PvIy1VZxW3BRvHYr8+YBtWwQr+JwhuFL8H
BwI7qIn7XflQ5V5t21h8aAgV7pVYZjtUriX2Edk7gb11axNXiM8BVhKC6pITzUmV
b+ioyT5i4Hys2kY4oNKTJ7jvjAZwlb182mXVqR5s/hAotbwv2UXYtDxcE/n2mKvf
5YM5JGTaCICF4liIFUIkqI4qCyFz4nUog3fG0688N7fx1mAzjn3+NvF4DqzMSz4S
/l57/IIRume1Coxcxt1v3/erJ1uk4hB/Qj7+hC6256iWKy6DOFGCk2Ed4XNUtG17
AwWyJ0H8zTNskg9SMXgPnZw5JdaX9l5SAaZr5t4eB3LMYHtoR3qDrKPI268kvBC4
Nw78YNnUTB0bMCe4knU0bUtPESKf0d4jj1YX58cEdHKWkyRRe22Fm7k0JS8yBsdU
ottJrcJmAGR4IfDr9Gb8ipNEcymNqdLeFvklhrmIKgrDCptKFWtukYzG8sa/jISi
ZYSjkC8UFrHeQD+sVWuK3VEeQ05ZcunfY3AW2kOeSK2i8OjYUiyaWSTf0smc2E/H
8cJ4P3U05DIQx8Zjt7KxFd9ajyzVA8XIuv6MS8Zj125fRe/ZqqAifb+1Xe/NuuD6
foUdRY2jREabhCgQ8LGvD60dcqP08PwSCjvNZaQtMUA/nVkaAa/LLvAfPw+9N7f4
kfknQWRAPc+eNvN+0qi7sVnxTdJjKmLaqXb6T92J04LPeuXt3cjeHUq19jWvzCOQ
XXRjFac1p/UqIm+NEBygMaI1DYo2RBcRz7i8j7Ywkj/m/oV4pG3tbRR/AkcG2HS8
WbR0v9fP7s+lQgOB5rWCc/5FNpXWaIfP2bP0Mt6g6e0IFK9j4gbx9pX5XNjaWNWU
CX4eJC4m+cM49rkvs++32p3/mrdzsyHlGn4GFulEX8s0awyOvz8gLcYP7kRKXjy/
XdStsqGUvn1yDX9vU+jcrgvAYdbjyZJN9Dh2piLXB8GNb+7u3E7lZ5QZQWzuunEB
bwQPlFt53CMwzoMSRWGcyrQIbJA1OTvO9mbMcaZCFIQjEp4q28Sr/EtKiTqRdrWY
B+GW6EDwugVORWnLeOLcoWJNEpEwW8Pemd2TgoCrIQv9X8XHGuh963Vu3RbQjl4P
v1s9bt/ESlDoKlji9JxRhssyck21ueUaA+4yy5MWqjdnaiyPBdslxRH4Ibxvwham
+Sfpu9zSXVGn2bISCuwsTwdc3+ko+eXZtuYDwaY0akjVFYK1VmSBrtAcG9evhXLx
6SYK5S8UlJ/F2MAHdZoUJ0dfr0u0bgolWOHmbSxV8bYonUF3+F9SdK1/R2J4sxM/
OTZBUl4qo6Mv/3yimnyiP5QQcy0n8mIi6UjD7jSGPfLsCJ5q6R+jtx61DcXh3xIN
n858uaepJ1tQbjOfaKj/w1taqDS3GC+75X9a+LV8dBvdju3zgNWJmptEcyQu1hxN
xz6Mn6AckNY+F03IbAjmhEf2/iMcgUPMaW8wTok9cpEC1/OJwa55VhVdqBNcmwA4
9Jud27VIJmzcOO63kNt7qRjgPUVXWocngRQxAlsACcHF/4Tc5xOEfRmDzngwgVKX
eydKwQ4w1Z8tYMpzI/mFlqBatHbYA6TpvfDqCvPxKzm2+/FKmYWJPLcEiYnF2scM
UaHDBUwtBQ6rUB0rCAn6mODHbBQWebQJALUfvyQDEPEBXInbSPKqagB3yD0zp2lB
dU2nRRAk/Zv0uMx67LWuZW+OlC1Izes5/nUwzCTR+0sGddKDX6ugH6CmjhSZZtwG
ywuVfDGzs6ZxayEsqzZKebvisZrK0FYMh1R76NnvguvjwruFKnkppkD9TZnaPGnb
M76HskV13yFev7nGwzEk6XnFLgWn9FUroc6D+QY1o0OYa5FfECZvDqE/i9WECfO5
NA2CRdjEzlgYZ8qlQk/yCzreLg0yAS/tA8BJU2AAJgyTYRpHb5xASljY0xMaAQwx
mjGZnAYKmUQQHxnlFViHAhMeQMtMJhoIzo8el8F+GozAZWrFQ4C/LKkQg96/wr7d
vdL6nOEY3BenCF9PSGjeiq7gODkojR8pijIr5cIPPuq6djo0GtOqqfeBiJx86Zxz
znMm5BvTaFLLaW5JLWS2Za+UhqiYF+lA8HoCQ7ZHS1IOATIdF92/u3ayCmTHdw5O
Yb+g7pcvob0YSyBXECEUE18qKQuSK2e0Ir+YIzojgymKy5Tz8ZS3rijtija1NNl5
UZ56eTHgQY4otgYllsI5BxPvJ87r2v0vyJo8gH1lP1bLFXQR7grgVfh5XzUGy0MG
KFIwNTSCRXDEAnZj00ZaWqX/maknHTpVw+d8AZ7CQzSJ5dRC8gNENAF9C4Lqn8MV
r8gIxwi2Rkbienext5xVijzBoKj/HNuI2gj1Ti9GKlAYjoLIkdJnipvhoPu2LyNW
R5Kse2qN8gJp5O7YvGQ68F+AsU010J+qEm4knsyUF5XstyK/7HvQzReCtZb84+Pd
goSpS6oIxj8yydxt7pk19bQ1n7BGVJ4fum6t3oN9Zbzhll/aU9sQUv9t92hbDvGC
M7Ff/RM4yMFqlY6MNImKjnSY6BK19Rq8eCrpEJyggErHq9dUSVZrb28TsglbmtML
j8+Mq/zNsb+WVOxSotJqOmtOlLGSKX7UiL/Z7IEmTKv4vwFn54l1uixLw4XHTlFb
W/IYpBtEVsw1esX4AQy+qf0ho5jrYIio9SjMD0JF2QWM8RPd8uHjozXvD3BtkpmU
d08Sp0WAr31zphmn0SUtu9Mlg0Dh7GzdMxhEOjBlYIrDOy/pMbHCYpcdWPvrPOKM
Msodou1F3jB0bb96u2vvrlhA1NgQONJo7vhng2fVJdhnicsPtUWOOrHisj93Gvay
Sngsa6mFFg9PIAQ+kccJ+ssxNYcnLmC9i3TTsZXAz53b9w7JRdUP7a7r0Qw3IVrv
jbn1hhUMnDlteABUvAAg1rMe8Ni3ho6rlKvMYPssXzwxgjaYXBdgrdBmPnWsw5+D
jnl73+AikVDkSXIPcH6eebaOo4vJTSmw71VNu9r79hG/FlNCbDGE7ji1gOsTEXq9
navT7qfSHkREHP93N02qcyOC6QRFKWtshbTg0K5V5m9cPnKP80ptl27AFS4EtGpN
TSoNSiDIeih3smZP/lXs6UQHlS2X1p8fTEvZa2iEMwJTJ19+RjLzjH7l9OFSUsAE
VnUZ02sy87Od8hvhHtPWKWEvtKbQ/z5u5SP75auKanHsNrxrh6Zf5paxTM/sZfx5
vdLfOobg4hqVDJQkOI/q24PSwYrTvo1tZB7fW/lc+osnt4U9zhKGUtbVDasMNMEk
d946cV1PI6K6c4MwEzBVA1KTVgpQtP557cF2jnfxy3TNAIu0nT6zHSt6+o9Q2RtF
G3DXiIVt+WAjjvRWu6RZ7Am9LH4zvqwWsfOsiC8VnAFc2TmghXJILtDaOY3ykFsV
AzeppzRBjixd+vwSSLOqb5HinzQ44BcwU1xoonQNBzBsEGcHC25rbWm7L8QfiZbN
1Kk2Ov7KpgcXrsYMi5tYJyhtdcT7qZdHPJOdm4fIuMpqS1CKXYJFMO2Zec16IU/k
G0LI17RYbOvlb6wYAJxnzmLJIC6Xn0fomgLVOry/kYunINIXMIXdNZHZ5Sq5hu5Z
td8Ssd61jTbgAXz6GN1yTvkY1IOZp/VS5Q1CDOt+052LRWY+AJrG9+zTaKby/nqy
7aI/xr6M3rwP7wjItIQisQl4LqMuIgI1yL8UzQ/zQWI7jyE2HLWd7H4/LWte52bF
Cy2fr0//cuI9k16jnqxwoe7wyq3zuPPT1vB93xrXwO4M2czVwsTUj1uGpblsryQy
b/yAT55TFjpf8uEtkuxNnWGk0KVQg3BM6mrthg8wtOUAvx5VAuzRJ9ULneN1zlPy
+LnM8X2PH24Zqd7H19+XVJyDpckpOcupb/ewIvy31jZvJBGT5XVS7MY1ocnT+A/Q
bnYeXGaHWcYuukD1tRx65R2lcd3oMDy3mGIrgevfJhBMov4nFcy3xsekPuXrz9Cs
s9q5x0Pq0frda65bbNiR7Q/A8pnl+oX0tQ4YM3E2uO/JoF4X/N9mHrx1oqr52XJl
fW0fq50nch8qRhMK2nGtEupDQkIj8KacfPKgI9Q1S3hvKw6KgBDVwYqZFKNmRie3
Mf4n4/hEiUFnm+AByzts7vUTmb5YnW9D7kFjjElEqOu7Vg0LWXahh84wMhvefz1B
GvOtrtihxMjCImfRoIakE7vCYppWPkgZMiRcIVsTgtj8E66aEgu943k/Tf7dU63g
Iyj7MzfOD4I7yOfYk7PW0J3ZiV26dnV2Del4nDxuSTW64bG1TnPf6aylqV9Rty+c
Tm8noWaDc851x5/orWCmLe2DqRgDVAXt79NFOaH651nFoSJfddf8927o7IQEosSa
oGDar68lNZqK+TTg4AKLZOhxjgn+0M8KgeXFeI3PVztbrSeZTOnS9M+SKMekjh2U
CGX6etB34LBxGe8VVh9OhkipUUZKVhYY9wvoccs9JBMJ7EFQlfFgBuGy4MHnaV9C
3037uJAUVipwpNR0yabsfvyN2seX9OWAnroEmPeDFkSmtddq9MNVzHwbRBAOSCqt
QyAFgoQh6MRI+EIaPLs2Lb333P0Hf5N1hgpRGNVEWIzW3qRkhKXpjpTQdBCCjqen
Rn1edwBg3uw3/42bjqveViUiGdaNoif086AsTmryiQ+BmnK8IlXVwNqBYHy6T1AG
Ddyu1NuraRBVxe8LAuH2jpsTAHxbJ2D/WVykKXWzxVhsQEj8Su4kv6P02vu+ZLn5
7E9A4E7SusSV1cXdmbkkp0PqQhXnxOc1K83UIFZ+S6RJiZEHyvK2E8V8gFAXA6oh
6h3Rk/Ojd2lpOB4B2bGNfcWkjhMKhMCiyealO7kP+VYiKAVPS2Mcz392kqCt5zOs
7yV7fVc3IjcL8sm98dAFlVmyn0rR0S/XoRp4uzbHEtuktrjriez6j0cn299rSmdd
LKsOs2C2zr4WL51oIHVCZq4fZ2C+uEC+00OajgsgEq1bCTMDppfywfwxHKYwoEpK
+tf3DHXMASw12Wlvrq7PMPiudycf4hbHH0gEYQc/X04dxWgwDV7TJiIsMcjV3TQh
HLl7l9OJhgosbEC/UFH7RCxHSq5PDIgp+rUSy6v7nGi4fFJ7NdNwJmPsUYZ03MB3
4ZktWT5tqKBUHgdS1LXeSxPlKRhrOv01yZaaiqQ/oDGJsSbnuEAKGFGAKt9B8PcM
b1NG6oXToRJ1QcU6kOcwih5AkHpCKWvjP8zWWSwRVNbkc8sec69QMfQCnQcEIZbw
uY2JqjV9VVmTxXe/ttvHyLINS6YhgGwW1rUDcVNo6G6+b8AY1dqZFZT8qPVN7dWz
DcvIFKHKvxl4/3QeUU/uNJtOjIwKaXZzp3WK3Own1Ba0cDl+6uzgJW/XZzDPmCsR
9iUW1iT3IL6Lk1Ojkxj7ZKXNeQ+45jNSkWWNpwNvmljUxOdzEyF0RwFo1jtvWq+7
H9vSYedLY6fagr8/CKYkHlMMFTbJBb6ClTs8vynOABlsOXxjJ4JA/IgRfF8Egbwy
HqTqpTLR3iAaPgiIwlA1+ST03hn92ypIyq6gfcKeM6wDzMW7doDkFz/vCL8lVmlT
wm7BnM66L0ArVFKU8ypnhepycPI1DfT/LkKz1LYwp+YihU6WLOm3yShPa77u05YB
z3kepjXbhUC8vitJUpKECGkcQ39MIT5lH6kDC++0bNddopzzxoUWosACR3UZE6vc
QeSIloMmdSwgsM/979+Ori8H9fzImlDqonSrjpdtgikOIbaa/rQMpFyw629Gh02U
AORPRzy61Oyruhz6Kdk79jHvgMk60D3AUVeY6mx4G/hbRJTRJ4QlKUyekt6Rx3Bg
aqk5ISbmd9ov8pTm7JVAHAY1vGCWb/iRFpxROtwSpVtTBn2oEWFZadzfoDEGAjAI
yp0rV2XbYT+NuYYPBnTUksC0ikAiKgGUAMcjmnT0zRj7/1XjqI3Ub6/NXn0+WBnh
u3kb4Clc6yj+6A9c+nGeFZiDRJqGvPqcsnpk8/J0Sq42NTZXFCTJMA7e3UV2m2rz
+voKRE6oWwRz5b7hkIh+U+OHZs819zM68TYYZRGK5gUP6day6BoVEzZU92ub4g0O
MbxsI3Vp8s+cw5bAwcKJfrgGjZba9GRz6BjiE3aaOLzONzmJoI3oEV9GJqyRdlHG
mWvimi/wZdGuEdwUi5lGNUF2CyYdv5HhuSn3hp5CYXv38YrTR8XaihbZJIS69FNw
Cei0H7Vcelyf/nM+m7dFAOktug5KpMnToxdRzsmrXaqkT55obRc1TB7c+DKAU2rj
2V6g65jxvxDVnmFvc48CcT58wX52ir4sntVyvGOSUKX0AUDmRq1xx6Ulaqg6AKna
lYoLLDZySBLaQ+kJRUFGE7KtqwzCokUpb152JLZv8Ad5o8w6WfF7MBN1FbeIAg/V
txu604p1WsY3xEV6Gth00Wk5TTJwKT/k3t8FfzMbCYlYivL088Q3QIZrH6sddJLH
DSUATatZHTLkH2xbUdx78PMeyKMBTgamutlbzpfbeB3UL8u0jriMDLHfO4dAhB8I
ASEPrTAEvlZSTI3RQzSAZfNG9AQ78DxrKtG3t86yWURPBl9ayOoAa22ZinchSO96
FvIH8bBgyjMyrvxE31l7NZigRCBpMe5u/usHnOm1D3R7w8tFj5vSEGHhwOHyAbB1
QWttLPTvgXHu6s1QVCGlSseikyT/E0/ZuzBgEX3iiHE9dubIvGHo6ImbDuWlr+cl
z3RyL2SfkDwrwFLWv9L6ZlpC8kB+uiHZKNLJ0778T6PmWy9qbTgdxrGGv4TV9WM2
b5Bt25Y5fDugj13X1RYlJ0zxAqp6zgukACiDbX1RFdyVXFXq1lH3KGdiob4az0pi
evwHgn+9w5lItBjjAxAXH8DV62sHB7JJ82l35ZGRGR/aDdxXfW9zQGaTBGw5SNwI
gV16o/M4w+WP8oYBvTypeeck3aU6AluztWHe1kAjXaXUQLSf8nZArEkR+TFmH6FZ
iCNACiDqbc+wYpFphSdauQkWmr+KbvfGzOg45wLwPGrVG0/dEZp5Pqw+ronm4AoP
xd180uB6LixYW0D/33vdFYOCKw7ycJKBhHQZ1xn7CKJrSrDxCD7u8FgawNBQ1jZM
EXqFz/75sybNEMMeIqBDqX8pkKhyZLZIE1XEviXAivTSBFGCdhaxX4FDTUT9Lg1z
Wg8Sn5f0gKfjWD5avWyvqmv1C6Hodm0nZK+JrPDrDwpwvZOQjm0ShqxYuasbDDbD
cCJ52EwQYOgOLqpVjbCj0ZceVi5Wk5EbaW1vkn5fIzOeAUSp14WJW5xkflY/5Jcu
4yK6frSl9hSoI5lPdPOqEX7a/0hOYzO3Gc1/JRC/3BDo0XwkChCO+updom2TnX45
silrm9CKjOURAXal8fF+cC4rXS0VkUgGgaCofiGZjXQLaXBjrZ/JgfWfyIjmDY/4
Cpcl6hIjZVO4GqVzFB8o8EjEV/BMKbBm4HN3ZHa+yGWDpcCypOCrCSbc9HsKKjQ1
wtcTuHl+vYMKaGfqMYPgeFwT32qVSIszDsZzg3c3YxOpDNoW6p2FGr5dvW5nuth/
MtKy354cnqeU1oSZ+dhJg0i+FqyFEjQMeQouczn1qkbk2e+dZrIQLZAc1Uof1smL
Ofb07t0YMjfjfiU3etOz2zaYAngzhTS9z1oNDcWIH0SX7FokKEZuP81Q9L988ddE
U9uMSCMlHUrcF6Bs0SYFLsSfSVhvBXdPkz3vJIWljj9p5dmmTzqhlZAfefeK2dbN
C5b5OaSY+ssKCg9EpLmIq34HNWduqVdntbtglZp9wFlDIVn2nFR92DoC/gFIrQdF
t6AAnJkCgEemAKmjbheXYqICJllM6Dufm6Ju/TStiU2nvGrj5ZarG+tuECKAO+yI
bDJAHoaUcMCJ2GP3Lzk8fSfqiHqbqSZ2XhIa4R5AUnujkwvCbo2cOTe2HK+odoWt
PxJHCj0y+YU9qHEZ2uCujfKVTl+KHYdraQTemIfzaUq51ri3kjeG3cI92alo0WWv
BnbrvPmgNTawBp/A3exuSBb3VG0gLnIOoHvcCBuBT/0QH0AW2RVouHZwQNYkgago
zD9lbEcLla5IAIAqrkcG05QM0v3t7rLRtvbXXHVqz9QBKeMhpZQ5kZJbWyFeO2lW
5vBanAk6pFpkhCsEF1fQ2fV1MF58mxtXdJo80bzQxMaTEmdbuyTQZlngsZL8+wVo
jYNLGz7RRK1ifekNkgb7eSn5axEjerYgoE8qDnW4cuDBYBdIMeK6VfrUx4J9Ow3k
oVzERGSwhpD4dM6NLzV988HkJ0LJW2EsYAGimPybSALdPSYHm77ie3wa9Boghzv4
T/cFCwvZ9FJcRu/YYfr20QaNxgzuyVHqE0hOuzqqu9y7h93vfTB2Cbj6yPk1DSNH
ovTIWyZ7vwBdPMdJQ3WG+3HoTT/4qEUAJsULvtjfDfhulFoMRTXvfTRD808+z2xy
I68qWP0n6wgDJmcm6P6e6plIvm46hOxUUpdvD/hr5RGuuIkAM8cMuncDVMiSsb0N
Y4FR414k/pvEJJNBiiF18VgzQBr3y1fd2inCWjS2pE3BUQb30yEplHgmlEE2aC0E
HqzIFP8f3L4LxS+CtCUmZzWrVyO/Y1B3HovdwZo4hPoUktP9hpnwiqElYa3Yh4Y7
KmqL3ASA5dNSyXrzoToSDMGCZJxcfVQwoFcCwlbm+7qg4GAa7KOIf4n6AQ37netJ
TdNhZDuAF2Ap0z3wyE0YN93ijWE7Bkxk/zsvta3D790dTw2BhAxU2Ag6IK1zwRgf
f/Iw+EHDdt/abhgm+q1UTPl0v0bS7s7fzJRAeTP3wYeRejKMjyfpIkEIvDauM4YF
8uDDjMoogPAtp/+Y+buTJdBVpe1MZ22AXDZMJdB5x7v4jFG/2t/KUV/smWt0TKRk
HbvuPx7SsZREYDSlS05G67qFoM1HeCrPOxoAvI/hUXLcg6x4iRMglEcxQsQIjxol
GriskFjM2IxWy9mP9lWhzFlMK7LtcvhX5D809hmdYOkrUnxYxr94grzt5BnuDGN0
fGtCk24PTiQKtEnaKUtQJy4QNC+aYTZw5hk5H2et7B+mV34g7Ohk9ktkkqoGwLlx
lI1huYzF063qZvxlsglxv0AAYgtha8/KzeG7TFF8vAaPKMAtDQcgtu0O1ip8scyE
/9rzD7Oy/7VogqW+GnJTUQrZz6geJilAi40ibj4Z7dbVulWSpfydBKobo9QtCOov
KhyfjDTo/8amaLhJCt9Fj/T+CVBhNS1VxmtrPph+sVYQyNLiVVON38PO2fZ2nrir
ILKJOoNG1GXQ3ivrsm0hE/BdIIRYvWXCfo/09TD5PXSVArAEBSRzRhta/LeKAbB/
9pxE2np0HjlpnryHcJesfkPTgGuhMjGRiUC6htVFJdLiDvBqWgY+L8+qhiBh2UzG
iTlWqagMavMnd8zSrdgwud2kOqpjB1hcon9AI0z1vgS5pLjMWWs36FTde66XmGSI
Wm6wOWbxv0MUl0cluZQzOOoamp/8/RIEBtdlY0ofHF5Hn8ul1vt9Ofq2ptD0+vkf
6YAPI/Nhi5Pz9JGWTuD2bDksJgqap4w4smrFXCAwsTOxhh2f9fUwkuhdon3u9+Tj
ykMVAedaQWcHPTaug7hGtFku69wbWTo123zYRb/1+Zy7MMCruAICrzYbS5hWai8W
pyGFBYvUTRr4QJKAX37qXnOqrV9pxzP4YhCY6AJjVz/tCSJSOgL7CLzzGglRMCou
TFhy/I8q8NMDAq4n/QzDprCwa3AbpKz0OmncF7GQJwOSddHHz5kU98UWVQTvGHut
D96er+0SfHciYGrslvF504Q0rAAjDTPfiULSfGpJOjuItrWGIFWFsiVxzbUbe1XL
p2HOxtzIh37wEEzv//PGCwlESJ2HsELLlm7sCsb/gLaHxJOwzp4N3n33t7HHN42/
8GQXwHpiNZnIIq7QyWKdwmTtxszrL+XvDsET+rxs8UciQYtMpCsS5+KxtxDVq7nj
WlmiAtzR1qXWCvrDDoP7mva8QgTuCgcIH1sfxALAUF+A8uzzzvFe4kGhQpHH6wTw
7AWPN0WTGoHXqtklzHTwoXFzZsZUYp6Gm8kv3GYCNFrPwQVndZjNcOdbywQbVP6M
lK0PEBvrNca7o82UJd8dbTHbCQ4vAXkGMM1/FqO8G6Ht8DcCbgFF5HBqtfcXaOL1
+cwF+HVaTGFhCHwm/C0mhyZfoSinKHWkxosNC0GAeWYnMCZEOxXbLB3L8GdYSiTu
HTAjPd+8tFve+uX7Xl9ODu6pFTukwNZfrBk/jsrppQoFbiyn/h8JIMcB+TmBVp3D
icMwE/fbQ6ykFqjpTSS+qMDPWNesVfgtZfUnGgy9gpkLVzmQKq2ZxsEtM07Z3URA
Z8rPmGdZ5AzjfceP4R5qb4+9JThVbeM3WuNVp1c853kgfU9UKzZ6N9ouAHOFefY2
aRhQHD/ffmH+mI8L2aSDcJ4WsWeOp31VR0I5l9wA9FHDFsgQ9t3zLGlOS07lrQcG
jdoXnHncfy30YloviAf6ijy32TtdevxHJmIpM1Nqg3wvqm2pOFun4iS/HzDnmtSS
LuhTEjKIprf3GHY1nj47J8aZMuyk159i9JZE/WwityMe6oEkQILuYCfFMryrOAdx
1nL44WNExd/LO2/zCrQu6BBUd4976IpqTM23dWplQ9KzSMM5XOzSJQGHK+ClBToy
K2mTQSnac+KOcNU6FdZKjdVXVE4okt0rZSIm2qSgGW6Ke0z/uIO2yeLXx+uYrd9f
rQpvnpFffiPX7HfHzTFipO4MFLDtdM33bHhfwPBvVDW0eX0WTE7MPKl2uYEz99GF
HkRnOQ7upGk3dElY+o9uU196mPhiuJu2PCS/igQ9qOK7iodPi9aqDpUakAPSvAk3
4exfNKXFn6eClS+dPtlH2rGNrLC7+cQykzcyqpd4+RJKRXRKOlB3sQVPFr/j1+zA
CdYIW3TzrX2sibcowbmCRZ94uaQUkLw+L68p5bX2/jNe5FUCMeNljbtOk6cChI8n
HDDTX2j+sO6NaJz8CXtoREt/vCAqIl1DXD8WJOqiTiFehpcrfL2eNbhe1YJkxbfw
C/8uC4qM3f2ls4M83VFwqL5FdcCzPL6AeFMgsTbUVf6rX9AUCRUh+zy8NF2nPqb6
IFsx/aZMCiY6JA+OfoKhsjc6fzj9U2B0FB6cQn2jiRf/WEB41i+w+WxvzAp0bAcB
oZ1vt7Vr/Q86BruqDhQorE0qWEbfJi0EhfYqUeYBLLdnRKwROiGynKq3XfbwuZpN
mhW9lICJkMFpGFjE0AT9wdfcISOWOlokV/LdK89i1Km06jNAlrU2F6GhiX/lOzBR
8aHPuz5MZjIA7Xttx33/U6GRNjUBoAl7HgLFHxaQMLUQtzRr6wGcwCXKD81trtmD
12xJ9AvIyKknUZLceoEmEUgla+8nN0ttIiihJmBL34jMMud8eS9iOaF07wpBbXOA
fBs2/+ANzMwH7aBn5Y0waLE0WuTT9+2AS84G4bC0OLiRK9tdG9YBLBLOwFzHDnxG
9VC+w1VRnaVF4bh9W4sQotcW/PbDYRYnRLk5kqFkK0RI17vCR8b65T0AUVRIpGta
qmgBqxP9XwqvSOBxng5GLqsyzn/zchETZz3UmwYXu1VXqWjLozaTVsXBk+gPfEAe
YfEHoKsl5j3/jHZtbrnjJdJcrW2/YtZQoHHcfwQR/EqKjxqnP6eJvcvFuk2tH5Wr
dKkyz2/ouZZWeNQFJaWO1uB6eVE5zPTB0Voecqb8f9nJegNnWFyS4+Don/GgrLZb
xPCwVmWxdz3qRKk+qkRdv1Ym72QXVObx+AkOlcotqhetwnqHwTT/MET4AR/1rOpe
+xk+CHLKEHFiypMNDNC9UtsGAGy/vcaqmAshRgwv2I7if+luJZE6WbTuVziWZ2Ya
i66qX03olBmOKxTHgc7NjjClaiYatMRxA0Vuc66Hcu1fBzvpfRLkGN3a2XmFRUhM
l6PzQwcckZ31dyYwaZqHNzk+rlcjKNJKNx2OXImCe6I9wC1YUfTYPXnh+IUW7XHm
xw7l1ilnZ/A32mIIc9sk7Gfqjrl6THTN1i8mOf5fJr6TYIQBRQ9NOCIhhjSOefnC
JMKklQ/EP1XGrZR0n80s6iMhrlIzXOBu39//gY1l6LrjKpzE+rRdjWrJIoCYauhz
8aoG1zGSzh8YyLjeODurM4IBqt5k1ZeKuNmBJaHNBmvFDEaJSZ4eZM5bolM36Nuz
9okogb5pIqGwdxqhxH5LeYhDOX1wbldqJ5mmU1z0Um1vD04D0LMCPZQcBdxYr72b
gqYnt4EBJ80L9kG3pFPYRT2x6JTxjgLyqxIYMOi1YkFoOYWPBxUickBdHzkwMOIq
07WiHHezm4rMR73rzMYWEpUeYPteLFx1dUFnVTAaPkL8jo/fCCuSuOmplQNcA3AL
3QBW5tVIxZSIAlHPk3lGrCFEH/T2KJkczBwyCVzi+YuGjUPWuB2iQ1wvugKTfwZR
/Sx6XyzL6WS7odY9bzlDp0LonSKM76lT3ACl3f92rrO9EpoatrW0MHubdA9fopxh
f3fCsLhurHG1TcozqMOWBlV4gFDFpTibN0jp6DHnQD1U9CWRCPKO0av0YEbUJc9j
LWROGzjJGfGjhPAwOidrJ6Poe/NnbeqZt+aYaGXXD+nvvOnURMUtiWeTl6fKzr1I
if9H29c58zXykp188rDk2+B4CJ0ZhT+EXJwUZdo7d3fyNtpQdwWCh0ww2QJCnzVN
bSQBGFPNcinV6UELRSxhAYWS9sLDjYois+fXCB0e6wgjxIwm/Z6P37GrHgM0rZA/
eLUT/IKD2wpWOnUTeNjIjA4hSwMu3mutAJtkOdRLLvWldb9zFktxduUs9KzrksF2
MiOk/yO+XXHRpSZcbrOOKW/zHob5hY1dmfSenejnB1V913/OKvg2AHXrrUnCsiLT
OU91iCoJ/ghV0wCd1hM7WlUDsv9uvjqwaCWa2FxCLBpWCe3gAenoL733kaDGnZR3
8wWtb1AXZyI0sQl0ouB13JRSXvktzzMUi7YdJAH68fUx0LcTxDlwnyK68qf1DMif
+AFeZBs5U58h+nx7gbGmzj7EfsAgZsvaFZnZXFaDYDDSO5kodsO39luyVo04HlGa
JJ6pDBiO1G9blRt9sjvySpiKAiY/TuBfoMvIIuVV8CjLOgZfajE1yCp4WhVBlB3q
ik1jEX9vtDbDae+qYQJPq0ppkYDlez0fsHpKH7jirsCfzZAhBbJ/DjjO9lzLJJFh
TRAK9j5zuyT6RmB15QZ5/NH4Kek9psWvAD1VH/gMKp0SEBW3dZDsCfzigYmzhdTT
QROoG3YoOuCROQdgYWNbuoCqOYy0ArXxlEwqP6QkZRwMy1T41YlFo4uE89s7mHjf
NFislUPlv7pl2UQTgNExWQ5yh5sK9bwvN7Oe4Wdu3NY1/u5drARwEslJv9Xvv93e
7pEQ4Npqfd2tWq3yZOyXM7pp0Nx8DXX6sGn9mq9GyoTTdhB4KoyQQmJGOekHEc9A
zelPJKHG0yH+tcZ3wwEr2vh9RfkuOaavqc20CSagJWbxkFoM1dsiIXhoiFlwS273
8Mwe7Ah5veiEg1Om/YBq/WADGGitaEpnbFTQNbqgkVINslTSofVeLc6spCofSIID
4JjdSru5UwTboEq+1NnIYPfkLsBFyyeFCikxo2fUSAPzTh5dwTAK6g108md0yCPq
4fg0TOB3PDFiZPfr8zLoId51AJK3hdRRU/wfziYlbnIFQWUdOq/Fi7afopLdp0gB
mkHO2q9GnATJ+3WpNxxAoM4ILf2GZeFs5ZuG+YR2h2GrhNG5xriNLN251qeNLSe6
LAX7WU67UlIcGKrrwpM7KZkoF6f67cEZxJlb2kOjM9KVm5zFYVyLdLpYJ8wR3jCy
pSVTVZgsETNw/Dq7TUIIRMh5hnxS/NKKsoL0V61NXD/8V//xs0ZicRiLV0gQlovJ
sfx2VplV0pexe1lCxcRdTmkfUH/M7nubxd8J7JcTajsAqTNL00rqCAZtVUQgQo63
mVi2+6uQqB8qiE6FUKxlBu9C6EcCICLkkp9RfKb5FCuBTjVaZCWc74dsIJn+tVxr
D2cRLdSUOYz844EvXlBiRv1IL++Zx8g8P/sIrZYNsvJBfD9sHWFRmPg2xf8xykDe
e7miJS+7gOUh3V2i9XrSJk4e7/0CsPd5QGFbkHhY12hgb0x1dCOBfaWBV9hrKwyB
d03oUXmbA5dtD7nBon0XeilgBZBibWmUuzKgQ2lVJX+NS4UzuomZxs6R4k9xCQX7
0amQL3W8nZKZjgo1wB5zNjLTCaSC5eaBofVM0vVhD18o5llHBRV7QeMqy5KCfVej
ZPIbigohLydYOjyFxp00ZKcMVn0t3LxjIonBaCD5VVyXCiQgJKBXmuA5jVihV+5i
LISQwPIbnrN5Z9RA0tAh6cndYT36nGfHg0o9AtZi07k2UrHsPODH0NK5bR18DVfG
GfpncpEWkSff6AYy1WhTx+tGZhyI/bYU0C9YtWHqaYnypInGJyptPblrJDaFJfL0
/drwWEV13BZ9Gt3P3+2SEjo2sUIZVmC0chqcJgquB+x/DByKC/6JHLsmmC2PFbYU
Y1Uw2G/9iylXLYKADfdVQF+x/fyQr/sKgFFgnrE8vFVsHlGRpo8yID5fiz85fkPp
xqIkDtcmVtKnvWgxguUNrloGVu/X6um8OJY9LW3bglTiF+wIKF93ooGVpMOzUVwv
E/1tDJ7uZK5ipfW5IsW6+P3fWEtSpmq9KBGMbKdt6iHyNzfUytFNK0cGx4vDlrU4
B6MmXCjPkAR8PC3vmMLsKTA+gtIfPFtK2Fz418jzvkCKMroL9BQjMcJVjyHB0ynq
VkY7IOdzoVZJtP7ZvtZ3CdxLJfPb/rFPYH47UhhcQ1RBlHNk/7Q6nJQNyQS2oz55
rF59hQLkLTgHvYTmp5UQ8ph7VrPWD2tc49jtr+klDQySwwwBAhUbA/BwPq6Yr7GW
kdLvvQ9DOXfYu2/vzBr3SzWuqyfdM7rIgvJETbdeuXlmciO5ZaBh7vaaiVajs8MI
U56iEYWYCRt6qT5qqm5ztLo966lKcsKvbehRW9c+8DMmqKrMwUxaTAD7c0NoYeR3
9/FOhpLJyMCWIHTvsqeRQoC6yqk6c9fYAFitU/62b8T6l4Rvr7EiTR/viQW6OmBh
Ovfas2b0YLC+ZR/poEpTCvmJd1hJtSvkPhZnNAAXNaJSbd6AjWrh0yOGX1NFbxCD
ufuEU+pBGhBUc1BdOEwPnfSZG4x5PggmeEHeFEZ1lth0mec9hZ08LN7XM13kFLRc
/YiHeCItHvu8nlJkYg7Xzbw6bo+BAL6uoeZjK5iSpKORHhNNulJPwtwr/WTBqReg
qbtuVCcsDP43oleewDttonxZeQRd4rQg9fc343ayL8ixqpeBDk+A3u2gN+W1zj+j
xTrkI9xKTQSckunNwGMNM5xEOfdByUFvzIWvgoRUgeike1SlQ6nJwCUcXgw6R7I4
0GQeuQVM3Kq0qUTVcZLM1YaxeULMdgCq7CLhEKsGkvUmz6d5yErdX8+Pcq+syROD
V000lV/4STIR84LTbgh9jS7xGCpXlAhY35qy/0vzH2YJPo9+FWi+qYo9Bks4SB4T
cTxLOZziP5/lCzVqAgk0ip6yy21M03RB0E1297IG0yE6Ev1GDJA8tHYTE6Z9kQBB
VfACC3UuVvzpn5eCksU4KNyuaKXKIHizFZSGpAcQ0krtAhJWKWOGS7keVExL5q8K
boZwODc90kGfS41XPJvbXPCkhbO3VIpqmglIPtVdRUF7aTRsWVct5+RuCNJg2WmC
RHRlcCucJpiONTa0q9WHs1Jp9foJsTgayi2/bQW++VkeW8VTR8SaqMZLJaiYjohw
CYFbHMJQLTguXy5T6Hf1LoWjn9wpVhCP5BTDLtdwCL59XFra7RCbsmt57192z0Lt
fdPzjwc+5GQNC2CKkLq7QGDluaO9CXFLscIQR17xrpqgIcg9TNTQqqHSLFKdWBIp
HcdbEpgB2ixGmu1TFwvulcr7r70f0T0FuGAFSpUBj0JDeJrE5S6PIQS/xjyjVA6n
anXtHoOLapaUp9Y/NbZF3Cjmf4C+vbLmYifRTGKAEz1eYGhFp6yJ2kGUeByFEQw/
PpBVIpHg9v81Wo9yv95/eimVzu+BRk0CpDOLkyvnZDQkUjo6305K/SQhgxHpIu0a
kgXDleQ0uQdzi8wpSUazuMQTmFUA2/zDiju27Hg9kOSvv3C7NGEXnWwaRu31OO6e
9s3iupwbo/g/8AHpblthCiF1/1+7Gr73GPB3DblNFNcNgqH0ryVebEtPK6ZKlFbO
ZigBQ/0iF476FOFl1wiAA8Hkw4vaZXQEI5Aevf43ZO3/0SoN6EKtVUWUul2wqflw
VBkeQX/brma48gKNVrffeFBl9F+gk0yW3QESxMUUO2fGjWE2OI2JE2ev0ibMVb2F
zSHLNWYUc29d5RbRvFl0Kt/UIft2rvb/Q9w25Sny6OGizUMFhC6pXGv0Tue1HW90
N7yZ+o6vSHRBP8NqMVkh5oBbRbMx5DZwneg3jKjpD7s8sQ9bui0hI6Bm1xZU2eHd
larja8156iHknSL/ZZb3uRDVl8AwZuCK5SOCVJEunZy0sorZDLexAKVVQFt8qxX2
gRnTH5Qq6hVDUnpXX2MQTbtu/FRmogdisFA9yqXjMO/lZUuYcDb7sZzPNwgdEf0e
DIn2QK6LzAreqDJYrhjON9eAFf5D5pVG9jqyCDz3nn/RGQEQSvZtv1UnfSjApBqU
rUG+kUvihGN0N9+Iyz9bVIIg0Mh0AliZW+eh7jwB2mVUdgy7XvJEXgzkD6evEw80
Ni/Wehv/Ywo7PTUL9i96Br5pATRhGtSta11F8v8BNZQLpstsiEVuLj0Vh1Opmw+O
Fs05BeG6QLzpg8ZE1OU6J1hb/TsUs5fGQ8uYinRQmDpIqCEFyZnds3UcIVf36JQI
2u66hEjE+VI4tJahsn1frR1Gp4TmzBRyJAWCzzzoKeigDjKpf1PXXNDDjWyR8NK7
MDq3ANUEoV1FCVVwTqGazLofmA0Tna8P91dptN7kvIBa4rNMXUsDpZ0ysPlByor4
5nrkf5sVlguc0fwoPNseB9H9VckhNQgJdk8FbfGwGP2or2So2sX4klmFB4qn7lTW
0qblg94IgYLhtupDnUsBHtfucKBjMGahtA5zdqtQkyYpW4p+mdnxlF88+sWg08Q9
U2xFcW5EseTJIBhsC1wC02gNpSqqYjeYdv5AL7kzgmwaDCe+/5M7DCnNppW4Mwbn
hDo/PIs59b4sCtZ0VIFqr6V37tuxdrxRrqlYSIiY6yd8AJNwBoLt7LFv4ZaX8gfC
aX4k672I8TCvbPNyeuWLsQ1SoidEqF9GP430mKJ+iLjH26lV7jGM1RkvSgU0ABis
Pt/5S6Xckf1R04ayqOmjf07H4vVNq+NQWUFUC/kw8bY3TePu3mpDtkeshP9pAV4A
8QAFAs9RtU6fv27zKWvwqZDDnaIMG83PUwzMh98E4R87ZnOE4sd4Hj55yiulKY+S
ZrBDEQkzTjtVzUnFM5TBMlPHp7QUnFV2FRmBO3k/191i9pE+ZuwVBdl3zf+1O2GG
tCMgSZu34HBhGc5lESm4dLDrrRBOhlptKdOGkLh3cGGXCR8eeZPk2R+fOvlVfBQI
mCbKU9t+vlDRVFB1f8tdER7FfV99ofrZ+4Hc591jZXKv+r8UyRCkHDOKo8mE3wIE
OFhDP5qbPYHP5kdFgcLClDHVbHHjyE4w5oimowZNvMHW/x0KqkDhw2vaxZhRxBga
B3xSQI4dlBT/dWfa+EQfzYDHsyjspSVdvE3J9F3jeRPeoSCjm0OHCQyeB7/dAhxq
e+pMEtAUdTVICMI6pYUsE3rdQiK5bjAMp190bjuvi1R4gJ8iDWFyoH7ruvvYpZJm
kAgpacemYUcsAk3e9MGlkZ+DwNvvbiUyTwYyoA/qIiv8xXdrZfzVUiDdKVqB51rL
kTrRezVKReRJKev+sYUoRIkBhfi4IwBPKCLI5W6aGdX3kQJZDYzJ8LXojvAmK63r
YrUPQmLM+WCmWf2lKnk0J2+Kaii/B3IQ+8iPEpjyWXLPT3A63q9sZQ9Air6n94Qo
PF83jWO1inAgmR6SobFH0p71gjsnA19+MZmOTEjI+7wvaCMkqwACOiq3FQMACJop
dkyYDLmPU+PwNNH/BlpkP96PByOg2B1FmvkKDuWeT8TYSKLgG1thhGeQuniNaAvJ
purypiNEQK9QvZoJ7+nLIsaYCDuSOo6oOwISymToD/OMTZV2wdQQIv5zNj5nr2TC
oO7XGO7YCoVRYpOIf3zXPxwXgE+DOntid9TnN8dREaVs/Z872pq3PkLkLhA0qQm1
nzEL0q95GXxfF8hbWCuEqu6fBJ/7B2yAzAlaJ9Rpnldn9gm8tAXFEUBrCtRZAT3e
ZdtE3qtA8165pmZqbvQXv6M4IWAfWC6Yy681lKLLIDc+P5TqnFSOUKJzpDdU4uam
NeYhR9RKWB7zVVYzPEeeWx/LQwppNi+2Y+03O/JdIQ7uHAvubmOIJlbqu0+CGcjp
PZO7UR0YwcgYVJtEBxzrwGHbRgYZwCQwzGdS1apyN15i2WhUPzEuDRavR44K5lK7
hmuBB7e9sIzlO42i0eXzg9HQhm8ytKoXlCLnS/lLC8WfrkNGMy8B1zG6AJ0aE6z3
5CckYGoBX9oMOr9J8QTpd145OCF+291gPfF0KsTepbe6/56zJ1X9QCBFdbf8mxYB
VLxc1mk+0Y62GPi1fJRCZUuHalxC+/J73O8hcE8igoVNUorboUcyjvfgYO+mNi7m
TzKPJ5dnNSKCjGd0ahq1s48iQckwnY0KJWN++7lB7EvBhvOB4YQfmE1MawKtcQeR
wZHvwOTKsIgGFhw5wZz6FyuVnYzh2W9OdbuyScV7RvPVjIsiZ9M4qDw4z9ECPI7+
9I5PzJC2/BtmwSycRv5FJgAB8U4UFV5NbxwLJ/sDiDfWYbHrEl5nOQ2kP1U02Qqx
3uuhJFwZDpq2ZVi4e8x3IlHiyvQ/+dQqKSbUKAxd7AIuBKfPcvkgkCaVMjJAVg6E
6GBXzJjIAu/Tv85CJNuY6gRceBRjVNLwv+UqrmLyCEFdyO2mNoNseirgeyg1DBSU
j/zQu+KyBx6NnDX1zG3f8jFYmBC0XzqurBDAZDT8ngwnucuJN+klDge63nVuc7cK
miHLkOHS5KYG6t5oqFQS1V1TKm4ah5xuL8gAEGdNG5VL40avvSE1f+ZeIpsYKRHc
YmsFqfB0mNM/NCEmx8JbeTgzlMMNHfwGWPIagQPCobREWqgsC1wPdJ+Z3vrgzAUr
Add4XdXzOOV/XZ639MSBo+UB5y23/ZwFkENyd6jnrx1tddq0OI5pH0VV28pe37hU
thFMwAmhrJ4FftwIVqHZrQ6NN9jw033RokZEEHtzWW5DsK6JjmmH91YgnkymOUTt
Cwskg1gkanaMlrFHLArvfW1sTo1ps8C7MzO0+Mk/Mp+T/k2Ywy4fB6rvshMNi1BD
xEuoWG213LukqWDMTa/RpXYFPc57V3mieZcj/CxhSJncnhFBqVpDDDW8XV5hHQsu
tGYtU+luNHDoHs3GThoOOXq8UP6Y084HXgK7JvuLC+9gQrL5kRcmVR4NLGradTr6
LouPuRXD2PoP1lS9cyYFQCBsSKt1p3eXJUe8YCXZfzmsjqqoa5Np8eYRwOp99eAc
TRvcNCwTGoFvd0qR+Qyf89PNh1kwvKZQPO68xnfdlfHduJDfsNIPFRnPlSqDY3Z2
IyxN0Jme/48fF9zeXiS64rk2czJvNbpi2EzaV7Pl1gW1JmJ7mDy5Gxyu3x9zoY2g
P9gdnJWynNpUgqXoCUhYZPN/VzS2QREJbxI6rhu45/4/K2c+Gfxb6Rtrdtf3hHYI
yx6ZR9/D1DgKOOabzKzZphkXJNFgRmyvofZAk+263TActwOuH/u5Uyz6PwrCdQfv
D4Wo3NmpT3B5QThooAs2u7aJuOJ+yesGcXC/JBB+K+3x5rs/CDxXvEEQS+zlxBzV
lunA64gOf68rvJOGkIOgHn7bx6nxwDg96zl8tiVzUKzgw34IeXAbCDkrFQl7x+In
6HzZpAummSyboGpNwVIKoU8wvJ4OSbQ18MYI5LwthxlJJf8CAMkHcPkKlkQTikR4
4Az6sPdp0XIjUvxKq6heJCCUS5xwS8RYEilO9U75hhHQhiEu/KlOi2Ka9J5xxVux
RHtuJ7VnmZszrqTkfUPTQb8FU7Fc8F8FSFZdePCkr6ZFruNcdGR30wfHY7p6Fn/l
BSBATa9ANkwDN47ts1KcE3iOmudHyM9lapSbWcOw7Frojxzzhj+qeOYgwQui3364
GWBIRakl4ohkKLMiPUbiDr9DTAu2ytHZoEPq/lL3/xbnoD9344kWsS4ydTFGGbVK
2igFSfUlUmSfQZOZ32agc2CSNY6+vdqp21mhHwGhLQzMoaV0ck1vBV0+IrYwR8S6
v63cfFYHl4paAj8synW7JwNW9+7UndxO1OEeeu4JGAUs3Jv4etKo2bVKhu0kJqwC
+uKEMjpk8XNUeUlWva6LvoCCynL9XRYE8d1buZY6bo+Cbm+RemORs8uqv+4gUMeI
KsX5p47GEt0NHpzO4YyrkW7HnlL3I7YlosChZRa8n3MOIkm6nNdwUu7z2AQ0kbqA
/PXSseGwf+tUcMA750d3GPpoZBYtEeYX55JFDIiwEs93UoWI0wVgiUGHVYh6rTWS
fCJ+jKr+1W7sGB6Ak+V/IPviDn+90e34hicqZBhBLEY1lAKNtZRxGSWcHtZre2vR
qH0dpw1OtpIqVh4famCGu6TNYvBojDH3bbatntWJDUGl365ihGQKLQtym+7aQalA
8cFrm07bFbnCU5cY3CKBlvfkJ4yysaqJYbBDigi/Lhj19juruCooOQzh7uhmcXZE
oyoIsrGxj90G3pO5OFldej7AmroQJdnHjOaH98agiGMiyh0ITdTWKdzJWlI6rpQa
gCocV00tC0KQaSGLabUFLXn48zyuBaijkZ2dQgsKKNpep41WbHcgGUKLLihkErwM
oFcAnZ0RYdKNYcfNl4EBNvCSHAAhN++cNYD1YWuLOjTYrzQEdWWCtARujl8T3Fnf
dUFp9StpOckIpjIFHpX4cmeRv72fNsl2so0SLKVkrs95pqRFLn9SkjriqBzUB7tC
thI6cYDGzHd+elPi91tWc3nnTxMP3sQkmSXHw9rAi5JOy+ZT4Hklw1mu3yVLRkRt
r1h22wPAok2iV8OLJPkirxYvcShfx2vg1b3aQvcyzWHwtMWbUxZ7Cu/tJ7haMPCS
yeLo08n4Bf0YqiKFmr6f2YYMmDyYGbp7SfLxlf74SR8J2Ms9QcMw0I8JSFItLz7U
6v7ul/oSEYUjt8jzN2cYDk8CgsA94rlFNdVIO0aoPqcwR+wR+Tbu81/5NVc9nEUW
qeRMHGSkl7filNbH5D4oi6MHVf43MHr+Fub+wQkbWtY+/D0cN/mbBZlFlX1kiGD4
KhtbcVXte5Jl0hzzpr4WMiXpB85kxVvAT8tuB3RgCetOa6FnzMo1dKTVCWPbeRcj
xMD4JgVBEsiph6/iGmwpbcHuEuIqs78yyVqeeVAF4FRMHg1j1w54F8Vqg/YJcOfm
VOWbhS5fUpBUHGaeI2lwPC9NsnFfALCcmUeJv24lkGhh4AwzH1w7GMakZ/OeNihx
61BrGE6u8Z9/QpnSIUqJMIc11w3f/sFGYqx/xkmy/yDCKfIq8LktjwoVdW0m4hww
xpeBEUHN+zbRnbBh0QTshkSMJ25m/Qubr82kZ8qiwmBZuYFjNh+hsJBQnJPZeqPT
9yGcUUd67Gj+2+2zTB8yjcdnE9tcgq2NMDZeltIWr+vExaGHhF1XAtIjaLu9wbch
2d34nwm8c7B9p6o2z6k/+rbZvRSyLLaZiAjtulSUqcfu3s6wbO+EQjyGu28qaIqw
Yqo6QoiCfBSOUSyddwo89SKFmXA4mkKCsjEogrfPNlokSxZXUpdG0PaF+eTF2GoW
Zb49nBdBXh0S6l+XoqWzP7yYrb0fxGnGCMnSsOp2UnKNMjWhiPM4E+tvucYRe7sN
u3WTfk/oWXcY31sDIg3aeVhSHJJqmgUgXj1OcS7e5ohLPu/8XP9EGPmcG41elFMR
w5MJqV1jNJgBiaUZtz16wPkmh/xMPKAPEWRT7VEFRAwRvzu4SIrCR60PTVjeOzoH
ZtMNHk6KZ/T1vxknuHCBi21QkV30FLT5fir+qxBF1L4mtg84RvwGwxukknTVAcYs
gTzp+TvIcYei/6qDYs5eEd2l/fF15UMi9iRcKz7qA4wnCUJEcLOK8XKM1IRJwi+C
lI83N28/AAzYk1m8YaYad+QmLJ5uRvR/aJHiTCnx8ahfLeYHypSVhBLhPnV1Jvwz
8IX+rPJ29mnaZ4/2uLChVeefM6tMH1+loDNoNO//gbya5Ox1toOWSxfbCTX+6UCX
YECPRin8ODMalh0AnnuIXUncT0w8Id2G7U+hiWWObp5gwBxTDnf+eyf8zZRPD3d0
PGreWwu6g/PMjARmVyLrN9AwEW3W03y8J/EV1bus3NryAbKr2MYF8jT38z75X5Et
iPFYj28lCAsmEPauyf9zMmgYC6K0c9K0GkJongZeQbx2wGGw0v1XmIUrUEH6m5lq
Cn3auS/fCP8OitFvMOX54OjoBWZFLUC200gcnB2JeEg4M9PxUUiPjaBbX/sDuxG0
+OV8E84C3AtuOIWy+VG1xpwHHy0R/5P5XUb3aiHo8vbolNnjawVbSTEzBPPphJk6
g9ijuSWM6TFTAh+zj4V0DdX1/KLU4Twdu0I2+Cjp0aTkVTZZbYfABrWvo2wO+PIT
8xSujgBMJlq3fN/lUHSOqEaPhC/wNF0M0JKReq+/3oRsXeI9fZb7JBkwNsasnj7J
nMoLBkKt2IMmJYlH20XFjkK5FB+C0uFy47NnefjNAEQ/K/66nuywo0YaWd2RouIC
Vfnz9usj0EVf5Bs8siPEbDkcLdcmW93ZYjJtXJW0B2Odv2bQwpVXhdYjaDtEAsW3
0gVx+x8wpF1pcvyO6tRp/KXBPNeiGoKaiEHmarFui5A0epufN2gcRfNYeUxg7pUx
PSzhw8foLXJZ5ehKlOY+Gjw2tc/q6BZopnPi6s0JBORD8+dLRwcSrOxlpYkX+Uas
ei7xqclOx6+CVzzosCOEmt7quyH1jj6+aMEyj1dGo7TEAEVDRMqV80Wrp9DEnnDD
heqXFTZ7IUDkxGJy0lNqMFLAYz4VAUS8KXe1PveNf3Kyz7hqwhU5jOM+1XikG+cF
Gzz5i8AL+t8lP6zlLYbLPdbnuQdWAWNk2VkYXSewQT4c9XGnyL5ffS0KVtgSb9jn
I8TjzNZHYGkKJMGa5zt0xZzNlxVVTeWF0F67WyiIfNOIMhz9SCfjRRJ9eDysvFsY
KtF8AhGBRWlD6xXzMiOAFGf3i1uojaFAmfgW/JDp9xruife1EkWlfd3257sqJDbk
z9BX0xQfnaueZaBFq/1VdUPmeyyjGZob0IR/QEveNAG5uU5IFpnAhElVhdHOLonP
P119KkfI1TcC4mX+ThqnfJ4gAzqccuAMHKe5a+FD6mo3tejBL1UIhpsNo2GeY48T
CG6w5Sufn23esSiVwQfO46sYZZeAhvSn4UY0YCSlpSKWg6+HQ0yMXkhi9CBLtLMw
skQOb9fr6xRRirzmYMqvA0ooNkoa6AiUvyGmdlaetAIiAmhi7JHra8YB+CS6kwt6
JFJ3/laYWXWJGkIDlo1Qo5JTw+dyMT3sfkdrwePX/iKo42H0Mu6ziKchbq6W5ajG
8Qk6/Ms0L7kM/d67AC4x9XYKw13LOz+2e9HlaISRSC2oVMqNKrIg5hy5+JssVmpR
rRyrpYIJWCSIJFb6ao38aGEDzkLCcuEif0Q5GpvkTb5LVG7//bXXnraKCgP28maM
SIkds1ZexxPK+jIiIZWK6x+bD7jQNX8ybyoY3lupNYx1BowiYM6oAJ8zCugCsQm6
Ggt6YuawMgLT7JOFn9o3TmlpCkvPW1wnCr6P2srWVThFgBPfYVkiJ1FxP+OBAmWH
fSUQVxYHtXYLC9LrbrE9qppJO6/aZzt1oHSUiJCvP69SpwzclfV/cpuw2JtCRnSN
coQeDciu53PpCpvhgx6qZtncz/Zd7nxsPRlB9OdPDZHq1Zc/kcAvKKsDudAdI9uq
IUrYzasOwdtqzBiMxirVzIMIAAughKiVLzxc5hfKqwSTE8B++bPYFIRnNiB+0jkT
VuNAU5frZdq//GupG9dH8QNSLrEIslQxjwjKq2/jMBltRILXNGMRB0sUyjSq+6Wh
VdE+/KT+vdP0cSb/OCuth4bNzG6Yrv6f7KHnqi81ehZWRqcSEH617cwEoH7+PFZc
7kmfhYT/7QOsMh1U25eMqHhff9M+agejOD/F0w0nohF/X29maO3+Wj+qmy/hAvMy
E1r9MqrfGil4otzwbW25rCvUXiXJz4itioxPb1mRc3+Fu8e767G4hshxjkhJQ1zZ
IPdTDhR4qrLD+lP5JhNOgWni2/1GC45F430+j8d5OCHmZ5zq2QLdDffkEoSklq4D
PvlCR/VHaHvDvNwFWnDKYp63rOr1rrCjqbs8hs9P0PGX7ar1Tf3TlF7G32HOsQvC
YR4O0L8N0NQoGjjzEP/zH4yhSWN6f5SVv9dqY73wCCIe+8hpvYdoM3jvmoLIiia4
CmaZS3vcSAhFYnJygkS/cDZOsxDzJo9MCkTVIKFVU2FJIDjowGwuprKdYuHLPuFU
l6tV3T98HlSq4BSZ0ENgG+Hvht+Uui1BG9B2Zp/7SHa5Ve75Ql+5wyt3FHRNAjVE
A/OEHK0UV+27l9uXlhmHdj80m5ukQNa7B/kjmWQ/XvYV1DdmgtrAqkEuERfocnia
EMieq6YbpZoogyOrHdn97GCH09pjoBKSMYFTpQgAO81yw7mkoc8xYtC10jSpNMZh
Nd0MKgnrIrcX0Z6VmkqM0UF/Q7b3gjQHp68zjMv7Br3kYbXzNGeTmnIn0Iw1BaSO
CTjcaiCOpMAUXj3Jte36uedYrdozhQIo5II+tWf9AW4tmNPSj86AgZHw+B3eiUlk
02yC5GXGe5GYDNiZsUCZ8uDPx9g7RUILSg3rhnqrah/qoZOY5ow6/3bNMMY0dLoy
UVa1xyrW1XsYCw7tveoXIU9FW/dmVq0XhXPvikRzk1RuiMb8gDwFK38kXvg5T/E3
aSSgZfgKYH1PQt8P3xg9oo4zSYQf+ZYQlORPSj4e13JBqtxgzqQtHvRW0ODPKqRC
yNOwQFkP+fsBNRPqStKyzrALDdBKF1KT/OqrsHeCg2scTokReZ5RUw1BOo+KosVf
ldY+/LjcOPCZaRms3aoS7rcyxSB4B71fzYoQUD/wdpuZkJBFIpNqa09YEYY0EGZS
H2F7ob8nIDDuBDuG7/Z7MooDd9VM23Qt37mGmBW/BP6+lPnET8GkD7hzpgEQzrSY
4dySYr/cMqkKalJgt4tQEWXO3BljRWVmRBoFvDQh6Pr5U2vLXaASjLek8n47TAK/
JNMsH3JopMW2QW+u/eXGkxCMdQIZu3wC0kCN2+RpkXfugtFkNNCmflERuyuqfdMk
/IDq8dT8cecdoLvsXP4iOMaghCR0jnV3pCKKJcR0PjnCbztBSXUfEIjtRCUKAFyd
HRHR1qXBxLjjM1LV1xy/y00DVCUya+evZSIYyZc1n/Ohlnj0ljAyG4t+bjjWs9ns
E1xrxfZvAuNY0sA9wbxgIIsN9wEL1IW9+ItXLpLdb2Nk/8QOM5JQxePPrG72FtJl
6eDp78mkrBtR93le2gMV+//53E6HmVThqt45ta4aQKHW0Cu6DEvam+FZSqwWQjYu
rmGGSDTJDDBoedS6O8zr70tn+voViVU02iBUZZg3L1nikPgpUzn0i8HAwwBQXYT9
7d0qV2YqwT50t92eACrapMZi/v4MGrg26WFdv4YlQicRRVGt4NOFdvsv9dlbeXuK
LpbDibcrQExgQvBqtvRktmlukv02UvWqzwhwzM1Ns+Jk/grR+eYbAoTD8RLON1NX
rKghrpiuX85r9ETLlKkP2vodwYdAcjFgoav5h/kZhVR/nEdQbL/H/x9G0JIRJJYK
ovGQqnkDLlMFMannUZkAheGfaJtlZPoF7pQ8K+xoStXUw+RHRIovdJqYR4qpz+nL
MHj93QO61rZd4X2LYpUCxdWEIyhJM41Gcdy2IsEhRGDxn0bGmpIP8zPCLjtyKOEX
KKLdauxRhaQPO/LA6gcMnjFn7uX5SV/UaKSZrZo6XBsoE4eLgc2AIRNPoQ+NaquX
/YXd3ddpFDBelbuuKBGBVzd2sksdfR7lQmFIDOh4LeOkSt8xpg4CYJ9XZ+4/1o9Y
nffkup0qFLYROoHlVmGY1RORJZ/swqFOm/ZrpBRZ6lT7gGApNMaGx4yOQZn5T+T3
pNm8hguPI1d37ESXXLxf3cZqofH8EOYuRveeCBBi79GY2W5B0BGjxAGi1Mjhp9S5
My66Lp0N+wvGcR+X3IDOjAoyJyqiM+7RDsBWArAT+b6pFiU0mUcL4A0Kg3LFyOgc
+2vr2CPSHMJgaechoaGfzaRo4RtPkY1s/ZFbFbJJ7HjP2ZKsmcD2mic0HoD1P/Uy
PtBgiwXJMt72d1o9+p5LSgoHvaJefST25RvcroTh9KUbbpHGOSEnARvwzgt0w8lb
WNb4jfaF27C8sBWhIXAo8Os1ny52UyoQxggsUisLuTIgbPAChsekz+KpP3h/lrGM
M7p6NlnKFxJ9BT0+fFCGEMOYrnBOTSIzhVesD9oKXI0reHWEZ8clIVKmSp2juXbm
aR2O3NGv63YFjIj1LCP/zrgeAOK4u0nMY+loEE/0TbN7OXHfWhRIwz+ykqvICXGJ
NWmV6I4Vp5oSGhcy3N3fBrQpGRtT+095wXY6v9OFRqaKvxfgPP9ExvUcM2vGj8CJ
ek5QoSiX4CI52CCqhvE40Bu/FKuxpww0NvNaE+x/i/VMKQc+buwhfg4nDsQQ0fR9
+e4kiZ5uw9T8W8WM+f8V55ql7eU7xVnHPooorJBRGav0qPsAk98T5uZOKvJg0kw5
Ocey7HDhtbJc+WIB4gfDA7QJlZYxMxa0LuI3Q5xRTaourEuRkMOKcq+tQcoIiyi9
CPdJ4ccVSpapM0fBTxLbFHhqAdnmPx0EDnCea+l8gU9X1fZ9dCV/kAeN2w6ltTDs
vEYmIBccjp+aoYcT3EdESqqqUK16X5OVjMAM9YA2Jh4x4Ot8o6pSEyQKfcqPMjP6
DLEi8Tc/22l1CaR3ZLxelIPEX2FMJTcSA644t/d1jFqYzsRoqubDXjUkYD9lPO8A
aSmUh+tQDQWH6QY6VgYJbcTlPSuTYRqTLKUYzZ5r5DXa3kW5tGstB4Y2kegwDHtf
p/IPZSJlnoYZg5K67EIeW3ILgoHeaoJqpxeoZLfvd5t6msvx+Sj/3pW8VJk4u3+N
k7h8b8sJ6mM//gFb/lMyBDwE0CFkbhq6kll7ytlvuqAor6g+21JpFLDA7eDJOdah
BgYLlF945S+mvWZW6IRwpPxhWMBTNbfpPZ/xzOzofl3P6ikqsoWHpSIgrBFRvaLK
XUbFtcmGyVyWdpkGEBuyb+BZsg3qVLBim9G/n7TEWHXZr+wyJBY5cOpBOypafvef
5/JZAACRffaptj//58YwvclqggjPp34p1lzRSua7zW9yIGahBiVoiP5BJedJfQ9h
xjDlH70LPOdKXXRZFlbd8yiery380qUwy7Rg8nXJUP2uCj06TgqvjjHUcrfHpXSl
26gLX7PRPAFgGD+YCo9wzr2kswzjmYJhgaW8b26f1trT9jOj/slsssQOELfLbBt7
x1xhD3aV0Xf8mxEzmRfIJl7fmsCGU5ImRrvcAx8dGMr1qU0gjdsnLKb5nDViRMQl
lNfM8XW9mVyZWiFy2hSCy+UoDt1JgwW7kprPQH7+do4X2aM6oosDq+VlzlA82zI3
0+cZsQgWG/ikUxoIO0cK26txcRjeMxvnUJzMA9DTNaoPhjdMKzmzh6WC1lm/GDNL
ZrFsYXrPE3mavanysJrWxN75OmDnhrUjc4BkJj1VYUXWEsS9LLp07U8yJqd3ZuJf
0Ox4mT4tkwPUcKzaITdn+hcykBmVSC+7Ty7v3oCaHMNobe567MkV7Co+YQeC7dCR
V4RxN9t90/olhSvYx9XmUkdQB2xSEtUh1k28VHSDhjnQ3ve0eBD0YAawgKx+z6fx
POtX+bWKDEK/bu83jExAVbp5udrIi5FeO/8qCVxIJxm9XcCsl6RZuht/b0Tmtvwb
RnaxXC7M42R7ABtqEJkQxMR4wvTfRIePUwiQeM3O7OqnUk8LG6k7Cjqln+nrmUyZ
ASoyIi1LmCwsJEn2iWh91vxX/kTt8f7iX9E1V9JBo/kNOe63RvQ+25gleUQg8Brr
gsNzhOPX02OIjpjskK4T9ApLoJRIM3Q+ZKXka6lWKWwXA0RtEy0ZGKysY9mMpMRr
/J6GoSvKJEWJ4pYsaGnvVgrb9fyMwc6i0rxjhCjc0nlHSH25sa1qqLeZvbdQ2cdF
npicrH0kgZ2jCr0gT6CuNs6n+y/pe7/OEBwkHp7XuhOoB2YDq6jcVWvZj0OXD5KF
7oGTFXvPsg+UEAhpOmQr6ZkHXmry2VpQyU9TQH54tcAXpf9/eU/h9ySkcSgNsMnJ
jjZntsKg0CQdsW3XymZDiaVt0u1B4kZ445n6fO89wqzqEYBFoE3QdIqyd5Ze/Mv3
FIPW6fThFY+XB3QxsgiIU28MDvQP/kpKkH0JnpjegNQHTCRjNZXOwdiLBPI38hxU
Ha+w6GfpkkFjoyS4p81dYLDNwUdEU2itIMYCOGk4Q+x+/GwtGbwYJF9FZOtYEAX/
/BsElbgAa020zPX+hy/B3ES08q2G6aB2X/2Q8JWfCT/SpTvRCzIREAjDybL0qYzn
oJmsk/q37XcshwqqY9R82N9cxuHAoqBo6lWmMc8GRpcwKrHjni1loRqZGFOPJ7Hz
3xBCwCLquCxrNIOBlBIxWE5pht/CP2Vr97PMGmrs4CEM8LGjrjHl6nuFhL/5MwS1
RWRFU89lWP/uvvNf6eTYmTMBXaW/nZqH+JCWHRU+p0VpHS0DERxajf14PCYraKHG
0gGrSiG3II2CAusS4fI1fiyzEClgPILupCF+M6SKTDGTe8oriim3lzXgPxM87kdg
ai19y0oHjXr723zwg4Ne8JqZq6Tmc6JSxUtbg+pe2X+f8n36UmRbZEm/ae9lAkzD
WJEcwCa2rmHpEkmzUdZhcXfcVAQKV/9uUqzm5i4Ew2tDFxg3KnTGiyob+y0GGZg9
PTRMqYBVvtlwPQpjbY+9/E+N7+n4mowjqzBjNiZ2vnMj7cMnwMtcWfjMLoWR0CJp
GcvbGmBjEFn2bw+6MyIr6rK5m6EdnFejcIVGhabaRKQYG/b+0GQCYd9Js6qtde9A
MougyoEOpz0qv0b+svRKL7S2Ureqhdn07M2j3nr8Y18AZh0wwsvw/M9+IRYLnjqP
UzUxn1IJQsb3nlZNhj4CHl/O0CARk0v25pG/PjQuv/KL74hhwtmfxFzo5BBnP60J
hD2h/h6L0sQLQ3O0uV/KBB9fUmb8MYFTeUyuFe8ohkxUmCsKsR4a98OK6OHnqoXs
s38EthWhKZ/XOMB3aoVz7xaiOKKmWfSMeYn8Ea+P4Ul6DpLBPjwyG6YuyCcZ454A
0kNaADV11+sn+JKbixeRjCUrBQjOpdJUZtV9SUpIHvq1YA3VXd1CAKBbk/YnnZZI
Bu9fDNepOfizFO0tT35Xi6EiuvDNwqL6etKN8EQbtvknCvCH8wch9WRbvVSfogDe
XqNnRlhbcldRgU1Mh9Y/2WTZadpIZRqoA2ftHatxkdaFaKK/zUD09l6S/Bz9P2lu
O5kxACQzRxSEIuzjtRMSQJOAZgehR2nTLIowSHFifJ6U0uhP5Td9qmrLWAoFtWRx
eI+EDdUOafUzUNMsA9N+OKSBm/08UqsuPnVLofFiidvIuuP6u9kznM1ztv6YL4XB
Gh+UiP2nNBsuQ69wpF7X1l24+mJ28Etk2xAPOXkh4NDzaWAxYE29noRtqQVcEPNS
MhWVCYo4jtmyW1qxiuwiuWrwoTFtdoRSuLly7d0TNl/1I0+ZbowIOtD7HiOts7e9
uGaH9ivxcD9rMl+Bqzhg+Z9Z5sBqrBNnUMHVJ1e4f62sv6TVRH7UTEdHp6BPRcXy
uLEQ/wFyedQQSfVDPZKYabe+sZ6vAhbf9VtJtQ2QM6w/8u7nOijAoz7Jmpb8kIJK
GCpwAwJEdI79TbkKoGiOODe5gvfq8or90mz9GxTUvttriCQl04O97miTBTdWWnM8
eM+Z59e6hI2xM5ffN4NwZ/qaaJedy8K3MF7lk+o6cCaIXBUF8EVhLqX2fUHSEefK
Ms1vENu6pM5Ga/h2s1qwuhls0eRuydMn2QLVAWyUrmC/O0T2GqVI/3kpGOucmOay
HKKW8kvFn7qCRm6hdoUY+5fTKxaIfqVYC3029LvtJLwcozsSoKqlZi+735AexLaO
6k9QulcmpmYf2E98AHbP2/4CM6qFRudtVRj1plqoes5yrVWnQnjNcLn8UozQfKOA
qinTSJlojfwX2xfyy1qADdnV9/Utfy0zqbWV6OGHqjHla5ItfnP8UfPM5jUstNwh
TVCjFVTSwhVm1fngnnb2b4wiQEWlZG8S/P57lZUrdx81/U68Nq1L1BYur3VOSB+4
ryZBOOYM3G87UZbGYWuDjIJMWqN/uq/EyOHMLzkoB33fh+qsMZdktBbXXVl04LvI
SfD7mIwI6advRP3yekEn4/l5vrnhGtLHqXQk/qfC2JhRMYIoz7BZTJyt6K5tVfQ0
bqItA+lAGuD7o+0B6BJkQgh0O+mIAT7whiX6fYA0iNDzGzcUNf9w8mdouF5KxZGP
snhxsp0QREQ6IoGCA+twRCI/QWAemFN2nSTrwPn1J3XozT64Itf7NZmu+Cqr6xEf
Jgk3pi9iJYa4FdODTdxXC1P4fNUWBwOBRXAVRm50VUsv5abt6IGCgsCKytoJA5J6
fzURE39RXUxE7Zv5LxmUMdTY9vN6+NiKslEaS9VZTFInUNjpvnZqspFLRGLkP5fE
p1qdLmrKAe1saUzdbMkpxIzXBbbDSAkjzz/W4jesNIRzJqvkkKyt/wGvs0DEs2sc
xGWElKpdBUPeA54a9yhC1IHq7ImBX8UeX5nugqF3QC4yIJViW6FdSQ3HMmvl88o2
oB5PMR6sVykJRkxduUtH16rj+sRHTjgJb78aeCgoSDzct0cyy1dLAPA7tww/RZs2
ljX4Gy9Gb1hQkcMSrk+JCUhG+R5hBYOJ+e92Kw9tUK214cQKcBwBszhmByqcw0j4
DlUJUiM+ZmMT2U4NguI7XgzRcfORDD4jTylQz4CRCtu+UpOBhwJvo/ShxYMtQuEk
Iz3AB13tNdhqgKiaZZFBRhTrDSL2Uzk0cDoF6MosO4jSS78Ml6msRUNEwHPuGDxi
YZ4pHO3n59vUwN8L86Cc/chLQQGOQWO/R2U31kdLt9gKZSJ1reRFdk7oGVRCiXz9
k6l0oHBh8RgayohymOoNiBpm+lavJGa2ArsCa3eYm9VqupwdIknC27yTQF3niHzO
KrQT7aTw3S/j1Q/Ol6/cIBU+MSfs7d0DeK5kalFU5R994y7HxKbKIPS23UkT/Y4Y
Fg6McUMky2eR6ejnNYaJXVQR5S20PDqRr3DatXzyNcgmxXYNfwKgKoCErLnUG21+
BXY0YP0UKWMTS6d3dn6maOa47n3s7265ngq1V7EbN3ZsLJecZt9T4SIaM0RcApHC
v6kpOZ7l7+ExgWJ16dmTDpgkoJJjU7kEilVcZjZiAHqKm5BThiUJQUg6LlMA1dFl
C/zMB5wK4ShAA8QQQjM4Ed54KcHSKKPHtMG66K7oWEuwRkNI3ZZkmatms0vAKB59
Y1IbvNP0ANlwPXJgnLVAcY0Yst4JqkPKqjpnwqp5vjUcE+cgFFQ+whR6pzr1XVg7
fe0CQTIuZi9zTRP18WfxSKJdVKwAWVDs3dKJkRnulCH6Qvywp8t3S1PTSj9G/6K0
6MVoC8cA3vpnEFYZ5SPUHGuvH7g63BNQJ2zZe2SNFUTZ6dtDR2Kv3vOhiEXwL9QD
sVe9LsS5mON4f5jqlb4ylkXwllEoIiuW8sLwNcrbm4STUTshyMkQhpTuGEtgjNnK
v7BmyiRhkLonOdVIyiGrVFNyOAyJXGZHgvV6bRBkF5s3XaLH2xStvC1+62qhr956
6dW/aVLbcQ3YMfdYnMLGfSnjaVyDCm+G9Q6CwztEX4kkukG2eHZU/TiPGgl39khN
c2Z4IupsFyIuutQ/fBFJ+XRlkk5kTYlpIu/Alb14XZTdCuCjQvQ2Yy/Ccn0PsxaP
lX85lbERYVJMyv0GVS9Dw1qg29vSCBw5lDFxOCk61j/yX0sPbu/xIfWL13ktPmf+
VkFkXbX/nTlCEFcjDvo2Rw4GeUI9hGin1S9gkBaGBp3TNrAJvx5DPJlcQfZIel/B
dkhWxcSIBFBwUkDrDG58RZDbM8X2gHR3lN9AWcgoKFxMezRr+/GoU9JolRy07LdG
ofMoo52yw8DNPKAgfjbc8xCVDPLt/kScyC6EsNlUtfWqiBsDZmWKUBg+I3/JjeD1
c9qqSajLijja7UNI34tzhSvsrcz91IGnBYE7fSdE8s41bHNAQJcUxZ9D0IL8kwSG
BNV2e3qtU+0wHNyH9g+2LAW165yxnJLsMMWWeg1t0OVOiImatdHpK87PkN8I9TuK
pLzeyGNn/McJ/neIgUK9yXkRgYMxgAblXt0jpoLaty0pC4p8p2qCMwOFdIDSO8aA
WYxaFPSmF2CpRTIF6uDPiK7t4WWh86PJ7ZEzBxMvj+ETk/5ZHAvX5j0KNezrNa9a
wcHT2PJXAnACn6XiAl53CZEnL73btDYSz7aCwFPWu/oeMEy4N7zh/pn2pk/7/1OF
PTndoESwio7DddhTNdPqQkA+RKIzfams46S/9ymiiQ9eTTaJweLbJ+1AXQGV0AWi
RuzWhyDYPtHS4PrbMbNg3lBflTKwJtjDqgfTxy5oV7SVFyitpqKUFBkB1o9GJ2yr
y+h/7ND4UCgamaL1R2pjyo4Oyx6GoYopMjRU0qMEhl3FD9rTq1aCkolY9Jji+R13
ei8IoClyl/edtmHl5d2rt6phsC8qfcjshpVIhdz2icFDY1V2A1wD26t9kCvndnMJ
N2Zr1WPYowIRVHorTRzP9hR0uIVQ+zXx3ZAFuxFroOBNPzW17//Qj6O33LrBVh5D
pr1DuOQMXUgaZzoEHt8qJLvuLtj6WznWJ672p39Nl52ewPqAM3BZ8p29Pm8tw9dT
764AFKRDt7MkEmdlNm1cHMs5BuhFpGpFMLtcEiWyhsR0M67RjUIDyfA1XY+TffJZ
l+nOVqLBbTNW+z7Hi7SzQF8fvKtn5ioiJ5+uVQt6/L0F8rhEBb4IggBEjKHp5gXt
3XSj+vwO1SMScrPM/PXB/NTJFD1p92ykRzNOjDsy3idqoV3H+myMTRa4SvR3Bw0y
c1aP4UXyrPHSxX9orHMlOmkr6WnTxJBFm6cJDiITw3XsHVbKROoTnUTbqGF/NtyT
9FFJvrozk5FZtrarMvn1ivIxflah9ReqXFmkA1qOKw0WCRugALqpGvo6Qn/ziOrB
+RCqIQs1hCk+4mef4YxYgxXnbmJXzOTBDdKifE+51p5UkKGuRwF/qeN9xyQlwPji
378uIdL+n32XIxs/Yr8ufnddhcVz/4qmmm5bF530Dv0tWFvIM2Ls7ZeQk9IskucY
MXgxl6g7SCiTWb56R2BddFRQEi2GRbcJ/82/D2CXOsvdk85qpxy96nuHcaRrDSV0
yTYB6EaNiJUnUSWD7NIvFDuJu154ftx4ayri8r/OzmGQDuIrZhbBqkeCN5N9ydxA
oNpi/jSjdaLEqrHn7j3eQqynDaavF12IGuB+/6IGqb/FWo1oSbaRoZ1T25MKNTJF
LK4cZRtFvG4IicaxoBOo32X/nkoXQOOkKY0mpUn6M1ounvDQKwyTA14txO1E8rYd
nYB8fqhAwQ0Un09dhU+K73yR0MDF2jRh3geRqpgBvT8iXE9xwrO0D635xsdeRzxW
aE3Qm6Mo0qWRChRwd0YoJM9P1RWD9Z6B3WBHO6ogZqqBdSocE/wZ1uPB6sX07dYN
6GMXlUsmWQM9ZRFRUSgFWL6j9x4UNy0c+ZstWQM39roiXRrY36bwRDdWekyDEswL
ZDxgM95yJQtDHG2Tvaj4r0oynBZnysPfdwDn5WRvK+xsYEzcevg6YBZnabWsXpIg
/qwauUtteljA2L+EA4PhEavtR+YbcUN6h5YfV73eW8qKu6L7r7nRPNcuJYly8BTg
AAxtglY8sx/sUCtUoDOXjvXaPbFWH4OtJPUBYYnL75DlsK9+osQZOvutDvNi4tOU
wUokHvwuMOsNNgOe4YYEthQFbrrWudjq/r6zvsfouqioIrk/s6va0K/oonijj4yp
QE7CyMiTAWXPoAo4jOX5CElTYACLbUws0oh8oMmIlPsGojKKW/L4NkN8Yl75wUcc
SCKmrnT1bBzsXImxR5foGmi7d+rOYJn9yr8EwU6rKkRAxnIa0esLsQhpPx7HhMjP
wrfH/DsmRgArN+5a1zRYmS7OVk9HNj7P4EP5D5NlPusU8Go++t3gjdEbdyTif94g
QkzI9R/jdXxV2af7Y76NRBvI7+8nhwv6KHOvGjiaekHxlJxt6V9ecg1f7XR9UnoO
aJCJhgPvsrLmBm7ii0hUDkdT3UIRojdVW/7YxEbWJFISHze6BsjxbwlzFj8eTZxG
u+sPhHlcWB/BUvRxprHsDO6oeuuexxIkhlNKs6KtXK8kxQx4dzDd7gEVIQGolvV6
+8pFrp4xDfTDxNv1PwyGLtVLUjcXWKSq5OlRgGADbyVVmlxu2IFMn/gGBvriGqQS
L5Rq+gRZaFmrvEyA8Gzq9wub2J8UPrBUKzTp/ILAEARGcyJzP7e3eb3eebplWkbg
geDkuw4hECMlW7j2RiCECKy894SFxYuGHlAhkWvjvMLmilQlnK7QdURhDk6NpgGY
w/ge98PBXs7nyAuJjhyM+NnOS3U5GVKKvsQ9g2F4Q0UJFM12NJTrMG7sum9O8evD
mgthauTHuVv6jYo8sVUu1SbhNZkFkzTHyOsaVWD3YMwB9+p34Gt/1WAZeoZ2AMF0
JGLt1pOB4VnSOD6PgR5sITFXfUxsaEaDp3bfXpR3ReMMOdqMsILLFKf8ht6rQDTY
peZwblYcAb3eghC2Hiq844Ovawr1RnvQ0ZX6cNinjt6ZJYXS479I5owrwj2uME7e
nSgYX/+GfAtz9elgt3u2WaqzZnw4bd+SFWYbD/f5e9i2R1MnwWxMVqdbxJCOxXkK
LYBdZ/eaFjNoyeOox617qV/DMDD5F0sw6KvyFShyvSOm+DuzuBGAKQl7HwsgT7F0
0PQZ4zXJefKbrOs9mqUlPMbv7rQMbDw+b9HAy64JT7+knFDXfUiaQHVKgHNqhHof
9Ze8avbKMKuuhP23qanfI2R1V3POehq0VBH5XtSnxnVMO5kVAjBeryg/Z0AcdvlC
xKOGHqAjNB8LL6FfDu2Y/CthpR8qU53jCS1oc/jzzMYHk+GUHSdE1bxg8ndxoSBZ
D09EI6dfsgpEwY+LkLWtUmN4fj+fahfDX7nEVPEVOk4z57UDX8bpLXycTkcnZaHJ
DoLL1YMYtunbXDK19OpuIWgB6BbSzs4nXktGBxOSc1fwlO9KB3RHlkDVQmsyC20g
5QewdEFSIvmNRGhlj/53/qcsVtuZHSpv0I2Kp2HpZ+9fHduObMmLV0hHmgpM4AeU
bkoh6e6Hs34CFnNECAGxHHNxTdVY5aAQZy2egu/gNWlrTZzX3S7Yx6iB8AjMRDV5
VhV2FRXcPYqZfhqfjiZGKANRPhrxQC44yUABNsrNlMGWX477GEJR9Lb/ufU5oBTj
LqPmGrnMyoGqQ22BqRbsSIAablWgCebzUeVl7/VuY/9lhCtf+8tjp2qQA4h4hGDr
nCkacv2ksTjRr/T6UcM5KecP4FV4KzotoEJ5tEXE4r5cWwCi2hEY1Q36VpWch3Ze
Lhi2z/aoU+yhM36p94JTul3eGhU/oEK3CZeKEUrhwP2JmZUEctTBQZW5YelNrvDB
hRaUKG+ReRbpH7IQ4SE96cAvMgMfV7eHtbLgB1b3O7yKrXBmKWoPLJh6xe+qf46N
NOCCHeVoyE2Fr5V7XcsVxAGb5WQ1aqrCvVV4b2i9ZKxfcoy/QFwXlGDSiU8sIHPG
xbyMgqEg1i+Om7nhgqQsHln3bEzpslWNY4+Ut6bT5n+G5/zVgsFDIKBNdOtt1iuw
Qf1Ez9ZIWDHSesWuJ+URd+MVBZQ47c2+fWL1gHXh/4icpp5IdJJE5iIg5T/jRqFw
4Msmxf4SC4p9HwbozH0veB17pgtJwoRL/54lj/ZUNURl8IbfO7DJ7zeehXMGJn9u
l8K3eEo9rUdjJNr+pE6X27+Ena19DKOu1qV2qfPGGrqOUdi5iAOS7wex8ZXs6PwX
XIiAPPgdU+ecMweaQihrE8twb45eDbG+pUduziu7fZrvX/jheIxBSMc9ZuVXlCei
QXlJ8dWhrUvdOW3AVc8t2CmUg3O9+89wjHLS+HFUpv1D43oBt3ItrfpH1UWOzMD6
90UAuVvKeLiGwzVdo3ecYOnk2H6lqbAQqjF4owRG5aTQ0940jAOlLfT85CcO1prS
vmfhmoc+pvadAgdwwWfwwg5ENBVVMXo9ZGsvKKVTCkWw5i211ObbFZZMYdDNDAz3
u6yySgp3ExhXfgOBTTtqRebzYaefHI7ydOo9YXb1uW0bLwkqxZWRCr7pckQK1K8N
1yoDj81RW9Knw34J9YLIiNbYiNqMOzz/DmBIBnFHvcKWxg+rk2ezgUL/ZAiE3uHh
d+O6qoJqIXMmSHY3salG0V3Ojtan5q42QN0FcxZdYVtaqimcGFdGGlGmaFzVkxmo
L52kjLVzM72dtFOYT6fNzV2JmZ8ZVjrNfyI1wMdEP/F/fG0sky2q53M9jSjJAjMb
ywe+C5Ud258eNR77+GM06TifgisMW0+FXoAjAZMIF+QrpuhgGnC2E3tdariuGCtX
vCxHhILh2lJc58/eBQH8BRbUgXP3rVP+N4dCgunbjsrcePQQJgYEwHj18Hj+zxaI
1sgZ+2zw+xPyl9KneFyGw/v3cNpHTg583q2zXw0UT+R49cviunoKh/RCiwPfiFwa
SxOQzKzk93CKgNUwWnAa6AhoJAgc2TrN35F1SfaJni6khXbsmliXzkPEioUYRDUZ
APiTpc+8reB2tpFMKzcO1i9WW15oUVfLFLWFZzMR4BFcvgYKtNPOnf5cqNnJYHDB
dtpj0WcfKYld1PwNyn6LNH5MKN2hAlgL1BhAYjQncy+IjRmA0Lk8TOpHgi1QKzGS
CPko8Wj6xASg/mnrZhcGrRLj61erTThgjsy2VgDrV1HdrmGhxxLqAowSkF9t+Q2F
lTVIoCzPQMXeY+6KeepvdAhD8WNrYCbf8wyd6iA6+Tf8cPcgEae2Nydh9NYAoRAG
I59ghfdFXHDKob3BKeT5OOEwowFVx9RGTRyuzKiGM/psVg7gQ3nHfJdQXVBIr5tM
l203Jlw1fewu72Q1C/5OrFnXgF41o/hbzV1zVvhxtL8mjGG55N6RNw+PLt5PRR2y
IFx9LMhRDtoJZuJ1MHjEAm0XZygjYuBblS61hqofigPBzd0G4WKWYqB46qxyu60l
l2I1Sq9wyN+xcbuLEyCT8gXfa+51ZTMBzvvPB+h3a9g4PniRiFKcpPdTUvP0JJYA
yaTgekVR03HvJ8d3XFGaT/SpPUO4jgofgDPX4PAEs10OK+iRUY95ZxKP+MjFU2yX
HDKUYgosxiAK2XE9pAvLXPSZ4HliB0N+mbAMUYB14C5HxDW6iDQDygABvrkwrnaO
J6vL+oYC9HE8WovCVgfz6b+1kP7Y50mwsPd6t8VXAeZQCa41HRZVSeoZIS2P7wDr
HHzqrOrgyNh38Ghoi4XYPjkIeleoDfR10Yn9ySN2D/1+dNqr4A5zHlRfzKIhMokr
ooJATY3qyhbWD2ANelUKGN8cpv6KOwIecHcnhlw7hUNg/8yB3/4r3+Yq1fEDAme5
RELm2dqbmxxv4cF4tPvtaczuwX4WNQb4aYyYUqWyYWcRQ7oBdUTbUGjNtBDBBdRx
/38Q08+EpNWOLD+3AKGNbMy+igcRuFRPXDK86OFoT2Hpk6bU4W7yEMFDAwyyXAZ2
FpEllEfdZGEyGAkS2qTGGzPnWM54GyTMNlRhnjSSflHkqX+MUNyDVoQYes1FINRE
sE2xZO6WM/ZmHJpkdp42ONvoupGx0MHGPmRi0/1s8y0poagiomLQCgUxVuTi3iMK
EEsn3C0ewIvJy+d9p8N4TbucrJrZCFJQBixKqvZqXqhuZLX9//FpnHDCEIajdVBL
/mhmN3sq/+85JndyZTT3RnwgrjpCwRPG0W/m4Grbtr5HqyMe+LbctfbxgCI4psHP
XkyAYbp+fuEoC5Ch0mSfzJcgKOs4n8fkX993mtOGsdfJ+/fbeYU0okTniD+av/VJ
GFbuiJf2wldfo9lXdBbpu5FLDYuw49Iu9fUc1KCuutb+89y9fge//6EH+/sXrW+D
3f5HEFGebDc7PH6huVb8F2JVXPgR1Frnrg7zZqb9iXt5hPv7RoOH9652956HVVAb
v/HDaH0bMFhpB+i2VtCzv1LIS2EyWEq+zp6RzNOK/ggUxHj1cOjOxspEuNux1seC
NWZhEy0IzX8L2TY2UT/P+Tko1m9DUgiMkNVrpgyn7B8Y1CG/8CBmQFv877I2MQx5
ULErDCbtPz6oGFWHsrUJi05SEfAFaMVq9rlraiS9C83Nqi7Q4i82S+DgUNky+4mL
YvwvtxviveiJ+5MUr5WHMmS5owQIAQgXapuYO4qwcvJ7sic5lmSQqCzdRrzxdwqM
ZGiVCislOZjaaM5KLjOjcHSZjaMqzIdd/hw76F0Ngo/zUEv2En9BIp2+g1wJr9vo
Jq1Kcmi5/xQGRS3J9voTDnUkP/VyQUCnX9goXFtLotl/geabHHlaP82O523Z0dV6
UnqSc5FM0Ej9hC30BIi0D52bROnsxgv5kAXFOcBxPt6RaS/jBBNl+acUIXTsMaKR
2Y1ZFe+yiJxQ44t0pCVw9vIW2utI0S4JDgI4mS6dxcgH9kXo7mEAt1PsZo9P5QwZ
SlaBfbbAZxbjRZn3Sji+QYXy0HgalYe6kGismwjQu3lDxIls7IeMx4qI1L3C7HnS
tIl2FRKzilM1AhQU0aWa5KuAtKvdUH+rCEyKgj3vRERQOrtiUzT5dyDrOLArD8d8
lt99uef0G0KvvIBZPU5Slc1UDezr5XVM3R08EngZlEhbYTw8k39IxeNx5aRNJwrC
fNoDTGH/7S94cZpgBtdqBRKO+bGCMnrGLOldkhc7gdmR7vkoGA3OvqRZarMi0bAs
mg0ptbFgGirYTFv3qNX8swMdCwJezwox08ITkXX1f1WRZ7r2+YGgktjFK/ksWV4b
VdMU1zygV7iVTF2gIyJ7s/+2W+him8iwAR9eQVUfnVYl46HALplp+0/n1sxC44oG
3DzJd6ufRkxYK+fL4+ubD7paAvNrP9b1jv2T4MXNeNs1NO3ZDU3OjiVee4dA28W7
wsjYtuzUN8denap6kT03UoNvgUYJJcJ5m5n1pr9f2pY9XcCkWV7JLxgIR1UwH4CW
f6a0DmnPmfMQIhGeFna1fFGIaWoc730XN9jIvogkZvAoZ6cdVGOdV407o1uJ+x5i
c+y1y54s/0HMtErCvrzzRYU+UF/BNMSTXPerAHFWFzEP+LiYgssXHEwtmZiVZtCV
O1vegQTDozoCJhURPtYdj/bVGgelT6hmbE8v4zVpG4hoo8JxBO5bPr2B5stY1LHb
KxBg91NfLNObupgFDnfdkhGFDDtKO5cZkalStglaxEFUCRHK6sW3szAfGoiON1lK
Lp7YT/JMU3md9HJ2leWQUJkEViRNctEE3qWt8tYQpOdnneJKX9xeWaAZeDvaDNmM
tlT2Q0lcY+PdhY92kN/U9hMQA44j1bDmwy2lJnr+W/Gx0/NAyYGORoYs4669Hnx6
sGmwWA8GBk/kb25lWgWfYE0/s4tLoKn0E9MvI6LnfbVIiYLk0+5smPsZfjKznIMM
pNkImNFqwfwSUHP/HnzCzvObybjVCZxdGOFlY18JfN61PDeD7uihPFKSJm5gYD2h
74dskmQaIwAp71MGTX61mqiYl/4y6+Jac2dcS6S+zdY3TWUQkB/AB7vGUxL3NcEm
ESakz5uyrzwuykPLavH2/QHgjt+uk2UrdqS44EgU8eR6d4B3Svr8qecD4ESLNRVT
nm97ioovcuURu4DtdsenNUzocc9wkPbNvyvHcG0ols86/+xpwCVTk6x41Jxk52fQ
BDaSQgwyk2iP2u54kJ/SfEL8q2BXY7f5ORK7eNnXlg+SDF+92pXJIljPmVrZ44c0
Fakiusu1mKxdjs+bs5ZGDdVrg7aOt/FlBNgWxFhRqHv/P+0g0ET3KtjbVQBW5544
3cgEyFxmLNKUcUhEI9tHEF2Dqts2zodtthUtCArAa+yXNhEVupoIxVGs850g+XVM
xo7iob1iKirZuPUOQtiyRt/FWarhxsEY7et7lcpmnfmjZ0TphZlmisNWsBWMin/V
z+4WK2gZieemWgV7k6eSPTaDtnP/7mq2reVgVZbGhThEBaoD+mTy3osgfX9sht6H
N4xawZdwPKrznC/8G8m6v1svxzj/n/JwLNv4mOZQ7udfl3ERNLB28zv16swE7eoY
cqNKvg9HnJaMM5AvjVFTIOFUr1hrJD4EsurjegmpGKlHDizyrY3hHnHKCFmJM8hv
Ssbj/FIBMu7mPuDZA36ui3ArxBWRHWZdMBtAtuOjEe5/1fDD3vHYrWlhmx3syFb2
Ta+fQ8nNzfXd7uDCNEI7X7wDEHu/68GFyAM7znT+jZYJVmg8dMMTDp1Ov8GaXGdT
oPrmg8T7ekbvR9GBxawwEtqW5JYep/7rj3JMrsfEJl/3Oy6LB+DmupYymAm7tZ/t
AjBeLfupSwkkv1yzZ042uh1iemBS7CZft7Gvlu4hj7BFj6tWean7CEvhPWOoR03d
ivUjPCHf/imLjR2fipKED+MCkaSTXHJf2GOlYIM+Kn8imrXbIpoLiodhuKWHj5Ex
opyQov1PTJGnHuHeXrzqCPwhl5RcjVyWjqZZN0NQAT1G47mzn8DIgcDCAA1tGbb4
jA4nZSuAZ0Yx5TA/EfWAUXg1vi5tEHwKead+T/9b+rWeiDfwKCtPJHsa/nfMf8Wm
1OqX0POcEEzkFjPkB65ERDJpDHdzkjdHlgiEhOC3nun90dHabG4q2Q+9ixNbXOgm
QTtSEVfRbpslLyEzSvx18/C1cj0w2azQTWU8FOCHL4if2+j+PH/9s+VxxR3lu1Xw
yTk0YDe+/g+8VcDWgb2zkzdBRHOJ2vWbFXs1OJzRJ7aeH1p82QRIY4caQE4jYoBt
PWE2V2fV2hQGUQkWXgEoIb1Mapz2AuPb2Yq0KtrN59rg9aU2SdeXdm/6wK28j0eq
4/ivfpvepQOerz9DMEYwgpC/cWnb4tiNMJcn8wktL+hhZkVsuw519wMW4yS1L3yy
lQ3bcdbCs9lAkVgpc3LMldB3FFtIqI1i7SclyOreJLqPAe1Ov/2lQOjbLO1buCiT
8XnbP5IAftQGofox59TZXPxpUS488qoElfQLDuCkP6rcfvAtjMzd/TwmFJXopCPq
WDJWGv9KwbOeG+mw+HVn/rC+tVYZy2nzh9VTF3Rdb96LpCq1gSlnKLGfOAc98BhY
aigvn8AFyNhpUkIPrXYgkrDoeVTgE+tKK0RMbKB3Twm8iUIkLaIbYkCp0AsS3Czt
jbVov4v82a0vzg/egA9o7l+DQeptaIAaDBOESOfOnNQjeE6oAjrU+EnxJNHA2nzy
ySEY6dxWa7FWMhStnGHSG1dAFeR6+fcCqLp/ZB+s+/ikvDYGpfPLjSdmLDLs8Jm9
rlzpTQu+IFkSUCBJ3TwhlbJTpf9cXopZrdLnBhMbrBlPQL6FrNbsRmPlh3CdVGU8
4FAlOMUHGZw90N+qpw6TqcUTcIGj8FX/a/XCOB5OxgSxpPF8ObIIEZSoAKx8fgsH
xzXwDegm3ihfjun0yN0i/j55h0TpxrC60Gyy9qUVVRORXCH+TjupnZN3E8291U3P
AVMsdtj5c/aEKrsMRFPy+Y90ZA7+HvufBatSWWJRcwVZ6LtrB4fN9QG2Oe21bige
CRZQDaDXziTBZTFl32Y24oZ9sj9jkokm0gsE9HrS2zbrPdRGMk0FwwjkxWIRs4ze
XoYL34cT39qoo58kRrY++2Hc4JeiJMZia0yAEXzjxqshlTBMYK+9DKsMj6gRgMqD
v3vFY1MVioWxGnUTi3/zM6E0AL+jaNs/0XkIc+YD+8/v2xXY9ooYtLTYMHwPriR1
NLw+C49UsXqlbxM4cOL8oBLSSLJP8cNw17JiuDMvtfPl59lBLS6k9coADtSBtZVy
I+2BhwuCFOXx6oP/JUR2ijBjo2PnkONlhozi/lZLjhWEo4LHOKqI4cvMLLRfi1LC
uzYU2Dpzeo8U1esQ4CS7F9e2bRVuGJAFldjUFgapLnq5igaGOk39PvKxdsgODPVy
JnTZOcaCwVAbIQNQsL6FLLiHhmOmDwNmjUmdU697qtMNCTVekEk3rVSHm+JJ8kRR
CWjwu8izNGUfSVTjPd0acCrZpehEsPLrIemKHZrHy3AyBaAQy+4B7ae4Qf1EideI
jHUqQ3uLTK2IYLKACRPjWpjvseEoKkdiPCz51NAaEGfrNIUe8zhyTVnndWbJvhh6
8cKvlXFflyqdLf1+mInEdoFtyanY2sKr6uD+iUmBBwVmevVXYEX1XC9nzK28xH8+
hNV4y5ZyoMjvZ2CiDixFDvVhiW41Oku6C7cXXYqHdRLadhWQYihKejZdwVW+ullL
dc0LgyXfKTk0ISCq7MmbBfcSqUPToYeAQnilkxodLj1HNkOFePshFyo85kie9HuH
HraGfS7vDr6L+AnabCD12dztmzaeReJC6vIugKnNCLlKN4BMAnEc0z2npzmZh4X5
TJuqly1FIocfZJtZ0EaECqHGr1GqJzmPsoTV+IgE+ackYbpS/JRhjA3+VORIVlGX
bklsr7P1zgwk6WJFkOPt/79sTXqmQrWMIycAmCdG+nKkdC0F2LkorBBW3UVwyHmW
B0c7B5qyMxOebd1NbezzQMCtSkp65Rtg53nKDC0qXjl2BZEQRWzUUvGxDNfOWpwB
mPtwAhV//cRmYrt1PA29Jl8QHEHvd20VgfLQTdJCykJCaLPWbIJZZPCASNcAgg45
HPAlIOSgvvLp/7xchD1baOvEMk0DzyMePY5llPPm9GqiIt5fXs3Z49vfVbez1mCw
7BtxP4Xw3mF4iSLQTcOGUScdWidiDQR+P8LwVe4u73Q3UX+eTXhFmD3aWQaXQDWg
UvkP3pisXxntta9vBviAEYv6O9+/9FODxL6Zi8FVpoC3BFvG0F/+xWdl3iNXmuww
5hOTH+GJN+9FIZjL8WLpyctYrqJdqg36A9cvAwRkhJYTx6PN2Stxv9x9T/RydB1s
xbNVvrx2Hk7LbYQ1MNHBlTf2nAi2ScWKB/q6Kb2huWOQbQSPQEEYU+MOIEvQBUpD
fokj8yGR0e9nxSP47Mtx0y5PD0uKaRHe49e2rz3u5OwX7MzezA7Ho7zoorgmpKde
SKxcNu0J5U2oCeHnYgoSmwxu8wU3ZWia7OpzeietB+G0rk/kUpIs0mzadQX2N8u3
wT2Tep2JvippgGhL17XDVp2axBIlxc8Vp1DFcoYXVUQumKm2p+6nGjr3pgpXKvDB
n+yf1HLLrHWrUzlQ4dKWKArD3fPIleM/w8z2huIYSJTrVPGVlbwfMxZjHMCRLpZh
OtVCws2zSf/JOSfgTrR7Un86RvpaJDoZo1laRCEDqAS5w9r5giD2iG8s6csuPqku
pyX+rN5zdQBJ5HFr2Bw2NkCtTXy3tSjK500yOt42qt+hVZy7ktJja7fkYe/x8vIz
aRNo3M9qiITCp5ZlA0qcZZC7ZMr9mo3QMeNhO8cd6xtQgjPAfPTvCKrsp54U1PLX
mjJpIdbw4ti1IfzDFNK6cpI382C7ko4xxnzIybivcqJDGHpo1DyM0KVvEV5nPnRt
VE58XOzRzCcITXuMAX1+DQLrONGNg8aoYNplViwMqmdspx4KsOuVycOAmeNq9yNy
U0mWzR0PMeEswphR3YpbC1RXFs55ggAofoIi2BmFThAIhbrgZshmhfU923xieRpC
G8iR1K68zvy5KP1rvytA+/fGlDYFU7rDz1YTXsbWqH6Zxua05ePkZocgBxXmKXwQ
rQGeJaQb5odrckzfz3NpMAWyS3m1soKPLE4OSfx07N7CyDY10mwZLznA0c5vSJb7
Nod6EBIB+XWKZZ0ysdH/lPCx5RjXF3F0HicsGMChd6ATafJQftq6t76U2Ki4m/1d
6sZvobVPJlMjiyepDRZq/d2Tssdzbqrb4/3BFseEkU0CZs9S2r/ircqAE09lCTFl
LdcCWan9yfZdZWFtA+v9EUCCpOT9x2x0bKh/lywb5mS3GAIKIrLCPrW4/GmBlSXi
HZvCbT9AmMg6kRKBhL7vO72oeci1a76gXsTsud2A3B2pXJ6E1ZlS46dFbgy2XF9Q
pqxErqGfDR5+BekFgQtWG12BA1LxysyYBzjma1SY/7TuNaWSbVafJpJv5A194ghM
GGRGfdnuRptkI+i3Fj/A7/mCu4TFWiKthmBI9YUUbr4YIl7keKUgt4cFU26CS9w/
MmNPulfTEwjwjEGqSQMSNDWofu2cZOvJUKzVjCzpn8ySTNQauBsI8I/nhHvrp6Qy
L5Mww13qQhJEK01sm22tZ6etlDNlcU0wsse9BQ9TYrMFKCh0/S/kCbtPvX8QSr7V
tdksXGZUMEDbEPpqeSwxRNonNrlDY79oPnL65ay9q5fcVR5OylV6yZLCAxXk3REV
Tz8/CNHEGbaAA/gr+LAWUF3KLjFK0JA+ikFZ5BMj5prYB8C1Kb62CjK0v76266hk
FlFYe3mSm+1hh8xba34XEY5FDQSrhu1bE0nTHjyGRRzTS5a37obNqIPMr3Sm/old
Di+0AscFkwGB6IvwoCglndoUQtY/ClSdxttnTbPurkglkwV5CcQFYH8wrx6d8RQg
V0O9LCuACvKxk3J8oJPbL0KivAXpOuRBal4WWs/AY0ZezNSuftYBUA93nJdlKyqU
j4FT8KY0J9dGA5hGYRkcCP3Np8WbSisAqNBLkeQArykfwgKDmaKCNp/Jc9w+HfcH
Hg3My5O7tnLNl1wiWQXvtY5llEGNCT4iLoxZsi9648ShhvMXFRurr6fHjn1SAK2j
SOa3nK/T3sTEvBzpB108GY54JmFRIEgPQsxseObOiSYoNU4rf0h+9svDoXl8haAx
pVXY6C12eWcpprmuWksvpTEiqPINECQ/P6x5ps01u2Z0yMz59rmdra+NpSeVd6ex
oOjsU+8eI93ZehzxE+8WrNGnRceoRdJgNTaYzigKz/EJVsxd2XUtkhQ0AyM2zEBO
krWWQHoSX1LWHgCqbQ3xsm+XJgq1uzTgiwMuyj+PWwMPn9L27ArF8Ua8q5XrlQ7+
m/5eketFCAsScN6mM6V/a6K59XlKNPmC69bm2EcexVJF+fAlx0gAYoOVsMkafq6j
corL35op6NoWIxgJvehRZM9bJqTQf5LUjXpCIneMMSLHRjf+bTip2eVBCCTOoUBP
GxPzrSO3NbmCsEYbwxAFPXIpjGxenE1hpXs2CJ8ZN9ipuIk+I3/KOa4CqwBjuBUb
bF2v6MUhp+wHQeU9dQvE7ZtpWe4OulNB46dVwE8HSQMXS/rvDrhvvaNnqA0VD1VY
hW3IRJce+OELRaV/pPIKMTiIBEKq8pFlZZM2QkXgfmmc/V/MG+Jl2aMDwlOTT26O
32U7R6ifpGGzuj7YsEQwaZYhuzOpFMn9RT2ff3lElAhd2eCsi3L829TWDGwOcZJ2
8B1lWGmA2L7QCvUtYnLBZVhE9za7dLH5mZG+9KuXzda5aICkq+WE0NkjtvfPHjVX
o/jWbT+gZj1Kxk1n415jo1edYViLyrhbIy879KYGcLqgqMgeR6J5Z2BUkJDyrDDf
7gL/or7p4CLtkwvdh5RMDbglQvlZRujsgzYFll8VYgiqJl9LE9sJ4S41HzEyd/9Q
BrfBM3KRRpfthaPfiOz7w4+SdGUjQB3TQHe08G77uEbsAyDaPbrv/Mt7aINweDIt
fxNSG4j2R0sxfIsiwjjFUK4S2hlDHoMTwBM80FPNKBBltpUq1xARscCmFkdlH/QH
CR8nHdLljvShM0XyN6dQ4wLKLkCCP9Lc4L4Q+smnieSmcOZtrpJm25CDa9Ae5N0N
SJblJ3xrYB8u0dysNfZZV1uJof9oLzfAWvfQwfUGhbBMGprV4zGR4pzqnuVtuFIi
LSx42XUjH6xf9nOhqYz0v+XOfv/ln+e/0y2NDfS5zrMbiDNEXOccu/GPsUOMk0Bw
dGR+44L55TB0GMaJF9MHMFdI2C/cUp16Dht8p9JVgd9kYpgmYn44O+UZBuA2bPq9
PWZhQfTRr1xDUlr/fmdXPvsPS+0antcQUiwGygdtIKWYWEOk1K0F3sC3kUZZu4Dt
6TX/rdUxdpEVBkKJxJON5dHxkuuBgfgRfBGjEhHm6R/JzwmMfo8PTlL5ah4GPcWY
7h4YcE2XGvsV4UgmxW4HaidnBlL24CaFwb6KXmeNvOTBAHHJujxMzEc72xjtECao
K4CIDIBUTQqGGxZpASgLsDSrQZVp1ZU4nTUSWm19v1DEsjT2xWv7FmT8WRWFZh/o
nsmY7HKi6AR4CbUbtK0ikSnURVcFGuiHiiOGoqPgKPzQVw36497yjOdGG0w3oJjW
X/RnSBb+iB/VlkJNqr1Mt542p7cxJgNnOiJF+jlJbSUY9yLsOKbGhn7AB9CjFYj3
kj61HKJq0/Om1v8eLhueGaBbz9dDfbwY3ITlhU88B2Dr23yvG6XCmRhy689c2BAQ
GWKjpIp98uPYxrCDKAE2KxwdJBzgoqXwdHpARJw7H19Ru7g1oZbE1J2whAtK+RKs
JCA4rfYOFQR5pk9beQTwFVrtOL9uZjvGFqQ5+fdX37T/25i0DthmXh5uVwJYvjl0
0BxK1uBFL9QfSrDxNv+ociATQL75QWArNb7PMyOjdzfhBYYelkOVAAigP8nJEmW+
dt28+Dq+brZL5qwcMEaeBjsxJcqMRm5ebjd1XinnCqybOtxdczhh/+jSrjwuba66
jBbXUxl56vgdM9axj0wQ9J7S5WEK0Jy0CQI83DQ7I0Sy1Iv5TtVHNtoz89B+Q6XU
xFsn3dfblfNN5LGuIUh82QA42smO7lyXxgy5xyg7EW9xVeC25Q8hBFfab4Mrkz0z
Yy1K16dvdv33v7CT7pYoEYIMfZTHWcCAvRk5/AqZrG4M3JhJmmBom/4IjH7xZ0eG
NtTQRed+dMwJEVB98EyEjsM+/THIFDEe8nv9d0XESvaaggvODqt0FO7l6xjthrRb
M+xNJCjdd2GQC7hZZxcBBHBDfxqtzjhX9rgNiHVhpwuYGxDyS92pwO+YYFcuhqID
OMuwHODbwtAUJAIFMDsnUCh3YCKK6fPbBJuUwH20MeNWtlM8ekkAA34KMmp1MNrS
mooPQnr7HP7YZZVNmN6K7k9W215dUpXYb5GHJ5zN95TYq9uvGdhFpAKkOkk7CTNj
HXpyvbJHaIXoXrwEYzJ/O5JIt/X0ISnDwWJB+eQA55LSkwoEuIEEFNkNlskuBV04
KqPAbv1wCeOF7W6OdpbUqyPiErH3gFGOjsQxkF5YvsUViL0vYnldXzTgegbiKmkH
LVIHmLEOeklt9qYDqUJtOQwWMkKjW9/lC5ESASohG/ge/mzMTBw0Pi47E9whu4Uo
12TSCcpcUOSn8JWnHSXOZIu7ykBcVS5zit415TqBi6ybmfwCneRrxmzgnqpCUxZR
lIwwIzx4I7JEoZCG/FxTgCcQm0yZ/EgWhtplnYQ6aqLmc4hZk7msvQGjcsPWV0yg
MBarQoCPXcZXzjcn1ESFRf9K7ickMhOZdjYoZn7UEypf7CftwPCbGm0Nz9Ii38Co
YILnWpQD0umcipfpofEhjCacUh3r9F71IRnTbev4I/29y7++wZzPBqiOtQA6ocni
PjdHwbNSQM1WaIjt/i1r3How6HpVez8YSJFJ3H/zUvWGq676QFuYXb3ADXEKWoi4
MYIIAYf7a2cA4OUz6CWPoKgCwvJGHLR/1kBA9EgpSDR8/VqVbLPYjg8FmBoPNo9/
mB7vOKZDQir9wteZeODOmgvJrCIoQ8yqJnzWHqQJ9uHi32Bf8uId0pwlBRJaWGUp
0DvpJY3VFSdVBX+ocLtidSEhnsujIAkKlg1RZ57vL6MKiDpudKvsp4iotQ19zdau
WETUv9Eu/9/Ea1tsx0CpoWUScJYb1pWZvKns2m2jCaPO+TrXHK5qC98D8hTLUjvM
QSx6ZoDRRj36OMUnFDuI/aKyBPnQRHE80mC2zp13xGbj0Z0tI6Tb2mj4YJVHm8p6
+80h5tPOGeQUDqzi+npPOsimauAr+jSnQTl+pgTjEJqUvSwXvEKtsrEJ6WTORzsX
cQB79RQxOPh02MWaOJitPxAy0r+H2PxIY8T5c32c40cDUz6F0xS0FARTO8HIRaCU
PnhL0HJWBNaB4WbmKZS8HOpqG7qseG/ReqWxzkEkTStSol0aEfuQBoY478bzEVDR
8UOiw9miovN06gPB23lEtrwO0EaZXucTVQwhK+D9OY+XEoAORX1N/+vatXP3AIhD
AH+RspwglUpBvlmW2oImCOFgS8cnp9HthAibQC4Vrr5T2JBYIy2YRbtfuC3OvPLT
WdEzgTtghrwXSgpdpoYnasuEScGaT66dyvz/4d121/AvMVG14l8f+wGIhx6zYSR3
fppseskfCfvZ49SLwnSuEjd8re7rOP582AaIQ2EuqgwfsFl6oCSsQY2LmRIHgA47
2fd45YcaTXoOFOv4u7Apv5GNYaDd7FAZvx3oxdzWDFCJr7IWbpJiOuBZvS8pxYky
1SOHh7LEi0JRH59yWRpoPUGyCXeuF0/IBDrkn7XMB6IQZ+fg/V+nDDV+Fcb0Hweg
8Lml30WBsO25/9N8WDejljYzHpT9VT5yCCUDK5lZLx4bMjuDdqbH/1IpJ42afFq/
5P8sTfTrIOJZoVnJAaGNzf7G0M3iV+2GnHrcTtyAvJaIBEaWiVvjmLTogZ020PkB
Nvfjw3lttPDzTAFhggnhEXbh6P28du9L2ZkMlf+9sros+E1rzUp1ACZiuFqNeBXH
Ywn2IRqWDoP/fhhf+RUbS3k6+lMREJEiPVJC5Ndm+Qtgfz3aycuJbkHbdWQYXKs4
9OOd/hdAmyEANIwNXSjXAo39+ja4zVUKwNDELvNPRM1m66yWqi3XdcW8nx5qDGaM
+wEFE2IUC4JQHhL/bS23zOvEsBXHSXVfU8wixZUorFVcehXeyA8YDNbR/UvBQqa4
OWDQ2/g3Cygd1TxFZRbORS63CGXwuXFACB8KBBCnGvsD2JAxLq0btBZ4tYySz0JG
XheS8KIR/2uFa/NqXVURfPnpKZmOD1gc2w0LwTriBVfkDbBp5kaqXYMPoJ2zQDgI
U+9umm2OD3X62L3QiO3ULB1T2IkWRKHYfdtEhGo7TbLbyySLyOS1NncjP8Es2V9U
tNn9xMOzhWNgB751SVvEqDRoDQLKgq2goDavK4D31jfZLJ6AnLuRm7AJ6h/ck8MT
aJGUPtsznW/ksmbMVPh7X9FYvAgouvM6x0wgK2FuJmhLInrVKks026tyCFI0Xgzu
xIbRf7qx6qeHtNLCuMQMNxG7M+t2NYTkQds/WGqLEllVWapo831fl0DOCAVd/Osc
WYDX4iNbjLu+AxOucF4eGe8s6fc47PUqc3GIXobQVKXZDe9Qc7zjzksV+1Ve4J/D
H+VZKtZQg4vliJnUwjR4ANLfnonHzETeJ+eXd30MEL3sXkAJxzo0A8lJ5844hTPn
i8O6DtzyFG/eA2tM6y16PKdGBpU1ROZYX4k2p6f2FNBVPhaJ1Z97PyAYbO4Vs/Nr
pqw7P0Tqkwsxns7WyYcr5nwd/BEeYTjaiWtvt6byDVriLulVGh3dQ/eTYhmi+vm5
yedmZBADCEwWkjZ/8ZMGZluqvOocwUCV2w4K3ZEJLpdCMd89mcRr4eHMpMp+Pmlz
DLKc54DzM1CIHdWJK41wUauJ/DAx2LhkzesG+JjpZIJiIvNzcHvv0iB0vBocuRmy
S5bWNELRFEYhNLE/htt1B6nTtM2xmon0Bly+baYzrNRBvDw/+afFSJW+8a+JqCH7
C222bUIhkPbnWOfLdBaFoQELx3F0EzYMu93uikIivAJN8NtglOiokNQd4DX7Wuk+
WOOUEq2olYG3lpNCiCaksYmV8d3U1azokO6EW6G44cKmAH/nXmIcYdsFwg3aJYj+
8bEWPk4LEjvSXLJOhUc+eurfMSqKU91I0oOv+VSs6xrm9WGswvd7AxvdOd5MeAmW
5Lxtp32hGekW5nvabHl/jvB9DgoXMzTkm4wgsTzspXx+L5mEGFP7cwlVzwwRtJ08
cus1HQayJtJuSbjf7KjVdkYkm1c6wB+fw63DPDnOEFceP3++OluEKe0OpqrKVgTD
ImZU9eDUvVb0k7sTBCbAYUMeo6m8NAffK+ny39TceFHzICPs1/zOReh1HeIqa+UO
jxgEWPCaXzgZ43jSZa+vyCNdXfzETMyTNBQdosASh/JVq1NcFIZxjfwXMDsjyGKY
yy2O5ctAjr950jexJ9TfOPn4Yk23C+AubwSWy7SWY3PQykOVi3FUEgJdmRHd/WN7
sYi//beJVrW2FFutzbWoLhSnkYkhqCXMX8fbNO/aiIji1oq9C6fW9iCUKeDecS9E
xpTVo3jXQGSbR1WJeHK1PCSto3iSLU4K/jKCJ6ToZVvCzkvieR4cHhXHIPkNUVx0
VShw0RBQH+uHSRr1X4+FTmdsMP3BzB4mb6/hMyv5qsk0WQVl6ZyabJEYwqbTVMM1
fMtxFwuHs/pkGf9k9atbw25MhTxmn0zJsieVpWabjIgq5okNI9tGcQKnjDz1KR2u
T7kZSLQ5TZ7KxzMSvfPTJmQpX0GKSu3JS4TFVIVdj9KG6xWqi/s0YlgGnG/DpPwS
sPP/nZNMBKJpCB3pAr/9xEmySTSfVyhDSJkVHwNx/Fmtx4BX4DgLbjkkRBHiiiS5
jvkyGe30RE9albqe+nzrhHNnuRTtjKm8qv1U3bIzKLyYtJod2CrUuuxBBRv6AYUh
AICDetVZPmbsUHU6axxMjqYQR7mPROILSLFS+Fgn0DweEraP6pi3JbPriNsM3mhO
4kQT5ZeWiytEs3nFBZ21wlO1shzgH5r7u8eTjfLXZmxgMI/RdxhEO9GIenrHJQuJ
zU1U1VskQE3321zc16j7uYtsrP/y7nNmH8d7t/YMj9OUjKwXk+GDBNfu5vFPQ7tM
saYIPCjY86oD7g33xirm2TRqR/0+srlCefSya3QtFoXSOTLyAtBk55Tk30drzZ7b
oBsLrvV9rCIURjBmj6wj2AudUGVvPFeRuehLZkTQObNqomtcc/JlyDuzHbERLRLV
NtpNzOz0rH0cENpuIySsQcUjZ0whhwIRNkhi41uWwgFM8JIG7ix90FIXvomqZJoq
1IR2KLuZPvIrM8WQ9jOAVjCZzZm7dR9Vr/CAXpC4WUh2ImCHCeUta2Pl/E8uqSCY
lyxxV/+A/ZgKQkfXEeA11jCIulvWtrzavKYOWKTr8+k358nljm2D+nBoOlx8/QvN
pbSbxqr9Dga7kjwS78ESjUWGUlw37DxgHdLNZMflg2De872KlH4RgHn0A9WcsZWg
y1fNI3oVkroMTtYzbK3sszIqlhE7nd8GNL2CG7RSNG9TUi8hJAmuci0HOYs4t1a4
40Q5+BUGYjzI8DrEK1ugD+9sxKj7KS3rYaA84XKac1WBc7fVxQwyHijX2rewEt3T
GGj9CTDLTWCewEu5uCLezOVY88kbJ1qi41JZSIC14MPtK7SvAeN4UYbwbPx5HUjw
ghIlP1mFgvBT9dqe1vFL9/IjcOfwhYwIIZgMqseXhvPNzGBw7Qc2nH9QS9mRlV8S
UvL1+WT7YL9pAG6zsvemmF9xfJwE74RB8XeoONmj8/Iyp6iJXKH6LM9+Sve2y2NZ
1FZdYyKtdL66qMbjc4Wo6sJP3JhFyv8CPlIaVbEJlq95+4ucPJl9KzSL8kQxo0vc
ijEmFxmrMpR5ydV6krDPXhgBH2n6hrFv1wkwvqDEUsC8D5cfEn6xPUfJDYvnNGo6
eAnxWY90EPrQ5ck1X0lIfaiaNWpkGqthrO248Af4h430tHgGIDbZ7p6cGFFxFqav
p0CcSdC7L0hqOlmRYqEbUfD39weTgcnLh8Ou3QsChGBfJSu+BHBJcru51bZ7ya6s
DWqlALmBy54dPgH6BKmsm6iuBEy+earRDZiuB1GfAC8u0PRmELcwSPyJdx/oEkAz
ENU0qPmolEHiAhYQ318qDuIvohCetNiYAYpBXffp8WSJVSjamr2zSBxe1yvH82n0
3OpqPN+ZH85Y4B9jE0NsdNhu8lBXVkJ7YYxzgGQ0TpQjeFw7H9q4Pf8HLKeMwmK7
yMeEVoQuvu+MAk3g0WafcZferFc5a0//nlPFlwtTzBQvZ0gRST/96oZs4KoUb7e8
/8MEAOn2mBzkHyvhzK5etPJdvzCeNMsfGNhWrwSzyn3dlX8ZCf1hr/1CwhgVkZmR
uS885kxjxFDUxc9QYfPLMH8eaAPGXa0IPCTi/XDkej4GHcz60gYPB3u2IcxWvKuQ
0yBqEvB5ZVKvZ4AIaSmHvezEJ/BKBdmJ/XHZ3fhB0ex+T1QR4ymYjuVVKP4XN8ZK
LyzSSLu0SPHCvu+ydSuk7wdGxWDmypW58RwXcz+JrK4U4kiaD5EBEwIgtor2NnWG
jytlJIec2MQ8j8PhJpTd4OLGFb5YCgcD0qnmzFC448mm9Yrd9lsB9ZGjiQnAGsAF
b0kNN5Mpt58HAhgnPJEy2iT28D0evgMFlpWjPrJki2G4eTTh6Knvkrd2LTQZxjbB
qqjbbBK3xNe5LbWYyApZgUtIWq4IoW0AxgMDpdgeiTuz7Y5sqSM3XphwQLjGWRSr
nL4unptZ5y4DKH30RvNJd23jv/dzG9i+GQnJDWL57wnsYXgawvJYgVYd8UM0LtWv
ex8lCMfLTDTNfCcwk8uoC05rkkMRIfq5rqWeXduJWoakB7q+B4K0Ix6ofgjpJL1Y
DGa61w+3CW4fcvR2+mhIIE5KfFkobS1VJVEMpuDQcIGboqi91lD9NbAR8LgAgeee
9BHRptoK18sFZDrRNsX4xzV/ifsICtNdRzY1wEdq6vBH9Ytf7ZQhfOvh3W9X4Hbh
9wWRrtDlbb9Y+jhnNt3Hkp9tN21pxsB1VsMM6hVfIgqjogWIls5DPa/DkdrYFdn4
bJtkWck/RTq8UcIl0cC8lB6Zfg+LeSXDygoJq76FFclEcb722UTQVedb5IwMiTku
aGDCvNFYgvQw2FON2mgw9Mx4WM7864Fv/WPjuPGnzP3Koq2wJjZce/dzxY4LUctt
4T78JapTNoDIKJ4XOX4cF7hWlWNtL3jy7FB+2t+cPTLWu2lfN8tIl7Mw6nxveVN9
8DU3eyANv9J1dY7Hx28lq/CluMuHA9DNHuVB3B895PUVmsF/6f5GbIN4useNZNXX
9HoPyieGN7UvVKrGQs+E+Zm3NgEMSDJTWZxav8nB7j1BQpRnYKspehppovcU9q6v
mQvt6mbz5oULU+k7CmEYh0M8+6O4/ixT142UzvuN9JBxZKGds/rqfsy5sqJRt7Vs
xhOkp3X8Z3XLu2bSr5+WV0R+krgrO3ZQNMUkxOEwQLRIen/APmW3v2BwM72pK+Sa
Zkym25GLiHs1t4snnAy7+pT91ylfYRp9oIgt39gFMrmpNV9h+INHYQeUUltXmP3r
m5uHNdbvy48Xu92EzoNdtAeSDe02hwvBEhwSL6Om4Q71Ha0oN50w+ozBdSYo2H95
fg8ekoYVyfQ23N4z8mt85JTlRZDTUNYSwUdrQ857DeUUrPpFLx/B90XMygZYsJc1
iLae0gOZtiI+M9rxqv9BpzfQAjAyh61kF4mxbxCsyLgyplEB7x49yd4tyN57HggX
IFV/jPgWs9thrOLHITb1c2KULO6WLymNu28FIHXs0a9XfvxxFTTERdpuY2ql65i7
r6bB+Hnt2wpSGC+OvaZDqC3peiK2GmR9K64Y1Rwn+d1bnxQsstk+dB0IH0H/st7J
svZsuP94f39c/CgdGHWXtEjM5zouW4LCHF+sk/pLOH6t3XVnWywHTwgzAJEXFlZj
dR02bUH1e5btqDyx0w8sU3c6JhgddONzmFcKVunpfOnDlCxHdHDA1Twz+A3VwQqd
z7WF2FhlPyhHHuTm/9f3aX8yALyo5TV4dQZ4MJjzR/RkvoCAY0owd4BZ4FEesIh5
jUrGB0WGcHeHJx9uT2bEIBJvXXVyPSPHuXI91mjJZ6I/Vtd0eM9DTxFJ//aCaoGW
lK/cV8X6Wv2U3XxD54cmkne1KHmdEyiBG3L+JAdWbUxy/E3Q7FSb5sNXUTW/qK1m
D99Xu1CvFPivKUHrLEuvtLBAnWncfWM030FYPRbj4yfuRZz37vYGtvbdflziRzBD
wdx3EXM4hEZ+wpdVfadlTgvDW6F4s1YR8VVUfqf990COkFXLX+9tzsGaFfbZpKnv
kvJWU5N+0qmpnR7Dk5l6xY+6PD9m6qwiKBGjxEOmX3HOQucYhLyGb4uhXH/JL4O5
jwtBbVdz+AFel+Jo+j2ytpVygw4jTZ/a/rjdYeXTpMegWhP7qISmSrBzd7CXL7Nn
Fmi/H0FHmE2vN30FZCJ7yGv4qqOD+IK0nPBiJyxkbZbIGKNgv4tO8ySK/Sj9GSl+
+qrP+IPPNDS5ad96+BgXU4ofFPeSdrReoZezRtZpj4DkLbOlwSOL9earSAn50I6l
wctBfnqJdR7mDffISBvJtKFnaFRHNv1rwyzO2GzOM+qh5FTpzFkZPUm2FPSsKQsx
hCsxHoDIwLP5TucMAfFy8DH0Djn54Bt2Dqqr5StMmq+rV36YK5MZDAJq9G9RzHr4
19STGTlIz44B9qBErQgdQt+tYZjYrjbFAvQSIq/K7BL++589vM92BwqApKcl2lO7
Nn8JA5rPcLMYh4FPxZ95gWUfvrnQjddV3XeWMkC9VZPpnjZ40GKnZMUOzLYYIABk
5VG3qZmFh3p+U63ii8uX/BpMw9hwl6u39vhLlcWYc3YSTSs/VNpmYi0qYvG5lp4n
xh/y17U0SVyIpV2DMSU8Io72IaSv9khcySZ1h8Fk3JV779iMiQLykpfV9W0k5s4H
6VROpKD3siyVodygv3kzgWQrJHzPrVO8rBZp0nHU+qJKFmvn8TecikBjDrwkmVFf
8Lqb85SG8NywSXDrbLG9wa6pHZ3jNKCczhzLE4lUIZSd/23l/4/axiucuvrXs5ie
1lFPURpiF8fQcygYkQ45B6gb9DSK0XAIaSyMVp0H491TXO1f1OhArJS9dvBRAaFl
T0XuXBQcOgBKrgAWoxb1GYtkJvuEQQQa7b+rrMmft3NnUOeMDgIS/6taDRAiPVGi
8qE+zF6fuAWoRPPL783Fw3zj2VJvc1Jx6VMe+DOWuTDjlPAYXuQPdX6WK3soIXlh
Yz080MrYRwSs379sKd5rUoM6tPfazRYIRyoh6xERMQWg1PdutmVYksYzbCSQGhqX
dgh1cKP7xXA1Nky225mOX3vd+0DCGs+sNG+EUESfOKfxDAmvdwwsMpT7XMPCvZs9
UGTD/CYNOkDPrYo4T7YUxaB0ELY5hmQ1tOP7vrcP8wJETx3nBn34oWf0THnWTiW6
rDCMp6eOu2kEre0ynNFkwnRrtXH0v+3q/RgbfNck6whIDfkPfIErAJoMyS9mhzOK
Prr2Pm4ew3EPkrip0LoGLG8nZwQIa66P5Y3OZbGvcgweBvfWCXjF+UBXnJcJqX2m
UbUH0bXplfeqrkr/hsLZ6NVJshUEZhYG78/jFykL7UqaQSk41xOChYfBElrLdozP
JWeM4r1DGaJi0eFVtl8qzxNpqQs5/mhNlLadX8eKtdQsh1LbBh28+WS6NyPxyzPK
3q8PYbxxpMq46+E8AcPlwAc5sPcnmP6BTNqqQ5x7XKWxBj8QrkdrcLENvC7R2Y4Q
7YkE/gQriA91GsupRnDEkmZbN6FRLF2B3bgSCCuGOKmcL/vFdRe5n22LvzJBM5w/
I8jMENWwR7ShNa8KEaimAFqkHQExDnYKejL7UVWogA4It6k7MiO5LfqQ+euEVg2d
EeaG32N1sFRniK5lrLKUz5Sz+uFktxzjid2AY6YxV0eWOkQQDjWaoDFrXxRZWqbm
5I1cbo/78FjH48OWmr9FYaF+HdfGursuacTE1i+UfluO0Ltp7cVRKsd5ypvjXN1j
ddYj5dw0o01EfGBlYoJOszxzBnDxQ8Z40vLHR1bIL2LnX47Ad/RbZDZM0B7QhSsT
neFl47z1BhWgZoS7SfE6TTy11am3MNVG2abrnaor/t23Dp6FB5hohNjh5xMc/Lx2
eYWqV/u9z8CEHQJ4BsVenca/H7iQtKy2/SEUE3aBWgIcxxGfZT4flxZtEq6K0QbF
3URAbyLCsg3t+UYJcxjLaLlooYcM9IXDw5Ph1Ul0hgzf7eYEqNQ+MUldGFJ/XBLW
/YKEO6RK1D8KfOWnSfWuAPv6/vk3d4sCZGEv7fC3gYUtnxeUEcXzmUUhjt91EL5c
ylnHh160vn+OQK4oWRtSIr0VE6A5HwyGInWDP3uWEXJ25GHK8pZJbATMbA/xWSu8
B4N+Li2C3Tkg/utaHN8iQKCCL6QfGhasCHo6onvlv51rj82aHCccbJ5WO6Qe34TU
DHxhUEtvLBdpJGRck1IvXtqX1pWckQc9MvK/J+wGlGHeN7OcowFmVVHQeiSD+OL/
YJFqFxyuZoEIc58POieakkLK70pv1bLee3zBR4Oi47Pr22L1uLemQDSIlVlwjSLe
/MYAxZj5Dk+KDfbjLeqJyBpo63QKZKMk+kI1EI89z16z2ld0U1pSl2N3d0gYyrz4
Vka6yF8dILLEvi9Rt0MKI+BYYBXm9QDsW8MDeDAEQgOLcTkqT1mUyzekmXjt2fLn
TqK5aI2/C9RsM5H3c3qn/2Uo/cCpsTp3jHcnvw6sGkI8spnoF1FbJyweco50ymPe
QQfKYIz048+m9KDUkl5RVvGUZRlXbNRWPw53AInL8+b1YsT1QZc1p2bioJPTRU8r
8pOE2NH7h8ekyk2TUG4IppqXnKseELhuJKR345mkIXUGhYUMD/btnfyRFFXbLimW
6mItB0cE19cbgkhbuRFCfhsBn+NqZwMn7TSH0kb7ztBrJ7Cmi1pisFwKj61tJbPi
D0AcegGP+7mOHaiSC0VhghDACXSsypl5WL+8wVPEp/ZifNbBLXmtH0bxDhO3/L7X
X7k7KvbOYnNu7IWU5qG0eagxsMbxrJIJ0iFBBGRZwrJpGTiEMaLNdrAuLevbOYL/
3kSgv6Vk0NI1kxmtlJ1rdByB3eI59ysG8eQuDRfDj9ZxaYhaM+AswIEucaBfAOR/
h2MouMkVSV4sW90HfHWO12FE5X4arQdDY1U1w9+MSCbgvfMMmu9oTuhU0+4mPpS3
s1yQmoLYgJzCasZaUstpROmBxVlSfQT745KfgX2MB1Y4wefm4mphveQXC2TT9xPW
QaXevaxa8MvCtuqvrwQWqWDZK5H/DERGre9VyskTeVUBDTdHxq2SOWLbeww2BSMU
K9XoAX4X53tUSvTtOrzDbcUHRPbmw1apAmBC8IAVnTuKb9Xb2ZSO7oJpuR7mR54g
om1af+9n7aHzlxKn4wv6LflNKKP6TtKLUxOgX5nyPaFCXXsPd6qRIb+mgu47jOwp
2Habdvy1Wvh+A650DmCYA3As5cdcRpYrl/ryENms5qmZoudmnsKz8Lr7HNqRsi9A
Fh17GT24HFl5BV+devHdA383NFtQrBr8S/+X+c4cvy1hXHs54a6XlqhP/fCYHi5j
0qLqm8rclUuJWuXghTjHN0hbWsRkIhY267sl1DfeKiyC8Zg/52ghsBcMC+/pIBi2
0l2lCc64OBemG9J9NwPtJFek6YDTe+vJ6AQ//7c6P8mTVsZm6Iooro2y273QHAGe
oOfhctZraDpR/4l3NzpHHv/n0bl2WNLlheKrfJoBVtF6Q8TYK3VLiMmpBwftjeqm
2uLrJxjUe1zYFFudQM2U2sttuKeTjIvQpMTpOMBXEm82cA+1fVPq66RVSigOainH
Zkwtd6ZX68K73O9OF/jc29stjopONaE6IvjF5xVAq5vEMkSTPAqXbOHVE8g0A8MU
34QVfDCswq3a+NMI5v9XTSI4e6nbBsjzpsKpF6dj2AYTwvr89bDq2UXN6+Jej78A
3pxmO6wt7mgEynfh9dvSlhkt9bn5XhAUMor1vVRJwQUJSuB8JZLFljmqCLlOUBEn
zFkdRCtSc0Fy1AYFqMVKf5fhtlqXhCUeafItw5N+Z8qTleenFS2PZn9zKLyyVsoc
LoFgcmXkWsBIGqZqR4hNhgYtqsgbNH2kT2SoC7oqaZKVlnJzocI6dpuI9XcLvKEi
Fb4i+/eyvrG7dCrQthzWPFXpJFeDPTKtzUqsY180rw3u1L0CojZjBddKkZ+lglS2
0+FmPoHk6QO0WlruBQrH47U7yrU0DgCkUTbwMmUS0fMXjDD0Mw/r9GfBcEjoN/xz
DY/4YEXY3qOW1ldS1SBy2op3qvzyGCFE6U9g80lYUN4TQTrchKkBjCda7hSJYEKi
1HH2XxOUXag1Utl5kNXAt4W26lnPYTerlhbgU6fcA7VT8Ixg6v1ul/Gs5zxZJVmX
XUcGunKQt3iT6oLCltWWZU9McV+wShqVAutx5OZ/a8g+cMnFLloygXt6DRu9MZpe
62A7e+g78P/gGG44r1gm0n06G+63nkO7c+lBVVR2jtroqptBfVVfqbUc/QdOi8St
2h6mY+PKDuC8DW6EpczVroY1ZfX069r1eZQDxPTjaW3lpCISZ0nF1oHddJYRBvbB
9uSMbJvplpkPfS9or+GIKVX5ouGM4t6Wz5yFpGI9TEh/Nsffns+k51flvVgOtQ0D
wNvTvsCkmgvkTxUqo8xjMPB6+4muwFfZ5YEAdW5EBKmjD/5GseG+Poz7M+4blnKQ
ij3NYv5XZOnF5RMhPBm26nb6ALeqG9pYgFSLxl3nO4Ft/s+hP7YieowNrJaZ488H
HXfosounxz1QyZLxUBkjngkhp3aplvUZDtELL9D6Pal7o4sGK8uPX50WlRgUh+ng
oyYkWPv0RdMmhx1ntYdnFw3RrxFF2jxspt7BnXILEt0FXn5kAqITYkY0v3npVx+B
D6wQUYMb3eg3/RZ6GKkqE9BIlrB0om6hfi24QxRYO/rSRxEhEPhaZ4RnCheYoh3M
SFVoHXQZyms0cHZDFJzoSbJVTXPkV3psTcNBmIhBYlvcHFvR9K66GN7UI4vGuvQ/
ojvQz6IHxh4JvWCKsKmcgz5EADjhyXV/lkczegEH8ObDS6LeXw491KSPd4K54yWw
CTwr9Q+bfiNeKbNC8fgi607if3HX7rdRBVPMuDq7H3Wy9Sv2h/JSbMuWePRWqS1H
5/DtPxc07PVn6BnCnbr9e4uBZfF34ipcO4Fc75TabARpJCtjDe9dBYyNDmk9S5kk
iI6k2qd2RrLQ7YbMxJi4NQ+rL8SOmdFAN/2g7nb+R/iNe0oNNR4lRdvXAllnC5As
QF7ib1mbLDXqPNIPGRUAL23ZGpTKMOJX6Bouby8Mbm0uM81l+VIyV909aJGznHIR
Se5GMozfy+A2eBnrpu+LKS8cM94IR2AZy2zubrOv2SbfhGFWrVDDsTge7xybarGG
I8JM0mPkvdg1hPkKcFITJNDY9fIvXiku9Ty1LAuTeQmEJJ+biK0ule7VKaE3a+98
iVgtTXffGcDb6Mn0ZM0q1E3MU83p/MOEur7Biwk5p897fc1fFAbdtdDj1LIqMU7N
Q4N25tG7NQGhTNDGMl/T+KG2IW0dp4W8BINK19zeK3ge3DBAJBjlCNKrqR9O2CRN
t/81YmsTkGiNZD4VAOEQxGV/ggdB63538EBzUD7puvXFq6T9ycxt/25E8yrZ82ci
+aU67AOS6/PtmmS09LUR/0d8a32BoMHG7fV/UOZo/yI01nCuMTZ+MwiURsQoY6+j
SMtFx7SUVQQTR7NcCGtNrSxebcmlKdxqQYV1x/WCnBqNH/rUaeOtVVq6Nv56h7SZ
YglgoWNhCEAyeExHZdlD4FPP5R2+Hrsf7kJx14oJ2QR6npkVooRCceqBT2+u+2S1
gkdS1yEbcZE1QZ4Hhon1U5cMPlkVD2MGeOrERhLuDCRjwFy68JwySgOL2T5t6zu1
PEnFODaedY3ejmCLrYsmsM9cOwmPRwgeJL60egOQgkr0LsKCd81wbqyNX3Go1SYS
tbeSl6SBphLl0yY+BmYL99VvVNObeqioo9X4k7IIziAr0B5O/6HgiDwtKKFzOlem
V0xyMVbxQDcHkh7dyl8Zx7P9HHrwDRs1f2x3/egUfdziDksjiCoW2f71sUymtOcq
8E7GA0L7OfAa6pQ0Jo5w03y372Mx4+CmusL/S8b7hDxsJxGED8T4JPbcc8D+4pCv
gxxcbu/MAUw+xlahv8EJqjPTjDPWaEbeXYVuMU9gxijw0+co+z/mkzgSDdfqpdUG
rXrtB6vLz3y592JFUmYqfSqbWGWHxEeSpKuVZNYBBhX3xqywjvCYXG0Wqmh1Oh58
HsWzja3ZqeF0yzmyPo0lu3HtgxnN9yTaJR6+1mD93McA9p+L7fR2jigwrfD2/f+I
CyDSw6B2Fo/UgOoxaQ8Yy2f1e4PQXkfwkycw/LDIVdpeVJ+sJMxW5bVLR6taeiul
lnYb5qXNtH/Sxmd7yH+hMcmd717lff1lP30XZpafY2rNIs4gVIWsGib7y6tSTJ1z
UebP8+qgycI1q0EzqK96eCHkvbd3gQU5hfUCDLyrq0BgARpzzpLQRcRi+ILzKEyr
2azyaX4AMFu/oxl2Dua5CETwmySrAXk1/yLTbZI/YIIcjwa2R4rhbuActR3hmMZF
Wkw3DnfOV2IgAlQDujoB1BmzXjk5U4qQvxwNbzDuQmmsKpVLy+ywX2rQgXVR+n4J
A7xphimzPcHqCxcKGo5+oTkA4m/Wj762I/vkUzBpMoCMbbmaDMdFLQWXyePUoIvU
1L/oAeUaAwEBCPLg2SzEyiHq1l51WB6LR1nf+8Bu+UxCz35WyFUIamUwiSQOd07s
YebwlddZMIPkKUaMEf73RhC4NsdlSsyDG0QGk7dTPGmP6bSUAd6o+MY0ZdKCuglw
a4wlKuvFhMlTThNNymuc2SvUvXp3fmEdH6TmtSqYpoqwfnf9xfaB4tukhi0mBiJY
EexhZ+Gdklx9GsTqFfPrZh38+WNUjKFqIGyEAquI2fQ7NWrzTa/lh/10AsSQ/yfr
Laj1fXLAWzvHpNXNbeA6O/Wh+/wVYGfw1YL3nQ8sA3enBMto2cIOOdimsMGgjJ4b
wY8y8rlG47+pJwZEFdMBla/ijeltrDikRcsk2YVTnyv0G8i7FkX450u3X9F/GapP
kuCQFPNPDc77pjaHVaT04ydY7fQuA8glatMQHXm+EIZqwj8O6mpztmn9YUEc+7/O
4xoIjItDyvDh7LI4GiZ3RRMwygQj5rUJTbTMdDBhRjBPx8/6JYFtxHHSznkiNHqn
Q0NiKobXK6ZO5MYo2wl9nGD5E5KsHUYsMCPXGJPdGfUhOdcll+jqpoFNbrxU/9j3
soXS40HVWQsmGfoYsT1m+uk0BZ6VbIEi5d7xrUq4oAfCvIbcHbO64ODvk4naUL2w
0qUOv2byTFWQS782V8u6GkhfAC4UeuYjOab7ugGSPhh305O9aj/Gkms9c1+92MHQ
RBTkf4YpUYBSaIv+/exKPxyt8nVbkB510OAxlkLBKc0Ao6OpDDbMv3QW+GB3E8LT
y4l2Dv90JZU7FAoXTOrL2QUCvCP2ixt7DPC6Nx0p5SU19HX7d9/hf5eArxULy1Wq
RtZKaD/iK84GTEcpBKkEF4IFycnlJmNG4CdxwEWjkWrFn3g8yvuMng1Zl2fEqfkM
QeF+4cvLsTYLsLADmvt/V+Ra25h1739JTOOFkf9TS+p+s6FOO9U08w4gAKabawLS
HkhojbTnLUyQpmPPwTrMqX4IJcbKyDzUWQvJm3jpBRZoDQI9CDAdR1G/xm/GE1Hp
YWLL9eXD9zL1X+0wKVjU7GZvbHODUZbof3/J1DAjxNg1/qcJhK1GaGKih/tK5E26
i46dFeSnzKjPjgQVfl7rr+p4DlqO8tsrM3xh2YJf+RmiObE2Ob93yXDnu35EZTV/
xlceUpdauxQu0g3HEeJ+qX2TT6pQIqBtDgsMOfCcpbFYtE7qgEUbjgFhT0UiqsY/
dFVnO9HRama5s1keTc+VEMRZwqBQMj5O3gH6vVu1UF8RI+HmK+lXmga8q/DhXyXy
qUHei8XT8nuqmFA5yQm7qDimskMsTppK+goz4U3IB49BJ+Yem+ijtsm7R1XISQ3r
uYZqgWz4qlbup+ht/BenSulcUuCd2gCDr6eVzQK7EH2OCxJbb8+h/uBdmNFzWdUc
qh3bDg4Qjo0AdqLux9EAG8ccdx/u5agYyrcLKUhTIrMHJBc2QWfvUf0CoiM8L2LE
6nEpMukBar2Edd/+9wAkC9dQGcslfh/osZG6OgP91Ju8Pie7n9f4oLVlVT1nYLmr
fEQivBSq7B5Z9SL5h6KV3MZhUMowyTRj8JSNMt8wvwxCLdgFS5gW3rqbiLoIcL/M
yuiJL2mZ/HU9vq32/ZKbGap8ACTURLXNPVdkmEsmBQFwKjPgCRi35CF+d+8CLSeA
tPILWEQcCNt9RD2GgPQLPX54kIFZerKGw7XFhfABv8K9sV2SWIsfm6GTgMAlzioq
10KRih8MulrFHwfAuOEiaDLG5g371/Bns+1wCBbEOVqVntAH0EGx5KfEEKspoka7
qWc6sjCK2JIZ955eBD6W7DCU1vsbz48Nu7moSUHLvzShB9CxozVe5J0/mbOvMvqr
YYMaMx5Pky4bAB2sj5+h4sVn/UwxkzsVf7bxzN//ZwVdTR7Rlb7LRflv917eOSOe
DzD5YdtLiyXuE/TI5b3gI1sviAdXlTu3AC98ACUs7iPQOa6cmqP2TsO+UutvLtvh
DqT/r1sTBEFSkS0H8mwSGYZj89XcdVICwviWLZNmZbUd83GXyk5LPOZ6zcPfYwQn
IsqwOuBy6pLWsqArqDOiv3/lOBRYi9XJzb5b6hRW2+bBG0nUxsGkPSVHaaB1JXiV
3Lq+idL70sR0ciy34veZDzWvFIBQ0aEKgh3VGsIfqPDj3nnoEy+r2N0mbM2wDEVT
4HAwdKsPOM0AF1cwuejivemGhRP7x/bedTkTWmDSjDj2R8YNKCtu2lb+tNL8jeBV
uDrbnZO9bdrlHh2H9uBnBZwrcXtqm8Q6z9PY1LTTKOBzuyUSW8uJWhAyVDRH511P
Ow4e/jN/zJMgRQYk9lOYTxW/zURk3FCIF1nq2fhV8sGs5bd/XNX9Emi27qR/jhbq
zPbHbA9Pyhl3cT/E8LbP7Z+SLixrefJL5Wes5T+lW2sEcC+73hmGjUaSlmtME0oK
63PB4bObbp8jw4bE4a3UoiHt4q2VyeE/5SBkVlbjIPBiEPtXvkP/5OkyCXy1AYOm
65xmnWUF5N8Dy9rdxY2PU9bA/ze48+ufWRaQW5jPDDWS32KyvawdGwEHQiQDB8uW
q72HwI3RfYRUc3+icmgjriZaboyt79NEccwg6JCRLzYM38NKnsReq1AFQ+/qEm9b
alniPfPdOIb7EJ1aT7DwFu6+Ap/hXPil5AG+AjmUfb73q6nu84WAJ1EOufXXzPFG
YLgp9RTisrtLBw8fNgAChked2PmjC9qDzhEO1G+jqWJImpw+eq7NWoKJc3rCPm8k
9RWUi0sJwTB3P+b4ZsTAHwa4iDFd7iVxsv/bGaea18anGiimcy1JNhqKFgluiU0V
m4WNQzUV8phpM5UM0mDlp2FAQDofUh/orhyQ4uOzy/kB1/cgrOsv5SUcNsxDhc2i
UCKAWB2T5j55hMBFq38/+c5mOhDRICydHlR6WbigmQ6gMhW2wx/amD7j5TYoJhBN
ivkc9fkFlojAcp6sTX/DXRoUOt0GKKyFrK+yPiAtXlld7tPbsns1AXiTl3MQepgI
+M2NRt+TDYzgQg8j959ChgzmQywrq2LSTBVJPGlMYhBYyg04q7yqqBn/0bckX6aP
ENYgCnkHqUfvqONnb1/lJOeP2zSRwl0njWeGypPiO/OTIAnYmeULvrNzUd7w4lz0
75LXKfd5zIGgEwxIAgMYSRRRAczmlknOgATQS7K5bhyw2jcXVcAt2GDgSInbAEHx
Oo1g+tpTzEJljKT+ypxGH97eYvd9V7nnWWSD8i5ESlZVjFTzbZ3mow8Lx7e8R4nD
kW/5pFvqaVac0rlpNMdK1EYYVKifIkvZhI51Ijdj+Mk30TDGMU2+ziYhSWuq9voN
H8khT52K8c48iglmwMRUz5fMtKckISLE0zxOHYPseqZVb06pIsjlS6fAfeSqmND3
qKykVby9rPC75ybnkaTYIfb/rq1CtHJBRJ7d4md3zvMvFo5Dse308NszW9F5Iqc3
XVIwxt/miUR4mCZ8tgCBRnpKeKSY2AUsDaLQbLF1Q3BCrksX2pxjoepmaj6dEskC
GsgbVZk44ovgamxgab7PYkPWamRtJam7Xwm/bbxE1Y99410NV5tuoQnF1sUQ1j4v
+xr1IOTIZiKD4c+sD6UftBiBCuhM62blEQNhH4KqiEjxSiWSnpy55C4qbfGbIb7h
oyX5YtdWAoGnGbllq8fvDQLvMqBLaVe5yDwoTv/yG2ebK/8Ue6FC7Wm1ybeG0JO2
SpSzIYDXU/JFZP3aUsDz317rT0xIhQKRlZ93Qw0OKlE9f+nexIBf5FKVIGvi+QQH
atSvUzEUbv/R8p6PNK/5SEJOtdV/cobJ5TbI4sKkAavwoSlMJol3HDkQin+UbEXe
5xQNFPMkOV7LM6ELS5P+12bD4YUgMYn+8NfCfDYZidLDJtETnlevt9Rcatc7E3+J
o0A3Jxc4kiGG6CAylCDHdP51YBJ0WHo0weith+uetItkS86rvRlDoNqatx/bWlrW
ePdGYa79XCvYlVIVIJflt7DRbHwQ2cqqFu8xaO5gcJgpBCrmzAIMleemZwEgR4oi
kGOFm/PlEUCaacsm9u/Pgb6aA5pzi7FxtaIQWakELMQfLFB/Qhu/dqD8bD5Xoryj
VwuGgYgyhiCevWkVGKEgdZ1uYWLetO3iiPXAHtieFXEoZtV/1WPjdIJ+n99jBTuk
IHB9tZvNX1w7xkMYUjBxAc2GeGLMAthj24bmZ4w4l9aoh3ILBZ1NxHEIl4R3Fyk8
T5G8eOhzRwRC0RDNM92BXAC6EfI2r1WX92JiNAlZeESv2Xsmkmdm/SQOxncyV4sK
Z8gYTmyu3gwMUGC5dg0/eJjAWdMk8dPeSf5juMOCwdTbcAswoJLfjzk7ko1zSiPM
1aM4i+uZKuClMwg0Rw5qi6OVTvLReymH4RF59UFbLZ2cGxafqUzojWKoN8pvHeKE
E9Gg7GgpGZpaHiKo3u/UYRLySNBzOJAKWgNKGAc3BfhXUipCUDpmHt8kc+t5Wgz/
3MHlZlqHgI8GRNuvek4qPpokZPqMNiuY/4MTpQzmM9vcxh+k5Xv4LthYOtwvOIY7
IOm1v/+S1oiPHiWBN9Gx0IFdj5rFXaGWrJJPYGvYBmIIlwgk4Yuz399x0iZVe2dO
Lk/ZRbX/igdcE4hZAL+TJ0zL/rChv0L0GyFO1dbvT13DiwQZNyIuFfT+kQ0VMkA9
uaTZk547hfX3fLqVOcc/SsanqvhIzEdT3ylkgnQZ70xwYC6GfoFW/oYqhFPfspvO
9OIq1x3dmcoBlVK6Ggt6Py4py40sOyF2EBT2TL5VO4Y+2csAGEJzKcuiyfzIzR1S
yZ4E9gfyBICjSMT4bSHn0S2uvNLGWvp3G27E9pva5Aj2Q6xCoYeSljICLsFhbnPP
OR2WVFt9Go1SDT3/jgYAGKdC3kX4SPr/LC0CYLme4LD8Ija6GtwZIuUddRvxG4ok
Ri3UPmeamOs1tFIiv8SD2CKtCizQ6eDN5sU9Dzg0+dw/mqiTJh5YjA2+0ea/pBHB
qWwEIx7dUm8ohr2bYZGEQsPZeHjLettlAAQRv/4OX+c+HwtpkgGQScYQIbuzui59
s3qv6bPQp7LfdGyChb4cdTY9HVMNx8Mac7Sau07Rz/MqpqXtD91oUjfDj0fxc2Hr
lPBoP4eY1JyYc6ys2JY45gI2WIyL8sXFDcSRZyQG3Ii8pVjVrGK5LAJ7h+U/bBvv
NqfFShPFVrBRJy1uKp0chcoRNpues1ww4A9O8/+lSVypD63KIKqvkpn5AfpXtw1y
Km9l4fTXpLreoeYJ5zD6Ap8iL/gLx4op9zUEPhutSyatEYk1DICqKsDYIdsaRprq
Ug9QtPD9K2prAFSVUaJkEFHGo5ajsdDlxtbOivewbH3N4gOax/oy4wZGezSHsdwo
pF3SoKhnAXnr+pX/ncyt/qKE9dihXxqY2lRpjOo5lQm8HO3dr/b/NRryaxacH1/I
k7Zzsy8c9ByCkNW42+n5lYVGmnhgZGtqiaCpGj1h2LBKNsX/VraENkovsnmfOzkN
MRAcB5wzmkksHXE9lLbg52fI01QZVipzuZUKmhmDjFUlvz4w3bn37M/FtbmuPDFC
vPWbGzjr/wpaKONSNqhTSJ7UVtpnG/TK0SaafNzq9k8BU0GOXeEqy5vVNa9P2B0d
2KzcdLsZUWoKdDj5K1BO7bZGBHNxZcO9jjqWWB8ywBJ0FKhmEa9McRaq7BvuG3F3
89epEwGFitfDSi//bIZ5F2h6iV7OlyVELVhNCRP6ob3Q03mjF1OtS4opbxC0d7Yz
lSJux3DdQdbMM4deUYv7A36vTklGOTmv3K5gzIuTEu5vodkoNC2odx5HFvbDbQC1
ZZDTt/1hzrGKN+O9mFlH6Mm4hAzkeOtdlc7jn2Ljfszv0bVaeRsWbVhFQgfsyLI6
pjn53qhpRmAvNRhflrBy71XIVTaNDIr3s7C2hmXIgq3e80I5NqvrVirOEfXYD9Uu
Lj+ARyWfQKi0+RZogNYWuzLUREl/NytVnto29hQZXmJmmcMx3GcET79mtqi+GDFw
z6ogaAO/CjV2JyRSh8x4/3nxC54iowFtbrIi4UkE34DPG2iBOLx9/5R8u1Me37qj
+W2WIj1BZSkTtyA+Cg/9XTfjFXfC9ZZdlIp22twNn2BpFMGHDEgrImSO07/hqLta
DFfcaeqh9PQ4wE0w3swOfEx/RheK6tW2g4CpRUZsAphpLkO9egrJT4oCw88aNrcN
Sv4wfaDhX6SXnkb+Nc1GudPhLMhnW2ZwweiBK4/TjQPIqz479Z1rFd9AlGR9Pjd4
3syd7cPz6q1bETdtF/9d19GBLpJ9aJVCku40545dWyucdRKaKMQzu0hUrAgrzxsB
HIynF30Ar/VjC4l13vwVhqYRRBhdvGhtT7uvqgpRJI3bU9aM4Dba/WnvQtQ3bbqe
N3Dz8NBlXG9tXIa/KhfUw2rLl4fgh0i+NxnISbfyDVAecMUvVqoCSduhFZFZldV5
So0DtYp1BbOyUyccHppsITG+2LndDSCrGuDiOd02nuK04kNedlcMSZlYhyhY+uB1
x7BM92URe/SFhBiOIsfZ5iy3DVHQrtP4gKhzVWRx3QmN7dWIEgDp0fkqBd+HP6gs
wthYmalGpyCoArU8Yz/aaLpvdgXKkRCtnf9Hrw2vjGIu/bdL3uvsLdnHv2aDLn8w
QeArItOoynLBxSpy5bjD2Ort1ibr+byPm6BQqkvUJQ7R/EXo1jYa9cBQRqPgS9K6
XljEFLoPKBOPqbGw/k1wC5cd/+ms++vvY4g1CGqvADF5lSN//a3YGgZb3mHcEbKD
mB+3lmpMOr14rlwKu9gmiAROIKhaca+GwLZHkVKDxoglAcWP6BvvtZYsR868sCy6
dlW+v4fPqZ0gQiwZHFSDkpU9O9cD12Xn1Ox32Z5/K5qQPb7eHpqiuxu1W/QFTnl0
6qF93Y7TZddfKBObPu1zltx+QldUEdVCUT5mDwxhqAleo+9H30DhxZWIt+38Z2ZY
oMSbH11prPyp0roHLaISo/dkAfcGMgrHbbLM3x66c+Gu3k6M3BtRF/Jbe9ZJZLm4
I+myzb8mI+7J6TZZboXSO9KzerqMmpD8T4DeN6slBeBkRlZ5sHGahdQ5oquIfiMJ
YumMRCqbUVy+D99CnB/gSNUIYEZT1Q4O2LTva1xei6Sph5hEgM8qiCtsceDLi3b8
au2OkYkmyBENlDVltTgt3GtdfZzfKkI6lTvJp2BMx5t7RX5vrvJCUUC+GVQtpW2m
EN05I4hekNwayEhD6DHr+MCFcUCfx1kqB6CJdiFdjZRqLOsJKRdYws2rMG3cAaH5
tk0rvVJ73RtOGzwxmCVL470x6DZvSyPiUvmiMktXB0QcTVK9ETsmDkI4Cj/v6u9B
WFeVlf6n12HwmpFAa0wra20b2sFYXiqklxNplnP7NsVcQngmehDsASSkjlIkaBWp
3UYvf4OiJ4MqBf3U7Mi6AYWhYQ/ASvLm75jAyM2lElOEw+k3czzGAhlfrrqMxavr
GYj3c7VIYa1xsCf3e4DMNUIOoj7GqM9aYHWgnME0KUKumGbIo8zInF7u9CeuXKfA
Ba4HYOMvBdVSYmZBedTwYzAcjs09LfNIAP2KjzVFtbNh9/ngpVitpI/P/e17edxg
Dnq1wBUJaritwEslD9cIpDRr0x/BFeTQkIVdgkQ/ZY42sPsjQdI77Omj/jP2Y6fC
Lmwha1Uj6NDpRKKKT9d8gtMmhQkVtnU7qXFl1caICAc7HN/Kf1UrcgGkiPIZNLCe
JVXL3KGpNFMyyIHLsATZqBmiCV0g2BGQslQc1o1cXuMZFpd+8jD6ZQH9N6AQeHH+
mF5YcwJJBcm9q/u4O0gz+OtsA9upWsTMnm9lYOxkJzfnNEppebYjQsYJwsLx6i57
spDaHI49SI7uFmqURLHhDl5ceUJTvUAJmwVwFZBxZRHfeOLiOOMn63hLlUDvedQs
CZfdUjGzy+j7R8EC6AXI0j8/eX33DjHKL1I+uM8iD6Rq18dM6q5GjiTKXCo7I7Pr
DGQObMvfJ3Pl4CDGsbGxB94soGSH8G2tOOs7qEuo+SOt0rSzSt/alg1oWnVm1jk8
wMmb/eGa+3rXJc/0hkrJ0nD3Jfc6P84YBiguN0j4abVyo0aV8EgQjJ1bYViTZYEV
7znmEv3Is+y6T+pv+bQwVVFId+ZSvb7X7C51IlHXi5X5UWXQptErviR5LtPzXg8Y
vXvxrOyhtSDv76K2FcFs3GQj4RhhwLtpFmvWJtu2xqT2TfSWUFMFCGSgF4MiLWTG
6KCDzPveN8RMTiWWesyAHHk3SUJisD2sj2Vq89ry5ktZBKC5q8TH9RF2G+o/1CWH
eOKv9CX8XKysjGH0Qpr5WBC/ClSdA3p8gsehSSwk82BVSsnqEjG0PJCDZ4yNgOKv
C+lCKdJAsC5jdhnBd6z0kmt8KzVhV6PdBCdVsbHagthZa/4mQ1rVfNJqj7J0EUVF
b7KgXcalNrxUQztzTV3dD4nS9qno9U5BZtrmclGtnlccdPBGksQMkxK52EXwWlmk
BCEbxxmZJO53sZ9xjppV5QLDN8lH8+rTFB+YsWYqanLgFicfI2/CwPLUCQachkJ1
36yQhoYh4u5FjaXYUAm+vYnmtvHWOdqO+QUq7fe2eNv+vnzFcOxMz3bAr8GF518o
SNn/O2o7LBm247LGkmDWLm8OtttvjWpYFLjrhNF6Clu1obYB5C+IBLE6i5M9BgeR
tYjMbggtJ2/m7YLkrJbaaWRev/p+1rAtPiixpQt5UmHmU/hD7bAzCrZVYNTU/seW
oLseOhl/XDUoqRfloBVKJcjFHW19LWG5X5xGfgL7q0DFik+7HoQ99CcLeoGX1nkA
mNoWAMBXHB2KvZe6Z8XcP1w016FliSXHgxv/Ms3wn+L49I3dIa1cmuWTODb1iBf1
CQigYR1vSMo2ZoL0EQm9/HxvauMcQqrn/nSI9rKB+ZpjoD4Rt6guoHYuP0tXvwVD
W7V/MR4rmdXAaZ8upfw8OdR4aiRNzSmX5keugURu0+4KrFt27Msfajv99wUn0aom
mAx/9eMVgjwNDkAyt9xnURTdpUX1BAs480tDew2meJ54XcCMDNBNhqsOXjC2KcXH
0SlZPdpoXyak0sD2MkrtsUiiEaYw74FIJAFYemHvEBSZDlAlWRiJqUTmEdXQ6gMz
lWVjD4FLuAb1RYCX/baVMTUFXb6l6619CkJHKwtBrseeOrK8ngq+izBkTTI+VxcM
mRhhyHkJEUEGzu36JedEEi0NsVge/U5LCWFxDEX9lwsa0mWRcZEsl7ko0UiJkn8V
NItm2wHRd/QgiQI3yCH47ecf8QGKpWBmk7lFQWhBt7MyOA/ugF4iQNmBJlSYcxT2
AzuF338e2N8X7KL3HH0vqiCMrcQ5y0NuE04F5fRkxirDEog0y8uV+yfhVLwbkWsw
4Vgu67zaV5ST7joxgTd2TZdZeokJ/j5Tz46vyGqk1cnwarN0gAnoiyuGeunhdhVV
83Vx9Un+HRqFJC/bIorjYW9CyyQ+zmUdHOHJUzteQ+tDiFiKhfkCWbvfcvg9neTf
zsasovCABWHPDxBw+JNzhUiibv88Dt/gC3suvUI3HtCnG02zhOHbU7I8uE96rsa/
Gh9QuhH2XRwBFKSwYH3YhXCnte4hqMyLtGWRBgZfZS6t4b0sjb/6r0q9Z9iCecQz
PA9SPEiU4xGZxEkvu4PJI97X1XYwEGcesNbdudyL2AAkKmR24OMhO66KZqOEE0eB
VwS3EhdThsUlxF2ZSogWIXzMgyblWPu6bthnwgymFhZK9SUSwvYrm97Ak0VgCbHY
+stqS5T35ihZ26Fs5WNfXpiEeZ+XX8PNq+TSsCG/sLQwTRjInY7Zve1B75Orp6pI
pe4k4+gIRsUHKZ2hKn0T+5WBAQRWBn+TrmxalupIJdw/uFSibICOgTYB28Ick8Ay
mreR7G9Bot8gHY3wb1KLhOITuqJoponMvEf3Ce5D+jR31H3aBwVs2LwSf49rIPa0
Gg+Fgdt5+22cESHwP/hMVF4Jobg6LPFM5gbAYxo8i+/tLERzVBzTk9JHYk3sz9cK
/NZr+Tn6/u0OU+x9xeRt4ftgTXIu4KC0Gl5HfTiF/yFMK4JtzNQdiThHxagIGyqV
D7otIE3ynFXX0zcA2bALAOmgQgKv+w69u9g06E84hLsWZi6AwGJ0OR5hXcqOi/3h
+7haqzDxg2wjVlzunDfJkvALi+IRWijJGbd7h4EM+ifKkNCSUHZdALJw2Go/pGEs
xRxPt6zws96xji+in3r1I+p+9zOERF1xB6swuPirchhe4mAqXhkLMjFdFZtaRB9m
ZYhYPBbZXw9g7p6UfQyT3cA0kRYEHVtXWMV22SUvP6lcmWvxQ7ShHdNkp2d95NOh
paqGzRBUmhPp0D5WIlI7GU6NziV5KCcDXf/A1xd0m1bILEFC5iDX6KMxT+V7liPb
k+fKMa1NTjps81Rn27fsaY3wnAPsYQn84YjK6Gz/NHcpmwsfw9js4eN5WkeqxCuW
0ByFVowlPxe3llvmftynbihI8mMTFuhQnZjfKf+ItvoSPm+nGtLpcNkoByRXluta
AglJYqNE1lZHB6V4AU5kl4z6KSomVELPl/49P1duTZqzufsRDXImuKbAD8IrbEhk
TBxj5nruMrWLGPxfOaFyY6r+GlPRgLS49EIFXuoEpJ1B0SD+KE857pDXaTeCRn8Q
IkFeF08qwZrrB5ihz7+H6O4QEZOKzAaMbHCi8+AtCiWeTYZZKzGnBOhYnV5GX/7i
FKdgCNaLIpMyu5+aHjxUzPdz9qJ8KMwaDAZdDk9FcCx5942cBYYnUIJ+hRf/19RK
2nPLrXXIiEJfv16EhD6Y/WydB/9zxtXBD7RunEE6K2RnyX/0LKqHbKVvcONb5fdW
Y1nZQiskHjKZ0+G34Eo5XMnsGmqOGS3BLZSWdIx6TBPNdOYj4+8oGcmfJhCWcEjA
lUHlet/nSBiCOJQ2nTdKV9bZiPA1gCsKoM7cgQ5t1LoAEzz0/SHCl6tsGr7xJq07
m3xo4ZLNSPnr6NyY6UAo6u1lMOeOOIaCLKoka/Kkeh+4OmAE0S9uoDiTc+Hm+dm/
N5F0sxsNQTRsBjGS93RlHlg/KWFSCMV52mTAFvsCbniU6jihWW4+BEDNuJXyAQRC
PthOHhlUzWdVUkqEjZZLJX6eYNZaY1o0D4acqyKVx+QsMdiaMY0JIdNiM5UFtnDN
bZxhzSt7v8wDqNMHhUEsBXhc18b4WxOW2NoWqHtNj5NAPz/9gSzLMaZ/QWntLLA5
X9Zdr2zj6f5q0I7B25oFS2ypvi/Jb87L0WsDoOmuPGGEB/rmTMeZcnupLuu/O6ft
pG26T7zu1r1OPFctiflSZoW9eEQ0abOfQsv5+2H//smFncNpQa5mDF9VOynMIsgH
FRxQeuJlcosCAHc9B4FlEgajeEpnIpbQoheDhAl0YnLjAwrw66UjFrFYzSsZ4l/h
pdcdT/a9lhnP2xLp+hVG3/rbl3tCXpCtucKBYWhZF3cPPxLz5bFpNrsAJXGEQb7H
anzkLnBJCb1VX5lgSogJBnZ/4ysTP9fCpQqjVLhaQ0hZyuZ6w0b5NRwNOloBGLbk
q8SyiiPoDvQdR9buwmyvFSOWWJF0Hasdz6C1Is3czityvj6hYILicseFJOD2fyJW
Ewavk9rG+tvc3CIcK+yQCCdrTwTl/6e2uNYYkpfs16BKghIoPviF2Rmwkd2pMM1X
jqhRzv/wXytuvqUs+40qMve/0T/A+UY+lU7xSH34b4o7kiH0W57i7ZCsGWZMaxmm
UZuAHqkCbdn95sUZ8feVod+86qHfyHKqb4D/19nO5DI1n2TqNTTayzL4sht48XZ9
HnDrPNhWn774gQJR78lVeE7hUSvAonEmiWAZ+vVcYfSLppDg8UEM/4muMtheXgf9
p9Hg+kHdPFb0OZoadCZ6y6mrv2PY7kkjqdm7zod13isGdrfP3AZEA9PmeBPGy7wc
pbCwgAt8c2iPb9elTea43LVjeHedwN7I4b4D2Q6MOzYNt8EUDTntDuOFK9hblMLH
3SmCdxtZ8MM2L+5JLUuXQHEcrR2nk3vG3RphqpHc5Nyjr7NDP3joQy+W+F5XsQzY
0PzYWdFxw1V+eekIIA1fFNsb/UM/EsBlDHJtfZxl+1QDElSwx/hgqshs89s+wSFx
JQd21VXuAlNb8TYF695hkO8gbffT06xKvapdbuGWhVowRjqLHPc7nTY3u1BlaP8M
bTEBS7Wc13rLO8o8SrwWsOYhqNX8TX465K0k3k9eIOdu9OFmlGMambHz8SN5IeZV
+LBHDZ6neZz2LwHC05u37j2sKs6g//KPKkCH4L9KgbLcVqfgX+p7K/R0PHtOlT8E
pBOv+6p+53HyeVndlvuAGBhs4QAF7Ceu1Uboqy0OKuuGGZv4o7/sZoSzD2Cx/rJ2
hxatmnhWuT7YcCcAFzo5Y+/22woJhEEEH3eO5p3yMWUTcLw2vxu6r4/0C4mHnwl0
s/u6fVVRq6NDpZp+MbE9RYkxwzwlr/K2TT4gbfcO3RVMMg1KBh+x2kuU7w4Pmwk4
XbYHNLgoCmvUxCtZ2OUNtqrqUJYawDsTcRnyvDhG1S6NYnXKcPg9fGbTWGFKWujl
tHXTUezD48xZZ/nNyQIjHIn995ZVKONCAx3BmgN8s5FwjEYJAJ3B9HX6p27hYiCY
M2ydUvUbUPM1pk/7AZAkGgEMEdZ0Y7YJAT3HBjloND+pxf8U6BtPN9kd/U5U4+Ga
264y8Z+PX+4c6Q2Jb+UFZ97d/bndS1G57WdioVP8DQgmAkoEGqX/ZrmhJFxGgjH+
aWLM2k32OfJ6IOLO2CeQI44xHEkOasT5am6y30WyPRdtv4+ByPo8JXHXyWym8Dpt
kdBqYa4hXZ89U5n9EbDmqSQzSD85ORCMlHKNggAd+nVTlUPHeNooIQtSYVXey8XX
3uJK8tA1T2jmA13HeWmFThwggGrMFmOICI4ecCupNeah5wKtSSKj8n+7cpx4A46m
wVVrDj1lhkXXjSog0J6wHDQDzl1q07Z7L8bywhDcy5AoJszp/0wZyfdzViuhoSv3
N3lR2r2g/HYTviEAPhvszhqBGATaEM0PpP7GVXAm5DrL9a+eO3spY2iyWDq0657H
pCBGykSuEZGa2AtHeLeDIPe2K/KEvsuzr1kl8QFtMEk/itwEuEh8ZfcYYN98Hsn7
mwFwLdpK94Jy8MUqh1JJeKQkM1HPGBWIg48c7DIWetq9R/g/PJUkaRi/88s/zdxT
OISYn0eGtcQi+vPIF2qza41NddUidSj/xDeUhr5C1zfK/XPqCDZrRZKznrAgj/jK
Jl90Byl8qGVh3/jEFKenuLhKJ+azH8PLV1SKmR2m/vsfp7bNPtJPGURh3XXX9uGN
Xqlzko2iSL8U7esKrZcYbHbvu35680LuSRXF0gcKf8OwPR8rb+Cg8bNiu4lP8hQY
u/wwHMvmM6GOp0DsAizNvvllBcuxfFAh6vX3cKmzY+s4xBgA+HUjj6ytZ+TQ779t
YoVISpD0mIBxWusrot5vtXpF2JCBn7JrdhEMqTj+MCNWk/eF8tQWF4UVwf7Bj4kb
+FBSkUKjKBpbLide4Z2xQLZ2+8WhNZAR/NzIFBQCQ5bnS8/omfYeK5NEjDaMaCQ8
vxmg/AuDijr3cNv1RJrjcUynxqhCVCXkQnN54Oea6/FQdPrK90DHIqEzCJedqC0e
Q1aCsphjXakgMWAt3S6bcSmFFlRzq0IriocYpRNTQ6V/bmqen1e5E9WmXJ6MOxm0
ltUjmlsHpZjEtDDN0kgZUmOQJGIUrOvkh9AUd9D679MbqhrY9duoZYIyEDkv0llG
q5F9yC4iSCeD+5QgqrjQhb5X5ukwqcne1DOgNaPMKbF6sXYZVtIad61i4ij0jjm4
wIzGTW7i3Qh/SJQC6qG3SxeLlgYBeRaYArjiCNfjHwlLYGP1tKL6CMYG5OGuoaHA
kzbUxQMIOUIOrkc3NjoeacZwFyryI+YRlcMKf30BV3kRgb70quforw6cMgylOgdn
t1Rq5xy/fwb0WevfAtDZo8EBMAQq0GhQGYGf9iEy65kDEpAfaf/NUTCgDsyPB8VN
Rez3oN9t4x50g4cr64BHPN+UMfIL83r6grK9LGccikzW4EgqKoPwaqfoQBqAvFE+
0yH1qL3O8+fI+ZN5hKB/imwqjqsbT0LXCT0TnD/wFKwlDuEMPxinNfjRU90hfGOO
zP7W+HX+K54W/sHpWABC52IdPRTIjB9wGb4AVgIPmQJkaxAj/AEAnpDIuE2i0r8q
enw8zomVcfawBQTcojB5iHR5rCm/ck8jV6XSAlcga7OYbQVmB7ebFZ7nVY8wFPX9
LD2OGO9SChYB6wg0/JTYkjSdg4hLldNu+uZEp+XmY6fSpBK3+AtYHPe6KCxOin2P
8NZQCPkoYd+3XQRXFAA5XRrIhKUgkGf4Sa+FbfKnQ1C202R8LbOnrChJZ87KAWKa
8sweJDd+ShnGCPLbmPJ1G5LXBReQoZfipvPp1Hymv6s16n1rbcKJreoUl/lJr4wy
5WMe761xWleEfqq7EIb/XEO4G4mLiu3MU12IQGCsyZfVj9jbQOUAqNyaU6kQxkcJ
p2PE7hyKOSDVFGOVTQPLKf4JPeeef0RBjM746sWkUgNli5tecSCOdugolhgSZ/CQ
Mopu7sSaNd5f8pqr/qZ4WLp5lOiavn3ZQYGNAWA4mYdOkeKKIDSwZoy1MITj8Kem
HPmo3mGmzDppsHxlwalG6F8hXQK87x+C9iRcTUoxCJxuw5xq9DMx3ahlUk4QWBJU
6ZGcMqpqrcDJhM2NQgO4YjDf9D5howYRKQeKPOkPw3svBkGuVEkgCgEKsD0QvVzu
q++OI+wfALjR9h9OkiqQ7EgP7nvZBRoTVAphli8kilukARuFCEdqf1i+c1n84ZZa
0ixkTRUraNcGwe8j/G4bCzGAINqLR932SChZq6PHz8BryrB261jd1gBhkcIMwXIM
xWlzVZF4yZDpDbqt1jyM62q4XvJvNJPDVIacDzEBW7PMd0gfkH93oz0D4rb1xRj8
AnBMozpCDUdPKfFotubMUdsQ2m/hICRNjeI8R0+MKIs12Tis6kXZ29C6MaE1WL12
HwYYdPGNZT2VRwpt+rVqvhSnEm5f2C2oPBHea1xzAI0t0CkGssVtCpJGMvJpvNE1
s5AfkTvyF3BpDPYboJOv3QIH5N3F92Z/bq5q7y2NdOKbN/uXsu3pgpjf9irtqJ01
iULhkCHUA9uOSHxH+o4XD+a6pCp+KmljRGu+BpTvH5iojVBYNas94cM58TkPcvwq
m6Q4+CpqWKtZxvXAPdB1Ao8uLfU6u7WKkLDewFauqQGLwjMls691vwk70QPN1oLM
x/IBwdATbn2Pv/SsaWnKQ72ZLA9DcAyR190VshGSzQwr3oSJQkIeebo3ZCddCAck
bAzpH2K79fHQZcVgTG7pFSXk9V3tksh27qLtpwMkNx3MLga3ZTCHya60j22uUaYi
F/qyxVEvbuRODiBvF1yQzljPw3Oj11ryju7hkCF/4qF6B2ESVWQ1tXrne1rZmt8Y
ZUqbRVRfxEwctc1F346dha/QOqafxxK2jid1S453uyG32uj7okWKv7fx5CxXFOGi
6ccqGphC6xWfPDB/fab5/NlXgDzX4riQmoZ6lR6JcuB08GlXYb5JdmFGQLIHmYL9
RZg/JWB0zmqtakxqovJeuyX6ju5MiXDWKnQb+jT7J2QazrgYFIzJqK32C3hXt3ur
XrdGmRQuVmECkym3lo37thxZ1IrxPxkjsrjnsCbOY4xnbaUtweHToek5z1xzq4vK
Lienz/Zv6M+vaLb21LRptk+PIMYG7Ku9GxM7SglzZxBr/wTGVRXzAqka4UjL1iDE
eDha0qCjjkjZ6hBjC6qGOXbBspPKf/+c5nBZh6z+qNjucoKmbxPs6huzKZ4vUbEU
ASbDydeuyzFkKb0qVwkl2DmTIXsUNx9A98nhConYXARGg1MX4GvIQN0+Ou4pamsD
9PmjiseJcNAU9txltovrpL0Kf4J22PztAau+cDc5LnmEF1pjtVYeBywbt403bjm4
9tFay+jHulPAiAf3NGK556kcZVHZhnwcft2vqF/sAgvfMcOxE5nOW9iMSffsG4Wv
Tg7XiPITGXAdvNnQrfZGO9/hajY/8HLGE0FPV/fsGF/1NlwfRr4b8jTfuNdOXAWf
Rwh9Z7a0rlLjSBXEZVm4pHO4s3FDclMu9P4CvGRJ3r4O8VHIzpTbKstjyL36bRxl
1N4umeEVAfdAwpWdAI5HIGZtREhq87MJ4Tku6KT8e3Aj2hjXnfXQ3HD00maTqtC1
sv2UIoqqk0fS82UsEVt/4Ch34l4EfnRxXzQBBQY99iosGu2sXRLAveHKPoeq740w
Xbr1qVpH5A+SUx+HWl/gigCjKMkjlo/r2exUpzS6lTvs7x5UfaA3civcfgjv55a5
5kRgisCcehZZDXQjlUwFDhWHA057VUgsT/znGSipMg2dKTemAfVuILFLNzmjMCEX
2Goj0Q0hCIB4yfjPUstcf7ZpHw0lbWAvpMv81k2CNscsv6zquV/GVtRSYoUEhegs
UCUtShYozfQgCoVfW5hwzV9bVPneocZm52OwcrxChgHC3jFkS2Z2duvhlO/1WB7+
q7OKzYBOnYW7iBZM0v2DOfs1YRFqXC1e93OKrE8RvJzxzOywICidNwM+B88EHCMG
NFMVhLXmbse18b0j48ODpPpA+YfzRUINgAq++Gi2EcJQ5tQZHJsB8DSYSAQ9eo7S
Z0BDieITpCqBDhtQKQfnWyEtj4kBWuwen1jJGohqt9pNpB5ZDA2nP72ZQkxzwZKO
TqXngqMUQqXvVnzZEOyWRKr2r7w1twVGf8lPZXslUD9v5TagcRPoJ3mJG5f4OE6P
rIcbAwj3tO6Vi4Fz7FLiKT6Yv5501GGkHsa/dWRl4Wrhzd05E4QAtaVtNy1lyaWa
uLUUwNcmxszkYhfCVFKHmr2yj0f4SyBWv0a4KW8AhStvPVWppHOIPruT+pjr/1Jt
+zxdm+mD7zgz48acWuZNG2U/Gyhi733pxS8EVMMebe74Em5Gz50ozTMrA27gUs/I
6PGl1cWoyNXQh/J9DcGCCHvjZIRt7JCOsungf5gFCc+jjxfkLuJRn+oP6GeCjUeV
lMuBCXyLkvs4G2BBHLw6z/N0TlmM16HnGzrW6MKK2S2LPqob4nPethMMOVEQIdmi
fueYRn31zjTgBQLNnacZauDD5UNPf9nAFTD+s8FQypbTJf9fch1dq0tmkXdzyk7T
UZeqldN9DmMsltAummR/41oHOAv7GahWaV4y6M17++EUs0o1lcbMQ1rB+T+V7aoS
YQ7dDthypMt8AlnspoVU5/tmFrt3xewpg0uJap9zymDODALZPdtZIzALf1v4hjdk
gHLSLyTLDX8s/M+DRrdTUJXC/QCaX9sI2fOAcsUpCsZyCfk/ATTT8vS75JaIfpx5
015BpkEB+DlnKqbsLy/qwWs/ktEccdeT3kZgPBQAfc1hpuq430g2wC6cWm38RVNa
lBQpM6YlzHZrTHLLLNwQTAWCWDxPNxZNJhwrX6xoU5Qk5K1YYyo6clLBl4g9ieqA
zvIIvta7FMjGmSBsZxoEzaufFzCaoITae/J7r6tM0oP9dbOZaOM224JW45qbcxod
LcmB1T0EA7rLITfzRGkWqESge7tMdCLtiSEZm5CK0s2yU4SK3lRHw9TzB/H6OYpD
utzBd5Pf51+UAZ7QPM6fBp8yAPZFAtC5mWu7f0VYtojFl3zrCs0+LGlaDsoCOCmj
eud2/+r964UF5VyWFI+gIw+KoeLEAs00DtfBqefd2cYG0JoKZMA22+HEVQqADuld
KmFtkxCLUJJ72/0d3mmFTR/HSxjeBU1v56dOZLfKhL7F5N7MmxdYj60sl7/HZC/A
IM/txeRd4oeo6RQDPHmpo7TpNMAGaHaQMRm316aKhiGRLesCGtz4XnrpECiTjnFF
O1Y8tH4n3QHTxWz8ziiIczcvHwsp9YRv8kmKPy6kVFklM2e8IPo8KDi1LUmFabBN
sHPhiccBwydKFh7WF/OZ/BNYZ4EVKetojg/vR1tllfvWQCmuys4/essWcXhTnlO7
qwmKg4SXPwQ6TsbWxq+5Uza3E+0VvZ1wxYAKp/uVenTv2yWjzWeZhIGyIE2ho4m5
kSeZj8BC168AVe7NehjeC2wvO/QSH+venamD3WeR75ZQRKchFtlro4hriWL45Pht
t0LTlgd76XrSV+2Fwzh+aHplH/mdTNAwMS8Fa5Opz1GDdyKMlB77l4lzOfmeB8b5
djlfQ4uAz3ysvThgp8i02NrTl5T9LI2w8kroyiS3nwgW6Y6tMDIqsmIy760A+gsd
8K1JR29rfxV4dQE4Ua0TXrfIXz8Ic/KDNQmWG5B2eUDztw0np0aY8sep3RZ0RxYI
sWkGthEX4u8RvqdMJKlngs3Xgae0JiW9wSZUaDNSZaCBJ4472RIqH5LOn6uqak7D
tzmTOXtZfo6Gawky7WaVGrrsQMVlMRnG8xZ4OGCoPDKZk5GAhHaClIEOiF+dBU3b
P9bB2xEr/DBVi7d4gpfbRqHwUt/9t8YDgkbi/BY8HlJu97FFaIXTFFnN8N1TP49X
PnQTCgbAjpu/K/vBwaF0rmsssQhsQKuKJs1h+qeZ5j82POK3UzDlm5bYvW5vISRp
k/n61iOD+NcDZkXEDU3zagnH6uHIMm/qrMyj37TLQ1BsnB/W8zq0fPp5ibsukxgm
5yeGdV90oj5DkLTPKaP8A/VRzJu8mVJZbxf+pSsRweT2cTkVjxhSxx9NHvT42PeG
gW21+0cgWH6xYm2qJKQzpdq8MhAF5o5fXhvh6Q8qq/MHlU8MRteDpbp4/5Z4WKBQ
jSTtJD25FQOi7hyrNSpmB0gcOXrLIlxX5TiCh5BtdoIgIW/uAH210Tf1/gBVsLqE
jLoBHVlQxM5UGg23TWGWLyIThucmZEFxSRW2OQ1WgbWqMF90PpGRyrDmM+BUJx0B
gxEVVvdz4RXhdbsRJD3NlDNe7LZtf0rXHL1Qn0fSV1TLmfQTQUfQiIljP3Ka7Ayy
h1Cd/VYu/UY1s7RPGGJzTHaw1D2MIUFb/y2k3KsCP7aeSPGKvHw10ZN1oblwk0a4
kV46SCcClhi7cs2XBv9MiqigrRBFwZ6xMzyFdb+SYe1IKl++L257B9b6YrXSjg+m
eK6wEyP6AbdwSQvVKrIVQ+zQg+GGZFyjtMWerwZOiLv7KXH/g9lnzvLD/AtALQfe
LWuYaSyj95ypj3mJyEC33MWTy6eWi2YkbEKqIre4YISwMNgWtyWm/C1xNnJSaDAK
X+YpWAzg/sbVuHU/VxFT1sfhKgMlawz9RpMJdP/lyMZM7tdmgLvdVbyXukhf5Ere
jJYWNbtqYvVllEGH90RQXLbmSzt49Rrx/rzOC3Phxk1tB4PXt/QRscZWPPR2OejW
d1qPJGF/G44t0ybLu95k2iJxgA/OGVneEwDea+Q+JvhHiTQE0XYAQe001O4A4qeq
MXP50j32uCFjlUzFQAYDlwhWKLNZMVPmhaoIIF3Xuo9vqrX7X7T/a3WEcrkU086X
YOJryStUti9akGDwe8Fioi7Qf9ZwwW78XQmC2NRbhDUXHLBD6fYMuczOyld5PpxH
6oEN8evyCqI2+mbS7LBwS9kG3lGhu8KJQGZai3zR8iwyLeyDwi70R48X2dAuPs78
gjc2u/yCrPiEYSsoReG3t3bBa9NrIlXn8WRsckkLNRSj8yFA0vubHiOXOy6CO2iw
fKKiTQTGlVNPpXn1/QrPFF1/P4kFun+eS3AsEigCu+4oARXkt0qanf08iZzMZvlz
br3Fye6yHmVCmRgaOJKTnlYkD5gpUqtq6+L00bAtZYfee+DnotiExyg2Kap90lG/
CuvGwhVIQpasUDnZjPekUTH6b+0NmjkYHAYowqFdn4kyzzOWOVRE3aMzGFkOf7Qp
nqv/YSLaooXzeZ+D30rXNaEoBt/puNzM02DuLF0C4NUcK09ZTuljqyjUx+hr5Zhx
FbtqUlA/NKzHceK7JnbAH3eLkjyWlbJJtWCbWSUn9xgn3Hg0S568sN+z61O9H3dG
0r1/co1AcH6u0IO+87bDoS66IaLaPiw2u006gH7D2dm2bRQH2uNYzyVa95MHbgbD
u9GbHhFxXrHO4E7sW/u+P1NIvoX068dVF+fOpZkuh4IpQn0LY220ao8PNFWz7z6y
fhhfbmiq5d3agTyKzhzC4moC/RpH9oCo8vGQKPY9k9fTOJsikT39g3F9bJhkUvZW
C2ZAWtQAq1HsCf4zRGjFmIhWGdA5+RaTmYI08CLbI9e1uCXabWNTtFbY1mIDghNv
TYHHI08xN9z1/GEXHS0xL+7jI0SGnRf8dZeydx3hRaoeQmXKkco1HmgkMlyNUW6k
xfU4jhg7pLJ7KayD9ztg7oqguYUGpM+Y7syiaoOXh0CxzczCW+iDsuTPWw2fVwHF
DI2llOqsW2YeiX6RaZWuLVChIDtWADvuyjz+t6nIFiq1t8SkXKYFsdBoMJuWiP4G
EHE39+CfdcKQTMqdFeaDnglQcewSym+wPDcaTIhoXjuY/J18dmp7atK4LSmGE5N7
ZUFzjUh9RtdTVxVEXQsi3EwYiI4Mrme6X3NnNy7TcHeBSHzMA5+TiIp1EKSIuCA3
2zzh4/HhDKActlZIbA0LvI7pTj7xfNDp8GKGaZRFR8NrA3nu1aaU0MzMkCG5io/X
3SQcqEHKG+lRo2hbWEUK5xRO5SyOHNfpfW4dHxSf0dc/cpvM1cg+3k6kvrpgVx06
4dZ2OjFsEdblciOhxORhEZRzwTH2y/86rGZZn5QFt8pHPIkZxL1xePn83T6fq5G0
unpjvTE3Nk5WETuysMPrC0/EFv0TocTMav5qqs7e/QUDBfcVQpztK5CmfyouTlWT
7F32ob0IWqnGB5MC5x1pJ3GXq4gtPZCWecQvEhg7OQl43sedXzAoU08ti/k7YQ/W
JJ5FaaF37DwsjvpxG8QoJkqTWwjsQLSY5RezaG2oTzEsYZSieJgNoc4vtXdDUnwA
pzliSl5tnOGfc3QHTiNH/sJLEQKAet34BxqM3deVqIv2heT2BZiAVQq19Ih/N49f
n1m5oLflTFcaKLtDbTTkDkYUGqYp0rj2MmljLXN0hCDCZtMMXlvDhsY3fpI/qCEk
Um3KwuTRs290zfETd6BAles/OPNW8Ymcrfxhu794roRCo118G0+5ypsusKwHxM7D
zk+T/5gz/Ohru2sFwcSZIYEOrU52DUpnlntX0a5g493bYhX6PMrwH6nZM90EUYXc
Ew5WmYfw8yYgls43+GRQFFLHFwumtHQs4eEiG0kFVkUiq+OjZivIPThLi2wLfcdF
ISS4SvW2v+5+Qk4CLd2P4heA+C6viModAjvJPGjGXxvkTTv6wNrBaDqzvflF7bu0
U3wEaY6K+TJeDnu6vfEmfROlNPy99Ltpo/yJxnrnduDh6N+AqU12Ul+mmlcT/cPJ
5St8NyVE7mXDgHhY4OP5BfM4ayFc36bEGP45zuOeQ/95obnuejrqN7qhdENONfsp
5FHONHi6vBKZn/cTm9a5flKyNgTWnydBv6sEBFWhoPJHDuCdG2wmZDNy9SbBY3+P
7Ey9+jYOWd0IvJfrp2HQ/1kRo/jNfUrg/IU5/CdjC5TtnDxzxDIRmKo7VDWqsl2g
5ii3/ja2uMThDk/IYlOqqOJggqD4pB/qhkiyIpxFCTL633DivvfXt8BBK19x8knv
IizCjW41dzi+cQwKGzy4kzyujRXrGRR5lhA+cwGOmwWnPHWkD6dET0/Z5MVFMDun
3yHultgDRg50mzkzvGg1ZbQ+u8AaEtFBb5cwZ732hUm0k+mcpv29mwNCVu3rZmQa
BZygHDzehUX55pANY8HCQFtPOcN1eB46gXZfQDlcPPGX1+gEV0Ht/HRrm2WSg27u
nRhcZoaESwDC/DCJjw02v1Fx54VL4cWWj6Whr9FUS6NQhNESP0LoX94Y6ImzhjWM
MiJRHMg8YTN5zxJKo2KJA2+q+wckAWt0cLYpQPJgFQpgBHqKEPOfgbwjc664T6Jd
47+u5cQ0nv16obGqjI3hwr4Y+0iseaVkwq23acuZtDaY1l53pUEcqpEe5WYHpdaz
dOxPgp0YA9N2Eeyut5qdGkBiICBFuMjyUia7iIH9mdMdBXK4OsFGInJSF7/+SHIJ
E7Gl30FapkrpBvRg1x2AXWNiZKkuXNe4JfqzBrT9u7Qy8fohgaAXywVm+aiqNqCF
hN81DFJHIihvh+LzsQ1TLkHcB3BBpOFPzVIUTvsr7MrbyDi+obWC/JTyT4EL+68t
GTifeCxEhrDBFf7aJsBhEHYKK/GkuR1RJjQWF9iuzaLCmyghY0QCRCETsqbFGd5w
t0ELS3WS5OL7I5Zb0jHsZXevYGtVZh8ZlUUB3Or+xDbJ3rj2AL9kjxK7fU8wLg4X
5w6y6/e2aaJjfBKJJTpQG09rkSSXfXn60WiN7YG+u8DzhudatZCeYOrCcdx7Ws53
qntG+kqOH4LNiE3ChWCJM3Sg/gRLc0sIRKk3ni2lRD2HC3GYBmmPewfkiPCQDzVB
HwiVq7MoX8Y5WBAMl0SrAl5RyVx5q1qGQeOf7Ek5jDH44t9IRoxW5Etmf0laMnKL
lOYwpioMCc1PQhrJsBEOiwuKtJWBPDlEGTclB23ZHVmNr20/PLPcmrsXP7AMLP/v
lPEXOR8hq8E9PeomNIDmUe6Fw82/oHm7xprB1RLDQerOnR0kecgy5DcHu+4R98ie
93MBdKdMW+OUy0jexubaZXDmcYuMD61W45Ch/8r0xz9/8r+h/EA8/KwmLx1AyYWY
uGPgRyQWdJvYfwNOi+IVqehYjNIpugcq0drlomm6YZq7SdaJIJsEfEDv7TLeY/mA
bF2c1hF+zZw28DF3d73Ou21jv2qrNmLWXYGHkWyEdUugzH0HPzrUPKEZXcToS0Tt
eLm73RT4nGZlYH9p+dQzI1RKJAPBAudjH301zTcj+wEkd8VqLlhOX9L6+tYgxYjc
8YSxRKCuu3BzmGbymaQ+hHcaXpCngBIVBdi446cJbU5iD+KTP8W9K+3q15krTjkQ
yoenZQoGiuuSagRuBubIx1O7tXPg6TTFU/OsQFXPf3MY8bUBAquajJ4/t0f/2sNl
hlm0OOK35uq3pYATVYbSkkqYSwZ/R/uC0C8A55oZEvzfTnmVMEyYAY7pzKY1YBGQ
TWgQyPA+G1vjgmq8YcIvkHJMtRbRvPeB2icaJlEbSOg1h35qe91rkEgFkYn5/ytU
m0lJju+uS7czKMWDN0LJctVKDtkMeG7Iwx9rp0sVCEsp2C3TtzVeMNq9AeLJS71Q
0IUX/1aNVCbG/sIlpvYYBX2a+2w3BBwIBxrHe97XCLRaHynTOaHWHwkggjBiqnGf
eTfrC1PTsR+I+I2OfOgjfxk5797Nphll/8qEkuK6zky5RQ/hQXbX6662DqCCPas9
SHBwiGyoaKelfH9S0XnFyAqkpxo9vUAeQaIVWobbInF721g/RMRmye9xU8suxlNS
UoSLp//W6xsJ9FXTvvV4/Ri/0a/0FRRILYnLJlxCIveDbyKiGkOF1dc4a8EEUDlT
bS+LlvBMPhmSl8TSWsKrlzgqRYEMWM3kQ+f0pb956f45pwfkDMdyD/nw6LABcGhO
g/59PntyzIBAXqxSGwE+h0oTICGDT17jwvdklaSsLlRP8bRmH5vz1ZykzGbYF56I
v1Tm5W5KwgutuQDUOhKP8DfP6p27OSzHhU0xTWcPmrqfn3ADvyB/Y8xwFItB5LXM
lwDrR0fvvmTfNgssiUzObwD6tvWrnkQ0YOhDy4WmJP7G3L4A7Y4O4PUlQdfwLhOz
TQhegO/lL9LmzPpUj1qmV54HLLP8g3zzr8KfFVvHRU2kmXplNbvSzdUf0r/ZgMaB
gaT5/SGDJznTpwJ/XVvzVllJmKe7jc2EI5VEgQxg6COi9/QxPWFTF+w2jsHHZ9AM
CZsS+rn1IHDIPJD6ce80p3LBSdzoR30NkZzEJrgdBcjsQl9ucmVRgayMAabcQ19R
XlG6iI4XKl0nKbOI6eorVz/gWugsYswnyedzcbQfkHBBoDmId2oySEte6mQtTSjU
Ihwgp3I6go4OfTp9gpcjMfKFoWebAcBitWbE8M7tHlwJBhnBjx6jkmPNz3AYrHEG
lbz2Zs4GeHctevJA5GsGhK0G9/k6bmorK/R4swxMB+5ibzRymFs7RRklzJbarJT9
W6hu3ID4HA5bBfL4AMsMCOkYqNzpPX9BjbiHovdokR0As2UPI2Tz7I47asYW+ZCW
F26TuNYbpvCFLE45ZYSg6W94sXY06OL61OmfjJypeVJtLd5ktHBd5VVBi+/cml1H
gRMW5ajPUQ+cFumqFVKh0138m50vHSTATRzMteeos5VrPCzGx7HbxOu+knXZm7Sc
y5EhWiiIyHNQeBD++UjEz0kz0xqUqxicRJu3LAyKxF5frlRH5SwOZgRNYKnh5/Wi
UA7rcy3OwoWQ72nKonQkRo0ziq0g0cpy5Wy/c+o0Tlye8XtuLV0MX1GAosf4sdlg
3oxdliwj0wM0l0zDMp2b2Y1+sy0GW6znOVSkbGCbMJu9cbPTHagEiG7uqmdnAU39
c4gAVfsDcLu2Tsznt/Z9IhBo29Iw7yD1Lc4xtRNN+QGv0I5lRvVfSxWBXli+K023
5Pq12oCEWZq3KNSONIbvOB+n006YH3WLejqvDgDasDnYtk31juPfng6a31YtsTIf
rxMW9iL38+i0Zwno8hVZuW7TrORXovn0rBzQpW5aqL+QQFDMz5v7t/MruPfTv+T/
Ln2cm4fRXcpD8qhRycyOLRybxb9ZfzjqDXawcPM02X1eku5pBoZWHVGExA4vGsae
qcLpX4sr85j53MNo3fc4f3z04HELdNJcQ+zpWANN8c3Cc/Eo54xpZr3C4ekdiigu
BX0WXAoAbonCLkBx9PR7FugNrYLI0Ldh/INXNrFLEqCAQeEVmVS1nJu5gmxvJCAH
jRiut0TSROzx2AV8bpjA16Zt39IoVZso70TXg2M8Svsa00Gw5DI/0vpFzOU8ozVG
53CLbI3+ayLesssk0T4+Iay1lfSU5/JctwiqHv0juZF0jpOcehD/TWQxj6Den4PQ
BgpSIy0sNtLOt7PCLveUiqCI0cQs3x3FjVOMmdFSTRJYkbJmO1+RMRYQwfRu7oSN
nH1U6v8eZvYwWbkXEU0GvvkQg5DQlKuGhzmXjry986I48QhVY+h+HobLYt5xTH2o
jPfqXa9z4jk1AF3IREJztj3Ewh7I2R69MODPx9PKDlIHqh1PznjxItV/PDkqIzP9
muWiBh0jIcQrmL/XV+VZb8Erb/gYTr6DEUBO1HvRB+uk19nN5NdfDifrO9PVAmwm
ZZEb4FVbTwjs32PAEbrjyfZdLBKou7w7/+scknp2n0KagdJ+vhdzWEv+/x8bxwaV
MdhK4HMt8FNSaVjDs9xBoP/F0Ph2fyJfCNmnynS0eZYgwqtVOdChRUZx0ccEXuob
3bcLMiJySkDh5cMs3/W9q//95K3XSKRnXrRGla4SgyaunfJiHREmcVShfQAjS2xc
wRvf9bCI2injrFDKUNmPrHIlHB4tRLmWqRMFAnb71HvfgUq9iT+Xso0lF2sxA4Sb
sDpurYExu3L7s0JHtWGKClEm8bE3coIlhEKMICI8eGb1P4e34kCyUHxGoD1yRvzl
L6EZk7P1NetVSAFuuyoyVgafnZ/CZNEdteQai+m67M3QQavAKlraGCfWKqOtmf+V
qZZowweum8dIMMEZ+GYHvzeSnNLnIhjJIKDxBc5dezwJsPY+IJhWYzELd/nnSQmF
U3/G7wibPHdyYCsGpE4u8r9oIYKZWFi6xgiafzm38Xf2YBT9WGw5cuaVIeC2jBep
FtQA0C6cvswzGbghZ+IjU0Xx3Ljo8ezm0L9uKQ451rkt0pkSfjAo1PdtCfocNbuh
udWrWLII9KLx/Xe2xQuLzOyWFa5twOtJNvVJKFgsTK7yMhqgRsEMpQ07oEXgsBBA
WQUUteR9VBsnSAUuQy2hA9x+4dviMMfPwv3nKbpabbS5bxTps2dtMNyMIkjmvVYx
TKf98WW3Xn9hHwhnmZ2pplJ4an1xh2R6oIboxg/ng3Ew/6oX492n/R98/IDL8w51
ldBO3w8QfGpXcEVgFfs4EB7osVy3YGNSX42iTwcgEMURM+j60+6pboOxiGHh3bIK
k3okwBr3g+GcXomNwDG0TVnjD4slysIMS+42CZx6GGjZUL7uCSLI8LE9sDF6OB5k
gd/pWamVAnl78A2bXUxh6DG2s48PCeNTM9cM0cV6CwbQMG2GJhyHF2T5Gu1Pwuma
sIK+zVn4izuaAV96NfjTdY6jm6JqyBOdQqewSFcFQCaExGIDBr555o+19ByDjxT8
ktrmiSFj1K9NbQPYEQkEoacYfd3MVaFQjnJQA86pAc1RpX40i1zSXChJDSOgbmIn
b8UST4G/1LEZT6rq2D6vXppKlAX3YNKj5i8S4WGkOILt7OTKkPFqJ94DGjb5PieI
Ie8wl38SWhmRugH44SPA3oyAacsNrYkbQwxSjRnVsnrOt3Gbzcd2bGi0kychtWGn
4etu+nMSz4/ed2uQeeBfOCyWM9HJUn9d8lXytHkCoDejyPQOE587Ju6ieL6P7QgW
o5hB8UvUvOQ9o/psIcIRo1Nob1e7c8X21fmk3+YRCUz0lWWrx1SXAyb12jVSGkjX
YDwQYUZNz9+Ip2qj6OGUXArQH03gPLe/FGZeVWC9t1sKStdLEi5l4PYK1WmTbzbB
mGRcV1TlWJ+ocuE0BkC16T7Gssyuzw3AzcB+5w8/PAyE7TKk9cf52ludrS/aZKxh
OkzwujvwFNqJZhX4P7i2ixvRkFGYo4tVmhuSlSOcQpMAtwZ+43GdG+sAvd3HCVzx
hfEY5LyujCQ2knJpV43cjNa8IWyG0O/FaBo7K2VTzHUM3vTyMUVyZeYPCHQyR17X
lYqfdhL01RDD/RTYA2dA4oEqItiwkh2YRj9uoe/3rVYg+RFSywZQKjWms2Qp9U8d
sZeNWktlXcbzb92q8uYK/x1mDYLWzs2UebPYogR0kLfln0aFcR6HFjEvGz0TQn5u
M3HY8PZbEYUQ1ePTYqJUch+miX/yQm4L4VSNcPWZELG7PEHvoFd1/m0YmtSZwp7f
95Y0lABjBNP37Mh5+I3gcJA3mXcaUXPCcTBGTjsm345Z6d0NVCHq5nZZuwyMw5bQ
3H9wupy6qryMJFJKFSg5M0AEqjckvtdGCGuGyEJQsu2Lse9g7KMUJBirV2BE7e7Q
0O4Om4Dysn4y8QfjY/VYxJkVe75A1FFlBa9ZqQcEZt2u1AYiT184XD5CNyxkpnwr
n8K1DqpXU2d/40nTz1cr5dMtON2gWd26CW3d3sKLFNeV8v89B5kspTBhGLcE26rl
oAeTo5+5rYoGdAwediEJO5XjhMBUckCUOHPr7U47nhR2t6XzBnkfMSHQeS1QAPWZ
aGmVpGB4n6W8m2pMcgSrrdL2JYmA01DuAqVOSgHOIRNHs9RsoSt68H7UUsYIfSQP
Cmg0z9ynRHBvlfeDOL9TMoAWTcSDhZgBYNoG89vTT2vSj8p6IlckrxRGczJ6FwN6
PYqVLhwrbNuNXKWPO395JSmz/VaCIB19/XE5Q63M1JNLY4lwCM0mjxh5N5ioKVqO
AaoqelubwGbZgyVSjdi/Ef5t7fj+FWL7d8EwWPTpMczRvTbQMAFEkA943/CdYULV
ab/Y0U3VuNz4V3wx9WUmIo+NhkelgNwhSaFQH/sn8wcHYafjjl/xRqU7HMwMqrON
mdeyVzpJ4aM0pc3Y15BcJ7IcN4M1F9xAGCx1OXUGdCoex9yEyvVbP0BrQaKwtIJh
YkNSQ7XnyW+LTEaMaZLmibsYa+D3oARSEKCxcDcFoRmvQN8uK7ru5k7gSnva93z9
x2EXOHVM0xM43KgK7rDF2OEt+IhnwDBJetLAmW08wUGNMIfeVStuqcnagNwt+IdU
4RVrtNanVBrLHJBcJSgVpc5laqfW4DJboS1D3zV85LhXb67DY8gyFgc7zAhZeHgK
ScBQJ2kPgxT4c6WESbaWYT3tKJZE4TSJAVEH8oalN/2ZVucLtTaRa0iSfSPYRTq+
YI0I7jhLsmllYGnILNAW0I/HV+IyIYiq/ylQkk91r1LHeyaiDYs7iQpyL6BWcWsE
kDr9VzxdAFelnRIyKSWYaatKdleSmyzKknDgDu5SDxudM+e4gQh8yaeJj/K8/MTI
PH6C6CDDeHGUKK11NwuiijwkP6rVBDPWqyRvZLwgtS33PBIs9R5L7kkdqtOKnTR1
6G9lmJamVpkJgrGSuVTXdQOnImiy7ID7DATUTbfB6lDty6WPFdEyG2sORC2qSOpA
NWkY+hh+gMf7mX+4dTMKhGi8SaSTZK5qhkyEVj4DsWFcqJ86yxD3FRmtGmdqRx+0
vhYQ3lzMBa9iQ/eLKWZ50bmr3WD0cP/J6Wkpo9kg8wtwLfAi8ExzkqLbwmXqoE/b
zqUXrhWqeO4E9IBdfRHta33IjvmGA/eqi+eXK6CISqh3mA/Dzaqn4IEY+tA4tLMW
XBLb+UFMVnnIq0JiC0EVsNq4r+ULcr82IbTep/lRyqPYys9+nopW0uhPpElrxfMc
mhZJu+W2A88UVSU9FqGKGbS7K9BvLd/WhtP7PHExDeUNs5Y5xDlFgnQBRGxkaOpc
uwxgFObhe5Q+SYkoVKfDJ8D6LXMOn2DhsZALtDfQkJZ6FcSCv1RN3oK14na9a+lv
j8E64epuk6vDoDt2Mjx20QKesgqSosEHNNLcXvh2R6GMsqVE9UdN4DEgYZII0JqD
pS2cf8iTLgDU9Qa6Xp7GHNgfIwOpF1PK3LoqOFXW7EXso2IZ46jyIjhdHvLrx9IU
DyLnww3kUChnl1IDLA3fs+ingbNiUOWcWdKtwckV0khLa2p/8TpVm/Ed4eqwgzCL
Ih/A9t8kgwC1NS4Sxc3OR1+xgJorpQG5sH4NJZZrOllneNbgn1EaWOwxWboE31VU
ar7Q7NzlFiQgt9WYlNTteJbLiQpaW64jbM3e5OeRD/wEXVBTwvcYISB5QxuFByne
6ATQrAvgc0tKfb1TmXkgfhc3yutpQ0E4fEJD6IQYIc1n4M0CEdVvBTnR1q8Y1Pem
NcoWVKwEB1Xsa1UgRLEkpmuyZpwhofsHPvUSoIYZnOQ9be786GAipDRJDLqGXdzq
VmU2+YCQraR1sUq3QcaxmUa0FzgrP4oQNIkNR19sJDejpTN/lI400/xAnMPeULhy
xTMy4HlYrVrJWiENH0Z/JLgobC+nwN3RJ3KAIwHmnTwJhQ7VhXCbAdJpIDwBYO4q
MJolk0AsW791Kx6he0PAr2OnnhymWDdsSWJYaGqgFn2Oyf5iNPgN/JcbO69/l27z
+WbhYm8KlumeC8MDNJIVSdXpSpYhych6R0Znit8o3TV4EKZWgbkVQ12qCQTU7wTe
GSyXhlWu97SLRH9SFHjzpwwIqfeZ/aMgMKfH1ewuK1yoyZ5dZNJIGfLQ40hXpy7q
vLotLb8bVC5GOQHAsbjHfXeOhBPHlE3XJ2Lx1HAFjzqf4W3tDuY2IUOoqNerOc2w
KEGyZLsCL3iYvYl9w/fkCyDg9ZKS2iag+yk8yStH8ebgeOLZrhIfQf3MOKr/Plks
pCbT/fdx14+NJB92G6TvSIdJKWGYLg3opWtWWotqWDUjXIzXSABOENOWoJDHIU3G
U3Ea1IofZu9WrqLHrhnatn7tIAwNro5BeMAdRqSEDifU5l2TN651VVymXywuOaWe
3kbrwmDymolix1LqKppqZpJHqbKA6cYgqsNJOFtku2lBacoC8PJ2e6FlczzRVkiE
XtxV1LK83bU11sQa6d9/lmfFiif/P/c7SuGPwfh66Hg/jzAIrChH64lewqZz01w+
xoLh5xEECpswOZDVa5dg2k9PapiNHPbjFflC84Ge8HTnJABQUPE6ywdbC3Z8wVNy
shy2SHPd48mteSmKwGTRioxSQ9SFiTzVNuURLRAQYgsTYd8isGhz9L7OtI7kDA8n
tzmEzBcOr0wwkw0vHxqRwQv/VcQPDNL95ecFGpwTcMqkhcBtwHXG7KjJZVSJ65c2
mNZvDJjQ9Clo0/qG8W9g6R7HgBNDfWaXKKnl72QjeUUCWgfHZe/ZhDxu4CkCNiaw
U2Cs5wFDHNXkvY5Lh5Iq3IJ32vaAi9hScnle6V6NPCiNLMeCA2GaSjWjhgGVDOQr
ge1csZwIt/2eSQHauNJ+wWdTfkwvRTLl2hNILa0Ic6FtjsgNJ0MYXwRGv2/SJb7K
ns2dEH1CxosxPHvcOqec9pCabt5YIXNCRAPjC1rDXb3y3hsLo7OVa4Ukqb0AFrdz
JjFkUUQeNm5BRAgyQnqDoYA3RuZjeqelVlP5kdoEkinE6seS7jgILi8LWdp4RMQB
3I1CejDIR4HVt7j5EvbOwKF9w9BsC0XrKaGvCJ2F1yQqLYMdZjy81XdGtLRsIri/
wTyRZUkVeNxdNQXD1a69B/b+dMPkrkEi0kdtp86avD5tFxUwRbUxVD92liC//a68
WlSjR4U630q8s6VX5QoOPeQUKAxmER716bdNnJrM+LpYpu90371ZJhtF2IqHYH/a
8DsBBmAa5+4f45dPrOGaGfjs89jaINB1BlB3EgeUYs1TKfvlbolgdhddbWg/WOp8
03Wmh9fGhtChAIttz9ehLRjMm6CJufaYQIPfix2XvTXG8vCPNoywQFgzESXedqa8
y7Tz/5fVrQuWq78R8bFSzuqCRfMTGyqR2xZCbi0BRvJoZ8ubhdAwbbKQ5Y8u5NQ6
Y6FTwMli4PEB5FTqdy7o/aUFCWjzoKOIGl4crp+LH6jUT4PWjUJ+DI9deWj1ABLt
88v0Q7cCDrDBt68x/lsNv2OmSkhfDFyoeaXA7PxgOvoR40q1E5KGjFnQP6XZSsxM
DWg8QnQFzQzxKKppqohhG7REL5YZAGrvsqal721xOf9E0VfXfS4iICxtrZQpm5bz
4lUmCxqnWfixjvoQneU7KSqVg3xm7JrtFzhB7Ef4/zbVFqRQuTCC6Vqk/hycn/uT
AXLr931d/1z4UjwznFY1Xm4LDxTZjHJ+k/kE3N/6hx2e0utKl/FuD/e2e0ZkNePe
Lo7il6gqBQtlcMdVVfryJHD7BsYWV/gBiaCbfr36Uog7iibgu55H6GtRxs5ArIVF
NReV4q69333g7XhhXZ3WSayNYuESTGCq887mqZDG6iyVec7//M+D4y5bbeNH/3X3
HZdIQj2lM0FCZYtceRzXj7J9KQs4H5Q7jeFdM4wsLm7WtF81kTtw2CFSuzJc2QsH
qBzbVHBIjKWj8eDEf6gytCC0X3eyjliM0J8ytx6TBQXzcysz2GnkNz9VSvH3/qLa
fdETPWDG4WTHt+iLMA7BgIOCAhCgA0uXjKcn/TUi7gZFGAyFhiLcs57wUmrWEqXI
1vrpn+y7XWmsFbk/jGpbarUaJgbUfe53ZkkVyxY3aA+/G86ceqmhSvSyK3h1Ugoz
fXi320WcFqYxB2+OJIXAitAF8FPvYmOZdw240wlwHDHXT0HLMpHeTBCbrxMuxPH+
oh3I0S2Snel4/uFXlJaSo2nU1LLggexa4F/gUpfWSlplu/Hje0soyjoXtWrjUc44
Xb8f3qTUALWiVaep8wFb398O2jdG8pkoG/BmPa+fq+kRchWrN1lvAgzlNXeMT4RL
iluHkjeDiydgIUrLJ7vUM9neU3eKvWTtSQBLluAA/fNvOeZa2/ItYxJJGXINxDt8
jxJoQBG0fEYsho8NrAbS3teYbxFTILBrBrspEWgcVJH343uxoloH6D5orhTOiFyd
nBA683BI7OjIgR6yQGAo7qi4WtiuPt5RkNHzAb5tc+Hy9x7UHuN7hHgowYuf79tK
r6SykgH5aMM4a+qLRLL0xzCfRswhnCRjnU/Ia/BQu742dE+n3t3aNzqqm1U0s4ee
c7aAcpeYCjQTf/RAI9LbT64M4ZHrGBIgIKZ0KS0r1HZEYfBsIA1ZE5ajUbA5mQ27
MIEAOAZxk+NyAeNd9pkDA0NMyTOlGfuFAvOZ+MQP4hCZeKdm0XbL3ERDB2xVWJcO
S2dMeikDDTONoJ2jnbqCPmmbBMxiRYTCqtiWhxR9QD32iNwChxD+8B5DTA6FtlKZ
eqFr7wkUczBwG2xd+8NsG1tnCuSYtjXFeXuqDykt4ZP6+vEodcSIH8zmzAmFK4Or
O/aPJsYY0+xqaSYvhXRH43f7iqtR13qQdCnt57MelxqYF2YeM3gGKYP3qskDQL0W
L2l9zwZ1yptR5o3vQIiVlVAKgIqWJDjlTEB9JIiycvmC1gnJWwHAH6dh3iAtVXcA
w9Gf286x41JHMiqypEh+km+MgLReedS5MuIUSSeJI5ZYGQtuBZSyeOOsPEeOmVBJ
Bmvm+jT7Mo4SckPBjVxF3pDe2spWtjZfBQy8/GrGk2QHcqdG9O2HMiz35fVLmn8e
zzriskz5fZQMaSU2RUSQ9akLTEh8ArUD/Uc+OtJkzqiAuLwpSjqqFIKgWCFHJdno
Buje4cdMwpWg05TqTqvLWhObJ7AX9KH2Pgm20arSTX8E2lwGxgCqljhi4Y02Psbp
zFIkaZi7oNIpyz0aV7qcM1+Sfiy38mF74bWiQ+sJ30nNDo3UHLsFPpOtHNS8HumW
kBaaXOqgPRIFDLd51w9kSHYur/eYmcYcTp/Hxo4gp949OB1UHAhK871gTWzYZocd
yYIrB1pEkz7n3YyKQmNc7tHfk/7/YR8P3c89cgRHnPrQzwViZfHKsnHI1RLsxeUR
qMXx585ZBwhMXiFsLQLbyrE/NSvavgU2UxFxPi1Rw0WeDZHb0jq78hWCqAOJlI+7
Bd8wWLRlUcsvuoU+2PAyGkxbuO/6jun8bNVACUMYBDCbTMFgmhMVZUoukoapaYhR
0x0xOvVGY+lqlp7je5SnVA68FwNnAr1temyg8BTPwMWwUu7455CLk4C23JlSVCND
fvZqmRF1lFOdu79CeX2cupwtGwcgvq9y11O3yrpu7R9MJT7g8Qsgj5u/171L8jZv
Kn7otgSNY+Ro11XKwXvsViTLADl+rxDwgy6bWqWePHn5NqTFfXXfsHSRudnhLhIv
6UjMmhiIWvaX/4VArH0JLZU7ube/FnGGMFa6uKjJ7nOuC3AoAB0sn4F9+6s4uQ4H
PfycOUo942RFrSyQ+VtlZrrvSu4rtntuaTJDIDlIzWjcQU9ujkA8rfx7TMtvFaEp
Y2FhfwG7x6sICE/4BzJqLogVdWje4IO2VqAQ5rFKHlXVWIXC+vEBU4lbxVv1211O
pMLxYHezDSabOGEVGlUQnjTKoBMprYDBSYkZpodGyJnfXJo5EumceEr8dWyv+TCk
LOWINSUVhFuaVnQhxX7zSx0D+0v06JPec1A/6kEVv5GfxSOr+Jt5HMe9vvqVDPwH
bHHKXWtITMQIPWDiaXnBl5ugAfsZNKICuVXBUCTxD0y7os73hGTX27DUCjPEZiTM
PH9atguxzXXrW6D3vbm5TKV+EZjWmnQgrIn7Ej5M4WX0P81kpO0gs8tSABiGxQvq
W8rB2QOIksZUTMXexxRyEmkCJka4Fui/WhIrbDSGslzMzTB7wsfjMUZ5Sge/T9dR
vvHMSwJkSiAWPMj5gbUuKFmBYPAs8JZgIp86X9Np5wOl2tHZtbUYKexHHVFziJhy
wb/RgMyy4T8W63qL8ZRgWq+oOW7yp10StT6wmtZeABqhK3cWDK47WJ4qMl1bmvGO
yvuCHqnbGXyT5PUNDTskZYgFHWHhnxu5+9UwUMGNUx86Rj9/8JYF739RX9IxnfSf
xZEzlGn6WRWoIMS6H/6Hdnanb0IKMwzWPqLETT1yhdw1sYOxFeGWyPT5OZDQs9dy
rT0Tztdg/wXyPnI+U/8EEe9d8dgtxHKFwdiHunrdFFs1w0LN6q9BFNYzHQMp1mrk
i1O3oWlbEh4F0PzJrzJjbyQZLoKrQxck7ZoCmLTcKaG4mDCVuengumApb9/U+qHC
L3JAnA4zuTqeAC8KArFoMmd4rdpLDbGSGo4zMdAObIrhEpRbZQtQwxw2TVJDAHCm
RerIsC/FpgG3Y/rRl5nyIX/fEXGvjuEBiE/pdsTKydPcMvAPOT10wOPzXL6SKMaG
aHsdLaZcs8rqh/tF+aF8J+Z2lxsN1Lnz+D2E7QejO2wgi1WCNBqRx6RndrUB4xWP
Iq6JF31Ajo06+hSw+/90yJEhbjMdKYhFMDZuwOQDLS/KkbYkUkMRL6hzSG8qFjmf
MVJV45mBCRpDiFmjcLgTrSvJ6UznBVS5WT9O3qxli5JZ5mEOIVShvL1jV56pxaq2
ijxGQyUjbz0OXk+sobbxNUFu8NSlCWUnqjd57S3MoWI37M2Y47cEAzbHscE2WTEi
u66Y8E/vJC8eFl/J02EPUe2NxLDzzzhVWcfwO6wsfLr0dzGU80q0phcVTT7g0nj8
YUAQ50E1La+xz2EgCg1UlxA0eWFDS5yd+s+jv4msi5ua4Og/Zhb8MgFRCNqzuEq9
+9mdmTFPzBBf6HgzQZzXSCzmhZQHQrQTJgo14RGzhHZ8+EcisZwF/bZ5GFf2FcEE
bO70sReIR9ulWzj9kYOuqnBL+roObPm547dwc/yj+etvNJlZ7JYfz74xyHPKsocK
lR5Ky1BQZ/WT3BkrLB8R94s7Z/qFTUFf8A3LcKWN7SkUfRGIWiwf9jgos+qLJqtZ
aNxtTG7byxtBEMDnaz4cPBwBhUv8kTk3QIofcS6pTWHQr5UOf5SjrBsxsHEiIqco
yXnis17GuIiVmhqC0Jv4ziN+0Hh9tyail4pJwtngXp6EPmXVAcqZb9vbi/s6W6cg
SV1lEkrbQVzQ9nfqE4Kr+W+F+BsoNKScWSCzn3fP2HAHnrX8ov2nqgHsrInrzPWn
8IQ43c5uiMOI3SJ8av7c0xfWydvRlqBKV7ZbtZo5ZjObWkyk1KcZXXGHPUr/Vz27
ZRO+kGCOjAbccQfviZBWtN2dhWrkG/Q4qJ7pNMbvv45sD3q9oppEzFcXtD/15fBT
XKqPvG21q7Jb3VKKITqBKprXA7qFo3c/LIlj+tRQLzNSHo9nA7aafZ9+N8SGQBzG
xBAMNzU2Dt8ngNjta22Zfl+xGH9TO2lGA2wsHem+1ELaDaQ1OgjhlAu8GNpvxYB+
ESqrcGwjoyfzeXK+yZqrwVpAvmbrFr4OPgU6evegd/61w+Fpu0oX3ttg+QwCGNa9
4rlpWkNY5zBzT9v7tg6Xa7eKIr18waUa9AE2LNMu/JxxNmhaqB0f4CXGODZWyq4W
O4qRXfgnshdOeqUNlIGKNmDQ21GLxO0W1S1cwHfIl39rWJw/Ul0I4jw+1eXa7ybk
OsEz9icF9ISclrPkql6lYAQKpnokY8/1CNM3dhQNIxwZ0rbsScHtGYW6nSbcnpMu
vk6XwSc+o2sj3iJF8EbEEseOTHOLb+IhoPK98o0I3QbEmmkM0OTNF+dR3ERnVS4Y
LdjYjPB9N60tOUoI7gRdKLWchWeE35DbDiBG2TLYe0icmYz2txgC522CTN/JNNph
M8cFYlDFY5M4RAPI2VoJaWTxTYGrB90y7MdP9oZXu3o3XZVNcuVYyHU9Z5HxX0Hd
0kgkFz5et/Pp9YT0o5yQlmli0W1qD7DPqLHcoUyWcpuOGLIAjxERxsIFnGEaMpJ1
0cFA/Pdi9+qs0PF6VG6gk8Ypo44ELRDW3buQdlJgu/TgE+L5zqJnQlFq/nxTTR79
prRVm3xs672yxbFNqtVBJV5t8LgB4VpAfy/m1hLfBnT2fHSfEjRJZ5cEFr24rQ8S
1Ec3K+oTmhvOBYNJVZKPSZw6G5w6AFkyjlc9i9YTO7HEqoz2P3KfiKcKLLHyoPYe
DjPEjDAV3HSHsGoqxRujch8ejpaZBbvMsT4YaHhlFYPH6meL9HZECv8kge3a4AKv
8/CbRpKk4cAcuPca1rtyRy8ODd+beAtNAcCPnDzRZliZoo1torHzis4RGsf6v2hY
DfDk8sarN9HXPxoQoA9qYUqmjnmVBWTHxZVrbvX5ZRmuXxGgI3IVinwylANve781
SdliUixY/NPzdptF/6DQbqN9adhf/U0UxYB/KJWLZ2VmZhQXtwGdyQp2VwXcsdQ8
tUdC6G+2mdPLIk4TuPj8QfrYL1nXNeUFVogrbeR4/RmYzGUJpRxOC63QEC7V5fUe
YLTeHeTNwdG4/ZDlFg903HAd8vvSpX+LbM0G+S+fssNVO4wKA0myKYybNiCT1zQj
VJflNbe1a3yNV/0t6vC3AptLa2KBaNlpWp1hi5duU7DSSa9IUUCGfhFTpwD+/imZ
E1chWmA6qaPYfYANAhluwOcBkkHV3PhjCIWQnKW4AHn1ICBuSRjlUZfIjQ9wukR8
oEIWSh68iQY6SS1yPDDS1n7bm4Dyy//mOsPlFEK+UXUp6Ijetx290d5FzvMRoWZV
opsnvq//LWIDQYv/IlETeY7yZz5qtgF1Z2E6WkO71ms37sWDa+TQrJr0ly2WQ5Mc
Oh9GTKEA2RfM4FXurqaqInU+5qD7/wrgaSAR8ofTxn3eOuYzKZGyOmctbzT3qKyZ
NXTaPgNdUc+dQjZWaJjMYndqQ0yM4UVHBb5Kh5cbUW+hE0G5CpZa5PRuOv/5fwka
owi5iVhqqug4nNuLVliFuLFOIZHQhPZgBeaBak+GVV2gkR3CyTaRaJPFBBz8h27X
XMhFRBDNvq8ipPfUM46kQ6InaQ1BzU15mjJsTQW/uLAiigCYrZx4pUJ7GU9XIhdv
ne/wzallBs09v/cJwyjtmqwqLQ0wovhkTvy+G949ufTbBNwJ/WmkVbKXcmQHMo0B
59nSIJu74eOrthvwaFlrCnZoEDVQ7uHWkZGBi9Xb2DVX/pgduBMNdTvaJhaOSfZ2
iGZWW4TT2y99vOmqjyM3EX+dSs4jm2w/Iu82g2YbiZk+0paL5kGg+LPcoNDnbYXN
dFoPfqC1mBbEDy2A7eLGmMsnbiF9vmQT+nUJEqzvKnNN/txat1epbWjOiklYKNat
Cg14GOj2rs8oFSYGToF+dmMY0pBqM/zj/SO/U4fnsjJXbaew5X4H4Wu66+nqrVhy
DYEehJYsgaVgWBP/G5vyD/yudo97uTQykkqcE6oXMZyFdvhUcxX7LCgvk6dV2A/g
qgP20VagWELksvsaQ8+E5fHM7I07sX0CO0MVQ8tnbIorsmhKOkXU320T9LSo0znM
HfZ0m3Bb+lZDzHSIAfTWoTesVWeC0W7jUy4foXEaInmu70X+rXHFdKewYb3VJBeI
HaYZWGq1va92BQj4E3quYfrGyRDxCikWa5q+SNE8kkFTBUm3aAQVLn5xtJ5UdC6o
R+1A2h6VUmQSpiKkPUp5X0whOALCaSwy4wo1AMufKSv4X8eTNfAaQ+KVZ6rjqZyh
KBk9XDaoLTf8Vw0z1QMnH4MHAp6MjKwsWd707eU9QjZ+NN0bCzUBFLiq6KnjK2Sn
eCEqx3Ig7Sglon794IV1p3YMjhTPbnx0QWvO4Mc2Nl05mOrVytkXKA5cfH9svjNJ
ys9lbrwPJf6HS/jIMSWyEbjR0qadgk0Kd8YZ/eibWzuHxbWgyfogwQUO0V4sfK1Q
snqpdiBjnj5UkAgX37nL9kRtgXHaad5vd3MSpqyhv5oiB57B+GhQ4VRuAe0Llf63
6Vwza9RvjefjN6Y+mUioz9l3hC63WN4Eu697FJBzGW60fJWJln9asIwZs54sKX+c
8GAWxXSlYqAq2V2cSOVhmF24a5t/7qXm6rpAmPMigKn8QWt+NzxwGTTRUB7+ic1c
2g+ssBpEYH6y/44YPEA5LAiqOb3E99Gm0EGMqErkk9aPsmeuntSULa4EQRVeFjwQ
pI2h56/ehupNtbPWqwXkuC8ZxLHed7PH1wAUetZAZp8/9AtOC1o8enQmaoxBHmD3
VeXF6GaDCvTcFwIPrajl1EKwDtVjGngEvID/tUX4FtzO9k+TJr7GmD7lR07vQQKa
bLajNdRbw2Grl7rosOHABw+YWroIfOg2dth7UMupqM3feiX7yPrgxAtmYru6PU6/
OqdHfDzI/6+9FiVfOJZPRgzXHwaBgof1nI3VjqrhEcrtbc8r/cABWtsnHDKnrJmM
D0RZHrwxI2QXomRYSk3OwICZlFaadeYZTLak/uSbsT9AJqyE5sheqYSEuQl0ysHw
R2LaDmj+3UZLmH+Li4TvUla3JwHBN6+4wrmvHd4vHIS0W4QLXqYF4kr7aJRx/TwH
qiCjJYl+5jYmtLiG9pHUseAWWKhmqFFYOwWp/cyGnT7Q8ha0szj5sCrLZTdqzpI7
qHp5RyzuUrV2g96r/2D58dtd2QcmA+lHGIXFV47r5SFab56qY9uHZjGQDxubniBy
u2FQPjUkw7R8PAt5ecvYCLIyMygz3e7iMVjHkYVAIMl79rl43ZRaiRSZXcxmOYtd
y0ffsBadml7BB31R9+DMv0o+1/QHsmNIe4du9vNFbXimfftqsomfBZAiZ33Qq9xn
nC6jv0kJHGGZIQQR9vmRte49hSL1eOxAcZf1S0tdm/BCFmRcoCKu/dksEAv/1IYq
NvVkexJUSZr5v78nrzVHaO770QVmxXaAR6ke1Qio8J3r7i3FOtXYTrgFC9E9Y3Xd
WTVZ4rb9JTUjH+7aEC2uWSKYH6T9JyR9CweYD7PPThQylIkAqCoXR5oJ7Xw4GZdm
Q2avITSL5pz/JDJs2w3QVzp8t2xUE1yiS4m8F7zwtwz5P1O4vUdlGmCKinOSW0Bv
HuSzhW49WJX8k/fVLq/oNtZgV9WbYj9vcnmjYqHOPPWAtCoDBBQvsq5PiUXESarW
AU7t73PIKkbaTZFzT0moG47z6L5P7XXSiDOt9jqfk6VjPgEuT2sQe1cF62R4cnyE
CVKnsDxWvUTljzo5HzajEsL/QiJtG25i28xMIdVtUsGr78BFnEKTUG2XU9nlRi9j
ojEACDCWR3Jidp5peuxw2cne9IyPK85dV0OrlvbiDUe4Q9uLGPxNRKeNKCBYkr3S
0A37feNUwux21hsTNZi5mnwPWE0wP5KosOPoYEHOl6bVbuoGZB+HtI/XuKxElL+J
aGw/jL/2F2JA/LGcpSMFHGWD1AxaPHAmEWmlkupzksukHH7VyZ1eRDtEV6Qw4LtP
5hiMmDbRjHjgYRlMWol2IvwSB+xp2SGKlv80jMstY/zgR51mrNtREomxKUpZw2O3
t6krlGB5/zyfhv1T7ocXgcnizxwH5tmjoDrbRmd0G2PAX3B4cNT6hfp8gl5UqCwn
8A/PxFjRwnqStPJbvVrC3+F2eVkQyTWmaLHvgbtQqH/GZPzyIugp4F3IYdugECwV
LmAh+nxYvbH5D4xLASlJBU39ZeX7FBt1zZoazlb2m01vTUtKbw/JIv9/AHhFqOLa
MP+72HLCzvGuC5lDtUMf9yFb8PsLQH+LTpy66AZTnQw0aAX7gFZW8iOctDWKX1Id
HNqgulqCB4XzQAFSVJHVN7xUqHekkmMbe0Wsh4jdpzm0eZ8FDfd3JozE5x6D73Ib
g4lxraWhRiAA+Emthpd8vnQu/M/eRwUolqutF903EzqB3skjqXWTiI4p9KWisTRZ
82BOCSe9vg89rQsmgjI8iQSMzDV8f/SbYaDUziuDisxSx+y6xJZvyQUksTZcsh6N
EWbMBuJLZtLwTdYRtjuCzLqFNrqz1Fv2DzOHl3ZZSHaOVa25zGwdkxQc0gYR5jeu
cneGr8OIx/Jks4mwLsRFiseVdTo365NT/uyeuyIvduieC58EMeYlKNx7/eUkKZDW
d4etdkrMCrT5/YYHSqUOgAd0BPMGJ9duvCghC5uIN8tz0H1W96m+L7rD4+/UQdww
2cEbDy5TdRkM+X8moKJWOBX4yN7R4ncGvsS/I3UTZXSLHA4c55RsuTiA++JRnIko
FDawimQVjmONP2tTlTf5P1vwx6sm2I8tqq2QynzrCAn0bt5E1q8jj15pT92r3zTe
09uaOIJOf52VsS2udkNIsCzwH207B2Mfi+ywbrWLFo0jR9afvnfze3CQcb1w0Z9W
hEH1hm2mEFvHPZwPYOzAlJ5CwaXNiGHryrefQnug9wdpn5ccSIulMf8qK3CpB7eZ
bI7yoMZNdfHMSjvaizVKkyNwf4UfnWqBuShWmSFUKm/GP4GxNU4QwT5ZkI1iL8qb
0Mi8GyLT9agdSc9dnT+bhdo9877naGbDc80tsYMvfkzH6DEMjXEip+fS0ipeOi26
JM5diF/VhQX0Yql/Ga/dXi1Tjh2D6SevMiYtNAAKDzz8zLDfz8S3yNdZD5QgPqyy
LDswNSCZIrmqpLWOcvHSRxiedbF35xVpbezSq225ohXEJ/DE5DW9xk0fUSlkfPwi
l1YXmmCrjvZLarHLZIHesasQzuH/pLPg41fGklms6LHcBBR3j794/QY5iARmBJFi
n7rOemDe6Ng4CBxSST+vQbykF2Eon3FF6BYcb9YA/jY1t/QDkjHglQHAJdXfqaFu
ATMRceFkVdBbNTnYDmoAH0UGGo6sCXn4VsdMgFmm3MX21b+1jnalenwuidAL03rk
Z/iJ+i29NOXXDhGik57XVthyLG6ZRZ73PT8fqfPaCLAmtEFzFst72NoagpZDwrUG
Q2XjrBPSEkmmTpLdhR61GDw+4nXwrr8B2d1wTrYZNO8erS34WdYlES1gzoUqOzxG
jKCc91+6NAqC4DlC7IVmUBkGJvL5M6PblG9sZj528nazVOcX2SU/qtb1q3iOUSsC
ZgRw7c8f+DMnEbPKgMmG+hQjzWZgwiPGe2uBHc9obPTmmI2m/qDUQIKV+x3NzMYK
VMxwlr03wxaaIcTrBDGBm9kowBSJ3h14ETcU55rBBwmfzpjI7n8yDZZZ65PJjJaE
ahvnFme5gbSPis5cRWjo2dNIdaIRrSGlBatu5cKvCq05Q79n5jlER9L6HEGCVsqZ
k4OrIxiTPoF+xMag4L6b1fDstqKBpsnWpcRRnmY2maWtDxwyS41EFeNqw09bzFCw
+ywgBtYBqcaLGjCh+K6Mam6uhVbI2mxIQZIKvDljMqNOPRYJxDzqHLPBPI6qDE9g
tUVKYhUGjm9GrRaYuM738rUZyOu1qj9l8X+DggQ55d9Y0XoLoduez65qZ3wJyzmw
00BGxLBHb9gUUypIhHClJueyX/0f9tvi01EEGkar3Z07ZVzVzBm9Fq/tOOydrIW7
IywWYdJ6H7/H3x4biHPdmdKLj3PZxEDPvrgqFobBr+wD/LNgY6fBWZxhDG7DxpfJ
nRgxep1O7p39KR0QqDShp9kSIRaGsWKp9p6VbvKC0X24VacnhffdXEkaR4ZMmriM
hLtZQ5zJ1E1m4r3rKvEW71jaRBUt7l5q3igWvysDJ0npwjIg/lTSUhS/QEtO0Ie6
0Ph06sodrruytsR6otlJjl+jDs+ypTqGmVLFmLl+wlHj7JeAzZJhlXmfMvpiQp75
SXHJJbf1GexmCc2tqvUTovL6ZPSmvgHVYQlBlq+Ytii2gQGMbIxRC+RjqiLeaGcI
hzw+je1BO0lQOrmbr5cMkgyKCEDvRp9M4y95Tb/sV8LKHepw7EFTJ7H5v8GxC1O+
VIIXQ9X4Tegj5fwNpHW4Vx4CyXLfAxmoYo2v9fI3OJJgHSi6ilHODLdPtkYQX8Yu
JGep1McvW75iRtMdSQn5N+R+5tkWHZ6ysG5j5SaZOQP7YXX+8xsKLBXPULwiysRr
qgLEP5VbwVn2RKr7xy+yLjTkeAMciSUrWvJWl/ODRZdYxuzzFbZCubocStirChjG
pc5xesSuAHb2LYjbgr1TFS6y7nnckEzl7/aMKfqeOfgmSfpBt4IC6SDE12pqpgjo
Y/hI5qQln4gI/ssS1qVwDF2oLkgfHkmyGxSXxH/UsPw0O37fofcvlE5lxanYFf5H
4l9ryVKiY+YkErQAJEbiWaKIlVYDKAAjHis3LxZUTUl2A6zHwAAfjAmUlJmAlFc8
pjXm8lv3bKLIhcK9cWvLCuBbyzHkWHnV0cdytLfa9P8xkhHuv2BuSGaJJNICaQyL
hdhDkI7qT39OqVv1oO8zvLFacnIfo0rYd0XFLcKpyxOAS4S4rurybQyRbFu8w/+3
iUJ7f942QazT5pfelVNqf57P4nZ9Y0UAUJsk1PkSoDqVePpamPdb1AH5Rh8yV/cu
cAyLeOGU0KDVVE26WguC3+VpQdoBWriIAUV8Xf1vZDDzpzZ3NucG04IjcBDXnrd5
2vwm1BvyrEoiciiuI9cTvW8rws47cnhnxN2GvspKXlo6kxx2FByieCAnJruIPpZy
DN4nP507gwDaudie7Yk/W4PZu+Z+VfDreXdeIQZQMdwgTQkJdGZQREmJC8Ur9vAz
7ApVJIi+cYSo1rSABrg3Z0gOR8ipL8tqqekXSMxJBtbc8q2aHsX3p3zTaDb3/18X
sd2TdD5NURt2f4+1t+RC0HPO4WCmofJHQpplG1q4NphUZJpmZvaoxt9r42UkuwVl
oER0R8GIC8bT0DVBIDr/GLfMHdj0Z7j9oFfkVYF6Zzq2J31ErB4AW4Zgpim5wOQD
rru6OD+OYo5Ae1h77kp8WW3ttv1DG/hxNSlLlK1dtUnjKXkcu5ZMa1zNraQ5mlpP
nPUyQAznp2QjHT9wTKCVnRSftpGdGePyZ5+KxVvJy799cTXbmOthqEn/uWje3S4E
X5ZV+f3chlMrK1iLAYcvCipZacJ6n7i/mtC9c4D++rp5DRGCJF6i+q+mHoIQd4Yk
CwriZgaWPIEgepkitduxTbOkK/aYQlCEMVAZ9S7zbpmFSmHJiY9zgFsFGCKaN3Qk
Ocp8r5D0Q9r2RSLrJc4rT1ILM145+MDI804HvT/MAekxzUMqO1i02aElwP06dqFE
57hV86hDFr+LPgkdeoWJEJmUHrvLSo9EpQO0oDmJAzpOWbMmERKS99woSlIxdxz0
IMm87wtbdP/M8CQuYfWxB/bi/s9DbJdfs2kx+5Uqj3j6J4Opgjg/SM1dNc4vdEL4
yPnrlqY743xyyLfMS2BIPk/jhtDzkjgvWddPRtImL5ViSZugu+we8ut9Px48Kg5/
v6LjGyD+aCTMX4JcNqT6JIkfnXL+yE8Gr96QUoD8Ru2OXCd2BEDv1Cb1ezONxG3Q
0q+YncI9ExQp0w+IdMDWRraHWcvFFxZCF+pTVYS6N/xwave6knyxj0RMIpWdfQ5x
SSLgOqWHQaNIDWUiFaiq9ZaUUsRq+YC1dWuLnXiAPIxiYW/fkGs+yfcFjBjS7hvO
tgcQN8mcbUBOGZoE9qX575mX4/P1MB7cNtHCqLz3jXSZ+9j+2a+ZJpTxwZkYbmku
So0S404L6hrSGtBfjlVE1tisEVGOCHbeVT++qYYyiNyV4QSh9abf/zXyqXzAspM6
kfuNQoYAVSeCjUdPGDHG3qEbxLtQ7EFzl6uD6EQmGNwVXkNCZNfwZDCrk0/kYp3B
+LLtfDx2sV9plb506EIw4X2ZrDLW5WpvaZCnLafnNZk3RKlNMM2D7RksbmqNeSKh
iWbPu4mEWbVSm/e2mGZhOF7Fxy9p+ARDWRWV9FZ7llIjVox/nToYTieLR5hzn3ZX
q65NoyzMGz0W8Ljdlwyk9/FwITKfHoBVIzJR0l0cddAKFtbDQrNOXtckYeBztKMH
4NXB6Lr1cfOq4/JNCixI8k+C8TYJEBVwNJaqJAWTecsfToql+PIF2FbkzaZOtml4
2sD/iKl57QZKTmqIcQl8XSxBF+n+GCAIcQftW57A9NynT2JAih3w1TggJcmWho8W
gEqBNreMrZpWEMd92VaSMJ/71iBXMKuysCgm5V+40bPoL7MR/DFGMkujWGKDbpQ3
HO4kqZEPp1kqfL8VazFPHVEnLy1RFiRmHbalm75ob+0ULmsRQAdIoCQDD+HCR3DJ
Bql4OFHW+XjfRx7EeFBJgyFlFLRBQZTHAiThfwDen15zFMv5jvCuYw5xKozIErbu
Uyb+rHZ9CLRA7X9mx9RbegTOVCJxl276XfFt4MdSUP6qTHCXouAo6YVfwbgTC5OL
k+8sHUbmBOR5zUisPyfQY0CUT0NzQTkGQ7o36nWpmRE1pU1KUKhTRu+6lnCIO5Z6
I9ZHtQCHolaz35vT57b39aXlOOV3jQVDnIySt0vhTLCCDyIDQe/kwnCqarqkOeaD
IA02isvLfuaGhTg9USVIz+EXWaw3rWMPwThEXQ3hEWN4Vq1d4VgHW+xc2Xd/T4C1
QmDO2Z5GxkmXZBIRvQI9NNqMHAOH96x6JyggChduFoM+XTP7Xn0ZBFn0CxZWaWLe
TDgmRE+VL8jJcrAjsz4Y/+SAHEcl2SkGzy6tXrv91pAguNPokjmKpw84n0A3TcWI
ttCFHdtfbltVD3odVI0T0XrQ9Km8uFla8zEsZrJNUYKExZA82OjGKi74uODOBoYT
V1m7snuty1Kt+kXj8sJAsOMjFSeIXvocXAW1K0NDcixCfkeeZ8XMTwKat4Tez9M4
U4kZxMpbEfKrbHzhm/I2t9YuXTrEm5pI3/nd1u7S7xW8hTW8wp15O4inrR3k4TD+
BEgpMPWOKNDicGqhSoK8BIc1OOxU7ROl4HdQbJpFntNlnm2qYgw95F8mPlf0iqz8
zAwNua/qOp9F8zKvUgyCWSVBQcswtjxcSt9ir/tfQmSovI0TGaureeUcB//Xqjg5
2I6H7UZdoTIztMKviTQhBM+0ztJpF5hh3LdfS9Hw2NjZFwIs3fpPbyB+fBgLWGB5
2vqijoEdQAtrPenvl/N0P8Ec32l9j5qK02GLnNr/absTgNXpSq9ca74eBSMKYmeo
I9OLVgya5fGl40gHqVpgpZyk/qilXl7dWOZHc7CkUlzKu36Wu0RLpHMsBzdh0zES
i2C8yZM/nCTJ7WScj7WKy3cXpPMLt+uo2HjGUDJaHGCj4IzCO3UiE5ZSc/uQADZ1
pNbzIlSaq1XmRA2o00csVdkYskCSjpT7fLpVnyQzxB58vuftv4bXpGFUGCneHL7u
h6cpSUv5F0LrUadBhb9zNJjB3H8ktRI3270BleUQ9i9jwCMTBDy3qewSjOHhovkg
vkcFdThhlnGfSeRKayL7hjOU/1crwjhaY2TWPrmzVkyzCqdQDwYoCbS0Vt70dl19
K8RCmKemGBqsw8Xh5axqx72DbD2NZ81xTLu/YI11+tlguvXziCLl/0dbRNgJTd0q
7peD+WNNGd8uUzkPYYW3eKCq+pVVVzQZNpaUGlj69oBM2RBJ39JkEkhepfGqYxwD
o2wrT3m7nWSP2MUkLe/KLr7lzqE7mU5UB53YFK7RojWD5W7ob6m28vFLxxGrmx3R
ZsyFolRQq9qJkStkRolDU5PVE8GIjWS0Qw8bKl5VYegxfwmAKSdHo22k58x4/BF5
sB2zlZtYzKcrp8XZxI/VU9ponI4pzVDazD+eagOt6Kojz+wUQ+L4ack+fDX9Ihk6
lixQA6qwm8DYTfSvil1REMLGtvX481Wd3mzOyxl43XYCTgWoparvPX8sANoYJezW
UxqXgN9CmKfRfBroRnA7J5/pbXJKB+obfeM7sVF378audsx49lbT6okUd8GhFNm8
sjlm5bzv/V0rQhgucusl/QE72yvNS4aybSOGckE0o/PmJ/U99Y45L1roq2rCLamN
IGnlL7SLTGKn0raJu5yFH6a+tisQ1b+8qdhYwz8qzsA7yZfCLhK1St4mVGsHL78r
0vkQ6oGTh98O/aqKKrWsJZAQDvDzj12yIZ+kpWd+PYu7ubM6+sXKMhzk9V4MJaCm
Syu2kUl9deuccVMv1p9DV4194DqDe0WaVihTNmkF7m9eQFqwnzUCrfqm2TOtcG0q
H5f/xwG591K8X1NI4+CLSDc/XeYq58yakmRYP/giL965yoD+5sjHQxB6G0xqtlUF
h35Qwuo/3TGr54ciac5d9S+O6ETYKzQ6WRjBOQE9P5D69Thd6+mkIW0wZ39g+K2l
CaeVEwFXTmuq+3vk+93l70eybkgyYTX11fa18RArtd7nHSAegF8Si8ePZw1KZcui
kJZCFvzO209w+jVdRyK8cW4SRbS4xvJcYVbkCqi8oWsqyobMuVqoIA01WNUDTZLe
4QBYZ61GHQfpgP6BccDAeBAK8bvpyQaP+IBe7IJR2x6BmNgZwWpwppEGaC8RwoNK
av6/5zYwdhEQab4jr2BdXlAEQClfHRgpRrpsn2/UUlJNLOuT4KBop8Ecux3TRBj9
ME81SazZYIpVTFcMClRBikgxnyC6ukvmYNImD28Ng/2BFTHVI6cIISnJilEkVaAn
sYs61YOaFF3ZsKSxe4+TeI/mgnFfrT0i4tNPeQchJOpUIVBaMqCcyiWyvTa08094
zyIOcpraKXJ38tYCZKIpfroisAYvW50eCoDGhLRZmgMyDbvNCBEL3ELsPfq8NC0N
CBUMgW9fC/dxmux9n1Q6bvAh7Ij/8eyT6Tw6DU+OKvNkB066KQTrLKH2xVFCMXCj
YFKjI6GSghFr6gaK6IqjEB5MI3dSAQxpFC3ZQcXZg7tJiJh+iR6/MZ2VmnsOHInz
PveMFaVKCM2kcx40Ar7RchoxRqpWZUTLkQmoKiIMboxThycT3L6ijzU9+wQ1PVeu
VLfCeAr/K+xaBe37URnULTW44UdvldTcgZtU9ViJiEkYcS7X2DguJcP+D88SjpE7
2FNRhH/nGR7BL+cjOw9T4MyQJLZsCtA1gsIIsZmc/1NvHf5U1r/zyVjJxruTUGYR
QwOhDacO8eHeQnOosjw8V/nVXZFd9uWGz7GVhDK3rhco4XwGq0Ekg5hyJ7Wh0OaZ
ncS8M8Jsl8k2saYFKzfiweayTVRQ2kccKOH8GTow78EbJTyzIGFNaSgnhHLH0URx
QIehaJ3MjbbuKzY3Jl+61Uc79HU3mreQuTMrlfHqGk/uqzyJ7JMDzNb2TvQusrhK
40UYYgfHh5K3ybskg+TxAz55LzOXezueuBR1stdCcNOb2+13qCWudyWrtE1Jb06/
Px527XXwD6CZUPPGf0ccA1pb6RBOSyA5Tk7Vi1BMYR3i6NcgU2sc7OjgVhPiHhJ1
pRY7LkH2PDG336z8EWG7q+6hGro0/XOeaWhps6UYewRlBYYOUPS2o5dqNnlQWH8X
UsdsETPM4bjuMt5K/PQXORG9I3t0j3zLk6l3MjlsU8X01J3Lt854xE0isAc3ws6H
KBZMdjyXR3vGt1uRBsjGgJthZEDpppNWTSKQ7hfhO0WkP+lps28hhsbmD+DEUUZM
Q1tycwe59T3CZCFUOJ/tveUZKw0f/CDxlp6v6LOEFHVZKYhzoV7s7LZYrFmcZ3v0
Qo79VJ0fBCg0pC+WfCiYNhF0PTRgsXtv7xOZKpWufKrInxN4Rhe/IXne4/j8rR5Z
FDXuheN5/WDfgv1gJRCATw9W4ywUGjV4l2h3otGkVXmabV6cvKq8LCBN6MpMG8Qq
+9+Y8ssYFCKv0NpOLzcsop+juChUHbZOVjs2XEXok9RPKfn/VmpMR+pk1Z7Dgilg
/ju6g6WE11//2ZJkWKzEGNyPfywJZgYem8m8lh7oTmrcQOG/5LtmrxcsdC3+YaKv
bd6HSWxrDUoQpMlu/aLqq/g2sdOmnJ4TYjQjV9xu0h6jUe/NQzRVNO4HDXP+Q2cQ
r2bsfhOxXCxV1d9iOLHD3f/OV2Ifp0ojtWVdLq8FT8H5rqLA/3GHaptA4MMpW7yP
OJECglVlYRCl9KMzxxA3Tbve3NejhfgpPMhqqgQDw8z5FspUBkDSWcTupeCr6eYy
K00CHDSDzlbYwsZb4OoJ9SXI3N+o/vC8Tnacx4U9mA/citlEMZVYWIhtrMoxG0cP
+2HuVl3p0RixR4W3BJAJ5E6HjaBKLpQ+hOHnQhKx+edGgzBFLa5PfpssHdDlmyVW
CKdGIAzKvCphIGtlLQk4oRZpEwiBfO8JNy69VXHjNg3hBYVIlC0bkEPtGrBd2Kli
bHBfN7GS9eUYa9fVjntygY9WiL1VRsUSokCaQT5Yzc5+suASbG5RNJCsyfCgQ+pw
S/bnNh1XlCE7/wdBAtN1fnQJT+5h51ze8YuVWWEgnLiRcfj7oxBGwbFy9i86K7JB
Ojth49LyM055OUtk2RWohMMK4Q4h9cegk5PWfS2oO4r39KmhnCbbWlsFTEQ+b8c6
iRZ9IPpCiBbsVJIxUcb+cNNrBIazpzOPA2Df/NgCchy5LZWEWdG0YljEs4P97VDQ
XgWK0wllJnUFb7IHo4wf5uU5JS8M9kjh5seR78JOJcJdQN8Ify4eQTZCGQhPHpo6
jAu/jqDVFzge3ZNxASFIDVr3X3PbBEXuR8dC2szBScZ0OYWf9SfNAa4LE7c5uUKj
edDT4TE5CCnSCAIChhl2AgTgxK18iVcDvish5U6IXWaImVyU+VghLZCtPHxIaggi
oNJQKhOS5FEH0vd4d1LXGrYOhC0bzz9EYpsyL/p0j5voIGly2gCTkoZ6n2Sm/1cW
vr9VH9tpGbr2czlQCCOM1ZtdZj8wKc/dGbNonISxuvT6s31Pn9ALjfALfyMS+TKf
KLoU6l09+0uJESye/nj9xUb0vBm3MRZLYlPz+nAHJtpccRPTpTb68hI+r6nZ8Ljh
Lr9GFL4NrC0yFK+r61tAXARpmqEkuCOors4qYnYCf2O1ruVoqOjqe+FSymcWCEUZ
jw6Ea3YCFxqh0NfEIqLhV9pIJFnsThF3z+CTFQvFn5p0EgF3oMuDJwLZC4dI2BAK
gxzhf9O0qpl2FaRA/e5+gGjx6E47TrvWxA5uosMRIleS8Jb8Y9eckHJ3KGy05mlz
bWBPC4XeuCK9sdKR2V2nkYlPR42gtgglxrbFhQedt/MHoXxfEk7bo4tKvcwrllLp
bwfaG2a9O156KmWylnx5eqFV2vzM0okjuJbfg2P9RpQS8ZRNXyOkqw6FCoFLwN0N
53E6jWa+NuFgLh1JNrhMZhEPI79oVmlRRdJluJhwpPab2QQAb8cbKaoQM3qBQgYo
b48/k02if0v8FYzYXCrTeoHf+8zmkDvbr9ykLEDolyGbQvCUX8vw5Ox7y07rI3YR
4qwrvMccUu98X3vvU9xdSPd02iQNDqHnx+rMbvN5NVbd3OdaS7HpidLfenJ1onOJ
PRE32/5GyxFwKcJ58oK8kWc/gk9jGxNNfXsbJpu8lQBKZAI88d/TifgDVn9Eom+2
Ri9LyJ8tVDVEbz6/Ats2zpKsVLScLQ4D7nD03tcNGoY0wOgDJDG4/PqOe3Hf198I
jpYfxC6bVJAjVUyzke8aHkf28JdLNk58YAELUmpVYsxRoQpKdhy3uDhReHlfzho5
v9Zn1zugypdNgwvE23OA5ILIWNoYpbFYwSmpCEUcXGv3nt+O4ucvoPPvWQthk8Ln
2Exsp4FzZhpR/QT4GfYdC13FbBFQr7ixysO8LHsCACskbsdWODHi2/bCZl4D6Dp5
pwLCaHXPQtu0DjDTV+wa33jQvzRa5uNEZBiuXVT/6dZlYQzoRJ+F/+g0DBVX0oNA
AibAaZ1yP/hzH67yVv2BgphBy9Po0XkeOKjbhRJl0DMCjlUh/dKqkNpf1Ki6SMbn
C2u/AyYwKeYzTIUXqYxU1ERbf5RmoHC8/CKNpTRM25MJaT6c+ZzdkranRSm+6VAK
r53TjGRk/dgOHixilKA+AZcXZo8qJP2R1JQ6LWHkYguc8DQgdM4b0tXf6ndh4avG
xqDRi58VWI96qDgRNOshW9tdHqKFZeXwFPmg4gdiTFPTxoHqowDRy6rRAxWxHWnD
5KobAJyeS2mpVBkPjRGRovIvthMB7Ckr9qoc4a0go5oTaFwTnRMWDx6SYlHbxtOY
ypi5HYkS5vgF3HQDGzzIYOhOF70llaLJ4V0KUxnUdiBAoWWpjWVmCeGCbkkoZdLW
T4avd3fSS1NhV9L6B1ZuFHFDkI/x6MLv/Y2c8390Mq0FOrm1tPQiFA4MHydO9/SN
QQWxIwIz4ZNPfkeN1f1+Y2sEKNASF2xC2F1S27M/B2f8x5qyofSfpwTZ6YDVMce8
1DOr43KGdP5fX35Iuh7Njo1+tupm57dC1CiG/m0xs5gilMV/BBDO1K+TJGwafhCD
dbVDebXZbi2NYRmPO/KXx0Z84H4zXgFhTLcVznclwfe2ZS0UL9fXRYlqYvDV8/Hh
JlO0uqNBFDoLPvwU9bcCVpePBS22uRCl2ygompKx8ZgFbpy/kVhvgN+HDIK/E1VJ
3VvhvWwDXngEBxeCbtUVSpYDEVoz7Gw6qnMOCwxaIFxErpmgTP/sk58OxqCKN/0m
m38Jxwo6oYOWG6jJ3qCvmL+Y/v+HDOu/1zqD+byC7YBvMTnNhHeNd5Ncpdt5pb0h
0c4a5ssRinx0SL9287VBzXqV8lLR4fmObtjMrf0oRKNfy9Ti6aJPp0QuzK3/SIe/
WeGZJqWsFpNi3MZpSW+z9/ClLqKBXO5wIwcNdF6mRErSyc+Bn9f1MJInlwpEDFAa
DulpSFO1ZOcMOQlpN/xV25FG7DuI4Fw1kC3pMnk+pynJV6bu61YNhlK8ae50FzFH
PwfLCpYzPHvEdYyayyThR1mFNCStuyP0ZysyDmr2Fvunapirlem3sSSOc6uYHosG
vbHAqw694tFaJa5TqKZEWlcAC+k8rBMO/Q+ofCHmiz3xLYyWYZ6808/zvyZEtmA+
pVssuzhML1iXFcLcqLVskszxsBltSUDnReMLwtUy0HQWcUjjmPOfvMLpyS62BvpE
YV79AaaENDnG3lpmhdd12E7pk/7aVedJIOa08RQCrHHC7fY9uV1BQ6KgltY6FKTl
VG/oyQODzuTfJgaLW6BplG6wwrm/sopxCASH3U/n65Spw0/H6agzqiK8rT/Tgh4f
2ZbgyNrJO4Q5n+xNFXxR1UZxibvdzg0pldlYMMypwc/QUeu3jmxHPDy5p042Hty+
qHgnUITz0CRJjd96xYclh+83pDjWun2TQYEhfTqpR4KH5Bbfe+OgAVpqOfVT5Uig
/6vRh/3CaVnyp7YorZWKz8619ehxZqARGtDyTB0Oq1Gd61qTR9IQDiic4Fle7byI
qjpHv3sckdeT+NNg52VIuTH9xuOoGVoXrVKIBrDZIk5jWqW1FN3+QTbLzJ4hyief
6tdmQau0IfNLG4aGruGVM+z65E3rkDoW1PMyJlQYKlj3pVp+79FPnwWq3ShMjjCo
RXC8jOaAbOlYqKBC/vldD9knB6xA2FpAdYSoYUQh+Y6Mq6Pp7MC8LAWzt3XjudkM
wtjsJ2a4Sfan8MqbQoFS5TLD4J81HitAouXyuRBPTE9jF/AuUnwlQZSoCw/DE71E
4uYZijVdGKT/9X9AAMe7l5nOv1HrQnbzSo5YhXAbgY2sf+j+u+XTYOgmmAmxW/Rg
UuVg6r2DyOn+OVS1H+FzyPw2oQtWjwhGCqtFQT7Kt/f5jbFVhGzLwh04Vq2RSdag
BkR9ZOwjxtLFDcIyGx+3C9D1M+AghPHRLZJrwLnivCG6vIJc+MoU4Tzp00Y9QCzP
CHBrYxn58KtKE0MDX3pBflBymV40tJUlCdkCCTnCbkHSZVPby+9YjBUySbEIEutT
oNtw9bq3d9FzECqUny6MTMhL8mMaRdzfz+XhSTOihedaWZe7KasSh7oSUfBcq/Wf
KZ0ZXRezcQ1mmaY4EjHUCxC3IF4Pxsv+6SAgmHUwLulJRNgyVjW7Cg5RPHhlEEOv
yJ7N21oOBZhhjj/+n5sKnOcBSTB+Nyu736YEVp8V6m+j6psY3euCr5P5ZL5umlWX
iusv7ZPmgZQcOEzm+ryBMT8Z0bg6bNh1xZuvG0zxOU7x97VOfEPUESxmkPUrfVu0
eqivL8+mIPeYQl3aXcr+mUW8osJ4WvyWLdUuWlisuuAzUMjaNai6MSmr9UMXQQPv
8zx4mI7EfV35Gohm0Y+XWwzXSrRIfVvDp9ug5M5hboaJtnDu+afvL9WZsyABG5CL
IgiQMwX0/VrWgnO8C5AigV+0zZlzw+6nB0H4yUNwDoFzwvKuKamnRNBtCkzpwaeU
QycWkPEDIBJmu7DNGKzRmE0gCLoF2uMwUojcj3E+GY093mDKY/0hZ93u5UBK1bKm
sD1CccaE1q3jysNkrYEZK7cnWe5MSO23B79JQpPFSaWxZI6ZChYeEcc/RXOMwpLI
7zLAm18aJOGHVj+H+ZQwfduDxBAKaa+uDU8BtfaQCeq+8GMuoGSXfj5e6bLYo4un
ufGqUPuWCtK83QsRRJwVJhP3uiuZb+a/a3jGskgixfsEbZxZD2MzSEHC+sRUrhgS
SHrf5G1A0oSWprHMhe0MnBALJ8WwrEbNt7VsirLLuOSTTsqrF6PrfCAj+toUMAu7
XHnloIlWVczbxkCoP2u+MYLesEuPeatDott7IqK5XNNFtlhjb9aBHz1nxhOSMsIl
BKuRC5xrnEmoyswVejCJQaNa0pV+SKrteEbp4RUiiwJinyaNI0NsILo3MAq+Y87z
UN2kMMzhaGSavBKBou9m8+Oa83oWXRDu1/R0Z+cjWQOYddorvBNup7y/WNrEixos
+3+53r2c7fnVPrVSx6Z8d2IxvFxZBXjZEo70LuTeWqAUCl5neoPI7vJdvyD81gXK
y2yzuWoU1KQc/8PkONlN/2oPgV1DpyG1WIIWHsycy7QLL+FOA4ZHY5mvXLb3ZVGS
Oo464WVn3Q+fFWdAEh56IqWISKuq4U2jbWSvRv9R0o9u5Fm8unaOlCMJp0l/0uCB
gGBeiXtirH8fORRAJSftlHRySXC5hi/IsMz6WSKnIkfP5zasxojBIzO0FEY1iXW2
Dt/OJW9uU4sFXpn00aq32vfzHqSnMJKhRJjyo6UDQmqQkEOZOOtUZLEYjaZeuGUk
2KrMs28gSoL0i9WZPq5TbD7DVMUzj/5ILBaI1/eDGnn6PSHZGixonJMJwx/NIcep
IT6Frcn5+Rgo+oC5QcGPeAc1mfv8TaGfoL/4Bouep2l56Z/ILGG2A5357g2/oziT
/wefwq2XSLcFzuEBK5ZAf/nDPUKUhF8nP7crpFMsBKRuIF5PEV508vH8ieQfcXf/
zdnXt1wRcNbVkMFx0k5qk0I90jNJGCEeqVsF00237Qi3Iq4J51nQDutbUvIfzwXk
JR74hyCL68zMS9mpoqCF/IA+1pvttydgeyJE8+1e0L6Z2gctzsRvIlrB0FyYhE/T
xzje3W4IAOv/Mox/1BpTeiFkJ4lm7I9ayni/lq2PW1OKDDpTyDcuPRwPhJ4cp9Av
9ly7Zk6bHI1maCAeQImR5VFWyXj0G+/Dd59rLkcKeYYUGXXX216C3QQKSgnAIwsh
rSwgGLhHQRbXXf2vvtUVBVl0wLCuU83ZSPGwQ78G7gaW4E36wYABSB29+qIKebV7
KqRn7u+JVUczhVw6n8D9MK/LqoJ+VfbUfkb7qVw+LCdZeZmq5euaqT7NioZgkQYo
AENHJBFcWkkuVIHg06mcbRmemTz2YjqV+dIK+F2gj1SdWK03FDdZ3RVZKGPOEA+U
Hl6Yqg+bd5APBzh+ezUXG5c9i6l9nJ6Z7Mkwx/xlad+QaP50BweZS8BBtq8LhVzL
DpEPyoqnhm51VQRHurFP4gQXf3FkeXGLADPGTwhqbCpi25ixfTc6mluBcEgt0aQN
N+pLGiQQbN0AnJLgm/W922peTOvyBWZmbdzzTYFms6QxdfrT1LI81xxAeRW1253k
rgHQFb6hlb6k6EUX+0pJDNNBlfMjcITajSo2vcDr0tfY3UhhMrW3juIF5t9ZP8jl
+QxL5Ou+EOzenZlDjee4AEAChNlQemz+oDAYsTrBJeoiWWvBTflbnAMqsP6xv9Bl
aZbYIXUNE+aVqsKqCEnwbvUxDMNRkmsGMmy1sMobFjmGe++W49kcf6xU7CPxWTKp
Ad3WlJtfkhI7IRQH5Hvhs4PAizU1AKI2Gug/n+mCeyJB33OBbqy+mZYWXeYJaOA/
TCeOg/Iyur5Pr2LOMQ21CwaWOHTjzWvX4hiuxcyP++TJo/FRz9aDcbG9uT9ns0q7
oUOhLRzquC2kbh0uWqVzJQNepSbYE5cP87UZ26Jpf39xfrSTzcmcHmcWRQlgTDor
WHZE6s44Ov4HMSamITTfbj/B4cy6SHWjdrIfa+PJJPCgMah2m3tdyWQaha/tob8J
91bAOeg38dKsIMMlbEMZXAn78TFGMPzduq+McLH5y77mtlW/SEAH8u2kwTg/FSsP
L4wZ+OT3t0L6TTs5YCBlbRbHopIiJkCPaBFXv3xu87YMQU7OdLkXCMehE/ukzROv
+iZMG7qIRFWkeZVp9aRzU+WBxKl+BFbqRtpSjv/oEzDApQiR2iz6qYruUSYr9k4p
M9lglQaDAvaZZ5gJcgeoIMbiztiWsDjyg5LaUO2sHXJw4C9Xj6GZJKHYPiC3jaQp
Eit1JAcz28HryJl1oNYsHl+Dfj+SuXUL0T3QgTFEkqD1WjvWL09lgrexo2y2aGbo
Vc/bETvHJ3/L4jxvNSLd+b2fKfFfSFxWfQhy4UZfA5SftP2r2oxed+6uMZ/zbXe6
86VH+0gGiXc7gxTnPX7klpDjf/NL2LBpI2KxxCWMosxgAjE0DO6OqPWvD4DRa5Cr
0LY6ZvcI+Xf+KLElEkDh4lAyq4Whp6aWZRPzrdBPqhNPobyF7dJWg09Py4c3zPOt
T3ImgK3bFbIPwlTwDtlSWtCWU3w4eYbngBuhEUy+m7CDeMb+UDX02ROHIBg4Nz5x
pSDZZEEZiJ1YF4Yc6SsalSK0tSW53ICGwdHZhuTAFOE6wd63mjA0/mgTJjPZfrUE
cIi1C5lo3e19HptOwRHNTaFnov8cdwPECJfjPi/TfRiWBJBzlx8+IcN4HVCYNVqy
jvaXM5cmRUsblhiwjv1b/ULZFBVnErgKXtgPTszQnotsohQ35zkL9OIW48ktiU0z
K8RZWQ1v/cp0HkDOqSXDU3EzKLvqydeZweMj0u7IN7UMqR7w3kNhKVG20D/b6Sg1
fxbl+I00XkC5FHO1f5/kS3NoyBhYRZabbUPPrMHVch7mAIw6Tb2AKWHghwtY6kpU
sbsJAMg/fpXqoAS1spnIpcm9fzvEiRXN/CbhsuhRLKgbtwXzRkM8hpgo82A3V+Dd
TTmAudKc4SA0Ror05AbWd4g016+6nUqhWUm1Ww0nEvIl+KZcruWDsKMvloK+W3AY
+9CLBBNJucjY5MwUq6lgKLVXtNXXswINkun3bQrozvKRH/J0SiiqerH4RD5vEtYh
EetaAOuQVX/MBQumqtCOkiXNoGYlmkdjbGvH++fyA9CKc8uhn6yPgrd15tok2C6n
89OjGXKU69t01XnM2EwNed6qhCIxUCJdO+xRZg6EIdBdW1jxtt2gOrvYyfQ69uAB
0RyAPT7eVPuJaB26iHLjwpPAvhO+WmfA78D2w7Zni+ZOne0qY5W/+KMkUfTGDqNg
9jIcSeaLFF2Nio1nACxJUhmTy+gEFdl+pviZDPA8V0BAT41q5P7/nOFdEKnrtr0m
ewtQI8o7NwZkDtEnNoicJvn5PHcmrRLwBvtBNwNlIZumQR2KuI59+1FNTHTv7h1Q
cCUfVeM1/LVUL+bBjmyrV3EiXd+b3/Z8iy4SqFaJg9pD2H/a3VQT/FQUv26WQ6Je
Lvyrhu3nUdyFywGdSUqSwhLe1cWl2PlqMXUK7XmNZseExGafF7KYwfA2pVxBD6iu
gOQ6DrRsJlLvOUcv/YFBo9C0TJi1JRfSU7zOsKuaU3CKs5VqPI/axfXDaaMooRNX
EXauKkEw6WTlFM+MguzRabFkQzubgSReEnsRXD6opaK2UTHv3GrHtUomdskWz9Ti
Xx3wpPF4TJarUhlJ/sqx+nXOcHchxTWeNYqfeIrMBOKLVaSzc2x+eXyRCGKd9uv9
FnbB1aN/San/+NuujknyOc/CuRhLKey2D8f33qH6C98KTQsH4OB1FrWcfGL2K4/3
kxsvO7vQ8vKsqO1MnZ2LJRPtkJ7zzREQcV+yKXvHnI3ezzbqoyyhNtMUkSboKhKE
6tSyx7YJV6ovOgtZhdXl5zoea3AjAOoab7hQc99d417vrBmHELNTnI8erCcbf4dX
8eCT6Qq0q8Uxpp1ZEv60GD5NixexclIlAI+Lcsq7kHig7UFphNMjJcHj0MhZ9dXe
0dG1C59BSONifPnyQd74qukrHObSMihWELLGK+NeBlEoGamTvkul2gcXXPPZxsIr
8zuSfrx67atS49tfkLQoOSWKBfLS0VZy7uQNbUdK0TAOrTkxS2agnKA3VpwuXn8+
oKONZ9HjcbHHJEAvLlFTTmGdBIdTo+0frJ3Fd0/oZ0zUIwxDl7ioXPP+DwrC60ry
kSaKw9F4+E4zRkTAAiJJipctHQxC1OayOIjHTz+778yao/WIqObVMcQNX6Prcbjj
2aRCUrG0hNAifovpLqBmk8J9fH949T2GBypAz8YzXoQiELIAOIlatrlEHP3rig8I
MTueJklYH+WhV60wHEQoudfagwuoquvyJQjDObQ8bmhmMPpFLd04LCHsa9QTTCXZ
nY4aSUxibHge8HEujhKAfF3tw3xMdqOPGsMMGRqAO0VIthEIQWkCfxQZTZce3UxB
Q1g5qlMWyFZQ+Ushid8ck42UlHg2BkhkSfAht0K9AmRqmh4laho9uRbJVO/jz/Ei
oR+Ok0HGuNt0YKjaspqwk6H0+buySS2ySLz2UEpGQlE5wqYoYo6YdMmUmOUudl8p
ZWBeUeTzrXHHPN4IYBF6cYr4oxe13HFuIwUqv1lZnMacn98DM79lLwISVMcRUyRh
fNih/9tUyRldhOX6WJKsNkWs4Mj5EvTNaBfh9Fdu2d8YqmHQU5C2JrtcvTOWYGGL
RCeOvlrl53+Z7+8OGT5eXV5GEoMxDUuQ8TLgFQrtYPim+wxprgFbxiSaGKNP2CcX
6X9WyppM+hKK94scEwxjx/qjzxgmK9kmSLDWZEjC2on6M0tn7QuclyP+OhkLTzlx
GPaCj/VXlFe+U97XzNy1yDzkr0jMWKe1ns+GQRmUGByO+O+pRY3VvTtMkbGkDQt+
n4P9QIDOrqv5pTYV9vo0V4riXKF21YNEzUghuWh2tgn8eup/Ae2GaB9rMSEF6bbn
KAkyOOBF7WNrHM/XmzKAjBVtEiWF9OrgITxu7+XSWwWc9XDagdXztNYjKJH44L+t
u21H/YPPbKWwv2oWLD7aCxd4eWJ3RWY+g1V/uL0pOfSRHBTQpKMweiucO4CFu6wv
EbmB9wDTEfJlI9PML43tS1aQTO6A/C0Sim8M/skd66FAzDxYyMzCn7apcAkD2SGZ
AXm24u79dLtAS1kcAtjH0YUQTSZ7o2/mSNLCaAGJ/CS4b4Q8Q9lrmuZXAGcYZ2Ci
Hw5HeIswYYrzSF799aR6jm0T1GdRJS+sSL3iGMkJ+obIh2P9cXxKggi+OZOBdtk2
I7UWyVqt7hAmAzg6dHcb8mGln7xrqVxDgJNRnXfmIw6k4wxA1naBW9kTF/SOmXIq
74wNYuIzRo8bQ4c75kb4zhIFsuPEBgRsIUAVOqxEFT0BWHRv3EH/5utlP2Ak652t
5uADnHhKg1qNAEsc9eXOL5zC7OBBHgKhgqmE1WIBOs55iu6RqkJO2bGAjl0sUnrK
hc2HDQPKxe9ZW4ufo1liwRWIl4t2bOel4JmPfP3HZtuvYp9zkhJdcm4hEOmOCGsl
lDMXymmt74vU6u0OWCbTIbjdPIZGnrRe838rJzOy5LD8xIsABpHQmJPi9HcZWN74
msXAOslzzyJQcep2T8h8N8zo69INeLzRBww2EsSBeFDIOX6JXKtquqaVES7B+UHV
QqgMxbUV9o5C4RYknyi2J9RjMa2M2v+WdTrDv+9wJXjweeJ3xMwc+e9PjXtljW3y
YJRV7eNtaCynqkoeLIASePY/jfNPGxYh4VV6iC8lWcs6vm09d/rtgFPTJhAj/iGu
6RrBd1SpUCSM0wt9RyAT6mjQcr+TbCAGxjZq8F4zwhFNg5Rwc0XhCkqTuWvW32cK
4WzEE51BYxbOxxIRDQIJ/zb0TtC3Iu3vS6TS0eMYnVLt9/y5gLOpDP2Tu9CIaTZE
Vs41uth2Tjxo//KpSMLmQaixQTCQBAWaSSvUYsZ/M0FDMvttEA2H4TWwe2Tpd7kq
2OAw6mQWnnep5e9Nr1gWtFETq1giYiHHdNEsN4SesUt0nQnCRDDoV5ocrDZ6PRPi
SFL2kl9ORS5P1cfVlBtw0EMsp+M2owQdmwWYwNhvK15WBOXwxLtp6yOrPgenqOsj
2959D9yLbHIc5fHBHDGS3lCONzgnsp4NI3O7YKmui4BpGZoq44OAgBF0iqMKoctL
HgQA1Hst2nk8EaizYLCnKThaXtizU4m81Y0DJPY4SChaB9Red6+V8NJVRRC4PGz3
Z9LNt12kg6IyrTt18pmAZDrXtd6qctlPhPVCFy5WlmIVzZv7UDPMpuI8hjui8hp1
pKJgwLITpp3/5cv7psxxMqszYjj7jonflTKzUdnmh7UAYQcMfx/bgfzS49N/sHJ6
BXwRocV/dvOPFhZVoEPa4ghEYEEw/99qWtcFVr7ASoSugZEFo9jQnAW3MQtwPquW
hbO3C2oj+uJ7dTwkk+jLj/1v/M81M5EdZSPpbPc5zduLNVMBiTRESp58jCszVERy
0t7ocrDqlQ51lii66nNJdFZphwF2tIuH9E1x3vW+pnhdkMf1Dml33svHOf2Jqwic
Fnuq/nKhhFaJBjtZz+3kkihu+UvAf5SrZr8aw3it8HsuaLU0Vdba3DMcM2DPhMS6
CmAEUTANU/0BmaQYHcqjFiP0LdGr+k15mk1fsRBK+OALrmK4V+MGuMV5lGYFN6K+
vW4n8n2Khw5tK2EPyoXg4Qvc6PXgMP6VGodLcZKJSsMR3xe+e8GIq6IHUgNci2FN
1nUO6lmtQMJ5c/s0h+I2JmaIhuC2xrr18E+CKJBhWyd1lYGhvtxjAOjvMUxEa1fA
TzWZc47QWlSxP+ykVwtVreoQWh5y3M+9aAhuxa5FcdyyhZr5Jnk5RQKGhCDcuq4K
i41w6Odl6u0K0R1Zx+rfEWHofXZBo0bJyKcpkP1qDeF7a31kilCEyr1mJU8OD173
/EtArsqHPvd9Dhs2ui/HXOUL5c6w+ddcJNolKqLXI/roj/UN0GL0DCrromY09JFt
/vUGABJ5XN5gquTP2/qHzGqh+kTv2em0WfTdlNJeuSHyo8t1F7oxrsXc5rgDsMgM
vSWPg/b9ETGN25qKhY5wXZpfjiv5Hj6Rpjg1LIY2CpZ6MThY8wYYS38LuyLxykj3
ipi/4knT4RZWVb6XoKPtnwlYtlcLKGRAjpPi6H562sW8zRzvxvBjEqLzrf5fhurZ
xOtIFzb/HmUykeEJPNTqgM2X1VpoaYEAANq3TQASvDj6iiih9cOY/+JL6rNMEtbV
5hWOBYrw+/HYpXWTbF0DbRV6rsMuFEXTqBV89aYtQoNJC7dafHZ1oGaTpw00ZF7T
fZks+q9Vl+HGK3ffMJIapKKJ+z6IL7uUro/b3SXVmDZf4fVOawMypYJ2sXghrAGf
9h3mHRrBOAg52ya1PpveWqyn3BZNFBRj/Cy8cbWu68KmmxwYlSzIfpibZYN1EWz+
P98p3exjYGEUdWmv8gA42yaMvp5CkTbV0Zw83sNEsqHUDaZ34JUMJIstsreBmRUD
9YK2FFuYFqYxSxbqX3mHEYoZdlluIDPAzoo9OY/DIQyvguXq/POQfhp7kV0oA2gT
PWEb7HhxM3TMshhl/GEBwH0i5sfTwAPsxmKne34o2HHCtkSIJweZ5RzsNJt7BQYO
o+lubBYObGi7VJcS/zbi4Y8ABTaWmIhHrFMPMsUpZxcKd7emEhwq2LXMavG+0HEb
X8Ic4AZwTMX31T4YaAFkKwvZLutTPYnLthYxLEwzOvjzBt633SD8iyCFWzDHGr3b
4nNdH5QHe7w7p5zPC+yYgQVB8QRqhQdhk4D2waw7DZ/vtJxGcPvy8nr0JbUMnOfE
ybsKnGkQHhxvR57sKudivZAd6ZQvSs0P2XxPve01bOca4IW5VuwvP3wL+SZ00kr2
ugWAN08wrRC03JlhCP6ZGzn8mMEdchWR1Hm9SNc1Juw+PZ+RpCRaWuWMnzgJHYdJ
GI9WhdiFmV7S7qWL0uFLOzPns/g4+hm7l9sZDlvD1Xcqozmj+J1LBVnWs8d1jtRO
1BKvlNK1M7TFCBYUv08y1pxBJ76FUS/+HGkdDOE6HyOhRB63kO/vy9aj/tbIzZHm
cut7660B7dGaWwgn8FF615/XiI2s3eZfVitHNwSsZHEB5wXNo/L3IuErqbgqqPM6
SM8x1lwfUNfZIxNlxMLXbuDaMUoKcW0E3bbI6biZdjQrr4lNG+s2rW05tZQ+8eYP
OQmY295uHAbbSB8cZ5WrXTNFwpxE5Bxua04gMKzgl0UFuytLUtFCmSFVQnN7fIKq
ATHlop6QoeWTQLG2NR6KZVubxGTtHrQmfHRh7nQFZki74tWBjOV/Sqla72tCWwuJ
/OSlQX59njNKL/rMtLOYgJofmNwWKJa5ckwqIpPEh3x7mG84uRrL/iBdqIGeYYtS
YapDl8YuKvrlboa11UNuMR06oGCZVyUDp1WUqZFGAGRZNvq3xBkRJybylzyoNbIJ
kYvnzn8ggMz0ttldr3L5otUUw9DsxtLPWBtqoHIAGF5t/CQV16Z+2S5gHl00xjdG
xKb9KY1/EP682vNUH8586mOxfQm5dSnfl3fNTulBCs5omBkDYHP/xS/wmwOiR6SF
QCQfccQ61EDPbDytGKNAIjFOl1A+OSr55Q/gJs1ReTKj2pTtD1sJU6bI7k/q/yvC
o/dM6AgwP/cX6DayLvoKqhHaetWzPxGM53RARoSrXy960S8qzALfuVcv25a/Uimc
w2xj2d+sh/8LpThGYujOnpQJ87UNsEOA4vLwvgAsz9D106d73LUIX2fLBrGz6Amo
ADwQpkczqfw++WrS+y7zOPwXvBaWB4q+MoDpiJm5B+r8A3XESvO/k7pzBp8PoTSe
jehE9zPos+OauU9wXVuV3lesrFCFSb1KOsb/tby5kdaUmEo+kRWvmLxaLppP/CLf
FQXekPVrUVyJS/x1UT8LL8JtgEFeGi+bwQkCe+2ZRlP6IR39kTcgbCT/srifV7pi
3GIh4yTGhLSQFOAekUVLV6J0b3RHbcSuFh3pR2dv2i9NchToFdimc5C1b8fQ54/Z
fNqNL3tx5vfOxPBwQ9m0VAvWejq+jG6N8LfsEFk67B4QJdRguS8vmkYF53Swvzz/
61YUK6NCsW9ux6OOl2QwBcI7zidslsSmrCrONund+K2cW1OTLN/E8lnHUXhBZBKo
E4s/O4r4kZ2915eHDADfYZPw7iAKBpYPu/G7BvxYFcGRNnLuOr0AInp/v8RJ3qjs
pX0XEeyjTfyEaAAFpuliBu9YnDYkEZ2RZzFNzCubgZMhf6iw9f7nbMyptHs6TTFr
ErNAt/ZO0H/WRiNqJGM67CnT3mJSWs/NvylcWlVNLHoLvtVxAUG36PSK7sHz4b6H
XMfmiVaGtIkdhFQR8cb8XvgcuJ08eJsnpYL0Ol4Rk1BL9+laJlx6VKG/q5Ffjcsq
yLRw0MqhkPYRzeZOS8nwVc6lKX9iPh7DHq8DzQwZSmr8lvtkL3kMoHEX1/zoMZtd
/SVHA0CUMyE8LmIgSW45fWtbr3+3CIe5gNJEoV01rywfj9+Yt64nwahegZDmZA+Q
qtNhm8u9lk/eOu6hJoMjaJhyIIHcrTDiZBWAVFk3cOtQ7TM7SKEFlrBlMIgQv25J
csUess3ue9GVQSjJdyD3aot+BwKDKCuZPjjGWVM4SDIrXQniThRsGcscDrtoms/6
six83r2My7d1iE2YmX+9XZD/dDOBRo5zqEHxDVm+24WzkKNmi7NwrLUccwaalacq
tSGal2Ik/EVoKrPq43cCf+JxVKj5vuEQvsZXyZp1TU34qKU+cLX9inG7qo7hFzp7
3ivh7QhJpE8h7BiskNga/3M4AIsRByW3KcSCm4tVFC6TSmHPk3WOI40XndhvgpC1
qki6yhRa60K3s6p6xiklgpl4ccFnzaKbTcyvZ01/S1OCm/ZTQRekDpTxXfuRmkVl
Ve83/1Iim3CQDrUs6KuR40rhogjIlSGQtI/IUTmNeqdY00o4H/RwTwwLHEHfB3ff
Wv+0VCxZZFscHIN2CrsDCY5otHv3DxfB+Neq6d9MWKf0vs9zTb4PSv3Bf4mCRYOo
G8OVcVHGRjpJ4n6xlFyCVxuOVAuFHlfJLiNnPX4JLhMSVD7Yr5tARl5dG2K3w2NF
9JiYMUwdY9WJ6Q6n3DeLF4ExMmM1UyUofBJVLy39cpUB15UOAoA1BJRkAFjaEZsx
fSAPiKCW9GsfP7vKtv7o8wJqAqGP6jl+o9yhgiYIUuVHrpS/thSWDT2TL1qttgDl
elAILkJjTkIGJMQHSGo3yq9UKTNLQ+FV7DrRy5WYDn5yRdy5WGLKizjmHpULW/Kk
ilgmmG7lNcVN0h8Wcpz+SwHHmW11wmyH4TcPVNObyPYp2JVBcF4qfdyxHWklU5XS
+zCh+3sN2WJEOrUNwOE5krLbvnbGbC4zzoazyFRJcT3JPvOUD5gVq6TrDoARSaDX
MBUr3+SGv5SMJ+jAvUqfi3rHuCi/EPo/J9e9KE5Km1N53Rs54EmsZv8viQ8B30el
Vb5TRwdhA8DjqxyHVYq5t/dBZ8ITY0vP7Nhjg0dWZVMEcmQ+ZFEPLcNW/PZ4HVFl
7a8xAsNMyFjhwjnHWCar2Ivb+8eY7jBUTLrrBsXAm6HXeJUpzJBzDNIUXc5bOAzR
PufXrYme9/Gxty5P7hMPOL6+px7HZMYritfRakWdVhdZigWkb9tUHRD/xFtJu5Ga
wUZgtBD1Lnl1BwW0ZY8JBgMgoWTQYWrnocbpdIWDboDmWcgbemv2Pw1j8D37cBxo
AOw6zH1NppgiRtuCWmJ/VNCNwjP0rYyO1Sc87QWJLwTeFnEBp4jIPIdbu8FXu5to
9l6PKGXa35kwKtdta5+QbxjT2IVRDWbSRvCT4iVRmnBMiomwhiF83y12W2jZinT4
ZrtCRW3lUzliDM4fZVP559VQ23rZg0pDIuN7Hwg3tpMXHRHIRSUkYrP5isgGEoCX
GpulGKVQW68ddxTBR1l9r5DqIDmqNgpoQv8Yiloz9PaYS8RVR4iPG9VKM3xlaq+4
BcrijOdFS9thKfOCC25lAprOwUGrlrc46u8Cy8gjUsAa5pMgdQRzLSGBcV5r4oEj
BTL6AiHPLSIkJsdzDJndXIPVlRtbeqVkl15io4Rc58KMG1gfCW+8yeK7WxHScOAW
g4WCErYfh6f1EzG/0xtq/yJIZXp7/kBK3SCUhE/gxwGkqCCpVJt4O99g04vPJEma
sya8FplTgwccxE2sr0xKrQgzzRtKqf3viBQ58YUwrmhpgXvHMTGZilN3irtrzi/o
FzcM6hTbuaFQKZr8I8IL4rTrlZWrmi5zsHV7ZYUIeN2KVehJTyuJmMGFwakJ3BUd
fL1X6uDlIM4/VuzlcdlSWi/IeIuGRkAnmVvtG73Zb59u4FNTccDTiOXP/9SiY4so
Wy0ORssnmFsHbK2Beg5Vkra5Cb/59ej7qlTmMxGScz5DO8nSHoqeQG32+OB+uyOl
TlDnObbwRW5ILoD5XH6DO5PktPqREEgwnt/zOUUaom1ytndtxT+0TEbKfdsYfIv6
EGACG/6lCU6fZ3mvxMw8lwK8aCAKOTwyuBmeLYXxXi4pPun9nvwfE18q0JJ8QEAt
L8tfEooGvJEcrrIfhap5FaDK3v/2na/B13HDRVUlbMC9fy90l0hsy3sXwNI86bxi
g7vz9ymZNQuBzx8ixbi3QrJHD7fSMq7wysWWbK2m+/q0opBLrkGoXhYMGkB0s8Zp
HcqAcMdKAM4YOPx680VUERIhddhyPzVDQLPZHuBKaflqDvaZrgOeYsICHAo+3YjP
JkGFhSejmLq/6gLObSY27qfETjS1a858XcZsa+32thUHA1Mxf88s7wFZNg30mqCX
eW0PGyZFh9V/cmhKQSiiMp4WO//H5dNvOG33ObYufBzFZ4lR6Z4KpaORfwb6PXmQ
ZMx504MhZU7sIgqo8+G3DN4OKvlnVysxO8c31+19nsQAeBBj/ZZJV01H2gmW9oFx
ZhEVGLWHdJBSVjq8xRCGtymPh0xX44vOfMtx7eyVVs4AnQ1PO/NmUU0v0Ep3vMrM
emERQJg0DMEZ4Vy7JR1nSSZUrc5wflTjYC75Q3foHcjkMRAwmkCulonqKIlO+IRX
nMKxJ8XQUumQ1OaRBA0LpkqDWo7YOsvWNhwBeNGwDmBKVNkKD7Wcmv30fnUzkhgI
MIDPXFYCiIrBIoIrEcFnWGHm7lvXqfghgkyiaYUUbllGTRY0k5ngrhw6rX3Idxoz
OG2+YZMySB9X75hir0m+KZOY6Kp/1CT1kQGMby85kpyWXxMp5THaPWX6b/Cfvk9C
MyR0h3E8QcgGDCjvAuzkfHQJvi1zk6wjlFk5EtqJJCbgGmNCAzTkrhJbGhU06AOw
kQEQ4U5FvfdPcVOku6vs2FSro8WLPQQ3cwgSVlZN5d1NlXuYchHC/bymw8JiRWYu
B9mvXyUWRX47WDLQPtX6B4EY+ym5YPgSgTutEYluBsIMqc0HAf59E/BMa26eNhBL
kSnIjCde5lNnvjFd+yIYAHfbnNKA1LnuGlYERz6xa7/Af2U4dgHVDOJSpCMHBQoJ
Hv/mH13I1z4W4GfiYiztWpuveNx9cYgyEX6wD+DvW9ZDMFpLZCBY0YlB7s77pHMN
c+DtCm0ydoEeTd+UCc1YT+hwt2bsUT2snUw9Wf5BArGilZmGYCvGSkGopgelW9ky
5sNV972aPkF+kXnLSjgjfeN//38cdA1EG8DUqqppFdU0AFChZIxRoaVZIpuoKhhd
V6Y048ZGXleGGUUPV+JLZvQp5XTs3yje6Vnl5ngP0h8xZoGtJw3HUKRpCOndEgl0
zhN8FrP8PVmBlPhYuaMT3q+YgSUIcu4Hta1ZybEEQ1J3S+l6jI9AAvFZW/fKT+3g
OcUK5CWGwUrcOVv45UBy3XtYU2YUj/q8Zi/Pj0XxeeKGzx+tbQl7MvljWZ6OmhQ0
ZWUENdXiuownDZUi2iAxi5XSXtsGSsZJ1cecZABw5vU6PYRvWmODnWdVVbN3cfO4
uQcvco4+y8NGAG8zJuDj1w3h9EzDcBakg4m3RiZsORVksiWP0GzuLamsXiTjN4ge
WoZ/T21LRqb9dYHhJIB1u+4/ZqrUeUY+cMsB24v0hYILklbhvZioycSRRIeWbzFC
b7ipYDDdyuMlDG9FpBqbx6+RHSl6cItLNB03rwsdo3GMKcwdcZ5ArqZjXhviKfKD
ayfSUtfxSV/WCklV7BXu0Qbgd45k6UgL8DMxXIpDAEdu30JEVNFm82gVjv4MiS2a
4HzKXx2O2gxjsltAHpYXbsANLo5WC5BByuwh7aXgpKWP16PNY5lK3o0iEEW41x5m
tgtyQ++o7bjrgi8ltv3i8DyXHdSQwFLYu/iM+Y4M0LZDI+kOBRYnPePiIlPzsce3
/V327uCAViO6AfsWf2BaCyXGSV6mGPhpUw6g1jjbTzbnmorf8rHaSvQNFcI8O4MX
oM+AEK8/s/4v1/9Pwz+MFAWKFM0fB15NWSMa2bMxifUeAc0eI1AbloZj8pgI90gV
eWE6ly2bdmZuIoj7KT5I4jdlYY9NvLIGerszIBW2yE28I+D8uF3mnli3UXV/81HA
yl6msS9sR6fBt4+KBr4CHjb0Gn5LiPB2HqKVUdNA8p8o0cTM/LsLcth52Szoh1HE
Gak812bp/TlIqEEGT+BkUeS2wvVVGBIzRLPNUsVznrbGHKyttBbrU90EgFXYGTxS
f7NBO66+OkHxrMMKU/MAlwKLsEz7eSQAj0rfVgUKyItu6KriaQTQ1oRunoV/bk6a
866TLQD2W+/jpz9LTJgkPygPvwkXIrulipLOe1f7RwoorP7ScJJ5DxxDg1NzXvNK
Wnf4owy9y6qUPJId8pF3RX4D7nD4gN+jobMmN34RaHCedUvkfgXqy2bxufigVUEE
CNIO+2yEnBBNmB16hgQ1BsjQLebxlT1B91TxjmlgCOW07qLvW0yXBYRF3dtelyFP
SktCriR4sYHS0atSzjc8CnV6V9IxVT9IDZ/VSz0mqZoJW2EldVzmwkcQwuhG0V4B
Pn7lpLDpYMbqW7gA3TaFq4/ZxR1UgqdravhR5gcOKPLVo6W6HgftuWFnr1Xo4/DN
dO2KefnJ67P/Q3DQfs2A1UIbquyRJXevzWgfPGDHEWMZp4y7V7vFK65cMxd5UWY0
sRxrZEso/mk6mgOnOJIfpbBjty5Zci5A1hNOpwbkv7bpyEzr/QFIGLTnzWwdyS6+
B53KVpg18MKsIAIWuaKTQmvjCvOCIa8LQUBxEXAYJZgnlqBzDMkajU8Y+qxSkHUF
0JM1p1rvy+Sy+QHYRVnb4XJlFFkGowgh6I/rOJ9uqebyIObw4JUjfBSsA9CBEhay
41+nYleF8ZYomdrp2i02+3wyRpvpHPsZUfU/rQw2bMlpbUUh9DYzPpcpNYE4sA3A
XyEfRlohcgysW2Jd2+mSIhdxVFb3/HQHGE0jNt6+sN9j2DglCBAA+4sjZvmwjo62
qoOi5NM94g11lfn1Csg5wXY/GOzQfXW0GOF6k2UzoH9Pky5jRYJTFLArMfQi1p5a
I6+WgnGrG+kBFDE1u398czIsVnkbUOz9vYcKkwaFhxUbbVfyisT0byGfgq26avJr
cGM/qWMQrIfckyZHqqCIbkHvctT4iF4uD4t5WRcToWz9tE2NeVNK9qv/Y2yCP1L5
xdHZEhN33VAFsDb9Y81yaUJJFgyR2KkKjcEIILP/0PEgyJ0RREeRUjP1UyzqndVF
+WIYa5C1w1+T0TSwU8XZUgeRV2G3gxWOp6l09PlJL1jYyiNmiJUjRawfbqlt7yYx
WZHuWke08tsxr1/arWFTrOqW9SyJy6F/lPU4pBuf3kF6+mlWj18exsxJQKDrdjcu
Vf8/CivGFEWmQcgGjanWlsgDL6iJeJfLCs/9ZrtUJERhp0cX+7mL5w0FApU15K99
Hj/61Cpb60PqgSqVL6jtkIco+iIxlSu2cJsl8yIcEtket+IOkVpr6gM8yeHgIiPJ
K2Bz8l229vXQVum3EhmDm9ZvBkYrwdEGBqkeFA4Z9AXuL5vrVqYQMrJ9PpxTa6S3
JJ8lv7MoYF6Jail147dPJfhuqmn1FnuHxoOs5Vd/M/xPOZrb5MXMBI2b0qweETM0
iY/8SDCFhW0FadoH39+EacDZDLv2ADmslA/n3VTCTkIUnxDgTxIyn1NUGS2tCbzU
RerLS0f7/ZUUmvJjxP44RRq3dTIAQbWV6oKL8qiIOeZRdAI7ubK3k3+9JEzJ+Psa
LS8QV3u0d/9Mqv/NAp0xR5LM9vaBjOilGkaxth3ogMVIngjKQ+dGS8mF5MKMl8G3
P61aaWBQpHMpsDA8g0J4nlXkMgsHUyAfBm4gK5cQaLNctYsmqJuBSfe5d6SiUtVM
it33fhzzaMKrOCNVHxsJHMAqP1eHMuQhmIGq5ofBwFL0skc1jWJQxsmFYJ6na3G1
BfNEWFRigQAdBJ/7ylugGX2sj65sh/kjlc/F8iaGlJlg/945F67QJh/L43RdhyEh
6lL70H6d2BWwv4xK36fkRtaabghrIdz24HvJZHvSsMY+BzRTH8QJTZHX4AtVkDcE
iG5JErM4p0D0wB/h1NtDqmvoZjpmyfVMIAUfEs3byOFqTxD24BoWekR/b+krpQXm
oyYG2OVraJXj7ihDJCLfWv5yUBMn3Gv1Y02eM/bdw8oB8ZSuG99pialzNOwbrVBT
0qCUuP5PAIFb5txIqEIJLigTS8tmhyRyFrNXnKCK0INlGoHicvkUIdphxrHZpbZp
uDEjGspanC0e1ae8GlEi9JXPKpE6U2iz+xQlwwC+oZ/PkwuvOrrtL5EN9973Ta30
L3QKPo+lMHMDfUDgGU1Sw6TGLwOO11NkFfPi/XBhyxBZcvdQ0vhburx3CswwRH8m
t6lfWHD55jkg/eQqlBsOWmMf8u7mq6VzvBF1aLwjZhNkarAu1V9Iq1aKdAt8WHoM
VTqLPnsBpSz7WrJARwe16cnLw3k/ukXycgfa0NdtqXfWLqRr8158PX4Pl3JHKvOw
ISlv/0y0nawZOc9lbgtlFlXKuDtW6HgndG+4AG0jn6QQH9ysHCg8KiMDWkuwfU+J
+Z9Fe9O30GQpSXzBB9BnAlAIp6o0x5lfsh9Wt9TVq06gRzo7aQy7qPb6qKlmpuU+
2GSD0eVwmgVtYGIZ8sU/K6QIHWH8julb4GThSnipo7ia7rSKIUugYkLlO0F9srZv
w12w+rrfMm2FqAI3q2KQtNS1PxM3p5RifGfyvqNz/Gu7H+mw7TvTRtvG40ErE4df
6YEcIMFr/N5QhyEqL7cUJLUcl9oCuRhW6YSNp5gZ5fSFRfn/yadHThDWjs8J/ijY
WPUBeXZgYZCAhnDPQtSUe4zryn/n2qVfhbu892iMlLaqqePMi7N3q5gM8Xc6L78a
3ai8Ak/vxhAuzN29tXO4zocXTwOjylHZwE2p0lr7WcuF2zQYnXQS4KXZ7tmo8eHa
W2rzymSoMFIOeMaxc/3AXtBb90fZa18PnL+Qs6ZNv8WxJhNXXr0wj1PkAvtT6v9T
m/NyquNoTj5x5IJZMOii2F4kdMK3ZEXug0QhXWvWpdqxdcaIs03llWmBQr5wCPID
hy6O2SYr9F9BHlTO+QiMCLwfLhVwPYebToaYOAcdG5Lkm1kv1DG9DcUK/n6MjHfr
Av0itI7kDkHwmTWgoV9H/udzusHNwECB7yGxBP9RjufhuWlGoOXaRoJmy2PRvFsr
4c8bKeeZI0NhCrBLhvFpWSi54xJ9GHvDs7Kql6vuBXmY17k8DRC17WYx03JF8SNe
QNspg6ceyBhyck2YjyB1qyAbOiOP7qYq1J7A/X4IloFPTom8vRHdtd7GDD8tSmE1
k7BvAJIRr2uzfzIPuz+0Giz6KfyMQ7Iy27sAtPtdlnd8appXN166o5whZFnLf4Ek
saHqP3RTtA3NeXGLX9pTdvo3Vl3MbljmuETSDxiJoYdcJMOrqfaUrEbnJwzWd9LR
ApP0kOOpc27G0ngNhNQwgC/BA1mWN/uMKfJJYVMvRPwCtC/jehRLFPyDbdmjgQjO
GwbWqIacRsEzglwYHbV8JDvehI6ugw3bA3VjarlWLDgnooSl+6Y/BkIKRug2JgRS
BtvolYkX9RqRolYNUGrcq4oyDa/1nfZAw9ZexVEmUzAkhnLpitmszgR7TkJmO9P6
kC20cYW5Y8HC3eFKj7jAvmM9hmHp22N5hjH7WjpuIgzLjjahQaqOFKw/kPajlpCA
nBx0LgzlNCgeF8jty77eyPozSA/rBvmPK+RliDwk/25O9glhHACN28amLDYlM68r
2HW2Gxl7MW5SjKUVszqA9HXfxaSoi4VIa5ztZRT1ywNYu2k/OGFSKmqMdFWL6jFc
KIPiK/g24ZVk6QWy/YVe7+QYIad2guCI1jn7mBxO/L4ovDSQX9HPDm/NLd1rI2K3
ZV6IWuYC7I9Vi/TdvIHILQ8dtfdwerkB2JJJ9JBxkpmTlSgMxmE5o57zhherpHE8
xjT9uiJtpCE6grgdz6D2uWT/1Y/KsFmdfHFD+LapPF5nZeHi2iF/V8w31fyRsJSB
rTefFQE8OZ36C+3ysOiQBIXIZ5mhy2WU1lkNtL2dydIfFWaI/kiEu2TxpKRaEu4J
sDKzKsx52RgYOD6yqaeSlymBdH21j/6nFtA5V7ZU8zLlhrvp4yVvFoY/Ndh8vcHb
vB1/nZ0UXIASCC00zPP7tHM4frDzWBKRJlzSRseWkwmaNGwQf5uopXka0mR9Zkph
go6ztIwrRJIf1n+JvHbwYtZnxqsDIfP+Mp7vlKC8PLSPmRp5gnlWpblxl8aVqyOS
QOY2ts/T+Ntcrqua7tT2WoXO+U+MYecJIViqYGi4zmCevEXPdgjcUGG5cg4MQx09
Up8gX4AqD9RFr0DSDSD7Zgdc9FgzqpwAn09wPwl7v+uBVaEYYTBKMRnqBQbRKnbc
x+SuwiTYcDFBNPOXmcRkgsWVd8zdnRLwJPaRW1dgv1w1zPE5Z8fwr0+j9tkAieUD
m51pE7km2KPqfyITkwifjgjYTzB7Lc6yBCmiUSXSZstVJSCEdMLdNdyoCFpc9/UO
FIMRJSPSRkuNjFhcyM3Qm/Y7Rr3CRKoCBLPwM/T38peOyc6dd6+aO4UN34SemBur
OEBMPgGrl1bUNx5EDqn2EboZySrLiMmLlWgWBxBohjIHVNIf5aAkYCqSpX7h/zuZ
l1Q3O5J0D7MnMZvITJaB5FzZt5xEqYnOlrw9M3KPPQXI/F5xVUi3W7Zn3eqkdnWs
UTh5NG+siUth4RH905D8A2q3WA5EWnZKXfcUqmh1T1FMLeok6yTyTt9HYOH392Dx
kuCHbf5ncJLj7oGCWC/btJqDCFemHiexwfH9mBYiXmEYRIo+LOcyQlvPkEjkMjhO
mq4eortpIojdLkejn7C8YUQMFrC8NXDwno6SQBlzjJ6P4PE5pUaaadGqyKikPDdP
2x69QcVA9Ux2qqykXBuFa1dR83QNRej8GxDA7HeMilpFTOM1nAtGEodnTyihC7aO
RWfZeq/2ZOBV10FRGOgLiygqoj+vOa40KaAsPLjzYHsIl2QROGRjdq+/zDnCqCfy
VlsrSmgmjVgtV3zTm3pg0dST5a2cdwgdELyab+04SRi9ZmUKgIVD8GgQFnPHFLy6
wf1ZjFGZO+h9DWbiMtLF2idRVjroz42zEcxnUO6oINadcnpKhi3Pm/Nfqm5c8eDv
t7sjQ1Av1RIpjTkalOjjig4Nlkgfzv6dnsBTOiM89g4f1FF3cJg6bccSnpmVviVJ
ELmrg9+xh1k1FAMP+8/f4GAblRnsHpGAizdwCZX03Yw4PGOp+nTSK54+tsNoTnI/
d0zRxRKjSH352NoR8rBE3E/9hhxX/nk1pUSeDgY5bbHbxlhzEfNUSPIjrHMCPVps
t5yKhNn+jVPtWcuNR6pwwlzm/jdSs0k/7K7A7J9Pjof+xtzFBjuOtXjMc/kJFk9G
gsKDAgXJlfeJEeCQjy9E2EfWal7hH738CGIwGSY8vhiS10KLllgTFCfT7VLNMXFL
1PFWi1yZ07kmW7oKhgAkpmYFPFNNXC8RLvDK/d6B9fd0cnzx3v1mg2Y8Lt/U0xu8
H/2HwAb1lpQNfLbQIs/ZHRE1oMjgtd+POHhNdFjDPjlvQpy7zgHWYLVpudP96xr3
5siJIBfTcVHmzTlez0kJvjYGjOL9hdiVchJCUj9lwkf+qdS8ZFQE39avZDSVwgHi
oqAwA7BR8YXQDWwGq/KMi3Ltr/Iw8uTn14Oe1FAf0BC/nP69ZhUv/OvPXrvgfJSN
Ku7h8cdcfgNF83ZuTw9qltQv4iYEW0BO0ojFzd7rj1jzxqxjEXygkbFBNNUvBF1R
F0qv6w4qleQ3YSR9efVY35e3BWQeuCm1HytHsFqPi1lojgS92efz3LExXhsVRvUZ
7tQSEWwC6dMuWq2ONqzeTKVcaqLpvII5mKrxaAShdvFkyu4KmvPE3FwsrjQcGKO5
HOAKSEbC+qPeP6QCSdI9NykRLc8WSNTBvdC6hmoqPAxY6bYoeqONqsKkOf9wSFLS
zeHcb3rLlAl1IHqYuknNhf2baaSsEUPO4MlB43zqA8gjpFOzQ+HegeCJdsWQAjRa
VK3PhR4FqnC0/8T4Ir3y/kyjwVzlazejC5hcUXmcTSvuKY1GuexVr6ZakDlNHMpP
FBL4UJp0HmaVsIcEOJyBWAunVBuOPVTH3dZmqv3WqwwoYkNYQP2zWQLt0hsTU8qT
fA+IYoeTgXQ53AkteYOlsiMKbkTyn7Ac922KsRN9L2yZZTKOxytt3K7mtjvwl/H3
m6vx/FvtepQ9spqLGrz8W80CdvRMQsnOEOfmANAYhB8b20uuQ2k6L2Xrqj40Kicc
iMWmuF5Q6h/nCGCTYO+tZw14Ei3n9lct1oGqlAvMUC/+vvn9lUNYoJ57RHyTAXdv
kIY0w6FS/YiOSvQDCsff7gPc/3x6cv18cWn5cchpF8KhUxKQrw+sjS0O9FGYYmx/
Jdvug8uQATxB1M51Q3q+zXw/D2oQUL1zT7qwJFF1LoVBACdM5LSZhhf64Datg/i8
/Y1au+r2/vLv/zus9IS9b2I1YBe2sfTpkctKDp7jzCiIrkO7mHP1rX3HTtiuD2Sr
333+Shn1a4HIP5qlBXBjbfpVmsdqF/t/4j/xvyn4ZQKU7aRtYzhtJTCBsKyuMh+o
X4bcy0a8G74Cb3OBvQQx3W3/V6jh4nlpIdWkbmE+kFUAM8R2y+HLpyOcyJ3/SzR3
clbdJkgVNBWfKntWPxENLT4u0b0x0Ct3g15twieU8PZUAttb3P9b9XHcVFHqI9/g
Sjg+A8nkRpW1FHclgiIws5PT5/eBwwQbIVlLY//2cRpgj8smsq60aJpW1Xpftrbl
/HAzM7xZTZ5QPiJM6wH5Eqzb7MTorECr/Eh7Cmi1OBIvbKNFVTGrN+8S2jz01hON
b0g8D7Pl1UA34xOSMbYbCCj/HZPv0RBbNKP7e3eakMxG3XhrhrKMtDNrsXMFbeK/
VthkfZJOuJqJMJ2bS8hUC8T+nPM49KntLzTk2pR1/ND1cbY/meMBB6n51I1nT7TB
eKJTjOqFY6959oCLF0fl65W7o50vJe5mfKJX+DW/Mh/ZpC0MlEzn0Mu4zI/qDrLu
Z0BexS9yEBAPRT6WCa8IIcnkbPoXWGaXJhaN4cY3YofxKw4fIZ9bQJb50k7Ha6xI
aaFS352sLJUA8+VdwIp39eyUEc4Nbg/KKCmK+QlGjWq60lwRNOhIR+UE++OY8FU7
/g7fH1J31C1JlizV/tVS/+2ex+HXFPlMXLTFPK7NjJuuscE23W8lfuMn6X7modj6
+Jwud55pgPDx8ReTRI9CReGM6l7FRPfPuZbpTUCnPUszUjPERMWs6dUTJeLlTi1J
gpIJUMNEMmj9E2odZ94q2nPdjJskcGn31jZuqz+hs6bw6oLIX61BJJ+Qwui4KciL
kRXenEnkh9FAAEqpKNrfcN2Dj3sJbMbeA8sECuvHeInYjh8W7hogHsKfPfwuGz9m
N9WUzyEKprhn50MuFYnYntovvNOwNeS7gr/djcShHLn6/C9/VFvDE/fLbUarAMCe
jKgov8dkLIy2UwzzJjbgfOPY2feil8dC2aQhe+Y3JszkQFhS8NiPQWuuT33MI6G7
nNgOPR86/rGel9ISpvYDcEr86yrALMqwecfz1nu0kPoxy71DLrOeMecVccnJH+B/
PNF/5XB76N1YY0ERB8J75syLavOkYNfhfrT0359UnkoDe8O9RJSY3e/SkkNBZ45I
5i4y3TWUiNQJ3QoSSMWvUdR/AsoVKvBb68HMgJ65MJdQI/9Px0oMOzkoTID25iuv
bj5qnPfeMQRyZPC466dK7aWcWk33/kaloWuwFIr5WXaRUqiGjnQS3WFU4C7VoWhA
TdC6OcrYhuUkX1k4++YYcvTwPOGXb33eKZVotSsZan2jewzQZJaUza8D9pcS+kqm
t3fdhepC7/9zU1g47DjSAYAcq1zUUDrdW/9SG+2/SSWDegAu9ccba9x0JiTgp9Wc
M69bg0aNHnYSEEEO/etmxEmTlXAPNXhomvDss32HVwY7AIgLR/aSo6LBE5ElCIGk
7DujYDOgZhhTEmj0CZyd4Xrf/qsh4mjYO1xqnFmvvsWxbR0boKsUhuiq9SyCbZF2
2Gz7PkAD3OJpr9hn9foeEa2ppCK9uYK1VIl+3x5sDmDHQ5w8O5WpBoOFSMSiYEK0
61dmYlgJIGW2CESoN8LSOfNHFCHVL+BVtHh4c5XzvTkC4uyogOUXs2AYgx1AuY+e
y6r+WNbiop4c7x0V9TYaT75dNEtE92kaldtNfsDk8bc4DBL7IvhgmpvAKV/I78HP
3QJ8OGe3GBNghnpya6ztUX67UCD+C+Xad+ptPcWTYzjtmuhnxvduaP/Pq56ahIm2
zFPGfMMzJRCIhcTcnE09tMU8u5cFxK7JOHTF+u2I8p4r7tk+uuBaRrNgQTWb2/Ts
pbEW4IvAJUI+9WOlDwn4Phf7qT2G2d3K8Cpuwkei9D7rQtRqJHmQqogU0UktaRrz
EFDsQtX6CLbpHmY4MiuAw61tv/kxvYxEdA1WOo/Muikp7qVK9mR2u+tdWQl2xmYP
7w60y7AHskAFs+9/ASsTyY8s/2AWXALCCYYVy+2lu6ZmV7UTSzVarmSPVkQx7cZk
ZJLifDAD76euxDoBnPKzyiUtUnf8uHdTc5sWiwUYJrRfJCZi4XFV9rGpJ9hp1sC+
nI25MvXq+0c9lcodFcUHmYhm0S9xcEZIsm72G5fDV8owuBj1p7+LVL/DI8y6PUBa
r9nGDbYzp5rvigzprFOEJDPKFN3iFJhSUa8C5Hw/XFcRQW09hHQB2IZcaM0WXHHL
IKUrzU/Vtdr+i+DTMIh1BArKxX6CPl/9dD718B3emDLZWp9HkF9kufNkWZ1DfUFK
9YpB5XS2Wxl0Lb4OIhs++l6kCUW/VNHtbuYIl851BFIRIavp1HQNuUmda0dPwRLo
6scAucK5hKW7Yy8CqQRrakjDEXKgO90LEXzoUQBiS1HjjDANe9bjKMH5fHKhDETk
guy+JmWZ7MuGy70CQlxynGl0TfSXUYyPVNCFt/9bQ5lvExl1pCGWGZVy3vhcWorJ
nDsyWqEIzVZBvRz0Gfw4MD+hGDT9/NpDGKyofFC1+fUBmE4gLEe3k6abQ1tL9r2N
t6Zpwmms9VfdxPL1LkAoYxxiGS6y3IfRzcTImHWaHjUFtyG+JszVjpI+9wCZiD26
6I10uxKWip1pIwLryw8Ovt+0BClydcun7efvs5YCOxrAGvPlsM4yvDznvTMYV6Wr
I15Ko2lPn/WSxIZHt5cfo/6pu2wfcrWZX0wA9PZ9BvnG9779icgl4GPeblQK8AJm
yxaBhvc2cmbINTVBQZLNnYHJgHk717flvXDE4LDgQpWRLbuVg4ccjv8PxJOf6LSJ
Ert6TzeqjzgO7BkVKkGal4n97V82IjB8YAx9iNUpRe3xXI+IlAcQS91I6ex/+mTw
VhLSaSQS4CHQkJ+gRvkr4ZESndmQYwiEZfg0SfOKhQv+KIi44Fp+FU0vi3EtS6nz
bgan52mvis/b4DFHOh/zwtk78AaCxvZ3feyWh4zXdNsXQiqJIKZzuAg36VWoH1TI
k4yLmOFz7xVF6Em9+934Hwiwo9r5xG34ATuvFemKViUhZBk2Jtp01X/RRAZQTtdr
DRifTgxUQOWF7OkuMk/e6r+d8muY/Im7BgW8wHqCQxgqgjjyX7hbDgx/AQDRWw5e
1TRBJlshSsbNy0lyhuHArMLHWLxNkKj4kM9bQ4FghFIaNIwnzc8tJ8amSDsB6ls4
XNfi3+6ixisHo/rrBIlwwot/CGu7FLqXPbD5bQ7vnbe1CD3Gp67d964A9IRY2QPP
+Xi2XNSPbZmFcpYq1XtEwoYLCp0ztA8ScKX6Jw+exI/lqvWwTwF1yjej1mMXt4fI
HEDJ5W8pnB+ZM8emI2wE6NRUDtSxMcDo9PXaEWYs8Qb1FOhP6LiipjSLomroG3x+
AR3RsCIwbODfWPvee3R+fciUsrdhdaSEnbODuBCtJwROTMIgf8BJdFsi/spEGgkB
dS7r9z7I73bIgRWonByaYoJIGMo7UdRSUJjDqNyMLan9HKmfONcwz90XClizYCeR
C1ZjmXjg+hLIsQIjNDY2ePThBQViF0h8bwFdS2DCaDfedI7Mwt0k5JVqzYbRSOYh
7E/bbxZb/5AsLQbfGNYfpfSTdw+NTXIKm6tcwPaa1CHKc+D5+UIRJXi7YGJSpqtX
oY4LgnsFodfDv5OGyjGsMtKJMs2hksjj+g2FCM853yuanGDC2GUv3lzKGvBsrrCa
QfzpC+5pOkdb9AzUzucyK7l1t0J2tvBmcWokn514XUcbkISH2hljMSW5Mw67f6qM
8ZFzkSkffyDOZ0tZQpfNzHY50ranZlEQ/Ml846mJswnkkBSgDnFylERuGdi7uZnB
Vf//ke+cwAgmGdtsse+wvGDJz4yxzfkxkQPIa62Nvkn0bjyU2WzPCaNN0xbefz/N
qhVkEJniVU2YzCgQbI8PYw1kUQ/fQjWjj5Q+8Kov0gkbIae8tIIDL43+sYOgL/qN
hBV/OH8QANwPWjFhrPBAe3d2661XkBS6hV8SOJ560+LrlTot+qIj0NX+4Gy2DsgX
2byH/Er/8/vup12MK25iN4C+1/2/kawq8SyH/QCK34lUMT+afeUn4xHVcUM2CtfM
fCjBGK09MIk3a+kRbgaJL2SQQFT2qs/KYFgAKYo/zi8NZi4uJlOFUan+OM6VAiXH
ZS/ioVh641oAMM2GX/pQ/NAuj2K6V9w1J245s816XF69IOMBksJXAGLYdyNwKWdN
gkZgoAxw3xAyx9DCOt8PY9IKvn7qweXvwKQpYQFOmW7CQul7KAkUvb0kLUuPohho
tyKn+0BcsfgAP+1z2PwZTmnpJsVQEmMF4nFDJ3uhlGzjQS61WB0cKw9o/v/roW9b
/saR1YQ4SuIqhU0JYP2G9UEH44Ixwjx33665r4oLRXtnMBnLCIpAeUXp51YHOFkV
FPjj3nWReLXMY/k6qwjdUFBi7VhNmyDgNAK2bXXyOAYPO+XmnHCQgY9KpXkejOay
G9EPj4MWR7xQMYsuCVw7uK7F4PnE8dymSrA0j+b/4SOXJDRLgo+0/ZHtN86mXFVk
y1ziwY6UzCEH1AKLlTH0/kwX4NDvgvEsDyPic8Nfec1zoLLAOZlh68xUrH5AhDz6
nX12gcZiLxsFHZc6KfIE0zMI1ocD1RkQc34WgEJbrBsKRiNXDmNZtksZ5MtjtHXg
kOxpZiJVbaZiYp3QbMZFS6CdWabznOf0vAAuNTqVWrP1tlz5sNC5HjnHDbTuA7TQ
I8kHZvkHSDLe4VJA/iroDv5PIKCgHnj2y+Kp9jZV2ZAyrTCcKLFvqxCE3rK/N1N5
Sq7a6GKsLMJ12UjqlVt5KJ9H8a4QfrLnvTG6zLx40O7O7BbKijJwFLzcJN1WYJSd
98tZ1cBKmvQhBJSpCJM7xkhmp0ZxHcXAyLfIwS5mD260kO4eeTWSH5G47H6V7Xvx
yW5HpJqPDjqCmF7APJ06spC1TUp2rK0bvanhoOucdMK3QppnpANAw/0RU41CpymK
EarQT5smJE8KiYDLMwR7JFF1tB0/1ScCMXelYggbUGiSHAp4mYjvKoxff5kFMNXX
g6dDbTdvWzZM+/B02jFwujaH4vCDFZvlNL/7DuAp5oEi7SZuXfwNEoqHukVRsgRg
qoJAHlbiTMiwa9KxjpRa9bOX089sxyAmeRRtNIu43r8QehHIJ2iBNXOIfczcS91R
7mmICJrhFg9cTb6TUtGXc/Cjr0lkh4sKjtSkmg3Yv/U0wKC3JnPrrjzZyUCWWVrF
yHdt07DnqTU8gUJCuTIADYqbgWH6Uw0JsElIQdqwXilX0vUSJ/lH1ql60uLdqk3V
MEPB3l5awwlc2K3EKSLzJu72pJnIZLzLB7Fzs3x5+cYNoGS3TGgautPyf+95Ndjx
URmZyWcrZiQrwm90iSQWtrw8fu07hOupg7P9tFTbUMzLockJXP5ToSiCe+rGr7uk
l1tBiGskOvz2v/3oaNj8u3z9iBD/q/lQcOZlulzyiELGwEGfETiOK9SdunSPBXLq
WZlE01wlaPxFtotrJxYUUJ6XSltY5aTowT5BB2hiiXNOonEfiYfUxlNmew0qfaWg
/LOSeSwvve9uiPqfpLomf6/3oeabsI6FRTcnblv+ROfju63uAL01cfKUv14Tjw7G
JHrxEiFFbFH1w1Wgu6nkV1Fw7D/qdUS4OPvUxCk2LnyVKC2fongFtgRqjsEgrF8/
9Jx9DmqwLM7v+E9g/DErmYDQCKtygNBvUeHz8kKvh/1LEPmhh0IFc3tucwh4ErZ1
n/1G/kG378XpESV1uFMGKQHii7wctuajS2BDWt5Ih9VOHEInUY/27ukHVyiTGAfF
2/0jfvyPzIbRdDOJQOxSkAhrrJlZlRFxV2nfldg8i7QT28gk1ULVekUYeXTP9xLw
Vg4AKarwNRUWAqslzX41OzLpJyWUq6YuL+YekE+AqUQR5kPxYKzH1Ik4Rd3BEAjs
sd0tLsXd0yeJyD6GX9THbWvdrUols4eR6nrrJ3y+F7OpCPDNFFKTFMHFgv1vrpZ5
GvcZ10lGp/iQ1xA7PjiW4FiKD45zTwgVX/5t2qmLT+YKbFgwwXqHRHWBZaoJpQFV
K2wMvWF18g2tpf+7LcvnSwzeh/wgdG+0lM04Uk+OKbTkgIZlzjq5Dbox8Ca9tIbv
HSDxfUS31d4xdJFU2juaMZaK2XnULIkdrNWpi3ymtMgNxPoyKKNPCLoX2gyn7fU2
tIyWO/tY5EsdKqrurlIEo+pkt9wOIJ974hTkX0idHegzJyZdY4xgwDdNt4q0NoRt
ZMXBTQclsuA+Jc4qM5bgQusjPvmUUvedZ76BsmwJvRTjeYFiF4idNtmDQgWlGR1S
KEcCce540YBYybdIkwGm9HWxfWP6UxgW8Jdl8/peZqAMB7uwNQ4V2G+70AIKiWr0
MyP/v8bP2/uVJXOFb9QfkXVTDb3AQNmH7lmzOl9jZAwstCdIdHu/91FcNJkv79/T
Q4pWz/MLyUG6IS8dq5ITnJi1+ExTiMF9rkm8d0DiKRkE7QZ1QhxDmYMcfWmIwMkV
uri9U1cNV0RehXxVzFBPnwBK6xvelclId1CGWCWCTzhXtWV1tT/sf7eFRYHLyvzW
L7grRkQ7Tw6BeHU1dYR95YlHG1BNqU5/UJnF1799VQIhmREbNuqTnmZEdl3oqRjj
vs1USfVPOYE2vnYoilkpo1xRC2uDeOMGoqf7Pn0O8T9KGgH23PQMD6CmW9/I4Hm3
jcJRHxnMaZwHA4sUd1ImQNx2QL81ASDY2+SEM0C3YWKgPDgQgaPpecYvNDc+v6sw
x5L20HwKULPz6z9SvIY7E+m6uCbxByQNnvw2QJE20sHnPyZsEO1EGjjZKJs5S8+M
J8kAvd8pv4fCPi9uVfgHxxpm06yIicg8JX/WgjPKTdcD3FFjuQokE+iTS2F+kQsV
Sd8yRY+l/a9yeSbR56ZnFJMXKK1fB7L5CAdk0StziJnc7UmqNZPCYXvxUzjXixvc
8KEKsmgRrv4xPNBsgbqZngfdwtqW+dvP+sR0istWu47x+uPezz+EyeZYeB8NVHYY
7gvN/xNi2+klgH8lBh0tGc9V0xdwHKMJ4QXxq6os7j8Lo7Zq+G0Nz0mTsjc8i/ct
CHTwYsAgH5csXvKnAeuZmI1R3KDhtwI6HPI/rMEPtVprQZC83oNkx8stgrOz6ark
KZqEuWXzXbF3FDQhdz/pDV2BAvYUobTFulwktrpF9shlnwiaCByZ4pTqsXe+7jyV
ptkC3KmpSFrQSUBakg5n2nTDHTB4esVa8UmalY7BZL7t9Hc+/4OZDjYBdQfmfnvQ
tsoPUqXZ+d+T5goZPXB64ZKmpUPgR6XS0kiH4Bz/KhNvYuGMenOXtpAEHL2Ip02N
mfG1pGzl2QNSTXIJdFTZIiSMEGWTS679ukYkFHCvoG/B3DBuoZeu3eoPoWSzBtnd
mEqzZDGo0zaSWJ98Vel2u0zbV+IfNMuiNHawxbtD3+r+anO0oqEpbp1GVOV+Cpdx
f35MZxIRrHwunqh2IbBJ6idgKyuRgSX/GMYV92HNTETgdRpl8iC5cUX/VOP1kSYH
PHE8Ew7S+0Bh/mFkawnsRgHSOXc9cQn8uDIb8L8xn8eZRr7dxB7iXhH0eZfWc6up
GXC7B4kc/fZ4x9pZivuY4aP8fWqh+7YNqk+FdkYzi+uVB4Go4uvS01SX/seKMV8i
AE5L5WTyRU6VGFXSNIEAXXb/WMDmrW3y4VVF4cWB/BysYhGH1MCZSgqy/fqP78/H
FaCfrck5UkWlpUiUmcf2yyAk6+sBMK+yN+KP3Kn79n8pyY/lyterYdquVjQ59Pr6
G4FOclHtvGMoA6eWn4Rt9x3LA0vR8QKliNQESac5k5t0N84k7pGTnwFZoO0kQqbu
LHo0MArLAv37Rx0DTqzqPChx0+85ZXxzFye5YXQjkRop1rSACgKghCIxKm1fB/8D
okkbv2fOtLMCqW1nCsstFo5syPm3lfr2VD0osI0AN14w/6GLHRdJcRstmvOVOMa/
bvrodczBx43ZB0IGSSqbFUT0jlkzD+ngGznJmadVN6TDSV4tjojgfOGKpNGkwtCi
5RIXlxfFlE7G7omzLIQkz0riiBUBDC9G3jNc70v83EIun40AZRxGr3+51mfie6GZ
5FhZYGZI8aGjFqCLhzdS+Kxq7QeqO1jILUptDmIu8UROuO0Aze2dN2nnM/6CJihs
DAh7qdd+WTckC71IbxPMTN/pNxCq9CYAOJFMR7eq20m/LFoE+rgghM87M8XOHlBX
McshQiNDad97g2BsKth7O28cRlgfURnjTEQEJ2TfXTa5vAkelhGxgwUFENt4Gwlw
tNJ6kl0PVAmRobeHe6c9r9VTw1JjstZRSlOKqy0kz/42HcnecH9Vn83gMnTdJInq
WYpZX6Cab8tqvNe/m35aer4gXnp41kjOU5xxN12mrjaCZAGAmnzdKy+92ZNgBPo9
UHLVzio3qS4Ka2P5BG8ipZ9M9e0DsbwZOAkUtVYGmLw1TfvDdfaYWD6jOWZZBNub
wGPw5c8++PWerHLs90hodO2Z8Lj0LEuukci0Psvg7qJByUc006+vT9o3yEtwp31a
u1B9Ww8GE1B9zoQnRBcV6XTdvNF4YwEhAKh7WCIv++6AakE9aCahfXa2LY49IvN2
MforwFvUVL3bqSbDheI5vTHCnsYwxPkG16CrzSgpYP8cae6scAr4tbECOayyK7Po
pxwjtwUkeSevDQK+/bvTLU3LSGwZgMA6QI5zb+udWr32BlNA5F5RxSFGV4q9nsFq
XV8gVJ2uAumJaHecPm1Ifd2knbWPILjzhyG0HSCbrthVyDNUKa5SKcyLy53K94jF
aceqICt44WJVzFnFrvXuxayaM5EBxG/NErRusThtX+4pwfUS/LudhsaTw1dssERB
JRzbOxUlLBvTrroHykoRHXfQ9nMcq1QBWXbHySqznPazYgf6ycy57A9tfoOdsuZl
5bfIT643WPPubmxHtMFfvTNMOtGqTvWeaCH7rvYA4Lxxo8Np6ad9OFeHD8cL+7mi
Dc/dxS1LbLKo8AekthnjqhBIBuwUYrnbPgR1KlCeLIJemwebWt0d+xToSmSHD4hm
bz45PdZVyjXi2uE0wrZaqzjF2mfcGOAWe1yLyn+HJlNpIkaw63QsfTTLqR84s1mt
xkDYsXuw9+yWqV4sLMvmZSd9VMUP76NESd09ImXAjVXsUevm2g49kSwZqPsMb7Dd
e+iDmDnOswwEU4ApCjVKSlBsUrrzUCQsqf6HrsEA1E9woW39QZTPZg2wIsHSZYAs
NnbxDYVnZfDIJgM3FItUv1+TRdrVpVAV3CEI9OWmS4rC5Dd8CPnGv4k/nXWiu3Np
9R9AyVxdyGKxON+P7IhMDhl8Rp++A8qOxAWE1vvCD1DLkRTlm8zwxQ7W/17HAagP
5YDbOXXeIvwWhVs7hHGT+XTTNCFvLMJS+6oh9LRBeoacXCJJhEJNLl8UmTenTQHN
E0jRskrjThJ6g6FFdglb0Kt3xBoZ8jxRkqEynq1LCtX9uhBNJ18GOAh6UdgHnr4C
19wOXM6IAQjzhxkj7WJ0486N+xLQ248WZ7e+idm9H/PZUGlrQg4shi7SQUAMAybW
s0ScvNsfLzGvBfFKd2K3eg0Xxcx2sIXy55x9UOI+6zDH1QlZex/dRUWCerb62LhI
XSm4r6okAIbiBLoIM7eS9hdLZU9txGPFzdPBqx6GnxbsRO5wU0UVPT4nzv3+jlrl
4rprX3CWVMjY6RsD1bDvJEzD7291G1ZD71FTT3rv3/AXGXH/2uz5si5+TYfld8v4
re4tnG6bCl0FeZvdz0gklAVdBmrTkuC0UtCadq4NaFzNg+lL+qJVKDYrYiwt0fY4
PizNOp4fj+kPaaoK+XNm2t32OQbq8BXoEukaZYvgkRy5XK1bPGnKgcYzTR/RUJIA
nlUhizMg9KnOpVCmZ4SGQSBm2oJiWEWxpwcWRsJsfUraz1E9YZDFlBR9m0ItEl7N
X99fcZtdiDZchEeqGjFiV2wqpqOlLTIZvcAYduuBe8CrJuitpzsGaclMCiSk5yHq
Y/kUIOSXNMr5d2HZIqxYttSTkFuVTKrdjWpdrMJJ/pcnNl4EK3IGAhrm2bxFci48
gYefcE1wikdxzPgG1xCzOg8uW2S8fQ8z8e1HAUXueyaSpNNa5Wtm9EH2P8dyVrJo
iy07XtDk6l8QbQ3cgHenCmZzWozCl5ul9G2HaBzilrfxdIHSUgfgbfrxudeiloKQ
bhjVSghJBCCyB2hTQFGcmt/NvuTPbBzsagNXb2oxJ0gVENbe/+7SDs1HKgcZ0/S1
32yWtZWsmGsBZBAIOAgXweuPQHbE9crGr0HXcaoHzj/KeN5TFjL7gG2WT8I8bCed
j9IPvvLAs20SK+Q8m1Wuus7/cW3nYC1+ajCieUakkSfhfzG/FOjcbzmn9KwWOsiA
bS1vI2kXY4vOhpaMTOE0F/mRH/ZKDBrjHKWfcMThZSRtXPx5jIyrsjhE2+nibnZY
rHJ4v4qenu7NP2TBDtyY74VXOzUv0WvMLOz1/ZgWSCQEuGakYic/4e8iMufBwJLL
q7kgVOE9MOhJDFIq3jbV0JzaTBOG8bKyFIVhhMnsdI/CwoZRXiGAnHzvOAqGCUJ8
+iRjD6IadeAimvsgQfFXEhk9PFHC/i9lQWSD1JRPzgqIeJniVqviDRTlNAcrGZZa
Rc1R1+TF8qq5B4aaxJqbhNAlgX7V76D9N/L8njVMYm6afl+9zKsUCw//nEYIZWqF
YSBIN4v9UPP1CcuUdDNO4mpjbfCsrlktFH+6/aXmuyu6ClT/Ao+5cIf6LAEVzIrE
X/rI+adhMC7us8Qij0rRMR6jBoe7dmKOsbsLkFmMgHTrmE7s458f/1zkTrT9oOtI
SJ6E7sRL9DeSchRWxsp7zvYqBp8VQkt8Zmx6pnGA6AycKIzsD8QIphflG/BugepQ
YBeturWlqz6UUO5zDbG5XWYrLhbaX/3EM0Dh7NsG1OUD7VXk7Vz2lfv/iegPcDNx
ZNPOR4tZUtnZKGW/VGtvhK6ZHKjQG9ZpxBbYS9PmHRY5IYOrUYIU0RU+uckumfbH
/mEcsJ/LalC+LNFqyHwvzG1ejkDcF2s/mRPxlOxMUGKlAepXRklKO5sXVSJJ9xye
1Rffwhn7XaNmIHIgxkjmogrfY/FU+Qu3B0I25dHm8bxOz2P5dBILJ2PrkwAM51m3
2abhnQgXEIl0FzoI4bNKXGBAlhHuy0pR1qWu8LixJj7fO54QLqYD2dK9Yk0HKArT
JkzqpB22X3GBq2Ni3O0Y7G58zwwtM8sCNjBX3/q5R37q201wv5vrZERnTIyBkSoz
w9mXo7ewpdB1E3Ht2Iri9VjtGQdGS+WGcVNY3gMc6K5BCxGiDfoyRySBp2CCmgTb
7+gGUDYipPObRu4mBuo+sC83nX62Lu8JPwbqxq7qLRIMTMtV0xdGubq6sZNGFOkN
jiH0rGq0Rxl++7e27x/iMJDklfZ4fqTUbFEe81og/bbNJRNON2i5LMwwjnfZ7QZW
WfLb1fUKlbUXyHbA7NDyeGBOnoFzSG7TWcUayWWGHwXnSMggFJs4mgi8U+mPY2KR
swx3IL76pu1F641DfBTvHOC+NRFOLgikEj1qp48cPMI8CXL0kdkewE1KO9NmJ8HM
Yx9tR5WpvNl6oFUPcbbhvVgIamqYq25p0nxgelfgbdIY7Bq44ze84a0OEN8Busq4
9yp0kxS7dVSFFgiJQqc8nZ1s0zxExBtejEeUAISfUjo5I9XsyAoV5z2BDnQ7vEm3
y7zV49XzhmXWZKzmk9ASRay3fFGiFl5US6S4WVMaFiL+o1LMp+QDVioW6w2HspXY
x9ZFD7dKukFg9oVn6oi5l545BqDkreya2awmNrh8CfP6LtKXJsvo0r33/5cd37lE
LWIL1ckZVzylq5uAK2+zDCZ/cM2zDxfZzQLJ2hXtYckWei/HH1CKwWwXRzqZiPdT
zUO5d343OhrHAJnuv87leOfSq3+VqZtYGWVVmLxHKF8DEvL+oriqRYTdNoAJuoKm
OXKC8jiR0LCNziLSxXD9WFyTsSkXfoBDqnmzOLhIA4uIk8sBPo/UtkSVbbF/J1SM
MDAvLmcjs975Uh6CsEXSZucjYMa/gr5WX4qPwd4xW8t2RMh3EuZxwMAeHqSB7oWi
mtyWrJuRMgnlO85bsbbLtc38Y0eBw6dh+OKdvq/W5hlxSCvVONj+1KvpAn0ZzBZr
ARPqm5dB3cDOkj6R578QabFOrK7VGqJNd1c6e9aj22FG0PV1bIS0xopuPwbBpNGE
xXFmLZ6+4fcWx9zpbOl07dsemAIeMw91gB71gmQpkMQ3FxpciUYnsHC4KqYQjSwn
Apny1x4+uJ/rmOgZ9eI66paBkrp0Ea8rZFrwGb+XOmFpyd087RciCHtVjq47kXUu
nfQiaJD1FZU6IwF4f/YrE3IGFdHZigUbwr6MmUXNLqZId8CpteZb6Ek8CsI2lO5I
PelyS94tzGgUTPRhf1WpmaSQMQyCSyaIU4qfqrtkEjAvlIvHZ24x2HVgedZk+6T0
a7kpy45segchVz8h4wsvVUdkJxFrY5kbYzllcjYGQ5E2zh+CKn0No+3ueGQnLkA1
zAOd73bpBp8uj/03lZOLD4b/tDnPtyu0b88aioAiJG6xKhjrUMOb/wqyh8m69i/Y
ck3tjNUWAKy6TKQY6GkJp+jJnNs9DYVQaTGTUJcZTTSDChWmWvri+mu6S6w1Eo7f
aoq0tVPCbzOELW5o8nMgt+y8M95TctObaqMtjDMov8q4rBas/jFs9N/v/J8t04Os
z93TaS1uT6SSy1auCxj80X8r5wNq2w9Gz2YDJhJvbensRBJUrC0FnjBgb6CIjqR2
CBa5Czy9wO+KrcDW+JHjYp80uLd5hDsp1i7AEemP/tx7c4nmNZJGHk0qIMzF24j9
LRWn8DrafOXturiS6Yrk/Tr8KVrsfq/6cH81c4m3Sr5BK3UFblsKMKsLD6pJbnzP
u5tzGNBy2lU4e/MBGz2fYZUmfh1HEqkhl/quY0AgL18dQyL/e44WqMPKT1kERZ6w
Sqy65GqfQ/euPWLCbCQ9b8W5pEM+wpCKPOR1xb11eXT0jqhCJQ0Z1t/rVD4MCFI9
oTZQ1nHjOUkLAlTYE/zyPcS2PAJjOYloufRujsa8aZlojE1sSuaLTY3yWd43tCYe
wAJvnhEWl+T3x830TgVufFcKEzG7Du+I2P+jAgQxCsJ9XGwa6hHLlC9cSWZMXALh
vts5VLdefEheZnWFn0X/PtD1TfVT6SGP3mlSrA1Brheow/iZUhh08rM3K8bp0sIF
v2cuqzHm2P8SUlNIZlf5PUSRTct6vEh5abbF7xi4uttT6NjhTT8CrQFd0V+kIFVi
3VFZ82LldgGbmY3PkLhQ+3GyVIjxp2XV0P6U072kC9RhpUHTZrILpfsw7wPy/nyj
rrBXvW+osz1l6zDnXjXE4aquSLK6tRGlkG9pcCipP7SLD5h5yrDTg9ByMTPzSWzQ
tEnWT4nDQNBb4RMaR4exQTqQa1Fssx/6YE0HTm+BIRUB951U8PUkiXFksPeoTUGT
jgGzYqotDST9xtIc7VZfUIdiKjwYkrYZF26052Mx1D1k8E4/sX3k3eGaai9K5up6
gKR/J1SD7VN2ELNvzqEhohuhuaWwn93WA8aAB1RtoRgpqP0BtBGprNF3znzn6IaP
/JNIBL1O7eqXhqSfd8maY4bBEC43e938vpi0kqylE0++lUDbT24I7ZNE5RfOgCFL
WGUjdigsxfbzDUyj521tP3stapf8sYZMelCBDAxmNgISUwHPtgpOn1VcBoI0Ed01
MYhqCZBt6BUPyPVbT6PlTG36zeF7MteuIoTePm+HIIRFpaZSYouB8Ze8BtSXNtEx
zpJP1UpPF91LN9XVJZf2/lS9VvIfE4LEmjaPomLE3jULYlFSJDicUjUNGrQlpRYS
46OeKDaiAxXxMMtpOoT2XLUBkIYc8dLegOaPR3QgRfsuWERELUI1imMCK15kutU+
i7k/kEllQ1KupHBuR7FOI0YFwWfkylkQ96ijkXR+ae07VRHSr4YbhfFzqufWiJd9
PvEoqoMAc9VtR7yHdF1vNHGfuocfJY+3GMwY+dxjyAfK7HMkMDt0p2fFq3aXWvd8
JlH8dYsm4WARrWJ6j8gkmsNHHEzdfx/2QO9aNoBSZkUsT7i/nisO+5CXSl9vJT2p
3PSxS6zpP1SFXXHFEUOio9h/rVn+i2lKFMhH4B9nTWFazbHPZnCdIZObvGKHf+jH
N4e4nqwURohyVNX/z95iCSMHQNOKxSFwXEtpzM6i6gMiIu2xd8dQXocx46vyhqb6
rJj4pHSQe1UpkiTJUByA/dLznMezvGGQzN1Gt+5e9mdXzHFglAy8v/P3A03LC1XS
SgWGWlTEY/qPNovvESMq6DdLcTjUDKyK2V+u+B5WdO14oB08Z8oFfSkNi95GMh7f
KM3cUSKI3T3VoMUVHRH4Tz21Oab1sB0DDFTSnF4FUdFDkZNszxyCyFnD0f0/UEgZ
XZHXGpPclJGwfU6E5UVVLLH01oY+PyPrX/ahqOMaPmPxZk3qrEkgXbOW01vq9c96
N2lfBGe/anYTKMXD562Q5FNBIwPQGRkGcc1nPbkEAVYzXHgdZZ8rLAPM1IbqBlf9
1IBqL74ZYLpjjwdjjienz3+apwqTBajBhy0CGAMxwi1hA59cCyHqpYE3C/nvE4Es
cniw5eNldBvMZEFSFjFzD8SysIRJIxiYkijclLPJnixTsyp+rZMIOPNQ5n3fINMC
qg9/yvpIENewVacJuo+a0TlMPKNcev5IKsiyWgsVpe6jgPnLDStsTW37LAHrxG48
UTQpH13Fe9zWE16JpMRm62g9Iz/nd/atzrqz0qsnAGrF/X3ugw2lZYGBZE3hVzB/
kmF9/p98zmsuUlRPX5wbYALMnkfvgYrfOLoLNBK1WVB4hIBETsPeuz1J5k0++vxV
pGIhfEgTB1tZqvTRoiMnJRA14Dm0pL+XvrzYXNxkWtfo+Tu8Me1nA4hQgyfo8f4F
d0lftRxMHADyrrR0hkrIiJrw7j4u47E7TtkFOfRw7HTBJilOd57zBx1HKuZKmio0
1ABFkLjjjXgzp4fo+q6oyNFHY4M9uc+TR5oD4/cM82KIef3ROf51ueymceBK9CDF
lTJbKck7B6YGFNmT8/vZHWS/Dtfq01GmM4sfbGF6Kp8Mv1rdgM9liEhgfaRdILux
FhnMDtNmj3HJNVApdnq5RlomWoSIH5AYgd6mkxPvqFN+szvB0Gnh8goLypkUGT2T
a16/iYrIR3cdcgpboz1wkiQCo0KhK04LEFRPjc3rzpADyO1+bP97H456bjqONs0z
NLzZDW6xXkd5e6M9YO//FSjropv7zNUnH69Yqo+ZoCj+8I43UBengt1Xd8l2L9Wa
QUc9fezCdr9mV3NIRrsxFzUZnJyZ6J65S9zAVCTCe8VPNi3UVjZ/g+fttSCBCYmf
93IjqiJj9//YJFFj8p7zpD3mpBsmfjNBi/UTGqEVfdMkJvJ0aKC2nJMSJdxo1RY3
i/987gDJ5+Bh1OVyOW67xrHfW+vLxkXSPtAbfef5UJoFYq36GTK62jOXy9p9d21m
P7+S+wQufST7LvIl5f6cP11RK7MLdvWFvaig3m9ff0pL1NMbqGOMGSX3uj9F7Tsm
0/gmeSsJy2nTd9pXRjvqCPZNjEJz5Dj28u8VFR4YrutFRR16fddf61vuMkx/J92D
2OK0qg7wtuW5tToz+tjSbWDmZqWnZqrn17hdeIbMT6elVxvygidZPZzITassrAyJ
KxAt2PU6+UWI05zVEfKdLDVskmefA0BDPmd4NRaSlY6Tyb9ZkKPuuviYiJV4lRCA
tfjR6Zfy5Nu5yuWx2RgzdZ0ImFWoykKD3P7YLqZIAk4DNArSj19yEXiyK+xkh14g
g09ov/aHcuOh1hBV6rjwHbU7iVw14ci6Dfo3PtHGak6k0mqy4QxYUe5VSFRtFPv4
gso3Vc5W0VEgYhr5GbJbPVopJ6iN0VhIXJEyi1DEQxboHIeUjEaUCtTcdk45NsuH
2kfRc8QxRxHXQxVLGIuzpHepBCux78wDpD+aXtLzKXL9N/JgIl+bIsxPYummS90i
fxWGmH+pr0+mnBLJr2NC9N85Fb0RIrYAPHoOnoUmtnXJ6rvvLhHdN7uyoqbCLY/k
K0Vz3CjU4JkMpscK5Wncc8ulLky8POhcMIiL7EtbXnlMaHWNAPZLfB4uebmz/61g
SsEonNVTzAS5bGRF39NXqcHpnkBEjBtmxHVYljezYI1gIaq4SuLo6dindpWp2oJ4
m3Yx2mu2hPBgMjPCIXPcxjxt/asNGW/bJ4x2046HysNWOPb2HfAxI+tVzXYRJuM1
BHChqv/DlEVhJRbRwJK6sIQ+rPx/WE5jzchqQePQWshdDpNRo0mIiq9BM6st5BfQ
SHMKPa2qsS374QWnle0XEkYNRAgJCwHBrB/dRv7kdZjS+Im6gxgMtDpoDc5U8MRj
6ZyUW+14Dm8LAbAidvnafgq5IAQMJi3nbZqsk80lQzjnWJjXyYjtogGfqgneBXLm
iks/yeZX5NSl2GVkFErfcUXs460nc0gTzRft6eufiv0uY+1z1QaUpx6+65h7EfCS
V4Gb+cJ1F64MlVQDegyasmK2JRoJNZEqz/4UgVh4xYI4V9zzNrShfWYc7pm0KAd3
zcTHvcAC0WJD1HTK/oKvBgJjof0i4rQe6w1RUUfkl2Zv+YJmAyiYdvcTui08lk5n
H34dzNyje8yg5I/BV88N3Lu+cc1GR2xB+/sL2NoU3FjXsUBGtgpvjseafry8gnz6
UdXB65cgqAQKP1+AUkd+LsG/gWfOvR2V1epubvbJN4mirfBRUmqigxF66ab1j0sa
LuPRCGyQsmpM05pLQnPZuy73K5kb6lA+t0dr5j/iibdPBnp7WN7WYi5UgQYuuvsW
O45xHaJJw8lYLM4ZlkjLkrUsy77+vxZ4Lt9/68bEJGy3Xr9ndnMZrHlTPYYGzlti
yq5HP+tklSqU/ejy31mCul4XnwpOVpXg108IC7G8nnZMIZHpB7iYyR5CHH6/79Wv
B4oRjziq/25hbrs1y34JGyDx7ep8uYLBYi87Qx1ZDoRQ9Cp44S7MtOu89zRK6WuW
r+aVwfHfBI3TVlz7BEFQbKlf9gR4EfmpWGlzrJ9kYteyVxIr8qgSHVWaWnDg41MM
wQaXVszV7yc5eEN8xl7PpwGYnuTRcg2gm6xY5byjOkce+daUHHJzgCiYQo5Yr1js
FDdO1H9lMgu0U9NrX+gnRcX5RLrSY067vlQ22YDzOS2nt1cAlhQvKM3HBnPd7boC
VfT1Lwcj1dBpw448JM+kjsLvMYqhXBEq2KQsUrJ0VJiKxdAFUO7Ys4KgCV+zhSSi
vN1MDwqEZJF7wRqcCLaI6OK5/sbgJBBL13pBbQDi9FkqlVcJuftZSLOM5i+Bn7RU
Qns5PZCL7xXC3SeggsJKRjF4Sf4a9XXcGNIyrP7RiZ3yjeA1G+O8naS5oQDa8Qt7
6ZtjpPid0HSjQ+HQYS8zk2khmNDVyYYZO2i63W3290uAi9IimOJhk9rZLa2HqJuj
Cxb2Ux4FXy0VM4G2v44JsAibdefbXqt5oPgO46CR/GXz5GWbj+3OyzvX4speTlfx
QuMPbnNwlvOWfMik/jASYEQBRRfy27Ni09jlxPK2FsBKX+3ZHl3q8+sAAe7GRIyz
YH0wUdKwcP3v/ZieR8QMYqgT6ytrSV67F9zme33Iy6o3toHdxY64b7cElKSfbMbW
jbKTU29MYykTRdhp2Inl/W5JRSmfR9zu+OyiW/6foi3p51+CBvWRLj7jD4xzy6cs
feqsHBzUgBoXvPaUHo1qKbTLbD3/JC2kcgSu5yfTv3tqy3rpsBeL2RXVXr7p3XYi
CN0kfgAV9HgGTk/Hhb00womt4ElFg9vxhXEpzVSLyL7nfk1vr1mmyWpYVZkRStHB
Pg/bCmUpq36c3gdi3r+dOJLWKQfsvXKynAIcBYTfVq2quSu+qTEtwygbieUtYuAD
WgXcupNIVV4hT7TXjBb6PFhlg3nZ77ksIBJzYUmNEvzxG1PgV5dAzeyWpm6RYTMe
q/gZAnbCDGf0tBcPaLWxOgoU6i7m2RL80YHcmiIwXvocZsT+uAbdzYST0gIpsrTp
JFFiHt62HZmg970Voj8iA9sn3b185CRQ5U7ktNVN5nI75pWwEM9scNRwUYwlamBu
V3G0ExYegiFBlPQoPwfMZ0agBaYw40DKDtNerNiepdTin4BjqeSeqrcMk5SP6rf1
vh3rNRli4FUgi0zWyj7sKfC58gEu40+rCY8i0YPHUXv2vfia9cHzOzkA9IvomieO
GooWybWVQUV1Wrs/jGCYMMvf7tbwpI4f63Dezs7IqzISEqY7Mo1hWrtWBUBCHcSU
8y8qVkUYmuF+Vu6L0mdsOEFCypJoh/AsVRTT/o9YY23B4Feadm+eJPjSnMf6C6pt
6V6m0ZckKncDykEEXsgLQKaX9sEZv4lCOcqSnrCTkDAI+Q9G9lDUmITiq7Y2oXqb
XmRwSeAZMNT0hKBUvRVjwtKneUdVSZHXyMr5ZMykurbFQciWfA2R2FTt6/wDqG1W
kiaM5HtD9YNJjqoFdPR9xlwYcHbzqFPj/xQn8WpxCRtIKC+Ft7MbDU15Dek90YV3
6ykHBmeJ8DX2P9geeO900WODkkMzrFmd2/3z9zMmSew2LWUxlBIfqLd2ba/gUr49
euYer+rFlm75lZDjOt2DCQ7xUK0bw9CxK3S3sBJewBB8ajoqs+jp12x+wxP6IF79
W44Qbq1bFVNygCZc6yezaatoRhw8FXZriASdPjV/eeU82JoSssjVawDTA4jMQ0x6
vi2+EeD7wLuGR9WALY9QfJQUVrQ2RZrCwkDbzhvD3BHTn/PMI4xEUo27kZ/8gUVq
5HkzFBPi3P/iZ4jlTyf6Jzw8PqDlJjbGhTrcw9GDRFV8NmyuRyytycBTykZ14WhQ
GRZ8XxJa7GSROhdsSfbzfX/kboTDiKxawgfFWdldUrM2Nt1QLFDRJK+uTQ97BtLm
DSMRrojOUZebzAsAwCYWpu7DLBJmLeXTW5KOnKezxL1FvHT5j/QrS6DbZvVSJjyB
unuRFL+8pGL6IAAA8SZlZANnMiGEhMi6WowAgxPam0qY4UBttNVsyI4i1Xh/rQ1e
5VTVRLEbub8WEneJvY3AJuqK8uoUUsQaXpJLxdWSa76tyNp23ALYB5zn0hBKfnS9
EBwf5QSAX4dgazCBQDJll44+E+xwBPAIYDnh67wlDYNQkrZyv5Czp+uwXoJBvPgF
OtFWHXi2S10CXV/y1oir0uBOyRQV+byom4Pt5UZzM6R5P2yLbfWuwDKBmej5sQN9
i7enXaX4AVgrDLPmLhtlGSsU8+qrQK9DZFhxLpsXGmQUcrgWfVh6/mHLWVMEjivu
Uc9gKm4hThEDXy/Cer5sv38vgMO5zathcZyf3DVi8wsNMmSl+/y94t5MSFrhwe7v
v5OLiteZaRoLws7/kQOWVswwr1rXgrYm6+v+mTsvAyYNQJQN7wisyPUVfDj8w8Ye
bMYlcb8c3Uk8FJZSrhb1d7gLlC1v3KtxCB9RmhzOTxI9zIEkOJT47MsZRtEKzujl
5LdLhUZuvLkaynKWndRQjdJAdSbUfTUOPnj3rHnwVlTmqvlDsmc6GIsHCrk0C1kP
Bn1n/j2CPd6Db+zfjbMhfwaw/yShP3LNdpjvTt93tqLj7SflPD9SBpCyVr26SZ3R
bNYuN9LpDSbtiyp+20IHxD0QNoBGnwOPm8LvjxLGdaHKrPabc9RQhP5LRvSq+SeF
wS5Z/1vDKxwfBYr1xI8kN2Rc9p9ltOQuWxsIynG5dhCuzWbP3dEHGOhkp5yq1vrR
5KsLOVc+ArPVsdHdDWCN40bDE9yXYULyHgWOCLO7+np2LMaRwtOjlky2/X0APSaz
tAwQIJIOR23pkkhXfHr8eQk0QQCmtZ/o6bSsmnUkPxo0yDeo293Z0smE9WodYkl1
2Br0YVzhqXXjdDPx+zJ6IQm6blmXWu3gQqg+37dgBWwct684sclHF+fOtcRgLp1Z
g4DP0gYV599rR/S9sRaXL8EeCaI4G2+w+SeKQP7/vXtsDIpLR2JXZJh1iyiyxktk
8uDbrWTwLOvKDqIGX+fyZ5fX2UHQBPPTcqyOXB6bjiFxvu027K9+073eTep3lVRd
qql7Ao6FPtWYxpkZkXqWsg/boL7u89oekyGrTnltHqDtFXmmeahKXWFNOV7e8IwO
TeiZgssgOLOMm9WKz0USk0Z8yL8+BcUCmBCjAgH8WXbVvJPYhyNwim23U12jLvPf
dvsrUaeS9Xi+NeG0wb3bDwjsUDMxhIUIuXzd2XRtMGPSRqCeBpjBZ8HtqAxpNBuU
7boVa6MWTiBnR0/4yJVA6pD1VC2gHCA+zjbgMqw0gk2zG/yMDuDSR//ql0uqHdki
W+FH2LTAKGYLcOwrbGbkp5uAkMLMCUoxDi20X1mGBZpBUDzcGyE5Dw+ig2ViDevY
zQGLXw8OjbjPVKVWFQ2VLi2jlrz5xCI34KsnNUEm1Lv8SJ2KkazNor8d2xAEk6HC
o+eRtDNOwm5JjwXgYMK3RHBrT5HZOeKhZCVJupcyzfguCE+81BegwgmgRWD8cGuk
aYXJ0/+/MltpBvNgnsz+tolNMim0ITrbiJF9G4RbRXmj3VpSepLrN4X8Vlc9tuqm
ZC/OY8FwldcgNx/+qRYP8MWR2vinHeXyIf1q4XDb2qtVhhzizVnULwVoTKfZh5Hu
mNZa2e+cvY9UbJOkp9kpLhWqugRGTJ7Ir0BwXIAOZPEgFkvlnbzST1/5unneobRd
O/3jh2QBx831th6LJQZRukzrz/etEuH7iEZKRQx7+ji1qe0o6V1R8RrFcC2PjxvB
8HMjprWEUYCXhDsIpEyr1obT/WkZZYKhc/DUTEGdcRiYtz7Ra1ZEl5O/0GQE/HDJ
q83nW9WlgHNrLw48LGhZfKj7mxRrrWEDmyWgahf5Nx9nsgcZ84EoOKx5eQk1ilrS
xJLiXD6+ffqACi3VE1QjgyAAFnGpntGsL1ECeew6IOwl/67AdCHOaqlqnCtfxKym
zzGzdTlZ77uQJr2sjAcptSLutWb8ho640/Uphe02dA3qxXQb9DHuOVMr9wJyoecS
LyRckXdQDbTves9GHjiGSFQ8xFOcTUE7GXyA4MveuGLAi9U0BDfzWU37Hd3iwQEX
DBx5nysgSoG3vFJJFZxl9RymIpgyNa5UyB+FttwwZabUswuTaI1KlIkWb3fp3BQL
P2LxtJrLGngW7EDtM24HNZFB0l9ZbQO9yIxPD7XMen1Bt+yOz3LdRkTqvDMBFCll
5ZtKtoXkKnQuv47KVWfavFt3nb8a5foIpXP/pCn652F3nx73Tf5E7pFHF7Ryvut1
4T87OvtpNodDHV7KnT2NdRjZmB0WfLdnRvZBBVyRytRYJ18Kn+X4e4wVFduS4kl3
D0+5DhX4LxLbsvFBgFAX18o/fr44xTUdppMcbPC0gERsX9vMnxHbBOunhZZgptJ0
/vX021GZjeblv9P5XmhJyknmVPxhwiyc/1MGKY7BCr6QTkwcN/yALfmlzVUknTfj
AdsIPc07E+lLgqtvEGRbKHR2CffA6bECD8mgOrYrIfmggd1FYXmeFT1fQZz/kTV2
OnKhAkuWvHGcC6VL0Sa34dm5zvNTxe9xqFTh4y9552Nwmt8DnX2mzryke163LmsN
q1bOuIL+jKKJCyH98wnLZ6z9yLUbhhIdp7eAV5P9edvxY6ktDRbh31FB625Idlx4
aVd/wS2/8URGBchKaksXMLwtjQ9+3S82j//muQB5c3TmsOMMbMS+E2q98/ylwThV
zLDPMU/jo+5hmDPcVkEntbh9aUL6ctqtYNxiKnUCnfvdMRcuCTr+UeLr5cwmqgQs
qDgTeHV7f58LZjXuw7uBSw69wb3mPluJQotQqSAfzDv7RnHQkvREt72Vb/xDmwoy
oPJ1HKopdvcPNdaJHkq1borlLOSguySlzJlTsLNQsogmh41bKyuD32bgjxs51JPQ
aQJu2mZL8i8/GQXA5Z1laik4aSNpw4lXPkROXEHKUk6UUjajkb1oD/xNRHBQB9RP
7KTB6i7MYlht4Dfi9pn4ZXcPsKitazxvq9MpIdFiZSzZR+8a/L46fDjGi/N3tCG1
0JLnPx8+qcylLwGtRy5NNOyhYiAWycJyJ05wD3QQKc15W0EaKhu/4uDbJI6CJ3um
dcwRnM0qTtI0qt39N30T69WnsqShPJWnBLT2OV9uEc6jSByZcvhexihHjy9TdCBM
0lkWfbY9WNR89BIRFpPkl+Y46mUTqtoM8SsLHwHMnZ+Ik8v8svzjipSGkeENpMlZ
peDGqwLIC7URJenk5ttzQeNCcY64pn8Zxe71fdV1hC5zS0XKcXDqZjBSugHnKow/
z14NhZZD4vb5xMXs6+wpKPk2KrbPCEFSpvEmrqwBdVW5/Br4FcLz0QsFri1KJiXi
5YGCYfmbnP5+X2ajWAfm+U+YeKwPtNhW2LD6uUIdpwHp4n05mBm19ujA3HX6bBBl
Gb8RuD8bhPd27iDzDFZ2Zwi23tUE9ML9El+27xBWePMcnAkdjcjA3/C3B7Lhsajk
fJzaXKbM7SIYPktqxsFTjTc40EuegAqTIlxsDJabLtXgUIMHiTbSjbNBZVf3z628
OcqBeJ69BlXGdq27/mLHYKkeReFH0Cmw+6/eFc562ksyfG/c0bdbn6YGHi+Br5op
g+Rfi8DwM+6rFby6XOuP5iW2ga70KjOc2tGAjvtw7T/wixBz11m6kOuMabl0VDW9
odiytFH9IDBPZBBzWtaRnKKqZrIqOud/kt1gabp+PJRwlV7qN5D0qDVsCwRzvCDE
c9HtvWkIEWSLYxvE8JpQMpBPUVnHThDNeSdV9AtIvrR0HwqKpOjhVWxcQc7sj3cX
xW8ktitP+q4FRYCaADi+hCGCwBWj+qYEdEh9yaXyG15xXNXV8yCeNQo9ugz661rF
AIaOFrU4+vK7n/ndbgcvSgc4Yjj5UxzXrq55ATpIa6ikBky+qbNTlxV7yOUjZswr
XCMyLJCOs8p9toaLti0ps+0wrBMxjLsOtoGLAapQqYZzKbsPsnD5pyFManRJjKRZ
YZjPW2hV2jhn1aO8FTdy0XRoYUDFI8LViofvg0M/pt5nptZUXpmXptPQspewSqsT
1F5ZfpTvPHg2bSRaKG/KXxX9nmxvq+CO/TtFEK/eNrfYXfhs4xDPs6SlAJU8q0JM
LWN4w9o/su3Vyy6RzhRRpua5jD37Ch34l6b+nHOnht526x7EurcUAPcNnre3DmmM
IBPFz1e9c9mOTmnlfDJihkxeTvEEdgvwufBoY3YPhg+iS6eb+C9xYnY/RAn/V83T
Id9Yrw6aRn9ewP5KMMqSD/6qmIhCcJ2bXl+2Zj/7jGXWWn0Bi04wshfUyaFfmxNW
UfVyI/BTgjJnafHbJqkJPXfEPRqmGdhNHLDG193PbGry4Y16FH4Jn/eGalOruYWe
GdpnbESLMxdFyexxB5Yh3KIgae4bHsbBSLP/cY1YEvswA1zvF/4+jHVOPAq2RCq6
e4B2NpCq7TB0QUqDAgVGE9CV8taQLd/0jDnWIcJFXBTt0Ttz9YLGVzzXO1QAXd93
E8PBpqMd1HcVwgUowApDX1LNM3nM61KAo9lmoJ5fATBewVws/2ceX6xft5VFmbIa
7T1JFj0//nAJj0Wek5RXPhSisHET6P/7j7d1PzumnWi0ZIul21q0G9XwIEwQHyDO
S087N19IOC6ELqlvCyJqbAb1NcR/J7IWdk+09M67SAOBYTMkEnzy/MURKJ0HsR98
Ix46rA26DJ90Dqeu2ThVbA+KcGVJrRw/29gThk5AJuIEr9kzjZ+gU5dVoM1lVPRd
3mnGhLmAucjQ+I2DQF39LJAK5Tu2xFGr0roK/uuKyXTp8BGHXISqsqhv9BVAck/D
TDZyH+I3jBu93fT1MvS1AjM9WHwiJPkI4dkAuo0wtO85qaqmKCVjD0Dal2uwi833
X+WqOydiBOQCM+LrdL3P4IQU1JIUFVTGQqJJUo2ikCbXzU513+FGqVw8gplcTdgS
f4ID7IpRorb10sA5Tw6ODNfRI0c/fEQuAEWhwatAibQZgLKJb7HymDaSxCShYasL
eTXuLkItSuhmO8eBrUaR4nOQ/wiYhGzaiEP3/kaHuZtO+Z1yEucWTHFpQcArHGTk
dbh0rxHe2MCApquSXlXWDzC6Ei2VqfakF4nRwZORLfdnDD9rAKbyfrhetgZRiRIt
ghBV59+aTxl/vp7eadyjPQcYGWalE9UzLh9LeA9/RtXe64Ty1K6s18R7Q22Ikn7o
VE+ewQhrpmvy6Cme1DcXBQM/RGUUhM9GKrIW9V+DJd56bwTSJimLKrGf+lfsNol2
SuHD74cEoycw3kSga2aYLdB8c2CTOQ0Yf/M7CWtd0VMFyiYAwy+EXbxZyVd39FK3
dDVHFgx3UZ9XPfTUfRgkfFUgLFQE+H5Ru4ndL2Lz8rEiQWSkbZgC2ZDpK+RqYihI
nZWnpMus3ECIAb3iNJ2fF1UAfRnrhir/p6sQ3VVPs3v48Fm5Jr33SN8VLZ+O6+pj
qQUCTjgFzwRKDErduUvPLgpOZKVmkYmJqS0glnMRFyvMRZLV+tjPnltp8W/ePnl+
vpLYCDp27QkgDZL6G2X0wbAjOzrl7XMECzPlw3KX1sT4dAo/QPLCokxXbu6C0fDM
QQaYr2U79YHq9Y0hbZyQPk0Q7gcWzivGu9FjZVLUQTAdvIUkdmXUr7rhBYx8UaRR
AY6avVMtRvbkUGPrLo+7dOd5bjXNc1w5n0Z0REYz2fLQGRnNaUEZoGglZzZvW0VM
Sli9/tgiCnoRrMSw7xuK9JaE9W2bcVIPk8CKMAlhKcQlY/ElI2r1V5vC40s24DV9
awnlsB25w1z2z9IXowvhya5DClmyWH1PtMFJLSgmVq4EiYOY1MU5A7zwKBjcCh39
qUVP+tJNIEAAwbpCTltwe6ILnxw/7AshJF5J5/3qYkagMA1wANoyKp7dKEqbDC7k
WgfwXu8G2XvvRHUa7O+OasMp4QS0Csu/kQXcTqIlnxNrMylKG1is9IsMbstSHKAQ
8/Vn7stuLU86Nb21xGo1brUlrBI9M5RknBDc/CHJzBAxpx9b1RMnICYaSBSWMRYA
/rv7tdsGZqgDNDsFluys/2euTSe39swIOETpyOyml9+xUoiOnBhQ9FScxHikC+BL
ne8hwrj7YhJFbGQJ3xgrUswoDuJIhpOrKXJsztQ3X3xGIhvplbCHRnXjErnPkwZG
+BEnfBk541IR4glQaMo9iMg21sF6/j/f5PUcTwgIKZWwkOKVAyxr8iSwt+1hbkKU
qVZZU38QHi4PFEcyZ1Os5d1bFmUu2+uusFJ1KHGpNreyAPZUp3XnUaS7PqX1ymze
TBSeHasiH0QLpPt9qaVgJa8xC3KxTDzA3kTk6/o5EDTJtnaieVybE0qOMsg5HRZA
67aJOU38k8wfESv5kz8aaLzkMRyjp3hs8em6iNRyuy0NHJu4ZX4np39OO38R29mm
sv39zO4U+YHKUu0+DZOEEOIFh6POx4ZOnqvm5sTbR4f1fRMIMr7H2mwEcj3TTBmm
LOyMykdQqJt30NcInxNxQLiI6m/tJIv0E5Fk6KkKZMWH+CvpYkPWCD2OXExZKqm2
F3q9qeXhM75tp4gm9RD+9RSh+amUTk2TlC+Nfzz/SO3pkBYoX2rLX9VYK4ZgwFtd
NvK4puRzgjfkyUkHyfjbl0qv7/EMp5uEfQhW5LKKMp7sSfnSdxExH8QABmd7LWdb
jJ9pthnxMn2loFxfyQojcXG2j4rXiaBwmtrsmtGBPVKIa8oOXpkj1kimBtQfCzVZ
+mBOyiY2piDiPI5PjcMNDUOkO3T9YXkqxHLjxLDK9C+V/oUmrJ+kW+L+01knUQ3P
4VmUi1ZZ83vfxHyZ30DwXg+jTFhzaBwxg/ZhZjVE7a+vjLVwR0Nr5e+fK2dmmuKb
rzVc2F/niTFPlElAgk3t044aed8XV4uxUktFdz0slRZ9KYyV3j16MW5unlrAk2Bs
Y5aI1Tqbg31+XJ5jQguT0tUaKZ1v1nkrxTVP278H0BkLGexVDAQKivG/zYIdL4M+
Ut23eZpT9GqCijTeIoGVBk/g9TGl/hJQOA+pntUFigIUozzwLOMTelCOieONCGm5
9nX37Hxy9idlWEEpLA7BC6tbbxEeH7GqwD0xlPYZpvTULg7HB7u29p4eq0GsNXod
2cKz9HIQrV3uGFEGFo5sbqP8FiIoJPZfLR44yPNUTAEzk6TzKUSibrwlMtrdQpl4
G0IgELGgVrkVNJcwAkkvYxyCmyiRQvA/YQcW5VFcJxuYOM0fFvgXjIWbszZJGQ8W
v0bq2w2BWGB/sjfkm8Z1uz+0dQLIariIDFva3mBRhZYgxwlwd4p/Nej9Jg3M0X4H
iXICyYLy3zu8mylEhLtVO1C1xmDFZcNAeONyVDOFClK681L6RuWou9admzxugymN
CetoM3l2IIuv79kLGrxC8qneQTpHO6fBcr88JYPEUJTI2FE44szQ9MtpgqZQFvMV
eFtAzF5kQ6y1Ucy1JpBBqdhtf0p9tyYv2XTJi00WJk6SdIgFoO3odV6CX/m026hL
WUUNOVFD/omOQ1NlRf1Og23QUyXmzu10K+kE5ZUqE09pnx7xhkDmg97MpSb426N6
SS4+B8iLF5FHqkkJsT5E6v71MTeIho2PJNb6/T2PDjI5WpIpx5iEOt+NzqOeCwUV
qHa2CiLt2/OFH+ZdHmvbGB/LBX2tS42828IwW7Ux1T5j1VrHR5rNwacla5Y/F9x9
abGzmmqinbXAXGA+aMWPGe9u+KvM7xaTGlY0/s6WWn+a4qT4+Hrwib4j9wi9R8EV
TyfGdLFgZd91Gkji8xnsHPxMMttOIiy1LaBU4d/jf94zBTvhC14KL+ke6CYsLaQy
8dsvGIAn7dHFUAo4I1JI1/bFkfC0nT6K1LK6Jp77yknxijN8Kq4cS2sIVA8Bu8iv
jwXHzkf1l8k1DVw7mdQjRMfb/n6wXteaeSod61Xr6dHID3iUwd/0eTcl/28rbB/U
0ws6UG4aWEtnBFveWKXutP6w+MKaD+geJfdHxRaE0xA09r5Np7bgsDAMv3wxXWmR
UcJ5wni9MWdaVVOSxw57QZb4WQu1ZvoVUar89GEVln6DNu0rj86c7IrLg64iY8C7
lCZczJrkk27mSatgOHy8d+oSAo29uK0m3r4TwPXapuzNZc/IHf8cvKVabsiy8iPF
8gaHLcLT7oFdWMSaBX1iDteH1rfBp5GpWu1lzTph7UAgbOhr5WlP97MyIY74K393
eGRnCYM8zqzK3kBYvXHdsSoOecvKUGxzpFw+8UfiLSg5GHNBjPQqUxnUaUuRPq3N
16THHMRYfGSEhIX0g5ZicWfXokEhQHUCDrVpbtDgO+I3BwroR1LyCl1iAwqBV++y
x2ZNoRENHyioS1S4eGkaU0Ez5R3CMZAt9igKqnwwvgl5Of5bhxQDYXMIydqW95NB
0F8rkxoY9nlIGBNhSbT2nj05xHxQ8E1GZsJyBh4oO8tbfJDTzzmC69w+VcB1fN4w
GkkHYQqsrrfGS1met5NbRJCvsmROzgP9clUOzsBmlXL3/EWwmx2L5X0Mdl2wLphZ
zzKosy4rxnDwe2/AYlrialtjb0Pj0NPHrvoxveoFg5ROuEpIM/gVE4V0WhfIiRrX
EIMV0MxkwVu3Jd4E8zkMz/0w3oyNylCPk4cMinEA3BNrNbY729bZg5ugAFo0UlMn
IEHRr1sE1wfj8/DdSM4lJ7EdqoRLkJJipp3BeCQ+bu/+jKDnIwcn9mPtjtpdDO/l
Idu8FHM8sNyHsupF3yuR8OBH+YH60b3MSpHNJ1Hyxg3XcmeUnmNhgimdSdn/fy62
gjdhWT4IUmKLibIyDWxUZ6Pl6QoF+I8mV07wIU2pgyUw1xerCkqFo+w4kJkD31MK
Vf26QwI5siLqlRSluwn9mfzZmRQZEWCFx17TL2DZ4nnX/PiLpYCVjRC/AAde9ruA
MAX89P2cWazxgNauEbMtwgnuLnLrx6JIDus4Nv/j5E4Ko7oOT1RRaNABZBynQOnp
BlryBTZMWAPcEywMoCRtoXuM+ncJ6CDH4NQh9XbSIysW3kTSyBjrXED/8aAbwXSr
U41tZPKDMtq61RpuULaZqaopO2K1AwpulIZUMzkV7pWrjnOU1yZ37KhHBhhaZWf6
vpjFL0voDs3byF75YnyuHnGvdpB2IZHvelmlwKtdpkL2w1oCUYonUGcaM94WjHnO
PzFdr2A0gT6oxNaxEYzmhwSXlYfxPYc5cnQaJzuqfCCGA20EjP7iRZmK8/PbMr1L
N+xDzUow4KIeLCYrFEs/xadrPYKzg+DIYo5l51fpN5iJq2fYgAABcawP80yCeLQh
x/6R0YXSpGx7ItUU2pEMiuB1jjbLRc7VCx1BJ483+2A0YHJU29UN0VjaB9lGkoP5
N6s02Me0QrgXODVQFMwWPIBnL2pERenHwQaQy0+pO1+iWqNt2giEAPxVk9rBFM2/
W50Ja6JTpv8sani3FTSOqO7YO1P4x4fGtBHiCSDm32V0avA6gw+no+eTDTVRF5tW
tMzv0c0d7z3SiEU/ZPKEfi+8OAy2dYHBZ80lEdYykxlDrrj2em1aKE6bnD30RMRM
bXhYaNuTAx3aEfoPW7GScbDZWzyYJge6YKSBw7YyHMQ/51jOnb0tWflezRbr2njH
5q2whN90MBii0IMlHKrmeaBEVj/kSk+0Det/s2u43m3pug2eVyxLpJZdtj/Vdcay
eblQK/ge6gml9e85PfcTfcuZalngnqFYHRkVpBuxog2P8nqFktWf9HLe/4xt0dze
fWig4KZ2ZBCnffhLnkrFEV+d6JwiTb+FryWXuKz4HJyJkLlho1ifrVNpODRF9R34
8KcY79JFIzr8hbMbl6trEzVnrEro+7y+4+/W1z7RcU9PLFzyJT45Pu3J+83dpqLD
k1mOahHc7JfruqJQJkiRESUudH5W/wr5FaACpyCiFbltPchd1ZepiagDyxW9c4RO
2KPqgdj2f127zKIkH8NL03QSYAW5NhmND0BpYBKJmLeQwdk57Z1nobD7lLuIUMBr
Q/AQoOITEGjAkM2LB1DS7TaEzJ+snKnmT5ZtQveN7QXio7Q0ZcRzdnnddmxoO74x
HUMDCKbTgxy5Qxo2OIy0oZPVxbenEg7yb+YPbfwKfRnT8FDB4xeXA3i5LOi8BQfh
HMWp/bonnRhVnci0vWRqsZEPeSn2N5wkompEEW1M76fuiPA3WPTkiiHrEZ92Ui1i
tCBsrIts6m6hK85umwztiGmXigV92Kxvfv/RMzzCHVJkowvBXKtua1n/tPIzA12k
b0MjN1dW5uO5WWSFpsSZC+/4IpyUVEQI5p/tIfFrnG9H2UKWWxS+L0NLbldNB36e
VH4DxnI60sj93EI8nnNVeVTmb2uDC/7ZenrYezJIMTFw3IV9LlJk1qMWjDD8Yz2r
88RpBq/PoY/b7LJhcAMpmOi4axn819Voam/HkYff7t7hI4vheEf7ekMDuW3BHImI
FAQ6vqCnZZs3GEaiqVxMFqeld5mNh6Q7bKgOTKk6T2pzk2ZsbRTT4rRELwfOHzrY
ioFSpUOO0pUIB5NFoDB6VlXrEGXAfb+bPC4TtQo0oktI6WJdDkcFLeZJcOXMfZ8k
tGnAswaW/C58dgw8FRO/4yRiyCMyYKeA/AvxxWBRBAQiJgAaSfq1kTCY3NTk7o7m
CDV0S7cP9hEO387oViRHOuemWuKUOm3cCr5k/MJsGcAlvCJXvmBUMXO9Z8L/bBV3
HMvB/NrWrht0PD+EX5RPwDKqqxWlXerB3gaByIdbfa1RFGJyXfrQnsRVNmFT1USv
vPVSSOapjnJixxje1RxaYLB7oKey2V8YHZCeaggRfAevD3SERGOxkOS7TMnMlJXt
Rp0e/Ki0ZfaFW/GB7rn2IsLMMtnfBah78eDBDPX9lFoaVWZdwzpazER1GK/Vftb2
5992xXM9wdJu0ElOJ/calQAKvW6DsY2dBG4SUybD2ejtBSrdCKAMrUh+3QqGIVr7
iuiIUMwtQHcDl1y09fhpXh6k248hwraFaHXhqoRF2gEYy+p2GnIX6xGN7St3gs0b
DQJClnMqX6sBS5LxHPl/e3KskNjLbUU7jzGv/d+h8/n88jICWksW2KJ+DEG+/cAU
suQ0vwEJUH9kqf8vA/Kr6QNA8os+IPK5hN2gUrWbrgG3z2q5vfww6XQMWciAFcOv
bIPjp49kpaM12UALNSv2zRyaB2UtXg+oOfYmZXu+FD+/mflU/wcE+md/a7lKTxMq
zJiQJZMUS8m8wkrB4bWkBbVqm1p+7vdkAuWiQTxaR3k+LW5N9xPhAeyZU2bzsNCF
5P+Yd1Bvi+X/oD5gE9IWZHIPB2w9JbUGe6VWoKUNqcfdSBSjJEiSwU0N6WckEo7m
kadpIg/ETMuGN1V76yt2CQM7sbsBtyz2bvnlv3bRu9910ATt9EnLEMwUBLHP6Qmq
Z+eD/p6ruBV1qKY/UunnGibJ9Rgo1cJDRMpTkMU5yfwHYORqm+MrPmTjsWmtBHS6
42xDzI3aNid2cuYazkF2TMnQelZkJpXu2oKmINRzhneEob8HXTdI6WKkZQyypJv7
WAw91cjJD7G0E4SIKgRdcT1zguGXj4EtY2JyRjLOWhSJZ7Kf//08mGpgtf6cnowA
223nliUj8RLJDPpuGSFQJ5GL1D1zYpH5wCxZOWDZbK3GJX+CgKlOjf7TH3Y/Z7Sp
Thsa3gdE/ygoqSOSJF9lKIvZ2fiBZZUbmS8kNO4s44htOXD2BT/kTCKSYcua6DZk
ni1GV+iDRnRhptzJiOLj1m1qYlbUdaK253pxzF3obn9h/2JuSX8aycx7aCU/ccs1
VBj2b4Qgrhd42/rDQUV6rPGXwgdpvixTtOHWMnuFXxtonFRyVTna4bEwQ/STsyNz
k2aO9zXRHcgoiDyDtkGmvIBXwJMyJeeO3OO0yCBFeosMiQFZorrXJ7MD2Ght1tZl
WeuTri8PSLGG2P8bAxbPJHkwAuXAHMVdriGDBPqf+GJSllQ3WN85VsOiR5jQos8e
a0JjlNlU4xlBUTGBMWjQsxE5fKhorj3r0AagbCc+NlTYOh9AQQ5LdpSWGl/+sU7O
rqJk8jcXEPxhy2T3aW9CzUxKKSj28RrKTLZYVx1UCGGnjOa46LEEW4rpaEiS5mn0
rM2TOpPT3G3vfrtzwCZjBrbYqep/9IdTiaVEirVH7qZ+LmyLstfjcZC6mRSOWD7N
37psM1elBIFEhRX2qLT4zJYcx2Qx6Qfjj0GVc7W3v+1esIEAqEk5ehFkMhM7CrcH
zZsjJb4iLbxcWcnHqb8b9/QUOR9ko4E2gRqrIxZNGx6iY2L2pprd3nnyNs1S5rA1
aYPLvTISF3S9QFFK0/QsInZLORwhwRCbZNMMzLHXP2KwwD1pRbk9LclpHc9jHNWt
omPDLtY4yhBGsY6L/82cFzuSu+cLJ3d0Nb2rDYqkcA4eWLAMxJwUGgm8Ug5Y+vI0
tE9Z7VMCxTqPHbkBngIVySEdFZBMzJPCis08L4gvuXVygkJcBB4x60gMJEmf5aez
EWQU4me6Cmew6NLb/bI+99bCi84VUrCCtX/nuMPptCVA0e6Btkc2vGYNpTXnRVk3
0p2mH25OTXJMdB/eZkKBKqjXyUuB4QhGtsvwwK1V5/0TKTZBJJMG7R0T9mPupxkY
ibeEsGpP01dkLT+NKYMH5bA8bkRaoMz/CKmQeOg0y+/ePNy3fM5EL6idRUK6Po7C
OmvGPr+l6aa4w7WPlqvd3dRE2pXuenicrclya1d7LfvT+8RW3Bd9VW35jdCX95et
f2txpRBbCXzP+K0IGwO39XN6XBLsAgJX2yWmQUC3WemwBP0joYvcqDfKLOBz/Nkr
1bS727RvJECwINizBMkUS+1SSzxbs5YdlEr/eZ31Jj9P1H65BWQTzD8XUXz1CD3e
tc+hKtZmiCiIc0QmKaHhE65JExv+HpW6ShOOcx8O+E0eU3tP6o1u8OTyJ6YXG5NP
US/mNnZqssoQuj+UPwACQIaoj336Sa7PttDbxmnF14LcUKV1CIDB/T5kl1rvs/CS
XyEK77TBD6wLwGdZ8r/dppTiSEZVuGqjweo9Dec5xaMN4asULXSNo2355WABRgQV
Vb06OhXJKRvvtiOQx2Tspu5gS1B014wfCLgC1zOfFJHi/dG9BAULrJTX4ww1OLUv
hBiUu9GpHi14TJDyMT68aacAcM+Zty82vgnVX+Ru2e7TCAuEUQl6GJljVGMm3XAf
qSvvdsxc8DcfYL85WWyn7e032GmvHnakIcj8+upbpmN41B/W6uNhbRPar9WgIvWa
2L7tHee5qo0y4wkz9olyJRFI/q0TEEXSL8BcB2y1nMUzrO5eoVkpkFEOp/9qMts/
iBTvFmVOJbmcG0/9otD+edkPP+MFnrfgvzfXcxG+cHsUcCBlaW0wZWKmoAMo/K/U
XE6uwbDlRKqACmGhzDLqsXHiK92T/H+YhxkpbKnO6SHKrj6t9F7MZ6i+qbOE+lyj
fiqmlea+MtVs6lmkqMhEWuKKPHvR4ece8TnvPZv+ovaWR5rRyz0rIHSUPA5ofZ86
+jMurMD2VjgHltksi2dBMLmtUUdsvCNeTfP0tulJut8P1jpM3nyK9/a9P4j6k9Ko
+Qmjf74mM1Gl59hu+I8Id3aExLrst2Pyn7Nu2UuLDnd7rxEgASgB3287dvBtdvpT
86Skqi0L5yUgl63fB+n0h8IRAS22zu9sHWTfSZMPj6T6eM2yvBiIAlEyhGqf+noq
naQWK/Z+1D7oVIXCgi+IK7EjmJOE/6KqHUXZerz8NzsMVgSziEFhXBI92Ed6/0wJ
CEu7IuNMBkOwoujILWLdnFGYGdZ+UGQnwrp2CRRaStg7fEL4Aa31696ssNs4zeK4
DgFJuKVqjZp24WGsBRrlqGoKQCKXuUB3M2qWHZWiyQuFDFAZh4eJ1ToxRt4B1FNW
sqjHUdea9N+Gu6nQ9V7DS3bIT3v4/KcPybSsOVcyjIc+B3OgmnmwZZ1knfPZ2xSZ
lUuBRB/J/KY9MTaWvlfnfHEYDl/8SYktDBWBf/zSdfdq8ErehY6s1Xgz3+6rgNHc
kViLwQmWYLaeTAjwtyEBv1DV/zGdFG6KpgnlEN+tjoRue5WBjZhbAcS5ZWdNIwDl
SDzyV6faTKcJ97OzaXn0SeK+f844w1AkroXZECPPk+54PAM2aPA6u1WT/udlVk1x
pYXxN0iTcuSg4Mex+Ip9C6TbvBWqituBFEgf1MefadPIthS0Ex0QS4UFu6HcoOJC
3n77JvLaq2tP3bo9Dd6eP9Zy56fSr+jsyt1sBDqPB/bi/gLsRyP+iWadXcuZUX0+
LRW9+wSAsMFqgxZ3hUE7iBEpQGv1D9QIL+GEgzI/mMr+UuUDFqf5x3wkz46ORJ5D
3BDK6Wgeoh0MmD75FPV078d2q73ShZcyPSb8rhoDKjC5hyKb0hkhMBXT/msnYLNi
lY4AVZjWEzaO4RlS4Bxie5Q9qhbBarRopmD5Te2hOUH1gCYVrzm1xksv838+OKZx
q5noKe5j3HiBrwDnRymbpzoJm5/s1Y8ZfG0+9rg+Tz4EZmSG548SpR6gpdeNibDk
LKqfRe2Omk5Cj4+HsBhhnoZeBUe+aesx2CEZf4TNgJgT3rpJ6ORi4oSoKMwe9+4W
bmGRg4qR6mrVxszWGF2wdMkaaxeG0Z5ZQFklwohHIDqzz0MXtnisuAWwHdEfz0nv
eLA6qkhpUhry1/f7aSVMYQb35ClDrRCyrMWDQ5DU1AdQQQJ3uaPQQQwy2LXHVg07
MzYkfkC7uhYHC4snuwquRTxqkRX1re247QG462jWS8Bvocd+7K8gYoffg4+tg3et
MMuaUBZ8IY+eHY0y0atSO0BoqVVRYb3Fj/UFVaTg3esITy8lAG55DreuWHotkJBA
X1kRe5gwQ5+mGks7UuDq6LlXVShx2MqZz5ov177oNICmbTGCGyie1fKwdpsbAGqE
IMVV5byjCt6E3hu3GaYfgl0Ud8ZS3TmBElPuDR4jgmWrez2MNP1cC8uosjKJPndH
TU3QW//5w1IWBBkM0EjOyChHeLrnvWalGtsXRMIN8bJsxKPA1tmiL/Cx4l/F60s7
vIpUPU+Naz0YJFl9FiID7kLWafWbbV5Ot1BZrWd8x16QHGfpjN1jSXIcSBQUEnfv
HVcuCQEIJCk5JiSWXDt5V2Gp/vbNgP3s8vAKqTqVqn8AFLZz++VPFonnVLnI6Lc/
+Xb1BJA64zHLo6qk/xT+toxZxWxvRwIxtm4K2+6Cv/PVBt/7TcXgczIi/pbQLLPP
WcMWhtjsk/Rv/lGj0xzyromr/Mymln447Ul+mWqScR6kBkAbvBqYBGVJK/OJA7C0
DHvHIiD+bXWaxhw6ervk8b+IBXnNk+nGWchM7Jr6nj2toIEAAGKw+BdnNEQHRL9I
4mHibKreAZqg8mAdZmDNvBopxvd/vo6N7Xxx357+wkM+4TsucfBUF5KAX5hzeDLv
pzDUcCLs1IFzIqWwZ/qcFGSx5hcoMsl5WS9Iv3LExoCsIlSewHOe+eg86lGMtT4X
M+eR58M6sJiR0viP1O0JpXGV8DWZ9WfDZTtKgnW3ZE2iLnPqRjPSi4RMMVLXpefN
W6Z9Angu2XMfgPmcE5Nzq/Zgvf+HAIY6xwFpw2Z9S40Cj908zNcnUlmxWI4TO8rQ
YZli9xClHe/mJxHDqEpwXjAPF8IizXJY0WCeWUJJesv6gNlACWpMHlmWjMBp5l0d
IKOQe9jtyg2dT9hPiH3ZXOjpCC64vGfsGOhJjORV1I5qApEU4rO1WKAAgV6wcmSI
EcXwDU8XBkrGSqk2A2RP/js4TnzzQCGEwmAJ3g57c+fCeakc5Qpd7uWbunqRuV3k
/I2hkMskiYi7kSW9d34YIayXCbqmmRle4zaqFtMn1/Hb6MbpZ3FeuEi5X8X4Sdxe
OYps6++FFV8A9IwyRNgPGTKdzL9i9io0fgfHHd19471v9AGZqIhemeu/6QRt1B6l
I7+WoUVGzYl2zvBhcpbur4BBjUeLtJlXyhTIpb81yvPrg/1v59T14y7bZK4DZeLq
nnbCI/4BSu09l1E51HuOw9IbFP+u9kec1rjRVnk0BiEqv3I0yTiX7AacL7yY/FEb
S+OAutt9N0gRq0SFtlxiO7Zyyr1xyZWq0a8Fg/lUXZypn5dBjBmVH+yRpnz9sJZk
suSqzq7Tvaxsy/ncI9yQU6YbzT4joOEVjy8Z+Hb7ANezbxkkuXki1+sFYdPebShh
tes3yA+560QPHALRcJ6J5Rdy42dmKL2dVK2qedowQANcEkLAce1Fo5YGKCpmMySy
WvlLdsNJj9Rwh4iiF/azA1gngpPr5fnMOq7Ua2olX/bJc+5ZArMeRkaBh2LrtptE
1Pn/tl1UtjD4UL+3D3QKvXe5wWILoou/NckheYyjodaDxrbn0moOiQjwnLvGp/9P
Y7Sxq2ZShORY3okAkuztWTxQ6PT6vCEtS5OtybaKy+5TiZqWoS0kRqV54m//31c+
z1zQ4I9roK8LjYm/F0QQlwPp2RDI223CN9brT3/ZpZEUp8InB02Ef6kFU8wJdIiy
OUXtFaKJSfxGc6LLD0z4erl5bwrQZ3E/V3uKMUAhl4HA6PC2DxbEGARF6yxiYjl8
lq1oVucovkK2gmQ5r3QuevStWZkUq3XZu7iI0q4K5zCkBb0klAA2P+TD0KEOef6J
GBjDawPRyfIs9IJYgimXRroyP1ZiA3XiQZ3qy4ldMELpygc3Kh6fIOKuh//3dl0V
fzWIMaVCqCCv4ytIgWgrugDFkM7hVH/WmHcstZhdIWIArMkzh8nrgqG7DaYyHF/P
fbwhU35dhUyOwzTmz0EZU+1eGRdcN2ntLO483ufPkVH15p/1lYyhB5o3dI4fhELT
9IyL+864pc3ADIVBfASx1toN9TTxhRezJeZHfp5yfHrrVrwuKgm6Xxm7ZSX3clIi
aZYNeM+ug3OQYfeRAWhDqL1Y2xy5MuCXlRGQ/fwdQmDx2PyZ46UVlYhrNWHst4y9
VMQeClE/JXVcXjUaYYNv0uiaJQIDiC44nywrWuThICkH8HY8ygAyo0yLA8ZloeXq
mp61X8umbnf7vH0AQtj8IjW0mZFaN3v1bFIw7/hYorOewg2vxh+AXFfJEMpBTkpj
Kp99GZbx2FU9Ua1/ZYhn/MK+BvPQox1cHMBDrmqeretGZylbBgMm4v/4cEzrLhN6
vi94L7mXNsuytK8l8E1awHqifTZnAGXBCrXO5mb6ZknX5Rc7kcB5ZfFaG1ZczM+F
PBL6xJ/BTMz27Y+YyFfT92zIzrBn82iKGP4l9jaix2OmTH7lLZKjNbCcOuikb6fF
Jt6FPS0D0GSvUQcaIgsUaEfZLaX735F04RcRXUyGaTSdH6nOD/+KkC3SC8o5c9vL
OWrkYlCPXxwzT63N8eWL+7UJtyOxYHED3pIaSpxZR2pveYTY3jQfy38gZhYcZZ/V
sVxlurMtarq5CUlKYZ9zb8fMKHqDZQkvHeRYAI3JCcyxGBqyaKaM/CI/ujr7A3/+
EZmWi8TBcZWHwRQKcHdIGr6rl0OpDscP05UWPqixOai4osrMtI1JM94pTWl5xozT
l1j/go8tBNECeBb3XCOz5sdUhby3J1vJYTzu6xybrAHxVffE4yPACrCI7FEBsoTj
yc3x8HU7UPH9taNkjBs3EDLosZrxrqKyBWJ7ZuFx7ZX9JgUD9aA6eOjxv5LkHATp
Q1Lc7V3q+9m4WFAZRuP/2acq+5jzxA2PZPYHL1+AXUgqu6AuUm3cvszQf2+wiWOM
k208wnGhOtHifJKiQIDxyHh4N1Vis5E8mxj0fUhtaFUOCFctZOKg46S7A1txYTtO
FKWg3rUHUjVleuCcSMctwDq8Jov67O5NHn3KQox5QqT1UjuXEltJxcGyQUzmxcg/
/EJM23fgX08WAxzVm6KFwEgeakf+xz+mcQacCGOzy7gHX19dIPO4cnIoijLCXhMJ
D/O8s8IEkySav5cCgx2EGdMpe1lzABO+WPrqpcuO4mXnGuWjatFo1i+0lmYS1UMN
uXTTtIXgVNsyaVKDgt59zVezgBgBeO6Yfngf3LlGpxWCZ+eCyn+Y01CgwNcIptAF
uwVaWO17xsHRKvsf5VsrhKAoGQ1s0SlvKK4rPvCZ8zZea7jzvpGOOELBb3oEYIOw
eoYpkpWa/38o8G2QNO7ynSRMRgOsGZiB/P19LsCCgTfvfD1vx/ldBhni0YYe62Zp
3Ay2zq6HGsp+ttZB0sTCXCVnWmeQbcTDoYbeN4qZ5yQ9TBncw8c04/7OcTI5G3gM
5LjPwyXvmiL8dC1a2u2lTFj7vVTV44BMtQxPSUUZ/0Xv40h+8v9bHpyrq1ArY+2L
/SHyR/8RAMjnXw4Mh98UL7Q81bFTrkj4M8zDlwKdOJVGxJr736HmBy8PxNdtbhrr
v2BYR4Ec7Sltc+mtDWTK8WjlZ3xd3nqO/4r/7uOEohWW6/EVUYlhsDJtH3quZR4K
huLakn/Pu1LXnWTmKEaZKFiZ/GesDpa63g/YGjK/vHQbVfsV5FjhIO4lWis6bfSm
rFJe+qQkn/wUbXELDQqdYRLBq4l33bmSdi5GbB0VE54FCj3ceEru7rcul/WhEJx4
lT20YG+B5oomprEVhuoUTNliqdUtyIJEwUeR+c3KT2cUE4/IuB/kEJlcUz5l5g3O
uykTWRWwWe2R4UQB0Mn9L2l3TpiUtltH8+z0StaNYfFWVm53V9A0Ouui6cnm1vFB
BMj2WdVxmYsER+Y5xTBqOiBiApaAWwh8JPnmxTu3PHrNhnmSYv/VwJccTrhYypkw
ZebJ9U9CBhe0B3y2BuNWuzkdvbzwm1OS+uB19SWCbO+SHE/wPRQZh/2iBoIwExj/
A0d00LhpmGNFIJV+4A+V2Az/58ML3XhYtlhndmqlkt1XEJEgwa/8VXNNjWr3bwNN
NfVcmtQGZFSaskj8InhOrVE0HRTl2JW9zvRCSTUfyq6/kssSMjOHbK4Uard9hVOz
DtDcUuSYUT3oJAlaHED+FEOFFyOGOgdoAlx+KVGLM6DtFpxFh05//OFRldDBLu6b
ODKLvOZjRDKYbdERNrc918pqAR0+oDSbo25xt+q0GlYeLLlk+nH0aW+QTTHKgV9c
0QqRafn0f+lkI3fWio3GHcbm9hYFhz0oGHt+TojTVCh++ShB/ABTYEWUpH52ajam
13LBAFIwyA9puao+V2Sxo3YveKtGDjNS0/n70o+Xd+ybBpruAWs4FbRpzoW3kSh8
4x014EIRIGn2+yv/BaOB1yFp3YAxAAx2m2i6t+QKxUIt0zla3ijLW8fxeop9chyj
QQ6q3DlFzwKfEoRoX1X4AmbGJIbpe+sCmc7FRiBhLH7/4vlJT+26RqvUP5heaJC4
YFg3YB4sK3i7V68cdoZRG59L7dUXk8DRER6F+VK0MywGDXTSYobeSdqXbRJlDvPs
eUrRo3RGkRUJhyDRYUHHa4VZtTmEKc4rZL0EuQW3Tr+fBqBK+v+clpYcGroch+WN
NlLUueJbefnbbU94IRFVDv+0ygnJ+5depH1nh14urbHx0tXK646weT+BL1e36CP1
bZBLvk8lSe7VvQKn/Eh9BRBs+nMtYM/umZqeeNK8wRT/b+Yu05ejUssFygpZkKT7
oTjXq+Wo2NGd/vusuSshTCJeRj4C+WSltBlaPtfIzsCz2CMIr6iAVMUQI8Jj6IMv
0LfsRyooGwt6TMofm4Kpc0wtHjMRxFghwXC2KTMpQ7ARm1clcL6J5P/AlNIeepPn
qHTDRlW0GuTI/Slk2oq1L/LAY3h9huBQT8ZmI/JhmTR/Pf9R3ZnG3lOTrTRlac64
8yVaSNNKZvNrGMzgBpJOPzipuX/rDlkVWHVwz3V2I4qMclG+Yckqe1ovUdt3VB1q
DTNfIb1lHgIIy9z6OtW8htqOkrRw27oSb2MH0kfU47MhKHDukD9iUO57PVLluLVC
vGLZndIcPn4SVVyIPuW/OirfvyPPJOxjBZ19bjHTowgZiP3PzoOh6nxtp5CGUeEG
xoPnm/VBW5CPssl8gK23NTrmP1fByfu1jyIwe4tA/CpSVAjJ6tsBfFRKz7vQKg+t
ig+hLpCoOpruue66bJNLZohlpiWoEECzeTrWcRS/3oSg2ZfTyw4BbdnxECHtfvmr
DmKwMp2jkKX/5n149ub6nFgrqNl7Tebo8GoUcgUEFNKo8Y8WsEyCoExHEK+oHphk
CSbe1oY3eTSNzKdr4FwkLOtP8pyBYLSc9nEiAqCqu6JHMWBUHyVSTma+tA7Yokii
qJ4TvuzSe3Z1N7tS94P+kkHJEBpHGKmY3aQ7g2rzBtnV3ykPyeW+rzKEPfmRuDX6
Hdy0y7YnxWvJZXt56IwBzhqpTRui65TVu9jyK20kxJXQQ2eRvpz82KSNDUX1b7AO
JEZjH6XO2FuCS+trxz5tEzF1JIqilOvFDPGcri3WjarMnExB5XHzY/1ucX0vyLov
the29svMbzy6doslR2NqMjrZvEBPZKDruY+4Up4nTwpoTED/d06gorB8vYRDrr5H
DBFj3WrnuAR6u6RcY0qNy8jjf9sP6N/NRwaOKxKzKVAJIgUNY8oc3Sjyx3mvygEq
S6AtjytSmb1pDa3gkE2dywvAtlTLaw2f5kPFoze7Kk1y9XKeIcbdgDTA8+pBfGCs
P3e3Ey0xoyXf4t1EdxAfkrfGgdFs/t1kpKydh5LDukC77XYsP0lfFWyAthQ/YF6j
W/PFnZ967ffIk3yeePjSk1IqUdDN62ym/4V1eF719AIx6Bfsz88E8V0Di9ftkB+w
81dQQPOijHd324PzmQzU0LtZWhboz4C4V+6bEInbahYrpVXcxYOddYFQx0FlPvCr
YPRrX/taiP3YhvQkT/PT1L0/HB7U3STxBj0fnWTd5s1JQj5FopCt/9IlgIKaDjyC
rwY2CIGN/DkYj7iOG8CMhCWR1yI6gIDowicchN/53jXMX42XOAryfCOz/id6K5RN
RcD4PSYzy+jtMNBCXc0f0/V4QZql63YntH493563Jvnw1Rm3cENYPryoABQGKPOd
x3RIkgIoA6LeA6U2j0OFzhuXPqWMrRAoeUW4mhBw20VYWTVhLA+jnbHcVe3szNgi
dhEfhr5e9tpNT4cdVoY7oAU6hW298PoPBhCZK6+HP71sRXMlG1sGLZclBk7f7Zzt
Np5Bp7IufImwMRdox23CpRAHm/ISNfHwOFxXkt3E9cLXizNtFXagY8BsSyIPgIjK
kpzvhgYMg0/ncVzkoX5ZxAnFetMSwzVbfPITWwAu/qO8gpandnlYbeU/Voe961i2
+J+UzsFqScdKRLgmgM0CFrsIsg6bu/Bl6/CxU1x3eTE9uFB1iHVAIk3ls7U9TUEA
o92Ye+5RjtEIlkz0zEty9WK0otEhbHKM9MT3yE2u0Gz+Dsg6jvQzz9rHBOQnWoPe
bv8wR4Rm+5/T2/w3IdibljVfpzrdai7oj3KSJuyQ8vNH4X7M9XuJDhok6zrOgmnK
e24hWbONe4g6eYQHB0DWP+hP64bc8IzZVD2vfx/11iIzBM5f2BxpBMcVDXUC2rid
/SU/r0CcNkiBWTmcKpLC1SL7HF5wBFCXSXa8XihH/TIhjLT4EzHJ/tEHhm/eh9PQ
dNez2CM4Ly7Z2KMLzO9dITKIDgaMfG7OqBrsjzP/KZLYEpejmYeLeosu6gS2sqhV
WGlnrpmx+lJmNEFTxob0PjU0Acre60jiTkSjiI9rHAHo/g+KvQB+DxY8Xwx2uOlU
2p5wJNqve5b6ao5I15aTIvJhSPmycFMc3sM4aYDuHil2eCtna90bo3TlAgXqnTfQ
EC9o3UJtT5JJ+43jS7k9dpkjDSwbugDfyVAOB4iGuWRnBUQylujE5yUUnSxj4jvi
OANHnkPW/ILOYw0EUOKppPE1gv6YoxqRFLKvaBlQTuuEmMBybBMf5Ft+bXZsLwoI
xj6ZoXXWAiU4gjPEaF9eH8DuHnev7ThkFkrc8C33QeC5/+FfUp+PxsN9iLmvjmrp
K3bqlgaV97iYFBeCZ2nKU5m2kJDf5Zj0NEbQYITctgnJmBxsrqeQz19lGJsF2W7V
8eeJPn0bjx+nIqGJKEZ+kaaVrOHcNx7TbgZdvM7R9XrKj3DTu6AdoKm/ZPfC9Yhv
2XHx4Fud/B5uCMJ7dHImWnTDHowcq5VT+jz2lMn26K7B8PmKqdxXtVh6dqA2dRb2
bDaGS1SV7iIoC9oukqb5HJtX7AnBqIjvUOQ2TkWsHC+hgz8lxUDrvX0o7j0b3bZs
2ceC9ioroI59sEv5cN7eON4lXMpxojvKxUsXw17kHztzhmtKrg70PEGxUi6Uuf/B
F6/Y0x/loh1bH/6O9wld4luX3RwK6K5ND3BRJJf+jgN16npsXIfVoQDV9pl6Hbvy
dKzFJNQCkH9KFC6IqXvwWZmKPF4krne4FOujranWCANaxXmuTrjf9nexUHLbOc+X
6IFB+qVCwpcsuqhMYFSDoiCaluSH8b3cyxpRAoLHKZes6TycFYfD+nL2Ave3RrDk
yzqMv975AOPWif8+PvkeAfTM6ynKnbjtOYtls8WIXF+nNS5SbhH9ZmO9FWoQU9iT
rn1pSL3emDsCI1Uh6AFkwvMoug+LaChYLzuLCXfBjJKpJCcrUc9tcZVnkKRR/YK2
zn90gvh+tYj05H319nLZQK9I2c5yQYShHoemYBJ8W95hYXmFCsFB2MndJpgpksLS
1le7NrMOa4zZpkqkRIJL93f6k+l6srzwKFFzsNTRijaDEGRmFnkHu2cqe+ABw6RO
/uYTQqkIBKo83nLanzj5uYFBUdMQQjZgx3rqGYgckMHvwzBhdWN+q0R4o5L5hAHb
MWwjDjGpCfTzrX/aDaS6pcGYHeqF+QY+/qgTAMhi7YmHHJ9Wj4KyD3txztd/NsLU
NIai2vWMtwiyzF8ILiOlkU54BhicwiYtdhN6wk+99jQyyYbgmYaVgCsqhkRkFEc2
231mSUm4DdQ56YYxpGhQDf764FRczQZG7wl4JFjovUD9pyUI1rR2ThCx4BnCSVQ+
udkyDnw+cAVqZOb1Hk+sVCVY09SWM4htv5lubzrbyi0af+ldeEtXMOlZoVT2sVay
VEqKzYb0AJrD3jK5ZcZlt38o3l1SIN2hPZxW8FZs5JWZ4k4C119NSMgx7d0jb9cN
TyjmKfCkjcVLHyoF8jKWLvc/Rc0skeLHj0JIZNyANYae7iiix06MN9yd0xIPrN5g
SUJr0kj5mf9SDhm2nerc4dw/QmUjrEFx5r2VTdEK0N85EOHmoP8KO+wfuDPaqiPQ
TULJNDLK6AtZOxPi8uZmVVa68CBRe/ux4y/q5wIeQ/P506y8ZyUAwvcUxByGZ+l0
0gG2Ww0rk5ZGpJZn8g3QL9vpd81Km9HuYv8LiyHiEwOUlr81iF4m3RN72CZCTftb
csm3UEXmCettB3bOU07FOPMwxHOWjk4mAjWd3+3xIjoypUk4g98R3Va2SiYck3Ty
FSsf0BAHDFMe4e4LCYiqLtQbvXKJk71aEyb6xpcmwWuQ4128D0++SywKGgXxt42a
I5CaIMs8xmCgAvP0jhN3junM2o3amalp2coHY3v9H6Fbt4ckyM/9/Mzf6C/ijMG+
paLAVXVk0vKDT2+SEh1JcKQJNUYDrReD2cEOIqZIh6B8pnQMOAutIjipyigzZ9wZ
fTiDYgOIrMPvPnDcIEIWNh0kkSoqEtaMugt0Z+oEhkQI3J/djFy6tBYbr9urAw4p
hLe2KGL1Hbed9oFiTpNjMbiUQMSLIR9eUSv8sGJ+wTGm0XSEdqJ0AvUStpHeQzJC
CAwVixThHNBzm8SAkvTbmsdPfkdXtoQOCCVBM4vD1ejGFWvhb7Pr0MVEymcfAYAI
mNKzRJw3pbMRg9D4Y2/WWF7dPErn+YD9Ye/l5akKQk4nIt4KxB7xaTYTzbt69jpS
Yeqz49DdUPMAbA+V3GYwP2oGuuEARRK7V9FiQubZOXEzXo7oOwoJtOo4Cis2+8d2
anK1V05SQp5mcyz/gffKZAFaKOxV0elG9sPPw6hUqYLDcl6HMK3is5Xi0GWIYrnu
26O1VqY3RFjhPvFxPvn607pXv9ynbIswhFKzORa/zowR4Plt1OxPBaQLoP4oqPlH
RQU6wY6Q2iSL524GRe3LgrA44CFnKd3EzwSsexDuPiMHWXhSx61pJHDynljhJJ4f
ujhV3QNUHuNJXlnQl3w5s0gQPcqkUYcUAM/KP5Y58ysBaDUCDJC8mffHIJaH3Hws
Euft7MujMmlB8sJHTljKk1/z5ehKYkhB70UXi+HGuOnXBBYk5IpGrQV3XckguYsG
9LueMNcqWjEqRPCbJYMRSKz4cfs4C7BjDox9LnJJc2XHxvTYCbF4mXtSet82eGoO
l9p+drMLz4uuZVPBjGv8AL4Gz8Zn9vYYflLxPcLFj99x0Sit38gM831U1b+PKe7m
BeQaMVOYWglizUZ2K2PfnDKns4/BlNsrmGDEV6Gmm5xEgFMJAcwSLgfwrmwSu7UK
C77aZcjMh34am9B0LZC4UFvPtZX4fZQmZbOMjecaMEkk4OZjGs20IpdkCVVd1r4c
U6MbbsK1hPCeULQkW+fQSLIKdjBNkGvGMjd3X/gFlHo2EvEIBDCe0bwVGSFmXDCS
jJlyKvRkDyzhJJamTc4MaZee7HTyQsZBWuYY9zWVMv9RPV2rmrYZzV77Gqf3bwUl
nojIyXGNyDdNiyp/pdSY5fymH7hP5xzoZsd0v6J4s+NPTN672vVuRZIelshzv34u
n2Y8XlxJuXDSd+RlZKyAkyiUKWTeBNzCGhOlwp2Kzmg+p2G1XwgiXAXplbFZ/VzU
B69bWET5qJ1ebx2bBzWL9o3KxOUsoOswsZGa1EaJ8EJ7ACHrulmfLaVaURMWiYDh
bXFbEM77KnQmdzwWsYgxw8UBb4zGicQaSbEsxwNqUwC1nlx2vFxTVcZcE4VACcw6
mbJ7tsAT2ZoMP+wAFWpSQHk4fvvHc8nVulgU0ETZZrLhXR0C2VGEWB3cI/a/XRhX
bUYvRf5xMCZ364YU6gu8aHjBDpW+mKZ4IfG2xD/Tsjb/on3+u7iCQmR4dDHvrEzR
kE3DGwAUxb8gq4d61Yd15oVviKPo031vLYB9mMgT+aCydIP5ihRtaGI9yjYTR/xk
LRqd04iFbHvdf36sc68m2j6QkM2N/Mo9y/OKaCfpWli6DeOZ5cmAzKjwUXM+mNq9
VofqfI0PDUMvGWzwX5CLDk3IDwbDPp4CQC2QxhwvBPWhDqqOu8XNbIwYJKHRodPL
kZXmr3/R4vi5iEzI+/Msgmdp4G9FtQk5FmOvaf2cATsK8BdEyoPObNcLE+8LvkYw
sIZBiuucS8U/PbVR449iqZLgr477clX6TNyGzInw5D1ullOmbK3KkBuj8mlfYl09
qmHKqFchXmQ+XQSoq9tguaUsqVfgMBHPjIBs6xAWc5bYoZlirnuV+FwYnCEuVDS3
WuNpQqB668OcaBpotGZqm8O1K3sYVJzv7IQrr/gYXpPkz5kzmVAxiKOgZyQLfxDS
ekdS12UnoL2TOlCeleEZ8FNGkN49AnbMLfkRfWWzLAS2McLWsrdTiu3mdBJrFWJD
5vhvDbXMMFd2fAuzcmjOs+65nXMcGckhwrPlqsWv1RLogBJYvDIfXNj2UF+1ahE1
JeexDtUAeqG7+QAQ7EzF21xve2GwKoyI8bRqKdunEsUpxMJ0NH8azuWJGoFrTp3F
7CCEo9Jp2ZRHihXLVACs0T7SZ+F3RAQ9K0Pkn8uTzIgSlICUsSwzUWjfnCgNI5U4
KNug5Pg6AbJkuQo76oNhJZzXBT0VNAa68DHjdYjRgzDd3irwVeiTmwK40xGpevDR
H5IeWiCfYNT47iyh+sWxXt1U176OuNKuCWO29BumZpAuhs+Sy4aEouUYSBlmC09G
84fjq6EV5y/0I7XfJ1KGhHfqR4/6aCdsozSQNSpnk0er2itBqQ4efACm4D9sjlaC
98aQsYz81RlTDhdZlDZWi8SoGesnDhgy6ZtSl1hRoNEBpdiyTFuRcwWT/vyUTkP9
W0ZkOEckUWQRMjnRfMB9TGlFw6RvoWhlfakcLv7huX6OJNxYBN7kxX/tV2cknIdW
Sy7Akdj8Fu1CHfHU7HLKPVTHzBQzomc/yZOjtnZf8ehdoQSta0cjuDwGuSOYH3Wl
cPSlOnbsqQUvgxPhkffbTFBKuzKWYnjqyvZBBfZW8Zhgvp4g70f1K9opg1OFdCE9
1vFzpIIazUIw80hGHJ1tW+QdDl4sMMyOtgFX2m+9/51T5d6HHVIDudkZvOIgVhDp
Ith5LaDRrk0h4GrZvMwDiuTl/RSMtd3CexWlKi3fMNCjNe9BXgITmlfrZhb7LPOE
r8CBpb269nVya+hzo+ogTYnARHtvoQR8bDX1Wc9Z1R0nl6m2EdaX9H6QHS5umwF9
dN6n/qRNFmIRcySERanCG176VLt3z3h5uVNrsNHcVl3OBgYpanICSVG1CMQRu0tx
cLlAR25HwHKhBIcdLq7jUDggF+V9EihCsv3dmK2yFXPbXFLdqJSYVZSCeDQkIIcV
Kd0Lfbadw71kuf0h2b91mEAxP9djR5pRg54UKKtPrFTVKNIIaXEwuxfXwemqg0ED
Bby+/1EfFixeiu4X+rG8ytiZQDJa4veZN3Yao5Jl7EcPPAqmuUVyq9e1crbBCci6
UMRAwNwOZqJtKV5Zu3dSn1sJwbLqRThC9QvWujXnLZihP8ae6w0GIWq1VAuE8Chq
XqT/ZjThnNbcwDgYT6+0+8/JZLgB3+3vrTZya+Zw9LzotAt+zbR8GokAcfEUvneC
LHqZGIxLeSv3yjQMfkih6yK1xRz2zVZ+f04FYAQkMYU8NISZFYthQ0wGEYaVob8T
gS/1ZWqNV33SFBZbQqs+QlsznGNLwIuP0DN4CaLZuA745uK5V9lxnhj8R5VLaPcR
lGoEnzIkjzDEXawIIgTO9yOPjYMsX1e4kPQh0nP/jXVzYSjXkfhSTS4tiqmT32RX
gcVUymoPAwmtZC7gLc3Myxj2UInL6OhPph4obLsX3UPe9Aj43h5eKYrl0ALs+39J
Mf+pV3xvN5gzl6WiZH9XF7M0GZzJtbJ2gIRG7c+HxP4YcPpuunVMNGnzM5IwquY3
nmcSJm438lYzbf0LBrjPOmP+eZWusywbwb1iVAKdVrtcAYfoJsUHanDXSR1C7fZ9
Fxro8CzCPU3kHdquF3anzITAy7axzJhXJoteMXzd/D/fAmyQ7z/uaTEXcDk1A99y
iUKHMcMNAt6i8awGA0xTFPBorA+N+Hx6+keamRyXHYfsOvOzJ8o2RFj3S55zNpBk
IURaX7lky+BTM1LuQ3izqWEvIRmItJfWrntrU6bZjTqxtL8sIaASWgtPrTRzbIVq
QDQSqfJdkeSNzUIlQVxQ8gzarcV/MeLTFmP4Hpb6WPtEQN5s2aFStk9UTrRJx/hf
AqxL6bH/sWBIouJgnLMZOyj3tBaMDira8HhZKefCERwQpw157QF71kuOXO8NVuE8
a25Dwj0Dq1LoqqavWmHBrCMKb02v+AUFufC9K9znAWBkSO/CPvait2HAl4ACBTHR
Y8Jv9vNbE3U7gYhGMKB64IgbOE/Oe+zEPHZytT3CkCm2iotvx8nLOpZtMuSW/CUs
VBgBFmLjyty9l8bbJ0TG3LeyEWNVZRhwqBZd8I0idoByn0HXV0NdzFySfWrECu0a
qelK3XwHwfgZIIkEPpYVS7I0K6RSRONPGObzpT5YNVxvNgyHHhLffL6Vlqk/DvzM
MVDM5Q6eYo/9y0PbR357vKCBmvQercfO0jndhNUdCBNwNBNxg+cORbuVnGoDWaqy
HXPd2u1hKm9xflQx3+3iyan14cTxwCmfhhVtBmP+aOzdJEEdj6hkF7+BIuxIUEht
zMNZTmRMBrTpq1B9IGAKqRXJbcw6WufTF3KVBqNEEeItsqmDJTHdo5aRO3y/x75C
YFERp760ZQVZ47zwba4ig2tC/qV/4gRTuQBkKu4tHYMmv9BKzGWBplBB6bq/wjxi
yDS7VuaGc84fpzVGOcJEiiSWjrkla2JI4sCee2BN08kylPeNSVaAPT07w8tV4B9E
pqZ9QLbs3eMlZZyyuHp6wsLDuEnmsS4EWwTaY2lqxoaWOhBvR2iaBStY6YBrfuV1
L7LogDRLUGh8K7Gp24ordlttNsnfbXVbQwPeCsQqPiS6Sk6eemZR3/h9qC9p+f8U
6n8e+MdMEeL44HsqvjWSQUxVv5QZLU/FtT7aEbzeudQxaw6q3f8aKpTsdmoFeW12
Z+IdO94nw135Vpt2v8Aoe3thXvVCNmumrVbvaWOBuJrsbiheeK6wAjGJ62FwSdgq
TctvIlYf9J6a+I45FoXSkg2+4MNmX/2O5zexkYYpydHf0l3R+IufEDPp+M2EAVR6
qBIYWbTF9Xhdy866SMSrZt2HTkbYl6XQRsu/Qv5TDleXUfjh8016p/daKuFBKnOy
AcXiw3ziVRpFZfKV3PG3maDdc306ZQDo2eL2EHu/EI/5z2X38vgZelPg1W0aHLPZ
f91NDDrUiSdnKx4JZduMQYkcNvqGUxFVKqjPyzGZI7npk3zjvzVInAeX3suih8j5
7EKatlZD18qGboyLgp0SJeF5qJmdJf3Xu1uEtpy66cnTSNkUnEIIJNnmKpF6IiTY
yn4WxjgBywR8mlX4dt44gprTR4wI+DBHyjRnMcWWuWsxrFGPvJCJU1gMyyFlS31d
EJR5Cqr4eHUR/zkKIHNVCDiv5WPl/0SccXhhrTYi4lFt8F1LiatjokZRF66y+LKd
03UvZmy4b8ED3nMRZ3oNr+57dCLSsLU6a9wp941+33ka4h6eHlQftWel+Q1rlSCc
ujo/LIt45nKcqRdI4YHcmhi33ssegimoHkwoSBlaw1EtL8l62ZhyHP7EmA/CWElP
J7B9AmkdnMp5ST3pn9SBDT892HdJMxSgo0fDQzpYKP5q9SfqaDJ1Bd0GXQOMy4kU
PvW4TE8lU9Yuqv77SWYeHKftTv7cExyuJ35oPAzyw60CmgCw//FSD/FNf5MUg5hu
imD19BIf2iGUVeHcpIcyyZKtrNAhFGzKVKf4b2giTU+SFmWiAX2f0TcYX95UKQXY
YjL4TFQRf4LAllf2n279sI0tqlV9HYdNGoi04PzSmRNF+KLA9xjS3rGpVWpyfcE/
1i4Zkz8htznj3D/6pCtdFLzx+PYx8s3FDOYaH2BqM//YTrdDZIDkzWwtUgf4hVOv
R0Upj4jF1C+B/53HvdfHHekSHtd7FHHWB/uUVAAG1IbnpXoy9Yj4egcq+tP7GkiT
UEMNAAX/1P4HF/ll66hdTdTVgPYtI3m3iS+1Epgo1tSaq8Vq5DncHYgM6zvA5HwR
AGx+bRNKRr4wI3eTyrt8H5JYdslQWm5wWVJUJl7DRf89cthntL2j+xgphXU1pXne
ZiG1i8IW3JbF7AfXukVP13/mJVUex+/cVf+/EDS78kh2/1avjp9NAhn8pYdEoPG4
de0lf8wN/gpakE3bRbS2P276oTYUddFNVcTRrO5ZzTAHXiIh+0sr80xTJPXhkRaX
GK7hwSmIAsnjTGRQKDtV4HlHhWcL/jc0iJJCSkexR6YsX6VBeDNtbdxtCeG33o5y
+cKOWsVz7ds+AcqniVhU1yxLD2Q7oIYc7dSNiGFhyP3pZkXtyTBV12TtnQEfxwKx
lt5azhOuSxVkmpligUg2GO6Zz+QEr24ksiBTYFe5vcMiHh2mNJsQXW5r/eJc+Cgi
hDerQ0jd+YlBe7P37I0++LeEMkqox0txqJYi2bjqNjnEq/XZUm/339oFg2679Vgj
7as6Wsw8yW7rtfhirWlZg+L7ea/sh++hXs3Ty7QaMUsm7ZdIrdgyMet8+SbF9dS0
hJH2o0+yeG/eQrmn210MWmtz5U3LWfgyBCIUuXiut3d3U+RbScsE47rCBXfGy9vm
RW4e9VFbSkE0oubP9/QWJfEjJZ2XG9o/pJvTrGJYtpaqr5VAzAOT5x9Selwgeq2H
n53uET2anKYVFMrpSq6fNb/sWohSYsrjWWbl2c+p3pJl6khfAcouNvzS25Ja3eaf
1gMyHj84WUxMR65O9byZTE9xC8tuK9DZsIf+4FWmjyRrOL0CwcP4BsMGK1Jx0KN1
Fma3MJLl3ppS6AgbcdWj0ajciaE54r2dUP4HOMIk/dj2VcW2LvL6NNQfpczopImX
N51iz3NQ6+Qj22FB+SLdfC682U2awy2vH+J2s95F3EuYof85r6VaQvZ55j/a6VD3
jiO1GlzaytO8vLxtt+0fvp8LbJe61FfkQPcFQ+1MinXuhCLXD8TbHd5zkneDDsEC
F1FrD2QDzG7+hVxwI78W4atlMKW+CVB8WjGgcL48c8KUppZMWXyDVQPUEwxxm2Je
beMCw8OA70Xe1Xr7Rrj9O4/4lAjIW6/XNx+m3gUBYmHKWD3NJWDcXW0c9bNbHhRJ
HWb4uNBqojL4AtD3Gmqwru6w/wGYSKvnvZKoV4xMYOY8BRdca/G5+FUuviFOerNi
CrKHMDWkx3T1jRfyh8o+bJ374jiYLWslgofZhXgq3M42Z3gdf+Pf16KTHg4/ph7x
EKz8Ts4xBaFfD4JwQ3v2L1G1qTZcx2/XVfHymX6OOYttzDrixJ9rxkMsUtw1t7I6
sOowVZ3C2SD9SiuIDR6RVk834UjjAWeMg5CJWkqiTPp2Fk59JKHBhKHqUGywuAv6
uEyVyr7zzDWnLwULWHLm3+GPL9AMwr/aHBiFpr1rKBv88q+4gLgZxdlBTpS/wRVU
bN3BT0j59EFWC28Z1nEPACF/6Rj1ZTx/7gqj00frBiXYZbJnib3MW+Ioxy2/qGrn
tszaRSwK86psB6ijppOD8MkIvscIy11gcg4YL4F5U8lptO0xBGOxfBm9APcyXh5B
S1op0cTHjkLX0pj0XxtGZYodU7wsimHX9vSXtKan16/YmLiaQmXFYxnvlDezx61H
tnpQLNISsmRZ1/EGNKkYKsOI2uI51kDHlFrbE0rdOqzxfb1YHmQado0J/4wlYk9n
6lriKYteXdJ42xqA1G7kjOdpGSV7ZaRsWqcrGwV9KhGVBAHXusF7ppK3H9IL/BNf
KB4vGzjpvHiqpuUR3t72nL/z3wMyZahfuI28XCtil0DQWPismoP2oUIkLChItOLW
v1BXClF6HJhGGK67ceppDQjSRvr1/OuJ2GsCW8SJihe8PobNBuobbMyAhPjIxHOs
/ZEA6umdbGWBC8n61Hb2ROrTTaE2lq9SDWp/S89Q1ZYyEGCoEH0kNqxD2YulqE04
vM91K4Gez6lq+NzYsD2aAResBQtSBwYKypy9v4IxhwWODEMIvXbZMoYpCQQjX+Oo
iKz5Iaf6eabPdBUd09NU2QWPc4UjcFY+va7Z5DQHtG3JnquposAYLWz/VwvZpap8
OjWHgFkDs29Nb94HVhQSE9cEU4IdBGIill1pHRh69tcks6lt+sn10b3gfdddGRnU
W9liH/hcR36coTTF2JdC11B3qnvVr8He7R34RZYgDNpJnVWmQeeUpLxTwBSfsT43
3LPEjsRpQiOBV1+ImuXCsE6VVRV933E38IJEA1+6IUJTFRRHk2t3LNkHHXQTr4EY
LTRTgNvWZH5mLg5qTZeXG+L3u9FRVXcmFuc/QfE9aJxmo9hdUhGGDndyZHZgPuNs
OayDQ/U9lG935jtQK3eZGqlF6tHt+WsnhrL7f+CD5hHp2pIhYogbid/kXZU1cUIL
EtoEKk+oBoOWoRQZEq0vmCOJOL+auHZ5nEhMBbX0ekVuPMNW4B3N9AAv5NWI/5+2
lyxFKRq3kjpZgmkDIB/As4+TBysxTCL1mF+J4JMUykoDwQZ3PVQEJdg3z4poHFnD
7YlLrZHrJRiCBMU4ebZ+FNwp9KdCp6Y7AC/hv1/ek1llUnpHfgGstDMbsvdiQIdy
c27jX9u1uacoRAN9aSydjCh+D7QbEiZvx8R+njj37HoHs33vvb9u38DhFe8Kkt4v
39FfIGAGFQ/406RoyTmATzv7G+aeZP1K6sMQkZiiWKZFbknRIwPy4YXDffwsjrAA
2PybyZl7HlaUrz46spdxJ3PjwJr0kjouH76iAkdVzuaM5xAdvv3ewh87o8OsAg4r
k2ozVnBinU2PtObTcDvOcifRY8TQUWv7cQSDF7mRb22zM3rneseKKS4d3xHP51s3
oxlI3jwoFGEl0JReMS1YlmsmNjtSmXTsmLhrexkoO36k6eDcmNMcMTdP8MSt7apg
PgUsMcHb8NGXP+x76BxQkpPApb2OrQukG5A0CJdVH1uNZV0Aea4c6cLWMa2En2fb
UIzjOM8dYKb0c19Ny/UPVudsSbuKj8Pli0l1P6aQoq4KHUSS98gjQfJQ0hUcmyQH
zRWpyPlHlJxdNaQrIXQZQamdQeYXSOyb1Soklg67JrSTdz4o73XQdpcJKL5oc3L7
W1thPbw5TL5rVifOsi7+bSSP7oI6UWWHf/YrEvmlsNtNV3dPC+ZPDo4aPZZS8ml/
rK6PLBaUVojS0YjV19FHeEL/fJNVNPA2jDVMaentmfqOzeA2BbF8XBGk4yUUgGOw
gVsnYpwK/ZS2rIqrwNTLHwYVwPt+UIFHS//pfABXv9BJuQGNNhSWpu5LBDdNsAdT
Lqx8/+PWsRrCJr1AB5+7xRUCjGXk+1Bq/LAHhz0bunLrrG92obf+u3ldc5QWvB1x
kJxZkDuWaT01Xo6qI9qq8cYnVC+iQjmJ8VMs+PTN2bFc2mF5d4dF/04gpzfy5wvG
gBA6tTCijac9aBGzm4ikWc6V20mM8bG7Mw5JeCsXuyOS5Cto0/GD+4rD2Cp9R/5z
OfkIvAiD5KDy2HB284SzYfJOu5ybo/K893wL4AI+wCx2Mv/9PcLqWTRAaDwGxRCw
YkP4xVKRw6XW4SIoQm6FjfIZeI2Dt8S5K5bjMWuTH+vKvai/PhFsiYTd7taBY2rG
vM6fFC9AQ/1efS5K/ks9vE3sKWBNX3KMxbzt1oKfx9AmzA7/jBGw83uxk070xyk9
KLudR2DyVCnI/NhqS+3fAfSrPdYWg9Eu35ft1fyp5+Q5cgfH+b9htCSOwC6VrnvI
6uzU/3swNnat2zJc9A/E/j0/GH0EiqnossdORLHTnHdY2wNUZGPOrMseCB73XQ4P
bN4NSWvSFeNiElZDgYc8nGprna5RlI3QbY1uh/KdIPMjNrBsLiEgG+P1+aqwOWES
MJBAcp2syjQFKac1Ts49z3Gi9ihJ7EURoK+B35CKR2ckWsW6OjgXPf8fU31b+xN7
2zgYVNZVSfNifxsEyB1fGTj+3JhKlSJI0J6l2Lpa1BRDNzDgNO7Zy/DZMkWaZesV
t1+fnIqw3OanVdJD/QJEsVmHHIhIhvCFEuY1A4NTrGXXt+OckzsOZfteqmisizjL
6tXAEk9aqR+P3f7+oYRYRAWwScZRZLmU0+ktWS79EbUQCimPAiV3V7fjLWELqIL7
e1v+cyYPI6G76YIHa883eZmdho3qwQsXxVJ3nglUfyX/DKC8gZKKyTbKCezDhnyZ
toqSsqRczcsVCfsc5QxBC/Wxsld1muL6TCyNc7jB6NehAizpfYRhffj5oLEg4brD
FzUuzsbtAycxjNeOKbfCLrwpMhway3341qx+G9EULPSbh2q0yt1pzLIoNpmET2F1
x/GOsX8hGW2ixglJz0NYtU+AcP/UoS6KxFvp695uNnmrHRg+LenhQiUb7BB5TD8K
E5XAXdRUFuMm5PAIgUZLqDBgxCHfsi2oE5VYeSiM1kX5DLwT8gPSZVPFWguZwyL1
Nmskeq+LAoXrouIVh95Q8/wh2VJ+60df73PqizQ8H3xdhDAE6NZObY9hcX3uqrX6
pvgc1/Sn1sly5DpjYsWxQEv2VQ/asCQlFwbNuDcLkXuuw9eZDiewDYXez3bblEqZ
cGnRRFKeCipUw8fO+Y1ACfAkdcgrBXX4gXhFtEZJgBsErGb/QxAEWOq7aylQmOZK
tbDRDTdaJMDu7b+EYUqsrk8TfPrMwU6DPihEjqnus068EAnrXM9EO0t5763Xtvno
i5YehM5MS69UttxkYMUjre5D6orMVHb+jdVeo81GPjkRe0D77TO7ZvLhedHmVR02
y7rQ6rAJV509uQJ0bZt4tZlAExEpZyv4L4UjtcpqpSe1UePjMTXPANNSk1VX/vJ9
Gn4T8P9hVRBz3CFwXvVgXxR1QSVmqL8JpXB9GUshzOQtLzQLkJ9S11DWZ8n4rIJc
31FyV6VQ8vs+A77oeYjodATA0Ez2wydGRkAoNJc8MPzlAtsRjlhRGmL2puaOX9ae
i5Dfx4NmJpiPfBvMrxxbJR2GXpiUTnec/NSLsnrFGw9f6pMkr5gaHcQsE/IIAvyb
KLk+/sHgEWORc3//r2ChBw8de+xea/0yaam3+yVofc2A9uMLrqkbV6lC5l7g4Egv
SPVqAGN+qJ5O/qX+h4XHVAEVBvfBDibaXvBEpvWHGbFT0UwMhWN5WFY0kI5yGdeo
2FRTVvB5yYbAtJhi6kilckCk+ip9+IPC09Emt01lqb7COEoe1bLjYF3jWaUxYPb8
aUye5d596pgMtSBgfQRMsL22bmL3IV0AdkkvEq9K1n4sFgFA9BATmyPEtSL/BU0I
lBN3aYrLxmzQdxdzHGfcDs5EHLLAMm8GACVp2w8fMjHlSsY4kmkRwfCJOyRvJ06x
Hx8V9QKw4BOiS2JQryS7tpibvk4WHYdks03bHCkfOAvqNGaOXbHIsfPypVYsE1Pe
+Ks8nmCndfiKCqmnofJFMsatrktaap085ZbUcyS1LZ7YE12KyuSYTG5KMAaH7ioo
4sgrLyM7TYExZIfUNCO4e41+UWdH4LYqp+MfwZizqqkMdvpTZBJcBvsYC8K0o146
s9/5PSUqXDSBKamCU+ir/HCSq/aaU8XvUvabE3O7WXBBXDbIuOMwQVthD5AANvD0
3frAyRyYvLmisCAnJTm5HOHgm8trcCfo4g37IR6FSR6lteYQ3WWYZS8pblKddExX
8SXDYN4h7t//TuR1GcxkiYvQlaF2V2KFfhe0d8LZUTbxMMWmEzgyrdMx7xf/soK+
18Z1k+bchSXRpyP5OeQMEtFm0pH7RlTF2oLFCWulZsW4bmRW8Vlp6oA8kewo7EFR
jIHwja2ynFmlIU8FICnrYJq8misk8BXqqCDLyya+6YMzu8CjA/vX2MHtD8g99fAD
jJpcu6EMvl7qGO5zHCUzwkpL/wUTi5TBcpYvZhe9e9OezWffZDgRisLgs4q/t1al
dcGyFjE0nBWVkGH1sqOhu0wVc0yJFtaYk7GKyS6GfZzmsqjEsLRGsIA4MmyO/jOY
Rmc0eWAv7grG6/tjkUyGpfpPBxeJuxQ+a9gNqQEb0ffBThdUky2+PRXkoI0IOVU0
pdWXk3nZqns+OsHzxIYluVyINB+kWi+NgDa2yjetS7KczJNOZnPm5QZ/dHG9ok7H
Cm1eqid5CEu4+nPzyieJTf8/6PflfI2zSVVCpO7hAxIUjwDpxLnYpgXkyI/lf7/D
Sl6z5YY0+1LxnaKwieoti6UCfL0/e8sTVPuuVr5aB2GKLpI9QFcP4jZleZ/oUIx1
w2O8GJtTdwI2efAZSdXt9aYm7FEmgLzC8UsWIa8lebqU08zi3OiRTHS39P0QiPAW
8npc7ImyISPLhf/+ihETnzdeWRHxQ9C254oW2zyJPLDWjnPaGDqKM7dzqp75M3SY
4pacPgXcplzN6VtVCFCgwboGF8YdDXJbeGLFbXhF5toeKRvTBfyR8qr1lRizb9ic
xy7Ux+spin1ytLTF48af0GJ6nfK3GWQ8FTzYRReOACzNXn52OOVQx4nkumzUzXH2
G4i20axltA2Jb2t3wjsVGXU0nAAEgZU+hXSdZ5TEj0heE9ZUrALZVxuSzTi3VdbC
rk/U8x+7rtaydAZUBbZ5HxIq50rGPdbR711b4I2X38XEzUtPBggrMyQROx2UzeDj
PNAlV9yrHvEVxpuCGb/zQ+08c1rbeGJaqUi/JcfQNAkKCGVz8rECRHlakVDdtcUX
T6zRF00nkl+pJ6+lzrlxW2iHpEa0xlQV91xbvu3MmiwuN5kWZBea13PUaI/8qQUc
oNUtKfQ/kaN3Hkj67aLjt8DrV5EUiWSOWrjhAkRlwtulmJK9jxeecGCam+fpGaP/
m8VNHwTK6ncFGx/Np0cMJbngcnum1DUh5kSQE9kbuqZhX7wPa8DJ+IvFxFv9wl55
JW/PdNYuG0mVtvCJnCbPy6Zeon+eWaO6umIn7rfLnKiQ5znhhqhi5X44Hp9m+t8H
yhFnVNEkIju/nF/Is6Cop6xiKJTyMO0qa53s70RTxUL6gryypzgwZlChTuEktOa5
OFeE8tyDO5vfLsop42y11DUwGXOn1Deb6El7o8CLvOO5C1mtnBu19DkuSnOrI4HR
NJqwCFgYyAS2yYtc2icx01OAevHCuUzUVakgywh38WXqCHW/31bPa//zMM4cBg2/
j01wLpHnar3jvwf8PBNI83mw3QVWSSF4xD1suDP9KMAV0dsntkhWqJnP/ixPUynB
EhuLkTS+CUYj7G+qVxG5dLI9IDLRltmQ+sq8Fe7xEaSCBp7ULN+zgr3OzkdDQ20f
1tSVOqee2RBFXwU+ioLu4stW05BJlET+DsYZN2UEvnJhzyPAUsjI0cmgYqWQreqe
dTD91/UHZ+TcJPFezEI7GAjDcp7OVpZ7i3pbVqilOxPaMGx52tP00CPUqYn7g3Bx
KCnuwOIS/0sGGCr3DKyyMxklNdWufUVryz+Aab5msgtlh7rYb1lrjti/VkA1kkch
3DB0oz4OpMpq2nRyW5oyZMQuZg02hLe2aHEcxQmjyZTIjI4x+nnLD1F9sWx+mzWr
fWyzsz8ucOVT2WcVufoTdS0WpIclfyhBgIyD4lhzLQxptR+19LX97irJPMrWGMco
kBXjV6garSqtPnRxRDX3fxjhoDAMynUjNvTqaR8OSN4xKkRutX7lZBpMexl5FNMD
Jf4VZpONi8CqCpNUxF8KJAb141HSJhg4hg6BSHXPD2XHAWqjxChgNkVCK0D5VRyQ
XUOUdrFjkv+v1mvW5YTeCDb7aL0Pr4ZLQpP4cvMLPFWGzlihRG34aR1ygD6ZiI/q
k73B9meE2lpoESbw1a4bGUxqhY1BH0ZUlc5IHu/grhDToRs8MNGDEHqlGKWy5wao
pUxErJGICJjkRfdrNRUUO/gc4dymkfrFRZdQu0T7Tp6OQQU5hIN94L5lyWn5jy5c
XWqMQ+fPJRmHPYvLifwUw9MDBF02NauzdVKzFGjfrIRK5tekZl9AZkaf/c6W9Az6
nKFhqrGuMOPiaBzjU7Ng3DWL7x5mLaA0O/u8BI/ewxxO8alHkBlvBc/D/SrjFZ6D
sOKszFzYDEyMhi7FtANdIpA0Z0jA+nhprw3L6vrWEd8/V71qY6rbSZa8W1CnJF3K
8dJzM7iQoJUhyPn/+lzwOkjcMoL+kQoR21wiwfEuw53WJ1DPRH1HEbnVN4QmqIhK
bw+ylVf1xaoDvP82AHI6t8x9Unih64KYVdz8+COdUYwlZSN1O94XavzR/S22NQKe
OeWlKqfL70M1x/OqLDyMm0umJmzO9ZqsmrRQgJv73jZXONyA5Tr3btoUtp22RylZ
fxgn/wpPJ4yZpEq9jYZdUZLa6YqEh0ig5KBlpAgO+aY46Xxc7RCHhg1It4q6EqT2
l6WEMS39Hzh9Hq0HrEAARKM/IN6oa/0RM0ZKDK1xFDlS2DmaqkH53qQ6cGTr642O
B/WR6su5r7F4bsvSI0rLHAVAaGgGT9LzAwEwdvqbuGvvwYzEEFmdYgDWVDlWfQT1
9mY3rplUVzEbTdKWucNcf5YAYMKjWgwTedVPurt9afv6vSyoYXITayKMmlMqTpbB
tE1TS/FLQwTLDIh8+tgiFb1or/stHh1rytoOwjNlyHicI0EgL8Wgx0YB/y42C22c
9GykQDHMdv0zGWG0/KilVZn1jy+NhfrIYt2Z50VZRdTE503LjTrCDygJhArI2FHM
ey5fb7Kf/IMDiahgwKvAn+Dpu8RqnOlYpuYnJVcLeasg/P7Db1HLI5TxKegviroc
IwdIT4H2VhLzh+sy7VY9pr/lAx6RHm6SzjXYGKyVCb2GrTJaIkz0kvN5LcHTIXjW
MiXuKH/TDSMibiNietAFLGUgaFKu2vQ0YDeuVPCP83bzrXJd9yYN9BpwaNTC16wO
ivoV4kpj1MCy2x1Nz+RC62P9dIvIHHlAZxwYLjFiuxy2nri8qNafBuyfFAeRUC9+
f3wwGLxQbpR9CyPW/G9AYZ94yE7dxyMmTblle4ksTQYlmbCth5j1yISBeQ5QiL+Z
L4V7Kr4GqWnMLjvoRMRREyXtzI4v2MCPCFFh0gnFeczjry9lP72OqxSElDNPysNC
Ne5GU+L1akhRrmRThGVYPJgfy/5PNKYR963dTW6dwX0dBmvNZOkeLo5IeDgyoBBO
gndqHfmrhJ9cR3vdfGvCiOheKGakxSrVBsW2acDN1w2mSrULB1z5HtrFNMF+fc50
vkWSq26dgYN/r0mHcvNDwyWHs0O3rGucyRPJVQNYE1gVunDJJfdsttckrxndIQxz
qCl2ZUJiHFQJ7Gh7hRjDPigbLLegIvY5HBo4hqu0tpKQ1ABGk3txqt8FwGLrNDk2
Mdqsm056L8i4pj6Foj4dHMOFG0Ae8j3u+7URpZcSxWusVmujKAyQuJVPTfiDLP91
sFoyMsvLwa2mJKSWeexHe/XRCgutRPSwUdntgu6g2mwHyuIW+dfzaJHrpyi04j9l
zo240KKumfRIhjDqbzPOPhbBBEyah61b4mFedKtTPUuT5SVfl24GFjgXyPqqJNpO
OZBvLQec42ejtUctEilnfaRAIaOLpxrBtCuMro4C56wAwJYgO5dAwq01TGpFxFvk
U7WEhVNgCUHJdzvGeK2+zeX8jtVEr7ZUFEhuHZW5O7/XatKoARvFEqTZkwgZPjwN
h2fAkueZCsD3960iT6kFOTS1Q+zbEfFImxkQAhAeWwnoXzRjUTskq7fJz4nNcSqG
SH2BuljHK4TelsQp6WASntpWZqGoP4Onie0E80ZLSRpZQ5YPW5TNoVQBp+m9Y+pE
siTxgQIROPyYrkl6zgNWIbIdCB1LBAtj/aQEfki0uJklN7CzxK63WlBXNvdT/Z/t
95EhuRxvEMe5sxN8ezqfu2iS6fFT/w/PID1N+1EfGGUi918GHPsoTPoA6d20uzbN
bbwt/51rOsVVtb7OBOcC3HrAfNmEK3uTSGlfM0XZBydABt2T7dqmAkQj94jnokfp
fPT0cYbtklI/33oSfogMx6hihzsxRl7VWEzWGV57mNqLAh3juoAcwScfOemRlL7j
6MPqsvi+8XaiN7wrEn8Dw9wyNwIZ1BV5HipD5Ig7J68qsLX0jvb/noNjpAzAyUai
1750kTLoI5G2iKv/8jVloi6/PSdt0h8cGrRKVvRKojoQDrVhZ/mVTGK6eWroO29h
H6xmTdGgBT+HOG/t/RU8qhcKEe1q3IOn6YX97DUQiyRKaRmEMraiZKTjnjKOfM/O
KVqbg2AcPi3XmlSHZzYs32Oo4MYyAjDhIDGGc+OC7s7XRJUF3zMVi+91gMOF5tl5
P2Mc3iyDGWXEAsTJ7RDahvbJasi7BiSl8tFqyyp+ZtwjBb/PEybKr0y/gfLwu8Fy
rQKPUMmSfkjuWm3HrXkZVZod5D39pB52ueK/rR6GCz+9g9MQaoxIhkXYWobHv57a
5HYgkSahig555+xRrnjOLtqCmunrb3XM4XZ7k3fCSzKTsmBsi+CERQwT++a50YVl
85Zrqhru/YyGBpRMWEhOJWHxD2LH6tgZh7AH3NmjhohicWpr2AWD5sHQQuGXagWk
yHm77EBGI24DlKvziTn29D/ClYrETquQgDHgAsD7heyS74XLe59b+BQKmJt/MfXw
ECip29R9jMAnNjjdWVbk4adFKHcBJb0rCsLIrOHDKqvh47j84mdZrE8HlPCoZ94k
/6zXPU48JuNgCLymWE0p1RkqkwfGoddLcIbUH433JIcgtn2qCGF94364hB5cFTX/
IxxWCUNec0vyIIDxfMXatyeF6caF8D38mxhqH62qoaqKoHQhHA4qMaWXqxaX3/cS
mbsxOW/pOzUPNaL1ajonO7K+hdWpP0/EQwQRt176ijOYcCM0grwNXawm48vRxq0a
oHrvAPDLkPPgUTJFD/VHjw/774/+f+vY/lIVHzaU1Ci21uwDbcPAr8Ob3VOBNl6r
3qPV8mtzQat7yHegZQVfeaf3fudm2AHaUKai1LcejBiVXNYv4iavurPZHzKplN4V
XAYHsvw8tUIfvAVykZHWfDCK9kFRd8la6L9DIxhUW6j4iK3UeCHw1otwfaCOli4v
yoEYIJKITGI9emWNp8cvG2Tsvtqy9NlN8zHdXefORljJX5caCcsUOVIkOhLfExm8
oOSpcRVdQbgjqjScpo1oRh/1cYrqtYR8osSrREVTvoxw6QYf5OfZKw8RQ7Npzu7Z
tCIcoAxPl+gsaVtZ/yMkfMggTo0tl685gxaVTb3EtBz2HdXOqkfEs+Yb/WhLE3LT
o9148J0pSAmX6HyaOarUHSFIIunaHwq9d4eFUcnyQxzo47O/W4lkQdl3mWpHCNGB
CgVzD78vn1yBYoowgi1PRzF0S2/o1Thd/F2jIQc/j3knXYz8koXK7MEYJu29faZG
7YncVTq7Awe9WFtG6kACSE+B9j5wd3LtrCgqgnjWFEBreGWOK53u+3SDY/bQHhHx
BRmUZOZFOp7o+jv2/U7gy8kGIq/4SOa910c2YQTzEgslXJI6TOSY8f++Its/w31r
diZozCYcCddCGMx5LbvCI6XosKrasVyrlwqXlTc8mCVrY/nhAhny6AJCGlTuJA7M
qmp576+MnlVUEFJA0XB4LcEpJ1SYZsUoN87rWzAqw4pK0AnE3s8nMUYJ2WkikzK7
braPFtWVEQxBXL8Inx1rLAe7MR53DUIibG0s9unke6/vo+P3JBS20M27E98Mg8jb
Q2uLMbAZRZirp6WRDG1Vo+GukqaB25/xnCNYOqcxcGZvUZkmkHV3fQlJI6PlgzWu
RiPRbdHFlNGofgwtxlLhp7QRpC5NsyLw5JzvUbTatGx3ld56FV+NHvvXwHnzGYuv
F7CSuoEpVAI42B6nObA04Iu3TO+lFAdBfY9jjI/gjb3FR2FakN4SpGRf0jMmvfdI
9oms++iy7UlqLNc8wjhoe/L+pNeZyhWGiGnYzH/DJbrqNyAE0uiKQ8Pi//HHkGJl
kiJkmdoBQnTO18aLXFhyEFhnz+GYgOn+mUkcTcAWAUZUnN5OZhikn6bVmp5hqKNS
iU0k+lPakllNGu6KG3SZSU0h+VPS35pDnA7Ez5vo4SW31mO9LtmLMvy81Y6c36tL
Y0erP2LyNz9Vo6GFxu1ho4xS7NpxWMdViEAn58JbfvC28vYCUeQP9a80SG7+8pxX
zuMXBvrwPXfbmHRIuHl2Y0nbR+JQXjAnrr3lVABh8QZsRl29WJ0Ax5lrUDYFdziP
i/feste6yLz+Ut70EYbsWfE1MrIgT2im2WjRmfNbqKfOcLKbg1gXNxva0EJOw+Ia
DvyT+ARSG5C1hDD90Nn7NNF8CGRVnltNm7arP6WWknGicaBnSuTbMFX5kfKl1QaB
UMrj0q1B0gjdA39tDahPkf2xSM08a2nzntYzebgVJpfWb58iM6axPHgVHQJ4rSVi
27JTK8Er8tASe/7wcwa5o60vhNFja2FJXqRQ7Eia9M0IaDTEdzrPw+e45/YdqV8n
UwTgXCqIhWBlAMjDPWcDMXLKkObXMuOHbbdm3B0Fs858SYCJt9t+p5IflGgIglKc
+P3qVnuJAKfbI51cQEVOh9jpqgHxw/AslTRLyRqaE0UxFXmpZC2PeEibTRxYG21n
+Hr9v4Gn5BMd9TL/doi6fOLIZ5zZWB5tpEkwUt1lPokln6hzPp4+At3r98oLF4yk
3edx7oIrUlo3x3w66XDBcYom8cnP6IBdwjw4SsMNrW2LumlDyNVclBK+x+LsZWYN
1SecoV5baAmQVYEcn2AgKcDazoKOWvz6JxrGvIxa9vX2xI1cOq/ZNYY3IJ8XPjH9
j0DhX+NAOqf/jccj5TRIIoWcCWsahNKcWU361ph9ajr6G7fxRKi3pwNsLwprjF2n
kQPdpr/nJu5lRzkd0SGR8X4jWwKX9GUqC+bU8r3eAWMVRvuYGjIF0dhRx9lGc2dN
YySgg4zSlA3PvXq6Ccpv5dF+/Fwh5BD39+ISA6CjXqhaScYXwmfulc+KXGm5Nv64
C8I0WCwnqWAYBVqXIJClxDnss7e4kZpAQBtyevMmlwI6j+M8/65g2S8k3ce9q/sC
gDc0jZl1nhidy9r9iyeOd1Ko880Rl4uvjT1f01Vkd3vJnamsaKiIeKZc/rpc8aNJ
KPCKFqmcMPt4d2pq1moSdoKdsTTiRv7F8llqA3LJcCVfOjdKgtwciJUOLdUWCtIc
N9C8F/3SAHi1+TnFDTDy36xOV/F0kkdgIuDUSUwmqVkPmhQk9idGG3ixTltdXYDS
YjekHqmBakLYIlXS4A48cEwrOUN3++HvKUTMhLzz3Y6AxVT/tAh1CITwD2wUUcVq
JmHpv7TDv2aBW1LKSLZo9LNPTpat8hu4+qcfeeQRmecRj3wNXC1ZvMNPR7sSuMSG
oYKea+hi7dUgp9BQM3g+Z5jLXYgH2Y28IE6xmO4S5ymvWgTv/Z3S3zimj/VsRAA8
B+xPVFW5FinMpRApFyk5ZqzDld8hqVmJPENQc6zC+sK9vzpIeTz/eMy1OBSmN38i
sTm089bYDBeK/1+1APMAOO4srnyG3IBP3YexqD/Fj8bpv9A6KaE/nfDu8DFDZXNj
G+4yKZxFBLRwIyRYGwmGhqKAzK3l0TxhQiGliHp+2UzQHuE+bVSYveqJ25N/kThk
dB4vdY17fT54KBog2QV9M/jju6GHi82hd0Dxb/vwTWt7+igwaLK4q9nM5OvJRANy
MAmE/NaD3oQxmmH8cGVOtPFpKIr7L8nxwC1MLqcWCbK7Ggn8Ym4oPGwc5yQyotRR
KW4WH2E+V4DWhsPTi5RNMAMnEolq2ovY6diAiboX5FERO14UD4e3D15KdGHqEfBM
E/RahUU/SnuaQa1vgKDSjur+fk01eIPR6NQ2UnWYOUXU2DddDy10RXs1R1lmPCUW
e6QKu7aiNDG6PxnJV6HlMwIv2GbHsN+QMx+IdamOacPrzCenShB4aIo7ZdcXOc3o
VX7Zc/d59a9BtwBiNA6URBjaM4rJJrwKYSn9pDztj4BZAO6c3BoAU2DaGIst71rV
TMiWUUNdrprVzp6wADaHqva2nXdvPq82jEJF9htVgCCoSFb2oxNVM0UXJrx12vBs
fZr5idvSVxVQNHSmG8OT91G1x0EScCtjQKlsdiQ5DoCBfI2ACyexywIZXaD4eHwq
r2iahRirvZK3qHazH20QmrvjHLCvZp8OR8KtZ7FZxz8jVS3aQekc7YGyVoxXyU9V
uaG8/f0496GXNTkmd4kktRSomrqh///KC4b0mphfRhOI8ORp6VXLhs4IAPHlSdoX
S6qxdHHoetHObHpm/40F+HmOamkpBEKZfXBNcLbGFCjGe612e0VK9hjskRcUQ5tW
LRSngzAjquf7TVL7kZmh8Aqu8vewCqYo7uDRgZtFjvQHBu+U+6e6w+1FnLu/iiSI
RnAIjLNHt+l0d/6kKrWE54u3vChgtfHYZn3M4lmkxOjtqMDwh1eJA/lsZKqiOwPT
2bRkiZxCCceFOGFAStfw7Z+BK3b5iGQ5ycB8w40Drd/7OpVMAya/027ZUjgEy2I1
Tn28caZyHElJ7WYcW0E5LDlEDO45Dy5cm7caXuqfG+hSJHy9E6xsH67d/U4FYN+q
2as8uMVOCdvTqlybdutaAj5Tx3fEHNL2KdNp5Iw9JX98bcSS/u8MBSfMlSh9aQ2I
QZIVHo1FdmnwwpzYZWUT+vzm/bceH9AhE2OCm9MLjPWiMDTwVGmvghwzYGSFaBg2
PMPCW0aH1D+bA+i2WRi2bMt4uQBIkgCCSNlnWYzbzQBXkG/uM76pbXSLwAlC6PZZ
m00l0MOxLdNX2Ic7cZjqNYyXlZ1YTSvjKqSA3aJmtFQ28d6sY8ZZXNxGpSFNIJrI
lym5B3g8lwBrqpBTR5hrgk3I15IZP6rR8kl0pVT8Q066+3hp3yyqM2sxKq0oHf5C
DetL7oXjXEJ7gPziihC4jD76XBuYCgUNYa3ZPTfq2MpRM/y70THchix2Y4hm09Aa
sjns+swdBFP8q7aNtpJUom/+bjbrDFgK2ufSKhwV5Lgc6MB0rJsCBUVtxvLJ/fgZ
n9ArX9rHGtXmaiOEXTmoxo7QsJeKqspgX5bM54kJNZO7HfgxS20WbjtaMGgV7YSI
PTliwVuhFSG4zLFAKFYiYNmd75i2+K98r/Z5L7b+q6HIDP3CMqKcA5YAdbiuC4cd
SURansq5EIzMlvHgo5+O+QWiB9E/90wXY3VrhR2o8ezs5d6U/NdfJ6d5wzAp+JoJ
rvWRHaz82RD+jWtAw+TL0n7GHDnhOT2U/Mam6y7T33yLLoVydnK0ybFqzGLnMju+
do6eMY06mCLU2OIh71tkIMTCeMP7UbyBs/ZYgkkQBRF7SfmDHBHNxtpHJbDXuhVE
RYJjUuyK9Y8Mjxy+CuQhTmvK8FoVF7SjLGXd2erGZIOk8RWNNFqAB6qd2RyLdEm/
waI/wOtSoDWyR60dd2IBbuvUK07PKg9fHLeHcaY3BxRtFhOhNzxrvgS/fOO/3iiu
NVjnjLFoXBJu7VAE3v9GbfH2hKNGFPCTcMoDte6O/6qY7t2woodlCeXLiz30RnJX
n1DaPMe4bCe0YKkgb+/6GE7sMxVAW/1B95C3GJbGKwRcWMTpVFNUmGsFBRtiwtlT
eigRsMN4cHxqXwnC8hnImB5OkL/x44dkQgWOf+TnsDsGRbRtJxSvJMGTzN8bIdtU
9+K/0h8PYDgOMvSUtZNGN1oRhfAQ3Srp23CkNcNglMI/8mIlE/uYUK1aNN501Dj+
T756RffYhzOlkagpjbEXjGavwNnczslupjIjmvUzh/XAIpo6NmDEoTOI6uYKLMij
3mE+RORHPY2DNo2nrh0qChdiqwc/8d8GWLJcCzH5mB1F1FhWrd1UZh22NWi/LL+5
88cfaKZfRBeunU2tNvTBs9xhX0QRq9IRvTFgVBsYDrGAo6fwPKrPDpLhx3dKgn3B
q4p+LVpuWbdYa17yeGQ+T5+DNQE93z7qFVO1dmGBCS2Fm878v47M43eoEJ/DArQC
xrGEWoOWf93u5pUYyxU3Syu1p03BHvS88S+H9gTscE6G4bbXMasQ3oAKhaH236Bm
fE1A4vWto2uBFna8xbGpKEvbubA3Lhk4srfe0vwzBA6wfBHws8FESZfumL61rM3g
06KnzxujlDhsCocQibsVb8GIOomMVUjZGxWynfZNv27CcAw7Ev+OZh8w/AeR8CWv
Glzmpbk+zU+R7weyX5gV2Qi/BBfCjr0Aqjquf0qvBXOBHm9IxgrgIZH/nm74bPHF
559kQxXOOyTpBfRC4GOwQnju3+dvcKRIoRkd+dvD5q76NrOMs+sIVtPC6gcy+8HF
zY7Yblc5N5dp9+WXWrD7rhxXY5A3mJYrqfWByD3Vv3WGRjgHs1h8vrkZrR4FeLx1
zdGHXRFOVetuin/fj1ud+oP4n3Y1onEyrHhdjZIZAdRmnBVU0uZr/4XsXho/vl81
h7uWunss3uNRI+NswdrBbw6s1xZAH+5Duy8vPdjzdBaKwSajM+emMlD8+xYwM0oB
+WuJsRn+N5SkISMI6cHLWNRaxfG94cNvWGjFEmnjblnxBAmk1h7LD5CY/z2L3LMB
vCX3zZlRSHJFfibjMrhPTxPZ9pBbX2hrME47XO3khB0Rwl84sbGHxKco2ay472SP
Cl1OEK5MfBcPh1V2HPzgaTx0xllWboVtd3mlv0vK2tUdGMIxHbfk+uBkLE5nbfM7
BnN3Ac0p9xOhJgdZ1Bh/IcWSo9/2dSO/cxMybWbSIw7xUOZtH3d5MiwYbBa+IY4N
9qoY2K0tvlIOCM0e18eKS3b4tUjZgW2z5+CjtrkPMzNSK5M9ZRhzK78gOPpSJeiA
GZ1h2VkTylKaNgg2115E0Ors+4hdpwATGKCJCVP9YHj9Dp1IILCmd0XQqg8fVGVG
WCL2+uCKcZg+JnFhQY9WV5yt9FKZRRUZ/vu7uSvq1VBwqK17QG2eRTfdFvvIqHTV
AW+5kRgfAzpxxwZ8MyeD1jv2qMc/EdRmdtdH7mhR3vAktOrKcn/Qk+bliOpLYSPM
qHJ8m/dK9xwk27VgfGmqrq5mA73HXKLThFq02TNi8HGhe6BtQepWVnoMrh0icsUR
sHTyBxav86VdzHHYCO3WXgktE07evtXxBriPg7B490Gnj7Dy3Hiq0xKcnFvaYwDX
505+zv2E624npnpSkU9p4Am5As400fkXQAkNV0d+vARlRN3PY/KQP5WC8tkspbnR
cYrKJ6g3ZluJAyveVVE5wgMQ0BnXuXFaU9dblauK6t4SNKygWq3NNghyYfaKfL60
AB0GPodCkQHgPLlmleP+MqUlyMH3OViHtPDNBFtyXJQmXyvELKR2gNZHqAfikAuZ
vnf0UI1xCAmDfPUKS6xO4hXuiLRZ41O2MbkMSIzsJwUCDny02o5W1/wnPmR6TS/2
3kmg4yEronuN2EYuBzF1trdmj9U046uxWmwCRmC5lUCcC/Um1+rCY5CWHTEq1zgq
uzdZ8ugqRMuZpFLShPuSW/9z/BuLSmCMravHt+SOMBbWiPvHnvz13bkk+y7ah/YU
5PS/QZm+OlVRvdksej1zK1LxI3zDo7Hi9nrRoxpsGgIkCjzROf1FHXBzXWPjNIfT
qyv8iYRtVcETrkdw85dDAdRBINxdq2JFwqhzWOB4rEqP1GHhktMuh55R/xmKujiF
9jEKlcQourgCGF5RK44R+QkTzv8Q/oWVpWJRrhkjrSSib6TpE8ooMpjfTzUSiBsu
wjgahgok22JzAOM0XaU3XqJpoR2rURu0Vgq+9ACm52nrrDasp/fy+9NTxheiO3AV
4J4ynmYmjjLaNY/94bBGc/5dFGOgpl3n0LBnmjymFR00sSi/+gFdGdh/mJhCICgL
9AsLR+WUvFMheOiyDY4CE2yuPHjqwZrxcUvX/8bf0DN7BcEdaCglpYTpUK7W4OFP
g++xuyym9004Vup36V1RZM/6mG55svJvYK5SJaeI7JGtDDQpTXqtAHrZdDaCOnm3
ARBqJd171Es1XPf7868hSB1xVv7VCu5HHrPUIxTAckUbcETQAzdFzeXc1lkXanVE
BM02FN/YTOR28AWxo1jx1lGh7YivKo+BSYBJdDV+/dobBxYxus0FpkCGslNGRDYZ
pQs3KMjC6t1eK+vSiaSDAK27+DzX276T2m47QU7x/fvrQdZ9FsnNIFYeriotQzBA
qEgzj8EpaCI62nnP+Oe521+1vZRSi3u80kWxQk9KGSPX2gXJTxBG+PNAU2QMunMQ
V0kXOjXvN66ghs5dN5h7JuGn5FDesdBUfKFxA4EpOn94JGV9maeGnICKOFpIrYpo
HqxjFbBQR5Rr9YARgPdAJb46wZf96L/npoh0tkC+prc8M9nAyl1Fidzm/zieqDM5
CVaMTcwjOVGGKHPOhbQ6pGpPXIUVWsa4pUNf9rWh4MztBFyklnCkreQsMekkulnr
2HH0qHuoNwF0H7MmGf/sGPlNiZ4DEOtTb4ayiRi4WDYL0DRJAlmYExUOPrW9GZiF
vv1PyrRL3EN9/6yOSEBJdWN/CQANV7RjxnicQE6ZRzResTgZRxsl6nnL1XZh1/MS
mZbRjM2d2usnRIVC+nBn1v2AC4sgvEbythRw8TxVs/RrCibcwj1emrYZyY91HUtr
0xXP4bKTT317C0+IO5shWwpZct1xjd9M6oA+RoEbn8PtJn6S+Nn9ZRJBe5ApOSl2
EodGKyuPhD8u4ad0GQwLqzUk6JdsmwaVsbpk5ojGwC9eIkfuRNg+2i1CDLifDsr0
0a/VdjpYkLIjZSSAlTLIC1I0qR8/J37qYeFxrWWk0ORsHI9BtzpLMMCoy1rdHlqN
3ow4CVh6C/7c0jdL932kYELkTzADXahIeCP+MDG12FuUEaObcfm9lcOs9QUc7PBK
G8P+fiMIQQDwOxLiN1Yi+Wl+y6NGkw8RPFZn/ZS/IVxExE3yWU6vljKeYR6vIpjm
EdjCi4krp77J883eSlggRgDkgFgetcCAB53lm/vLPwv94Gf0bn/78Oa8g6k1XH4K
oEY+rFvpQkFhRXUO8lPxC7T4j6N8xBEaVscaGtFx2SXdYWHKRD7wFKmMxKDFGLzs
LoVdjuXER2+x2hGDxAYiYEM52n1liYHFUP8+RDk51YPZk88JA6EG3wmsGXSQI8YO
dE78zz8vD434fK5GHQ6oT3wmiVtAz07zuS8qTyHahgHBTVUQmJKYTY2W7MWU9IxB
iej8axQBY9m/Bz//dABheo05rskBUhXqxOWYt38VqF7FXdTz8MtxMYMknX0W/wdi
9kBPVZe9xa5oHVc/MdbAUUJNZ3TOw8VMDth6j/qS5BmvFIYOq2Z0XLkXAKKF65Rf
cfYF5uCcvJzjWgix7R3+/ibUeJangYUQf4yXKtlmY5hjEN4klE1E0MGhb6vwJHqv
oI+SjnkEepkm5G+3tg+C0x4Tvpj0jdH3qfMYXxalZN3P4IT1fLMhVmRRyhS7NY+t
4bSGF0aP9fHGuBNs6mzqfOTOd8WAWWQG//hsif1Z/Qh7yi5Yeru5HRNGOTv7WfoJ
ibFYndbN+/WnHo3dXGy+PZHJXoRUUAc5KHYmZejTyRZsEnFBdgc3N2LPPu6nYGwk
MP4IdC90X8/uN14v+DZ22L6Ps1SQ0LPVjsBlKujISrZZLXXmVmhBG71mHc1w/ggs
uBAgx4I7Z4nHv96eUQGWcz9ldQGr6lNGQ1TBhQT4jnaUIK4eSg03fAqxQKrAnRGH
+Bd440KEGAXqMxO8JBU7bXhD5TXdsIOM4WUAiLEgMWe40/4JLmd/TwR9RXauRUD5
w1imghy++fN5ft7MHfCTQfT6LDO+T5i4Mt6ibShemrEx7BLTv9xm2sYO+HLaTm5Z
1DqFB0StQc7K0vmzeRxY+/RTWVDFhT5eZdFZpScsADH3BsaZ38K6/+twdkIC1wji
/HD8F4TjU5cq4//tld3Zu2PjzR1z+vxiqrqvfj4hJd3JtgVIgTDL/+GQmnQntX5A
BHG3D4i7uZfb9buHVCrfIPcf/cbWxP3RitzdGZN19QRNfGnMKLL8UL82Q/Pm8WVw
U4GaGlOqe2upN69SBeyxYI6RQGCL1wa6oJGIJbRkLbIS8u8mHDMZku2KNpDzHN55
RRzWABeLQCwYY2YAdoPk93hbdk9lfjeuIfA75OAy81ZnBz2TcLD+7ThDLZTmsd1b
nuZuDliyWAArp8dBDPJYcZs1D7pmS0aOFA4tiUo5Zvbjdm3ip9hKgP3KTtDbsntA
4WNkfD7rdtJDjvONmP5LCNfYmptE1zV8y5iIBL5iHACVVmntfe3oHM6qyH+H2kpO
XDyWyskEgbM5d1ein5Bnb9Ag4T73kkw6Lv6aDC89DS/M2PoAa/ChS5CxZVby9O/v
qJL125ev6BLmkP5X7c+5y4/gJgKIkPvHR/ocvdFq6Zdf7JqSFpN2mAn7kE8x+zIj
lcEMUeljYK+xmc2k5+8SzKBa8PA3066MACgO6S9HHAvfLQduLrtgKG7Zo+ArtYv6
7lhEKAwkdS3xaBwpLAzIhXej6lfRpc+H0PNmCf30nwwBuA8ryDuerhtvVEMJsehs
jeesMYqFbaZ6ZlMSpgrZJW9C4xcaY8ffHyPwG0DKOhIa1r8BDMdZua8oAaRkWLQt
qM5tsFBKSxuE9yYQFuJcitMB2agqi9itXYa1vnqQ799b/pVuKO+nEESroPoViIFN
u8fej82VOjuOiEdRo2JchfohrPTqFMQdKY85q+Bvwp6JKqFLOAMHw+kxjiH115gf
na9XHcZqBCZ4QugE6svlIYcBzXX8JGhzdjnR1DyGFT6l8YYMz6SyIN4KVF+pJPMp
owVxhcx7jaPfLmRfmNJhjeiQZLt06hqg3Yvcpj+vSMd/hNdbjAz+Blp8hBMBUMlK
wO8A9THkF88bMW1YN/gHo2g+zEUvSFS/MhvrJOhvZyxlxsyHJOh9GUA966g1Bjfk
N8xGTqLXROT3PjXOs8NYaaRKW9PHiGFJ7A6GXlBwzXyR0LrB/zZwKRImNeJHnmNj
VD/VVlwwzGaCE+PdKgZnZVxP2ZUY6hV2z0Vjts5kvoNSOUptaw3oasuTEjr45wKG
S78pGsKCWnZHo6dxblxYR+4jIi9xmdkAtPbFt7e2PqUluHlSURgv+/9OgZUkxMqq
gsjsIP3nIlT99npvqZCGDfV8AyUAVoN74eIH/osp25g7kQhDzIRYIb5BKXkHP+kV
iv08YTSHb0KO0IlUeL3qtJJzY1yotu+V0/Se1H0VxyQDNdo+n/yoEE4qH71lrFve
rJnrNgl4a6wU6VVgJptjd21/l1Wfe/jLzsJAKZLflz2KPqNlb7AOL6YGUMuHEg7I
SzwZ+mnq2J88/LdYmMRjh3lnmh59KCGb8E0qkK/pbBtlMF6LeWVuwYrryjv8vbqG
8YkaHvlXuK1Fx4uKYJ5EiTcaW6s5aG1SSzQqSgmBUcS4gLZ02jRvt7GPlEgHLN3O
A9uUHCTgBTYRivvuhLtjSvBQh3zl2OtLHTMEaIz0wupuQ/0ZgVoDrYAuV1aob8eB
FvZAE9p0BwvTi3ypr6FCDHxzGsZlMtShUQX68KyEyRhG9CYhZqdWqhDiQxuYBGb7
GOn3bTITfNNRzOTNVG2eAd4FfYpJdORnnImEdUzh2+QMaBLqwoRe6Y6jOST/sDqX
7jZmLpsB1nJUPHfl8tA8AK5p1clusJQavsjJe8/d6aOfnM0joB9A3VKzD6Wpz3hh
HRRw2I1O3/vELiv3d+EbU2wFuX/5cqD855qXM4h5pnJ2A6W8ZKmLQcw5En4B+wkS
HeixcQq3Chrl3GZqHJ+6d1msWkS9HseewEDWXmiY+cIgkHXYH/ZarAMNzjVUenBz
OTB7V4ltgBWBdhbqdAeOZ7jnfZEUKaGMEd4+YrPLjwVdIB4xO2nhlzoGZtEXPaCd
5MU1I6juO5sll9nxhWrcsbviefAgf32j1Pd8GOBTYBpfrgbtpmZ1YoV4MitmPHog
A/QxtuNpBxVyKSetRULiMMtKxu/oFcBJurE2nrO9bpFHA0E/l8BYemBYxsLpLhiD
jhDiU/j1QU86M+n1ZR23mCq+/W0JIVVcVmJc6LeQNyJ7tDUVzf0e/ShwJ+7Fu0le
8Zk+efZUxiySs+0m6494clolKTl3tFd0ySK4/tG6ihGosY2gZIz1yvltM9i6H4Tb
RT1CiCxW/EZPdsQyD86xP2hYVQ5iWBdnCgGNU7AkoBAVjdxaxu4fO7JO++dveKmO
6eOH8noyp9sIWinl1WPxvFNwQIdENpIQHc2LgVNnfihvuj0mYFWvLTL2+E9Cx1fV
0ezOvHDqj5Fu/Z0R7eIROf4aPTKBy4LYZLc8P7kXJ+capSgAXBwBB3N98HTi+adF
ZVMUQt6cfHFVYZj56Hk09PRLVA4mmjQ9jmwLGCr/MSkiC0wS5RrJCq46i8UrjmBr
LEoVPM75aW5eZjmnN3jW979ShtUekrt25TA8u9rrAXKrrIUSQpzPdZF8wZTk4Kox
znxAt9hwuYw/GX67HRMc0XEXc+9RSMjoOHSrWhXU+i9aUOzH70EdiZWD8ii8UsZJ
/MuTU88TWCQvwtdea+uqC0ljZhBbG+5ry7BK7PyWE/G3Qx8EE4Xs1zuJiYJRIyUD
iK7gdlxvInHVE+OzKrroOVyxpd3QWyUr3d+IQPsPqb47p2oheWNx1xvhXwmi/I98
BEEzTZZeg1PIAwrkie+TsiQG7w6U4ogrpsLXH/Tz0WFgoqm3gUpknA/YkZ8gt0Ds
KnU+GjGboDmx8r7cb2va7WLCaCkgWD/rZXCQ9p7+RPhjDU7+yXM6UKZVU4WEfghg
oW8Fj/Ex971RbJeQuru1wFH4jijlT1L+zKuOVMT6vvu2VQ73Ga2AQIMW4cu/Jj9B
CVzksxlCeoGsmD6Nfos2usCtYgXAB24ajDX5oX7jPmDy+jcMszPHf1S1deGP/mdt
zQTIOmERYjWtnB0aapQA/8J9ua4OoIn/3IqkneYI0bve/Xu69BBkjwyxqKrXJaik
vPP9stYSc8+KwlZU7DrKmNpw0Pg8/BaUF362XSSyNOTJkT8lhEV3zrQvVHtP+Hs0
5wrUAYXSZey2a/iiKA0Vaf3PPHVduhasFRiWIyhz5MijJ8vnVlqM7sHL6LRElPOX
I4zX2GKx4G5YBUGUCm0ZOZSoXgkXnCPagswFa119XgwHTbZqCwpKKmbyarMELmp3
uJkBPYNHsCXtng9m6wXgoxTbn0LXHlLcjE2B1G+0GvtaXeEMT0b74XaSfnZYEXQM
Q3aRUWSSmkZZZCjpk6pZs2oX8dM62SMqtWtYxk0xpIUPCQazUiN2EuBqu5ZjLaT6
Tvn+8ECJAhErWyITamwbTfdP+TsMhZ0NUnSyEdSbwymiS4TMKSy2RHbapBt5fWr3
g5QjwAYhCx/QUOqUFaoBrnroxLKQ24n7qEPgqhpRS1Lj4HqZwsxMwgkIwVQukjhB
0w/uc1mde7TA9pow+jEbBRw6mb8Fi8FwgdBUsSJQ8nK8ti676C9m6/Jfn9MMBEfb
M845IXjMbsn3cc4xzI8JZMnw01t/6CYrkmswp+5GhsUt81zFFw55XqQKTCi87M/Y
B8sB62vL0WoHKF1pEWVyy62ptF4Wdq563kdWCGGQurqoptpq2g8julaS1zgJ7Oyz
+G+XD1+u5mqNl3WregtykAIb8V385K7lmjT6OhjB3Pdqv3YN4kyQtCDDePQqcbut
82P3r6vTDNXvgmCbNHsgMDSFqtpVpls/YkL2BVEzNDrHNBz6+tw+06cbeSb+HyqY
KMCcoT76Gja7mLz2DiBmuc1nEX4d64RxNQoNN7n6yEvqMeK5TajQxtdRAflPTzpG
0tcRxowqkhPpC5DV7eakXCN3rg210doIdBLHuIZgAxBpslIhRAlUmtU2GFhmldpu
xKsRAcq8bEw6TdoCiwsEiycGcaGZAFZsSbq8u8WQMSWlasYT9bhlt/1J1I4+BFhU
5TV7lpeJGWw9YczX8G3kM9UfU9zJutCB8y/2PmhSr8xek1cuMh0PQX8SjSFrIoGE
fZoRUQcJlpd4QVvn6WR/vPIRzHswcCrongCOL34+UJd0ejyd8ZNcghEUVnITEFgO
qRnA3gPmJD1uC6EfOmbMtMDD+3dLIi79XVs7hRTCNxbJ6bQ/BWGBPdegoG7vU19/
y06ldeRSWXKlLh+oBJ2HhtaDveRbgz90/QHM00949xTv+ktVfegwRvPP5W+/Rswd
fjhzGpYPT+Me0ND0MWpeja3wFuX/utPltlCHR6EHO8nTT5vXvKuNzp0M0Aycks3h
dfafuMoJ6Dm3UfAAQ76ag7THYVml1odhSbuXYP5pTHTSecbI+H9QwpYms2lZG5zL
bl7mc9UFU/KoidEtZJePTNo6kb2rd0l87XDEVkB+0Zml7zycaYIwM9OTyVNwOP4M
9N3d+QcU+nGTh1txKmkE6kAkq3ezw5Zd15OetHu9Oy5Mr7cNm2aigElsKzd37nH0
XzdNA5EPVaGjrKDAwdjvtqtn/OtWCeA7/MmWmrWJIW2OLw5gk5wvh8KzYq9tAQDx
ZsPf1z9bL89V7Qig67QXBS4Q+jE6jDc/m2sVasIuQxur/f8eRPG0BgQb3MWqZowf
Vbr/D6YFA5Xs6hnKn834cWzUcD0XOw9T4i9IoDtsszt9OSckP+suKMWW6pJydfuM
IFxlLo71rjt9W4g0lqdmdMHEvnv3PMr3TZC4v79ZyK8e7cn5OWJ1xl/1ZbD/fClt
pjQYe++TP4W2fxR42RUFz+Dx8WIgix1EBNfN9veXgHICJOdsw+a+e+e8RmPBdv45
inDtKqhEKThSoSIvwB4Q4icl6aGROc8RZvknJWe2B8rhOx6NvBwKjDMSJZPSCfoe
KEZALsk/GQfEfMV0y9w9+R1xY0qsC935MF0VYOZUZv6vVNU0iFxozyxWipoHvMOC
l4BaLCBF3yzD35E7H9r8sYR7p3ePy2Moj70jvSa9BoZ4CCzfLsSRzdgvB4vyvNeN
je2H3xHZxNBSR5KTa61MAMye3LIbHOQFAY0GgekjliPoZxjBq9ZoyVJc7kGeLzdX
BvPfPoMZQXi40+tJ+f6lRZN7AEkWo+tntXDgjXgfhXUtSzSKdszpU5xmBEmdW/3C
dX3D4busEXPfQ21VzPwoqnqp15qG8XhYqdvUhfchZ3PlbyQdc6TlXQapu0RK/41Q
h+IoIXwvvVUm4CbPlxJZQlFuUfCKW1z48OifCvg8lqTJRObl4NHQPTq1P8zUJ1HE
FwqPaCr80F5RVcJOehUVGWhPoWWueZKl8u3mp03+oRQ5y/g6O7WLVLaQ0GgMrg/p
4mHHmeBXMdb+qJCq1SDDR403ucf1cH4Whxxr4SSePhqbOetdcSJp3Qfw89YeNLpu
PfokFpGXrqtlT4u0gh+e2vG07sao8+Ycb+uRurE2/RxrWQAH0nXRmn7F7a+YnjrY
bqdgXotIUiVumVoQDMOcu3he4qF6fdDFifsrJ12Fplzm5A8fl1Mps5COFpS8HVBO
PpbdyjlGbZYIWU4WlivzNe926OFhRtFIu3eQn59Dt7wf+zVECKUwyeo7YX7HVQoM
OTctE+vYBLCWL95qnuAngwNHVlqehBD4ELXzKJTrlpYpgeBBXtrGDqtTkIEQH71+
77rggeSATbEcDqtrIB94j4emjsi0Mgn6aqm/PlyK51BpN1onlo5PYSVlnP396ScF
U0mCKO4saBJJXhO4J9HWwOuZsVcQHwXf8C033djE1a/CEPI9Cux3UkqwxbTEv88F
ipqLtyvISm/m6ZWTeZaSQXgMyFJJuELk24AA3EvjhhqfqoUyhc/z1E4xFb3edOi3
0o+knvxYvl3oMheitf5EM1532OKIM5Qappl9zTKl9WYOZXboW+cmhJ4yTs4pzY9d
RU3AgqYK7ImV/V/K3jHMFtnmPIhal5F/vdJoPARiE0gO4ArWmJHk4n0SiVsSdo8w
VoK12OD+wwswReKGInsDpcAcrrl8U0zIxX2ryTVhXS+0BkU5LBGQhQi5/cvw1nBx
g2VY2rCRnfWwiCh1pRvnnTUT92rs6C44H6OCwRGgd8FTV8G1P6yWfjOLAefFMEHJ
+zoTQvVCuVutMyTib6CGgx1v7ve+jw0lhrEgPpJM6LToFddxrz/I6wdETl347tO1
82YrH5pKYWVx2BRVXgNwobrZtzLXuSxbWIeg2pWoJ0vQraf/BTkfet3J3Di0Dpdm
eTVxIyvTod7L+uIav6JMBL7HEtuB049QmY3cFXwlGYAs1rIYOX0YCKOkqU1r/Ue3
ioJDqLGmW61z/yOCHehnYQSTmZYhw7TyQhv06czo9i63Rgy7VeBO0tA5YippUisH
fJR9dVqSDpj79MUviR5J28rYN81M0h493xApb9jy958Lie4AujLrRKUhx4oydQol
H2BmqPuAwIRYOHXbG3wTr/YHjQ/CmInidnVmll5n+e+lYyfKHQLeW8yhUi32BVi/
SNnkLSfX0Z4PftytIWbgbEPsjD85x4Xfy0PwORIwEU34BKngtcH0zDQaDtcfZ52n
yjX6eXif31qComqZ8KClelvzYAl9H/vzyLc/U1+7QsQgRv+O/FAw+7wc8PeYzWZa
RhgUBou4ZA8L/6rkChyWbx5QSIx/D8/zIofnkilRsSuf1DWCRo+Y4YcFwtJzUyiO
rBWWn5s3Os3CrmRYM6RlTtS2TGj2NP9Rp+7yW4nrbE+sH+vwm3BtqTVXGtOZKh/t
+p4hzN0e0gjSWmF4QBiWtHTkr0z54L3aePyVxxlXsitNSoGjnMY6iMREnp4mn+F5
dWfc4TkX1YsavmKHcO4j1uIYmS2o+5KfxKvv93gBVFVQY75SD7PIKMfKsUocO1Mw
geG6YkEUO1fQfXM3UPH6NOfZpj2bVIEcelg1JAlNrto1qq5TxRD4eUBZ5c4R0px3
pJPB0HF8nk0pzX9yN3CC+ym2AARNZGLYcUW8zfqAjo1pDn9RoqNC5EUWZLg+YnKn
m66guV0EIJqm+c0QW2RRVHw3CO3D2HwWM+Bm6cMu/b8NzR6T0Qe+x19GpT+TAFI4
DsBVmjX5ea1Y5+KqjDLrxk9ISlaGgXUyuGNpQ1YG2Vr7miv+JYFY9wM8ufvehVaE
c2ZW2TXCbceRFePU1fxXKs5WSj7Y3WQM/oABfP+5yJjIWwFbpwpoCsnetPzlA8v5
eRgCUMZ83ClYFWUyn8Po6hpEKUYYx59Q1vATrOkWMAasV7YO7pzItAxlG8Gp0Pie
z8+/gh9wfIxOupu4NKTJ3aiNbD6E/BC+pvFjdbys/pPSdmGoFT7x8pPCmYDtO6Mz
cclUMh6BV0EdiFfM4awtcevdmpthObzky/xH7Vi+6LmH3iI8qDPE4OP4NeXBWQrZ
MuerwtBjmhcaDN/UoM1T6BuOP3ZN4gYH+C9Qohifu8EkDpPpRHH5dq8iwqNsq/oJ
kiEvQQykOaLHUrgYIEJqkRh5xpZ18M6a985ufDTQjl+t5g5uZnO4jorzr7hkRRwW
CQ8K+citZBaQR96p25gJR+sg/6/qJ9NMzesuwVS2qHA5gEnrUp4bzsJ9qgk2/St1
rZmgwcNI08kUyt1OTOBJcDj98blNpDOczB767zTkf10mwY57NmHS8J1GFV+ru/bb
kbwWRWJfn9gWm6YpH87I/Nve45MeFL1JqyKG4IZuXReDjonnuj40yx2fG/0M0aXl
KJoNBtB/AlzmgYb5SD31Mbd4W3Lv4KVI3ZwM+wOhoVE57l/VSdjdPzdZimeg0qFJ
jewHzbws0AbjIyoF7g0O9tUBPxVjAF9cD5QqXm7ycD8kkmTzLLKekhga8zXWoLRa
wkpxdXSu/9GFNPQTaU1u6kBBYJmZmY06YJ7+HTBFBbT2XG3DxvCopTu/sICh9HjE
mMgWHP+zwDWtPK4rbLL9Y3MSb4OwvnWlx+MjKWAq+Dk9PuU+PVfGyITYfeXUxRXU
ip98miE0UQOO7EbYwdi6wq8cnqzWaWYsZWdutwH+GgBHbsif5XEa2E73GGKbe7hf
+HTZbQPdrtQ91d8Kb57CEyNw7pnnK0U0MoH0StBSwS6le+bYWlKLVf+dqLSCZkin
+dnDjIIFzAjL+TiePAMvlIw2312SObWqxYraeICj52OVL5fw6xTUeqThWC3+G7LU
9WTvtptkpbrzqJCabWDsuY/8ES8pr8JQ2ba94DKCdWppca+Xl5xTQWsehJI+LvFu
eusqas3p8hUDXa3Q5zXzKpBDlyNQX6VigbKmqmkQEKVN1FiTYIBHoYHHLaDZBcnX
ckMzUKlNy4SXNASm4bc5P2Lcv7AB2rMF1uaMfIupsskQcqEwIxfEiy6FXKR2b5IS
IudAFylSYNgII7RsbZDMktJylc0nhw5ewyikZ21y6xz3BGfZrjrfQj3tUvsGR/hn
t7bzJLOPXWKIqzDbjse0P3V/4YH/egJRE16p4cJSwJ+ocI0lgyxpwGE8ofwjlMa+
Xg2tNz27CbzG1n57v+bbnsj+WTQlQEbcQI4Wa5g8oLDXNBrchMF6eu5F/YIt7Yrk
QmvrOdmPMXF4aWTtPdrmv0tx5aOnFrh7O+oPWlVI149LlTGrBXgV1MC8FwREzz87
G/ZY5mZKcIWF4S/0IAr2L9cfCNrog4i0NXvkW55BE5Rb2TtmSANzRetLxuWDwcJ5
8sQvR5cXOkZEy2g1epId7z7tjM1ycezsVCbvSqbYOry1xxq5CIj7CWBsimC+w1o3
k1Kvt5YZfcP2rmcRCtDUzeVQupP28nvY1ER4YbzZWHJXFd8exJRexypDMNJBJc3q
qoT5YG1b+GPApe/qUWCH3tg7Xg98sgtAfBj8jJd7j6uN9JshbVrDvDl8kFXZDkuf
53gbLUVMwRJxgrJtrootWqvvkuGBUrmtIDoiGoStMQPfF6OjKANFYERx/60WRD2I
mfx2Byxggk7dtixYWBgikcAFhPN2EfVPKVXzKxvFc5/SBWiXv/HwVWMfLqdXQkhq
vBlMnwUbfjyq1+9j508JD3rrUQiDd6BvvdRieaPkTvfJKPeEk3OH3HtLBlI1+mcM
midIFmZgYECQD3lwkRjkp0Vq6GgwQeGXkrl5om3AUT9BemGVY+HjGijcvft0szEy
i8NO3fxmt1VMUtXSPqLVqF1fhq2+KAhHt859hEukW+hcFuuEKrQff5cNc2/rzhOP
cDuMeD+tn8Y6f2ezFqJnKIE2Ei2Cdz+UOgngOuk7t5hXsQKdrOXO4tm7ulM6xGce
W2bWD+SvFgYtxcjIkzqZKULR6SUqCGETVABidChUqG8BvtQNIwp9jyzWaxNRkacV
I1+2WGb69BF2RZXN2vm6HkV6sg78ZneYr8T/Hlshlwi8uYTJZFVC6U/+rLBO9gp4
YVEnM1HSB6cYSimMfhL/oA3jDCgkpnImWI9NQyY8fjJT5uf9I8TZvNdVKd1kfyEP
ctgIHy3euYh+NU1tgW2gwUhfa34QQlhcyLHNH7EODthHHy/oHtvqhkyFpX6m5J9/
fUW5zPlkaPLVwWPC5KwS3rbilsSH/mmfYNldBrxN7PMqYsTnuSRclVbXIiaER0QP
qY5S6L3Xd+s8JoG6SIOKsa0/4EKXpfIHUutyavmrxFXW7+gpYn/v9emVrLsa3UAu
ouPneFsV54tpxiwirEmXDvwJBLD30xic903j7QQ3pR/WumBTMS/yp/Sf3SL68Ss1
boi49fSUXXoL6MLq6QW9Px8K1cgcID5q4U2YTLRp94TBI1IiCIZjX7DLjCfM3WCQ
nuSfOb+oKbxY6Tw/dZoy7Y5v5IzLghZtA4SUnvfiiitw057Ry5W80gNctXhPWyX4
be06+NdkVvaNc2kSCI0avLeCrNuBd1kJ0jdDIQBlEC7mPt9eO+fW3wxzHP/Q99+N
sjcWV0HQNFPRQzgkTqbaPVOr8rWLi1bF541w7qw7wayYns/SRoCrRu0MGCtUqKsY
EsVxrtgVHjDuiAkj+j6q6eh0dd75YFwzARr4D2JhKADkTU1V8iiZDskhbACtfz5b
bFcw5S6R0xSBhjU0Dq7/c2DzVZX+hO5e3TK9+M6+7fh8J22XKHMJKlGjkQT5Rw5g
7rDyRyaJsCVTAFxbNN7Xe353X99fYeHarv/tPh/VTm/3Uu3d8nX9oF6zMY2I0bZs
S8cv77j3ZKxguVA5NQaUW6TbsEE5rnyUL8fZpBocYu5mWbb5UAa+mpj8l+7igkjr
K2YPyUE5sSOvh5m3KZSl3OJt2dMXUBQQVDQeBLXCmobjeSpBUxpoTfCHNnktydaW
ZcLnl1auhWNC07lkwYeuOQEBYMC5xdUIFByLmxXzWCs3yRKYzigFAS8kSIF8qgYH
hd+AfegDqCxhToFHl19qEjQk224yHpJhpPBHBS2LtE1+bYjgCMp694e/2lqcQw7L
vHSpOi1I6w2FQcu1oTLPdetuOTCV2MWJOAQ00hH8/4WcV7fy4psyXfBqkMBaHD/j
LPb/w2zHSaQqVL8wWoMk/RjzlhonBs+9h23S5h1BGKKiJQ3WfJ/GZ7mBuxbLQpIN
TyZvSG24Ikki/CPbtv3sMoEG9eyrC7duEoXX/uCx1OTmmKGGWFkFuwf7z+5u5LYQ
p6+Zj1SYldoPWi1elnbd0t1/djX0gWbKslsro6r0oYHYKaM/lR1HEtM3H46ckIe8
NfSWmuOQkYS93tr8wBEVW6fuBkZZZb+UqZmVMc+ytSh8SswMtf0+b0GzCKeuF2J+
SyT9Ag6dZTmJErB8rLFeE35clrHnDU8oIfuih/ROhGwSzb9hRWG3OJm7i7VqaJen
qwR9N/RGcYy/RnnpEO53itCRG92FbSK5dQziq5PBirqUT6SOnnqjzA+WvcKu65ae
riUiURQmTrch+dYFj0ednsSMh1JkD1h9rByk6xD3f2VG9FAHjw5abcGv5ymbM8Qv
mv/VaCSvnrZCrx/jA8wdZ17XGlLpXLVgFnnwpSSFirNsyCzOneh+Y5ZZ4OR6BoMm
FIo9/K5VAQBHEQJMNbf/wKoE6Km19p+l1R3cqGOi4dc2Q3wJw6HcPZVkwR64HNKQ
alAcOtC0kpLnoAXSDgP9HHfUlHIDRgt/CKUOeDa3DIG131q5tlgee0ae74oAfFBM
G35PEpPqZS2WQM5d2SzyhgOb+yFlU5U0So5eM7jHz5QhBB2uVlqck9PBkqKYYkX4
e68lITpbkyQjNGTGUqS6OLgSD7sg3FdlfuxxwTyxPB18MaEu4nBEqU4MObUYZ273
VHzdZollupPrtPILAkIVnCfdhCzFaymymBLwtZQ8b3x/nvd8INK4sqTCrTYJEm+I
y9iK91M8wAvO44S2ZACi9n/1jwDlC8Z5XmeqOl0owoQl3mRB9h8O1pDT0Oh3jKwV
WuUHKlOHJRRLXTYPSsx140A00/UTIeEZpv4gB0+zjm2zUAtKbVbEEvkwuJTdNziJ
yahl1xWBX35w66W70bwr8PsHJndfQIBEg83uhW4ln1eG4cVQjX1ccdf+VSne/Qob
ckzi4KSA8chVk+hAtQ7p72383ISBjAPsTVp7IPNLNo36In151Gx5GCR2vERo+DBJ
eY6e+lvwb7xUUhyQvhjdanbkn9Q/WqrzNLJsW6rlPocreL+wFUdux7ly8YdJ/4k0
9o2xBN9vlkcDUroEZeAl1HvQmDBnJPMtSltb6E8lOoONydlLqZe3c/hKddSj1v0t
MUMyeYygcCAYpkdFjHrOznam4kXaJx9TH8i0LdENWhmp7VcB7h3L5JjVaYxwH1QJ
jIrkuQVNfC/o3iOaJsUVH5lXV2COR+GX+KLHp76aVeF/3f8e/G5xAZSkHc3BXYzF
3/cGJKjqHN0S+DRKahnS0pU+L54vBgm1VfHl8ZgnMiriAAfIFZ2U85wYojxYcYHs
iiXOuhgRe7nhhPtZvnKneQkJWyQ0XKH14+K0CGKicpIGBIpnCNhI5gql/wNLVcaN
SEJ2/lPkKVr6+UDdzDcKZpU7LgJlLl1gopEVdnezOHbVmdGc+ybnwNN1tflJQ+3Q
K9XYwYLXtrY6xQTgZu7mSvPsyHkjAdNgtm73O1ukynZtmDaV3vCDUoE3onRns4Tk
/T+sTmv0bGYb/hOyyINy6bIUiAwG7iO1wwcZf9ENvXaEID5EoQUDotdJklH0WQs7
c+ZOGXdKUearS8JylB19F9PS1D5tuKEk12K1xrFURe/yx5FnNrTfKks3l2Ajo+7P
GM7Rwc8a+5j1ReG7d+HmrkUdHwrG7NTOzbaFFgyq/0+qe5L2MAAc/zjyAxRMCZMX
U0rKxD7pR8hOWUAJa1stXKnTltyLAPI040ebOtL5JgPkdxzvuyz9YCKSqdQW5vPf
D8CkwM0VItJ21UZDsKKNY0InRp6ChWI09rW2k+OhUjdT9qXo86QNA5MLqOhuY9n0
rU1BfrOkZ1N6pAbtqK78J7oe1lMYVKiNoUwWkjWP7aIgDunpUy8EcerjBkxOGp3q
7TcSOXTKUlAP0FNeJsNFin0qgOHEtykMHpqJFGzoh7gjO3rdsE08lzZP5S17vZTq
AyFkg6sD3vJWI/Y4HN5YEtm+JpAUXrUy4syJjDbyR/qiv0FTrSm7i+534lmE7ZHo
OfRkUpF77JcvqgtYUFEsrTpNi1plnVfQr7gehNtPd3I6I/euJZxb7HyRykLBbxsP
xXfz3Ntxr2ljE7E1gbevYslOiPruM6i7MLXI7OTZrzBMJjxF79trAwr7aosL5a1C
plhDtLE6azwmusuWqfddYyAwCKMmZT0ux9iVAzG05gBx+E1xwiFZMJXeVHN+LVgX
afRWq0/VFpgwMkVwHWobXCeiJ7EQxeFFc3yZjStGNBZhc4PrgezilPR6IBYrP5TF
6e/2VA2n3KFDcKl/p3bdw7RpunDGfg5ImTPu6kbbdSFxpbxMuxTjt8ozA6zxB2cZ
4IhLUNGMmbmbLDcnNOxDN3gp8Y+yODYSqVSAwJH5bMAqFvVILObp7P2MuaohXza1
KLYiVrRIqBdXnn7ir9R+H5vFCD2S5JBs6uIZMZJmHtu/7aMNWPjn2/Wupxdkkglw
78lpmv3wTvE+FwdqIOzAqtByHM0zIU3MSnX7gjBnp3uQn86XGzXnZo9Iux7PfJB7
2VaELEEJy8lC3SCePV5HaCUOLlQTWbpTtplP92SIXuVw0mE6s6/Pfh4LvV8m/6lm
dM23n+jnLuk8B3OALyDxun7tIC4/ClkhSgn9qmoFfBbtR7R8mqY/1/K2rhR/bVl8
qn3uLk55uZk/Fj5ztT7WS26XvlakC2Jcf/l1r3C/scKivIKmP1pw4uhuCMvGxphg
PIfkhwMONoFawCIo5Y+Cn2oFg3IMKPijg2QWTyWd4MoZsYFtwQ9Kd22s4D38jTWt
MwQSFi4VnDEOoCKF7Giuw2UigKz9262aPKvbHpzqNCCv1QmjpDvEusxoYEluGt7h
tacjV0k7cQc9cs+rtVbmahx4BZOa11bzMkgJW6KgbTrQ1u418RaHmfC3neLqZup6
LHfZkjfAad2ZG1f+UgkersgbiNOHrFaUhZERN0U+gn2ke2W8z348eX3hEzg4VrfR
A0XNssa9aIOpWRcAok7RmbE84D782cTXDfHTEmJGT+V2Ys8X4wWomzrORAFTuLYQ
M8r/0nTazbZ7tdzezTSgq8STXzizuI47wMJCDqHj1x1sudkrn3P9Uo2fw3HpQsEb
jDRoQzItGAQZ58Qbg0sJEyWyveWrL1yUY5OVwa8vlr6ZSBYZ8LinZlQFqe3wQOix
0bJgT3nMW5Lq3IxKmWqYmtaZVZXjFeOladMZD1A5B4NkfYbc3PgRxvwoAxoPalZs
Maz6DrvIcygchy+AWFHHSlQfDyK5ck7l49GEPNtKXy6LkyZnDSEZcXkr1q3zoeY3
n2yJXCs6nPSjTHxv77iR0MpoeBmlzB9clfcIJGQqku18RpsldboUVwqs8F20V2AY
H+pBP3b6oE36iBec73vXcwd6HfHpBoRqhD80L9yRL/XeDu0PuwW2oq06tmkU6NEB
Ga/jgwH4FDLmwe+lSggWKdddIEE8mNiPb84p/73L3vyWByjy7UesNwP5LuISHFmy
oYY+bwFuCKSXje7W4j1lzfLm2VTYtvMNdrxsE68vMOzzyElVg8vK2erYKBB09XO0
ZEkfHWN3WtSNc93l/RCnZpUFRaL5GiT4ayY10Z4RZl62BqjA19hdRxTXkgQy/DCf
uOURabzab8wevLTyASJz1YsQxFniHOAP8jEjcGdBQCz/e3BzFxLKcJ6K/gNZrxg2
Awfpdo809Pz5nJemGOwCHiZkb0BoszqCX8BxEdUcycnqI5uqRMjSO3Mriuin4ejM
ACT0xvTLpfxErNYoyqNPRO3VAHxCbG/8lCCUbKAoPYcZSNNRosDCCjPn+rp9WfgQ
gTof93CsiBwKF3UzJeegU30wWpOTnxoC57mZwRIREbQKYwVtSMFVJM2DSjLMqrBz
0f4EQwA49VsavDhl60NS4uxNfMCbt2IUkW5mRh3vpZle0qrS6BYlJQy/5GL8Q6nT
ecSmXT3+5bPX1bFT/7wfQAjXLxkX45JdmhTmy0N7kDRvCkUNCSsvieo9AlzoYmIN
isOQ5YgkvJL1+vgZsN31zoBuE/uWUq9e7ap+Sj25r1v87UQ2wi3PdAslJ3VJD6xA
LGufA6+zng65LjxUzT20y/pjzf5zCPOkGaOGQELf2d9GXhpXxBFj6wrzrPsnnLYK
8JGKcfypQwiX5lNHaNI1G9FX2UOFN8e9BdEa/oYpjB4wGPmaQad3bjuf9Wpo5rr8
edlrSP9tjHi/y5Qvei1mmqx1ke39W0U0xpxRdy4yNxTfTvW8YGSLtmL7uCExyukm
r3VRkT0+2eh/kv9/vySDThltlAYqbh9fjJonBu+c8W19fPftfnOxtvymeXpQrddi
Cj20vDT5JxA3OO8mhW/qZl0Lm+ku0D5YcZoPHz0B8yrBvCuCuTzVSog9gaPyCYHg
ZGo+w0+wKp/3hsULdwu6ki2CbyYUsRfC/5QSqTf8mqK9mvx0XYuCFITmyWkHz8ZR
MKuODNJMkLVrtoIYzEa56C4dP1iLhfEvGiA4XfIEsH1bbvGR9GhMFRvGybKsT75Q
XYMk8E2QNvNewe2lhJIf6MjKd/OyMVJc6G+j4oxWd9LaFzeiFGunX+ZuP50brm/G
zrEWR6lrcQnWEHIqJ+zLjQq9HZEG1KleXmTLZ4xAHrS4KmC9eVg3srAkwzsbaDiN
HAx1nNVi6IdSxOsPxH9t4nCqr+rNb/Pmih8go/Yi5DCIwbfHFNF3VwLEF14poVpx
HiRlFhWZaooeJyZ8VTTTgfEbfQAE4I/DwiM/c0fjA1W1B3v4OdIe4D7VSf3WgF1n
T1HclYQNH6TfEot2/uS1/AutuZCbU9EPk11HwoADHiOcHKd1KEKZ9VO/7KaIpun6
oAYHW4xrYx50xI0BAw1HsySvs/+LLFwyH/jB3iN+bHhNOc4utuVgeq+5I5OJFJXJ
/iZ0aYsMlWM/95eiwB5VH9xm0MVenjdKE1spU7S4Zp3aKwb+RhZcv6HlQV27D2Jt
mZp59b6bv5QvRuqqN58H4vj9gKnrU4HGsSa03bsufYgV4GfwaIqhtoOdKbZLhavU
UJvrc2pPei+ZO0zapb4oMQSOq6mMPlXygeh3nFmo5uKkLpl3T/Zwy4eoptUaLDW3
eMKOnv2OfqKgiIXiJO6P8fFObyvFJVxshBiG6iTOa1wzk54ltsKpVkuYy+1tAUkm
EiVYa6Ga/jCG2yZJaCnIkNblYod/d8f/DajrhJ8a1M/tTWvfi8BYAsm+UIkGgzaf
S3iG8BJvaV4pcD8XWm6lnD2Namku6+6zC6LSI2fD1/ynOJUxgcMnis06DaOH2baT
2HXlLk6MEhjyReYKWLhpQarWdSF0sLteqGI5UEM/QvsFCPCAJc9h7xVTqiN9uIEs
Vbu+hQY4+aUS4GUKw8xpNJzGbtKx+DxH/ATvG29sclpCT4Nj6PbeZQ/8mNLhMTXz
qlFaZ2oWBD+2ntikqsCH1f+QcLg7Vqm65xcV7tFcwQ74983Bs8+O2suB1dtVo4Yb
YsyZ3RC6LvUxeu7yGWFgXqcMrINbPKPO0ay8wyMytk+xW6rlkgV23UYdgmgJvgEG
ABtBJm5ufb5IijeELPIMqhhfKAYtRkfuwigoehFCIzzhON5WJBWAfOt4C8rGpGPz
jYHKNm8b/j4EMR4RyTFjrDODVTvx9G4hzxagtbTQziMLtOqLHKFj3bYlxsN65rVH
xepKQmAt32Dwwj+8NzSd3dy8peGq6NW+7mDmmeDVZHlja2xTQt5Z7bYCDjci90kz
ot6wBc17opu2M/QB5EBo2upm5T8R4zNTT33ZVu6iqab1ydAg3EIdxESWh640z/fI
0dfdsx6AEkLWXCrZj37ZaePxAs90YUoCPg02nF+mWH7o5iBx28NZjaZLSXGC0sgA
cLIxtGpaJXQwvUCpGXsx7MNgy0BmUG0iVHZ+e1IL5Ak/YCSRgQPxXXOBw0hXHUAi
FkH5mfI9ySJ+tyupF5D9UVfyyun1mOTBgGtWT6Uy1N5bgTcEwTGFs3uw/cjUPRkU
nA3nMIsMzpdbFLaR4CorDAmy1KZLci0XJWR9ZI/uArj0ZXVCyMEE6r5XZe+PaN7N
uxLrj4wThoNh503rn+q8+wxpxdqV8ZYYvqMJtpeupGD1P+e84jWtpOayGxJHIFzg
R5d8S8DnPSSLXFzEPwixF/LX7zlMolpcOLoJB+lfnnTdRqmvQ/IZdQdtxVRxr4/e
BayYQWncOv9zDgysPc9IX1fsBHPoMhJTF1RqweYDWBgxe5cSJrli/XRRnyDkUaF8
D+OkVBb3Pal9PSe/3KWba3vt6dAL3mhon7IM+6iHPu0Xml/oBBxqMQP6gLhTWFzG
YgT6ut3mdfEKgxeFAiAxS+b1V+gsom4h4zdCKBoPtmjrz+OTUyvKP6d480OCDAAZ
hwNpksjxPhBvgZxox8N+e8hZpAZO3X41QPsXxpbo1/nVjb4opQIjsQ7V8OXqHMwY
C+3H7DhQHzQon+PcArjT1FJibqBUKmJPSjpa+646H2txX1D1qe1Vt1uLSf0z2tGI
ZhzWNLSmS05DVYgCsgmSdsWLArDu8M7K7U1EMppB4U1P8uwxTfIQsDKiAnENvnwc
nI8UtVAZrWDwo+8bGnBcc2y9HMDUtb+7FNRouHZ4P2+hjReNQpB2bGanCpK+lvkN
1TUVJM/VeySSDry68y7/tepyCwv7/EMZJTK7iI2t6BDDNYHKaspPfyb7Q9H8XbmT
`pragma protect end_protected
