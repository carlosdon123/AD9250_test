
module core_pll (
	locked,
	outclk_0,
	outclk_1,
	refclk,
	rst,
	outclk_2);	

	output		locked;
	output		outclk_0;
	output		outclk_1;
	input		refclk;
	input		rst;
	output		outclk_2;
endmodule
