// jesd204b.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module jesd204b (
		input  wire        alldev_lane_aligned,        //       alldev_lane_aligned.export
		output wire [4:0]  csr_cf,                     //                    csr_cf.export
		output wire [1:0]  csr_cs,                     //                    csr_cs.export
		output wire [7:0]  csr_f,                      //                     csr_f.export
		output wire        csr_hd,                     //                    csr_hd.export
		output wire [4:0]  csr_k,                      //                     csr_k.export
		output wire [4:0]  csr_l,                      //                     csr_l.export
		output wire [1:0]  csr_lane_powerdown,         //        csr_lane_powerdown.export
		output wire [7:0]  csr_m,                      //                     csr_m.export
		output wire [4:0]  csr_n,                      //                     csr_n.export
		output wire [4:0]  csr_np,                     //                    csr_np.export
		output wire [3:0]  csr_rx_testmode,            //           csr_rx_testmode.export
		output wire [4:0]  csr_s,                      //                     csr_s.export
		output wire        dev_lane_aligned,           //          dev_lane_aligned.export
		output wire        dev_sync_n,                 //                dev_sync_n.export
		input  wire        jesd204_rx_avs_chipselect,  //            jesd204_rx_avs.chipselect
		input  wire [7:0]  jesd204_rx_avs_address,     //                          .address
		input  wire        jesd204_rx_avs_read,        //                          .read
		output wire [31:0] jesd204_rx_avs_readdata,    //                          .readdata
		output wire        jesd204_rx_avs_waitrequest, //                          .waitrequest
		input  wire        jesd204_rx_avs_write,       //                          .write
		input  wire [31:0] jesd204_rx_avs_writedata,   //                          .writedata
		input  wire        jesd204_rx_avs_clk,         //        jesd204_rx_avs_clk.clk
		input  wire        jesd204_rx_avs_rst_n,       //      jesd204_rx_avs_rst_n.reset_n
		input  wire [63:0] jesd204_rx_dlb_data,        //       jesd204_rx_dlb_data.export
		input  wire [1:0]  jesd204_rx_dlb_data_valid,  // jesd204_rx_dlb_data_valid.export
		input  wire [7:0]  jesd204_rx_dlb_disperr,     //    jesd204_rx_dlb_disperr.export
		input  wire [7:0]  jesd204_rx_dlb_errdetect,   //  jesd204_rx_dlb_errdetect.export
		input  wire [7:0]  jesd204_rx_dlb_kchar_data,  // jesd204_rx_dlb_kchar_data.export
		input  wire        jesd204_rx_frame_error,     //    jesd204_rx_frame_error.export
		output wire        jesd204_rx_int,             //            jesd204_rx_int.irq
		output wire [63:0] jesd204_rx_link_data,       //           jesd204_rx_link.data
		output wire        jesd204_rx_link_valid,      //                          .valid
		input  wire        jesd204_rx_link_ready,      //                          .ready
		input  wire        pll_ref_clk,                //               pll_ref_clk.clk
		input  wire [1:0]  rx_analogreset,             //            rx_analogreset.rx_analogreset
		output wire [1:0]  rx_cal_busy,                //               rx_cal_busy.rx_cal_busy
		input  wire [1:0]  rx_digitalreset,            //           rx_digitalreset.rx_digitalreset
		output wire [1:0]  rx_islockedtodata,          //         rx_islockedtodata.rx_is_lockedtodata
		input  wire [1:0]  rx_serial_data,             //            rx_serial_data.rx_serial_data
		input  wire        rxlink_clk,                 //                rxlink_clk.clk
		input  wire        rxlink_rst_n_reset_n,       //              rxlink_rst_n.reset_n
		output wire [1:0]  rxphy_clk,                  //                 rxphy_clk.export
		output wire [3:0]  sof,                        //                       sof.export
		output wire [3:0]  somf,                       //                      somf.export
		input  wire        sysref                      //                    sysref.export
	);

	jesd204b_altera_jesd204_161_zta4dmq #(
		.DEVICE_FAMILY            ("Arria 10"),
		.SUBCLASSV                (1),
		.PCS_CONFIG               ("JESD_PCS_CFG1"),
		.L                        (2),
		.M                        (2),
		.F                        (2),
		.N                        (14),
		.N_PRIME                  (16),
		.S                        (1),
		.K                        (16),
		.SCR                      (1),
		.CS                       (0),
		.CF                       (0),
		.HD                       (0),
		.ECC_EN                   (0),
		.DLB_TEST                 (0),
		.PHADJ                    (0),
		.ADJCNT                   (0),
		.ADJDIR                   (0),
		.OPTIMIZE                 (0),
		.DID                      (0),
		.BID                      (0),
		.LID0                     (0),
		.FCHK0                    (0),
		.LID1                     (1),
		.FCHK1                    (0),
		.LID2                     (2),
		.FCHK2                    (0),
		.LID3                     (3),
		.FCHK3                    (0),
		.LID4                     (4),
		.FCHK4                    (0),
		.LID5                     (5),
		.FCHK5                    (0),
		.LID6                     (6),
		.FCHK6                    (0),
		.LID7                     (7),
		.FCHK7                    (0),
		.JESDV                    (1),
		.PMA_WIDTH                (32),
		.SER_SIZE                 (4),
		.FK                       (32),
		.RES1                     (0),
		.RES2                     (0),
		.BIT_REVERSAL             (0),
		.BYTE_REVERSAL            (0),
		.ALIGNMENT_PATTERN        (658812),
		.PULSE_WIDTH              (2),
		.LS_FIFO_DEPTH            (32),
		.LS_FIFO_WIDTHU           (5),
		.UNUSED_TX_PARALLEL_WIDTH (92),
		.UNUSED_RX_PARALLEL_WIDTH (72),
		.XCVR_PLL_LOCKED_WIDTH    (2),
		.RECONFIG_ADDRESS_WIDTH   (11)
	) jesd204_0 (
		.pll_ref_clk                (pll_ref_clk),                //               pll_ref_clk.clk
		.rxlink_clk                 (rxlink_clk),                 //                rxlink_clk.clk
		.rxlink_rst_n_reset_n       (rxlink_rst_n_reset_n),       //              rxlink_rst_n.reset_n
		.jesd204_rx_avs_clk         (jesd204_rx_avs_clk),         //        jesd204_rx_avs_clk.clk
		.jesd204_rx_avs_rst_n       (jesd204_rx_avs_rst_n),       //      jesd204_rx_avs_rst_n.reset_n
		.jesd204_rx_avs_chipselect  (jesd204_rx_avs_chipselect),  //            jesd204_rx_avs.chipselect
		.jesd204_rx_avs_address     (jesd204_rx_avs_address),     //                          .address
		.jesd204_rx_avs_read        (jesd204_rx_avs_read),        //                          .read
		.jesd204_rx_avs_readdata    (jesd204_rx_avs_readdata),    //                          .readdata
		.jesd204_rx_avs_waitrequest (jesd204_rx_avs_waitrequest), //                          .waitrequest
		.jesd204_rx_avs_write       (jesd204_rx_avs_write),       //                          .write
		.jesd204_rx_avs_writedata   (jesd204_rx_avs_writedata),   //                          .writedata
		.jesd204_rx_link_data       (jesd204_rx_link_data),       //           jesd204_rx_link.data
		.jesd204_rx_link_valid      (jesd204_rx_link_valid),      //                          .valid
		.jesd204_rx_link_ready      (jesd204_rx_link_ready),      //                          .ready
		.jesd204_rx_dlb_data        (jesd204_rx_dlb_data),        //       jesd204_rx_dlb_data.export
		.jesd204_rx_dlb_data_valid  (jesd204_rx_dlb_data_valid),  // jesd204_rx_dlb_data_valid.export
		.jesd204_rx_dlb_kchar_data  (jesd204_rx_dlb_kchar_data),  // jesd204_rx_dlb_kchar_data.export
		.jesd204_rx_dlb_errdetect   (jesd204_rx_dlb_errdetect),   //  jesd204_rx_dlb_errdetect.export
		.jesd204_rx_dlb_disperr     (jesd204_rx_dlb_disperr),     //    jesd204_rx_dlb_disperr.export
		.alldev_lane_aligned        (alldev_lane_aligned),        //       alldev_lane_aligned.export
		.sysref                     (sysref),                     //                    sysref.export
		.jesd204_rx_frame_error     (jesd204_rx_frame_error),     //    jesd204_rx_frame_error.export
		.jesd204_rx_int             (jesd204_rx_int),             //            jesd204_rx_int.irq
		.csr_rx_testmode            (csr_rx_testmode),            //           csr_rx_testmode.export
		.dev_lane_aligned           (dev_lane_aligned),           //          dev_lane_aligned.export
		.dev_sync_n                 (dev_sync_n),                 //                dev_sync_n.export
		.sof                        (sof),                        //                       sof.export
		.somf                       (somf),                       //                      somf.export
		.csr_f                      (csr_f),                      //                     csr_f.export
		.csr_k                      (csr_k),                      //                     csr_k.export
		.csr_l                      (csr_l),                      //                     csr_l.export
		.csr_m                      (csr_m),                      //                     csr_m.export
		.csr_n                      (csr_n),                      //                     csr_n.export
		.csr_s                      (csr_s),                      //                     csr_s.export
		.csr_cf                     (csr_cf),                     //                    csr_cf.export
		.csr_cs                     (csr_cs),                     //                    csr_cs.export
		.csr_hd                     (csr_hd),                     //                    csr_hd.export
		.csr_np                     (csr_np),                     //                    csr_np.export
		.csr_lane_powerdown         (csr_lane_powerdown),         //        csr_lane_powerdown.export
		.rxphy_clk                  (rxphy_clk),                  //                 rxphy_clk.export
		.rx_serial_data             (rx_serial_data),             //            rx_serial_data.rx_serial_data
		.rx_analogreset             (rx_analogreset),             //            rx_analogreset.rx_analogreset
		.rx_digitalreset            (rx_digitalreset),            //           rx_digitalreset.rx_digitalreset
		.rx_islockedtodata          (rx_islockedtodata),          //         rx_islockedtodata.rx_is_lockedtodata
		.rx_cal_busy                (rx_cal_busy)                 //               rx_cal_busy.rx_cal_busy
	);

endmodule
